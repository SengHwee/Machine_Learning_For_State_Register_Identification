
module aes_core(\bus_in[0] , \bus_in[1] , \bus_in[2] , \bus_in[3] , \bus_in[4] , \bus_in[5] , \bus_in[6] , \bus_in[7] , \bus_in[8] , \bus_in[9] , \bus_in[10] , \bus_in[11] , \bus_in[12] , \bus_in[13] , \bus_in[14] , \bus_in[15] , \bus_in[16] , \bus_in[17] , \bus_in[18] , \bus_in[19] , \bus_in[20] , \bus_in[21] , \bus_in[22] , \bus_in[23] , \bus_in[24] , \bus_in[25] , \bus_in[26] , \bus_in[27] , \bus_in[28] , \bus_in[29] , \bus_in[30] , \bus_in[31] , \iv_en[0] , \iv_en[1] , \iv_en[2] , \iv_en[3] , \iv_sel_rd[0] , \iv_sel_rd[1] , \iv_sel_rd[2] , \iv_sel_rd[3] , \key_en[0] , \key_en[1] , \key_en[2] , \key_en[3] , \key_sel_rd[0] , \key_sel_rd[1] , \data_type[0] , \data_type[1] , \addr[0] , \addr[1] , \op_mode[0] , \op_mode[1] , \aes_mode[0] , \aes_mode[1] , start, disable_core, write_en, read_en, first_block, rst_n, clk, \col_out[0] , \col_out[1] , \col_out[2] , \col_out[3] , \col_out[4] , \col_out[5] , \col_out[6] , \col_out[7] , \col_out[8] , \col_out[9] , \col_out[10] , \col_out[11] , \col_out[12] , \col_out[13] , \col_out[14] , \col_out[15] , \col_out[16] , \col_out[17] , \col_out[18] , \col_out[19] , \col_out[20] , \col_out[21] , \col_out[22] , \col_out[23] , \col_out[24] , \col_out[25] , \col_out[26] , \col_out[27] , \col_out[28] , \col_out[29] , \col_out[30] , \col_out[31] , \key_out[0] , \key_out[1] , \key_out[2] , \key_out[3] , \key_out[4] , \key_out[5] , \key_out[6] , \key_out[7] , \key_out[8] , \key_out[9] , \key_out[10] , \key_out[11] , \key_out[12] , \key_out[13] , \key_out[14] , \key_out[15] , \key_out[16] , \key_out[17] , \key_out[18] , \key_out[19] , \key_out[20] , \key_out[21] , \key_out[22] , \key_out[23] , \key_out[24] , \key_out[25] , \key_out[26] , \key_out[27] , \key_out[28] , \key_out[29] , \key_out[30] , \key_out[31] , \iv_out[0] , \iv_out[1] , \iv_out[2] , \iv_out[3] , \iv_out[4] , \iv_out[5] , \iv_out[6] , \iv_out[7] , \iv_out[8] , \iv_out[9] , \iv_out[10] , \iv_out[11] , \iv_out[12] , \iv_out[13] , \iv_out[14] , \iv_out[15] , \iv_out[16] , \iv_out[17] , \iv_out[18] , \iv_out[19] , \iv_out[20] , \iv_out[21] , \iv_out[22] , \iv_out[23] , \iv_out[24] , \iv_out[25] , \iv_out[26] , \iv_out[27] , \iv_out[28] , \iv_out[29] , \iv_out[30] , \iv_out[31] , end_aes);
  wire AES_CORE_CONTROL_UNIT__abc_10818_n109;
  wire AES_CORE_CONTROL_UNIT__abc_10818_n112;
  wire AES_CORE_CONTROL_UNIT__abc_10818_n118;
  wire AES_CORE_CONTROL_UNIT__abc_10818_n12;
  wire AES_CORE_CONTROL_UNIT__abc_10818_n122;
  wire AES_CORE_CONTROL_UNIT__abc_10818_n24;
  wire AES_CORE_CONTROL_UNIT__abc_10818_n29;
  wire AES_CORE_CONTROL_UNIT__abc_10818_n303;
  wire AES_CORE_CONTROL_UNIT__abc_10818_n306;
  wire AES_CORE_CONTROL_UNIT__abc_10818_n307;
  wire AES_CORE_CONTROL_UNIT__abc_10818_n310;
  wire AES_CORE_CONTROL_UNIT__abc_10818_n4;
  wire AES_CORE_CONTROL_UNIT__abc_10818_n41;
  wire AES_CORE_CONTROL_UNIT__abc_10818_n59;
  wire AES_CORE_CONTROL_UNIT__abc_10818_n79;
  wire AES_CORE_CONTROL_UNIT__abc_10818_n97;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n100;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n101_1;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n103;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n104;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n105;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n106_1;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n107;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n108;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n109_1;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n110_1;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n111;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n112;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n113;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n114_1;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n115;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n117_1;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n118;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n119;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n121;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n122;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n123;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n124_1;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n125;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n127;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n128;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n130_1;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n131;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n132;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n134;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n135;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n137;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n138;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n140;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n141_1;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n142;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n143;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n144;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n145;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n148;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n149;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n151;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n152;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n154;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n155_1;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n156;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n158;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n159;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n160;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n163;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n164;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n165;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n166;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n168;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n169;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n170;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n171_1;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n173;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n174;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n175_1;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n176;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n178;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n179_1;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n180;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n181_1;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n183_1;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n184_1;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n185;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n186;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n188;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n189_1;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n190;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n193;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n195;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n196;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n197_1;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n198;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n199;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n200_1;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n201;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n203_1;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n204;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n206_1;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n207_1;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n209_1;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n210_1;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n211_1;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n212_1;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n213;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n214;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n215;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n216;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n217;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n218;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n219;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n220;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n221;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n222;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n223;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n225;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n226;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n227;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n228;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n229;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n230;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n231;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n232;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n236;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n238;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n239;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n241;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n242;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n244;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n245;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n247;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n248;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n249;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n73;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n75;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n76_1;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n77;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n78;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n79_1;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n81_1;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n82_1;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n84_1;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n85;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n86_1;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n87_1;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n88;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n89_1;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n90;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n91;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n92;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n93_1;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n94;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n95;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n96_1;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n97;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n98;
  wire AES_CORE_CONTROL_UNIT__abc_15841_n99_1;
  wire AES_CORE_CONTROL_UNIT_bypass_key_en;
  wire AES_CORE_CONTROL_UNIT_bypass_rk;
  wire AES_CORE_CONTROL_UNIT_bypass_rk_bF_buf0;
  wire AES_CORE_CONTROL_UNIT_bypass_rk_bF_buf1;
  wire AES_CORE_CONTROL_UNIT_bypass_rk_bF_buf2;
  wire AES_CORE_CONTROL_UNIT_bypass_rk_bF_buf3;
  wire AES_CORE_CONTROL_UNIT_col_en_0_;
  wire AES_CORE_CONTROL_UNIT_col_en_1_;
  wire AES_CORE_CONTROL_UNIT_col_en_2_;
  wire AES_CORE_CONTROL_UNIT_col_en_3_;
  wire AES_CORE_CONTROL_UNIT_col_sel_0_;
  wire AES_CORE_CONTROL_UNIT_col_sel_1_;
  wire AES_CORE_CONTROL_UNIT_encrypt_decrypt;
  wire AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf0;
  wire AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf1;
  wire AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf10;
  wire AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf11;
  wire AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf12;
  wire AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf13;
  wire AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf14;
  wire AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf2;
  wire AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf3;
  wire AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf4;
  wire AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf5;
  wire AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf6;
  wire AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf7;
  wire AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf8;
  wire AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf9;
  wire AES_CORE_CONTROL_UNIT_iv_cnt_en;
  wire AES_CORE_CONTROL_UNIT_key_derivation_en;
  wire AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf0;
  wire AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf1;
  wire AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf10;
  wire AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf2;
  wire AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf3;
  wire AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf4;
  wire AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf5;
  wire AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf6;
  wire AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf7;
  wire AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf8;
  wire AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf9;
  wire AES_CORE_CONTROL_UNIT_key_en_0_;
  wire AES_CORE_CONTROL_UNIT_key_en_1_;
  wire AES_CORE_CONTROL_UNIT_key_en_2_;
  wire AES_CORE_CONTROL_UNIT_key_en_3_;
  wire AES_CORE_CONTROL_UNIT_key_gen;
  wire AES_CORE_CONTROL_UNIT_key_out_sel_0_;
  wire AES_CORE_CONTROL_UNIT_key_out_sel_1_;
  wire AES_CORE_CONTROL_UNIT_key_sel;
  wire AES_CORE_CONTROL_UNIT_last_round;
  wire AES_CORE_CONTROL_UNIT_last_round_bF_buf0;
  wire AES_CORE_CONTROL_UNIT_last_round_bF_buf1;
  wire AES_CORE_CONTROL_UNIT_last_round_bF_buf2;
  wire AES_CORE_CONTROL_UNIT_last_round_bF_buf3;
  wire AES_CORE_CONTROL_UNIT_last_round_bF_buf4;
  wire AES_CORE_CONTROL_UNIT_last_round_bF_buf5;
  wire AES_CORE_CONTROL_UNIT_mode_cbc;
  wire AES_CORE_CONTROL_UNIT_mode_cbc_bF_buf0;
  wire AES_CORE_CONTROL_UNIT_mode_cbc_bF_buf1;
  wire AES_CORE_CONTROL_UNIT_mode_cbc_bF_buf2;
  wire AES_CORE_CONTROL_UNIT_mode_cbc_bF_buf3;
  wire AES_CORE_CONTROL_UNIT_mode_cbc_bF_buf4;
  wire AES_CORE_CONTROL_UNIT_mode_ctr;
  wire AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf0;
  wire AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf1;
  wire AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf2;
  wire AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf3;
  wire AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf4;
  wire AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf5;
  wire AES_CORE_CONTROL_UNIT_rd_count_0_;
  wire AES_CORE_CONTROL_UNIT_rd_count_0__FF_INPUT;
  wire AES_CORE_CONTROL_UNIT_rd_count_1_;
  wire AES_CORE_CONTROL_UNIT_rd_count_1__FF_INPUT;
  wire AES_CORE_CONTROL_UNIT_rd_count_2_;
  wire AES_CORE_CONTROL_UNIT_rd_count_2__FF_INPUT;
  wire AES_CORE_CONTROL_UNIT_rd_count_3_;
  wire AES_CORE_CONTROL_UNIT_rd_count_3__FF_INPUT;
  wire AES_CORE_CONTROL_UNIT_rk_sel_0_;
  wire AES_CORE_CONTROL_UNIT_rk_sel_1_;
  wire AES_CORE_CONTROL_UNIT_sbox_sel_0_;
  wire AES_CORE_CONTROL_UNIT_sbox_sel_1_;
  wire AES_CORE_CONTROL_UNIT_sbox_sel_2_;
  wire AES_CORE_CONTROL_UNIT_state_0_;
  wire AES_CORE_CONTROL_UNIT_state_11_;
  wire AES_CORE_CONTROL_UNIT_state_12_;
  wire AES_CORE_CONTROL_UNIT_state_13_;
  wire AES_CORE_CONTROL_UNIT_state_14_;
  wire AES_CORE_CONTROL_UNIT_state_15_;
  wire AES_CORE_CONTROL_UNIT_state_1_;
  wire AES_CORE_CONTROL_UNIT_state_2_;
  wire AES_CORE_CONTROL_UNIT_state_3_;
  wire AES_CORE_CONTROL_UNIT_state_4_;
  wire AES_CORE_CONTROL_UNIT_state_6_;
  wire AES_CORE_CONTROL_UNIT_state_7_;
  wire AES_CORE_CONTROL_UNIT_state_8_;
  wire AES_CORE_CONTROL_UNIT_state_9_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1000;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1001;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1003;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1004;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1006;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1007;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1008;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1010;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1011;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1013;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1014;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1015;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1017;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1018;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1020;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1021;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1022;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1024;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1025;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1027;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1028;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1029;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1031;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1032;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1034;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1035;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1036;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1038;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1039;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1041;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1042;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1043;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1045;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1046;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1048;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1049;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1050;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1052;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1053;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1054;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1056;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1057;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1058;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1060;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1061;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1062;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1064;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1065;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1066;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1068;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1069;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1070;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1072;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1073;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1074;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1076;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1077;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1078;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1080;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1081;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1082;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1084;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1085;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1086;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1088;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1089;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1090;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1092;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1093;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1094;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1096;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1097;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1098;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1100;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1101;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1102;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1104;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1105;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1106;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1108;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1109;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1110;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1112;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1113;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1114;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1116;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1117;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1118;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1120;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1121;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1122;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1124;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1125;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1126;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1128;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1129;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1130;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1132;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1133;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1134;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1136;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1137;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1138;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1140;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1141;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1142;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1144;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1145;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1146;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1147;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1149;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1150;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1151;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1153;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1154;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1155;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1157;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1158;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1159;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1160;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1162;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1163;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1164;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1166;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1167;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1168;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1170;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1171;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1172;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1174;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1175;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1176;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1178;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1179;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1180;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1182;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1183;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1184;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1186;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1187;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1188;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1190;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1191;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1192;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1194;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1195;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1196;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1198;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1199;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1200;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1202;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1203;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1204;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1206;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1207;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1208;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1210;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1211;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1212;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1214;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1215;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1216;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1218;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1219;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1220;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1222;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1223;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1224;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1226;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1227;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1228;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1230;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1231;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1232;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1234;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1235;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1236;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1238;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1239;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1240;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1242;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1243;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1244;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1246;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1247;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1248;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1250;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1251;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1252;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1254;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1255;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1256;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1258;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1259;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1260;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1262;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1263;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1264;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1266;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1267;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1268;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1270;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1271;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1272;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1274;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1275;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1276;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1278;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1279;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1280;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1282;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1283;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1284;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1286;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1287;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1288;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1290;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1291;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1292;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1294;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1295;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1296;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1298;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1299;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1300;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1302;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1303;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1304;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n327_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n328_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n329_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n330_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n331_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n332_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n333_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n334_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n335_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n336_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n338_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n339_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n340_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n341_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n342_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n343_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n344_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n345_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n346_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n347_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n349_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n350_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n351_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n352_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n353_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n354_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n355_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n356_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n357_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n358_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n360_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n361_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n362_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n363_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n364_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n365_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n366_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n367_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n368_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n369_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n371_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n372_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n373_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n374_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n375_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n376_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n377_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n378_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n379_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n380_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n382_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n383_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n384_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n385_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n386_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n387_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n388_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n389_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n390_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n391_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n393_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n394_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n395_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n396_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n397_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n398_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n399_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n400_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n401_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n402_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n404_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n405_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n406_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n407_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n408_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n409_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n410_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n411_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n412_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n413_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n415_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n416_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n417_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n418_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n419_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n420_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n421_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n422_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n423_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n424_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n426_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n427_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n428_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n429_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n430_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n431_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n432_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n433_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n434_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n435_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n437_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n438_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n439_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n440_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n441_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n442_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n443_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n444_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n445_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n446_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n448_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n449_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n450_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n451_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n452_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n453_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n454_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n455_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n456_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n457_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n459_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n460_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n461_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n462_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n463_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n464_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n465_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n466_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n467_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n468_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n470_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n471_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n472_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n473_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n474_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n475_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n476_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n477_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n478_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n479_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n481_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n482_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n483_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n484_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n485_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n486_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n487_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n488_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n489_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n490_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n492_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n493_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n494_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n495_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n496_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n497_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n498_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n499_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n500_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n501_1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n503;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n504;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n505;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n506;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n507;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n508;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n509;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n510;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n511;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n512;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n514;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n515;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n516;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n517;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n518;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n519;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n520;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n521;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n522;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n523;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n525;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n526;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n527;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n528;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n529;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n530;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n531;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n532;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n533;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n534;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n536;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n537;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n538;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n539;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n540;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n541;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n542;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n543;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n544;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n545;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n547;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n548;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n549;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n550;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n551;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n552;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n553;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n554;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n555;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n556;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n558;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n559;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n560;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n561;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n562;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n563;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n564;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n565;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n566;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n567;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n569;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n570;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n571;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n572;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n573;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n574;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n575;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n576;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n577;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n578;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n580;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n581;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n582;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n583;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n584;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n585;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n586;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n587;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n588;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n589;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n591;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n592;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n593;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n594;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n595;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n596;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597_bF_buf0;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597_bF_buf1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597_bF_buf2;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597_bF_buf3;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597_bF_buf4;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n598;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n599;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n600;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n601;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n602;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n603;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n604;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n605;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n606;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n607;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n608;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n609;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n610;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n611;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n612;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n613;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n614;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n615;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n617;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n618;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n619;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n620;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n621;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n622;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n623;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n624;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n625;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n626;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n627;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n628;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n629;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n630;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n631;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n632;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n633;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n634;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n635;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n636;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n637;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n638;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n639;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n640;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n641;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n642;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n643;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n644;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n645;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n646;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n647;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n648;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n650;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n651;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n652;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n653;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n654;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n655;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n656;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n657;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n658;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n659;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n660;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n661;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n662;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n663;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n664;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n665;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n666;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n667;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n668;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n669;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n670;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n671;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n672;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n673;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n674;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n675;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n676;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n677;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n678;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n679;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n680;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n681;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n682;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n683;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n684;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n685;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n686;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n687;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n688;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n690;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n691;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n692;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n693;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n694;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n695;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n696;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n697;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n698;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n699;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n700;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n701;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n702;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n703;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n704;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n705;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n706;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n707;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n708;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n709;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n711;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n712;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n713;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n714;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n715;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n716;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n717;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n718;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n719;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n720;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n721;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n722;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n723;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n724;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n725;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n726;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n727;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n728;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n729;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n730;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n731;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n732;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n733;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n734;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n735;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n736;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n737;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n738;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n740;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n741;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n742;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n743;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n744;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n745;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n746;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n747;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n748;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n749;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n750;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n751;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n752;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n753;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n754;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n755;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n756;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n757;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n758;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n759;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n760;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n761;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n762;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n763;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n764;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n765;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n766;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n768;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n769;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n770;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n771;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n772;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n773;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n774;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n775;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n776;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n777;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n778;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n779;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n780;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n781;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n782;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n783;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n784;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n785;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n786;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n787;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n788;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n789;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n790;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n791;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n792;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n793;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n794;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n795;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n796;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n797;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n798;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n800;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n801;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n802;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n803;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n804;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n805;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n806;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n807;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n808;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n809;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n810;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n811;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n812;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n813;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n814;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n815;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n816;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n817;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n818;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n819;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n820;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n821;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n822;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n824;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n825;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n826;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n828;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n829;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n831;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n832;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n833;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n835;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n836;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n838;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n839;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n840;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n842;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n843;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n845;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n846;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n847;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n849;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n850;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n852;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n853;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n854;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n856;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n857;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n859;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n860;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n861;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n863;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n864;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n866;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n867;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n868;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n870;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n871;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n873;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n874;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n875;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n877;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n878;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n880;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n881;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n882;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n884;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n885;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n887;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n888;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n889;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n891;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n892;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n894;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n895;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n896;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n898;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n899;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n901;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n902;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n903;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n905;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n906;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n908;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n909;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n910;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n912;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n913;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n915;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n916;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n917;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n919;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n920;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n922;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n923;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n924;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n926;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n927;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n929;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n930;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n931;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n933;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n934;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n936;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n937;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n938;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n940;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n941;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n943;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n944;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n945;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n947;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n948;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n950;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n951;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n952;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n954;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n955;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n957;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n958;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n959;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n961;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n962;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n964;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n965;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n966;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n968;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n969;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n971;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n972;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n973;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n975;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n976;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n978;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n979;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n980;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n982;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n983;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n985;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n986;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n987;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n989;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n990;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n992;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n993;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n994;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n996;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n997;
  wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n999;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out_bF_buf0;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out_bF_buf1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out_bF_buf2;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out_bF_buf3;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out_bF_buf4;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf0;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf1;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf2;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf3;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf4;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf5;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf6;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf7;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_0_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_10_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_11_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_12_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_13_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_14_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_15_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_16_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_17_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_18_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_19_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_1_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_20_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_21_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_22_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_23_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_2_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_3_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_4_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_5_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_6_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_7_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_8_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_9_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_0_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_10_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_11_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_12_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_13_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_14_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_15_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_16_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_17_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_18_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_19_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_1_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_20_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_21_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_22_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_23_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_24_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_25_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_26_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_27_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_28_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_29_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_2_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_30_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_31_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_3_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_4_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_5_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_6_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_7_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_8_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_9_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_out_24_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_out_25_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_out_26_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_out_27_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_out_28_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_out_29_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_out_30_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_g_out_31_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__0_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__10_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__11_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__12_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__13_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__14_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__15_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__16_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__17_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__18_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__19_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__1_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__20_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__21_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__22_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__23_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__24_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__25_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__26_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__27_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__28_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__29_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__2_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__30_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__31_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__3_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__4_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__5_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__6_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__7_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__8_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__9_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__0_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__10_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__11_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__12_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__13_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__14_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__15_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__16_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__17_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__18_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__19_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__1_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__20_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__21_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__22_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__23_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__24_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__25_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__26_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__27_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__28_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__29_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__2_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__30_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__31_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__3_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__4_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__5_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__6_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__7_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__8_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__9_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__0_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__10_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__11_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__12_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__13_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__14_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__15_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__16_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__17_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__18_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__19_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__1_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__20_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__21_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__22_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__23_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__24_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__25_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__26_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__27_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__28_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__29_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__2_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__30_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__31_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__3_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__4_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__5_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__6_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__7_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__8_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__9_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__0_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__10_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__11_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__12_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__13_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__14_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__15_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__16_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__17_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__18_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__19_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__1_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__20_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__21_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__22_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__23_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__24_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__25_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__26_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__27_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__28_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__29_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__2_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__30_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__31_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__3_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__4_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__5_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__6_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__7_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__8_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__9_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_0_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_100_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_101_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_102_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_103_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_104_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_105_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_106_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_107_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_108_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_109_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_10_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_110_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_111_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_112_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_113_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_114_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_115_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_116_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_117_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_118_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_119_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_11_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_120_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_121_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_122_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_123_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_124_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_125_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_126_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_127_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_12_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_13_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_14_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_15_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_16_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_17_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_18_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_19_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_1_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_20_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_21_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_22_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_23_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_24_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_25_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_26_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_27_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_28_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_29_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_2_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_30_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_31_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_32_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_33_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_34_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_35_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_36_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_37_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_38_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_39_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_3_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_40_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_41_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_42_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_43_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_44_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_45_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_46_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_47_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_48_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_49_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_4_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_50_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_51_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_52_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_53_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_54_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_55_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_56_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_57_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_58_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_59_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_5_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_60_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_61_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_62_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_63_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_64_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_65_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_66_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_67_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_68_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_69_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_6_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_70_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_71_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_72_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_73_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_74_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_75_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_76_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_77_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_78_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_79_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_7_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_80_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_81_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_82_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_83_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_84_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_85_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_86_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_87_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_88_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_89_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_8_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_90_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_91_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_92_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_93_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_94_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_95_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_96_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_97_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_98_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_99_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_9_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_round_0_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_round_1_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_round_2_;
  wire AES_CORE_DATAPATH_KEY_EXPANDER_round_3_;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n100;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n101;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n102;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n103;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n104;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n105_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n106;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n107;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n108;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n109_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n110;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n111;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n112;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n113;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n114;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n115_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n116;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n117;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n119_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n120;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n121;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n122;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n123_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n124;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n125;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n126;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n127_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n128;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n129_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n130;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n131;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n132;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n133;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n134_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n135;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n136_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n137;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n138;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n139;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n140_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n141;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n142_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n143;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n144;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n145;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n146;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n147_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n148;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n149_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n150;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n151;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n152;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n153;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n154_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n155;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n156_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n157;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n159;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n160_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n161;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n162_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n163;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n164;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n165;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n166_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n167;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n168_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n169;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n170;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n171;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n172_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n173;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n174_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n175;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n176_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n177_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n178;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n179;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n180_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n181_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n182;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n183_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n185;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n186;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n187_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n188_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n189;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n190;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n191_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n192_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n193;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n194_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n195_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n196;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n197_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n198_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n199;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n200_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n201_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n202;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n203_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n204_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n205;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n206;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n207_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n208_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n209;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n210_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n211_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n212;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n213;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n214_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n215_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n216;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n217;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n218_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n219_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n221_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n222_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n223;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n224_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n225_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n226;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n227_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n228_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n229;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n230;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n231;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n232;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n233;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n234;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n235;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n236;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n237;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n239;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n240;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n241;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n242;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n243;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n244;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n245;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n246;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n247;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n248;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n249;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n250;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n251;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n252;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n253;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n254;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n255;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n256;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n257;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n258;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n259;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n260;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n261;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n262;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n263;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n264;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n265;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n266;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n267;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n268;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n269;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n270;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n271;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n272;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n273;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n274;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n276;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n277;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n278;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n279;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n280;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n281;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n282;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n283;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n284;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n285;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n286;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n287;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n288;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n289;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n290;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n291;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n292;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n293;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n294;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n295;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n296;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n297;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n298;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n300;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n301;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n302;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n303;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n304;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n305;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n306;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n307;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n308;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n309;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n310;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n311;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n312;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n313;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n314;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n315;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n316;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n317;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n318;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n319;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n320;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n321;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n322;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n323;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n324;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n325;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n326;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n327;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n328;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n329;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n330;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n331;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n332;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n333;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n334;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n335;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n336;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n337;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n339;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n340;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n341;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n342;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n343;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n344;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n345;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n346;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n347;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n348;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n349;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n350;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n351;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n352;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n353;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n354;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n355;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n356;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n357;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n358;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n359;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n360;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n361;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n363;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n364;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n365;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n366;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n367;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n368;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n369;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n370;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n371;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n372;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n373;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n374;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n375;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n376;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n377;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n378;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n379;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n380;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n381;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n382;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n383;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n384;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n385;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n386;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n387;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n388;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n389;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n390;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n391;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n392;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n393;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n394;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n395;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n396;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n397;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n398;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n399;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n401;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n402;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n403;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n404;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n405;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n406;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n407;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n408;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n409;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n410;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n411;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n412;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n414;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n415;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n416;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n417;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n418;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n419;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n420;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n421;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n422;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n423;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n424;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n425;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n426;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n427;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n428;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n429;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n430;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n431;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n432;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n433;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n434;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n435;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n436;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n437;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n438;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n439;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n440;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n441;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n442;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n444;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n445;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n446;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n447;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n448;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n449;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n450;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n451;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n452;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n453;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n454;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n455;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n456;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n457;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n459;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n460;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n461;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n462;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n463;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n464;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n465;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n466;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n467;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n468;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n469;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n470;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n471;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n472;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n473;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n474;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n475;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n476;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n477;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n479;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n480;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n481;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n482;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n483;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n484;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n485;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n486;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n487;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n488;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n490;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n491;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n492;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n493;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n494;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n495;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n496;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n497;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n498;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n499;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n500;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n502;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n503;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n504;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n505;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n506;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n507;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n508;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n509;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n510;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n511;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n513;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n514;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n515;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n516;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n517;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n518;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n519;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n521;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n522;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n523;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n524;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n525;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n526;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n527;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n528;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n529;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n530;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n531;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n532;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n533;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n534;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n535;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n537;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n538;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n539;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n540;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n541;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n542;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n544;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n545;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n546;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n547;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n548;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n549;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n550;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n551;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n552;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n553;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n555;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n556;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n557;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n558;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n559;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n560;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n561;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n563;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n564;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n565;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n566;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n567;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n568;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n569;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n570;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n571;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n572;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n573;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n574;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n575;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n576;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n578;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n579;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n580;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n581;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n582;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n583;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n584;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n585;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n586;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n588;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n589;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n590;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n591;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n592;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n593;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n594;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n595;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n596;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n597;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n598;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n599;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n600;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n601;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n603;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n604;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n605;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n606;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n607;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n608;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n609;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n610;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n611;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n613;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n614;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n615;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n616;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n617;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n618;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n619;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n620;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n621;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n622;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n624;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n625;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n626;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n627;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n628;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n629;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n630;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n631;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n632;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n634;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n635;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n636;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n637;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n638;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n639;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n640;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n641;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n642;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n643;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n644;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n646;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n647;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n648;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n649;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n650;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n651;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n653;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n654;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n655;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n656;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n657;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n658;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n659;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n660;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n661;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n662;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n663;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n664;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n665;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n666;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n667;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n669;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n670;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n671;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n672;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n673;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n674;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n676;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n677;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n678;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n679;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n680;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n681;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n682;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n683;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n684;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n685;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n687;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n688;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n689;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n691;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n692;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n693;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n694;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n695;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n696;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n697;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n698;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n699;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n700;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n701;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n702;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n703;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n704;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n705;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n707;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n708;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n710;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n711;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n712;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n713;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n714;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n715;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n716;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n717;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n718;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n719;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n721;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n722;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n723;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n725;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n726;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n727;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n728;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n729;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n730;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n731;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n732;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n733;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n734;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n735;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n736;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n737;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n739;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n740;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n741;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n743;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n744;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n745;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n746;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n747;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n748;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n749;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n750;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n751;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n752;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n753;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n754;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n755;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n756;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n757;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n759;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n760;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n762;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n763;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n764;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n765;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n766;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n767;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n768;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n769;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n770;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n771;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n772;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n774;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n775;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n777;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n778;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n779;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n780;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n781;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n782;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n783;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n784;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n785;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n786;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n788;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n789;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n790;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n792;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n793;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n794;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n795;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n796;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n797;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n798;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n799;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n800;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n801;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n802;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n804;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n805;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n807;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n808;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n809;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n810;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n811;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n812;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n814;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n815;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n816;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n818;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n819;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n820;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n821;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n822;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n823;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n824;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n825;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n826;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n827;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n828;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n829;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n830;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n831;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n832;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n834;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n835;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n837;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n838;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n839;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n840;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n841;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n842;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n843;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n844;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n845;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n846;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n847;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n849;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n850;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n852;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n853;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n854;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n855;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n856;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n857;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n858;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n859;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n860;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n861;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n862;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n863;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n864;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n865;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n867;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n868;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n869;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n871;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n872;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n873;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n874;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n875;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n876;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n877;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n878;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n879;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n880;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n881;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n882;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n883;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n884;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n885;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n887;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n888;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n890;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n891;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n892;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n893;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n894;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n895;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n896;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n897;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n898;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n899;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n900;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n902;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n903;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n905;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n906;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n907;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n908;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n909;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n910;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n911;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n912;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n913;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n914;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n916;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n917;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n918;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n920;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n921;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n922;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n923;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n924;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n925;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n926;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n928;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n929;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n97_1;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n98;
  wire AES_CORE_DATAPATH_MIX_COL__abc_25501_n99;
  wire AES_CORE_DATAPATH_MIX_COL_col_0__0_;
  wire AES_CORE_DATAPATH_MIX_COL_col_0__1_;
  wire AES_CORE_DATAPATH_MIX_COL_col_0__2_;
  wire AES_CORE_DATAPATH_MIX_COL_col_0__3_;
  wire AES_CORE_DATAPATH_MIX_COL_col_0__4_;
  wire AES_CORE_DATAPATH_MIX_COL_col_0__5_;
  wire AES_CORE_DATAPATH_MIX_COL_col_0__6_;
  wire AES_CORE_DATAPATH_MIX_COL_col_0__7_;
  wire AES_CORE_DATAPATH_MIX_COL_col_1__0_;
  wire AES_CORE_DATAPATH_MIX_COL_col_1__1_;
  wire AES_CORE_DATAPATH_MIX_COL_col_1__2_;
  wire AES_CORE_DATAPATH_MIX_COL_col_1__3_;
  wire AES_CORE_DATAPATH_MIX_COL_col_1__4_;
  wire AES_CORE_DATAPATH_MIX_COL_col_1__5_;
  wire AES_CORE_DATAPATH_MIX_COL_col_1__6_;
  wire AES_CORE_DATAPATH_MIX_COL_col_1__7_;
  wire AES_CORE_DATAPATH_MIX_COL_col_2__0_;
  wire AES_CORE_DATAPATH_MIX_COL_col_2__1_;
  wire AES_CORE_DATAPATH_MIX_COL_col_2__2_;
  wire AES_CORE_DATAPATH_MIX_COL_col_2__3_;
  wire AES_CORE_DATAPATH_MIX_COL_col_2__4_;
  wire AES_CORE_DATAPATH_MIX_COL_col_2__5_;
  wire AES_CORE_DATAPATH_MIX_COL_col_2__6_;
  wire AES_CORE_DATAPATH_MIX_COL_col_2__7_;
  wire AES_CORE_DATAPATH_MIX_COL_col_3__0_;
  wire AES_CORE_DATAPATH_MIX_COL_col_3__1_;
  wire AES_CORE_DATAPATH_MIX_COL_col_3__2_;
  wire AES_CORE_DATAPATH_MIX_COL_col_3__3_;
  wire AES_CORE_DATAPATH_MIX_COL_col_3__4_;
  wire AES_CORE_DATAPATH_MIX_COL_col_3__5_;
  wire AES_CORE_DATAPATH_MIX_COL_col_3__6_;
  wire AES_CORE_DATAPATH_MIX_COL_col_3__7_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_0_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_10_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_11_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_12_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_13_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_14_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_15_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_16_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_17_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_18_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_19_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_1_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_20_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_21_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_22_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_23_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_24_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_25_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_26_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_27_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_28_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_29_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_2_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_30_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_31_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_3_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_4_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_5_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_6_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_7_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_8_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_9_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_0_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_10_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_11_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_12_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_13_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_14_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_15_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_16_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_17_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_18_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_19_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_1_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_20_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_21_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_22_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_23_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_24_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_25_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_26_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_27_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_28_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_29_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_2_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_30_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_31_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_3_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_4_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_5_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_6_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_7_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_8_;
  wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_9_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n100;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n101_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n102;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n103;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n104_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n105;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n106;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n107;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n108;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n109;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n110;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n111;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n112;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n113;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n114;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n116;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n117;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n118;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n119;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n120;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n121_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n122;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n123;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n124;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n125;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n126_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n128;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n129;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n130;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n131;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n132;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n133;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n134;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n135;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n136;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n138;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n139_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n140;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n142;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n143_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n144;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n145_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n146_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n147;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n148_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n149;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n150_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n151_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n152_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n153_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n154;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n156;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n157;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n158;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n159;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n160;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n161;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n162;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n163;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n164;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n165;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n166_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n167;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n168;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n169;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n170;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n171;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n172;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n173;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n174;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n175;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n176_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n177;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n178;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n179;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n180;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n181;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n182_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n183;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n184;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n185;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n186;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n187_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n188_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n189_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n190_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n191;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n192;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n193;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n194;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n195;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n196;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n197;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n198;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n199;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n200;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n201;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n202;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n203;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n204;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n205;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n206;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n207;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n208;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n209;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n210;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n211;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n212;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n213;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n214;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n215;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n216;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n217;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n218;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n219;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n220;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n221;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n222;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n223;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n224;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n225;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n226;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n227;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n228;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n229;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n230;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n231;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n232;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n233;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n234;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n235;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n236;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n237;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n238;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n239;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n240;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n241;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n242;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n243;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n244;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n245;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n246;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n247;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n248;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n249;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n250;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n251;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n252;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n253;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n254;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n255;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n256;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n257;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n258;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n259;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n260;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n261;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n262;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n263;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n264;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n265;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n266;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n267;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n268;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n269;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n270;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n271;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n272;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n273;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n274;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n275;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n276;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n277;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n278;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n279;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n280;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n281;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n282;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n283;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n284;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n285;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n286;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n287;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n288;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n289;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n290;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n291;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n292;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n293;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n294;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n295;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n296;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n297;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n298;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n299;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n300;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n301;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n302;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n303;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n304;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n305;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n306;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n307;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n308;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n309;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n310;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n311;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n312;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n313;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n314;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n315;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n316;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n317;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n318;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n319;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n321;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n322;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n323;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n324;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n325;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n326;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n327;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n328;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n329;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n330;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n331;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n332;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n333;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n334;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n335;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n336;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n337;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n338;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n339;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n340;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n342;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n343;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n344;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n345;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n346;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n347;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n348;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n349;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n350;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n351;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n352;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n353;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n354;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n355;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n356;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n358;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n359;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n360;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n361;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n362;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n363;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n364;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n365;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n366;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n367;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n368;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n369;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n370;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n371;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n372;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n373;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n374;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n375;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n376;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n377;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n378;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n379;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n380;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n381;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n382;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n383;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n384;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n385;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n386;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n387;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n388;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n389;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n390;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n391;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n392;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n393;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n394;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n395;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n396;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n397;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n398;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n399;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n401;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n402;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n403;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n404;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n405;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n406;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n407;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n408;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n409;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n410;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n412;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n413;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n414;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n415;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n416;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n417;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n418;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n419;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n420;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n421;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n422;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n423;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n424;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n425;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n426;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n427;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n429;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n430;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n431;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n432;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n433;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n434;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n435;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n436;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n437;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n439;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n441;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n442;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n443;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n444;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n445;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n447;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n448;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n449;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n450;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n451;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n452;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n453;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n454;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n456;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n457;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n459;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n460;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n461;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n463;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n464;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n466;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n467;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n468;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n469;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n470;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n471;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n472;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n473;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n474;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n475;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n476;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n477;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n478;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n479;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n480;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n481;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n482;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n483;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n484;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n485;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n486;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n487;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n488;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n489;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n490;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n491;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n492;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n493;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n494;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n495;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n496;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n497;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n498;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n499;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n50;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n500;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n501;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n502;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n503;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n504;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n505;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n506;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n507;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n508;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n510;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n511;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n512;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n513;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n514;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n515;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n516;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n517;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n518;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n519;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n51_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n52;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n520;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n521;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n522;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n523;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n524;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n525;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n526;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n527;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n528;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n529;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n530;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n531;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n532;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n533;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n534;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n535;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n536;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n537;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n538;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n539;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n53_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n540;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n541;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n542;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n543;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n544;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n545;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n546;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n548;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n549;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n54_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n55;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n550;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n551;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n552;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n553;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n554;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n555;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n556;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n557;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n558;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n559;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n56;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n560;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n561;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n562;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n563;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n564;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n565;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n567;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n568;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n569;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n57;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n570;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n571;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n572;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n573;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n574;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n575;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n576;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n577;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n578;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n579;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n58;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n580;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n582;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n583;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n584;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n586;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n587;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n589;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n59;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n590;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n60;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n61;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n62;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n63;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n64;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n65;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n66_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n67;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n68;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n69;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n70;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n71_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n72;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n73;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n74;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n75;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n76;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n78;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n79;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n80;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n81;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n82;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n83;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n84_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n85;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n86_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n87;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n89;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n90;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n91;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n92;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n93;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n94_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n95;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n96;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n97_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n98;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_0_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_1_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_2_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_3_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_4_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_5_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_6_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_7_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_0_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_1_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_2_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_3_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_4_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_5_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_6_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_7_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_1_2_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_stage1_0_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_stage1_1_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_stage1_2_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_stage1_3_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_0_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_1_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_2_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_3_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_0_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_1_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_2_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_3_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_4_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_5_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_6_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_7_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_1_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_2_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_3_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_4_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_5_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_6_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_7_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n100;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n101_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n102;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n103;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n104_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n105;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n106;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n107;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n108;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n109;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n110;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n111;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n112;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n113;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n114;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n116;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n117;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n118;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n119;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n120;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n121_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n122;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n123;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n124;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n125;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n126_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n128;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n129;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n130;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n131;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n132;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n133;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n134;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n135;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n136;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n138;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n139_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n140;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n142;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n143_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n144;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n145_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n146_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n147;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n148_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n149;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n150_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n151_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n152_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n153_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n154;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n156;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n157;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n158;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n159;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n160;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n161;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n162;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n163;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n164;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n165;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n166_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n167;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n168;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n169;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n170;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n171;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n172;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n173;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n174;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n175;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n176_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n177;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n178;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n179;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n180;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n181;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n182_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n183;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n184;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n185;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n186;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n187_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n188_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n189_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n190_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n191;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n192;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n193;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n194;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n195;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n196;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n197;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n198;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n199;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n200;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n201;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n202;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n203;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n204;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n205;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n206;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n207;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n208;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n209;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n210;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n211;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n212;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n213;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n214;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n215;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n216;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n217;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n218;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n219;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n220;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n221;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n222;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n223;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n224;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n225;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n226;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n227;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n228;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n229;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n230;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n231;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n232;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n233;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n234;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n235;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n236;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n237;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n238;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n239;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n240;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n241;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n242;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n243;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n244;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n245;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n246;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n247;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n248;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n249;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n250;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n251;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n252;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n253;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n254;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n255;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n256;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n257;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n258;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n259;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n260;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n261;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n262;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n263;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n264;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n265;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n266;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n267;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n268;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n269;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n270;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n271;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n272;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n273;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n274;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n275;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n276;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n277;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n278;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n279;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n280;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n281;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n282;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n283;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n284;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n285;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n286;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n287;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n288;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n289;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n290;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n291;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n292;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n293;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n294;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n295;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n296;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n297;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n298;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n299;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n300;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n301;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n302;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n303;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n304;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n305;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n306;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n307;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n308;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n309;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n310;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n311;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n312;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n313;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n314;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n315;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n316;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n317;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n318;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n319;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n321;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n322;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n323;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n324;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n325;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n326;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n327;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n328;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n329;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n330;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n331;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n332;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n333;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n334;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n335;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n336;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n337;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n338;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n339;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n340;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n342;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n343;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n344;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n345;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n346;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n347;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n348;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n349;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n350;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n351;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n352;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n353;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n354;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n355;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n356;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n358;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n359;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n360;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n361;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n362;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n363;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n364;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n365;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n366;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n367;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n368;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n369;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n370;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n371;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n372;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n373;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n374;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n375;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n376;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n377;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n378;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n379;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n380;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n381;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n382;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n383;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n384;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n385;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n386;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n387;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n388;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n389;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n390;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n391;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n392;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n393;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n394;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n395;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n396;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n397;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n398;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n399;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n401;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n402;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n403;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n404;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n405;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n406;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n407;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n408;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n409;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n410;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n412;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n413;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n414;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n415;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n416;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n417;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n418;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n419;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n420;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n421;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n422;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n423;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n424;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n425;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n426;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n427;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n429;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n430;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n431;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n432;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n433;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n434;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n435;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n436;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n437;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n439;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n441;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n442;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n443;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n444;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n445;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n447;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n448;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n449;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n450;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n451;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n452;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n453;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n454;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n456;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n457;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n459;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n460;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n461;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n463;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n464;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n466;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n467;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n468;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n469;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n470;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n471;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n472;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n473;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n474;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n475;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n476;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n477;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n478;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n479;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n480;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n481;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n482;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n483;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n484;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n485;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n486;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n487;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n488;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n489;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n490;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n491;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n492;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n493;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n494;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n495;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n496;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n497;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n498;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n499;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n50;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n500;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n501;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n502;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n503;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n504;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n505;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n506;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n507;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n508;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n510;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n511;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n512;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n513;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n514;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n515;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n516;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n517;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n518;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n519;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n51_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n52;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n520;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n521;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n522;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n523;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n524;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n525;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n526;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n527;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n528;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n529;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n530;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n531;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n532;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n533;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n534;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n535;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n536;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n537;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n538;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n539;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n53_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n540;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n541;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n542;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n543;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n544;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n545;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n546;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n548;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n549;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n54_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n55;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n550;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n551;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n552;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n553;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n554;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n555;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n556;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n557;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n558;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n559;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n56;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n560;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n561;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n562;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n563;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n564;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n565;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n567;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n568;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n569;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n57;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n570;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n571;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n572;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n573;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n574;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n575;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n576;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n577;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n578;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n579;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n58;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n580;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n582;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n583;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n584;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n586;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n587;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n589;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n59;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n590;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n60;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n61;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n62;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n63;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n64;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n65;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n66_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n67;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n68;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n69;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n70;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n71_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n72;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n73;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n74;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n75;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n76;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n78;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n79;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n80;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n81;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n82;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n83;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n84_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n85;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n86_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n87;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n89;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n90;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n91;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n92;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n93;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n94_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n95;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n96;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n97_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n98;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_0_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_1_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_2_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_3_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_4_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_5_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_6_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_7_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_0_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_1_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_2_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_3_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_4_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_5_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_6_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_7_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_1_2_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_stage1_0_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_stage1_1_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_stage1_2_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_stage1_3_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_0_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_1_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_2_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_3_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_0_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_1_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_2_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_3_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_4_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_5_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_6_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_7_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_1_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_2_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_3_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_4_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_5_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_6_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_7_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n100;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n101_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n102;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n103;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n104_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n105;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n106;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n107;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n108;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n109;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n110;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n111;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n112;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n113;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n114;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n116;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n117;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n118;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n119;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n120;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n121_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n122;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n123;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n124;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n125;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n126_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n128;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n129;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n130;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n131;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n132;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n133;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n134;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n135;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n136;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n138;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n139_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n140;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n142;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n143_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n144;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n145_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n146_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n147;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n148_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n149;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n150_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n151_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n152_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n153_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n154;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n156;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n157;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n158;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n159;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n160;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n161;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n162;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n163;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n164;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n165;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n166_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n167;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n168;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n169;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n170;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n171;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n172;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n173;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n174;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n175;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n176_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n177;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n178;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n179;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n180;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n181;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n182_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n183;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n184;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n185;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n186;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n187_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n188_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n189_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n190_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n191;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n192;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n193;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n194;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n195;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n196;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n197;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n198;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n199;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n200;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n201;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n202;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n203;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n204;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n205;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n206;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n207;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n208;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n209;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n210;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n211;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n212;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n213;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n214;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n215;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n216;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n217;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n218;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n219;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n220;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n221;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n222;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n223;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n224;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n225;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n226;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n227;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n228;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n229;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n230;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n231;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n232;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n233;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n234;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n235;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n236;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n237;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n238;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n239;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n240;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n241;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n242;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n243;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n244;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n245;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n246;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n247;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n248;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n249;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n250;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n251;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n252;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n253;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n254;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n255;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n256;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n257;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n258;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n259;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n260;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n261;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n262;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n263;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n264;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n265;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n266;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n267;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n268;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n269;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n270;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n271;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n272;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n273;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n274;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n275;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n276;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n277;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n278;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n279;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n280;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n281;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n282;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n283;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n284;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n285;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n286;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n287;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n288;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n289;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n290;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n291;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n292;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n293;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n294;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n295;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n296;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n297;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n298;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n299;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n300;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n301;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n302;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n303;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n304;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n305;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n306;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n307;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n308;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n309;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n310;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n311;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n312;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n313;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n314;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n315;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n316;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n317;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n318;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n319;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n321;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n322;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n323;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n324;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n325;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n326;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n327;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n328;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n329;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n330;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n331;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n332;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n333;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n334;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n335;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n336;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n337;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n338;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n339;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n340;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n342;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n343;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n344;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n345;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n346;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n347;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n348;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n349;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n350;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n351;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n352;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n353;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n354;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n355;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n356;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n358;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n359;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n360;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n361;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n362;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n363;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n364;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n365;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n366;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n367;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n368;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n369;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n370;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n371;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n372;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n373;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n374;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n375;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n376;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n377;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n378;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n379;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n380;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n381;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n382;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n383;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n384;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n385;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n386;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n387;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n388;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n389;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n390;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n391;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n392;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n393;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n394;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n395;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n396;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n397;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n398;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n399;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n401;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n402;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n403;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n404;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n405;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n406;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n407;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n408;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n409;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n410;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n412;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n413;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n414;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n415;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n416;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n417;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n418;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n419;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n420;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n421;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n422;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n423;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n424;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n425;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n426;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n427;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n429;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n430;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n431;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n432;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n433;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n434;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n435;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n436;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n437;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n439;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n441;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n442;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n443;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n444;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n445;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n447;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n448;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n449;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n450;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n451;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n452;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n453;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n454;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n456;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n457;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n459;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n460;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n461;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n463;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n464;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n466;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n467;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n468;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n469;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n470;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n471;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n472;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n473;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n474;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n475;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n476;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n477;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n478;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n479;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n480;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n481;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n482;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n483;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n484;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n485;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n486;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n487;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n488;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n489;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n490;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n491;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n492;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n493;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n494;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n495;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n496;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n497;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n498;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n499;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n50;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n500;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n501;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n502;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n503;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n504;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n505;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n506;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n507;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n508;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n510;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n511;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n512;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n513;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n514;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n515;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n516;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n517;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n518;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n519;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n51_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n52;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n520;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n521;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n522;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n523;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n524;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n525;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n526;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n527;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n528;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n529;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n530;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n531;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n532;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n533;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n534;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n535;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n536;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n537;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n538;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n539;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n53_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n540;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n541;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n542;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n543;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n544;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n545;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n546;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n548;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n549;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n54_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n55;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n550;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n551;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n552;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n553;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n554;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n555;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n556;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n557;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n558;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n559;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n56;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n560;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n561;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n562;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n563;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n564;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n565;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n567;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n568;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n569;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n57;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n570;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n571;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n572;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n573;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n574;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n575;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n576;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n577;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n578;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n579;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n58;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n580;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n582;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n583;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n584;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n586;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n587;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n589;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n59;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n590;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n60;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n61;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n62;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n63;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n64;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n65;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n66_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n67;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n68;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n69;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n70;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n71_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n72;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n73;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n74;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n75;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n76;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n78;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n79;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n80;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n81;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n82;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n83;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n84_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n85;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n86_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n87;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n89;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n90;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n91;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n92;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n93;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n94_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n95;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n96;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n97_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n98;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_0_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_1_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_2_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_3_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_4_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_5_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_6_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_7_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_0_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_1_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_2_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_3_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_4_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_5_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_6_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_7_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_1_2_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_stage1_0_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_stage1_1_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_stage1_2_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_stage1_3_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_0_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_1_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_2_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_3_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_0_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_1_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_2_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_3_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_4_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_5_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_6_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_7_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_1_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_2_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_3_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_4_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_5_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_6_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_7_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n100;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n101_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n102;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n103;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n104_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n105;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n106;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n107;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n108;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n109;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n110;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n111;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n112;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n113;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n114;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n116;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n117;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n118;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n119;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n120;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n121_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n122;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n123;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n124;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n125;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n126_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n128;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n129;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n130;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n131;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n132;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n133;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n134;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n135;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n136;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n138;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n139_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n140;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n142;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n143_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n144;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n145_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n146_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n147;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n148_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n149;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n150_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n151_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n152_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n153_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n154;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n156;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n157;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n158;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n159;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n160;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n161;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n162;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n163;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n164;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n165;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n166_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n167;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n168;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n169;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n170;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n171;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n172;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n173;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n174;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n175;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n176_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n177;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n178;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n179;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n180;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n181;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n182_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n183;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n184;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n185;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n186;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n187_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n188_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n189_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n190_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n191;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n192;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n193;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n194;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n195;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n196;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n197;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n198;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n199;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n200;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n201;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n202;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n203;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n204;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n205;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n206;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n207;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n208;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n209;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n210;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n211;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n212;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n213;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n214;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n215;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n216;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n217;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n218;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n219;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n220;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n221;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n222;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n223;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n224;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n225;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n226;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n227;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n228;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n229;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n230;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n231;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n232;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n233;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n234;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n235;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n236;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n237;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n238;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n239;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n240;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n241;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n242;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n243;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n244;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n245;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n246;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n247;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n248;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n249;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n250;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n251;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n252;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n253;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n254;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n255;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n256;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n257;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n258;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n259;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n260;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n261;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n262;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n263;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n264;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n265;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n266;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n267;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n268;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n269;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n270;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n271;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n272;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n273;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n274;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n275;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n276;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n277;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n278;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n279;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n280;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n281;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n282;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n283;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n284;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n285;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n286;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n287;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n288;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n289;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n290;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n291;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n292;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n293;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n294;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n295;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n296;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n297;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n298;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n299;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n300;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n301;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n302;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n303;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n304;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n305;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n306;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n307;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n308;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n309;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n310;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n311;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n312;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n313;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n314;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n315;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n316;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n317;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n318;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n319;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n321;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n322;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n323;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n324;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n325;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n326;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n327;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n328;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n329;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n330;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n331;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n332;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n333;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n334;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n335;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n336;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n337;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n338;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n339;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n340;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n342;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n343;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n344;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n345;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n346;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n347;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n348;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n349;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n350;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n351;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n352;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n353;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n354;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n355;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n356;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n358;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n359;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n360;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n361;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n362;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n363;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n364;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n365;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n366;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n367;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n368;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n369;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n370;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n371;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n372;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n373;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n374;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n375;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n376;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n377;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n378;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n379;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n380;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n381;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n382;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n383;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n384;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n385;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n386;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n387;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n388;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n389;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n390;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n391;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n392;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n393;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n394;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n395;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n396;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n397;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n398;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n399;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n401;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n402;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n403;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n404;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n405;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n406;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n407;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n408;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n409;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n410;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n412;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n413;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n414;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n415;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n416;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n417;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n418;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n419;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n420;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n421;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n422;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n423;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n424;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n425;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n426;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n427;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n429;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n430;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n431;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n432;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n433;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n434;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n435;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n436;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n437;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n439;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n441;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n442;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n443;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n444;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n445;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n447;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n448;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n449;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n450;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n451;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n452;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n453;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n454;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n456;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n457;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n459;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n460;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n461;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n463;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n464;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n466;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n467;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n468;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n469;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n470;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n471;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n472;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n473;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n474;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n475;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n476;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n477;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n478;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n479;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n480;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n481;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n482;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n483;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n484;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n485;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n486;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n487;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n488;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n489;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n490;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n491;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n492;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n493;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n494;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n495;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n496;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n497;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n498;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n499;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n50;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n500;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n501;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n502;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n503;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n504;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n505;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n506;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n507;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n508;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n510;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n511;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n512;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n513;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n514;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n515;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n516;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n517;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n518;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n519;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n51_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n52;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n520;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n521;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n522;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n523;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n524;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n525;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n526;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n527;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n528;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n529;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n530;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n531;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n532;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n533;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n534;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n535;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n536;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n537;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n538;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n539;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n53_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n540;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n541;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n542;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n543;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n544;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n545;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n546;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n548;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n549;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n54_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n55;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n550;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n551;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n552;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n553;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n554;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n555;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n556;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n557;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n558;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n559;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n56;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n560;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n561;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n562;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n563;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n564;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n565;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n567;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n568;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n569;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n57;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n570;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n571;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n572;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n573;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n574;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n575;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n576;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n577;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n578;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n579;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n58;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n580;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n582;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n583;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n584;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n586;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n587;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n589;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n59;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n590;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n60;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n61;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n62;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n63;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n64;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n65;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n66_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n67;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n68;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n69;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n70;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n71_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n72;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n73;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n74;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n75;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n76;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n78;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n79;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n80;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n81;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n82;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n83;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n84_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n85;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n86_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n87;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n89;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n90;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n91;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n92;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n93;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n94_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n95;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n96;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n97_1;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n98;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_0_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_1_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_2_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_3_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_4_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_5_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_6_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_7_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_0_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_1_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_2_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_3_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_4_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_5_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_6_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_7_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_1_2_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_stage1_0_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_stage1_1_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_stage1_2_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_stage1_3_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_0_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_1_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_2_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_3_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_0_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_1_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_2_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_3_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_4_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_5_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_6_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_7_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_1_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_2_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_3_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_4_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_5_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_6_;
  wire AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_7_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_0_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_100_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_101_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_102_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_103_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_104_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_105_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_106_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_107_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_108_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_109_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_10_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_110_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_111_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_112_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_113_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_114_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_115_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_116_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_117_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_118_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_119_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_11_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_120_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_121_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_122_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_123_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_124_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_125_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_126_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_127_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_12_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_13_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_14_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_15_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_16_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_17_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_18_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_19_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_1_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_20_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_21_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_22_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_23_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_24_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_25_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_26_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_27_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_28_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_29_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_2_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_30_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_31_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_32_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_33_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_34_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_35_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_36_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_37_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_38_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_39_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_3_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_40_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_41_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_42_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_43_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_44_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_45_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_46_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_47_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_48_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_49_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_4_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_50_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_51_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_52_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_53_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_54_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_55_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_56_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_57_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_58_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_59_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_5_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_60_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_61_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_62_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_63_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_64_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_65_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_66_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_67_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_68_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_69_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_6_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_70_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_71_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_72_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_73_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_74_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_75_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_76_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_77_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_78_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_79_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_7_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_80_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_81_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_82_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_83_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_84_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_85_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_86_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_87_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_88_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_89_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_8_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_90_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_91_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_92_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_93_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_94_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_95_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_96_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_97_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_98_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_99_;
  wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_9_;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n101_1;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n102_1;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n103;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n104;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n105;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n106_1;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n108;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n109;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n110_1;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n111;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n112;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n113;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n115;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n116;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n117;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n118_1;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n119;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n120;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n122_1;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n123;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n124;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n125;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n126_1;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n127;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n129;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n130_1;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n131;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n132;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n133;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n134_1;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n136;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n137;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n138_1;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n139;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n140;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n141;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n143;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n144;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n145;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n146_1;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n147;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n148;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n150_1;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n151;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n152;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n153;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n154_1;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n155;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n157;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n158_1;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n159;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n160;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n161;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n162_1;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n164;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n165;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n166_1;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n167;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n168;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n169;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n171;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n172;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n173;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n174;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n175;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n176;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n178;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n179;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n180;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n181;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n182;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n183;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n185;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n186;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n187;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n188;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n189;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n190;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n192;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n193;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n194;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n195;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n196;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n197;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n199;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n200;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n201;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n202;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n203;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n204;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n206;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n207;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n208;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n209;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n210;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n211;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n213;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n214;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n215;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n216;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n217;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n218;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n220;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n221;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n222;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n223;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n224;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n225;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n227;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n228;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n229;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n230;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n231;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n232;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n234;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n235;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n236;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n237;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n238;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n239;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n241;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n242;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n243;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n244;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n245;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n246;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n248;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n249;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n250;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n251;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n252;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n253;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n255;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n256;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n257;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n258;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n259;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n260;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n262;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n263;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n264;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n265;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n266;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n267;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n269;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n270;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n271;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n272;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n273;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n274;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n276;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n277;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n278;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n279;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n280;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n281;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n283;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n284;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n285;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n286;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n287;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n288;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n290;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n291;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n292;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n293;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n294;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n295;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1_bF_buf0;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1_bF_buf1;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1_bF_buf2;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1_bF_buf3;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1_bF_buf4;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n68;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n69;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70_bF_buf0;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70_bF_buf1;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70_bF_buf2;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70_bF_buf3;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70_bF_buf4;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n71_1;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n72_1;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n73;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74_bF_buf0;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74_bF_buf1;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74_bF_buf2;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74_bF_buf3;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74_bF_buf4;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n75;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1_bF_buf0;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1_bF_buf1;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1_bF_buf2;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1_bF_buf3;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1_bF_buf4;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n77_1;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n78;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n80;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n81_1;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n82_1;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n83;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n84;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n85;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n87_1;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n88;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n89;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n90;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n91_1;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n92_1;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n94;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n95;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n96_1;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n97_1;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n98;
  wire AES_CORE_DATAPATH_SWAP_IN__abc_16028_n99;
  wire AES_CORE_DATAPATH_SWAP_IN_data_swap_0_;
  wire AES_CORE_DATAPATH_SWAP_IN_data_swap_10_;
  wire AES_CORE_DATAPATH_SWAP_IN_data_swap_11_;
  wire AES_CORE_DATAPATH_SWAP_IN_data_swap_12_;
  wire AES_CORE_DATAPATH_SWAP_IN_data_swap_13_;
  wire AES_CORE_DATAPATH_SWAP_IN_data_swap_14_;
  wire AES_CORE_DATAPATH_SWAP_IN_data_swap_15_;
  wire AES_CORE_DATAPATH_SWAP_IN_data_swap_16_;
  wire AES_CORE_DATAPATH_SWAP_IN_data_swap_17_;
  wire AES_CORE_DATAPATH_SWAP_IN_data_swap_18_;
  wire AES_CORE_DATAPATH_SWAP_IN_data_swap_19_;
  wire AES_CORE_DATAPATH_SWAP_IN_data_swap_1_;
  wire AES_CORE_DATAPATH_SWAP_IN_data_swap_20_;
  wire AES_CORE_DATAPATH_SWAP_IN_data_swap_21_;
  wire AES_CORE_DATAPATH_SWAP_IN_data_swap_22_;
  wire AES_CORE_DATAPATH_SWAP_IN_data_swap_23_;
  wire AES_CORE_DATAPATH_SWAP_IN_data_swap_24_;
  wire AES_CORE_DATAPATH_SWAP_IN_data_swap_25_;
  wire AES_CORE_DATAPATH_SWAP_IN_data_swap_26_;
  wire AES_CORE_DATAPATH_SWAP_IN_data_swap_27_;
  wire AES_CORE_DATAPATH_SWAP_IN_data_swap_28_;
  wire AES_CORE_DATAPATH_SWAP_IN_data_swap_29_;
  wire AES_CORE_DATAPATH_SWAP_IN_data_swap_2_;
  wire AES_CORE_DATAPATH_SWAP_IN_data_swap_30_;
  wire AES_CORE_DATAPATH_SWAP_IN_data_swap_31_;
  wire AES_CORE_DATAPATH_SWAP_IN_data_swap_3_;
  wire AES_CORE_DATAPATH_SWAP_IN_data_swap_4_;
  wire AES_CORE_DATAPATH_SWAP_IN_data_swap_5_;
  wire AES_CORE_DATAPATH_SWAP_IN_data_swap_6_;
  wire AES_CORE_DATAPATH_SWAP_IN_data_swap_7_;
  wire AES_CORE_DATAPATH_SWAP_IN_data_swap_8_;
  wire AES_CORE_DATAPATH_SWAP_IN_data_swap_9_;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n101_1;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n102_1;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n103;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n104;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n105;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n106_1;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n108;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n109;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n110_1;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n111;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n112;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n113;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n115;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n116;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n117;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n118_1;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n119;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n120;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n122_1;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n123;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n124;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n125;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n126_1;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n127;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n129;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n130_1;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n131;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n132;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n133;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n134_1;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n136;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n137;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n138_1;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n139;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n140;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n141;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n143;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n144;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n145;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n146_1;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n147;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n148;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n150_1;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n151;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n152;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n153;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n154_1;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n155;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n157;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n158_1;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n159;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n160;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n161;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n162_1;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n164;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n165;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n166_1;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n167;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n168;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n169;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n171;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n172;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n173;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n174;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n175;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n176;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n178;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n179;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n180;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n181;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n182;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n183;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n185;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n186;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n187;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n188;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n189;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n190;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n192;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n193;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n194;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n195;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n196;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n197;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n199;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n200;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n201;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n202;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n203;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n204;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n206;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n207;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n208;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n209;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n210;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n211;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n213;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n214;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n215;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n216;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n217;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n218;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n220;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n221;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n222;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n223;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n224;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n225;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n227;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n228;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n229;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n230;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n231;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n232;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n234;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n235;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n236;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n237;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n238;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n239;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n241;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n242;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n243;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n244;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n245;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n246;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n248;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n249;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n250;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n251;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n252;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n253;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n255;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n256;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n257;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n258;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n259;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n260;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n262;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n263;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n264;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n265;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n266;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n267;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n269;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n270;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n271;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n272;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n273;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n274;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n276;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n277;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n278;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n279;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n280;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n281;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n283;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n284;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n285;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n286;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n287;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n288;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n290;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n291;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n292;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n293;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n294;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n295;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1_bF_buf0;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1_bF_buf1;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1_bF_buf2;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1_bF_buf3;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1_bF_buf4;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n68;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n69;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70_bF_buf0;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70_bF_buf1;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70_bF_buf2;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70_bF_buf3;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70_bF_buf4;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n71_1;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n72_1;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n73;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74_bF_buf0;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74_bF_buf1;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74_bF_buf2;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74_bF_buf3;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74_bF_buf4;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n75;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1_bF_buf0;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1_bF_buf1;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1_bF_buf2;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1_bF_buf3;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1_bF_buf4;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n77_1;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n78;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n80;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n81_1;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n82_1;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n83;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n84;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n85;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n87_1;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n88;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n89;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n90;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n91_1;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n92_1;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n94;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n95;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n96_1;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n97_1;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n98;
  wire AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n99;
  wire AES_CORE_DATAPATH__0bkp_0__31_0__0_;
  wire AES_CORE_DATAPATH__0bkp_0__31_0__10_;
  wire AES_CORE_DATAPATH__0bkp_0__31_0__11_;
  wire AES_CORE_DATAPATH__0bkp_0__31_0__12_;
  wire AES_CORE_DATAPATH__0bkp_0__31_0__13_;
  wire AES_CORE_DATAPATH__0bkp_0__31_0__14_;
  wire AES_CORE_DATAPATH__0bkp_0__31_0__15_;
  wire AES_CORE_DATAPATH__0bkp_0__31_0__16_;
  wire AES_CORE_DATAPATH__0bkp_0__31_0__17_;
  wire AES_CORE_DATAPATH__0bkp_0__31_0__18_;
  wire AES_CORE_DATAPATH__0bkp_0__31_0__19_;
  wire AES_CORE_DATAPATH__0bkp_0__31_0__1_;
  wire AES_CORE_DATAPATH__0bkp_0__31_0__20_;
  wire AES_CORE_DATAPATH__0bkp_0__31_0__21_;
  wire AES_CORE_DATAPATH__0bkp_0__31_0__22_;
  wire AES_CORE_DATAPATH__0bkp_0__31_0__23_;
  wire AES_CORE_DATAPATH__0bkp_0__31_0__24_;
  wire AES_CORE_DATAPATH__0bkp_0__31_0__25_;
  wire AES_CORE_DATAPATH__0bkp_0__31_0__26_;
  wire AES_CORE_DATAPATH__0bkp_0__31_0__27_;
  wire AES_CORE_DATAPATH__0bkp_0__31_0__28_;
  wire AES_CORE_DATAPATH__0bkp_0__31_0__29_;
  wire AES_CORE_DATAPATH__0bkp_0__31_0__2_;
  wire AES_CORE_DATAPATH__0bkp_0__31_0__30_;
  wire AES_CORE_DATAPATH__0bkp_0__31_0__31_;
  wire AES_CORE_DATAPATH__0bkp_0__31_0__3_;
  wire AES_CORE_DATAPATH__0bkp_0__31_0__4_;
  wire AES_CORE_DATAPATH__0bkp_0__31_0__5_;
  wire AES_CORE_DATAPATH__0bkp_0__31_0__6_;
  wire AES_CORE_DATAPATH__0bkp_0__31_0__7_;
  wire AES_CORE_DATAPATH__0bkp_0__31_0__8_;
  wire AES_CORE_DATAPATH__0bkp_0__31_0__9_;
  wire AES_CORE_DATAPATH__0bkp_1_0__31_0__0_;
  wire AES_CORE_DATAPATH__0bkp_1_0__31_0__10_;
  wire AES_CORE_DATAPATH__0bkp_1_0__31_0__11_;
  wire AES_CORE_DATAPATH__0bkp_1_0__31_0__12_;
  wire AES_CORE_DATAPATH__0bkp_1_0__31_0__13_;
  wire AES_CORE_DATAPATH__0bkp_1_0__31_0__14_;
  wire AES_CORE_DATAPATH__0bkp_1_0__31_0__15_;
  wire AES_CORE_DATAPATH__0bkp_1_0__31_0__16_;
  wire AES_CORE_DATAPATH__0bkp_1_0__31_0__17_;
  wire AES_CORE_DATAPATH__0bkp_1_0__31_0__18_;
  wire AES_CORE_DATAPATH__0bkp_1_0__31_0__19_;
  wire AES_CORE_DATAPATH__0bkp_1_0__31_0__1_;
  wire AES_CORE_DATAPATH__0bkp_1_0__31_0__20_;
  wire AES_CORE_DATAPATH__0bkp_1_0__31_0__21_;
  wire AES_CORE_DATAPATH__0bkp_1_0__31_0__22_;
  wire AES_CORE_DATAPATH__0bkp_1_0__31_0__23_;
  wire AES_CORE_DATAPATH__0bkp_1_0__31_0__24_;
  wire AES_CORE_DATAPATH__0bkp_1_0__31_0__25_;
  wire AES_CORE_DATAPATH__0bkp_1_0__31_0__26_;
  wire AES_CORE_DATAPATH__0bkp_1_0__31_0__27_;
  wire AES_CORE_DATAPATH__0bkp_1_0__31_0__28_;
  wire AES_CORE_DATAPATH__0bkp_1_0__31_0__29_;
  wire AES_CORE_DATAPATH__0bkp_1_0__31_0__2_;
  wire AES_CORE_DATAPATH__0bkp_1_0__31_0__30_;
  wire AES_CORE_DATAPATH__0bkp_1_0__31_0__31_;
  wire AES_CORE_DATAPATH__0bkp_1_0__31_0__3_;
  wire AES_CORE_DATAPATH__0bkp_1_0__31_0__4_;
  wire AES_CORE_DATAPATH__0bkp_1_0__31_0__5_;
  wire AES_CORE_DATAPATH__0bkp_1_0__31_0__6_;
  wire AES_CORE_DATAPATH__0bkp_1_0__31_0__7_;
  wire AES_CORE_DATAPATH__0bkp_1_0__31_0__8_;
  wire AES_CORE_DATAPATH__0bkp_1_0__31_0__9_;
  wire AES_CORE_DATAPATH__0bkp_1_1__31_0__0_;
  wire AES_CORE_DATAPATH__0bkp_1_1__31_0__10_;
  wire AES_CORE_DATAPATH__0bkp_1_1__31_0__11_;
  wire AES_CORE_DATAPATH__0bkp_1_1__31_0__12_;
  wire AES_CORE_DATAPATH__0bkp_1_1__31_0__13_;
  wire AES_CORE_DATAPATH__0bkp_1_1__31_0__14_;
  wire AES_CORE_DATAPATH__0bkp_1_1__31_0__15_;
  wire AES_CORE_DATAPATH__0bkp_1_1__31_0__16_;
  wire AES_CORE_DATAPATH__0bkp_1_1__31_0__17_;
  wire AES_CORE_DATAPATH__0bkp_1_1__31_0__18_;
  wire AES_CORE_DATAPATH__0bkp_1_1__31_0__19_;
  wire AES_CORE_DATAPATH__0bkp_1_1__31_0__1_;
  wire AES_CORE_DATAPATH__0bkp_1_1__31_0__20_;
  wire AES_CORE_DATAPATH__0bkp_1_1__31_0__21_;
  wire AES_CORE_DATAPATH__0bkp_1_1__31_0__22_;
  wire AES_CORE_DATAPATH__0bkp_1_1__31_0__23_;
  wire AES_CORE_DATAPATH__0bkp_1_1__31_0__24_;
  wire AES_CORE_DATAPATH__0bkp_1_1__31_0__25_;
  wire AES_CORE_DATAPATH__0bkp_1_1__31_0__26_;
  wire AES_CORE_DATAPATH__0bkp_1_1__31_0__27_;
  wire AES_CORE_DATAPATH__0bkp_1_1__31_0__28_;
  wire AES_CORE_DATAPATH__0bkp_1_1__31_0__29_;
  wire AES_CORE_DATAPATH__0bkp_1_1__31_0__2_;
  wire AES_CORE_DATAPATH__0bkp_1_1__31_0__30_;
  wire AES_CORE_DATAPATH__0bkp_1_1__31_0__31_;
  wire AES_CORE_DATAPATH__0bkp_1_1__31_0__3_;
  wire AES_CORE_DATAPATH__0bkp_1_1__31_0__4_;
  wire AES_CORE_DATAPATH__0bkp_1_1__31_0__5_;
  wire AES_CORE_DATAPATH__0bkp_1_1__31_0__6_;
  wire AES_CORE_DATAPATH__0bkp_1_1__31_0__7_;
  wire AES_CORE_DATAPATH__0bkp_1_1__31_0__8_;
  wire AES_CORE_DATAPATH__0bkp_1_1__31_0__9_;
  wire AES_CORE_DATAPATH__0bkp_1_2__31_0__0_;
  wire AES_CORE_DATAPATH__0bkp_1_2__31_0__10_;
  wire AES_CORE_DATAPATH__0bkp_1_2__31_0__11_;
  wire AES_CORE_DATAPATH__0bkp_1_2__31_0__12_;
  wire AES_CORE_DATAPATH__0bkp_1_2__31_0__13_;
  wire AES_CORE_DATAPATH__0bkp_1_2__31_0__14_;
  wire AES_CORE_DATAPATH__0bkp_1_2__31_0__15_;
  wire AES_CORE_DATAPATH__0bkp_1_2__31_0__16_;
  wire AES_CORE_DATAPATH__0bkp_1_2__31_0__17_;
  wire AES_CORE_DATAPATH__0bkp_1_2__31_0__18_;
  wire AES_CORE_DATAPATH__0bkp_1_2__31_0__19_;
  wire AES_CORE_DATAPATH__0bkp_1_2__31_0__1_;
  wire AES_CORE_DATAPATH__0bkp_1_2__31_0__20_;
  wire AES_CORE_DATAPATH__0bkp_1_2__31_0__21_;
  wire AES_CORE_DATAPATH__0bkp_1_2__31_0__22_;
  wire AES_CORE_DATAPATH__0bkp_1_2__31_0__23_;
  wire AES_CORE_DATAPATH__0bkp_1_2__31_0__24_;
  wire AES_CORE_DATAPATH__0bkp_1_2__31_0__25_;
  wire AES_CORE_DATAPATH__0bkp_1_2__31_0__26_;
  wire AES_CORE_DATAPATH__0bkp_1_2__31_0__27_;
  wire AES_CORE_DATAPATH__0bkp_1_2__31_0__28_;
  wire AES_CORE_DATAPATH__0bkp_1_2__31_0__29_;
  wire AES_CORE_DATAPATH__0bkp_1_2__31_0__2_;
  wire AES_CORE_DATAPATH__0bkp_1_2__31_0__30_;
  wire AES_CORE_DATAPATH__0bkp_1_2__31_0__31_;
  wire AES_CORE_DATAPATH__0bkp_1_2__31_0__3_;
  wire AES_CORE_DATAPATH__0bkp_1_2__31_0__4_;
  wire AES_CORE_DATAPATH__0bkp_1_2__31_0__5_;
  wire AES_CORE_DATAPATH__0bkp_1_2__31_0__6_;
  wire AES_CORE_DATAPATH__0bkp_1_2__31_0__7_;
  wire AES_CORE_DATAPATH__0bkp_1_2__31_0__8_;
  wire AES_CORE_DATAPATH__0bkp_1_2__31_0__9_;
  wire AES_CORE_DATAPATH__0bkp_1_3__31_0__0_;
  wire AES_CORE_DATAPATH__0bkp_1_3__31_0__10_;
  wire AES_CORE_DATAPATH__0bkp_1_3__31_0__11_;
  wire AES_CORE_DATAPATH__0bkp_1_3__31_0__12_;
  wire AES_CORE_DATAPATH__0bkp_1_3__31_0__13_;
  wire AES_CORE_DATAPATH__0bkp_1_3__31_0__14_;
  wire AES_CORE_DATAPATH__0bkp_1_3__31_0__15_;
  wire AES_CORE_DATAPATH__0bkp_1_3__31_0__16_;
  wire AES_CORE_DATAPATH__0bkp_1_3__31_0__17_;
  wire AES_CORE_DATAPATH__0bkp_1_3__31_0__18_;
  wire AES_CORE_DATAPATH__0bkp_1_3__31_0__19_;
  wire AES_CORE_DATAPATH__0bkp_1_3__31_0__1_;
  wire AES_CORE_DATAPATH__0bkp_1_3__31_0__20_;
  wire AES_CORE_DATAPATH__0bkp_1_3__31_0__21_;
  wire AES_CORE_DATAPATH__0bkp_1_3__31_0__22_;
  wire AES_CORE_DATAPATH__0bkp_1_3__31_0__23_;
  wire AES_CORE_DATAPATH__0bkp_1_3__31_0__24_;
  wire AES_CORE_DATAPATH__0bkp_1_3__31_0__25_;
  wire AES_CORE_DATAPATH__0bkp_1_3__31_0__26_;
  wire AES_CORE_DATAPATH__0bkp_1_3__31_0__27_;
  wire AES_CORE_DATAPATH__0bkp_1_3__31_0__28_;
  wire AES_CORE_DATAPATH__0bkp_1_3__31_0__29_;
  wire AES_CORE_DATAPATH__0bkp_1_3__31_0__2_;
  wire AES_CORE_DATAPATH__0bkp_1_3__31_0__30_;
  wire AES_CORE_DATAPATH__0bkp_1_3__31_0__31_;
  wire AES_CORE_DATAPATH__0bkp_1_3__31_0__3_;
  wire AES_CORE_DATAPATH__0bkp_1_3__31_0__4_;
  wire AES_CORE_DATAPATH__0bkp_1_3__31_0__5_;
  wire AES_CORE_DATAPATH__0bkp_1_3__31_0__6_;
  wire AES_CORE_DATAPATH__0bkp_1_3__31_0__7_;
  wire AES_CORE_DATAPATH__0bkp_1_3__31_0__8_;
  wire AES_CORE_DATAPATH__0bkp_1_3__31_0__9_;
  wire AES_CORE_DATAPATH__0bkp_1__31_0__0_;
  wire AES_CORE_DATAPATH__0bkp_1__31_0__10_;
  wire AES_CORE_DATAPATH__0bkp_1__31_0__11_;
  wire AES_CORE_DATAPATH__0bkp_1__31_0__12_;
  wire AES_CORE_DATAPATH__0bkp_1__31_0__13_;
  wire AES_CORE_DATAPATH__0bkp_1__31_0__14_;
  wire AES_CORE_DATAPATH__0bkp_1__31_0__15_;
  wire AES_CORE_DATAPATH__0bkp_1__31_0__16_;
  wire AES_CORE_DATAPATH__0bkp_1__31_0__17_;
  wire AES_CORE_DATAPATH__0bkp_1__31_0__18_;
  wire AES_CORE_DATAPATH__0bkp_1__31_0__19_;
  wire AES_CORE_DATAPATH__0bkp_1__31_0__1_;
  wire AES_CORE_DATAPATH__0bkp_1__31_0__20_;
  wire AES_CORE_DATAPATH__0bkp_1__31_0__21_;
  wire AES_CORE_DATAPATH__0bkp_1__31_0__22_;
  wire AES_CORE_DATAPATH__0bkp_1__31_0__23_;
  wire AES_CORE_DATAPATH__0bkp_1__31_0__24_;
  wire AES_CORE_DATAPATH__0bkp_1__31_0__25_;
  wire AES_CORE_DATAPATH__0bkp_1__31_0__26_;
  wire AES_CORE_DATAPATH__0bkp_1__31_0__27_;
  wire AES_CORE_DATAPATH__0bkp_1__31_0__28_;
  wire AES_CORE_DATAPATH__0bkp_1__31_0__29_;
  wire AES_CORE_DATAPATH__0bkp_1__31_0__2_;
  wire AES_CORE_DATAPATH__0bkp_1__31_0__30_;
  wire AES_CORE_DATAPATH__0bkp_1__31_0__31_;
  wire AES_CORE_DATAPATH__0bkp_1__31_0__3_;
  wire AES_CORE_DATAPATH__0bkp_1__31_0__4_;
  wire AES_CORE_DATAPATH__0bkp_1__31_0__5_;
  wire AES_CORE_DATAPATH__0bkp_1__31_0__6_;
  wire AES_CORE_DATAPATH__0bkp_1__31_0__7_;
  wire AES_CORE_DATAPATH__0bkp_1__31_0__8_;
  wire AES_CORE_DATAPATH__0bkp_1__31_0__9_;
  wire AES_CORE_DATAPATH__0bkp_2__31_0__0_;
  wire AES_CORE_DATAPATH__0bkp_2__31_0__10_;
  wire AES_CORE_DATAPATH__0bkp_2__31_0__11_;
  wire AES_CORE_DATAPATH__0bkp_2__31_0__12_;
  wire AES_CORE_DATAPATH__0bkp_2__31_0__13_;
  wire AES_CORE_DATAPATH__0bkp_2__31_0__14_;
  wire AES_CORE_DATAPATH__0bkp_2__31_0__15_;
  wire AES_CORE_DATAPATH__0bkp_2__31_0__16_;
  wire AES_CORE_DATAPATH__0bkp_2__31_0__17_;
  wire AES_CORE_DATAPATH__0bkp_2__31_0__18_;
  wire AES_CORE_DATAPATH__0bkp_2__31_0__19_;
  wire AES_CORE_DATAPATH__0bkp_2__31_0__1_;
  wire AES_CORE_DATAPATH__0bkp_2__31_0__20_;
  wire AES_CORE_DATAPATH__0bkp_2__31_0__21_;
  wire AES_CORE_DATAPATH__0bkp_2__31_0__22_;
  wire AES_CORE_DATAPATH__0bkp_2__31_0__23_;
  wire AES_CORE_DATAPATH__0bkp_2__31_0__24_;
  wire AES_CORE_DATAPATH__0bkp_2__31_0__25_;
  wire AES_CORE_DATAPATH__0bkp_2__31_0__26_;
  wire AES_CORE_DATAPATH__0bkp_2__31_0__27_;
  wire AES_CORE_DATAPATH__0bkp_2__31_0__28_;
  wire AES_CORE_DATAPATH__0bkp_2__31_0__29_;
  wire AES_CORE_DATAPATH__0bkp_2__31_0__2_;
  wire AES_CORE_DATAPATH__0bkp_2__31_0__30_;
  wire AES_CORE_DATAPATH__0bkp_2__31_0__31_;
  wire AES_CORE_DATAPATH__0bkp_2__31_0__3_;
  wire AES_CORE_DATAPATH__0bkp_2__31_0__4_;
  wire AES_CORE_DATAPATH__0bkp_2__31_0__5_;
  wire AES_CORE_DATAPATH__0bkp_2__31_0__6_;
  wire AES_CORE_DATAPATH__0bkp_2__31_0__7_;
  wire AES_CORE_DATAPATH__0bkp_2__31_0__8_;
  wire AES_CORE_DATAPATH__0bkp_2__31_0__9_;
  wire AES_CORE_DATAPATH__0bkp_3__31_0__0_;
  wire AES_CORE_DATAPATH__0bkp_3__31_0__10_;
  wire AES_CORE_DATAPATH__0bkp_3__31_0__11_;
  wire AES_CORE_DATAPATH__0bkp_3__31_0__12_;
  wire AES_CORE_DATAPATH__0bkp_3__31_0__13_;
  wire AES_CORE_DATAPATH__0bkp_3__31_0__14_;
  wire AES_CORE_DATAPATH__0bkp_3__31_0__15_;
  wire AES_CORE_DATAPATH__0bkp_3__31_0__16_;
  wire AES_CORE_DATAPATH__0bkp_3__31_0__17_;
  wire AES_CORE_DATAPATH__0bkp_3__31_0__18_;
  wire AES_CORE_DATAPATH__0bkp_3__31_0__19_;
  wire AES_CORE_DATAPATH__0bkp_3__31_0__1_;
  wire AES_CORE_DATAPATH__0bkp_3__31_0__20_;
  wire AES_CORE_DATAPATH__0bkp_3__31_0__21_;
  wire AES_CORE_DATAPATH__0bkp_3__31_0__22_;
  wire AES_CORE_DATAPATH__0bkp_3__31_0__23_;
  wire AES_CORE_DATAPATH__0bkp_3__31_0__24_;
  wire AES_CORE_DATAPATH__0bkp_3__31_0__25_;
  wire AES_CORE_DATAPATH__0bkp_3__31_0__26_;
  wire AES_CORE_DATAPATH__0bkp_3__31_0__27_;
  wire AES_CORE_DATAPATH__0bkp_3__31_0__28_;
  wire AES_CORE_DATAPATH__0bkp_3__31_0__29_;
  wire AES_CORE_DATAPATH__0bkp_3__31_0__2_;
  wire AES_CORE_DATAPATH__0bkp_3__31_0__30_;
  wire AES_CORE_DATAPATH__0bkp_3__31_0__31_;
  wire AES_CORE_DATAPATH__0bkp_3__31_0__3_;
  wire AES_CORE_DATAPATH__0bkp_3__31_0__4_;
  wire AES_CORE_DATAPATH__0bkp_3__31_0__5_;
  wire AES_CORE_DATAPATH__0bkp_3__31_0__6_;
  wire AES_CORE_DATAPATH__0bkp_3__31_0__7_;
  wire AES_CORE_DATAPATH__0bkp_3__31_0__8_;
  wire AES_CORE_DATAPATH__0bkp_3__31_0__9_;
  wire AES_CORE_DATAPATH__0col_0__31_0__0_;
  wire AES_CORE_DATAPATH__0col_0__31_0__10_;
  wire AES_CORE_DATAPATH__0col_0__31_0__11_;
  wire AES_CORE_DATAPATH__0col_0__31_0__12_;
  wire AES_CORE_DATAPATH__0col_0__31_0__13_;
  wire AES_CORE_DATAPATH__0col_0__31_0__14_;
  wire AES_CORE_DATAPATH__0col_0__31_0__15_;
  wire AES_CORE_DATAPATH__0col_0__31_0__16_;
  wire AES_CORE_DATAPATH__0col_0__31_0__17_;
  wire AES_CORE_DATAPATH__0col_0__31_0__18_;
  wire AES_CORE_DATAPATH__0col_0__31_0__19_;
  wire AES_CORE_DATAPATH__0col_0__31_0__1_;
  wire AES_CORE_DATAPATH__0col_0__31_0__20_;
  wire AES_CORE_DATAPATH__0col_0__31_0__21_;
  wire AES_CORE_DATAPATH__0col_0__31_0__22_;
  wire AES_CORE_DATAPATH__0col_0__31_0__23_;
  wire AES_CORE_DATAPATH__0col_0__31_0__24_;
  wire AES_CORE_DATAPATH__0col_0__31_0__25_;
  wire AES_CORE_DATAPATH__0col_0__31_0__26_;
  wire AES_CORE_DATAPATH__0col_0__31_0__27_;
  wire AES_CORE_DATAPATH__0col_0__31_0__28_;
  wire AES_CORE_DATAPATH__0col_0__31_0__29_;
  wire AES_CORE_DATAPATH__0col_0__31_0__2_;
  wire AES_CORE_DATAPATH__0col_0__31_0__30_;
  wire AES_CORE_DATAPATH__0col_0__31_0__31_;
  wire AES_CORE_DATAPATH__0col_0__31_0__3_;
  wire AES_CORE_DATAPATH__0col_0__31_0__4_;
  wire AES_CORE_DATAPATH__0col_0__31_0__5_;
  wire AES_CORE_DATAPATH__0col_0__31_0__6_;
  wire AES_CORE_DATAPATH__0col_0__31_0__7_;
  wire AES_CORE_DATAPATH__0col_0__31_0__8_;
  wire AES_CORE_DATAPATH__0col_0__31_0__9_;
  wire AES_CORE_DATAPATH__0col_1__31_0__0_;
  wire AES_CORE_DATAPATH__0col_1__31_0__10_;
  wire AES_CORE_DATAPATH__0col_1__31_0__11_;
  wire AES_CORE_DATAPATH__0col_1__31_0__12_;
  wire AES_CORE_DATAPATH__0col_1__31_0__13_;
  wire AES_CORE_DATAPATH__0col_1__31_0__14_;
  wire AES_CORE_DATAPATH__0col_1__31_0__15_;
  wire AES_CORE_DATAPATH__0col_1__31_0__16_;
  wire AES_CORE_DATAPATH__0col_1__31_0__17_;
  wire AES_CORE_DATAPATH__0col_1__31_0__18_;
  wire AES_CORE_DATAPATH__0col_1__31_0__19_;
  wire AES_CORE_DATAPATH__0col_1__31_0__1_;
  wire AES_CORE_DATAPATH__0col_1__31_0__20_;
  wire AES_CORE_DATAPATH__0col_1__31_0__21_;
  wire AES_CORE_DATAPATH__0col_1__31_0__22_;
  wire AES_CORE_DATAPATH__0col_1__31_0__23_;
  wire AES_CORE_DATAPATH__0col_1__31_0__24_;
  wire AES_CORE_DATAPATH__0col_1__31_0__25_;
  wire AES_CORE_DATAPATH__0col_1__31_0__26_;
  wire AES_CORE_DATAPATH__0col_1__31_0__27_;
  wire AES_CORE_DATAPATH__0col_1__31_0__28_;
  wire AES_CORE_DATAPATH__0col_1__31_0__29_;
  wire AES_CORE_DATAPATH__0col_1__31_0__2_;
  wire AES_CORE_DATAPATH__0col_1__31_0__30_;
  wire AES_CORE_DATAPATH__0col_1__31_0__31_;
  wire AES_CORE_DATAPATH__0col_1__31_0__3_;
  wire AES_CORE_DATAPATH__0col_1__31_0__4_;
  wire AES_CORE_DATAPATH__0col_1__31_0__5_;
  wire AES_CORE_DATAPATH__0col_1__31_0__6_;
  wire AES_CORE_DATAPATH__0col_1__31_0__7_;
  wire AES_CORE_DATAPATH__0col_1__31_0__8_;
  wire AES_CORE_DATAPATH__0col_1__31_0__9_;
  wire AES_CORE_DATAPATH__0col_2__31_0__0_;
  wire AES_CORE_DATAPATH__0col_2__31_0__10_;
  wire AES_CORE_DATAPATH__0col_2__31_0__11_;
  wire AES_CORE_DATAPATH__0col_2__31_0__12_;
  wire AES_CORE_DATAPATH__0col_2__31_0__13_;
  wire AES_CORE_DATAPATH__0col_2__31_0__14_;
  wire AES_CORE_DATAPATH__0col_2__31_0__15_;
  wire AES_CORE_DATAPATH__0col_2__31_0__16_;
  wire AES_CORE_DATAPATH__0col_2__31_0__17_;
  wire AES_CORE_DATAPATH__0col_2__31_0__18_;
  wire AES_CORE_DATAPATH__0col_2__31_0__19_;
  wire AES_CORE_DATAPATH__0col_2__31_0__1_;
  wire AES_CORE_DATAPATH__0col_2__31_0__20_;
  wire AES_CORE_DATAPATH__0col_2__31_0__21_;
  wire AES_CORE_DATAPATH__0col_2__31_0__22_;
  wire AES_CORE_DATAPATH__0col_2__31_0__23_;
  wire AES_CORE_DATAPATH__0col_2__31_0__24_;
  wire AES_CORE_DATAPATH__0col_2__31_0__25_;
  wire AES_CORE_DATAPATH__0col_2__31_0__26_;
  wire AES_CORE_DATAPATH__0col_2__31_0__27_;
  wire AES_CORE_DATAPATH__0col_2__31_0__28_;
  wire AES_CORE_DATAPATH__0col_2__31_0__29_;
  wire AES_CORE_DATAPATH__0col_2__31_0__2_;
  wire AES_CORE_DATAPATH__0col_2__31_0__30_;
  wire AES_CORE_DATAPATH__0col_2__31_0__31_;
  wire AES_CORE_DATAPATH__0col_2__31_0__3_;
  wire AES_CORE_DATAPATH__0col_2__31_0__4_;
  wire AES_CORE_DATAPATH__0col_2__31_0__5_;
  wire AES_CORE_DATAPATH__0col_2__31_0__6_;
  wire AES_CORE_DATAPATH__0col_2__31_0__7_;
  wire AES_CORE_DATAPATH__0col_2__31_0__8_;
  wire AES_CORE_DATAPATH__0col_2__31_0__9_;
  wire AES_CORE_DATAPATH__0col_3__31_0__0_;
  wire AES_CORE_DATAPATH__0col_3__31_0__10_;
  wire AES_CORE_DATAPATH__0col_3__31_0__11_;
  wire AES_CORE_DATAPATH__0col_3__31_0__12_;
  wire AES_CORE_DATAPATH__0col_3__31_0__13_;
  wire AES_CORE_DATAPATH__0col_3__31_0__14_;
  wire AES_CORE_DATAPATH__0col_3__31_0__15_;
  wire AES_CORE_DATAPATH__0col_3__31_0__16_;
  wire AES_CORE_DATAPATH__0col_3__31_0__17_;
  wire AES_CORE_DATAPATH__0col_3__31_0__18_;
  wire AES_CORE_DATAPATH__0col_3__31_0__19_;
  wire AES_CORE_DATAPATH__0col_3__31_0__1_;
  wire AES_CORE_DATAPATH__0col_3__31_0__20_;
  wire AES_CORE_DATAPATH__0col_3__31_0__21_;
  wire AES_CORE_DATAPATH__0col_3__31_0__22_;
  wire AES_CORE_DATAPATH__0col_3__31_0__23_;
  wire AES_CORE_DATAPATH__0col_3__31_0__24_;
  wire AES_CORE_DATAPATH__0col_3__31_0__25_;
  wire AES_CORE_DATAPATH__0col_3__31_0__26_;
  wire AES_CORE_DATAPATH__0col_3__31_0__27_;
  wire AES_CORE_DATAPATH__0col_3__31_0__28_;
  wire AES_CORE_DATAPATH__0col_3__31_0__29_;
  wire AES_CORE_DATAPATH__0col_3__31_0__2_;
  wire AES_CORE_DATAPATH__0col_3__31_0__30_;
  wire AES_CORE_DATAPATH__0col_3__31_0__31_;
  wire AES_CORE_DATAPATH__0col_3__31_0__3_;
  wire AES_CORE_DATAPATH__0col_3__31_0__4_;
  wire AES_CORE_DATAPATH__0col_3__31_0__5_;
  wire AES_CORE_DATAPATH__0col_3__31_0__6_;
  wire AES_CORE_DATAPATH__0col_3__31_0__7_;
  wire AES_CORE_DATAPATH__0col_3__31_0__8_;
  wire AES_CORE_DATAPATH__0col_3__31_0__9_;
  wire AES_CORE_DATAPATH__0iv_0__31_0__0_;
  wire AES_CORE_DATAPATH__0iv_0__31_0__10_;
  wire AES_CORE_DATAPATH__0iv_0__31_0__11_;
  wire AES_CORE_DATAPATH__0iv_0__31_0__12_;
  wire AES_CORE_DATAPATH__0iv_0__31_0__13_;
  wire AES_CORE_DATAPATH__0iv_0__31_0__14_;
  wire AES_CORE_DATAPATH__0iv_0__31_0__15_;
  wire AES_CORE_DATAPATH__0iv_0__31_0__16_;
  wire AES_CORE_DATAPATH__0iv_0__31_0__17_;
  wire AES_CORE_DATAPATH__0iv_0__31_0__18_;
  wire AES_CORE_DATAPATH__0iv_0__31_0__19_;
  wire AES_CORE_DATAPATH__0iv_0__31_0__1_;
  wire AES_CORE_DATAPATH__0iv_0__31_0__20_;
  wire AES_CORE_DATAPATH__0iv_0__31_0__21_;
  wire AES_CORE_DATAPATH__0iv_0__31_0__22_;
  wire AES_CORE_DATAPATH__0iv_0__31_0__23_;
  wire AES_CORE_DATAPATH__0iv_0__31_0__24_;
  wire AES_CORE_DATAPATH__0iv_0__31_0__25_;
  wire AES_CORE_DATAPATH__0iv_0__31_0__26_;
  wire AES_CORE_DATAPATH__0iv_0__31_0__27_;
  wire AES_CORE_DATAPATH__0iv_0__31_0__28_;
  wire AES_CORE_DATAPATH__0iv_0__31_0__29_;
  wire AES_CORE_DATAPATH__0iv_0__31_0__2_;
  wire AES_CORE_DATAPATH__0iv_0__31_0__30_;
  wire AES_CORE_DATAPATH__0iv_0__31_0__31_;
  wire AES_CORE_DATAPATH__0iv_0__31_0__3_;
  wire AES_CORE_DATAPATH__0iv_0__31_0__4_;
  wire AES_CORE_DATAPATH__0iv_0__31_0__5_;
  wire AES_CORE_DATAPATH__0iv_0__31_0__6_;
  wire AES_CORE_DATAPATH__0iv_0__31_0__7_;
  wire AES_CORE_DATAPATH__0iv_0__31_0__8_;
  wire AES_CORE_DATAPATH__0iv_0__31_0__9_;
  wire AES_CORE_DATAPATH__0iv_1__31_0__0_;
  wire AES_CORE_DATAPATH__0iv_1__31_0__10_;
  wire AES_CORE_DATAPATH__0iv_1__31_0__11_;
  wire AES_CORE_DATAPATH__0iv_1__31_0__12_;
  wire AES_CORE_DATAPATH__0iv_1__31_0__13_;
  wire AES_CORE_DATAPATH__0iv_1__31_0__14_;
  wire AES_CORE_DATAPATH__0iv_1__31_0__15_;
  wire AES_CORE_DATAPATH__0iv_1__31_0__16_;
  wire AES_CORE_DATAPATH__0iv_1__31_0__17_;
  wire AES_CORE_DATAPATH__0iv_1__31_0__18_;
  wire AES_CORE_DATAPATH__0iv_1__31_0__19_;
  wire AES_CORE_DATAPATH__0iv_1__31_0__1_;
  wire AES_CORE_DATAPATH__0iv_1__31_0__20_;
  wire AES_CORE_DATAPATH__0iv_1__31_0__21_;
  wire AES_CORE_DATAPATH__0iv_1__31_0__22_;
  wire AES_CORE_DATAPATH__0iv_1__31_0__23_;
  wire AES_CORE_DATAPATH__0iv_1__31_0__24_;
  wire AES_CORE_DATAPATH__0iv_1__31_0__25_;
  wire AES_CORE_DATAPATH__0iv_1__31_0__26_;
  wire AES_CORE_DATAPATH__0iv_1__31_0__27_;
  wire AES_CORE_DATAPATH__0iv_1__31_0__28_;
  wire AES_CORE_DATAPATH__0iv_1__31_0__29_;
  wire AES_CORE_DATAPATH__0iv_1__31_0__2_;
  wire AES_CORE_DATAPATH__0iv_1__31_0__30_;
  wire AES_CORE_DATAPATH__0iv_1__31_0__31_;
  wire AES_CORE_DATAPATH__0iv_1__31_0__3_;
  wire AES_CORE_DATAPATH__0iv_1__31_0__4_;
  wire AES_CORE_DATAPATH__0iv_1__31_0__5_;
  wire AES_CORE_DATAPATH__0iv_1__31_0__6_;
  wire AES_CORE_DATAPATH__0iv_1__31_0__7_;
  wire AES_CORE_DATAPATH__0iv_1__31_0__8_;
  wire AES_CORE_DATAPATH__0iv_1__31_0__9_;
  wire AES_CORE_DATAPATH__0iv_2__31_0__0_;
  wire AES_CORE_DATAPATH__0iv_2__31_0__10_;
  wire AES_CORE_DATAPATH__0iv_2__31_0__11_;
  wire AES_CORE_DATAPATH__0iv_2__31_0__12_;
  wire AES_CORE_DATAPATH__0iv_2__31_0__13_;
  wire AES_CORE_DATAPATH__0iv_2__31_0__14_;
  wire AES_CORE_DATAPATH__0iv_2__31_0__15_;
  wire AES_CORE_DATAPATH__0iv_2__31_0__16_;
  wire AES_CORE_DATAPATH__0iv_2__31_0__17_;
  wire AES_CORE_DATAPATH__0iv_2__31_0__18_;
  wire AES_CORE_DATAPATH__0iv_2__31_0__19_;
  wire AES_CORE_DATAPATH__0iv_2__31_0__1_;
  wire AES_CORE_DATAPATH__0iv_2__31_0__20_;
  wire AES_CORE_DATAPATH__0iv_2__31_0__21_;
  wire AES_CORE_DATAPATH__0iv_2__31_0__22_;
  wire AES_CORE_DATAPATH__0iv_2__31_0__23_;
  wire AES_CORE_DATAPATH__0iv_2__31_0__24_;
  wire AES_CORE_DATAPATH__0iv_2__31_0__25_;
  wire AES_CORE_DATAPATH__0iv_2__31_0__26_;
  wire AES_CORE_DATAPATH__0iv_2__31_0__27_;
  wire AES_CORE_DATAPATH__0iv_2__31_0__28_;
  wire AES_CORE_DATAPATH__0iv_2__31_0__29_;
  wire AES_CORE_DATAPATH__0iv_2__31_0__2_;
  wire AES_CORE_DATAPATH__0iv_2__31_0__30_;
  wire AES_CORE_DATAPATH__0iv_2__31_0__31_;
  wire AES_CORE_DATAPATH__0iv_2__31_0__3_;
  wire AES_CORE_DATAPATH__0iv_2__31_0__4_;
  wire AES_CORE_DATAPATH__0iv_2__31_0__5_;
  wire AES_CORE_DATAPATH__0iv_2__31_0__6_;
  wire AES_CORE_DATAPATH__0iv_2__31_0__7_;
  wire AES_CORE_DATAPATH__0iv_2__31_0__8_;
  wire AES_CORE_DATAPATH__0iv_2__31_0__9_;
  wire AES_CORE_DATAPATH__0iv_3__31_0__0_;
  wire AES_CORE_DATAPATH__0iv_3__31_0__10_;
  wire AES_CORE_DATAPATH__0iv_3__31_0__11_;
  wire AES_CORE_DATAPATH__0iv_3__31_0__12_;
  wire AES_CORE_DATAPATH__0iv_3__31_0__13_;
  wire AES_CORE_DATAPATH__0iv_3__31_0__14_;
  wire AES_CORE_DATAPATH__0iv_3__31_0__15_;
  wire AES_CORE_DATAPATH__0iv_3__31_0__16_;
  wire AES_CORE_DATAPATH__0iv_3__31_0__17_;
  wire AES_CORE_DATAPATH__0iv_3__31_0__18_;
  wire AES_CORE_DATAPATH__0iv_3__31_0__19_;
  wire AES_CORE_DATAPATH__0iv_3__31_0__1_;
  wire AES_CORE_DATAPATH__0iv_3__31_0__20_;
  wire AES_CORE_DATAPATH__0iv_3__31_0__21_;
  wire AES_CORE_DATAPATH__0iv_3__31_0__22_;
  wire AES_CORE_DATAPATH__0iv_3__31_0__23_;
  wire AES_CORE_DATAPATH__0iv_3__31_0__24_;
  wire AES_CORE_DATAPATH__0iv_3__31_0__25_;
  wire AES_CORE_DATAPATH__0iv_3__31_0__26_;
  wire AES_CORE_DATAPATH__0iv_3__31_0__27_;
  wire AES_CORE_DATAPATH__0iv_3__31_0__28_;
  wire AES_CORE_DATAPATH__0iv_3__31_0__29_;
  wire AES_CORE_DATAPATH__0iv_3__31_0__2_;
  wire AES_CORE_DATAPATH__0iv_3__31_0__30_;
  wire AES_CORE_DATAPATH__0iv_3__31_0__31_;
  wire AES_CORE_DATAPATH__0iv_3__31_0__3_;
  wire AES_CORE_DATAPATH__0iv_3__31_0__4_;
  wire AES_CORE_DATAPATH__0iv_3__31_0__5_;
  wire AES_CORE_DATAPATH__0iv_3__31_0__6_;
  wire AES_CORE_DATAPATH__0iv_3__31_0__7_;
  wire AES_CORE_DATAPATH__0iv_3__31_0__8_;
  wire AES_CORE_DATAPATH__0iv_3__31_0__9_;
  wire AES_CORE_DATAPATH__0key_0__31_0__0_;
  wire AES_CORE_DATAPATH__0key_0__31_0__10_;
  wire AES_CORE_DATAPATH__0key_0__31_0__11_;
  wire AES_CORE_DATAPATH__0key_0__31_0__12_;
  wire AES_CORE_DATAPATH__0key_0__31_0__13_;
  wire AES_CORE_DATAPATH__0key_0__31_0__14_;
  wire AES_CORE_DATAPATH__0key_0__31_0__15_;
  wire AES_CORE_DATAPATH__0key_0__31_0__16_;
  wire AES_CORE_DATAPATH__0key_0__31_0__17_;
  wire AES_CORE_DATAPATH__0key_0__31_0__18_;
  wire AES_CORE_DATAPATH__0key_0__31_0__19_;
  wire AES_CORE_DATAPATH__0key_0__31_0__1_;
  wire AES_CORE_DATAPATH__0key_0__31_0__20_;
  wire AES_CORE_DATAPATH__0key_0__31_0__21_;
  wire AES_CORE_DATAPATH__0key_0__31_0__22_;
  wire AES_CORE_DATAPATH__0key_0__31_0__23_;
  wire AES_CORE_DATAPATH__0key_0__31_0__24_;
  wire AES_CORE_DATAPATH__0key_0__31_0__25_;
  wire AES_CORE_DATAPATH__0key_0__31_0__26_;
  wire AES_CORE_DATAPATH__0key_0__31_0__27_;
  wire AES_CORE_DATAPATH__0key_0__31_0__28_;
  wire AES_CORE_DATAPATH__0key_0__31_0__29_;
  wire AES_CORE_DATAPATH__0key_0__31_0__2_;
  wire AES_CORE_DATAPATH__0key_0__31_0__30_;
  wire AES_CORE_DATAPATH__0key_0__31_0__31_;
  wire AES_CORE_DATAPATH__0key_0__31_0__3_;
  wire AES_CORE_DATAPATH__0key_0__31_0__4_;
  wire AES_CORE_DATAPATH__0key_0__31_0__5_;
  wire AES_CORE_DATAPATH__0key_0__31_0__6_;
  wire AES_CORE_DATAPATH__0key_0__31_0__7_;
  wire AES_CORE_DATAPATH__0key_0__31_0__8_;
  wire AES_CORE_DATAPATH__0key_0__31_0__9_;
  wire AES_CORE_DATAPATH__0key_1__31_0__0_;
  wire AES_CORE_DATAPATH__0key_1__31_0__10_;
  wire AES_CORE_DATAPATH__0key_1__31_0__11_;
  wire AES_CORE_DATAPATH__0key_1__31_0__12_;
  wire AES_CORE_DATAPATH__0key_1__31_0__13_;
  wire AES_CORE_DATAPATH__0key_1__31_0__14_;
  wire AES_CORE_DATAPATH__0key_1__31_0__15_;
  wire AES_CORE_DATAPATH__0key_1__31_0__16_;
  wire AES_CORE_DATAPATH__0key_1__31_0__17_;
  wire AES_CORE_DATAPATH__0key_1__31_0__18_;
  wire AES_CORE_DATAPATH__0key_1__31_0__19_;
  wire AES_CORE_DATAPATH__0key_1__31_0__1_;
  wire AES_CORE_DATAPATH__0key_1__31_0__20_;
  wire AES_CORE_DATAPATH__0key_1__31_0__21_;
  wire AES_CORE_DATAPATH__0key_1__31_0__22_;
  wire AES_CORE_DATAPATH__0key_1__31_0__23_;
  wire AES_CORE_DATAPATH__0key_1__31_0__24_;
  wire AES_CORE_DATAPATH__0key_1__31_0__25_;
  wire AES_CORE_DATAPATH__0key_1__31_0__26_;
  wire AES_CORE_DATAPATH__0key_1__31_0__27_;
  wire AES_CORE_DATAPATH__0key_1__31_0__28_;
  wire AES_CORE_DATAPATH__0key_1__31_0__29_;
  wire AES_CORE_DATAPATH__0key_1__31_0__2_;
  wire AES_CORE_DATAPATH__0key_1__31_0__30_;
  wire AES_CORE_DATAPATH__0key_1__31_0__31_;
  wire AES_CORE_DATAPATH__0key_1__31_0__3_;
  wire AES_CORE_DATAPATH__0key_1__31_0__4_;
  wire AES_CORE_DATAPATH__0key_1__31_0__5_;
  wire AES_CORE_DATAPATH__0key_1__31_0__6_;
  wire AES_CORE_DATAPATH__0key_1__31_0__7_;
  wire AES_CORE_DATAPATH__0key_1__31_0__8_;
  wire AES_CORE_DATAPATH__0key_1__31_0__9_;
  wire AES_CORE_DATAPATH__0key_2__31_0__0_;
  wire AES_CORE_DATAPATH__0key_2__31_0__10_;
  wire AES_CORE_DATAPATH__0key_2__31_0__11_;
  wire AES_CORE_DATAPATH__0key_2__31_0__12_;
  wire AES_CORE_DATAPATH__0key_2__31_0__13_;
  wire AES_CORE_DATAPATH__0key_2__31_0__14_;
  wire AES_CORE_DATAPATH__0key_2__31_0__15_;
  wire AES_CORE_DATAPATH__0key_2__31_0__16_;
  wire AES_CORE_DATAPATH__0key_2__31_0__17_;
  wire AES_CORE_DATAPATH__0key_2__31_0__18_;
  wire AES_CORE_DATAPATH__0key_2__31_0__19_;
  wire AES_CORE_DATAPATH__0key_2__31_0__1_;
  wire AES_CORE_DATAPATH__0key_2__31_0__20_;
  wire AES_CORE_DATAPATH__0key_2__31_0__21_;
  wire AES_CORE_DATAPATH__0key_2__31_0__22_;
  wire AES_CORE_DATAPATH__0key_2__31_0__23_;
  wire AES_CORE_DATAPATH__0key_2__31_0__24_;
  wire AES_CORE_DATAPATH__0key_2__31_0__25_;
  wire AES_CORE_DATAPATH__0key_2__31_0__26_;
  wire AES_CORE_DATAPATH__0key_2__31_0__27_;
  wire AES_CORE_DATAPATH__0key_2__31_0__28_;
  wire AES_CORE_DATAPATH__0key_2__31_0__29_;
  wire AES_CORE_DATAPATH__0key_2__31_0__2_;
  wire AES_CORE_DATAPATH__0key_2__31_0__30_;
  wire AES_CORE_DATAPATH__0key_2__31_0__31_;
  wire AES_CORE_DATAPATH__0key_2__31_0__3_;
  wire AES_CORE_DATAPATH__0key_2__31_0__4_;
  wire AES_CORE_DATAPATH__0key_2__31_0__5_;
  wire AES_CORE_DATAPATH__0key_2__31_0__6_;
  wire AES_CORE_DATAPATH__0key_2__31_0__7_;
  wire AES_CORE_DATAPATH__0key_2__31_0__8_;
  wire AES_CORE_DATAPATH__0key_2__31_0__9_;
  wire AES_CORE_DATAPATH__0key_3__31_0__0_;
  wire AES_CORE_DATAPATH__0key_3__31_0__10_;
  wire AES_CORE_DATAPATH__0key_3__31_0__11_;
  wire AES_CORE_DATAPATH__0key_3__31_0__12_;
  wire AES_CORE_DATAPATH__0key_3__31_0__13_;
  wire AES_CORE_DATAPATH__0key_3__31_0__14_;
  wire AES_CORE_DATAPATH__0key_3__31_0__15_;
  wire AES_CORE_DATAPATH__0key_3__31_0__16_;
  wire AES_CORE_DATAPATH__0key_3__31_0__17_;
  wire AES_CORE_DATAPATH__0key_3__31_0__18_;
  wire AES_CORE_DATAPATH__0key_3__31_0__19_;
  wire AES_CORE_DATAPATH__0key_3__31_0__1_;
  wire AES_CORE_DATAPATH__0key_3__31_0__20_;
  wire AES_CORE_DATAPATH__0key_3__31_0__21_;
  wire AES_CORE_DATAPATH__0key_3__31_0__22_;
  wire AES_CORE_DATAPATH__0key_3__31_0__23_;
  wire AES_CORE_DATAPATH__0key_3__31_0__24_;
  wire AES_CORE_DATAPATH__0key_3__31_0__25_;
  wire AES_CORE_DATAPATH__0key_3__31_0__26_;
  wire AES_CORE_DATAPATH__0key_3__31_0__27_;
  wire AES_CORE_DATAPATH__0key_3__31_0__28_;
  wire AES_CORE_DATAPATH__0key_3__31_0__29_;
  wire AES_CORE_DATAPATH__0key_3__31_0__2_;
  wire AES_CORE_DATAPATH__0key_3__31_0__30_;
  wire AES_CORE_DATAPATH__0key_3__31_0__31_;
  wire AES_CORE_DATAPATH__0key_3__31_0__3_;
  wire AES_CORE_DATAPATH__0key_3__31_0__4_;
  wire AES_CORE_DATAPATH__0key_3__31_0__5_;
  wire AES_CORE_DATAPATH__0key_3__31_0__6_;
  wire AES_CORE_DATAPATH__0key_3__31_0__7_;
  wire AES_CORE_DATAPATH__0key_3__31_0__8_;
  wire AES_CORE_DATAPATH__0key_3__31_0__9_;
  wire AES_CORE_DATAPATH__0key_host_0__31_0__0_;
  wire AES_CORE_DATAPATH__0key_host_0__31_0__10_;
  wire AES_CORE_DATAPATH__0key_host_0__31_0__11_;
  wire AES_CORE_DATAPATH__0key_host_0__31_0__12_;
  wire AES_CORE_DATAPATH__0key_host_0__31_0__13_;
  wire AES_CORE_DATAPATH__0key_host_0__31_0__14_;
  wire AES_CORE_DATAPATH__0key_host_0__31_0__15_;
  wire AES_CORE_DATAPATH__0key_host_0__31_0__16_;
  wire AES_CORE_DATAPATH__0key_host_0__31_0__17_;
  wire AES_CORE_DATAPATH__0key_host_0__31_0__18_;
  wire AES_CORE_DATAPATH__0key_host_0__31_0__19_;
  wire AES_CORE_DATAPATH__0key_host_0__31_0__1_;
  wire AES_CORE_DATAPATH__0key_host_0__31_0__20_;
  wire AES_CORE_DATAPATH__0key_host_0__31_0__21_;
  wire AES_CORE_DATAPATH__0key_host_0__31_0__22_;
  wire AES_CORE_DATAPATH__0key_host_0__31_0__23_;
  wire AES_CORE_DATAPATH__0key_host_0__31_0__24_;
  wire AES_CORE_DATAPATH__0key_host_0__31_0__25_;
  wire AES_CORE_DATAPATH__0key_host_0__31_0__26_;
  wire AES_CORE_DATAPATH__0key_host_0__31_0__27_;
  wire AES_CORE_DATAPATH__0key_host_0__31_0__28_;
  wire AES_CORE_DATAPATH__0key_host_0__31_0__29_;
  wire AES_CORE_DATAPATH__0key_host_0__31_0__2_;
  wire AES_CORE_DATAPATH__0key_host_0__31_0__30_;
  wire AES_CORE_DATAPATH__0key_host_0__31_0__31_;
  wire AES_CORE_DATAPATH__0key_host_0__31_0__3_;
  wire AES_CORE_DATAPATH__0key_host_0__31_0__4_;
  wire AES_CORE_DATAPATH__0key_host_0__31_0__5_;
  wire AES_CORE_DATAPATH__0key_host_0__31_0__6_;
  wire AES_CORE_DATAPATH__0key_host_0__31_0__7_;
  wire AES_CORE_DATAPATH__0key_host_0__31_0__8_;
  wire AES_CORE_DATAPATH__0key_host_0__31_0__9_;
  wire AES_CORE_DATAPATH__0key_host_1__31_0__0_;
  wire AES_CORE_DATAPATH__0key_host_1__31_0__10_;
  wire AES_CORE_DATAPATH__0key_host_1__31_0__11_;
  wire AES_CORE_DATAPATH__0key_host_1__31_0__12_;
  wire AES_CORE_DATAPATH__0key_host_1__31_0__13_;
  wire AES_CORE_DATAPATH__0key_host_1__31_0__14_;
  wire AES_CORE_DATAPATH__0key_host_1__31_0__15_;
  wire AES_CORE_DATAPATH__0key_host_1__31_0__16_;
  wire AES_CORE_DATAPATH__0key_host_1__31_0__17_;
  wire AES_CORE_DATAPATH__0key_host_1__31_0__18_;
  wire AES_CORE_DATAPATH__0key_host_1__31_0__19_;
  wire AES_CORE_DATAPATH__0key_host_1__31_0__1_;
  wire AES_CORE_DATAPATH__0key_host_1__31_0__20_;
  wire AES_CORE_DATAPATH__0key_host_1__31_0__21_;
  wire AES_CORE_DATAPATH__0key_host_1__31_0__22_;
  wire AES_CORE_DATAPATH__0key_host_1__31_0__23_;
  wire AES_CORE_DATAPATH__0key_host_1__31_0__24_;
  wire AES_CORE_DATAPATH__0key_host_1__31_0__25_;
  wire AES_CORE_DATAPATH__0key_host_1__31_0__26_;
  wire AES_CORE_DATAPATH__0key_host_1__31_0__27_;
  wire AES_CORE_DATAPATH__0key_host_1__31_0__28_;
  wire AES_CORE_DATAPATH__0key_host_1__31_0__29_;
  wire AES_CORE_DATAPATH__0key_host_1__31_0__2_;
  wire AES_CORE_DATAPATH__0key_host_1__31_0__30_;
  wire AES_CORE_DATAPATH__0key_host_1__31_0__31_;
  wire AES_CORE_DATAPATH__0key_host_1__31_0__3_;
  wire AES_CORE_DATAPATH__0key_host_1__31_0__4_;
  wire AES_CORE_DATAPATH__0key_host_1__31_0__5_;
  wire AES_CORE_DATAPATH__0key_host_1__31_0__6_;
  wire AES_CORE_DATAPATH__0key_host_1__31_0__7_;
  wire AES_CORE_DATAPATH__0key_host_1__31_0__8_;
  wire AES_CORE_DATAPATH__0key_host_1__31_0__9_;
  wire AES_CORE_DATAPATH__0key_host_2__31_0__0_;
  wire AES_CORE_DATAPATH__0key_host_2__31_0__10_;
  wire AES_CORE_DATAPATH__0key_host_2__31_0__11_;
  wire AES_CORE_DATAPATH__0key_host_2__31_0__12_;
  wire AES_CORE_DATAPATH__0key_host_2__31_0__13_;
  wire AES_CORE_DATAPATH__0key_host_2__31_0__14_;
  wire AES_CORE_DATAPATH__0key_host_2__31_0__15_;
  wire AES_CORE_DATAPATH__0key_host_2__31_0__16_;
  wire AES_CORE_DATAPATH__0key_host_2__31_0__17_;
  wire AES_CORE_DATAPATH__0key_host_2__31_0__18_;
  wire AES_CORE_DATAPATH__0key_host_2__31_0__19_;
  wire AES_CORE_DATAPATH__0key_host_2__31_0__1_;
  wire AES_CORE_DATAPATH__0key_host_2__31_0__20_;
  wire AES_CORE_DATAPATH__0key_host_2__31_0__21_;
  wire AES_CORE_DATAPATH__0key_host_2__31_0__22_;
  wire AES_CORE_DATAPATH__0key_host_2__31_0__23_;
  wire AES_CORE_DATAPATH__0key_host_2__31_0__24_;
  wire AES_CORE_DATAPATH__0key_host_2__31_0__25_;
  wire AES_CORE_DATAPATH__0key_host_2__31_0__26_;
  wire AES_CORE_DATAPATH__0key_host_2__31_0__27_;
  wire AES_CORE_DATAPATH__0key_host_2__31_0__28_;
  wire AES_CORE_DATAPATH__0key_host_2__31_0__29_;
  wire AES_CORE_DATAPATH__0key_host_2__31_0__2_;
  wire AES_CORE_DATAPATH__0key_host_2__31_0__30_;
  wire AES_CORE_DATAPATH__0key_host_2__31_0__31_;
  wire AES_CORE_DATAPATH__0key_host_2__31_0__3_;
  wire AES_CORE_DATAPATH__0key_host_2__31_0__4_;
  wire AES_CORE_DATAPATH__0key_host_2__31_0__5_;
  wire AES_CORE_DATAPATH__0key_host_2__31_0__6_;
  wire AES_CORE_DATAPATH__0key_host_2__31_0__7_;
  wire AES_CORE_DATAPATH__0key_host_2__31_0__8_;
  wire AES_CORE_DATAPATH__0key_host_2__31_0__9_;
  wire AES_CORE_DATAPATH__0key_host_3__31_0__0_;
  wire AES_CORE_DATAPATH__0key_host_3__31_0__10_;
  wire AES_CORE_DATAPATH__0key_host_3__31_0__11_;
  wire AES_CORE_DATAPATH__0key_host_3__31_0__12_;
  wire AES_CORE_DATAPATH__0key_host_3__31_0__13_;
  wire AES_CORE_DATAPATH__0key_host_3__31_0__14_;
  wire AES_CORE_DATAPATH__0key_host_3__31_0__15_;
  wire AES_CORE_DATAPATH__0key_host_3__31_0__16_;
  wire AES_CORE_DATAPATH__0key_host_3__31_0__17_;
  wire AES_CORE_DATAPATH__0key_host_3__31_0__18_;
  wire AES_CORE_DATAPATH__0key_host_3__31_0__19_;
  wire AES_CORE_DATAPATH__0key_host_3__31_0__1_;
  wire AES_CORE_DATAPATH__0key_host_3__31_0__20_;
  wire AES_CORE_DATAPATH__0key_host_3__31_0__21_;
  wire AES_CORE_DATAPATH__0key_host_3__31_0__22_;
  wire AES_CORE_DATAPATH__0key_host_3__31_0__23_;
  wire AES_CORE_DATAPATH__0key_host_3__31_0__24_;
  wire AES_CORE_DATAPATH__0key_host_3__31_0__25_;
  wire AES_CORE_DATAPATH__0key_host_3__31_0__26_;
  wire AES_CORE_DATAPATH__0key_host_3__31_0__27_;
  wire AES_CORE_DATAPATH__0key_host_3__31_0__28_;
  wire AES_CORE_DATAPATH__0key_host_3__31_0__29_;
  wire AES_CORE_DATAPATH__0key_host_3__31_0__2_;
  wire AES_CORE_DATAPATH__0key_host_3__31_0__30_;
  wire AES_CORE_DATAPATH__0key_host_3__31_0__31_;
  wire AES_CORE_DATAPATH__0key_host_3__31_0__3_;
  wire AES_CORE_DATAPATH__0key_host_3__31_0__4_;
  wire AES_CORE_DATAPATH__0key_host_3__31_0__5_;
  wire AES_CORE_DATAPATH__0key_host_3__31_0__6_;
  wire AES_CORE_DATAPATH__0key_host_3__31_0__7_;
  wire AES_CORE_DATAPATH__0key_host_3__31_0__8_;
  wire AES_CORE_DATAPATH__0key_host_3__31_0__9_;
  wire AES_CORE_DATAPATH__abc_16259_n10000;
  wire AES_CORE_DATAPATH__abc_16259_n10001;
  wire AES_CORE_DATAPATH__abc_16259_n10002;
  wire AES_CORE_DATAPATH__abc_16259_n10003;
  wire AES_CORE_DATAPATH__abc_16259_n10005;
  wire AES_CORE_DATAPATH__abc_16259_n10006;
  wire AES_CORE_DATAPATH__abc_16259_n10007;
  wire AES_CORE_DATAPATH__abc_16259_n10008;
  wire AES_CORE_DATAPATH__abc_16259_n10009;
  wire AES_CORE_DATAPATH__abc_16259_n10010;
  wire AES_CORE_DATAPATH__abc_16259_n10011;
  wire AES_CORE_DATAPATH__abc_16259_n10013;
  wire AES_CORE_DATAPATH__abc_16259_n10014;
  wire AES_CORE_DATAPATH__abc_16259_n10015;
  wire AES_CORE_DATAPATH__abc_16259_n10016;
  wire AES_CORE_DATAPATH__abc_16259_n10017;
  wire AES_CORE_DATAPATH__abc_16259_n10018;
  wire AES_CORE_DATAPATH__abc_16259_n10019;
  wire AES_CORE_DATAPATH__abc_16259_n10021;
  wire AES_CORE_DATAPATH__abc_16259_n10022;
  wire AES_CORE_DATAPATH__abc_16259_n10023;
  wire AES_CORE_DATAPATH__abc_16259_n10024;
  wire AES_CORE_DATAPATH__abc_16259_n10025;
  wire AES_CORE_DATAPATH__abc_16259_n10026;
  wire AES_CORE_DATAPATH__abc_16259_n10027;
  wire AES_CORE_DATAPATH__abc_16259_n10029;
  wire AES_CORE_DATAPATH__abc_16259_n10030;
  wire AES_CORE_DATAPATH__abc_16259_n10031;
  wire AES_CORE_DATAPATH__abc_16259_n10032;
  wire AES_CORE_DATAPATH__abc_16259_n10033;
  wire AES_CORE_DATAPATH__abc_16259_n10034;
  wire AES_CORE_DATAPATH__abc_16259_n10035;
  wire AES_CORE_DATAPATH__abc_16259_n10036;
  wire AES_CORE_DATAPATH__abc_16259_n10038;
  wire AES_CORE_DATAPATH__abc_16259_n10039;
  wire AES_CORE_DATAPATH__abc_16259_n10040;
  wire AES_CORE_DATAPATH__abc_16259_n10041;
  wire AES_CORE_DATAPATH__abc_16259_n10042;
  wire AES_CORE_DATAPATH__abc_16259_n10043;
  wire AES_CORE_DATAPATH__abc_16259_n10044;
  wire AES_CORE_DATAPATH__abc_16259_n10046;
  wire AES_CORE_DATAPATH__abc_16259_n10047;
  wire AES_CORE_DATAPATH__abc_16259_n10048;
  wire AES_CORE_DATAPATH__abc_16259_n10049;
  wire AES_CORE_DATAPATH__abc_16259_n10050;
  wire AES_CORE_DATAPATH__abc_16259_n10051;
  wire AES_CORE_DATAPATH__abc_16259_n10052;
  wire AES_CORE_DATAPATH__abc_16259_n10054;
  wire AES_CORE_DATAPATH__abc_16259_n10055;
  wire AES_CORE_DATAPATH__abc_16259_n10056;
  wire AES_CORE_DATAPATH__abc_16259_n10057;
  wire AES_CORE_DATAPATH__abc_16259_n10058;
  wire AES_CORE_DATAPATH__abc_16259_n10059;
  wire AES_CORE_DATAPATH__abc_16259_n10060;
  wire AES_CORE_DATAPATH__abc_16259_n10062;
  wire AES_CORE_DATAPATH__abc_16259_n10063;
  wire AES_CORE_DATAPATH__abc_16259_n10064;
  wire AES_CORE_DATAPATH__abc_16259_n10065;
  wire AES_CORE_DATAPATH__abc_16259_n10066;
  wire AES_CORE_DATAPATH__abc_16259_n10067;
  wire AES_CORE_DATAPATH__abc_16259_n10068;
  wire AES_CORE_DATAPATH__abc_16259_n10070;
  wire AES_CORE_DATAPATH__abc_16259_n10071;
  wire AES_CORE_DATAPATH__abc_16259_n10072;
  wire AES_CORE_DATAPATH__abc_16259_n10073;
  wire AES_CORE_DATAPATH__abc_16259_n10074;
  wire AES_CORE_DATAPATH__abc_16259_n10075;
  wire AES_CORE_DATAPATH__abc_16259_n10076;
  wire AES_CORE_DATAPATH__abc_16259_n10078;
  wire AES_CORE_DATAPATH__abc_16259_n10079;
  wire AES_CORE_DATAPATH__abc_16259_n10080;
  wire AES_CORE_DATAPATH__abc_16259_n10081;
  wire AES_CORE_DATAPATH__abc_16259_n10082;
  wire AES_CORE_DATAPATH__abc_16259_n10083;
  wire AES_CORE_DATAPATH__abc_16259_n10084;
  wire AES_CORE_DATAPATH__abc_16259_n10086;
  wire AES_CORE_DATAPATH__abc_16259_n10087;
  wire AES_CORE_DATAPATH__abc_16259_n10088;
  wire AES_CORE_DATAPATH__abc_16259_n10089;
  wire AES_CORE_DATAPATH__abc_16259_n10090;
  wire AES_CORE_DATAPATH__abc_16259_n10091;
  wire AES_CORE_DATAPATH__abc_16259_n10092;
  wire AES_CORE_DATAPATH__abc_16259_n10094;
  wire AES_CORE_DATAPATH__abc_16259_n10095;
  wire AES_CORE_DATAPATH__abc_16259_n10096;
  wire AES_CORE_DATAPATH__abc_16259_n10097;
  wire AES_CORE_DATAPATH__abc_16259_n10098;
  wire AES_CORE_DATAPATH__abc_16259_n10099;
  wire AES_CORE_DATAPATH__abc_16259_n10100;
  wire AES_CORE_DATAPATH__abc_16259_n10102;
  wire AES_CORE_DATAPATH__abc_16259_n10103;
  wire AES_CORE_DATAPATH__abc_16259_n10104;
  wire AES_CORE_DATAPATH__abc_16259_n10105;
  wire AES_CORE_DATAPATH__abc_16259_n10106;
  wire AES_CORE_DATAPATH__abc_16259_n10107;
  wire AES_CORE_DATAPATH__abc_16259_n10108;
  wire AES_CORE_DATAPATH__abc_16259_n10110;
  wire AES_CORE_DATAPATH__abc_16259_n10111;
  wire AES_CORE_DATAPATH__abc_16259_n10112;
  wire AES_CORE_DATAPATH__abc_16259_n10113;
  wire AES_CORE_DATAPATH__abc_16259_n10114;
  wire AES_CORE_DATAPATH__abc_16259_n10115;
  wire AES_CORE_DATAPATH__abc_16259_n10116;
  wire AES_CORE_DATAPATH__abc_16259_n10118;
  wire AES_CORE_DATAPATH__abc_16259_n10119;
  wire AES_CORE_DATAPATH__abc_16259_n10119_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n10119_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n10119_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n10119_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n10119_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n10120;
  wire AES_CORE_DATAPATH__abc_16259_n10122;
  wire AES_CORE_DATAPATH__abc_16259_n10123;
  wire AES_CORE_DATAPATH__abc_16259_n10125;
  wire AES_CORE_DATAPATH__abc_16259_n10126;
  wire AES_CORE_DATAPATH__abc_16259_n10128;
  wire AES_CORE_DATAPATH__abc_16259_n10129;
  wire AES_CORE_DATAPATH__abc_16259_n10131;
  wire AES_CORE_DATAPATH__abc_16259_n10132;
  wire AES_CORE_DATAPATH__abc_16259_n10134;
  wire AES_CORE_DATAPATH__abc_16259_n10135;
  wire AES_CORE_DATAPATH__abc_16259_n10137;
  wire AES_CORE_DATAPATH__abc_16259_n10138;
  wire AES_CORE_DATAPATH__abc_16259_n10140;
  wire AES_CORE_DATAPATH__abc_16259_n10141;
  wire AES_CORE_DATAPATH__abc_16259_n10143;
  wire AES_CORE_DATAPATH__abc_16259_n10144;
  wire AES_CORE_DATAPATH__abc_16259_n10146;
  wire AES_CORE_DATAPATH__abc_16259_n10147;
  wire AES_CORE_DATAPATH__abc_16259_n10149;
  wire AES_CORE_DATAPATH__abc_16259_n10150;
  wire AES_CORE_DATAPATH__abc_16259_n10152;
  wire AES_CORE_DATAPATH__abc_16259_n10153;
  wire AES_CORE_DATAPATH__abc_16259_n10155;
  wire AES_CORE_DATAPATH__abc_16259_n10156;
  wire AES_CORE_DATAPATH__abc_16259_n10158;
  wire AES_CORE_DATAPATH__abc_16259_n10159;
  wire AES_CORE_DATAPATH__abc_16259_n10161;
  wire AES_CORE_DATAPATH__abc_16259_n10162;
  wire AES_CORE_DATAPATH__abc_16259_n10164;
  wire AES_CORE_DATAPATH__abc_16259_n10165;
  wire AES_CORE_DATAPATH__abc_16259_n10167;
  wire AES_CORE_DATAPATH__abc_16259_n10168;
  wire AES_CORE_DATAPATH__abc_16259_n10170;
  wire AES_CORE_DATAPATH__abc_16259_n10171;
  wire AES_CORE_DATAPATH__abc_16259_n10173;
  wire AES_CORE_DATAPATH__abc_16259_n10174;
  wire AES_CORE_DATAPATH__abc_16259_n10176;
  wire AES_CORE_DATAPATH__abc_16259_n10177;
  wire AES_CORE_DATAPATH__abc_16259_n10179;
  wire AES_CORE_DATAPATH__abc_16259_n10180;
  wire AES_CORE_DATAPATH__abc_16259_n10182;
  wire AES_CORE_DATAPATH__abc_16259_n10183;
  wire AES_CORE_DATAPATH__abc_16259_n10185;
  wire AES_CORE_DATAPATH__abc_16259_n10186;
  wire AES_CORE_DATAPATH__abc_16259_n10188;
  wire AES_CORE_DATAPATH__abc_16259_n10189;
  wire AES_CORE_DATAPATH__abc_16259_n10191;
  wire AES_CORE_DATAPATH__abc_16259_n10192;
  wire AES_CORE_DATAPATH__abc_16259_n10194;
  wire AES_CORE_DATAPATH__abc_16259_n10195;
  wire AES_CORE_DATAPATH__abc_16259_n10197;
  wire AES_CORE_DATAPATH__abc_16259_n10198;
  wire AES_CORE_DATAPATH__abc_16259_n10200;
  wire AES_CORE_DATAPATH__abc_16259_n10201;
  wire AES_CORE_DATAPATH__abc_16259_n10203;
  wire AES_CORE_DATAPATH__abc_16259_n10204;
  wire AES_CORE_DATAPATH__abc_16259_n10206;
  wire AES_CORE_DATAPATH__abc_16259_n10207;
  wire AES_CORE_DATAPATH__abc_16259_n10209;
  wire AES_CORE_DATAPATH__abc_16259_n10210;
  wire AES_CORE_DATAPATH__abc_16259_n10212;
  wire AES_CORE_DATAPATH__abc_16259_n10213;
  wire AES_CORE_DATAPATH__abc_16259_n10215;
  wire AES_CORE_DATAPATH__abc_16259_n10216;
  wire AES_CORE_DATAPATH__abc_16259_n10217;
  wire AES_CORE_DATAPATH__abc_16259_n10217_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n10217_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n10217_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n10217_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n10217_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n10217_bF_buf5;
  wire AES_CORE_DATAPATH__abc_16259_n10217_bF_buf6;
  wire AES_CORE_DATAPATH__abc_16259_n10217_bF_buf7;
  wire AES_CORE_DATAPATH__abc_16259_n10218;
  wire AES_CORE_DATAPATH__abc_16259_n10218_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n10218_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n10218_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n10218_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n10218_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n10218_bF_buf5;
  wire AES_CORE_DATAPATH__abc_16259_n10218_bF_buf6;
  wire AES_CORE_DATAPATH__abc_16259_n10219;
  wire AES_CORE_DATAPATH__abc_16259_n10220;
  wire AES_CORE_DATAPATH__abc_16259_n10222;
  wire AES_CORE_DATAPATH__abc_16259_n10223;
  wire AES_CORE_DATAPATH__abc_16259_n10225;
  wire AES_CORE_DATAPATH__abc_16259_n10226;
  wire AES_CORE_DATAPATH__abc_16259_n10228;
  wire AES_CORE_DATAPATH__abc_16259_n10229;
  wire AES_CORE_DATAPATH__abc_16259_n10231;
  wire AES_CORE_DATAPATH__abc_16259_n10232;
  wire AES_CORE_DATAPATH__abc_16259_n10234;
  wire AES_CORE_DATAPATH__abc_16259_n10235;
  wire AES_CORE_DATAPATH__abc_16259_n10237;
  wire AES_CORE_DATAPATH__abc_16259_n10238;
  wire AES_CORE_DATAPATH__abc_16259_n10240;
  wire AES_CORE_DATAPATH__abc_16259_n10241;
  wire AES_CORE_DATAPATH__abc_16259_n10243;
  wire AES_CORE_DATAPATH__abc_16259_n10244;
  wire AES_CORE_DATAPATH__abc_16259_n10246;
  wire AES_CORE_DATAPATH__abc_16259_n10247;
  wire AES_CORE_DATAPATH__abc_16259_n10249;
  wire AES_CORE_DATAPATH__abc_16259_n10250;
  wire AES_CORE_DATAPATH__abc_16259_n10251;
  wire AES_CORE_DATAPATH__abc_16259_n10253;
  wire AES_CORE_DATAPATH__abc_16259_n10254;
  wire AES_CORE_DATAPATH__abc_16259_n10255;
  wire AES_CORE_DATAPATH__abc_16259_n10257;
  wire AES_CORE_DATAPATH__abc_16259_n10258;
  wire AES_CORE_DATAPATH__abc_16259_n10260;
  wire AES_CORE_DATAPATH__abc_16259_n10261;
  wire AES_CORE_DATAPATH__abc_16259_n10262;
  wire AES_CORE_DATAPATH__abc_16259_n10264;
  wire AES_CORE_DATAPATH__abc_16259_n10265;
  wire AES_CORE_DATAPATH__abc_16259_n10267;
  wire AES_CORE_DATAPATH__abc_16259_n10268;
  wire AES_CORE_DATAPATH__abc_16259_n10269;
  wire AES_CORE_DATAPATH__abc_16259_n10271;
  wire AES_CORE_DATAPATH__abc_16259_n10272;
  wire AES_CORE_DATAPATH__abc_16259_n10274;
  wire AES_CORE_DATAPATH__abc_16259_n10275;
  wire AES_CORE_DATAPATH__abc_16259_n10276;
  wire AES_CORE_DATAPATH__abc_16259_n10278;
  wire AES_CORE_DATAPATH__abc_16259_n10279;
  wire AES_CORE_DATAPATH__abc_16259_n10281;
  wire AES_CORE_DATAPATH__abc_16259_n10282;
  wire AES_CORE_DATAPATH__abc_16259_n10284;
  wire AES_CORE_DATAPATH__abc_16259_n10285;
  wire AES_CORE_DATAPATH__abc_16259_n10287;
  wire AES_CORE_DATAPATH__abc_16259_n10288;
  wire AES_CORE_DATAPATH__abc_16259_n10289;
  wire AES_CORE_DATAPATH__abc_16259_n10291;
  wire AES_CORE_DATAPATH__abc_16259_n10292;
  wire AES_CORE_DATAPATH__abc_16259_n10294;
  wire AES_CORE_DATAPATH__abc_16259_n10295;
  wire AES_CORE_DATAPATH__abc_16259_n10297;
  wire AES_CORE_DATAPATH__abc_16259_n10298;
  wire AES_CORE_DATAPATH__abc_16259_n10300;
  wire AES_CORE_DATAPATH__abc_16259_n10301;
  wire AES_CORE_DATAPATH__abc_16259_n10303;
  wire AES_CORE_DATAPATH__abc_16259_n10304;
  wire AES_CORE_DATAPATH__abc_16259_n10306;
  wire AES_CORE_DATAPATH__abc_16259_n10307;
  wire AES_CORE_DATAPATH__abc_16259_n10309;
  wire AES_CORE_DATAPATH__abc_16259_n10310;
  wire AES_CORE_DATAPATH__abc_16259_n10312;
  wire AES_CORE_DATAPATH__abc_16259_n10313;
  wire AES_CORE_DATAPATH__abc_16259_n10315;
  wire AES_CORE_DATAPATH__abc_16259_n10316;
  wire AES_CORE_DATAPATH__abc_16259_n10318;
  wire AES_CORE_DATAPATH__abc_16259_n10319;
  wire AES_CORE_DATAPATH__abc_16259_n10321;
  wire AES_CORE_DATAPATH__abc_16259_n10322;
  wire AES_CORE_DATAPATH__abc_16259_n10323;
  wire AES_CORE_DATAPATH__abc_16259_n10324;
  wire AES_CORE_DATAPATH__abc_16259_n10325;
  wire AES_CORE_DATAPATH__abc_16259_n10326;
  wire AES_CORE_DATAPATH__abc_16259_n10327;
  wire AES_CORE_DATAPATH__abc_16259_n10329;
  wire AES_CORE_DATAPATH__abc_16259_n10330;
  wire AES_CORE_DATAPATH__abc_16259_n10331;
  wire AES_CORE_DATAPATH__abc_16259_n10332;
  wire AES_CORE_DATAPATH__abc_16259_n10333;
  wire AES_CORE_DATAPATH__abc_16259_n10334;
  wire AES_CORE_DATAPATH__abc_16259_n10335;
  wire AES_CORE_DATAPATH__abc_16259_n10337;
  wire AES_CORE_DATAPATH__abc_16259_n10338;
  wire AES_CORE_DATAPATH__abc_16259_n10339;
  wire AES_CORE_DATAPATH__abc_16259_n10340;
  wire AES_CORE_DATAPATH__abc_16259_n10341;
  wire AES_CORE_DATAPATH__abc_16259_n10342;
  wire AES_CORE_DATAPATH__abc_16259_n10343;
  wire AES_CORE_DATAPATH__abc_16259_n10345;
  wire AES_CORE_DATAPATH__abc_16259_n10346;
  wire AES_CORE_DATAPATH__abc_16259_n10347;
  wire AES_CORE_DATAPATH__abc_16259_n10348;
  wire AES_CORE_DATAPATH__abc_16259_n10349;
  wire AES_CORE_DATAPATH__abc_16259_n10350;
  wire AES_CORE_DATAPATH__abc_16259_n10351;
  wire AES_CORE_DATAPATH__abc_16259_n10353;
  wire AES_CORE_DATAPATH__abc_16259_n10354;
  wire AES_CORE_DATAPATH__abc_16259_n10355;
  wire AES_CORE_DATAPATH__abc_16259_n10356;
  wire AES_CORE_DATAPATH__abc_16259_n10357;
  wire AES_CORE_DATAPATH__abc_16259_n10358;
  wire AES_CORE_DATAPATH__abc_16259_n10359;
  wire AES_CORE_DATAPATH__abc_16259_n10361;
  wire AES_CORE_DATAPATH__abc_16259_n10362;
  wire AES_CORE_DATAPATH__abc_16259_n10363;
  wire AES_CORE_DATAPATH__abc_16259_n10364;
  wire AES_CORE_DATAPATH__abc_16259_n10365;
  wire AES_CORE_DATAPATH__abc_16259_n10366;
  wire AES_CORE_DATAPATH__abc_16259_n10367;
  wire AES_CORE_DATAPATH__abc_16259_n10369;
  wire AES_CORE_DATAPATH__abc_16259_n10370;
  wire AES_CORE_DATAPATH__abc_16259_n10371;
  wire AES_CORE_DATAPATH__abc_16259_n10372;
  wire AES_CORE_DATAPATH__abc_16259_n10373;
  wire AES_CORE_DATAPATH__abc_16259_n10374;
  wire AES_CORE_DATAPATH__abc_16259_n10375;
  wire AES_CORE_DATAPATH__abc_16259_n10377;
  wire AES_CORE_DATAPATH__abc_16259_n10378;
  wire AES_CORE_DATAPATH__abc_16259_n10379;
  wire AES_CORE_DATAPATH__abc_16259_n10380;
  wire AES_CORE_DATAPATH__abc_16259_n10381;
  wire AES_CORE_DATAPATH__abc_16259_n10382;
  wire AES_CORE_DATAPATH__abc_16259_n10383;
  wire AES_CORE_DATAPATH__abc_16259_n10385;
  wire AES_CORE_DATAPATH__abc_16259_n10386;
  wire AES_CORE_DATAPATH__abc_16259_n10387;
  wire AES_CORE_DATAPATH__abc_16259_n10388;
  wire AES_CORE_DATAPATH__abc_16259_n10389;
  wire AES_CORE_DATAPATH__abc_16259_n10390;
  wire AES_CORE_DATAPATH__abc_16259_n10391;
  wire AES_CORE_DATAPATH__abc_16259_n10393;
  wire AES_CORE_DATAPATH__abc_16259_n10394;
  wire AES_CORE_DATAPATH__abc_16259_n10395;
  wire AES_CORE_DATAPATH__abc_16259_n10396;
  wire AES_CORE_DATAPATH__abc_16259_n10397;
  wire AES_CORE_DATAPATH__abc_16259_n10398;
  wire AES_CORE_DATAPATH__abc_16259_n10399;
  wire AES_CORE_DATAPATH__abc_16259_n10401;
  wire AES_CORE_DATAPATH__abc_16259_n10402;
  wire AES_CORE_DATAPATH__abc_16259_n10403;
  wire AES_CORE_DATAPATH__abc_16259_n10404;
  wire AES_CORE_DATAPATH__abc_16259_n10405;
  wire AES_CORE_DATAPATH__abc_16259_n10406;
  wire AES_CORE_DATAPATH__abc_16259_n10407;
  wire AES_CORE_DATAPATH__abc_16259_n10408;
  wire AES_CORE_DATAPATH__abc_16259_n10410;
  wire AES_CORE_DATAPATH__abc_16259_n10411;
  wire AES_CORE_DATAPATH__abc_16259_n10412;
  wire AES_CORE_DATAPATH__abc_16259_n10413;
  wire AES_CORE_DATAPATH__abc_16259_n10414;
  wire AES_CORE_DATAPATH__abc_16259_n10415;
  wire AES_CORE_DATAPATH__abc_16259_n10416;
  wire AES_CORE_DATAPATH__abc_16259_n10417;
  wire AES_CORE_DATAPATH__abc_16259_n10419;
  wire AES_CORE_DATAPATH__abc_16259_n10420;
  wire AES_CORE_DATAPATH__abc_16259_n10421;
  wire AES_CORE_DATAPATH__abc_16259_n10422;
  wire AES_CORE_DATAPATH__abc_16259_n10423;
  wire AES_CORE_DATAPATH__abc_16259_n10424;
  wire AES_CORE_DATAPATH__abc_16259_n10425;
  wire AES_CORE_DATAPATH__abc_16259_n10427;
  wire AES_CORE_DATAPATH__abc_16259_n10428;
  wire AES_CORE_DATAPATH__abc_16259_n10429;
  wire AES_CORE_DATAPATH__abc_16259_n10430;
  wire AES_CORE_DATAPATH__abc_16259_n10431;
  wire AES_CORE_DATAPATH__abc_16259_n10432;
  wire AES_CORE_DATAPATH__abc_16259_n10433;
  wire AES_CORE_DATAPATH__abc_16259_n10434;
  wire AES_CORE_DATAPATH__abc_16259_n10436;
  wire AES_CORE_DATAPATH__abc_16259_n10437;
  wire AES_CORE_DATAPATH__abc_16259_n10438;
  wire AES_CORE_DATAPATH__abc_16259_n10439;
  wire AES_CORE_DATAPATH__abc_16259_n10440;
  wire AES_CORE_DATAPATH__abc_16259_n10441;
  wire AES_CORE_DATAPATH__abc_16259_n10442;
  wire AES_CORE_DATAPATH__abc_16259_n10444;
  wire AES_CORE_DATAPATH__abc_16259_n10445;
  wire AES_CORE_DATAPATH__abc_16259_n10446;
  wire AES_CORE_DATAPATH__abc_16259_n10447;
  wire AES_CORE_DATAPATH__abc_16259_n10448;
  wire AES_CORE_DATAPATH__abc_16259_n10449;
  wire AES_CORE_DATAPATH__abc_16259_n10450;
  wire AES_CORE_DATAPATH__abc_16259_n10451;
  wire AES_CORE_DATAPATH__abc_16259_n10453;
  wire AES_CORE_DATAPATH__abc_16259_n10454;
  wire AES_CORE_DATAPATH__abc_16259_n10455;
  wire AES_CORE_DATAPATH__abc_16259_n10456;
  wire AES_CORE_DATAPATH__abc_16259_n10457;
  wire AES_CORE_DATAPATH__abc_16259_n10458;
  wire AES_CORE_DATAPATH__abc_16259_n10459;
  wire AES_CORE_DATAPATH__abc_16259_n10461;
  wire AES_CORE_DATAPATH__abc_16259_n10462;
  wire AES_CORE_DATAPATH__abc_16259_n10463;
  wire AES_CORE_DATAPATH__abc_16259_n10464;
  wire AES_CORE_DATAPATH__abc_16259_n10465;
  wire AES_CORE_DATAPATH__abc_16259_n10466;
  wire AES_CORE_DATAPATH__abc_16259_n10467;
  wire AES_CORE_DATAPATH__abc_16259_n10468;
  wire AES_CORE_DATAPATH__abc_16259_n10470;
  wire AES_CORE_DATAPATH__abc_16259_n10471;
  wire AES_CORE_DATAPATH__abc_16259_n10472;
  wire AES_CORE_DATAPATH__abc_16259_n10473;
  wire AES_CORE_DATAPATH__abc_16259_n10474;
  wire AES_CORE_DATAPATH__abc_16259_n10475;
  wire AES_CORE_DATAPATH__abc_16259_n10476;
  wire AES_CORE_DATAPATH__abc_16259_n10478;
  wire AES_CORE_DATAPATH__abc_16259_n10479;
  wire AES_CORE_DATAPATH__abc_16259_n10480;
  wire AES_CORE_DATAPATH__abc_16259_n10481;
  wire AES_CORE_DATAPATH__abc_16259_n10482;
  wire AES_CORE_DATAPATH__abc_16259_n10483;
  wire AES_CORE_DATAPATH__abc_16259_n10484;
  wire AES_CORE_DATAPATH__abc_16259_n10486;
  wire AES_CORE_DATAPATH__abc_16259_n10487;
  wire AES_CORE_DATAPATH__abc_16259_n10488;
  wire AES_CORE_DATAPATH__abc_16259_n10489;
  wire AES_CORE_DATAPATH__abc_16259_n10490;
  wire AES_CORE_DATAPATH__abc_16259_n10491;
  wire AES_CORE_DATAPATH__abc_16259_n10492;
  wire AES_CORE_DATAPATH__abc_16259_n10494;
  wire AES_CORE_DATAPATH__abc_16259_n10495;
  wire AES_CORE_DATAPATH__abc_16259_n10496;
  wire AES_CORE_DATAPATH__abc_16259_n10497;
  wire AES_CORE_DATAPATH__abc_16259_n10498;
  wire AES_CORE_DATAPATH__abc_16259_n10499;
  wire AES_CORE_DATAPATH__abc_16259_n10500;
  wire AES_CORE_DATAPATH__abc_16259_n10501;
  wire AES_CORE_DATAPATH__abc_16259_n10503;
  wire AES_CORE_DATAPATH__abc_16259_n10504;
  wire AES_CORE_DATAPATH__abc_16259_n10505;
  wire AES_CORE_DATAPATH__abc_16259_n10506;
  wire AES_CORE_DATAPATH__abc_16259_n10507;
  wire AES_CORE_DATAPATH__abc_16259_n10508;
  wire AES_CORE_DATAPATH__abc_16259_n10509;
  wire AES_CORE_DATAPATH__abc_16259_n10511;
  wire AES_CORE_DATAPATH__abc_16259_n10512;
  wire AES_CORE_DATAPATH__abc_16259_n10513;
  wire AES_CORE_DATAPATH__abc_16259_n10514;
  wire AES_CORE_DATAPATH__abc_16259_n10515;
  wire AES_CORE_DATAPATH__abc_16259_n10516;
  wire AES_CORE_DATAPATH__abc_16259_n10517;
  wire AES_CORE_DATAPATH__abc_16259_n10519;
  wire AES_CORE_DATAPATH__abc_16259_n10520;
  wire AES_CORE_DATAPATH__abc_16259_n10521;
  wire AES_CORE_DATAPATH__abc_16259_n10522;
  wire AES_CORE_DATAPATH__abc_16259_n10523;
  wire AES_CORE_DATAPATH__abc_16259_n10524;
  wire AES_CORE_DATAPATH__abc_16259_n10525;
  wire AES_CORE_DATAPATH__abc_16259_n10527;
  wire AES_CORE_DATAPATH__abc_16259_n10528;
  wire AES_CORE_DATAPATH__abc_16259_n10529;
  wire AES_CORE_DATAPATH__abc_16259_n10530;
  wire AES_CORE_DATAPATH__abc_16259_n10531;
  wire AES_CORE_DATAPATH__abc_16259_n10532;
  wire AES_CORE_DATAPATH__abc_16259_n10533;
  wire AES_CORE_DATAPATH__abc_16259_n10535;
  wire AES_CORE_DATAPATH__abc_16259_n10536;
  wire AES_CORE_DATAPATH__abc_16259_n10537;
  wire AES_CORE_DATAPATH__abc_16259_n10538;
  wire AES_CORE_DATAPATH__abc_16259_n10539;
  wire AES_CORE_DATAPATH__abc_16259_n10540;
  wire AES_CORE_DATAPATH__abc_16259_n10541;
  wire AES_CORE_DATAPATH__abc_16259_n10543;
  wire AES_CORE_DATAPATH__abc_16259_n10544;
  wire AES_CORE_DATAPATH__abc_16259_n10545;
  wire AES_CORE_DATAPATH__abc_16259_n10546;
  wire AES_CORE_DATAPATH__abc_16259_n10547;
  wire AES_CORE_DATAPATH__abc_16259_n10548;
  wire AES_CORE_DATAPATH__abc_16259_n10549;
  wire AES_CORE_DATAPATH__abc_16259_n10551;
  wire AES_CORE_DATAPATH__abc_16259_n10552;
  wire AES_CORE_DATAPATH__abc_16259_n10553;
  wire AES_CORE_DATAPATH__abc_16259_n10554;
  wire AES_CORE_DATAPATH__abc_16259_n10555;
  wire AES_CORE_DATAPATH__abc_16259_n10556;
  wire AES_CORE_DATAPATH__abc_16259_n10557;
  wire AES_CORE_DATAPATH__abc_16259_n10559;
  wire AES_CORE_DATAPATH__abc_16259_n10560;
  wire AES_CORE_DATAPATH__abc_16259_n10561;
  wire AES_CORE_DATAPATH__abc_16259_n10562;
  wire AES_CORE_DATAPATH__abc_16259_n10563;
  wire AES_CORE_DATAPATH__abc_16259_n10564;
  wire AES_CORE_DATAPATH__abc_16259_n10565;
  wire AES_CORE_DATAPATH__abc_16259_n10567;
  wire AES_CORE_DATAPATH__abc_16259_n10568;
  wire AES_CORE_DATAPATH__abc_16259_n10569;
  wire AES_CORE_DATAPATH__abc_16259_n10570;
  wire AES_CORE_DATAPATH__abc_16259_n10571;
  wire AES_CORE_DATAPATH__abc_16259_n10572;
  wire AES_CORE_DATAPATH__abc_16259_n10573;
  wire AES_CORE_DATAPATH__abc_16259_n10575;
  wire AES_CORE_DATAPATH__abc_16259_n10576;
  wire AES_CORE_DATAPATH__abc_16259_n10577;
  wire AES_CORE_DATAPATH__abc_16259_n10578;
  wire AES_CORE_DATAPATH__abc_16259_n10579;
  wire AES_CORE_DATAPATH__abc_16259_n10580;
  wire AES_CORE_DATAPATH__abc_16259_n10581;
  wire AES_CORE_DATAPATH__abc_16259_n10583;
  wire AES_CORE_DATAPATH__abc_16259_n10584;
  wire AES_CORE_DATAPATH__abc_16259_n10584_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n10584_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n10584_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n10584_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n10584_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n10585;
  wire AES_CORE_DATAPATH__abc_16259_n10587;
  wire AES_CORE_DATAPATH__abc_16259_n10588;
  wire AES_CORE_DATAPATH__abc_16259_n10590;
  wire AES_CORE_DATAPATH__abc_16259_n10591;
  wire AES_CORE_DATAPATH__abc_16259_n10593;
  wire AES_CORE_DATAPATH__abc_16259_n10594;
  wire AES_CORE_DATAPATH__abc_16259_n10596;
  wire AES_CORE_DATAPATH__abc_16259_n10597;
  wire AES_CORE_DATAPATH__abc_16259_n10599;
  wire AES_CORE_DATAPATH__abc_16259_n10600;
  wire AES_CORE_DATAPATH__abc_16259_n10602;
  wire AES_CORE_DATAPATH__abc_16259_n10603;
  wire AES_CORE_DATAPATH__abc_16259_n10605;
  wire AES_CORE_DATAPATH__abc_16259_n10606;
  wire AES_CORE_DATAPATH__abc_16259_n10608;
  wire AES_CORE_DATAPATH__abc_16259_n10609;
  wire AES_CORE_DATAPATH__abc_16259_n10611;
  wire AES_CORE_DATAPATH__abc_16259_n10612;
  wire AES_CORE_DATAPATH__abc_16259_n10614;
  wire AES_CORE_DATAPATH__abc_16259_n10615;
  wire AES_CORE_DATAPATH__abc_16259_n10617;
  wire AES_CORE_DATAPATH__abc_16259_n10618;
  wire AES_CORE_DATAPATH__abc_16259_n10620;
  wire AES_CORE_DATAPATH__abc_16259_n10621;
  wire AES_CORE_DATAPATH__abc_16259_n10623;
  wire AES_CORE_DATAPATH__abc_16259_n10624;
  wire AES_CORE_DATAPATH__abc_16259_n10626;
  wire AES_CORE_DATAPATH__abc_16259_n10627;
  wire AES_CORE_DATAPATH__abc_16259_n10629;
  wire AES_CORE_DATAPATH__abc_16259_n10630;
  wire AES_CORE_DATAPATH__abc_16259_n10632;
  wire AES_CORE_DATAPATH__abc_16259_n10633;
  wire AES_CORE_DATAPATH__abc_16259_n10635;
  wire AES_CORE_DATAPATH__abc_16259_n10636;
  wire AES_CORE_DATAPATH__abc_16259_n10638;
  wire AES_CORE_DATAPATH__abc_16259_n10639;
  wire AES_CORE_DATAPATH__abc_16259_n10641;
  wire AES_CORE_DATAPATH__abc_16259_n10642;
  wire AES_CORE_DATAPATH__abc_16259_n10644;
  wire AES_CORE_DATAPATH__abc_16259_n10645;
  wire AES_CORE_DATAPATH__abc_16259_n10647;
  wire AES_CORE_DATAPATH__abc_16259_n10648;
  wire AES_CORE_DATAPATH__abc_16259_n10650;
  wire AES_CORE_DATAPATH__abc_16259_n10651;
  wire AES_CORE_DATAPATH__abc_16259_n10653;
  wire AES_CORE_DATAPATH__abc_16259_n10654;
  wire AES_CORE_DATAPATH__abc_16259_n10656;
  wire AES_CORE_DATAPATH__abc_16259_n10657;
  wire AES_CORE_DATAPATH__abc_16259_n10659;
  wire AES_CORE_DATAPATH__abc_16259_n10660;
  wire AES_CORE_DATAPATH__abc_16259_n10662;
  wire AES_CORE_DATAPATH__abc_16259_n10663;
  wire AES_CORE_DATAPATH__abc_16259_n10665;
  wire AES_CORE_DATAPATH__abc_16259_n10666;
  wire AES_CORE_DATAPATH__abc_16259_n10668;
  wire AES_CORE_DATAPATH__abc_16259_n10669;
  wire AES_CORE_DATAPATH__abc_16259_n10671;
  wire AES_CORE_DATAPATH__abc_16259_n10672;
  wire AES_CORE_DATAPATH__abc_16259_n10674;
  wire AES_CORE_DATAPATH__abc_16259_n10675;
  wire AES_CORE_DATAPATH__abc_16259_n10677;
  wire AES_CORE_DATAPATH__abc_16259_n10678;
  wire AES_CORE_DATAPATH__abc_16259_n10680;
  wire AES_CORE_DATAPATH__abc_16259_n10681;
  wire AES_CORE_DATAPATH__abc_16259_n10683;
  wire AES_CORE_DATAPATH__abc_16259_n10684;
  wire AES_CORE_DATAPATH__abc_16259_n10686;
  wire AES_CORE_DATAPATH__abc_16259_n10687;
  wire AES_CORE_DATAPATH__abc_16259_n10689;
  wire AES_CORE_DATAPATH__abc_16259_n10690;
  wire AES_CORE_DATAPATH__abc_16259_n10692;
  wire AES_CORE_DATAPATH__abc_16259_n10693;
  wire AES_CORE_DATAPATH__abc_16259_n10695;
  wire AES_CORE_DATAPATH__abc_16259_n10696;
  wire AES_CORE_DATAPATH__abc_16259_n10698;
  wire AES_CORE_DATAPATH__abc_16259_n10699;
  wire AES_CORE_DATAPATH__abc_16259_n10701;
  wire AES_CORE_DATAPATH__abc_16259_n10702;
  wire AES_CORE_DATAPATH__abc_16259_n10704;
  wire AES_CORE_DATAPATH__abc_16259_n10705;
  wire AES_CORE_DATAPATH__abc_16259_n10707;
  wire AES_CORE_DATAPATH__abc_16259_n10708;
  wire AES_CORE_DATAPATH__abc_16259_n10710;
  wire AES_CORE_DATAPATH__abc_16259_n10711;
  wire AES_CORE_DATAPATH__abc_16259_n10713;
  wire AES_CORE_DATAPATH__abc_16259_n10714;
  wire AES_CORE_DATAPATH__abc_16259_n2457_1;
  wire AES_CORE_DATAPATH__abc_16259_n2458;
  wire AES_CORE_DATAPATH__abc_16259_n2459_1;
  wire AES_CORE_DATAPATH__abc_16259_n2460;
  wire AES_CORE_DATAPATH__abc_16259_n2461_1;
  wire AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf5;
  wire AES_CORE_DATAPATH__abc_16259_n2462;
  wire AES_CORE_DATAPATH__abc_16259_n2462_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n2462_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n2462_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n2462_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n2462_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n2462_bF_buf5;
  wire AES_CORE_DATAPATH__abc_16259_n2462_bF_buf6;
  wire AES_CORE_DATAPATH__abc_16259_n2462_bF_buf7;
  wire AES_CORE_DATAPATH__abc_16259_n2463_1;
  wire AES_CORE_DATAPATH__abc_16259_n2464;
  wire AES_CORE_DATAPATH__abc_16259_n2465_1;
  wire AES_CORE_DATAPATH__abc_16259_n2466;
  wire AES_CORE_DATAPATH__abc_16259_n2467_1;
  wire AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf5;
  wire AES_CORE_DATAPATH__abc_16259_n2468;
  wire AES_CORE_DATAPATH__abc_16259_n2469_1;
  wire AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf5;
  wire AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf6;
  wire AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf7;
  wire AES_CORE_DATAPATH__abc_16259_n2470;
  wire AES_CORE_DATAPATH__abc_16259_n2471_1;
  wire AES_CORE_DATAPATH__abc_16259_n2472;
  wire AES_CORE_DATAPATH__abc_16259_n2473_1;
  wire AES_CORE_DATAPATH__abc_16259_n2474;
  wire AES_CORE_DATAPATH__abc_16259_n2474_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n2474_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n2474_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n2474_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n2474_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n2474_bF_buf5;
  wire AES_CORE_DATAPATH__abc_16259_n2475_1;
  wire AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf5;
  wire AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf6;
  wire AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf7;
  wire AES_CORE_DATAPATH__abc_16259_n2476;
  wire AES_CORE_DATAPATH__abc_16259_n2477_1;
  wire AES_CORE_DATAPATH__abc_16259_n2478;
  wire AES_CORE_DATAPATH__abc_16259_n2479_1;
  wire AES_CORE_DATAPATH__abc_16259_n2480;
  wire AES_CORE_DATAPATH__abc_16259_n2481_1;
  wire AES_CORE_DATAPATH__abc_16259_n2482;
  wire AES_CORE_DATAPATH__abc_16259_n2482_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n2482_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n2482_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n2482_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n2482_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n2482_bF_buf5;
  wire AES_CORE_DATAPATH__abc_16259_n2483_1;
  wire AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf5;
  wire AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf6;
  wire AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf7;
  wire AES_CORE_DATAPATH__abc_16259_n2484;
  wire AES_CORE_DATAPATH__abc_16259_n2484_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n2484_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n2484_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n2484_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n2484_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n2484_bF_buf5;
  wire AES_CORE_DATAPATH__abc_16259_n2484_bF_buf6;
  wire AES_CORE_DATAPATH__abc_16259_n2484_bF_buf7;
  wire AES_CORE_DATAPATH__abc_16259_n2485_1;
  wire AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf5;
  wire AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf6;
  wire AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf7;
  wire AES_CORE_DATAPATH__abc_16259_n2486;
  wire AES_CORE_DATAPATH__abc_16259_n2487_1;
  wire AES_CORE_DATAPATH__abc_16259_n2488;
  wire AES_CORE_DATAPATH__abc_16259_n2489_1;
  wire AES_CORE_DATAPATH__abc_16259_n2491_1;
  wire AES_CORE_DATAPATH__abc_16259_n2492_1;
  wire AES_CORE_DATAPATH__abc_16259_n2493;
  wire AES_CORE_DATAPATH__abc_16259_n2494_1;
  wire AES_CORE_DATAPATH__abc_16259_n2495;
  wire AES_CORE_DATAPATH__abc_16259_n2496;
  wire AES_CORE_DATAPATH__abc_16259_n2497_1;
  wire AES_CORE_DATAPATH__abc_16259_n2498;
  wire AES_CORE_DATAPATH__abc_16259_n2500;
  wire AES_CORE_DATAPATH__abc_16259_n2501_1;
  wire AES_CORE_DATAPATH__abc_16259_n2502;
  wire AES_CORE_DATAPATH__abc_16259_n2503_1;
  wire AES_CORE_DATAPATH__abc_16259_n2504_1;
  wire AES_CORE_DATAPATH__abc_16259_n2505;
  wire AES_CORE_DATAPATH__abc_16259_n2506_1;
  wire AES_CORE_DATAPATH__abc_16259_n2507;
  wire AES_CORE_DATAPATH__abc_16259_n2509_1;
  wire AES_CORE_DATAPATH__abc_16259_n2510;
  wire AES_CORE_DATAPATH__abc_16259_n2511_1;
  wire AES_CORE_DATAPATH__abc_16259_n2512;
  wire AES_CORE_DATAPATH__abc_16259_n2513_1;
  wire AES_CORE_DATAPATH__abc_16259_n2514_1;
  wire AES_CORE_DATAPATH__abc_16259_n2515;
  wire AES_CORE_DATAPATH__abc_16259_n2516_1;
  wire AES_CORE_DATAPATH__abc_16259_n2518_1;
  wire AES_CORE_DATAPATH__abc_16259_n2519_1;
  wire AES_CORE_DATAPATH__abc_16259_n2520;
  wire AES_CORE_DATAPATH__abc_16259_n2521_1;
  wire AES_CORE_DATAPATH__abc_16259_n2522;
  wire AES_CORE_DATAPATH__abc_16259_n2523_1;
  wire AES_CORE_DATAPATH__abc_16259_n2524_1;
  wire AES_CORE_DATAPATH__abc_16259_n2525;
  wire AES_CORE_DATAPATH__abc_16259_n2527;
  wire AES_CORE_DATAPATH__abc_16259_n2528_1;
  wire AES_CORE_DATAPATH__abc_16259_n2529_1;
  wire AES_CORE_DATAPATH__abc_16259_n2530;
  wire AES_CORE_DATAPATH__abc_16259_n2531_1;
  wire AES_CORE_DATAPATH__abc_16259_n2532;
  wire AES_CORE_DATAPATH__abc_16259_n2533_1;
  wire AES_CORE_DATAPATH__abc_16259_n2534_1;
  wire AES_CORE_DATAPATH__abc_16259_n2536_1;
  wire AES_CORE_DATAPATH__abc_16259_n2537;
  wire AES_CORE_DATAPATH__abc_16259_n2538_1;
  wire AES_CORE_DATAPATH__abc_16259_n2539_1;
  wire AES_CORE_DATAPATH__abc_16259_n2540;
  wire AES_CORE_DATAPATH__abc_16259_n2541_1;
  wire AES_CORE_DATAPATH__abc_16259_n2542;
  wire AES_CORE_DATAPATH__abc_16259_n2543_1;
  wire AES_CORE_DATAPATH__abc_16259_n2545;
  wire AES_CORE_DATAPATH__abc_16259_n2546_1;
  wire AES_CORE_DATAPATH__abc_16259_n2547;
  wire AES_CORE_DATAPATH__abc_16259_n2548_1;
  wire AES_CORE_DATAPATH__abc_16259_n2549_1;
  wire AES_CORE_DATAPATH__abc_16259_n2550;
  wire AES_CORE_DATAPATH__abc_16259_n2551_1;
  wire AES_CORE_DATAPATH__abc_16259_n2552;
  wire AES_CORE_DATAPATH__abc_16259_n2554_1;
  wire AES_CORE_DATAPATH__abc_16259_n2555;
  wire AES_CORE_DATAPATH__abc_16259_n2556_1;
  wire AES_CORE_DATAPATH__abc_16259_n2557;
  wire AES_CORE_DATAPATH__abc_16259_n2558_1;
  wire AES_CORE_DATAPATH__abc_16259_n2559_1;
  wire AES_CORE_DATAPATH__abc_16259_n2560;
  wire AES_CORE_DATAPATH__abc_16259_n2561_1;
  wire AES_CORE_DATAPATH__abc_16259_n2563_1;
  wire AES_CORE_DATAPATH__abc_16259_n2564_1;
  wire AES_CORE_DATAPATH__abc_16259_n2565;
  wire AES_CORE_DATAPATH__abc_16259_n2566_1;
  wire AES_CORE_DATAPATH__abc_16259_n2567;
  wire AES_CORE_DATAPATH__abc_16259_n2568_1;
  wire AES_CORE_DATAPATH__abc_16259_n2569_1;
  wire AES_CORE_DATAPATH__abc_16259_n2570;
  wire AES_CORE_DATAPATH__abc_16259_n2572;
  wire AES_CORE_DATAPATH__abc_16259_n2573_1;
  wire AES_CORE_DATAPATH__abc_16259_n2574_1;
  wire AES_CORE_DATAPATH__abc_16259_n2575;
  wire AES_CORE_DATAPATH__abc_16259_n2576_1;
  wire AES_CORE_DATAPATH__abc_16259_n2577;
  wire AES_CORE_DATAPATH__abc_16259_n2578_1;
  wire AES_CORE_DATAPATH__abc_16259_n2579_1;
  wire AES_CORE_DATAPATH__abc_16259_n2581_1;
  wire AES_CORE_DATAPATH__abc_16259_n2582;
  wire AES_CORE_DATAPATH__abc_16259_n2583_1;
  wire AES_CORE_DATAPATH__abc_16259_n2584_1;
  wire AES_CORE_DATAPATH__abc_16259_n2585;
  wire AES_CORE_DATAPATH__abc_16259_n2586_1;
  wire AES_CORE_DATAPATH__abc_16259_n2587;
  wire AES_CORE_DATAPATH__abc_16259_n2588_1;
  wire AES_CORE_DATAPATH__abc_16259_n2590;
  wire AES_CORE_DATAPATH__abc_16259_n2591_1;
  wire AES_CORE_DATAPATH__abc_16259_n2592;
  wire AES_CORE_DATAPATH__abc_16259_n2593_1;
  wire AES_CORE_DATAPATH__abc_16259_n2594_1;
  wire AES_CORE_DATAPATH__abc_16259_n2595;
  wire AES_CORE_DATAPATH__abc_16259_n2596_1;
  wire AES_CORE_DATAPATH__abc_16259_n2597;
  wire AES_CORE_DATAPATH__abc_16259_n2599_1;
  wire AES_CORE_DATAPATH__abc_16259_n2600;
  wire AES_CORE_DATAPATH__abc_16259_n2601_1;
  wire AES_CORE_DATAPATH__abc_16259_n2602;
  wire AES_CORE_DATAPATH__abc_16259_n2603_1;
  wire AES_CORE_DATAPATH__abc_16259_n2604_1;
  wire AES_CORE_DATAPATH__abc_16259_n2605;
  wire AES_CORE_DATAPATH__abc_16259_n2606_1;
  wire AES_CORE_DATAPATH__abc_16259_n2608_1;
  wire AES_CORE_DATAPATH__abc_16259_n2609_1;
  wire AES_CORE_DATAPATH__abc_16259_n2610;
  wire AES_CORE_DATAPATH__abc_16259_n2611_1;
  wire AES_CORE_DATAPATH__abc_16259_n2612;
  wire AES_CORE_DATAPATH__abc_16259_n2613_1;
  wire AES_CORE_DATAPATH__abc_16259_n2614_1;
  wire AES_CORE_DATAPATH__abc_16259_n2615;
  wire AES_CORE_DATAPATH__abc_16259_n2617;
  wire AES_CORE_DATAPATH__abc_16259_n2618_1;
  wire AES_CORE_DATAPATH__abc_16259_n2619_1;
  wire AES_CORE_DATAPATH__abc_16259_n2620;
  wire AES_CORE_DATAPATH__abc_16259_n2621_1;
  wire AES_CORE_DATAPATH__abc_16259_n2622;
  wire AES_CORE_DATAPATH__abc_16259_n2623_1;
  wire AES_CORE_DATAPATH__abc_16259_n2624_1;
  wire AES_CORE_DATAPATH__abc_16259_n2626_1;
  wire AES_CORE_DATAPATH__abc_16259_n2627;
  wire AES_CORE_DATAPATH__abc_16259_n2628_1;
  wire AES_CORE_DATAPATH__abc_16259_n2629_1;
  wire AES_CORE_DATAPATH__abc_16259_n2630;
  wire AES_CORE_DATAPATH__abc_16259_n2631_1;
  wire AES_CORE_DATAPATH__abc_16259_n2632;
  wire AES_CORE_DATAPATH__abc_16259_n2633_1;
  wire AES_CORE_DATAPATH__abc_16259_n2635;
  wire AES_CORE_DATAPATH__abc_16259_n2636_1;
  wire AES_CORE_DATAPATH__abc_16259_n2637;
  wire AES_CORE_DATAPATH__abc_16259_n2638_1;
  wire AES_CORE_DATAPATH__abc_16259_n2639_1;
  wire AES_CORE_DATAPATH__abc_16259_n2640;
  wire AES_CORE_DATAPATH__abc_16259_n2641_1;
  wire AES_CORE_DATAPATH__abc_16259_n2642;
  wire AES_CORE_DATAPATH__abc_16259_n2644_1;
  wire AES_CORE_DATAPATH__abc_16259_n2645;
  wire AES_CORE_DATAPATH__abc_16259_n2646_1;
  wire AES_CORE_DATAPATH__abc_16259_n2647;
  wire AES_CORE_DATAPATH__abc_16259_n2648_1;
  wire AES_CORE_DATAPATH__abc_16259_n2649_1;
  wire AES_CORE_DATAPATH__abc_16259_n2650;
  wire AES_CORE_DATAPATH__abc_16259_n2651_1;
  wire AES_CORE_DATAPATH__abc_16259_n2653_1;
  wire AES_CORE_DATAPATH__abc_16259_n2654_1;
  wire AES_CORE_DATAPATH__abc_16259_n2655;
  wire AES_CORE_DATAPATH__abc_16259_n2656_1;
  wire AES_CORE_DATAPATH__abc_16259_n2657;
  wire AES_CORE_DATAPATH__abc_16259_n2658_1;
  wire AES_CORE_DATAPATH__abc_16259_n2659;
  wire AES_CORE_DATAPATH__abc_16259_n2660;
  wire AES_CORE_DATAPATH__abc_16259_n2662;
  wire AES_CORE_DATAPATH__abc_16259_n2663_1;
  wire AES_CORE_DATAPATH__abc_16259_n2664;
  wire AES_CORE_DATAPATH__abc_16259_n2665_1;
  wire AES_CORE_DATAPATH__abc_16259_n2666;
  wire AES_CORE_DATAPATH__abc_16259_n2667_1;
  wire AES_CORE_DATAPATH__abc_16259_n2668;
  wire AES_CORE_DATAPATH__abc_16259_n2669_1;
  wire AES_CORE_DATAPATH__abc_16259_n2671_1;
  wire AES_CORE_DATAPATH__abc_16259_n2672;
  wire AES_CORE_DATAPATH__abc_16259_n2673_1;
  wire AES_CORE_DATAPATH__abc_16259_n2674;
  wire AES_CORE_DATAPATH__abc_16259_n2675_1;
  wire AES_CORE_DATAPATH__abc_16259_n2676;
  wire AES_CORE_DATAPATH__abc_16259_n2677_1;
  wire AES_CORE_DATAPATH__abc_16259_n2678;
  wire AES_CORE_DATAPATH__abc_16259_n2680;
  wire AES_CORE_DATAPATH__abc_16259_n2681_1;
  wire AES_CORE_DATAPATH__abc_16259_n2682;
  wire AES_CORE_DATAPATH__abc_16259_n2683_1;
  wire AES_CORE_DATAPATH__abc_16259_n2684;
  wire AES_CORE_DATAPATH__abc_16259_n2685_1;
  wire AES_CORE_DATAPATH__abc_16259_n2686;
  wire AES_CORE_DATAPATH__abc_16259_n2687_1;
  wire AES_CORE_DATAPATH__abc_16259_n2689_1;
  wire AES_CORE_DATAPATH__abc_16259_n2690;
  wire AES_CORE_DATAPATH__abc_16259_n2691_1;
  wire AES_CORE_DATAPATH__abc_16259_n2692;
  wire AES_CORE_DATAPATH__abc_16259_n2693_1;
  wire AES_CORE_DATAPATH__abc_16259_n2694;
  wire AES_CORE_DATAPATH__abc_16259_n2695_1;
  wire AES_CORE_DATAPATH__abc_16259_n2696;
  wire AES_CORE_DATAPATH__abc_16259_n2698;
  wire AES_CORE_DATAPATH__abc_16259_n2699_1;
  wire AES_CORE_DATAPATH__abc_16259_n2700;
  wire AES_CORE_DATAPATH__abc_16259_n2701_1;
  wire AES_CORE_DATAPATH__abc_16259_n2702;
  wire AES_CORE_DATAPATH__abc_16259_n2703_1;
  wire AES_CORE_DATAPATH__abc_16259_n2704;
  wire AES_CORE_DATAPATH__abc_16259_n2705_1;
  wire AES_CORE_DATAPATH__abc_16259_n2707_1;
  wire AES_CORE_DATAPATH__abc_16259_n2708;
  wire AES_CORE_DATAPATH__abc_16259_n2709_1;
  wire AES_CORE_DATAPATH__abc_16259_n2710;
  wire AES_CORE_DATAPATH__abc_16259_n2711_1;
  wire AES_CORE_DATAPATH__abc_16259_n2712;
  wire AES_CORE_DATAPATH__abc_16259_n2713_1;
  wire AES_CORE_DATAPATH__abc_16259_n2714;
  wire AES_CORE_DATAPATH__abc_16259_n2716;
  wire AES_CORE_DATAPATH__abc_16259_n2717_1;
  wire AES_CORE_DATAPATH__abc_16259_n2718;
  wire AES_CORE_DATAPATH__abc_16259_n2719_1;
  wire AES_CORE_DATAPATH__abc_16259_n2720;
  wire AES_CORE_DATAPATH__abc_16259_n2721_1;
  wire AES_CORE_DATAPATH__abc_16259_n2722;
  wire AES_CORE_DATAPATH__abc_16259_n2723_1;
  wire AES_CORE_DATAPATH__abc_16259_n2725;
  wire AES_CORE_DATAPATH__abc_16259_n2726;
  wire AES_CORE_DATAPATH__abc_16259_n2727_1;
  wire AES_CORE_DATAPATH__abc_16259_n2728;
  wire AES_CORE_DATAPATH__abc_16259_n2729;
  wire AES_CORE_DATAPATH__abc_16259_n2730;
  wire AES_CORE_DATAPATH__abc_16259_n2731_1;
  wire AES_CORE_DATAPATH__abc_16259_n2732;
  wire AES_CORE_DATAPATH__abc_16259_n2734;
  wire AES_CORE_DATAPATH__abc_16259_n2735_1;
  wire AES_CORE_DATAPATH__abc_16259_n2736;
  wire AES_CORE_DATAPATH__abc_16259_n2737_1;
  wire AES_CORE_DATAPATH__abc_16259_n2738;
  wire AES_CORE_DATAPATH__abc_16259_n2739;
  wire AES_CORE_DATAPATH__abc_16259_n2740;
  wire AES_CORE_DATAPATH__abc_16259_n2741;
  wire AES_CORE_DATAPATH__abc_16259_n2743;
  wire AES_CORE_DATAPATH__abc_16259_n2744;
  wire AES_CORE_DATAPATH__abc_16259_n2745;
  wire AES_CORE_DATAPATH__abc_16259_n2746_1;
  wire AES_CORE_DATAPATH__abc_16259_n2747;
  wire AES_CORE_DATAPATH__abc_16259_n2748;
  wire AES_CORE_DATAPATH__abc_16259_n2749;
  wire AES_CORE_DATAPATH__abc_16259_n2750;
  wire AES_CORE_DATAPATH__abc_16259_n2752_1;
  wire AES_CORE_DATAPATH__abc_16259_n2753_1;
  wire AES_CORE_DATAPATH__abc_16259_n2754;
  wire AES_CORE_DATAPATH__abc_16259_n2755_1;
  wire AES_CORE_DATAPATH__abc_16259_n2756_1;
  wire AES_CORE_DATAPATH__abc_16259_n2757;
  wire AES_CORE_DATAPATH__abc_16259_n2758;
  wire AES_CORE_DATAPATH__abc_16259_n2759;
  wire AES_CORE_DATAPATH__abc_16259_n2761;
  wire AES_CORE_DATAPATH__abc_16259_n2762_1;
  wire AES_CORE_DATAPATH__abc_16259_n2763;
  wire AES_CORE_DATAPATH__abc_16259_n2764_1;
  wire AES_CORE_DATAPATH__abc_16259_n2765;
  wire AES_CORE_DATAPATH__abc_16259_n2766;
  wire AES_CORE_DATAPATH__abc_16259_n2767;
  wire AES_CORE_DATAPATH__abc_16259_n2768;
  wire AES_CORE_DATAPATH__abc_16259_n2770;
  wire AES_CORE_DATAPATH__abc_16259_n2771_1;
  wire AES_CORE_DATAPATH__abc_16259_n2772_1;
  wire AES_CORE_DATAPATH__abc_16259_n2773;
  wire AES_CORE_DATAPATH__abc_16259_n2774;
  wire AES_CORE_DATAPATH__abc_16259_n2774_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n2774_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n2774_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n2774_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n2774_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n2775_1;
  wire AES_CORE_DATAPATH__abc_16259_n2776;
  wire AES_CORE_DATAPATH__abc_16259_n2777_1;
  wire AES_CORE_DATAPATH__abc_16259_n2778;
  wire AES_CORE_DATAPATH__abc_16259_n2778_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n2778_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n2778_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n2778_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n2778_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n2779_1;
  wire AES_CORE_DATAPATH__abc_16259_n2780;
  wire AES_CORE_DATAPATH__abc_16259_n2781_1;
  wire AES_CORE_DATAPATH__abc_16259_n2782;
  wire AES_CORE_DATAPATH__abc_16259_n2782_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n2782_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n2782_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n2782_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n2782_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n2783;
  wire AES_CORE_DATAPATH__abc_16259_n2784;
  wire AES_CORE_DATAPATH__abc_16259_n2785;
  wire AES_CORE_DATAPATH__abc_16259_n2786;
  wire AES_CORE_DATAPATH__abc_16259_n2786_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n2786_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n2786_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n2786_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n2786_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n2787;
  wire AES_CORE_DATAPATH__abc_16259_n2788;
  wire AES_CORE_DATAPATH__abc_16259_n2789;
  wire AES_CORE_DATAPATH__abc_16259_n2789_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n2789_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n2789_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n2789_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n2789_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n2790;
  wire AES_CORE_DATAPATH__abc_16259_n2791;
  wire AES_CORE_DATAPATH__abc_16259_n2792;
  wire AES_CORE_DATAPATH__abc_16259_n2793_1;
  wire AES_CORE_DATAPATH__abc_16259_n2794;
  wire AES_CORE_DATAPATH__abc_16259_n2796;
  wire AES_CORE_DATAPATH__abc_16259_n2796_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n2796_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n2796_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n2796_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n2796_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n2796_bF_buf5;
  wire AES_CORE_DATAPATH__abc_16259_n2796_bF_buf6;
  wire AES_CORE_DATAPATH__abc_16259_n2796_bF_buf7;
  wire AES_CORE_DATAPATH__abc_16259_n2797;
  wire AES_CORE_DATAPATH__abc_16259_n2798;
  wire AES_CORE_DATAPATH__abc_16259_n2798_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n2798_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n2798_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n2798_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n2798_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n2799;
  wire AES_CORE_DATAPATH__abc_16259_n2800_1;
  wire AES_CORE_DATAPATH__abc_16259_n2801_1;
  wire AES_CORE_DATAPATH__abc_16259_n2802;
  wire AES_CORE_DATAPATH__abc_16259_n2802_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n2802_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n2802_bF_buf10;
  wire AES_CORE_DATAPATH__abc_16259_n2802_bF_buf11;
  wire AES_CORE_DATAPATH__abc_16259_n2802_bF_buf12;
  wire AES_CORE_DATAPATH__abc_16259_n2802_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n2802_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n2802_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n2802_bF_buf5;
  wire AES_CORE_DATAPATH__abc_16259_n2802_bF_buf6;
  wire AES_CORE_DATAPATH__abc_16259_n2802_bF_buf7;
  wire AES_CORE_DATAPATH__abc_16259_n2802_bF_buf8;
  wire AES_CORE_DATAPATH__abc_16259_n2802_bF_buf9;
  wire AES_CORE_DATAPATH__abc_16259_n2803;
  wire AES_CORE_DATAPATH__abc_16259_n2803_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n2803_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n2803_bF_buf10;
  wire AES_CORE_DATAPATH__abc_16259_n2803_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n2803_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n2803_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n2803_bF_buf5;
  wire AES_CORE_DATAPATH__abc_16259_n2803_bF_buf6;
  wire AES_CORE_DATAPATH__abc_16259_n2803_bF_buf7;
  wire AES_CORE_DATAPATH__abc_16259_n2803_bF_buf8;
  wire AES_CORE_DATAPATH__abc_16259_n2803_bF_buf9;
  wire AES_CORE_DATAPATH__abc_16259_n2804_1;
  wire AES_CORE_DATAPATH__abc_16259_n2804_1_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n2804_1_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n2804_1_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n2804_1_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n2804_1_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n2805;
  wire AES_CORE_DATAPATH__abc_16259_n2806_1;
  wire AES_CORE_DATAPATH__abc_16259_n2807;
  wire AES_CORE_DATAPATH__abc_16259_n2807_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n2807_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n2807_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n2807_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n2807_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n2807_bF_buf5;
  wire AES_CORE_DATAPATH__abc_16259_n2808_1;
  wire AES_CORE_DATAPATH__abc_16259_n2809;
  wire AES_CORE_DATAPATH__abc_16259_n2810_1;
  wire AES_CORE_DATAPATH__abc_16259_n2811;
  wire AES_CORE_DATAPATH__abc_16259_n2812;
  wire AES_CORE_DATAPATH__abc_16259_n2813;
  wire AES_CORE_DATAPATH__abc_16259_n2814;
  wire AES_CORE_DATAPATH__abc_16259_n2815;
  wire AES_CORE_DATAPATH__abc_16259_n2816;
  wire AES_CORE_DATAPATH__abc_16259_n2817;
  wire AES_CORE_DATAPATH__abc_16259_n2818;
  wire AES_CORE_DATAPATH__abc_16259_n2819;
  wire AES_CORE_DATAPATH__abc_16259_n2820;
  wire AES_CORE_DATAPATH__abc_16259_n2821;
  wire AES_CORE_DATAPATH__abc_16259_n2822_1;
  wire AES_CORE_DATAPATH__abc_16259_n2823;
  wire AES_CORE_DATAPATH__abc_16259_n2824_1;
  wire AES_CORE_DATAPATH__abc_16259_n2825;
  wire AES_CORE_DATAPATH__abc_16259_n2826;
  wire AES_CORE_DATAPATH__abc_16259_n2826_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n2826_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n2826_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n2826_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n2826_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n2827;
  wire AES_CORE_DATAPATH__abc_16259_n2828;
  wire AES_CORE_DATAPATH__abc_16259_n2829_1;
  wire AES_CORE_DATAPATH__abc_16259_n2830_1;
  wire AES_CORE_DATAPATH__abc_16259_n2830_1_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n2830_1_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n2830_1_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n2830_1_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n2830_1_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n2831;
  wire AES_CORE_DATAPATH__abc_16259_n2832;
  wire AES_CORE_DATAPATH__abc_16259_n2833_1;
  wire AES_CORE_DATAPATH__abc_16259_n2834;
  wire AES_CORE_DATAPATH__abc_16259_n2835_1;
  wire AES_CORE_DATAPATH__abc_16259_n2836;
  wire AES_CORE_DATAPATH__abc_16259_n2837_1;
  wire AES_CORE_DATAPATH__abc_16259_n2837_1_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n2837_1_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n2837_1_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n2837_1_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n2837_1_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n2838;
  wire AES_CORE_DATAPATH__abc_16259_n2839_1;
  wire AES_CORE_DATAPATH__abc_16259_n2840;
  wire AES_CORE_DATAPATH__abc_16259_n2841;
  wire AES_CORE_DATAPATH__abc_16259_n2841_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n2841_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n2841_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n2841_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n2841_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n2842;
  wire AES_CORE_DATAPATH__abc_16259_n2844;
  wire AES_CORE_DATAPATH__abc_16259_n2845;
  wire AES_CORE_DATAPATH__abc_16259_n2846;
  wire AES_CORE_DATAPATH__abc_16259_n2847;
  wire AES_CORE_DATAPATH__abc_16259_n2848;
  wire AES_CORE_DATAPATH__abc_16259_n2849;
  wire AES_CORE_DATAPATH__abc_16259_n2850;
  wire AES_CORE_DATAPATH__abc_16259_n2851_1;
  wire AES_CORE_DATAPATH__abc_16259_n2852;
  wire AES_CORE_DATAPATH__abc_16259_n2853_1;
  wire AES_CORE_DATAPATH__abc_16259_n2853_1_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n2853_1_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n2853_1_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n2853_1_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n2853_1_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n2854;
  wire AES_CORE_DATAPATH__abc_16259_n2855;
  wire AES_CORE_DATAPATH__abc_16259_n2855_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n2855_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n2855_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n2855_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n2855_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n2856;
  wire AES_CORE_DATAPATH__abc_16259_n2857;
  wire AES_CORE_DATAPATH__abc_16259_n2857_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n2857_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n2857_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n2857_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n2857_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n2858_1;
  wire AES_CORE_DATAPATH__abc_16259_n2859_1;
  wire AES_CORE_DATAPATH__abc_16259_n2860;
  wire AES_CORE_DATAPATH__abc_16259_n2861;
  wire AES_CORE_DATAPATH__abc_16259_n2862_1;
  wire AES_CORE_DATAPATH__abc_16259_n2863;
  wire AES_CORE_DATAPATH__abc_16259_n2864_1;
  wire AES_CORE_DATAPATH__abc_16259_n2864_1_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n2864_1_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n2864_1_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n2864_1_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n2864_1_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n2865;
  wire AES_CORE_DATAPATH__abc_16259_n2866_1;
  wire AES_CORE_DATAPATH__abc_16259_n2867;
  wire AES_CORE_DATAPATH__abc_16259_n2868_1;
  wire AES_CORE_DATAPATH__abc_16259_n2869;
  wire AES_CORE_DATAPATH__abc_16259_n2870;
  wire AES_CORE_DATAPATH__abc_16259_n2872;
  wire AES_CORE_DATAPATH__abc_16259_n2873;
  wire AES_CORE_DATAPATH__abc_16259_n2874;
  wire AES_CORE_DATAPATH__abc_16259_n2875;
  wire AES_CORE_DATAPATH__abc_16259_n2876;
  wire AES_CORE_DATAPATH__abc_16259_n2877;
  wire AES_CORE_DATAPATH__abc_16259_n2878;
  wire AES_CORE_DATAPATH__abc_16259_n2879;
  wire AES_CORE_DATAPATH__abc_16259_n2880_1;
  wire AES_CORE_DATAPATH__abc_16259_n2881;
  wire AES_CORE_DATAPATH__abc_16259_n2882_1;
  wire AES_CORE_DATAPATH__abc_16259_n2883;
  wire AES_CORE_DATAPATH__abc_16259_n2885;
  wire AES_CORE_DATAPATH__abc_16259_n2886;
  wire AES_CORE_DATAPATH__abc_16259_n2887_1;
  wire AES_CORE_DATAPATH__abc_16259_n2887_1_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n2887_1_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n2887_1_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n2887_1_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n2887_1_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n2888_1;
  wire AES_CORE_DATAPATH__abc_16259_n2889;
  wire AES_CORE_DATAPATH__abc_16259_n2890;
  wire AES_CORE_DATAPATH__abc_16259_n2891_1;
  wire AES_CORE_DATAPATH__abc_16259_n2892;
  wire AES_CORE_DATAPATH__abc_16259_n2894;
  wire AES_CORE_DATAPATH__abc_16259_n2895_1;
  wire AES_CORE_DATAPATH__abc_16259_n2896;
  wire AES_CORE_DATAPATH__abc_16259_n2897_1;
  wire AES_CORE_DATAPATH__abc_16259_n2898;
  wire AES_CORE_DATAPATH__abc_16259_n2899;
  wire AES_CORE_DATAPATH__abc_16259_n2900;
  wire AES_CORE_DATAPATH__abc_16259_n2901;
  wire AES_CORE_DATAPATH__abc_16259_n2902;
  wire AES_CORE_DATAPATH__abc_16259_n2903;
  wire AES_CORE_DATAPATH__abc_16259_n2904;
  wire AES_CORE_DATAPATH__abc_16259_n2905;
  wire AES_CORE_DATAPATH__abc_16259_n2906;
  wire AES_CORE_DATAPATH__abc_16259_n2907;
  wire AES_CORE_DATAPATH__abc_16259_n2908;
  wire AES_CORE_DATAPATH__abc_16259_n2909_1;
  wire AES_CORE_DATAPATH__abc_16259_n2910;
  wire AES_CORE_DATAPATH__abc_16259_n2911_1;
  wire AES_CORE_DATAPATH__abc_16259_n2913;
  wire AES_CORE_DATAPATH__abc_16259_n2914;
  wire AES_CORE_DATAPATH__abc_16259_n2915;
  wire AES_CORE_DATAPATH__abc_16259_n2916_1;
  wire AES_CORE_DATAPATH__abc_16259_n2917_1;
  wire AES_CORE_DATAPATH__abc_16259_n2918;
  wire AES_CORE_DATAPATH__abc_16259_n2919;
  wire AES_CORE_DATAPATH__abc_16259_n2920_1;
  wire AES_CORE_DATAPATH__abc_16259_n2921;
  wire AES_CORE_DATAPATH__abc_16259_n2922_1;
  wire AES_CORE_DATAPATH__abc_16259_n2923;
  wire AES_CORE_DATAPATH__abc_16259_n2924_1;
  wire AES_CORE_DATAPATH__abc_16259_n2926_1;
  wire AES_CORE_DATAPATH__abc_16259_n2927;
  wire AES_CORE_DATAPATH__abc_16259_n2928;
  wire AES_CORE_DATAPATH__abc_16259_n2929;
  wire AES_CORE_DATAPATH__abc_16259_n2930;
  wire AES_CORE_DATAPATH__abc_16259_n2931;
  wire AES_CORE_DATAPATH__abc_16259_n2932;
  wire AES_CORE_DATAPATH__abc_16259_n2934;
  wire AES_CORE_DATAPATH__abc_16259_n2935;
  wire AES_CORE_DATAPATH__abc_16259_n2936;
  wire AES_CORE_DATAPATH__abc_16259_n2937;
  wire AES_CORE_DATAPATH__abc_16259_n2938_1;
  wire AES_CORE_DATAPATH__abc_16259_n2939;
  wire AES_CORE_DATAPATH__abc_16259_n2940_1;
  wire AES_CORE_DATAPATH__abc_16259_n2941;
  wire AES_CORE_DATAPATH__abc_16259_n2942;
  wire AES_CORE_DATAPATH__abc_16259_n2943;
  wire AES_CORE_DATAPATH__abc_16259_n2944;
  wire AES_CORE_DATAPATH__abc_16259_n2945_1;
  wire AES_CORE_DATAPATH__abc_16259_n2946_1;
  wire AES_CORE_DATAPATH__abc_16259_n2947;
  wire AES_CORE_DATAPATH__abc_16259_n2948;
  wire AES_CORE_DATAPATH__abc_16259_n2949_1;
  wire AES_CORE_DATAPATH__abc_16259_n2950;
  wire AES_CORE_DATAPATH__abc_16259_n2951_1;
  wire AES_CORE_DATAPATH__abc_16259_n2953_1;
  wire AES_CORE_DATAPATH__abc_16259_n2954;
  wire AES_CORE_DATAPATH__abc_16259_n2955_1;
  wire AES_CORE_DATAPATH__abc_16259_n2956;
  wire AES_CORE_DATAPATH__abc_16259_n2957;
  wire AES_CORE_DATAPATH__abc_16259_n2958;
  wire AES_CORE_DATAPATH__abc_16259_n2959;
  wire AES_CORE_DATAPATH__abc_16259_n2960;
  wire AES_CORE_DATAPATH__abc_16259_n2961;
  wire AES_CORE_DATAPATH__abc_16259_n2962;
  wire AES_CORE_DATAPATH__abc_16259_n2963;
  wire AES_CORE_DATAPATH__abc_16259_n2964;
  wire AES_CORE_DATAPATH__abc_16259_n2966;
  wire AES_CORE_DATAPATH__abc_16259_n2967_1;
  wire AES_CORE_DATAPATH__abc_16259_n2968;
  wire AES_CORE_DATAPATH__abc_16259_n2969_1;
  wire AES_CORE_DATAPATH__abc_16259_n2970;
  wire AES_CORE_DATAPATH__abc_16259_n2971;
  wire AES_CORE_DATAPATH__abc_16259_n2972;
  wire AES_CORE_DATAPATH__abc_16259_n2974_1;
  wire AES_CORE_DATAPATH__abc_16259_n2975_1;
  wire AES_CORE_DATAPATH__abc_16259_n2976;
  wire AES_CORE_DATAPATH__abc_16259_n2977;
  wire AES_CORE_DATAPATH__abc_16259_n2978_1;
  wire AES_CORE_DATAPATH__abc_16259_n2979;
  wire AES_CORE_DATAPATH__abc_16259_n2980_1;
  wire AES_CORE_DATAPATH__abc_16259_n2981;
  wire AES_CORE_DATAPATH__abc_16259_n2982_1;
  wire AES_CORE_DATAPATH__abc_16259_n2983;
  wire AES_CORE_DATAPATH__abc_16259_n2984_1;
  wire AES_CORE_DATAPATH__abc_16259_n2985;
  wire AES_CORE_DATAPATH__abc_16259_n2986;
  wire AES_CORE_DATAPATH__abc_16259_n2987;
  wire AES_CORE_DATAPATH__abc_16259_n2988;
  wire AES_CORE_DATAPATH__abc_16259_n2989;
  wire AES_CORE_DATAPATH__abc_16259_n2990;
  wire AES_CORE_DATAPATH__abc_16259_n2991;
  wire AES_CORE_DATAPATH__abc_16259_n2993;
  wire AES_CORE_DATAPATH__abc_16259_n2994;
  wire AES_CORE_DATAPATH__abc_16259_n2995;
  wire AES_CORE_DATAPATH__abc_16259_n2996_1;
  wire AES_CORE_DATAPATH__abc_16259_n2997;
  wire AES_CORE_DATAPATH__abc_16259_n2998_1;
  wire AES_CORE_DATAPATH__abc_16259_n2999;
  wire AES_CORE_DATAPATH__abc_16259_n3000;
  wire AES_CORE_DATAPATH__abc_16259_n3001;
  wire AES_CORE_DATAPATH__abc_16259_n3002;
  wire AES_CORE_DATAPATH__abc_16259_n3003_1;
  wire AES_CORE_DATAPATH__abc_16259_n3004_1;
  wire AES_CORE_DATAPATH__abc_16259_n3006;
  wire AES_CORE_DATAPATH__abc_16259_n3007_1;
  wire AES_CORE_DATAPATH__abc_16259_n3008;
  wire AES_CORE_DATAPATH__abc_16259_n3009_1;
  wire AES_CORE_DATAPATH__abc_16259_n3010;
  wire AES_CORE_DATAPATH__abc_16259_n3011_1;
  wire AES_CORE_DATAPATH__abc_16259_n3012;
  wire AES_CORE_DATAPATH__abc_16259_n3014;
  wire AES_CORE_DATAPATH__abc_16259_n3015;
  wire AES_CORE_DATAPATH__abc_16259_n3016;
  wire AES_CORE_DATAPATH__abc_16259_n3017;
  wire AES_CORE_DATAPATH__abc_16259_n3018;
  wire AES_CORE_DATAPATH__abc_16259_n3019;
  wire AES_CORE_DATAPATH__abc_16259_n3020;
  wire AES_CORE_DATAPATH__abc_16259_n3021;
  wire AES_CORE_DATAPATH__abc_16259_n3022;
  wire AES_CORE_DATAPATH__abc_16259_n3023;
  wire AES_CORE_DATAPATH__abc_16259_n3024;
  wire AES_CORE_DATAPATH__abc_16259_n3025_1;
  wire AES_CORE_DATAPATH__abc_16259_n3026;
  wire AES_CORE_DATAPATH__abc_16259_n3027_1;
  wire AES_CORE_DATAPATH__abc_16259_n3028;
  wire AES_CORE_DATAPATH__abc_16259_n3029;
  wire AES_CORE_DATAPATH__abc_16259_n3030;
  wire AES_CORE_DATAPATH__abc_16259_n3031;
  wire AES_CORE_DATAPATH__abc_16259_n3033_1;
  wire AES_CORE_DATAPATH__abc_16259_n3034;
  wire AES_CORE_DATAPATH__abc_16259_n3035;
  wire AES_CORE_DATAPATH__abc_16259_n3036_1;
  wire AES_CORE_DATAPATH__abc_16259_n3037;
  wire AES_CORE_DATAPATH__abc_16259_n3038_1;
  wire AES_CORE_DATAPATH__abc_16259_n3039;
  wire AES_CORE_DATAPATH__abc_16259_n3040_1;
  wire AES_CORE_DATAPATH__abc_16259_n3041;
  wire AES_CORE_DATAPATH__abc_16259_n3042_1;
  wire AES_CORE_DATAPATH__abc_16259_n3043;
  wire AES_CORE_DATAPATH__abc_16259_n3044;
  wire AES_CORE_DATAPATH__abc_16259_n3046;
  wire AES_CORE_DATAPATH__abc_16259_n3047;
  wire AES_CORE_DATAPATH__abc_16259_n3048;
  wire AES_CORE_DATAPATH__abc_16259_n3049;
  wire AES_CORE_DATAPATH__abc_16259_n3050;
  wire AES_CORE_DATAPATH__abc_16259_n3051;
  wire AES_CORE_DATAPATH__abc_16259_n3052;
  wire AES_CORE_DATAPATH__abc_16259_n3054_1;
  wire AES_CORE_DATAPATH__abc_16259_n3055;
  wire AES_CORE_DATAPATH__abc_16259_n3056_1;
  wire AES_CORE_DATAPATH__abc_16259_n3057;
  wire AES_CORE_DATAPATH__abc_16259_n3058;
  wire AES_CORE_DATAPATH__abc_16259_n3059;
  wire AES_CORE_DATAPATH__abc_16259_n3060;
  wire AES_CORE_DATAPATH__abc_16259_n3061_1;
  wire AES_CORE_DATAPATH__abc_16259_n3062_1;
  wire AES_CORE_DATAPATH__abc_16259_n3063;
  wire AES_CORE_DATAPATH__abc_16259_n3064;
  wire AES_CORE_DATAPATH__abc_16259_n3065_1;
  wire AES_CORE_DATAPATH__abc_16259_n3066;
  wire AES_CORE_DATAPATH__abc_16259_n3067_1;
  wire AES_CORE_DATAPATH__abc_16259_n3068;
  wire AES_CORE_DATAPATH__abc_16259_n3069_1;
  wire AES_CORE_DATAPATH__abc_16259_n3070;
  wire AES_CORE_DATAPATH__abc_16259_n3071_1;
  wire AES_CORE_DATAPATH__abc_16259_n3073;
  wire AES_CORE_DATAPATH__abc_16259_n3074;
  wire AES_CORE_DATAPATH__abc_16259_n3075;
  wire AES_CORE_DATAPATH__abc_16259_n3076;
  wire AES_CORE_DATAPATH__abc_16259_n3077;
  wire AES_CORE_DATAPATH__abc_16259_n3078;
  wire AES_CORE_DATAPATH__abc_16259_n3079;
  wire AES_CORE_DATAPATH__abc_16259_n3080;
  wire AES_CORE_DATAPATH__abc_16259_n3081;
  wire AES_CORE_DATAPATH__abc_16259_n3082;
  wire AES_CORE_DATAPATH__abc_16259_n3083_1;
  wire AES_CORE_DATAPATH__abc_16259_n3084;
  wire AES_CORE_DATAPATH__abc_16259_n3086;
  wire AES_CORE_DATAPATH__abc_16259_n3087;
  wire AES_CORE_DATAPATH__abc_16259_n3088;
  wire AES_CORE_DATAPATH__abc_16259_n3089;
  wire AES_CORE_DATAPATH__abc_16259_n3090_1;
  wire AES_CORE_DATAPATH__abc_16259_n3091_1;
  wire AES_CORE_DATAPATH__abc_16259_n3092;
  wire AES_CORE_DATAPATH__abc_16259_n3094_1;
  wire AES_CORE_DATAPATH__abc_16259_n3095;
  wire AES_CORE_DATAPATH__abc_16259_n3096_1;
  wire AES_CORE_DATAPATH__abc_16259_n3097;
  wire AES_CORE_DATAPATH__abc_16259_n3098_1;
  wire AES_CORE_DATAPATH__abc_16259_n3099;
  wire AES_CORE_DATAPATH__abc_16259_n3100_1;
  wire AES_CORE_DATAPATH__abc_16259_n3101;
  wire AES_CORE_DATAPATH__abc_16259_n3102;
  wire AES_CORE_DATAPATH__abc_16259_n3103;
  wire AES_CORE_DATAPATH__abc_16259_n3104;
  wire AES_CORE_DATAPATH__abc_16259_n3105;
  wire AES_CORE_DATAPATH__abc_16259_n3106;
  wire AES_CORE_DATAPATH__abc_16259_n3107;
  wire AES_CORE_DATAPATH__abc_16259_n3108;
  wire AES_CORE_DATAPATH__abc_16259_n3109;
  wire AES_CORE_DATAPATH__abc_16259_n3110;
  wire AES_CORE_DATAPATH__abc_16259_n3111;
  wire AES_CORE_DATAPATH__abc_16259_n3113;
  wire AES_CORE_DATAPATH__abc_16259_n3114_1;
  wire AES_CORE_DATAPATH__abc_16259_n3115;
  wire AES_CORE_DATAPATH__abc_16259_n3116;
  wire AES_CORE_DATAPATH__abc_16259_n3117;
  wire AES_CORE_DATAPATH__abc_16259_n3118;
  wire AES_CORE_DATAPATH__abc_16259_n3119_1;
  wire AES_CORE_DATAPATH__abc_16259_n3120_1;
  wire AES_CORE_DATAPATH__abc_16259_n3121;
  wire AES_CORE_DATAPATH__abc_16259_n3122;
  wire AES_CORE_DATAPATH__abc_16259_n3123_1;
  wire AES_CORE_DATAPATH__abc_16259_n3124;
  wire AES_CORE_DATAPATH__abc_16259_n3126;
  wire AES_CORE_DATAPATH__abc_16259_n3127_1;
  wire AES_CORE_DATAPATH__abc_16259_n3128;
  wire AES_CORE_DATAPATH__abc_16259_n3129_1;
  wire AES_CORE_DATAPATH__abc_16259_n3130;
  wire AES_CORE_DATAPATH__abc_16259_n3131;
  wire AES_CORE_DATAPATH__abc_16259_n3132;
  wire AES_CORE_DATAPATH__abc_16259_n3134;
  wire AES_CORE_DATAPATH__abc_16259_n3135;
  wire AES_CORE_DATAPATH__abc_16259_n3136;
  wire AES_CORE_DATAPATH__abc_16259_n3137;
  wire AES_CORE_DATAPATH__abc_16259_n3138;
  wire AES_CORE_DATAPATH__abc_16259_n3139;
  wire AES_CORE_DATAPATH__abc_16259_n3140;
  wire AES_CORE_DATAPATH__abc_16259_n3141_1;
  wire AES_CORE_DATAPATH__abc_16259_n3142;
  wire AES_CORE_DATAPATH__abc_16259_n3143_1;
  wire AES_CORE_DATAPATH__abc_16259_n3144;
  wire AES_CORE_DATAPATH__abc_16259_n3145;
  wire AES_CORE_DATAPATH__abc_16259_n3146;
  wire AES_CORE_DATAPATH__abc_16259_n3147;
  wire AES_CORE_DATAPATH__abc_16259_n3148_1;
  wire AES_CORE_DATAPATH__abc_16259_n3149_1;
  wire AES_CORE_DATAPATH__abc_16259_n3150;
  wire AES_CORE_DATAPATH__abc_16259_n3151;
  wire AES_CORE_DATAPATH__abc_16259_n3153;
  wire AES_CORE_DATAPATH__abc_16259_n3154_1;
  wire AES_CORE_DATAPATH__abc_16259_n3155;
  wire AES_CORE_DATAPATH__abc_16259_n3156_1;
  wire AES_CORE_DATAPATH__abc_16259_n3157;
  wire AES_CORE_DATAPATH__abc_16259_n3158_1;
  wire AES_CORE_DATAPATH__abc_16259_n3159;
  wire AES_CORE_DATAPATH__abc_16259_n3160;
  wire AES_CORE_DATAPATH__abc_16259_n3161;
  wire AES_CORE_DATAPATH__abc_16259_n3162;
  wire AES_CORE_DATAPATH__abc_16259_n3163;
  wire AES_CORE_DATAPATH__abc_16259_n3164;
  wire AES_CORE_DATAPATH__abc_16259_n3166;
  wire AES_CORE_DATAPATH__abc_16259_n3167;
  wire AES_CORE_DATAPATH__abc_16259_n3168;
  wire AES_CORE_DATAPATH__abc_16259_n3169;
  wire AES_CORE_DATAPATH__abc_16259_n3170_1;
  wire AES_CORE_DATAPATH__abc_16259_n3171;
  wire AES_CORE_DATAPATH__abc_16259_n3172_1;
  wire AES_CORE_DATAPATH__abc_16259_n3174;
  wire AES_CORE_DATAPATH__abc_16259_n3175;
  wire AES_CORE_DATAPATH__abc_16259_n3176;
  wire AES_CORE_DATAPATH__abc_16259_n3177_1;
  wire AES_CORE_DATAPATH__abc_16259_n3178_1;
  wire AES_CORE_DATAPATH__abc_16259_n3179;
  wire AES_CORE_DATAPATH__abc_16259_n3180;
  wire AES_CORE_DATAPATH__abc_16259_n3181_1;
  wire AES_CORE_DATAPATH__abc_16259_n3182;
  wire AES_CORE_DATAPATH__abc_16259_n3183_1;
  wire AES_CORE_DATAPATH__abc_16259_n3184;
  wire AES_CORE_DATAPATH__abc_16259_n3185_1;
  wire AES_CORE_DATAPATH__abc_16259_n3186;
  wire AES_CORE_DATAPATH__abc_16259_n3187_1;
  wire AES_CORE_DATAPATH__abc_16259_n3188;
  wire AES_CORE_DATAPATH__abc_16259_n3189;
  wire AES_CORE_DATAPATH__abc_16259_n3190;
  wire AES_CORE_DATAPATH__abc_16259_n3191;
  wire AES_CORE_DATAPATH__abc_16259_n3193;
  wire AES_CORE_DATAPATH__abc_16259_n3194;
  wire AES_CORE_DATAPATH__abc_16259_n3195;
  wire AES_CORE_DATAPATH__abc_16259_n3196;
  wire AES_CORE_DATAPATH__abc_16259_n3197;
  wire AES_CORE_DATAPATH__abc_16259_n3198;
  wire AES_CORE_DATAPATH__abc_16259_n3199_1;
  wire AES_CORE_DATAPATH__abc_16259_n3200;
  wire AES_CORE_DATAPATH__abc_16259_n3201_1;
  wire AES_CORE_DATAPATH__abc_16259_n3202;
  wire AES_CORE_DATAPATH__abc_16259_n3203;
  wire AES_CORE_DATAPATH__abc_16259_n3204;
  wire AES_CORE_DATAPATH__abc_16259_n3206_1;
  wire AES_CORE_DATAPATH__abc_16259_n3207_1;
  wire AES_CORE_DATAPATH__abc_16259_n3208;
  wire AES_CORE_DATAPATH__abc_16259_n3209;
  wire AES_CORE_DATAPATH__abc_16259_n3210_1;
  wire AES_CORE_DATAPATH__abc_16259_n3211;
  wire AES_CORE_DATAPATH__abc_16259_n3212_1;
  wire AES_CORE_DATAPATH__abc_16259_n3214_1;
  wire AES_CORE_DATAPATH__abc_16259_n3215;
  wire AES_CORE_DATAPATH__abc_16259_n3216_1;
  wire AES_CORE_DATAPATH__abc_16259_n3217;
  wire AES_CORE_DATAPATH__abc_16259_n3218;
  wire AES_CORE_DATAPATH__abc_16259_n3219;
  wire AES_CORE_DATAPATH__abc_16259_n3220;
  wire AES_CORE_DATAPATH__abc_16259_n3221;
  wire AES_CORE_DATAPATH__abc_16259_n3222;
  wire AES_CORE_DATAPATH__abc_16259_n3223;
  wire AES_CORE_DATAPATH__abc_16259_n3224;
  wire AES_CORE_DATAPATH__abc_16259_n3225;
  wire AES_CORE_DATAPATH__abc_16259_n3226;
  wire AES_CORE_DATAPATH__abc_16259_n3227;
  wire AES_CORE_DATAPATH__abc_16259_n3228_1;
  wire AES_CORE_DATAPATH__abc_16259_n3229;
  wire AES_CORE_DATAPATH__abc_16259_n3230_1;
  wire AES_CORE_DATAPATH__abc_16259_n3231;
  wire AES_CORE_DATAPATH__abc_16259_n3233;
  wire AES_CORE_DATAPATH__abc_16259_n3234;
  wire AES_CORE_DATAPATH__abc_16259_n3235_1;
  wire AES_CORE_DATAPATH__abc_16259_n3236_1;
  wire AES_CORE_DATAPATH__abc_16259_n3237;
  wire AES_CORE_DATAPATH__abc_16259_n3238;
  wire AES_CORE_DATAPATH__abc_16259_n3239_1;
  wire AES_CORE_DATAPATH__abc_16259_n3240;
  wire AES_CORE_DATAPATH__abc_16259_n3241_1;
  wire AES_CORE_DATAPATH__abc_16259_n3242;
  wire AES_CORE_DATAPATH__abc_16259_n3243_1;
  wire AES_CORE_DATAPATH__abc_16259_n3244;
  wire AES_CORE_DATAPATH__abc_16259_n3246;
  wire AES_CORE_DATAPATH__abc_16259_n3247;
  wire AES_CORE_DATAPATH__abc_16259_n3248;
  wire AES_CORE_DATAPATH__abc_16259_n3249;
  wire AES_CORE_DATAPATH__abc_16259_n3250;
  wire AES_CORE_DATAPATH__abc_16259_n3251;
  wire AES_CORE_DATAPATH__abc_16259_n3252;
  wire AES_CORE_DATAPATH__abc_16259_n3254;
  wire AES_CORE_DATAPATH__abc_16259_n3255;
  wire AES_CORE_DATAPATH__abc_16259_n3256;
  wire AES_CORE_DATAPATH__abc_16259_n3257_1;
  wire AES_CORE_DATAPATH__abc_16259_n3258;
  wire AES_CORE_DATAPATH__abc_16259_n3259_1;
  wire AES_CORE_DATAPATH__abc_16259_n3260;
  wire AES_CORE_DATAPATH__abc_16259_n3261;
  wire AES_CORE_DATAPATH__abc_16259_n3262;
  wire AES_CORE_DATAPATH__abc_16259_n3263;
  wire AES_CORE_DATAPATH__abc_16259_n3264_1;
  wire AES_CORE_DATAPATH__abc_16259_n3265_1;
  wire AES_CORE_DATAPATH__abc_16259_n3266;
  wire AES_CORE_DATAPATH__abc_16259_n3267;
  wire AES_CORE_DATAPATH__abc_16259_n3268_1;
  wire AES_CORE_DATAPATH__abc_16259_n3269;
  wire AES_CORE_DATAPATH__abc_16259_n3270_1;
  wire AES_CORE_DATAPATH__abc_16259_n3271;
  wire AES_CORE_DATAPATH__abc_16259_n3273;
  wire AES_CORE_DATAPATH__abc_16259_n3274_1;
  wire AES_CORE_DATAPATH__abc_16259_n3275;
  wire AES_CORE_DATAPATH__abc_16259_n3276;
  wire AES_CORE_DATAPATH__abc_16259_n3277;
  wire AES_CORE_DATAPATH__abc_16259_n3278;
  wire AES_CORE_DATAPATH__abc_16259_n3279;
  wire AES_CORE_DATAPATH__abc_16259_n3280;
  wire AES_CORE_DATAPATH__abc_16259_n3281;
  wire AES_CORE_DATAPATH__abc_16259_n3282;
  wire AES_CORE_DATAPATH__abc_16259_n3283;
  wire AES_CORE_DATAPATH__abc_16259_n3284;
  wire AES_CORE_DATAPATH__abc_16259_n3286_1;
  wire AES_CORE_DATAPATH__abc_16259_n3287;
  wire AES_CORE_DATAPATH__abc_16259_n3288_1;
  wire AES_CORE_DATAPATH__abc_16259_n3289;
  wire AES_CORE_DATAPATH__abc_16259_n3290;
  wire AES_CORE_DATAPATH__abc_16259_n3291;
  wire AES_CORE_DATAPATH__abc_16259_n3292;
  wire AES_CORE_DATAPATH__abc_16259_n3294_1;
  wire AES_CORE_DATAPATH__abc_16259_n3295;
  wire AES_CORE_DATAPATH__abc_16259_n3296;
  wire AES_CORE_DATAPATH__abc_16259_n3297_1;
  wire AES_CORE_DATAPATH__abc_16259_n3298;
  wire AES_CORE_DATAPATH__abc_16259_n3299_1;
  wire AES_CORE_DATAPATH__abc_16259_n3300;
  wire AES_CORE_DATAPATH__abc_16259_n3301_1;
  wire AES_CORE_DATAPATH__abc_16259_n3302;
  wire AES_CORE_DATAPATH__abc_16259_n3303_1;
  wire AES_CORE_DATAPATH__abc_16259_n3304;
  wire AES_CORE_DATAPATH__abc_16259_n3305;
  wire AES_CORE_DATAPATH__abc_16259_n3306;
  wire AES_CORE_DATAPATH__abc_16259_n3307;
  wire AES_CORE_DATAPATH__abc_16259_n3308;
  wire AES_CORE_DATAPATH__abc_16259_n3309;
  wire AES_CORE_DATAPATH__abc_16259_n3310;
  wire AES_CORE_DATAPATH__abc_16259_n3311;
  wire AES_CORE_DATAPATH__abc_16259_n3313;
  wire AES_CORE_DATAPATH__abc_16259_n3314;
  wire AES_CORE_DATAPATH__abc_16259_n3315_1;
  wire AES_CORE_DATAPATH__abc_16259_n3316;
  wire AES_CORE_DATAPATH__abc_16259_n3317_1;
  wire AES_CORE_DATAPATH__abc_16259_n3318;
  wire AES_CORE_DATAPATH__abc_16259_n3319;
  wire AES_CORE_DATAPATH__abc_16259_n3320;
  wire AES_CORE_DATAPATH__abc_16259_n3321;
  wire AES_CORE_DATAPATH__abc_16259_n3322_1;
  wire AES_CORE_DATAPATH__abc_16259_n3323_1;
  wire AES_CORE_DATAPATH__abc_16259_n3324;
  wire AES_CORE_DATAPATH__abc_16259_n3326_1;
  wire AES_CORE_DATAPATH__abc_16259_n3327;
  wire AES_CORE_DATAPATH__abc_16259_n3328_1;
  wire AES_CORE_DATAPATH__abc_16259_n3329;
  wire AES_CORE_DATAPATH__abc_16259_n3330_1;
  wire AES_CORE_DATAPATH__abc_16259_n3331;
  wire AES_CORE_DATAPATH__abc_16259_n3332_1;
  wire AES_CORE_DATAPATH__abc_16259_n3334;
  wire AES_CORE_DATAPATH__abc_16259_n3335;
  wire AES_CORE_DATAPATH__abc_16259_n3336;
  wire AES_CORE_DATAPATH__abc_16259_n3337;
  wire AES_CORE_DATAPATH__abc_16259_n3338;
  wire AES_CORE_DATAPATH__abc_16259_n3339;
  wire AES_CORE_DATAPATH__abc_16259_n3340;
  wire AES_CORE_DATAPATH__abc_16259_n3341;
  wire AES_CORE_DATAPATH__abc_16259_n3342;
  wire AES_CORE_DATAPATH__abc_16259_n3343;
  wire AES_CORE_DATAPATH__abc_16259_n3344_1;
  wire AES_CORE_DATAPATH__abc_16259_n3345;
  wire AES_CORE_DATAPATH__abc_16259_n3346_1;
  wire AES_CORE_DATAPATH__abc_16259_n3347;
  wire AES_CORE_DATAPATH__abc_16259_n3348;
  wire AES_CORE_DATAPATH__abc_16259_n3349;
  wire AES_CORE_DATAPATH__abc_16259_n3350;
  wire AES_CORE_DATAPATH__abc_16259_n3351_1;
  wire AES_CORE_DATAPATH__abc_16259_n3353;
  wire AES_CORE_DATAPATH__abc_16259_n3354;
  wire AES_CORE_DATAPATH__abc_16259_n3355_1;
  wire AES_CORE_DATAPATH__abc_16259_n3356;
  wire AES_CORE_DATAPATH__abc_16259_n3357_1;
  wire AES_CORE_DATAPATH__abc_16259_n3358;
  wire AES_CORE_DATAPATH__abc_16259_n3359_1;
  wire AES_CORE_DATAPATH__abc_16259_n3360;
  wire AES_CORE_DATAPATH__abc_16259_n3361_1;
  wire AES_CORE_DATAPATH__abc_16259_n3362;
  wire AES_CORE_DATAPATH__abc_16259_n3363;
  wire AES_CORE_DATAPATH__abc_16259_n3364;
  wire AES_CORE_DATAPATH__abc_16259_n3366;
  wire AES_CORE_DATAPATH__abc_16259_n3367;
  wire AES_CORE_DATAPATH__abc_16259_n3368;
  wire AES_CORE_DATAPATH__abc_16259_n3369;
  wire AES_CORE_DATAPATH__abc_16259_n3370;
  wire AES_CORE_DATAPATH__abc_16259_n3371;
  wire AES_CORE_DATAPATH__abc_16259_n3372;
  wire AES_CORE_DATAPATH__abc_16259_n3374;
  wire AES_CORE_DATAPATH__abc_16259_n3375_1;
  wire AES_CORE_DATAPATH__abc_16259_n3376;
  wire AES_CORE_DATAPATH__abc_16259_n3377;
  wire AES_CORE_DATAPATH__abc_16259_n3378;
  wire AES_CORE_DATAPATH__abc_16259_n3379;
  wire AES_CORE_DATAPATH__abc_16259_n3380_1;
  wire AES_CORE_DATAPATH__abc_16259_n3381_1;
  wire AES_CORE_DATAPATH__abc_16259_n3382;
  wire AES_CORE_DATAPATH__abc_16259_n3383;
  wire AES_CORE_DATAPATH__abc_16259_n3384_1;
  wire AES_CORE_DATAPATH__abc_16259_n3385;
  wire AES_CORE_DATAPATH__abc_16259_n3386_1;
  wire AES_CORE_DATAPATH__abc_16259_n3387;
  wire AES_CORE_DATAPATH__abc_16259_n3388_1;
  wire AES_CORE_DATAPATH__abc_16259_n3389;
  wire AES_CORE_DATAPATH__abc_16259_n3390_1;
  wire AES_CORE_DATAPATH__abc_16259_n3391;
  wire AES_CORE_DATAPATH__abc_16259_n3393;
  wire AES_CORE_DATAPATH__abc_16259_n3394;
  wire AES_CORE_DATAPATH__abc_16259_n3395;
  wire AES_CORE_DATAPATH__abc_16259_n3396;
  wire AES_CORE_DATAPATH__abc_16259_n3397;
  wire AES_CORE_DATAPATH__abc_16259_n3398;
  wire AES_CORE_DATAPATH__abc_16259_n3399;
  wire AES_CORE_DATAPATH__abc_16259_n3400;
  wire AES_CORE_DATAPATH__abc_16259_n3401;
  wire AES_CORE_DATAPATH__abc_16259_n3402_1;
  wire AES_CORE_DATAPATH__abc_16259_n3403;
  wire AES_CORE_DATAPATH__abc_16259_n3404_1;
  wire AES_CORE_DATAPATH__abc_16259_n3406;
  wire AES_CORE_DATAPATH__abc_16259_n3407;
  wire AES_CORE_DATAPATH__abc_16259_n3408;
  wire AES_CORE_DATAPATH__abc_16259_n3409_1;
  wire AES_CORE_DATAPATH__abc_16259_n3410_1;
  wire AES_CORE_DATAPATH__abc_16259_n3411;
  wire AES_CORE_DATAPATH__abc_16259_n3412;
  wire AES_CORE_DATAPATH__abc_16259_n3414;
  wire AES_CORE_DATAPATH__abc_16259_n3415_1;
  wire AES_CORE_DATAPATH__abc_16259_n3416;
  wire AES_CORE_DATAPATH__abc_16259_n3417_1;
  wire AES_CORE_DATAPATH__abc_16259_n3418;
  wire AES_CORE_DATAPATH__abc_16259_n3419_1;
  wire AES_CORE_DATAPATH__abc_16259_n3420;
  wire AES_CORE_DATAPATH__abc_16259_n3421;
  wire AES_CORE_DATAPATH__abc_16259_n3422;
  wire AES_CORE_DATAPATH__abc_16259_n3423;
  wire AES_CORE_DATAPATH__abc_16259_n3424;
  wire AES_CORE_DATAPATH__abc_16259_n3425;
  wire AES_CORE_DATAPATH__abc_16259_n3426;
  wire AES_CORE_DATAPATH__abc_16259_n3427;
  wire AES_CORE_DATAPATH__abc_16259_n3428;
  wire AES_CORE_DATAPATH__abc_16259_n3429;
  wire AES_CORE_DATAPATH__abc_16259_n3430;
  wire AES_CORE_DATAPATH__abc_16259_n3431_1;
  wire AES_CORE_DATAPATH__abc_16259_n3433_1;
  wire AES_CORE_DATAPATH__abc_16259_n3434;
  wire AES_CORE_DATAPATH__abc_16259_n3435;
  wire AES_CORE_DATAPATH__abc_16259_n3436;
  wire AES_CORE_DATAPATH__abc_16259_n3437;
  wire AES_CORE_DATAPATH__abc_16259_n3438_1;
  wire AES_CORE_DATAPATH__abc_16259_n3439_1;
  wire AES_CORE_DATAPATH__abc_16259_n3440;
  wire AES_CORE_DATAPATH__abc_16259_n3441;
  wire AES_CORE_DATAPATH__abc_16259_n3442_1;
  wire AES_CORE_DATAPATH__abc_16259_n3443;
  wire AES_CORE_DATAPATH__abc_16259_n3444_1;
  wire AES_CORE_DATAPATH__abc_16259_n3446_1;
  wire AES_CORE_DATAPATH__abc_16259_n3447;
  wire AES_CORE_DATAPATH__abc_16259_n3448_1;
  wire AES_CORE_DATAPATH__abc_16259_n3449;
  wire AES_CORE_DATAPATH__abc_16259_n3450;
  wire AES_CORE_DATAPATH__abc_16259_n3451;
  wire AES_CORE_DATAPATH__abc_16259_n3452;
  wire AES_CORE_DATAPATH__abc_16259_n3454;
  wire AES_CORE_DATAPATH__abc_16259_n3455;
  wire AES_CORE_DATAPATH__abc_16259_n3456;
  wire AES_CORE_DATAPATH__abc_16259_n3457;
  wire AES_CORE_DATAPATH__abc_16259_n3458;
  wire AES_CORE_DATAPATH__abc_16259_n3459;
  wire AES_CORE_DATAPATH__abc_16259_n3460_1;
  wire AES_CORE_DATAPATH__abc_16259_n3461;
  wire AES_CORE_DATAPATH__abc_16259_n3462_1;
  wire AES_CORE_DATAPATH__abc_16259_n3463;
  wire AES_CORE_DATAPATH__abc_16259_n3464;
  wire AES_CORE_DATAPATH__abc_16259_n3465;
  wire AES_CORE_DATAPATH__abc_16259_n3466;
  wire AES_CORE_DATAPATH__abc_16259_n3467_1;
  wire AES_CORE_DATAPATH__abc_16259_n3468_1;
  wire AES_CORE_DATAPATH__abc_16259_n3469;
  wire AES_CORE_DATAPATH__abc_16259_n3470;
  wire AES_CORE_DATAPATH__abc_16259_n3471_1;
  wire AES_CORE_DATAPATH__abc_16259_n3473_1;
  wire AES_CORE_DATAPATH__abc_16259_n3474;
  wire AES_CORE_DATAPATH__abc_16259_n3475_1;
  wire AES_CORE_DATAPATH__abc_16259_n3476;
  wire AES_CORE_DATAPATH__abc_16259_n3477_1;
  wire AES_CORE_DATAPATH__abc_16259_n3478;
  wire AES_CORE_DATAPATH__abc_16259_n3479;
  wire AES_CORE_DATAPATH__abc_16259_n3480;
  wire AES_CORE_DATAPATH__abc_16259_n3481;
  wire AES_CORE_DATAPATH__abc_16259_n3482;
  wire AES_CORE_DATAPATH__abc_16259_n3483;
  wire AES_CORE_DATAPATH__abc_16259_n3484;
  wire AES_CORE_DATAPATH__abc_16259_n3486;
  wire AES_CORE_DATAPATH__abc_16259_n3487;
  wire AES_CORE_DATAPATH__abc_16259_n3488;
  wire AES_CORE_DATAPATH__abc_16259_n3489_1;
  wire AES_CORE_DATAPATH__abc_16259_n3490;
  wire AES_CORE_DATAPATH__abc_16259_n3491_1;
  wire AES_CORE_DATAPATH__abc_16259_n3492;
  wire AES_CORE_DATAPATH__abc_16259_n3494;
  wire AES_CORE_DATAPATH__abc_16259_n3495;
  wire AES_CORE_DATAPATH__abc_16259_n3496_1;
  wire AES_CORE_DATAPATH__abc_16259_n3497_1;
  wire AES_CORE_DATAPATH__abc_16259_n3498;
  wire AES_CORE_DATAPATH__abc_16259_n3499;
  wire AES_CORE_DATAPATH__abc_16259_n3500_1;
  wire AES_CORE_DATAPATH__abc_16259_n3501;
  wire AES_CORE_DATAPATH__abc_16259_n3502_1;
  wire AES_CORE_DATAPATH__abc_16259_n3503;
  wire AES_CORE_DATAPATH__abc_16259_n3504_1;
  wire AES_CORE_DATAPATH__abc_16259_n3505;
  wire AES_CORE_DATAPATH__abc_16259_n3506_1;
  wire AES_CORE_DATAPATH__abc_16259_n3507;
  wire AES_CORE_DATAPATH__abc_16259_n3508;
  wire AES_CORE_DATAPATH__abc_16259_n3509;
  wire AES_CORE_DATAPATH__abc_16259_n3510;
  wire AES_CORE_DATAPATH__abc_16259_n3511;
  wire AES_CORE_DATAPATH__abc_16259_n3513;
  wire AES_CORE_DATAPATH__abc_16259_n3514;
  wire AES_CORE_DATAPATH__abc_16259_n3515;
  wire AES_CORE_DATAPATH__abc_16259_n3516;
  wire AES_CORE_DATAPATH__abc_16259_n3517;
  wire AES_CORE_DATAPATH__abc_16259_n3518_1;
  wire AES_CORE_DATAPATH__abc_16259_n3519;
  wire AES_CORE_DATAPATH__abc_16259_n3520_1;
  wire AES_CORE_DATAPATH__abc_16259_n3521;
  wire AES_CORE_DATAPATH__abc_16259_n3522;
  wire AES_CORE_DATAPATH__abc_16259_n3523;
  wire AES_CORE_DATAPATH__abc_16259_n3524;
  wire AES_CORE_DATAPATH__abc_16259_n3526_1;
  wire AES_CORE_DATAPATH__abc_16259_n3527;
  wire AES_CORE_DATAPATH__abc_16259_n3528;
  wire AES_CORE_DATAPATH__abc_16259_n3529_1;
  wire AES_CORE_DATAPATH__abc_16259_n3530;
  wire AES_CORE_DATAPATH__abc_16259_n3531_1;
  wire AES_CORE_DATAPATH__abc_16259_n3532;
  wire AES_CORE_DATAPATH__abc_16259_n3534;
  wire AES_CORE_DATAPATH__abc_16259_n3535_1;
  wire AES_CORE_DATAPATH__abc_16259_n3536;
  wire AES_CORE_DATAPATH__abc_16259_n3537;
  wire AES_CORE_DATAPATH__abc_16259_n3538;
  wire AES_CORE_DATAPATH__abc_16259_n3539;
  wire AES_CORE_DATAPATH__abc_16259_n3540;
  wire AES_CORE_DATAPATH__abc_16259_n3541;
  wire AES_CORE_DATAPATH__abc_16259_n3542;
  wire AES_CORE_DATAPATH__abc_16259_n3543;
  wire AES_CORE_DATAPATH__abc_16259_n3544;
  wire AES_CORE_DATAPATH__abc_16259_n3545;
  wire AES_CORE_DATAPATH__abc_16259_n3546;
  wire AES_CORE_DATAPATH__abc_16259_n3547_1;
  wire AES_CORE_DATAPATH__abc_16259_n3548;
  wire AES_CORE_DATAPATH__abc_16259_n3549_1;
  wire AES_CORE_DATAPATH__abc_16259_n3550;
  wire AES_CORE_DATAPATH__abc_16259_n3551;
  wire AES_CORE_DATAPATH__abc_16259_n3553;
  wire AES_CORE_DATAPATH__abc_16259_n3554_1;
  wire AES_CORE_DATAPATH__abc_16259_n3555_1;
  wire AES_CORE_DATAPATH__abc_16259_n3556;
  wire AES_CORE_DATAPATH__abc_16259_n3557;
  wire AES_CORE_DATAPATH__abc_16259_n3558_1;
  wire AES_CORE_DATAPATH__abc_16259_n3559;
  wire AES_CORE_DATAPATH__abc_16259_n3560_1;
  wire AES_CORE_DATAPATH__abc_16259_n3561;
  wire AES_CORE_DATAPATH__abc_16259_n3562_1;
  wire AES_CORE_DATAPATH__abc_16259_n3563;
  wire AES_CORE_DATAPATH__abc_16259_n3564_1;
  wire AES_CORE_DATAPATH__abc_16259_n3566;
  wire AES_CORE_DATAPATH__abc_16259_n3567;
  wire AES_CORE_DATAPATH__abc_16259_n3568;
  wire AES_CORE_DATAPATH__abc_16259_n3569;
  wire AES_CORE_DATAPATH__abc_16259_n3570;
  wire AES_CORE_DATAPATH__abc_16259_n3571;
  wire AES_CORE_DATAPATH__abc_16259_n3572;
  wire AES_CORE_DATAPATH__abc_16259_n3574;
  wire AES_CORE_DATAPATH__abc_16259_n3575;
  wire AES_CORE_DATAPATH__abc_16259_n3576_1;
  wire AES_CORE_DATAPATH__abc_16259_n3577;
  wire AES_CORE_DATAPATH__abc_16259_n3578_1;
  wire AES_CORE_DATAPATH__abc_16259_n3579;
  wire AES_CORE_DATAPATH__abc_16259_n3580;
  wire AES_CORE_DATAPATH__abc_16259_n3581;
  wire AES_CORE_DATAPATH__abc_16259_n3582;
  wire AES_CORE_DATAPATH__abc_16259_n3583_1;
  wire AES_CORE_DATAPATH__abc_16259_n3584_1;
  wire AES_CORE_DATAPATH__abc_16259_n3585;
  wire AES_CORE_DATAPATH__abc_16259_n3586;
  wire AES_CORE_DATAPATH__abc_16259_n3587_1;
  wire AES_CORE_DATAPATH__abc_16259_n3588;
  wire AES_CORE_DATAPATH__abc_16259_n3589_1;
  wire AES_CORE_DATAPATH__abc_16259_n3590;
  wire AES_CORE_DATAPATH__abc_16259_n3591_1;
  wire AES_CORE_DATAPATH__abc_16259_n3593_1;
  wire AES_CORE_DATAPATH__abc_16259_n3594;
  wire AES_CORE_DATAPATH__abc_16259_n3595;
  wire AES_CORE_DATAPATH__abc_16259_n3596;
  wire AES_CORE_DATAPATH__abc_16259_n3597;
  wire AES_CORE_DATAPATH__abc_16259_n3598;
  wire AES_CORE_DATAPATH__abc_16259_n3599;
  wire AES_CORE_DATAPATH__abc_16259_n3600;
  wire AES_CORE_DATAPATH__abc_16259_n3601;
  wire AES_CORE_DATAPATH__abc_16259_n3602;
  wire AES_CORE_DATAPATH__abc_16259_n3603;
  wire AES_CORE_DATAPATH__abc_16259_n3604;
  wire AES_CORE_DATAPATH__abc_16259_n3606;
  wire AES_CORE_DATAPATH__abc_16259_n3607_1;
  wire AES_CORE_DATAPATH__abc_16259_n3608;
  wire AES_CORE_DATAPATH__abc_16259_n3609;
  wire AES_CORE_DATAPATH__abc_16259_n3610;
  wire AES_CORE_DATAPATH__abc_16259_n3611;
  wire AES_CORE_DATAPATH__abc_16259_n3612_1;
  wire AES_CORE_DATAPATH__abc_16259_n3614;
  wire AES_CORE_DATAPATH__abc_16259_n3615;
  wire AES_CORE_DATAPATH__abc_16259_n3616_1;
  wire AES_CORE_DATAPATH__abc_16259_n3617;
  wire AES_CORE_DATAPATH__abc_16259_n3618_1;
  wire AES_CORE_DATAPATH__abc_16259_n3619;
  wire AES_CORE_DATAPATH__abc_16259_n3620_1;
  wire AES_CORE_DATAPATH__abc_16259_n3621;
  wire AES_CORE_DATAPATH__abc_16259_n3622_1;
  wire AES_CORE_DATAPATH__abc_16259_n3623;
  wire AES_CORE_DATAPATH__abc_16259_n3624;
  wire AES_CORE_DATAPATH__abc_16259_n3625;
  wire AES_CORE_DATAPATH__abc_16259_n3626;
  wire AES_CORE_DATAPATH__abc_16259_n3627;
  wire AES_CORE_DATAPATH__abc_16259_n3628;
  wire AES_CORE_DATAPATH__abc_16259_n3629;
  wire AES_CORE_DATAPATH__abc_16259_n3630;
  wire AES_CORE_DATAPATH__abc_16259_n3631;
  wire AES_CORE_DATAPATH__abc_16259_n3633;
  wire AES_CORE_DATAPATH__abc_16259_n3634_1;
  wire AES_CORE_DATAPATH__abc_16259_n3635;
  wire AES_CORE_DATAPATH__abc_16259_n3636_1;
  wire AES_CORE_DATAPATH__abc_16259_n3637;
  wire AES_CORE_DATAPATH__abc_16259_n3638;
  wire AES_CORE_DATAPATH__abc_16259_n3639;
  wire AES_CORE_DATAPATH__abc_16259_n3640;
  wire AES_CORE_DATAPATH__abc_16259_n3641_1;
  wire AES_CORE_DATAPATH__abc_16259_n3642_1;
  wire AES_CORE_DATAPATH__abc_16259_n3643;
  wire AES_CORE_DATAPATH__abc_16259_n3644;
  wire AES_CORE_DATAPATH__abc_16259_n3646;
  wire AES_CORE_DATAPATH__abc_16259_n3647_1;
  wire AES_CORE_DATAPATH__abc_16259_n3648;
  wire AES_CORE_DATAPATH__abc_16259_n3649_1;
  wire AES_CORE_DATAPATH__abc_16259_n3650;
  wire AES_CORE_DATAPATH__abc_16259_n3651_1;
  wire AES_CORE_DATAPATH__abc_16259_n3652;
  wire AES_CORE_DATAPATH__abc_16259_n3654;
  wire AES_CORE_DATAPATH__abc_16259_n3655;
  wire AES_CORE_DATAPATH__abc_16259_n3656;
  wire AES_CORE_DATAPATH__abc_16259_n3657;
  wire AES_CORE_DATAPATH__abc_16259_n3658;
  wire AES_CORE_DATAPATH__abc_16259_n3659;
  wire AES_CORE_DATAPATH__abc_16259_n3660;
  wire AES_CORE_DATAPATH__abc_16259_n3661;
  wire AES_CORE_DATAPATH__abc_16259_n3662;
  wire AES_CORE_DATAPATH__abc_16259_n3663_1;
  wire AES_CORE_DATAPATH__abc_16259_n3664;
  wire AES_CORE_DATAPATH__abc_16259_n3665_1;
  wire AES_CORE_DATAPATH__abc_16259_n3666;
  wire AES_CORE_DATAPATH__abc_16259_n3667;
  wire AES_CORE_DATAPATH__abc_16259_n3668;
  wire AES_CORE_DATAPATH__abc_16259_n3669;
  wire AES_CORE_DATAPATH__abc_16259_n3670_1;
  wire AES_CORE_DATAPATH__abc_16259_n3671_1;
  wire AES_CORE_DATAPATH__abc_16259_n3673_1;
  wire AES_CORE_DATAPATH__abc_16259_n3674;
  wire AES_CORE_DATAPATH__abc_16259_n3675;
  wire AES_CORE_DATAPATH__abc_16259_n3676;
  wire AES_CORE_DATAPATH__abc_16259_n3677;
  wire AES_CORE_DATAPATH__abc_16259_n3678_1;
  wire AES_CORE_DATAPATH__abc_16259_n3679_1;
  wire AES_CORE_DATAPATH__abc_16259_n3680;
  wire AES_CORE_DATAPATH__abc_16259_n3681_1;
  wire AES_CORE_DATAPATH__abc_16259_n3682;
  wire AES_CORE_DATAPATH__abc_16259_n3683;
  wire AES_CORE_DATAPATH__abc_16259_n3684;
  wire AES_CORE_DATAPATH__abc_16259_n3686_1;
  wire AES_CORE_DATAPATH__abc_16259_n3687_1;
  wire AES_CORE_DATAPATH__abc_16259_n3688;
  wire AES_CORE_DATAPATH__abc_16259_n3689_1;
  wire AES_CORE_DATAPATH__abc_16259_n3690;
  wire AES_CORE_DATAPATH__abc_16259_n3691;
  wire AES_CORE_DATAPATH__abc_16259_n3692;
  wire AES_CORE_DATAPATH__abc_16259_n3694_1;
  wire AES_CORE_DATAPATH__abc_16259_n3695_1;
  wire AES_CORE_DATAPATH__abc_16259_n3696;
  wire AES_CORE_DATAPATH__abc_16259_n3697_1;
  wire AES_CORE_DATAPATH__abc_16259_n3698;
  wire AES_CORE_DATAPATH__abc_16259_n3699;
  wire AES_CORE_DATAPATH__abc_16259_n3700;
  wire AES_CORE_DATAPATH__abc_16259_n3701;
  wire AES_CORE_DATAPATH__abc_16259_n3702_1;
  wire AES_CORE_DATAPATH__abc_16259_n3703_1;
  wire AES_CORE_DATAPATH__abc_16259_n3704;
  wire AES_CORE_DATAPATH__abc_16259_n3705_1;
  wire AES_CORE_DATAPATH__abc_16259_n3706;
  wire AES_CORE_DATAPATH__abc_16259_n3707;
  wire AES_CORE_DATAPATH__abc_16259_n3708;
  wire AES_CORE_DATAPATH__abc_16259_n3709;
  wire AES_CORE_DATAPATH__abc_16259_n3710_1;
  wire AES_CORE_DATAPATH__abc_16259_n3711_1;
  wire AES_CORE_DATAPATH__abc_16259_n3713_1;
  wire AES_CORE_DATAPATH__abc_16259_n3714;
  wire AES_CORE_DATAPATH__abc_16259_n3715;
  wire AES_CORE_DATAPATH__abc_16259_n3716;
  wire AES_CORE_DATAPATH__abc_16259_n3717;
  wire AES_CORE_DATAPATH__abc_16259_n3718_1;
  wire AES_CORE_DATAPATH__abc_16259_n3719_1;
  wire AES_CORE_DATAPATH__abc_16259_n3720;
  wire AES_CORE_DATAPATH__abc_16259_n3721_1;
  wire AES_CORE_DATAPATH__abc_16259_n3722;
  wire AES_CORE_DATAPATH__abc_16259_n3723;
  wire AES_CORE_DATAPATH__abc_16259_n3724;
  wire AES_CORE_DATAPATH__abc_16259_n3726_1;
  wire AES_CORE_DATAPATH__abc_16259_n3727_1;
  wire AES_CORE_DATAPATH__abc_16259_n3728;
  wire AES_CORE_DATAPATH__abc_16259_n3729_1;
  wire AES_CORE_DATAPATH__abc_16259_n3730;
  wire AES_CORE_DATAPATH__abc_16259_n3731;
  wire AES_CORE_DATAPATH__abc_16259_n3732;
  wire AES_CORE_DATAPATH__abc_16259_n3734_1;
  wire AES_CORE_DATAPATH__abc_16259_n3735_1;
  wire AES_CORE_DATAPATH__abc_16259_n3736;
  wire AES_CORE_DATAPATH__abc_16259_n3737_1;
  wire AES_CORE_DATAPATH__abc_16259_n3738;
  wire AES_CORE_DATAPATH__abc_16259_n3739;
  wire AES_CORE_DATAPATH__abc_16259_n3740;
  wire AES_CORE_DATAPATH__abc_16259_n3741;
  wire AES_CORE_DATAPATH__abc_16259_n3742_1;
  wire AES_CORE_DATAPATH__abc_16259_n3743_1;
  wire AES_CORE_DATAPATH__abc_16259_n3744;
  wire AES_CORE_DATAPATH__abc_16259_n3745_1;
  wire AES_CORE_DATAPATH__abc_16259_n3746;
  wire AES_CORE_DATAPATH__abc_16259_n3747;
  wire AES_CORE_DATAPATH__abc_16259_n3748;
  wire AES_CORE_DATAPATH__abc_16259_n3749;
  wire AES_CORE_DATAPATH__abc_16259_n3750_1;
  wire AES_CORE_DATAPATH__abc_16259_n3751_1;
  wire AES_CORE_DATAPATH__abc_16259_n3753_1;
  wire AES_CORE_DATAPATH__abc_16259_n3754;
  wire AES_CORE_DATAPATH__abc_16259_n3755;
  wire AES_CORE_DATAPATH__abc_16259_n3756;
  wire AES_CORE_DATAPATH__abc_16259_n3757;
  wire AES_CORE_DATAPATH__abc_16259_n3758_1;
  wire AES_CORE_DATAPATH__abc_16259_n3759_1;
  wire AES_CORE_DATAPATH__abc_16259_n3760;
  wire AES_CORE_DATAPATH__abc_16259_n3761_1;
  wire AES_CORE_DATAPATH__abc_16259_n3762;
  wire AES_CORE_DATAPATH__abc_16259_n3763;
  wire AES_CORE_DATAPATH__abc_16259_n3764;
  wire AES_CORE_DATAPATH__abc_16259_n3766_1;
  wire AES_CORE_DATAPATH__abc_16259_n3767_1;
  wire AES_CORE_DATAPATH__abc_16259_n3768;
  wire AES_CORE_DATAPATH__abc_16259_n3769_1;
  wire AES_CORE_DATAPATH__abc_16259_n3770;
  wire AES_CORE_DATAPATH__abc_16259_n3771;
  wire AES_CORE_DATAPATH__abc_16259_n3772;
  wire AES_CORE_DATAPATH__abc_16259_n3774_1;
  wire AES_CORE_DATAPATH__abc_16259_n3775_1;
  wire AES_CORE_DATAPATH__abc_16259_n3776;
  wire AES_CORE_DATAPATH__abc_16259_n3777_1;
  wire AES_CORE_DATAPATH__abc_16259_n3778;
  wire AES_CORE_DATAPATH__abc_16259_n3779;
  wire AES_CORE_DATAPATH__abc_16259_n3780;
  wire AES_CORE_DATAPATH__abc_16259_n3781;
  wire AES_CORE_DATAPATH__abc_16259_n3782_1;
  wire AES_CORE_DATAPATH__abc_16259_n3783_1;
  wire AES_CORE_DATAPATH__abc_16259_n3784;
  wire AES_CORE_DATAPATH__abc_16259_n3785_1;
  wire AES_CORE_DATAPATH__abc_16259_n3786;
  wire AES_CORE_DATAPATH__abc_16259_n3787;
  wire AES_CORE_DATAPATH__abc_16259_n3788;
  wire AES_CORE_DATAPATH__abc_16259_n3789;
  wire AES_CORE_DATAPATH__abc_16259_n3790_1;
  wire AES_CORE_DATAPATH__abc_16259_n3791_1;
  wire AES_CORE_DATAPATH__abc_16259_n3793_1;
  wire AES_CORE_DATAPATH__abc_16259_n3794;
  wire AES_CORE_DATAPATH__abc_16259_n3795;
  wire AES_CORE_DATAPATH__abc_16259_n3796;
  wire AES_CORE_DATAPATH__abc_16259_n3797;
  wire AES_CORE_DATAPATH__abc_16259_n3798_1;
  wire AES_CORE_DATAPATH__abc_16259_n3799_1;
  wire AES_CORE_DATAPATH__abc_16259_n3800;
  wire AES_CORE_DATAPATH__abc_16259_n3801_1;
  wire AES_CORE_DATAPATH__abc_16259_n3802;
  wire AES_CORE_DATAPATH__abc_16259_n3803;
  wire AES_CORE_DATAPATH__abc_16259_n3804;
  wire AES_CORE_DATAPATH__abc_16259_n3806_1;
  wire AES_CORE_DATAPATH__abc_16259_n3807_1;
  wire AES_CORE_DATAPATH__abc_16259_n3808;
  wire AES_CORE_DATAPATH__abc_16259_n3809_1;
  wire AES_CORE_DATAPATH__abc_16259_n3810;
  wire AES_CORE_DATAPATH__abc_16259_n3811;
  wire AES_CORE_DATAPATH__abc_16259_n3812;
  wire AES_CORE_DATAPATH__abc_16259_n3814_1;
  wire AES_CORE_DATAPATH__abc_16259_n3815_1;
  wire AES_CORE_DATAPATH__abc_16259_n3816;
  wire AES_CORE_DATAPATH__abc_16259_n3817_1;
  wire AES_CORE_DATAPATH__abc_16259_n3818;
  wire AES_CORE_DATAPATH__abc_16259_n3819;
  wire AES_CORE_DATAPATH__abc_16259_n3820;
  wire AES_CORE_DATAPATH__abc_16259_n3821;
  wire AES_CORE_DATAPATH__abc_16259_n3822_1;
  wire AES_CORE_DATAPATH__abc_16259_n3823_1;
  wire AES_CORE_DATAPATH__abc_16259_n3824;
  wire AES_CORE_DATAPATH__abc_16259_n3825_1;
  wire AES_CORE_DATAPATH__abc_16259_n3826;
  wire AES_CORE_DATAPATH__abc_16259_n3827;
  wire AES_CORE_DATAPATH__abc_16259_n3828;
  wire AES_CORE_DATAPATH__abc_16259_n3829;
  wire AES_CORE_DATAPATH__abc_16259_n3830_1;
  wire AES_CORE_DATAPATH__abc_16259_n3831_1;
  wire AES_CORE_DATAPATH__abc_16259_n3833_1;
  wire AES_CORE_DATAPATH__abc_16259_n3834;
  wire AES_CORE_DATAPATH__abc_16259_n3835;
  wire AES_CORE_DATAPATH__abc_16259_n3836;
  wire AES_CORE_DATAPATH__abc_16259_n3837;
  wire AES_CORE_DATAPATH__abc_16259_n3838_1;
  wire AES_CORE_DATAPATH__abc_16259_n3839_1;
  wire AES_CORE_DATAPATH__abc_16259_n3840;
  wire AES_CORE_DATAPATH__abc_16259_n3841_1;
  wire AES_CORE_DATAPATH__abc_16259_n3842;
  wire AES_CORE_DATAPATH__abc_16259_n3843;
  wire AES_CORE_DATAPATH__abc_16259_n3844;
  wire AES_CORE_DATAPATH__abc_16259_n3846_1;
  wire AES_CORE_DATAPATH__abc_16259_n3847_1;
  wire AES_CORE_DATAPATH__abc_16259_n3848;
  wire AES_CORE_DATAPATH__abc_16259_n3849_1;
  wire AES_CORE_DATAPATH__abc_16259_n3850;
  wire AES_CORE_DATAPATH__abc_16259_n3851;
  wire AES_CORE_DATAPATH__abc_16259_n3852;
  wire AES_CORE_DATAPATH__abc_16259_n3854_1;
  wire AES_CORE_DATAPATH__abc_16259_n3855_1;
  wire AES_CORE_DATAPATH__abc_16259_n3856;
  wire AES_CORE_DATAPATH__abc_16259_n3857_1;
  wire AES_CORE_DATAPATH__abc_16259_n3858;
  wire AES_CORE_DATAPATH__abc_16259_n3859;
  wire AES_CORE_DATAPATH__abc_16259_n3860;
  wire AES_CORE_DATAPATH__abc_16259_n3861;
  wire AES_CORE_DATAPATH__abc_16259_n3862_1;
  wire AES_CORE_DATAPATH__abc_16259_n3863_1;
  wire AES_CORE_DATAPATH__abc_16259_n3864;
  wire AES_CORE_DATAPATH__abc_16259_n3865_1;
  wire AES_CORE_DATAPATH__abc_16259_n3866;
  wire AES_CORE_DATAPATH__abc_16259_n3867;
  wire AES_CORE_DATAPATH__abc_16259_n3868;
  wire AES_CORE_DATAPATH__abc_16259_n3869;
  wire AES_CORE_DATAPATH__abc_16259_n3870_1;
  wire AES_CORE_DATAPATH__abc_16259_n3871_1;
  wire AES_CORE_DATAPATH__abc_16259_n3873_1;
  wire AES_CORE_DATAPATH__abc_16259_n3874;
  wire AES_CORE_DATAPATH__abc_16259_n3875;
  wire AES_CORE_DATAPATH__abc_16259_n3876;
  wire AES_CORE_DATAPATH__abc_16259_n3877;
  wire AES_CORE_DATAPATH__abc_16259_n3878_1;
  wire AES_CORE_DATAPATH__abc_16259_n3879_1;
  wire AES_CORE_DATAPATH__abc_16259_n3880;
  wire AES_CORE_DATAPATH__abc_16259_n3881_1;
  wire AES_CORE_DATAPATH__abc_16259_n3882;
  wire AES_CORE_DATAPATH__abc_16259_n3883;
  wire AES_CORE_DATAPATH__abc_16259_n3884;
  wire AES_CORE_DATAPATH__abc_16259_n3886_1;
  wire AES_CORE_DATAPATH__abc_16259_n3887_1;
  wire AES_CORE_DATAPATH__abc_16259_n3888;
  wire AES_CORE_DATAPATH__abc_16259_n3889_1;
  wire AES_CORE_DATAPATH__abc_16259_n3890;
  wire AES_CORE_DATAPATH__abc_16259_n3891;
  wire AES_CORE_DATAPATH__abc_16259_n3892;
  wire AES_CORE_DATAPATH__abc_16259_n3894_1;
  wire AES_CORE_DATAPATH__abc_16259_n3895_1;
  wire AES_CORE_DATAPATH__abc_16259_n3896;
  wire AES_CORE_DATAPATH__abc_16259_n3897_1;
  wire AES_CORE_DATAPATH__abc_16259_n3898;
  wire AES_CORE_DATAPATH__abc_16259_n3899;
  wire AES_CORE_DATAPATH__abc_16259_n3900;
  wire AES_CORE_DATAPATH__abc_16259_n3901;
  wire AES_CORE_DATAPATH__abc_16259_n3902_1;
  wire AES_CORE_DATAPATH__abc_16259_n3903_1;
  wire AES_CORE_DATAPATH__abc_16259_n3904;
  wire AES_CORE_DATAPATH__abc_16259_n3905_1;
  wire AES_CORE_DATAPATH__abc_16259_n3906;
  wire AES_CORE_DATAPATH__abc_16259_n3907;
  wire AES_CORE_DATAPATH__abc_16259_n3908;
  wire AES_CORE_DATAPATH__abc_16259_n3909;
  wire AES_CORE_DATAPATH__abc_16259_n3910_1;
  wire AES_CORE_DATAPATH__abc_16259_n3911_1;
  wire AES_CORE_DATAPATH__abc_16259_n3913_1;
  wire AES_CORE_DATAPATH__abc_16259_n3914;
  wire AES_CORE_DATAPATH__abc_16259_n3915;
  wire AES_CORE_DATAPATH__abc_16259_n3916;
  wire AES_CORE_DATAPATH__abc_16259_n3917;
  wire AES_CORE_DATAPATH__abc_16259_n3918_1;
  wire AES_CORE_DATAPATH__abc_16259_n3919_1;
  wire AES_CORE_DATAPATH__abc_16259_n3920;
  wire AES_CORE_DATAPATH__abc_16259_n3921_1;
  wire AES_CORE_DATAPATH__abc_16259_n3922;
  wire AES_CORE_DATAPATH__abc_16259_n3923;
  wire AES_CORE_DATAPATH__abc_16259_n3924;
  wire AES_CORE_DATAPATH__abc_16259_n3926_1;
  wire AES_CORE_DATAPATH__abc_16259_n3927_1;
  wire AES_CORE_DATAPATH__abc_16259_n3928;
  wire AES_CORE_DATAPATH__abc_16259_n3929_1;
  wire AES_CORE_DATAPATH__abc_16259_n3930;
  wire AES_CORE_DATAPATH__abc_16259_n3931;
  wire AES_CORE_DATAPATH__abc_16259_n3932;
  wire AES_CORE_DATAPATH__abc_16259_n3934_1;
  wire AES_CORE_DATAPATH__abc_16259_n3935_1;
  wire AES_CORE_DATAPATH__abc_16259_n3936;
  wire AES_CORE_DATAPATH__abc_16259_n3937_1;
  wire AES_CORE_DATAPATH__abc_16259_n3938;
  wire AES_CORE_DATAPATH__abc_16259_n3939;
  wire AES_CORE_DATAPATH__abc_16259_n3940;
  wire AES_CORE_DATAPATH__abc_16259_n3941;
  wire AES_CORE_DATAPATH__abc_16259_n3942_1;
  wire AES_CORE_DATAPATH__abc_16259_n3943_1;
  wire AES_CORE_DATAPATH__abc_16259_n3944;
  wire AES_CORE_DATAPATH__abc_16259_n3945_1;
  wire AES_CORE_DATAPATH__abc_16259_n3946;
  wire AES_CORE_DATAPATH__abc_16259_n3947;
  wire AES_CORE_DATAPATH__abc_16259_n3948;
  wire AES_CORE_DATAPATH__abc_16259_n3949;
  wire AES_CORE_DATAPATH__abc_16259_n3950_1;
  wire AES_CORE_DATAPATH__abc_16259_n3951_1;
  wire AES_CORE_DATAPATH__abc_16259_n3953_1;
  wire AES_CORE_DATAPATH__abc_16259_n3954;
  wire AES_CORE_DATAPATH__abc_16259_n3955;
  wire AES_CORE_DATAPATH__abc_16259_n3956;
  wire AES_CORE_DATAPATH__abc_16259_n3957;
  wire AES_CORE_DATAPATH__abc_16259_n3958_1;
  wire AES_CORE_DATAPATH__abc_16259_n3959_1;
  wire AES_CORE_DATAPATH__abc_16259_n3960;
  wire AES_CORE_DATAPATH__abc_16259_n3961_1;
  wire AES_CORE_DATAPATH__abc_16259_n3962;
  wire AES_CORE_DATAPATH__abc_16259_n3963;
  wire AES_CORE_DATAPATH__abc_16259_n3964;
  wire AES_CORE_DATAPATH__abc_16259_n3966_1;
  wire AES_CORE_DATAPATH__abc_16259_n3967_1;
  wire AES_CORE_DATAPATH__abc_16259_n3968;
  wire AES_CORE_DATAPATH__abc_16259_n3969_1;
  wire AES_CORE_DATAPATH__abc_16259_n3970;
  wire AES_CORE_DATAPATH__abc_16259_n3971;
  wire AES_CORE_DATAPATH__abc_16259_n3972;
  wire AES_CORE_DATAPATH__abc_16259_n3974_1;
  wire AES_CORE_DATAPATH__abc_16259_n3975_1;
  wire AES_CORE_DATAPATH__abc_16259_n3976;
  wire AES_CORE_DATAPATH__abc_16259_n3977_1;
  wire AES_CORE_DATAPATH__abc_16259_n3978;
  wire AES_CORE_DATAPATH__abc_16259_n3979;
  wire AES_CORE_DATAPATH__abc_16259_n3980;
  wire AES_CORE_DATAPATH__abc_16259_n3981;
  wire AES_CORE_DATAPATH__abc_16259_n3982_1;
  wire AES_CORE_DATAPATH__abc_16259_n3983_1;
  wire AES_CORE_DATAPATH__abc_16259_n3984;
  wire AES_CORE_DATAPATH__abc_16259_n3985_1;
  wire AES_CORE_DATAPATH__abc_16259_n3986;
  wire AES_CORE_DATAPATH__abc_16259_n3987;
  wire AES_CORE_DATAPATH__abc_16259_n3988;
  wire AES_CORE_DATAPATH__abc_16259_n3989;
  wire AES_CORE_DATAPATH__abc_16259_n3990_1;
  wire AES_CORE_DATAPATH__abc_16259_n3991_1;
  wire AES_CORE_DATAPATH__abc_16259_n3993_1;
  wire AES_CORE_DATAPATH__abc_16259_n3994;
  wire AES_CORE_DATAPATH__abc_16259_n3995;
  wire AES_CORE_DATAPATH__abc_16259_n3996;
  wire AES_CORE_DATAPATH__abc_16259_n3997;
  wire AES_CORE_DATAPATH__abc_16259_n3998_1;
  wire AES_CORE_DATAPATH__abc_16259_n3999_1;
  wire AES_CORE_DATAPATH__abc_16259_n4000;
  wire AES_CORE_DATAPATH__abc_16259_n4001_1;
  wire AES_CORE_DATAPATH__abc_16259_n4002;
  wire AES_CORE_DATAPATH__abc_16259_n4003;
  wire AES_CORE_DATAPATH__abc_16259_n4004;
  wire AES_CORE_DATAPATH__abc_16259_n4006_1;
  wire AES_CORE_DATAPATH__abc_16259_n4007_1;
  wire AES_CORE_DATAPATH__abc_16259_n4008;
  wire AES_CORE_DATAPATH__abc_16259_n4009_1;
  wire AES_CORE_DATAPATH__abc_16259_n4010;
  wire AES_CORE_DATAPATH__abc_16259_n4011;
  wire AES_CORE_DATAPATH__abc_16259_n4012;
  wire AES_CORE_DATAPATH__abc_16259_n4014_1;
  wire AES_CORE_DATAPATH__abc_16259_n4015_1;
  wire AES_CORE_DATAPATH__abc_16259_n4016;
  wire AES_CORE_DATAPATH__abc_16259_n4017_1;
  wire AES_CORE_DATAPATH__abc_16259_n4018;
  wire AES_CORE_DATAPATH__abc_16259_n4019;
  wire AES_CORE_DATAPATH__abc_16259_n4020;
  wire AES_CORE_DATAPATH__abc_16259_n4021;
  wire AES_CORE_DATAPATH__abc_16259_n4022_1;
  wire AES_CORE_DATAPATH__abc_16259_n4023_1;
  wire AES_CORE_DATAPATH__abc_16259_n4024;
  wire AES_CORE_DATAPATH__abc_16259_n4025_1;
  wire AES_CORE_DATAPATH__abc_16259_n4026;
  wire AES_CORE_DATAPATH__abc_16259_n4027;
  wire AES_CORE_DATAPATH__abc_16259_n4028;
  wire AES_CORE_DATAPATH__abc_16259_n4029;
  wire AES_CORE_DATAPATH__abc_16259_n4030_1;
  wire AES_CORE_DATAPATH__abc_16259_n4031_1;
  wire AES_CORE_DATAPATH__abc_16259_n4033_1;
  wire AES_CORE_DATAPATH__abc_16259_n4034;
  wire AES_CORE_DATAPATH__abc_16259_n4035;
  wire AES_CORE_DATAPATH__abc_16259_n4036;
  wire AES_CORE_DATAPATH__abc_16259_n4037;
  wire AES_CORE_DATAPATH__abc_16259_n4038_1;
  wire AES_CORE_DATAPATH__abc_16259_n4039_1;
  wire AES_CORE_DATAPATH__abc_16259_n4040;
  wire AES_CORE_DATAPATH__abc_16259_n4041_1;
  wire AES_CORE_DATAPATH__abc_16259_n4042;
  wire AES_CORE_DATAPATH__abc_16259_n4043;
  wire AES_CORE_DATAPATH__abc_16259_n4044;
  wire AES_CORE_DATAPATH__abc_16259_n4046_1;
  wire AES_CORE_DATAPATH__abc_16259_n4047_1;
  wire AES_CORE_DATAPATH__abc_16259_n4048;
  wire AES_CORE_DATAPATH__abc_16259_n4049_1;
  wire AES_CORE_DATAPATH__abc_16259_n4050;
  wire AES_CORE_DATAPATH__abc_16259_n4051;
  wire AES_CORE_DATAPATH__abc_16259_n4052;
  wire AES_CORE_DATAPATH__abc_16259_n4054_1;
  wire AES_CORE_DATAPATH__abc_16259_n4055_1;
  wire AES_CORE_DATAPATH__abc_16259_n4056;
  wire AES_CORE_DATAPATH__abc_16259_n4057_1;
  wire AES_CORE_DATAPATH__abc_16259_n4058;
  wire AES_CORE_DATAPATH__abc_16259_n4059;
  wire AES_CORE_DATAPATH__abc_16259_n4060;
  wire AES_CORE_DATAPATH__abc_16259_n4061;
  wire AES_CORE_DATAPATH__abc_16259_n4062_1;
  wire AES_CORE_DATAPATH__abc_16259_n4063_1;
  wire AES_CORE_DATAPATH__abc_16259_n4064;
  wire AES_CORE_DATAPATH__abc_16259_n4065_1;
  wire AES_CORE_DATAPATH__abc_16259_n4066;
  wire AES_CORE_DATAPATH__abc_16259_n4067;
  wire AES_CORE_DATAPATH__abc_16259_n4068;
  wire AES_CORE_DATAPATH__abc_16259_n4069;
  wire AES_CORE_DATAPATH__abc_16259_n4070_1;
  wire AES_CORE_DATAPATH__abc_16259_n4071_1;
  wire AES_CORE_DATAPATH__abc_16259_n4073_1;
  wire AES_CORE_DATAPATH__abc_16259_n4074;
  wire AES_CORE_DATAPATH__abc_16259_n4075;
  wire AES_CORE_DATAPATH__abc_16259_n4076;
  wire AES_CORE_DATAPATH__abc_16259_n4077;
  wire AES_CORE_DATAPATH__abc_16259_n4078_1;
  wire AES_CORE_DATAPATH__abc_16259_n4079_1;
  wire AES_CORE_DATAPATH__abc_16259_n4080;
  wire AES_CORE_DATAPATH__abc_16259_n4081_1;
  wire AES_CORE_DATAPATH__abc_16259_n4082;
  wire AES_CORE_DATAPATH__abc_16259_n4083;
  wire AES_CORE_DATAPATH__abc_16259_n4084;
  wire AES_CORE_DATAPATH__abc_16259_n4086_1;
  wire AES_CORE_DATAPATH__abc_16259_n4087_1;
  wire AES_CORE_DATAPATH__abc_16259_n4088;
  wire AES_CORE_DATAPATH__abc_16259_n4089_1;
  wire AES_CORE_DATAPATH__abc_16259_n4090;
  wire AES_CORE_DATAPATH__abc_16259_n4091;
  wire AES_CORE_DATAPATH__abc_16259_n4092;
  wire AES_CORE_DATAPATH__abc_16259_n4094_1;
  wire AES_CORE_DATAPATH__abc_16259_n4095_1;
  wire AES_CORE_DATAPATH__abc_16259_n4096;
  wire AES_CORE_DATAPATH__abc_16259_n4097_1;
  wire AES_CORE_DATAPATH__abc_16259_n4098;
  wire AES_CORE_DATAPATH__abc_16259_n4099;
  wire AES_CORE_DATAPATH__abc_16259_n4100;
  wire AES_CORE_DATAPATH__abc_16259_n4101;
  wire AES_CORE_DATAPATH__abc_16259_n4102_1;
  wire AES_CORE_DATAPATH__abc_16259_n4103_1;
  wire AES_CORE_DATAPATH__abc_16259_n4104;
  wire AES_CORE_DATAPATH__abc_16259_n4105_1;
  wire AES_CORE_DATAPATH__abc_16259_n4106;
  wire AES_CORE_DATAPATH__abc_16259_n4107;
  wire AES_CORE_DATAPATH__abc_16259_n4108;
  wire AES_CORE_DATAPATH__abc_16259_n4109;
  wire AES_CORE_DATAPATH__abc_16259_n4110_1;
  wire AES_CORE_DATAPATH__abc_16259_n4111_1;
  wire AES_CORE_DATAPATH__abc_16259_n4113_1;
  wire AES_CORE_DATAPATH__abc_16259_n4114;
  wire AES_CORE_DATAPATH__abc_16259_n4116;
  wire AES_CORE_DATAPATH__abc_16259_n4117;
  wire AES_CORE_DATAPATH__abc_16259_n4119_1;
  wire AES_CORE_DATAPATH__abc_16259_n4120;
  wire AES_CORE_DATAPATH__abc_16259_n4122;
  wire AES_CORE_DATAPATH__abc_16259_n4123;
  wire AES_CORE_DATAPATH__abc_16259_n4125;
  wire AES_CORE_DATAPATH__abc_16259_n4126_1;
  wire AES_CORE_DATAPATH__abc_16259_n4128;
  wire AES_CORE_DATAPATH__abc_16259_n4129_1;
  wire AES_CORE_DATAPATH__abc_16259_n4131;
  wire AES_CORE_DATAPATH__abc_16259_n4132;
  wire AES_CORE_DATAPATH__abc_16259_n4134_1;
  wire AES_CORE_DATAPATH__abc_16259_n4135_1;
  wire AES_CORE_DATAPATH__abc_16259_n4137_1;
  wire AES_CORE_DATAPATH__abc_16259_n4138;
  wire AES_CORE_DATAPATH__abc_16259_n4140;
  wire AES_CORE_DATAPATH__abc_16259_n4141;
  wire AES_CORE_DATAPATH__abc_16259_n4143_1;
  wire AES_CORE_DATAPATH__abc_16259_n4144;
  wire AES_CORE_DATAPATH__abc_16259_n4146;
  wire AES_CORE_DATAPATH__abc_16259_n4147;
  wire AES_CORE_DATAPATH__abc_16259_n4149;
  wire AES_CORE_DATAPATH__abc_16259_n4150_1;
  wire AES_CORE_DATAPATH__abc_16259_n4152;
  wire AES_CORE_DATAPATH__abc_16259_n4153_1;
  wire AES_CORE_DATAPATH__abc_16259_n4155;
  wire AES_CORE_DATAPATH__abc_16259_n4156;
  wire AES_CORE_DATAPATH__abc_16259_n4158_1;
  wire AES_CORE_DATAPATH__abc_16259_n4159_1;
  wire AES_CORE_DATAPATH__abc_16259_n4161_1;
  wire AES_CORE_DATAPATH__abc_16259_n4162;
  wire AES_CORE_DATAPATH__abc_16259_n4164;
  wire AES_CORE_DATAPATH__abc_16259_n4165;
  wire AES_CORE_DATAPATH__abc_16259_n4167_1;
  wire AES_CORE_DATAPATH__abc_16259_n4168;
  wire AES_CORE_DATAPATH__abc_16259_n4170;
  wire AES_CORE_DATAPATH__abc_16259_n4171;
  wire AES_CORE_DATAPATH__abc_16259_n4173;
  wire AES_CORE_DATAPATH__abc_16259_n4174_1;
  wire AES_CORE_DATAPATH__abc_16259_n4176;
  wire AES_CORE_DATAPATH__abc_16259_n4177_1;
  wire AES_CORE_DATAPATH__abc_16259_n4179;
  wire AES_CORE_DATAPATH__abc_16259_n4180;
  wire AES_CORE_DATAPATH__abc_16259_n4182_1;
  wire AES_CORE_DATAPATH__abc_16259_n4183_1;
  wire AES_CORE_DATAPATH__abc_16259_n4185_1;
  wire AES_CORE_DATAPATH__abc_16259_n4186;
  wire AES_CORE_DATAPATH__abc_16259_n4188;
  wire AES_CORE_DATAPATH__abc_16259_n4189;
  wire AES_CORE_DATAPATH__abc_16259_n4191_1;
  wire AES_CORE_DATAPATH__abc_16259_n4192;
  wire AES_CORE_DATAPATH__abc_16259_n4194;
  wire AES_CORE_DATAPATH__abc_16259_n4195;
  wire AES_CORE_DATAPATH__abc_16259_n4197;
  wire AES_CORE_DATAPATH__abc_16259_n4198_1;
  wire AES_CORE_DATAPATH__abc_16259_n4200;
  wire AES_CORE_DATAPATH__abc_16259_n4201_1;
  wire AES_CORE_DATAPATH__abc_16259_n4203;
  wire AES_CORE_DATAPATH__abc_16259_n4204;
  wire AES_CORE_DATAPATH__abc_16259_n4206_1;
  wire AES_CORE_DATAPATH__abc_16259_n4207_1;
  wire AES_CORE_DATAPATH__abc_16259_n4209_1;
  wire AES_CORE_DATAPATH__abc_16259_n4210;
  wire AES_CORE_DATAPATH__abc_16259_n4211;
  wire AES_CORE_DATAPATH__abc_16259_n4212;
  wire AES_CORE_DATAPATH__abc_16259_n4213;
  wire AES_CORE_DATAPATH__abc_16259_n4214_1;
  wire AES_CORE_DATAPATH__abc_16259_n4215_1;
  wire AES_CORE_DATAPATH__abc_16259_n4217_1;
  wire AES_CORE_DATAPATH__abc_16259_n4218;
  wire AES_CORE_DATAPATH__abc_16259_n4219;
  wire AES_CORE_DATAPATH__abc_16259_n4220;
  wire AES_CORE_DATAPATH__abc_16259_n4221;
  wire AES_CORE_DATAPATH__abc_16259_n4222_1;
  wire AES_CORE_DATAPATH__abc_16259_n4223_1;
  wire AES_CORE_DATAPATH__abc_16259_n4225_1;
  wire AES_CORE_DATAPATH__abc_16259_n4226;
  wire AES_CORE_DATAPATH__abc_16259_n4227;
  wire AES_CORE_DATAPATH__abc_16259_n4228;
  wire AES_CORE_DATAPATH__abc_16259_n4229;
  wire AES_CORE_DATAPATH__abc_16259_n4230_1;
  wire AES_CORE_DATAPATH__abc_16259_n4231_1;
  wire AES_CORE_DATAPATH__abc_16259_n4233_1;
  wire AES_CORE_DATAPATH__abc_16259_n4234;
  wire AES_CORE_DATAPATH__abc_16259_n4235;
  wire AES_CORE_DATAPATH__abc_16259_n4236;
  wire AES_CORE_DATAPATH__abc_16259_n4237;
  wire AES_CORE_DATAPATH__abc_16259_n4238_1;
  wire AES_CORE_DATAPATH__abc_16259_n4239_1;
  wire AES_CORE_DATAPATH__abc_16259_n4241_1;
  wire AES_CORE_DATAPATH__abc_16259_n4242;
  wire AES_CORE_DATAPATH__abc_16259_n4243;
  wire AES_CORE_DATAPATH__abc_16259_n4244;
  wire AES_CORE_DATAPATH__abc_16259_n4245;
  wire AES_CORE_DATAPATH__abc_16259_n4246_1;
  wire AES_CORE_DATAPATH__abc_16259_n4247_1;
  wire AES_CORE_DATAPATH__abc_16259_n4249_1;
  wire AES_CORE_DATAPATH__abc_16259_n4250;
  wire AES_CORE_DATAPATH__abc_16259_n4251;
  wire AES_CORE_DATAPATH__abc_16259_n4252;
  wire AES_CORE_DATAPATH__abc_16259_n4253;
  wire AES_CORE_DATAPATH__abc_16259_n4254_1;
  wire AES_CORE_DATAPATH__abc_16259_n4255_1;
  wire AES_CORE_DATAPATH__abc_16259_n4257_1;
  wire AES_CORE_DATAPATH__abc_16259_n4258;
  wire AES_CORE_DATAPATH__abc_16259_n4259;
  wire AES_CORE_DATAPATH__abc_16259_n4260;
  wire AES_CORE_DATAPATH__abc_16259_n4261;
  wire AES_CORE_DATAPATH__abc_16259_n4262_1;
  wire AES_CORE_DATAPATH__abc_16259_n4263_1;
  wire AES_CORE_DATAPATH__abc_16259_n4265_1;
  wire AES_CORE_DATAPATH__abc_16259_n4266;
  wire AES_CORE_DATAPATH__abc_16259_n4267;
  wire AES_CORE_DATAPATH__abc_16259_n4268;
  wire AES_CORE_DATAPATH__abc_16259_n4269;
  wire AES_CORE_DATAPATH__abc_16259_n4270_1;
  wire AES_CORE_DATAPATH__abc_16259_n4271_1;
  wire AES_CORE_DATAPATH__abc_16259_n4273_1;
  wire AES_CORE_DATAPATH__abc_16259_n4274;
  wire AES_CORE_DATAPATH__abc_16259_n4275;
  wire AES_CORE_DATAPATH__abc_16259_n4276;
  wire AES_CORE_DATAPATH__abc_16259_n4277;
  wire AES_CORE_DATAPATH__abc_16259_n4278_1;
  wire AES_CORE_DATAPATH__abc_16259_n4279_1;
  wire AES_CORE_DATAPATH__abc_16259_n4281_1;
  wire AES_CORE_DATAPATH__abc_16259_n4282;
  wire AES_CORE_DATAPATH__abc_16259_n4283;
  wire AES_CORE_DATAPATH__abc_16259_n4284;
  wire AES_CORE_DATAPATH__abc_16259_n4285;
  wire AES_CORE_DATAPATH__abc_16259_n4286_1;
  wire AES_CORE_DATAPATH__abc_16259_n4287_1;
  wire AES_CORE_DATAPATH__abc_16259_n4289_1;
  wire AES_CORE_DATAPATH__abc_16259_n4290;
  wire AES_CORE_DATAPATH__abc_16259_n4291;
  wire AES_CORE_DATAPATH__abc_16259_n4292;
  wire AES_CORE_DATAPATH__abc_16259_n4293;
  wire AES_CORE_DATAPATH__abc_16259_n4294_1;
  wire AES_CORE_DATAPATH__abc_16259_n4295_1;
  wire AES_CORE_DATAPATH__abc_16259_n4297_1;
  wire AES_CORE_DATAPATH__abc_16259_n4298;
  wire AES_CORE_DATAPATH__abc_16259_n4299;
  wire AES_CORE_DATAPATH__abc_16259_n4300;
  wire AES_CORE_DATAPATH__abc_16259_n4301;
  wire AES_CORE_DATAPATH__abc_16259_n4302_1;
  wire AES_CORE_DATAPATH__abc_16259_n4303_1;
  wire AES_CORE_DATAPATH__abc_16259_n4305_1;
  wire AES_CORE_DATAPATH__abc_16259_n4306;
  wire AES_CORE_DATAPATH__abc_16259_n4307;
  wire AES_CORE_DATAPATH__abc_16259_n4308;
  wire AES_CORE_DATAPATH__abc_16259_n4309;
  wire AES_CORE_DATAPATH__abc_16259_n4310_1;
  wire AES_CORE_DATAPATH__abc_16259_n4311_1;
  wire AES_CORE_DATAPATH__abc_16259_n4313_1;
  wire AES_CORE_DATAPATH__abc_16259_n4314;
  wire AES_CORE_DATAPATH__abc_16259_n4315;
  wire AES_CORE_DATAPATH__abc_16259_n4316;
  wire AES_CORE_DATAPATH__abc_16259_n4317;
  wire AES_CORE_DATAPATH__abc_16259_n4318_1;
  wire AES_CORE_DATAPATH__abc_16259_n4319_1;
  wire AES_CORE_DATAPATH__abc_16259_n4321_1;
  wire AES_CORE_DATAPATH__abc_16259_n4322;
  wire AES_CORE_DATAPATH__abc_16259_n4323;
  wire AES_CORE_DATAPATH__abc_16259_n4324;
  wire AES_CORE_DATAPATH__abc_16259_n4325;
  wire AES_CORE_DATAPATH__abc_16259_n4326_1;
  wire AES_CORE_DATAPATH__abc_16259_n4327_1;
  wire AES_CORE_DATAPATH__abc_16259_n4329_1;
  wire AES_CORE_DATAPATH__abc_16259_n4330;
  wire AES_CORE_DATAPATH__abc_16259_n4331;
  wire AES_CORE_DATAPATH__abc_16259_n4332;
  wire AES_CORE_DATAPATH__abc_16259_n4333;
  wire AES_CORE_DATAPATH__abc_16259_n4334_1;
  wire AES_CORE_DATAPATH__abc_16259_n4335_1;
  wire AES_CORE_DATAPATH__abc_16259_n4337_1;
  wire AES_CORE_DATAPATH__abc_16259_n4338;
  wire AES_CORE_DATAPATH__abc_16259_n4339;
  wire AES_CORE_DATAPATH__abc_16259_n4340;
  wire AES_CORE_DATAPATH__abc_16259_n4341;
  wire AES_CORE_DATAPATH__abc_16259_n4342_1;
  wire AES_CORE_DATAPATH__abc_16259_n4343_1;
  wire AES_CORE_DATAPATH__abc_16259_n4345_1;
  wire AES_CORE_DATAPATH__abc_16259_n4346;
  wire AES_CORE_DATAPATH__abc_16259_n4347;
  wire AES_CORE_DATAPATH__abc_16259_n4348;
  wire AES_CORE_DATAPATH__abc_16259_n4349;
  wire AES_CORE_DATAPATH__abc_16259_n4350_1;
  wire AES_CORE_DATAPATH__abc_16259_n4351_1;
  wire AES_CORE_DATAPATH__abc_16259_n4353_1;
  wire AES_CORE_DATAPATH__abc_16259_n4354;
  wire AES_CORE_DATAPATH__abc_16259_n4355;
  wire AES_CORE_DATAPATH__abc_16259_n4356;
  wire AES_CORE_DATAPATH__abc_16259_n4357;
  wire AES_CORE_DATAPATH__abc_16259_n4358_1;
  wire AES_CORE_DATAPATH__abc_16259_n4359_1;
  wire AES_CORE_DATAPATH__abc_16259_n4361_1;
  wire AES_CORE_DATAPATH__abc_16259_n4362;
  wire AES_CORE_DATAPATH__abc_16259_n4363;
  wire AES_CORE_DATAPATH__abc_16259_n4364;
  wire AES_CORE_DATAPATH__abc_16259_n4365;
  wire AES_CORE_DATAPATH__abc_16259_n4366_1;
  wire AES_CORE_DATAPATH__abc_16259_n4367_1;
  wire AES_CORE_DATAPATH__abc_16259_n4369_1;
  wire AES_CORE_DATAPATH__abc_16259_n4370;
  wire AES_CORE_DATAPATH__abc_16259_n4371;
  wire AES_CORE_DATAPATH__abc_16259_n4372;
  wire AES_CORE_DATAPATH__abc_16259_n4373;
  wire AES_CORE_DATAPATH__abc_16259_n4374_1;
  wire AES_CORE_DATAPATH__abc_16259_n4375_1;
  wire AES_CORE_DATAPATH__abc_16259_n4377_1;
  wire AES_CORE_DATAPATH__abc_16259_n4378;
  wire AES_CORE_DATAPATH__abc_16259_n4379;
  wire AES_CORE_DATAPATH__abc_16259_n4380;
  wire AES_CORE_DATAPATH__abc_16259_n4381;
  wire AES_CORE_DATAPATH__abc_16259_n4382_1;
  wire AES_CORE_DATAPATH__abc_16259_n4383_1;
  wire AES_CORE_DATAPATH__abc_16259_n4385_1;
  wire AES_CORE_DATAPATH__abc_16259_n4386;
  wire AES_CORE_DATAPATH__abc_16259_n4387;
  wire AES_CORE_DATAPATH__abc_16259_n4388;
  wire AES_CORE_DATAPATH__abc_16259_n4389;
  wire AES_CORE_DATAPATH__abc_16259_n4390_1;
  wire AES_CORE_DATAPATH__abc_16259_n4391_1;
  wire AES_CORE_DATAPATH__abc_16259_n4393_1;
  wire AES_CORE_DATAPATH__abc_16259_n4394;
  wire AES_CORE_DATAPATH__abc_16259_n4395;
  wire AES_CORE_DATAPATH__abc_16259_n4396;
  wire AES_CORE_DATAPATH__abc_16259_n4397;
  wire AES_CORE_DATAPATH__abc_16259_n4398_1;
  wire AES_CORE_DATAPATH__abc_16259_n4399_1;
  wire AES_CORE_DATAPATH__abc_16259_n4401_1;
  wire AES_CORE_DATAPATH__abc_16259_n4402;
  wire AES_CORE_DATAPATH__abc_16259_n4403;
  wire AES_CORE_DATAPATH__abc_16259_n4404;
  wire AES_CORE_DATAPATH__abc_16259_n4405;
  wire AES_CORE_DATAPATH__abc_16259_n4406_1;
  wire AES_CORE_DATAPATH__abc_16259_n4407_1;
  wire AES_CORE_DATAPATH__abc_16259_n4409_1;
  wire AES_CORE_DATAPATH__abc_16259_n4410;
  wire AES_CORE_DATAPATH__abc_16259_n4411;
  wire AES_CORE_DATAPATH__abc_16259_n4412;
  wire AES_CORE_DATAPATH__abc_16259_n4413;
  wire AES_CORE_DATAPATH__abc_16259_n4414_1;
  wire AES_CORE_DATAPATH__abc_16259_n4415_1;
  wire AES_CORE_DATAPATH__abc_16259_n4417_1;
  wire AES_CORE_DATAPATH__abc_16259_n4418;
  wire AES_CORE_DATAPATH__abc_16259_n4419;
  wire AES_CORE_DATAPATH__abc_16259_n4420;
  wire AES_CORE_DATAPATH__abc_16259_n4421;
  wire AES_CORE_DATAPATH__abc_16259_n4422_1;
  wire AES_CORE_DATAPATH__abc_16259_n4423_1;
  wire AES_CORE_DATAPATH__abc_16259_n4425_1;
  wire AES_CORE_DATAPATH__abc_16259_n4426;
  wire AES_CORE_DATAPATH__abc_16259_n4427;
  wire AES_CORE_DATAPATH__abc_16259_n4428;
  wire AES_CORE_DATAPATH__abc_16259_n4429;
  wire AES_CORE_DATAPATH__abc_16259_n4430_1;
  wire AES_CORE_DATAPATH__abc_16259_n4431_1;
  wire AES_CORE_DATAPATH__abc_16259_n4433_1;
  wire AES_CORE_DATAPATH__abc_16259_n4434;
  wire AES_CORE_DATAPATH__abc_16259_n4435;
  wire AES_CORE_DATAPATH__abc_16259_n4436;
  wire AES_CORE_DATAPATH__abc_16259_n4437;
  wire AES_CORE_DATAPATH__abc_16259_n4438_1;
  wire AES_CORE_DATAPATH__abc_16259_n4439;
  wire AES_CORE_DATAPATH__abc_16259_n4441;
  wire AES_CORE_DATAPATH__abc_16259_n4442;
  wire AES_CORE_DATAPATH__abc_16259_n4443_1;
  wire AES_CORE_DATAPATH__abc_16259_n4444_1;
  wire AES_CORE_DATAPATH__abc_16259_n4445_1;
  wire AES_CORE_DATAPATH__abc_16259_n4446_1;
  wire AES_CORE_DATAPATH__abc_16259_n4447_1;
  wire AES_CORE_DATAPATH__abc_16259_n4449_1;
  wire AES_CORE_DATAPATH__abc_16259_n4450_1;
  wire AES_CORE_DATAPATH__abc_16259_n4451_1;
  wire AES_CORE_DATAPATH__abc_16259_n4452_1;
  wire AES_CORE_DATAPATH__abc_16259_n4453_1;
  wire AES_CORE_DATAPATH__abc_16259_n4454_1;
  wire AES_CORE_DATAPATH__abc_16259_n4455_1;
  wire AES_CORE_DATAPATH__abc_16259_n4457_1;
  wire AES_CORE_DATAPATH__abc_16259_n4458_1;
  wire AES_CORE_DATAPATH__abc_16259_n4459_1;
  wire AES_CORE_DATAPATH__abc_16259_n4460_1;
  wire AES_CORE_DATAPATH__abc_16259_n4461_1;
  wire AES_CORE_DATAPATH__abc_16259_n4462_1;
  wire AES_CORE_DATAPATH__abc_16259_n4463_1;
  wire AES_CORE_DATAPATH__abc_16259_n4466_1;
  wire AES_CORE_DATAPATH__abc_16259_n4467_1;
  wire AES_CORE_DATAPATH__abc_16259_n4468_1;
  wire AES_CORE_DATAPATH__abc_16259_n4468_1_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n4468_1_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n4468_1_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n4468_1_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n4468_1_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n4469_1;
  wire AES_CORE_DATAPATH__abc_16259_n4470_1;
  wire AES_CORE_DATAPATH__abc_16259_n4471_1;
  wire AES_CORE_DATAPATH__abc_16259_n4472_1;
  wire AES_CORE_DATAPATH__abc_16259_n4473_1;
  wire AES_CORE_DATAPATH__abc_16259_n4474_1;
  wire AES_CORE_DATAPATH__abc_16259_n4474_1_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n4474_1_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n4474_1_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n4474_1_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n4474_1_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n4475_1;
  wire AES_CORE_DATAPATH__abc_16259_n4475_1_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n4475_1_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n4475_1_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n4475_1_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n4475_1_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n4476_1;
  wire AES_CORE_DATAPATH__abc_16259_n4477_1;
  wire AES_CORE_DATAPATH__abc_16259_n4478_1;
  wire AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf10;
  wire AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf5;
  wire AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf6;
  wire AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf7;
  wire AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf8;
  wire AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf9;
  wire AES_CORE_DATAPATH__abc_16259_n4479_1;
  wire AES_CORE_DATAPATH__abc_16259_n4480_1;
  wire AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf10;
  wire AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf5;
  wire AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf6;
  wire AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf7;
  wire AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf8;
  wire AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf9;
  wire AES_CORE_DATAPATH__abc_16259_n4481_1;
  wire AES_CORE_DATAPATH__abc_16259_n4482_1;
  wire AES_CORE_DATAPATH__abc_16259_n4483_1;
  wire AES_CORE_DATAPATH__abc_16259_n4484_1;
  wire AES_CORE_DATAPATH__abc_16259_n4485_1;
  wire AES_CORE_DATAPATH__abc_16259_n4486_1;
  wire AES_CORE_DATAPATH__abc_16259_n4487_1;
  wire AES_CORE_DATAPATH__abc_16259_n4489_1;
  wire AES_CORE_DATAPATH__abc_16259_n4490_1;
  wire AES_CORE_DATAPATH__abc_16259_n4491_1;
  wire AES_CORE_DATAPATH__abc_16259_n4492_1;
  wire AES_CORE_DATAPATH__abc_16259_n4493_1;
  wire AES_CORE_DATAPATH__abc_16259_n4494_1;
  wire AES_CORE_DATAPATH__abc_16259_n4495_1;
  wire AES_CORE_DATAPATH__abc_16259_n4496_1;
  wire AES_CORE_DATAPATH__abc_16259_n4498_1;
  wire AES_CORE_DATAPATH__abc_16259_n4499_1;
  wire AES_CORE_DATAPATH__abc_16259_n4500_1;
  wire AES_CORE_DATAPATH__abc_16259_n4501_1;
  wire AES_CORE_DATAPATH__abc_16259_n4502_1;
  wire AES_CORE_DATAPATH__abc_16259_n4503_1;
  wire AES_CORE_DATAPATH__abc_16259_n4504_1;
  wire AES_CORE_DATAPATH__abc_16259_n4505_1;
  wire AES_CORE_DATAPATH__abc_16259_n4507;
  wire AES_CORE_DATAPATH__abc_16259_n4508;
  wire AES_CORE_DATAPATH__abc_16259_n4509;
  wire AES_CORE_DATAPATH__abc_16259_n4510_1;
  wire AES_CORE_DATAPATH__abc_16259_n4511;
  wire AES_CORE_DATAPATH__abc_16259_n4512;
  wire AES_CORE_DATAPATH__abc_16259_n4513_1;
  wire AES_CORE_DATAPATH__abc_16259_n4514;
  wire AES_CORE_DATAPATH__abc_16259_n4516_1;
  wire AES_CORE_DATAPATH__abc_16259_n4517;
  wire AES_CORE_DATAPATH__abc_16259_n4518;
  wire AES_CORE_DATAPATH__abc_16259_n4519_1;
  wire AES_CORE_DATAPATH__abc_16259_n4520;
  wire AES_CORE_DATAPATH__abc_16259_n4521;
  wire AES_CORE_DATAPATH__abc_16259_n4522_1;
  wire AES_CORE_DATAPATH__abc_16259_n4523;
  wire AES_CORE_DATAPATH__abc_16259_n4525_1;
  wire AES_CORE_DATAPATH__abc_16259_n4526;
  wire AES_CORE_DATAPATH__abc_16259_n4527;
  wire AES_CORE_DATAPATH__abc_16259_n4528_1;
  wire AES_CORE_DATAPATH__abc_16259_n4529;
  wire AES_CORE_DATAPATH__abc_16259_n4530;
  wire AES_CORE_DATAPATH__abc_16259_n4531_1;
  wire AES_CORE_DATAPATH__abc_16259_n4532;
  wire AES_CORE_DATAPATH__abc_16259_n4534_1;
  wire AES_CORE_DATAPATH__abc_16259_n4535;
  wire AES_CORE_DATAPATH__abc_16259_n4536;
  wire AES_CORE_DATAPATH__abc_16259_n4537_1;
  wire AES_CORE_DATAPATH__abc_16259_n4538;
  wire AES_CORE_DATAPATH__abc_16259_n4539;
  wire AES_CORE_DATAPATH__abc_16259_n4540_1;
  wire AES_CORE_DATAPATH__abc_16259_n4541;
  wire AES_CORE_DATAPATH__abc_16259_n4543_1;
  wire AES_CORE_DATAPATH__abc_16259_n4544;
  wire AES_CORE_DATAPATH__abc_16259_n4545;
  wire AES_CORE_DATAPATH__abc_16259_n4546_1;
  wire AES_CORE_DATAPATH__abc_16259_n4547;
  wire AES_CORE_DATAPATH__abc_16259_n4548;
  wire AES_CORE_DATAPATH__abc_16259_n4549_1;
  wire AES_CORE_DATAPATH__abc_16259_n4550;
  wire AES_CORE_DATAPATH__abc_16259_n4552_1;
  wire AES_CORE_DATAPATH__abc_16259_n4553;
  wire AES_CORE_DATAPATH__abc_16259_n4554;
  wire AES_CORE_DATAPATH__abc_16259_n4555_1;
  wire AES_CORE_DATAPATH__abc_16259_n4556;
  wire AES_CORE_DATAPATH__abc_16259_n4557;
  wire AES_CORE_DATAPATH__abc_16259_n4558_1;
  wire AES_CORE_DATAPATH__abc_16259_n4559;
  wire AES_CORE_DATAPATH__abc_16259_n4561_1;
  wire AES_CORE_DATAPATH__abc_16259_n4562;
  wire AES_CORE_DATAPATH__abc_16259_n4563;
  wire AES_CORE_DATAPATH__abc_16259_n4564_1;
  wire AES_CORE_DATAPATH__abc_16259_n4565;
  wire AES_CORE_DATAPATH__abc_16259_n4566;
  wire AES_CORE_DATAPATH__abc_16259_n4567_1;
  wire AES_CORE_DATAPATH__abc_16259_n4568;
  wire AES_CORE_DATAPATH__abc_16259_n4570_1;
  wire AES_CORE_DATAPATH__abc_16259_n4571;
  wire AES_CORE_DATAPATH__abc_16259_n4572;
  wire AES_CORE_DATAPATH__abc_16259_n4573_1;
  wire AES_CORE_DATAPATH__abc_16259_n4574;
  wire AES_CORE_DATAPATH__abc_16259_n4575;
  wire AES_CORE_DATAPATH__abc_16259_n4576_1;
  wire AES_CORE_DATAPATH__abc_16259_n4577;
  wire AES_CORE_DATAPATH__abc_16259_n4579_1;
  wire AES_CORE_DATAPATH__abc_16259_n4580;
  wire AES_CORE_DATAPATH__abc_16259_n4581;
  wire AES_CORE_DATAPATH__abc_16259_n4582_1;
  wire AES_CORE_DATAPATH__abc_16259_n4583;
  wire AES_CORE_DATAPATH__abc_16259_n4584;
  wire AES_CORE_DATAPATH__abc_16259_n4585_1;
  wire AES_CORE_DATAPATH__abc_16259_n4586;
  wire AES_CORE_DATAPATH__abc_16259_n4588_1;
  wire AES_CORE_DATAPATH__abc_16259_n4589;
  wire AES_CORE_DATAPATH__abc_16259_n4590;
  wire AES_CORE_DATAPATH__abc_16259_n4591_1;
  wire AES_CORE_DATAPATH__abc_16259_n4592;
  wire AES_CORE_DATAPATH__abc_16259_n4593;
  wire AES_CORE_DATAPATH__abc_16259_n4594_1;
  wire AES_CORE_DATAPATH__abc_16259_n4595;
  wire AES_CORE_DATAPATH__abc_16259_n4597_1;
  wire AES_CORE_DATAPATH__abc_16259_n4598;
  wire AES_CORE_DATAPATH__abc_16259_n4599;
  wire AES_CORE_DATAPATH__abc_16259_n4600_1;
  wire AES_CORE_DATAPATH__abc_16259_n4601;
  wire AES_CORE_DATAPATH__abc_16259_n4602;
  wire AES_CORE_DATAPATH__abc_16259_n4603_1;
  wire AES_CORE_DATAPATH__abc_16259_n4604_1;
  wire AES_CORE_DATAPATH__abc_16259_n4606;
  wire AES_CORE_DATAPATH__abc_16259_n4607_1;
  wire AES_CORE_DATAPATH__abc_16259_n4608;
  wire AES_CORE_DATAPATH__abc_16259_n4609;
  wire AES_CORE_DATAPATH__abc_16259_n4610;
  wire AES_CORE_DATAPATH__abc_16259_n4611_1;
  wire AES_CORE_DATAPATH__abc_16259_n4612;
  wire AES_CORE_DATAPATH__abc_16259_n4613;
  wire AES_CORE_DATAPATH__abc_16259_n4615;
  wire AES_CORE_DATAPATH__abc_16259_n4616_1;
  wire AES_CORE_DATAPATH__abc_16259_n4617;
  wire AES_CORE_DATAPATH__abc_16259_n4618;
  wire AES_CORE_DATAPATH__abc_16259_n4619;
  wire AES_CORE_DATAPATH__abc_16259_n4620;
  wire AES_CORE_DATAPATH__abc_16259_n4621;
  wire AES_CORE_DATAPATH__abc_16259_n4622_1;
  wire AES_CORE_DATAPATH__abc_16259_n4624;
  wire AES_CORE_DATAPATH__abc_16259_n4625;
  wire AES_CORE_DATAPATH__abc_16259_n4626;
  wire AES_CORE_DATAPATH__abc_16259_n4627;
  wire AES_CORE_DATAPATH__abc_16259_n4628_1;
  wire AES_CORE_DATAPATH__abc_16259_n4629;
  wire AES_CORE_DATAPATH__abc_16259_n4630;
  wire AES_CORE_DATAPATH__abc_16259_n4631;
  wire AES_CORE_DATAPATH__abc_16259_n4633;
  wire AES_CORE_DATAPATH__abc_16259_n4634;
  wire AES_CORE_DATAPATH__abc_16259_n4635_1;
  wire AES_CORE_DATAPATH__abc_16259_n4636;
  wire AES_CORE_DATAPATH__abc_16259_n4637;
  wire AES_CORE_DATAPATH__abc_16259_n4638;
  wire AES_CORE_DATAPATH__abc_16259_n4639;
  wire AES_CORE_DATAPATH__abc_16259_n4640;
  wire AES_CORE_DATAPATH__abc_16259_n4642;
  wire AES_CORE_DATAPATH__abc_16259_n4643;
  wire AES_CORE_DATAPATH__abc_16259_n4644;
  wire AES_CORE_DATAPATH__abc_16259_n4645;
  wire AES_CORE_DATAPATH__abc_16259_n4646;
  wire AES_CORE_DATAPATH__abc_16259_n4647;
  wire AES_CORE_DATAPATH__abc_16259_n4648_1;
  wire AES_CORE_DATAPATH__abc_16259_n4649;
  wire AES_CORE_DATAPATH__abc_16259_n4651;
  wire AES_CORE_DATAPATH__abc_16259_n4652;
  wire AES_CORE_DATAPATH__abc_16259_n4653;
  wire AES_CORE_DATAPATH__abc_16259_n4654_1;
  wire AES_CORE_DATAPATH__abc_16259_n4655;
  wire AES_CORE_DATAPATH__abc_16259_n4656;
  wire AES_CORE_DATAPATH__abc_16259_n4657;
  wire AES_CORE_DATAPATH__abc_16259_n4658;
  wire AES_CORE_DATAPATH__abc_16259_n4660;
  wire AES_CORE_DATAPATH__abc_16259_n4661;
  wire AES_CORE_DATAPATH__abc_16259_n4662_1;
  wire AES_CORE_DATAPATH__abc_16259_n4663;
  wire AES_CORE_DATAPATH__abc_16259_n4664;
  wire AES_CORE_DATAPATH__abc_16259_n4665;
  wire AES_CORE_DATAPATH__abc_16259_n4666;
  wire AES_CORE_DATAPATH__abc_16259_n4667;
  wire AES_CORE_DATAPATH__abc_16259_n4669;
  wire AES_CORE_DATAPATH__abc_16259_n4670;
  wire AES_CORE_DATAPATH__abc_16259_n4671;
  wire AES_CORE_DATAPATH__abc_16259_n4672;
  wire AES_CORE_DATAPATH__abc_16259_n4673;
  wire AES_CORE_DATAPATH__abc_16259_n4674;
  wire AES_CORE_DATAPATH__abc_16259_n4675_1;
  wire AES_CORE_DATAPATH__abc_16259_n4676;
  wire AES_CORE_DATAPATH__abc_16259_n4678;
  wire AES_CORE_DATAPATH__abc_16259_n4679;
  wire AES_CORE_DATAPATH__abc_16259_n4680;
  wire AES_CORE_DATAPATH__abc_16259_n4681_1;
  wire AES_CORE_DATAPATH__abc_16259_n4682;
  wire AES_CORE_DATAPATH__abc_16259_n4683;
  wire AES_CORE_DATAPATH__abc_16259_n4684;
  wire AES_CORE_DATAPATH__abc_16259_n4685;
  wire AES_CORE_DATAPATH__abc_16259_n4687;
  wire AES_CORE_DATAPATH__abc_16259_n4688;
  wire AES_CORE_DATAPATH__abc_16259_n4689_1;
  wire AES_CORE_DATAPATH__abc_16259_n4690;
  wire AES_CORE_DATAPATH__abc_16259_n4691;
  wire AES_CORE_DATAPATH__abc_16259_n4692;
  wire AES_CORE_DATAPATH__abc_16259_n4693;
  wire AES_CORE_DATAPATH__abc_16259_n4694;
  wire AES_CORE_DATAPATH__abc_16259_n4696;
  wire AES_CORE_DATAPATH__abc_16259_n4697;
  wire AES_CORE_DATAPATH__abc_16259_n4698;
  wire AES_CORE_DATAPATH__abc_16259_n4699;
  wire AES_CORE_DATAPATH__abc_16259_n4700;
  wire AES_CORE_DATAPATH__abc_16259_n4701;
  wire AES_CORE_DATAPATH__abc_16259_n4702_1;
  wire AES_CORE_DATAPATH__abc_16259_n4703;
  wire AES_CORE_DATAPATH__abc_16259_n4705;
  wire AES_CORE_DATAPATH__abc_16259_n4706;
  wire AES_CORE_DATAPATH__abc_16259_n4707;
  wire AES_CORE_DATAPATH__abc_16259_n4708_1;
  wire AES_CORE_DATAPATH__abc_16259_n4709;
  wire AES_CORE_DATAPATH__abc_16259_n4710;
  wire AES_CORE_DATAPATH__abc_16259_n4711;
  wire AES_CORE_DATAPATH__abc_16259_n4712;
  wire AES_CORE_DATAPATH__abc_16259_n4714;
  wire AES_CORE_DATAPATH__abc_16259_n4715;
  wire AES_CORE_DATAPATH__abc_16259_n4716;
  wire AES_CORE_DATAPATH__abc_16259_n4717_1;
  wire AES_CORE_DATAPATH__abc_16259_n4718;
  wire AES_CORE_DATAPATH__abc_16259_n4719;
  wire AES_CORE_DATAPATH__abc_16259_n4720;
  wire AES_CORE_DATAPATH__abc_16259_n4721;
  wire AES_CORE_DATAPATH__abc_16259_n4723_1;
  wire AES_CORE_DATAPATH__abc_16259_n4724;
  wire AES_CORE_DATAPATH__abc_16259_n4725;
  wire AES_CORE_DATAPATH__abc_16259_n4726;
  wire AES_CORE_DATAPATH__abc_16259_n4727;
  wire AES_CORE_DATAPATH__abc_16259_n4728;
  wire AES_CORE_DATAPATH__abc_16259_n4729;
  wire AES_CORE_DATAPATH__abc_16259_n4730_1;
  wire AES_CORE_DATAPATH__abc_16259_n4732;
  wire AES_CORE_DATAPATH__abc_16259_n4733;
  wire AES_CORE_DATAPATH__abc_16259_n4734;
  wire AES_CORE_DATAPATH__abc_16259_n4735;
  wire AES_CORE_DATAPATH__abc_16259_n4736_1;
  wire AES_CORE_DATAPATH__abc_16259_n4737;
  wire AES_CORE_DATAPATH__abc_16259_n4738;
  wire AES_CORE_DATAPATH__abc_16259_n4739;
  wire AES_CORE_DATAPATH__abc_16259_n4741;
  wire AES_CORE_DATAPATH__abc_16259_n4742;
  wire AES_CORE_DATAPATH__abc_16259_n4743;
  wire AES_CORE_DATAPATH__abc_16259_n4744_1;
  wire AES_CORE_DATAPATH__abc_16259_n4745;
  wire AES_CORE_DATAPATH__abc_16259_n4746;
  wire AES_CORE_DATAPATH__abc_16259_n4747;
  wire AES_CORE_DATAPATH__abc_16259_n4748;
  wire AES_CORE_DATAPATH__abc_16259_n4750_1;
  wire AES_CORE_DATAPATH__abc_16259_n4751;
  wire AES_CORE_DATAPATH__abc_16259_n4752;
  wire AES_CORE_DATAPATH__abc_16259_n4753;
  wire AES_CORE_DATAPATH__abc_16259_n4754;
  wire AES_CORE_DATAPATH__abc_16259_n4755;
  wire AES_CORE_DATAPATH__abc_16259_n4756;
  wire AES_CORE_DATAPATH__abc_16259_n4757_1;
  wire AES_CORE_DATAPATH__abc_16259_n4759;
  wire AES_CORE_DATAPATH__abc_16259_n4760;
  wire AES_CORE_DATAPATH__abc_16259_n4761;
  wire AES_CORE_DATAPATH__abc_16259_n4762;
  wire AES_CORE_DATAPATH__abc_16259_n4763_1;
  wire AES_CORE_DATAPATH__abc_16259_n4764;
  wire AES_CORE_DATAPATH__abc_16259_n4765;
  wire AES_CORE_DATAPATH__abc_16259_n4766;
  wire AES_CORE_DATAPATH__abc_16259_n4768;
  wire AES_CORE_DATAPATH__abc_16259_n4769;
  wire AES_CORE_DATAPATH__abc_16259_n4769_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n4769_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n4769_bF_buf10;
  wire AES_CORE_DATAPATH__abc_16259_n4769_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n4769_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n4769_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n4769_bF_buf5;
  wire AES_CORE_DATAPATH__abc_16259_n4769_bF_buf6;
  wire AES_CORE_DATAPATH__abc_16259_n4769_bF_buf7;
  wire AES_CORE_DATAPATH__abc_16259_n4769_bF_buf8;
  wire AES_CORE_DATAPATH__abc_16259_n4769_bF_buf9;
  wire AES_CORE_DATAPATH__abc_16259_n4770;
  wire AES_CORE_DATAPATH__abc_16259_n4772_1;
  wire AES_CORE_DATAPATH__abc_16259_n4773;
  wire AES_CORE_DATAPATH__abc_16259_n4775;
  wire AES_CORE_DATAPATH__abc_16259_n4776;
  wire AES_CORE_DATAPATH__abc_16259_n4778_1;
  wire AES_CORE_DATAPATH__abc_16259_n4779;
  wire AES_CORE_DATAPATH__abc_16259_n4781;
  wire AES_CORE_DATAPATH__abc_16259_n4782;
  wire AES_CORE_DATAPATH__abc_16259_n4784;
  wire AES_CORE_DATAPATH__abc_16259_n4785_1;
  wire AES_CORE_DATAPATH__abc_16259_n4787;
  wire AES_CORE_DATAPATH__abc_16259_n4788;
  wire AES_CORE_DATAPATH__abc_16259_n4790;
  wire AES_CORE_DATAPATH__abc_16259_n4791_1;
  wire AES_CORE_DATAPATH__abc_16259_n4793;
  wire AES_CORE_DATAPATH__abc_16259_n4794;
  wire AES_CORE_DATAPATH__abc_16259_n4796;
  wire AES_CORE_DATAPATH__abc_16259_n4797;
  wire AES_CORE_DATAPATH__abc_16259_n4799_1;
  wire AES_CORE_DATAPATH__abc_16259_n4800;
  wire AES_CORE_DATAPATH__abc_16259_n4802;
  wire AES_CORE_DATAPATH__abc_16259_n4803;
  wire AES_CORE_DATAPATH__abc_16259_n4805_1;
  wire AES_CORE_DATAPATH__abc_16259_n4806;
  wire AES_CORE_DATAPATH__abc_16259_n4808;
  wire AES_CORE_DATAPATH__abc_16259_n4809;
  wire AES_CORE_DATAPATH__abc_16259_n4811;
  wire AES_CORE_DATAPATH__abc_16259_n4812_1;
  wire AES_CORE_DATAPATH__abc_16259_n4814;
  wire AES_CORE_DATAPATH__abc_16259_n4815;
  wire AES_CORE_DATAPATH__abc_16259_n4817;
  wire AES_CORE_DATAPATH__abc_16259_n4818_1;
  wire AES_CORE_DATAPATH__abc_16259_n4820_1;
  wire AES_CORE_DATAPATH__abc_16259_n4821_1;
  wire AES_CORE_DATAPATH__abc_16259_n4823_1;
  wire AES_CORE_DATAPATH__abc_16259_n4824_1;
  wire AES_CORE_DATAPATH__abc_16259_n4826_1;
  wire AES_CORE_DATAPATH__abc_16259_n4827_1;
  wire AES_CORE_DATAPATH__abc_16259_n4829_1;
  wire AES_CORE_DATAPATH__abc_16259_n4830_1;
  wire AES_CORE_DATAPATH__abc_16259_n4832_1;
  wire AES_CORE_DATAPATH__abc_16259_n4833_1;
  wire AES_CORE_DATAPATH__abc_16259_n4835_1;
  wire AES_CORE_DATAPATH__abc_16259_n4836_1;
  wire AES_CORE_DATAPATH__abc_16259_n4838_1;
  wire AES_CORE_DATAPATH__abc_16259_n4839_1;
  wire AES_CORE_DATAPATH__abc_16259_n4841_1;
  wire AES_CORE_DATAPATH__abc_16259_n4842_1;
  wire AES_CORE_DATAPATH__abc_16259_n4844_1;
  wire AES_CORE_DATAPATH__abc_16259_n4845_1;
  wire AES_CORE_DATAPATH__abc_16259_n4847_1;
  wire AES_CORE_DATAPATH__abc_16259_n4848_1;
  wire AES_CORE_DATAPATH__abc_16259_n4850_1;
  wire AES_CORE_DATAPATH__abc_16259_n4851_1;
  wire AES_CORE_DATAPATH__abc_16259_n4853_1;
  wire AES_CORE_DATAPATH__abc_16259_n4854_1;
  wire AES_CORE_DATAPATH__abc_16259_n4856_1;
  wire AES_CORE_DATAPATH__abc_16259_n4857_1;
  wire AES_CORE_DATAPATH__abc_16259_n4859_1;
  wire AES_CORE_DATAPATH__abc_16259_n4860_1;
  wire AES_CORE_DATAPATH__abc_16259_n4862_1;
  wire AES_CORE_DATAPATH__abc_16259_n4863_1;
  wire AES_CORE_DATAPATH__abc_16259_n4865_1;
  wire AES_CORE_DATAPATH__abc_16259_n4866_1;
  wire AES_CORE_DATAPATH__abc_16259_n4867_1;
  wire AES_CORE_DATAPATH__abc_16259_n4867_1_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n4867_1_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n4867_1_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n4867_1_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n4867_1_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n4868_1;
  wire AES_CORE_DATAPATH__abc_16259_n4869_1;
  wire AES_CORE_DATAPATH__abc_16259_n4870_1;
  wire AES_CORE_DATAPATH__abc_16259_n4871_1;
  wire AES_CORE_DATAPATH__abc_16259_n4872_1;
  wire AES_CORE_DATAPATH__abc_16259_n4872_1_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n4872_1_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n4872_1_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n4872_1_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n4872_1_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n4873_1;
  wire AES_CORE_DATAPATH__abc_16259_n4873_1_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n4873_1_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n4873_1_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n4873_1_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n4873_1_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n4874_1;
  wire AES_CORE_DATAPATH__abc_16259_n4875_1;
  wire AES_CORE_DATAPATH__abc_16259_n4876_1;
  wire AES_CORE_DATAPATH__abc_16259_n4877_1;
  wire AES_CORE_DATAPATH__abc_16259_n4878_1;
  wire AES_CORE_DATAPATH__abc_16259_n4879_1;
  wire AES_CORE_DATAPATH__abc_16259_n4880_1;
  wire AES_CORE_DATAPATH__abc_16259_n4881_1;
  wire AES_CORE_DATAPATH__abc_16259_n4883_1;
  wire AES_CORE_DATAPATH__abc_16259_n4884;
  wire AES_CORE_DATAPATH__abc_16259_n4885;
  wire AES_CORE_DATAPATH__abc_16259_n4886_1;
  wire AES_CORE_DATAPATH__abc_16259_n4887;
  wire AES_CORE_DATAPATH__abc_16259_n4888;
  wire AES_CORE_DATAPATH__abc_16259_n4889_1;
  wire AES_CORE_DATAPATH__abc_16259_n4890;
  wire AES_CORE_DATAPATH__abc_16259_n4892_1;
  wire AES_CORE_DATAPATH__abc_16259_n4893;
  wire AES_CORE_DATAPATH__abc_16259_n4894;
  wire AES_CORE_DATAPATH__abc_16259_n4895_1;
  wire AES_CORE_DATAPATH__abc_16259_n4896;
  wire AES_CORE_DATAPATH__abc_16259_n4897;
  wire AES_CORE_DATAPATH__abc_16259_n4898_1;
  wire AES_CORE_DATAPATH__abc_16259_n4899;
  wire AES_CORE_DATAPATH__abc_16259_n4901_1;
  wire AES_CORE_DATAPATH__abc_16259_n4902;
  wire AES_CORE_DATAPATH__abc_16259_n4903;
  wire AES_CORE_DATAPATH__abc_16259_n4904_1;
  wire AES_CORE_DATAPATH__abc_16259_n4905;
  wire AES_CORE_DATAPATH__abc_16259_n4906;
  wire AES_CORE_DATAPATH__abc_16259_n4907_1;
  wire AES_CORE_DATAPATH__abc_16259_n4908;
  wire AES_CORE_DATAPATH__abc_16259_n4910_1;
  wire AES_CORE_DATAPATH__abc_16259_n4911;
  wire AES_CORE_DATAPATH__abc_16259_n4912;
  wire AES_CORE_DATAPATH__abc_16259_n4913_1;
  wire AES_CORE_DATAPATH__abc_16259_n4914;
  wire AES_CORE_DATAPATH__abc_16259_n4915;
  wire AES_CORE_DATAPATH__abc_16259_n4916_1;
  wire AES_CORE_DATAPATH__abc_16259_n4917;
  wire AES_CORE_DATAPATH__abc_16259_n4919_1;
  wire AES_CORE_DATAPATH__abc_16259_n4920;
  wire AES_CORE_DATAPATH__abc_16259_n4921;
  wire AES_CORE_DATAPATH__abc_16259_n4922_1;
  wire AES_CORE_DATAPATH__abc_16259_n4923;
  wire AES_CORE_DATAPATH__abc_16259_n4924;
  wire AES_CORE_DATAPATH__abc_16259_n4925_1;
  wire AES_CORE_DATAPATH__abc_16259_n4926;
  wire AES_CORE_DATAPATH__abc_16259_n4928_1;
  wire AES_CORE_DATAPATH__abc_16259_n4929;
  wire AES_CORE_DATAPATH__abc_16259_n4930;
  wire AES_CORE_DATAPATH__abc_16259_n4931_1;
  wire AES_CORE_DATAPATH__abc_16259_n4932;
  wire AES_CORE_DATAPATH__abc_16259_n4933;
  wire AES_CORE_DATAPATH__abc_16259_n4934_1;
  wire AES_CORE_DATAPATH__abc_16259_n4935;
  wire AES_CORE_DATAPATH__abc_16259_n4937_1;
  wire AES_CORE_DATAPATH__abc_16259_n4938;
  wire AES_CORE_DATAPATH__abc_16259_n4939;
  wire AES_CORE_DATAPATH__abc_16259_n4940_1;
  wire AES_CORE_DATAPATH__abc_16259_n4941;
  wire AES_CORE_DATAPATH__abc_16259_n4942;
  wire AES_CORE_DATAPATH__abc_16259_n4943_1;
  wire AES_CORE_DATAPATH__abc_16259_n4944;
  wire AES_CORE_DATAPATH__abc_16259_n4946_1;
  wire AES_CORE_DATAPATH__abc_16259_n4947;
  wire AES_CORE_DATAPATH__abc_16259_n4948;
  wire AES_CORE_DATAPATH__abc_16259_n4949_1;
  wire AES_CORE_DATAPATH__abc_16259_n4950;
  wire AES_CORE_DATAPATH__abc_16259_n4951;
  wire AES_CORE_DATAPATH__abc_16259_n4952_1;
  wire AES_CORE_DATAPATH__abc_16259_n4953;
  wire AES_CORE_DATAPATH__abc_16259_n4955_1;
  wire AES_CORE_DATAPATH__abc_16259_n4956;
  wire AES_CORE_DATAPATH__abc_16259_n4957;
  wire AES_CORE_DATAPATH__abc_16259_n4958_1;
  wire AES_CORE_DATAPATH__abc_16259_n4959;
  wire AES_CORE_DATAPATH__abc_16259_n4960;
  wire AES_CORE_DATAPATH__abc_16259_n4961_1;
  wire AES_CORE_DATAPATH__abc_16259_n4962;
  wire AES_CORE_DATAPATH__abc_16259_n4964_1;
  wire AES_CORE_DATAPATH__abc_16259_n4965;
  wire AES_CORE_DATAPATH__abc_16259_n4966;
  wire AES_CORE_DATAPATH__abc_16259_n4967_1;
  wire AES_CORE_DATAPATH__abc_16259_n4968;
  wire AES_CORE_DATAPATH__abc_16259_n4969;
  wire AES_CORE_DATAPATH__abc_16259_n4970_1;
  wire AES_CORE_DATAPATH__abc_16259_n4971;
  wire AES_CORE_DATAPATH__abc_16259_n4973_1;
  wire AES_CORE_DATAPATH__abc_16259_n4974;
  wire AES_CORE_DATAPATH__abc_16259_n4975;
  wire AES_CORE_DATAPATH__abc_16259_n4976_1;
  wire AES_CORE_DATAPATH__abc_16259_n4977;
  wire AES_CORE_DATAPATH__abc_16259_n4978;
  wire AES_CORE_DATAPATH__abc_16259_n4979_1;
  wire AES_CORE_DATAPATH__abc_16259_n4980_1;
  wire AES_CORE_DATAPATH__abc_16259_n4982_1;
  wire AES_CORE_DATAPATH__abc_16259_n4983_1;
  wire AES_CORE_DATAPATH__abc_16259_n4984_1;
  wire AES_CORE_DATAPATH__abc_16259_n4985_1;
  wire AES_CORE_DATAPATH__abc_16259_n4986_1;
  wire AES_CORE_DATAPATH__abc_16259_n4987_1;
  wire AES_CORE_DATAPATH__abc_16259_n4988_1;
  wire AES_CORE_DATAPATH__abc_16259_n4989_1;
  wire AES_CORE_DATAPATH__abc_16259_n4991_1;
  wire AES_CORE_DATAPATH__abc_16259_n4992_1;
  wire AES_CORE_DATAPATH__abc_16259_n4993_1;
  wire AES_CORE_DATAPATH__abc_16259_n4994_1;
  wire AES_CORE_DATAPATH__abc_16259_n4995_1;
  wire AES_CORE_DATAPATH__abc_16259_n4996_1;
  wire AES_CORE_DATAPATH__abc_16259_n4997_1;
  wire AES_CORE_DATAPATH__abc_16259_n4998_1;
  wire AES_CORE_DATAPATH__abc_16259_n5000_1;
  wire AES_CORE_DATAPATH__abc_16259_n5001_1;
  wire AES_CORE_DATAPATH__abc_16259_n5002_1;
  wire AES_CORE_DATAPATH__abc_16259_n5003_1;
  wire AES_CORE_DATAPATH__abc_16259_n5004_1;
  wire AES_CORE_DATAPATH__abc_16259_n5005_1;
  wire AES_CORE_DATAPATH__abc_16259_n5006_1;
  wire AES_CORE_DATAPATH__abc_16259_n5007_1;
  wire AES_CORE_DATAPATH__abc_16259_n5009_1;
  wire AES_CORE_DATAPATH__abc_16259_n5010_1;
  wire AES_CORE_DATAPATH__abc_16259_n5011_1;
  wire AES_CORE_DATAPATH__abc_16259_n5012_1;
  wire AES_CORE_DATAPATH__abc_16259_n5013;
  wire AES_CORE_DATAPATH__abc_16259_n5014_1;
  wire AES_CORE_DATAPATH__abc_16259_n5015_1;
  wire AES_CORE_DATAPATH__abc_16259_n5016_1;
  wire AES_CORE_DATAPATH__abc_16259_n5018_1;
  wire AES_CORE_DATAPATH__abc_16259_n5019_1;
  wire AES_CORE_DATAPATH__abc_16259_n5020_1;
  wire AES_CORE_DATAPATH__abc_16259_n5021_1;
  wire AES_CORE_DATAPATH__abc_16259_n5022_1;
  wire AES_CORE_DATAPATH__abc_16259_n5023_1;
  wire AES_CORE_DATAPATH__abc_16259_n5024_1;
  wire AES_CORE_DATAPATH__abc_16259_n5025_1;
  wire AES_CORE_DATAPATH__abc_16259_n5027_1;
  wire AES_CORE_DATAPATH__abc_16259_n5028_1;
  wire AES_CORE_DATAPATH__abc_16259_n5029_1;
  wire AES_CORE_DATAPATH__abc_16259_n5030_1;
  wire AES_CORE_DATAPATH__abc_16259_n5031_1;
  wire AES_CORE_DATAPATH__abc_16259_n5032_1;
  wire AES_CORE_DATAPATH__abc_16259_n5033_1;
  wire AES_CORE_DATAPATH__abc_16259_n5034_1;
  wire AES_CORE_DATAPATH__abc_16259_n5036_1;
  wire AES_CORE_DATAPATH__abc_16259_n5037_1;
  wire AES_CORE_DATAPATH__abc_16259_n5038_1;
  wire AES_CORE_DATAPATH__abc_16259_n5039_1;
  wire AES_CORE_DATAPATH__abc_16259_n5040_1;
  wire AES_CORE_DATAPATH__abc_16259_n5041_1;
  wire AES_CORE_DATAPATH__abc_16259_n5042_1;
  wire AES_CORE_DATAPATH__abc_16259_n5043_1;
  wire AES_CORE_DATAPATH__abc_16259_n5045_1;
  wire AES_CORE_DATAPATH__abc_16259_n5046_1;
  wire AES_CORE_DATAPATH__abc_16259_n5047_1;
  wire AES_CORE_DATAPATH__abc_16259_n5048_1;
  wire AES_CORE_DATAPATH__abc_16259_n5049_1;
  wire AES_CORE_DATAPATH__abc_16259_n5050_1;
  wire AES_CORE_DATAPATH__abc_16259_n5051_1;
  wire AES_CORE_DATAPATH__abc_16259_n5052_1;
  wire AES_CORE_DATAPATH__abc_16259_n5054_1;
  wire AES_CORE_DATAPATH__abc_16259_n5055_1;
  wire AES_CORE_DATAPATH__abc_16259_n5056_1;
  wire AES_CORE_DATAPATH__abc_16259_n5057_1;
  wire AES_CORE_DATAPATH__abc_16259_n5058_1;
  wire AES_CORE_DATAPATH__abc_16259_n5059_1;
  wire AES_CORE_DATAPATH__abc_16259_n5060_1;
  wire AES_CORE_DATAPATH__abc_16259_n5061_1;
  wire AES_CORE_DATAPATH__abc_16259_n5063_1;
  wire AES_CORE_DATAPATH__abc_16259_n5064_1;
  wire AES_CORE_DATAPATH__abc_16259_n5065_1;
  wire AES_CORE_DATAPATH__abc_16259_n5066_1;
  wire AES_CORE_DATAPATH__abc_16259_n5067_1;
  wire AES_CORE_DATAPATH__abc_16259_n5068_1;
  wire AES_CORE_DATAPATH__abc_16259_n5069_1;
  wire AES_CORE_DATAPATH__abc_16259_n5070_1;
  wire AES_CORE_DATAPATH__abc_16259_n5072_1;
  wire AES_CORE_DATAPATH__abc_16259_n5073_1;
  wire AES_CORE_DATAPATH__abc_16259_n5074_1;
  wire AES_CORE_DATAPATH__abc_16259_n5075_1;
  wire AES_CORE_DATAPATH__abc_16259_n5076_1;
  wire AES_CORE_DATAPATH__abc_16259_n5077_1;
  wire AES_CORE_DATAPATH__abc_16259_n5078;
  wire AES_CORE_DATAPATH__abc_16259_n5079;
  wire AES_CORE_DATAPATH__abc_16259_n5081;
  wire AES_CORE_DATAPATH__abc_16259_n5082;
  wire AES_CORE_DATAPATH__abc_16259_n5083_1;
  wire AES_CORE_DATAPATH__abc_16259_n5084;
  wire AES_CORE_DATAPATH__abc_16259_n5085;
  wire AES_CORE_DATAPATH__abc_16259_n5086_1;
  wire AES_CORE_DATAPATH__abc_16259_n5087;
  wire AES_CORE_DATAPATH__abc_16259_n5088;
  wire AES_CORE_DATAPATH__abc_16259_n5090;
  wire AES_CORE_DATAPATH__abc_16259_n5091;
  wire AES_CORE_DATAPATH__abc_16259_n5092_1;
  wire AES_CORE_DATAPATH__abc_16259_n5093;
  wire AES_CORE_DATAPATH__abc_16259_n5094;
  wire AES_CORE_DATAPATH__abc_16259_n5095_1;
  wire AES_CORE_DATAPATH__abc_16259_n5096;
  wire AES_CORE_DATAPATH__abc_16259_n5097;
  wire AES_CORE_DATAPATH__abc_16259_n5099;
  wire AES_CORE_DATAPATH__abc_16259_n5100;
  wire AES_CORE_DATAPATH__abc_16259_n5101_1;
  wire AES_CORE_DATAPATH__abc_16259_n5102;
  wire AES_CORE_DATAPATH__abc_16259_n5103;
  wire AES_CORE_DATAPATH__abc_16259_n5104_1;
  wire AES_CORE_DATAPATH__abc_16259_n5105;
  wire AES_CORE_DATAPATH__abc_16259_n5106;
  wire AES_CORE_DATAPATH__abc_16259_n5108;
  wire AES_CORE_DATAPATH__abc_16259_n5109;
  wire AES_CORE_DATAPATH__abc_16259_n5110_1;
  wire AES_CORE_DATAPATH__abc_16259_n5111;
  wire AES_CORE_DATAPATH__abc_16259_n5112;
  wire AES_CORE_DATAPATH__abc_16259_n5113_1;
  wire AES_CORE_DATAPATH__abc_16259_n5114;
  wire AES_CORE_DATAPATH__abc_16259_n5115;
  wire AES_CORE_DATAPATH__abc_16259_n5117;
  wire AES_CORE_DATAPATH__abc_16259_n5118;
  wire AES_CORE_DATAPATH__abc_16259_n5119_1;
  wire AES_CORE_DATAPATH__abc_16259_n5120;
  wire AES_CORE_DATAPATH__abc_16259_n5121;
  wire AES_CORE_DATAPATH__abc_16259_n5122_1;
  wire AES_CORE_DATAPATH__abc_16259_n5123;
  wire AES_CORE_DATAPATH__abc_16259_n5124;
  wire AES_CORE_DATAPATH__abc_16259_n5126;
  wire AES_CORE_DATAPATH__abc_16259_n5127;
  wire AES_CORE_DATAPATH__abc_16259_n5128_1;
  wire AES_CORE_DATAPATH__abc_16259_n5129;
  wire AES_CORE_DATAPATH__abc_16259_n5130;
  wire AES_CORE_DATAPATH__abc_16259_n5131_1;
  wire AES_CORE_DATAPATH__abc_16259_n5132;
  wire AES_CORE_DATAPATH__abc_16259_n5133;
  wire AES_CORE_DATAPATH__abc_16259_n5135;
  wire AES_CORE_DATAPATH__abc_16259_n5136;
  wire AES_CORE_DATAPATH__abc_16259_n5137_1;
  wire AES_CORE_DATAPATH__abc_16259_n5138;
  wire AES_CORE_DATAPATH__abc_16259_n5139;
  wire AES_CORE_DATAPATH__abc_16259_n5140_1;
  wire AES_CORE_DATAPATH__abc_16259_n5141;
  wire AES_CORE_DATAPATH__abc_16259_n5142;
  wire AES_CORE_DATAPATH__abc_16259_n5144;
  wire AES_CORE_DATAPATH__abc_16259_n5145;
  wire AES_CORE_DATAPATH__abc_16259_n5146_1;
  wire AES_CORE_DATAPATH__abc_16259_n5147;
  wire AES_CORE_DATAPATH__abc_16259_n5148;
  wire AES_CORE_DATAPATH__abc_16259_n5149_1;
  wire AES_CORE_DATAPATH__abc_16259_n5150;
  wire AES_CORE_DATAPATH__abc_16259_n5151;
  wire AES_CORE_DATAPATH__abc_16259_n5153;
  wire AES_CORE_DATAPATH__abc_16259_n5154;
  wire AES_CORE_DATAPATH__abc_16259_n5155_1;
  wire AES_CORE_DATAPATH__abc_16259_n5156;
  wire AES_CORE_DATAPATH__abc_16259_n5157;
  wire AES_CORE_DATAPATH__abc_16259_n5158_1;
  wire AES_CORE_DATAPATH__abc_16259_n5159;
  wire AES_CORE_DATAPATH__abc_16259_n5160;
  wire AES_CORE_DATAPATH__abc_16259_n5162;
  wire AES_CORE_DATAPATH__abc_16259_n5163;
  wire AES_CORE_DATAPATH__abc_16259_n5165;
  wire AES_CORE_DATAPATH__abc_16259_n5166;
  wire AES_CORE_DATAPATH__abc_16259_n5168;
  wire AES_CORE_DATAPATH__abc_16259_n5169;
  wire AES_CORE_DATAPATH__abc_16259_n5171;
  wire AES_CORE_DATAPATH__abc_16259_n5172;
  wire AES_CORE_DATAPATH__abc_16259_n5174_1;
  wire AES_CORE_DATAPATH__abc_16259_n5175_1;
  wire AES_CORE_DATAPATH__abc_16259_n5177_1;
  wire AES_CORE_DATAPATH__abc_16259_n5178_1;
  wire AES_CORE_DATAPATH__abc_16259_n5180_1;
  wire AES_CORE_DATAPATH__abc_16259_n5181_1;
  wire AES_CORE_DATAPATH__abc_16259_n5183_1;
  wire AES_CORE_DATAPATH__abc_16259_n5184_1;
  wire AES_CORE_DATAPATH__abc_16259_n5186_1;
  wire AES_CORE_DATAPATH__abc_16259_n5187_1;
  wire AES_CORE_DATAPATH__abc_16259_n5189_1;
  wire AES_CORE_DATAPATH__abc_16259_n5190_1;
  wire AES_CORE_DATAPATH__abc_16259_n5192_1;
  wire AES_CORE_DATAPATH__abc_16259_n5193_1;
  wire AES_CORE_DATAPATH__abc_16259_n5195_1;
  wire AES_CORE_DATAPATH__abc_16259_n5196_1;
  wire AES_CORE_DATAPATH__abc_16259_n5198_1;
  wire AES_CORE_DATAPATH__abc_16259_n5199_1;
  wire AES_CORE_DATAPATH__abc_16259_n5201_1;
  wire AES_CORE_DATAPATH__abc_16259_n5202_1;
  wire AES_CORE_DATAPATH__abc_16259_n5204_1;
  wire AES_CORE_DATAPATH__abc_16259_n5205_1;
  wire AES_CORE_DATAPATH__abc_16259_n5207;
  wire AES_CORE_DATAPATH__abc_16259_n5208_1;
  wire AES_CORE_DATAPATH__abc_16259_n5210_1;
  wire AES_CORE_DATAPATH__abc_16259_n5211_1;
  wire AES_CORE_DATAPATH__abc_16259_n5213_1;
  wire AES_CORE_DATAPATH__abc_16259_n5214_1;
  wire AES_CORE_DATAPATH__abc_16259_n5216_1;
  wire AES_CORE_DATAPATH__abc_16259_n5217_1;
  wire AES_CORE_DATAPATH__abc_16259_n5219_1;
  wire AES_CORE_DATAPATH__abc_16259_n5220_1;
  wire AES_CORE_DATAPATH__abc_16259_n5222_1;
  wire AES_CORE_DATAPATH__abc_16259_n5223_1;
  wire AES_CORE_DATAPATH__abc_16259_n5225_1;
  wire AES_CORE_DATAPATH__abc_16259_n5226_1;
  wire AES_CORE_DATAPATH__abc_16259_n5228_1;
  wire AES_CORE_DATAPATH__abc_16259_n5229_1;
  wire AES_CORE_DATAPATH__abc_16259_n5231_1;
  wire AES_CORE_DATAPATH__abc_16259_n5232_1;
  wire AES_CORE_DATAPATH__abc_16259_n5234_1;
  wire AES_CORE_DATAPATH__abc_16259_n5235_1;
  wire AES_CORE_DATAPATH__abc_16259_n5237_1;
  wire AES_CORE_DATAPATH__abc_16259_n5238_1;
  wire AES_CORE_DATAPATH__abc_16259_n5240_1;
  wire AES_CORE_DATAPATH__abc_16259_n5241_1;
  wire AES_CORE_DATAPATH__abc_16259_n5243_1;
  wire AES_CORE_DATAPATH__abc_16259_n5244_1;
  wire AES_CORE_DATAPATH__abc_16259_n5246_1;
  wire AES_CORE_DATAPATH__abc_16259_n5247_1;
  wire AES_CORE_DATAPATH__abc_16259_n5249_1;
  wire AES_CORE_DATAPATH__abc_16259_n5250_1;
  wire AES_CORE_DATAPATH__abc_16259_n5252_1;
  wire AES_CORE_DATAPATH__abc_16259_n5253_1;
  wire AES_CORE_DATAPATH__abc_16259_n5255_1;
  wire AES_CORE_DATAPATH__abc_16259_n5256_1;
  wire AES_CORE_DATAPATH__abc_16259_n5258_1;
  wire AES_CORE_DATAPATH__abc_16259_n5259_1;
  wire AES_CORE_DATAPATH__abc_16259_n5260_1;
  wire AES_CORE_DATAPATH__abc_16259_n5260_1_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n5260_1_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n5260_1_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n5260_1_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n5260_1_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n5261_1;
  wire AES_CORE_DATAPATH__abc_16259_n5262_1;
  wire AES_CORE_DATAPATH__abc_16259_n5263_1;
  wire AES_CORE_DATAPATH__abc_16259_n5264_1;
  wire AES_CORE_DATAPATH__abc_16259_n5265_1;
  wire AES_CORE_DATAPATH__abc_16259_n5265_1_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n5265_1_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n5265_1_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n5265_1_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n5265_1_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n5266_1;
  wire AES_CORE_DATAPATH__abc_16259_n5266_1_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n5266_1_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n5266_1_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n5266_1_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n5266_1_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n5267_1;
  wire AES_CORE_DATAPATH__abc_16259_n5268_1;
  wire AES_CORE_DATAPATH__abc_16259_n5269_1;
  wire AES_CORE_DATAPATH__abc_16259_n5270_1;
  wire AES_CORE_DATAPATH__abc_16259_n5271_1;
  wire AES_CORE_DATAPATH__abc_16259_n5272;
  wire AES_CORE_DATAPATH__abc_16259_n5273;
  wire AES_CORE_DATAPATH__abc_16259_n5274_1;
  wire AES_CORE_DATAPATH__abc_16259_n5276;
  wire AES_CORE_DATAPATH__abc_16259_n5277_1;
  wire AES_CORE_DATAPATH__abc_16259_n5278;
  wire AES_CORE_DATAPATH__abc_16259_n5279;
  wire AES_CORE_DATAPATH__abc_16259_n5280_1;
  wire AES_CORE_DATAPATH__abc_16259_n5281;
  wire AES_CORE_DATAPATH__abc_16259_n5282;
  wire AES_CORE_DATAPATH__abc_16259_n5283_1;
  wire AES_CORE_DATAPATH__abc_16259_n5285;
  wire AES_CORE_DATAPATH__abc_16259_n5286_1;
  wire AES_CORE_DATAPATH__abc_16259_n5287;
  wire AES_CORE_DATAPATH__abc_16259_n5288;
  wire AES_CORE_DATAPATH__abc_16259_n5289_1;
  wire AES_CORE_DATAPATH__abc_16259_n5290;
  wire AES_CORE_DATAPATH__abc_16259_n5291;
  wire AES_CORE_DATAPATH__abc_16259_n5292_1;
  wire AES_CORE_DATAPATH__abc_16259_n5294;
  wire AES_CORE_DATAPATH__abc_16259_n5295_1;
  wire AES_CORE_DATAPATH__abc_16259_n5296;
  wire AES_CORE_DATAPATH__abc_16259_n5297;
  wire AES_CORE_DATAPATH__abc_16259_n5298_1;
  wire AES_CORE_DATAPATH__abc_16259_n5299;
  wire AES_CORE_DATAPATH__abc_16259_n5300;
  wire AES_CORE_DATAPATH__abc_16259_n5301_1;
  wire AES_CORE_DATAPATH__abc_16259_n5303;
  wire AES_CORE_DATAPATH__abc_16259_n5304_1;
  wire AES_CORE_DATAPATH__abc_16259_n5305;
  wire AES_CORE_DATAPATH__abc_16259_n5306;
  wire AES_CORE_DATAPATH__abc_16259_n5307_1;
  wire AES_CORE_DATAPATH__abc_16259_n5308;
  wire AES_CORE_DATAPATH__abc_16259_n5309;
  wire AES_CORE_DATAPATH__abc_16259_n5310_1;
  wire AES_CORE_DATAPATH__abc_16259_n5312;
  wire AES_CORE_DATAPATH__abc_16259_n5313_1;
  wire AES_CORE_DATAPATH__abc_16259_n5314;
  wire AES_CORE_DATAPATH__abc_16259_n5315;
  wire AES_CORE_DATAPATH__abc_16259_n5316_1;
  wire AES_CORE_DATAPATH__abc_16259_n5317;
  wire AES_CORE_DATAPATH__abc_16259_n5318;
  wire AES_CORE_DATAPATH__abc_16259_n5319_1;
  wire AES_CORE_DATAPATH__abc_16259_n5321;
  wire AES_CORE_DATAPATH__abc_16259_n5322_1;
  wire AES_CORE_DATAPATH__abc_16259_n5323;
  wire AES_CORE_DATAPATH__abc_16259_n5324;
  wire AES_CORE_DATAPATH__abc_16259_n5325_1;
  wire AES_CORE_DATAPATH__abc_16259_n5326;
  wire AES_CORE_DATAPATH__abc_16259_n5327;
  wire AES_CORE_DATAPATH__abc_16259_n5328_1;
  wire AES_CORE_DATAPATH__abc_16259_n5330;
  wire AES_CORE_DATAPATH__abc_16259_n5331_1;
  wire AES_CORE_DATAPATH__abc_16259_n5332;
  wire AES_CORE_DATAPATH__abc_16259_n5333;
  wire AES_CORE_DATAPATH__abc_16259_n5334_1;
  wire AES_CORE_DATAPATH__abc_16259_n5335;
  wire AES_CORE_DATAPATH__abc_16259_n5336;
  wire AES_CORE_DATAPATH__abc_16259_n5337_1;
  wire AES_CORE_DATAPATH__abc_16259_n5339;
  wire AES_CORE_DATAPATH__abc_16259_n5340_1;
  wire AES_CORE_DATAPATH__abc_16259_n5341;
  wire AES_CORE_DATAPATH__abc_16259_n5342;
  wire AES_CORE_DATAPATH__abc_16259_n5343_1;
  wire AES_CORE_DATAPATH__abc_16259_n5344;
  wire AES_CORE_DATAPATH__abc_16259_n5345;
  wire AES_CORE_DATAPATH__abc_16259_n5346_1;
  wire AES_CORE_DATAPATH__abc_16259_n5348;
  wire AES_CORE_DATAPATH__abc_16259_n5349_1;
  wire AES_CORE_DATAPATH__abc_16259_n5350;
  wire AES_CORE_DATAPATH__abc_16259_n5351;
  wire AES_CORE_DATAPATH__abc_16259_n5352_1;
  wire AES_CORE_DATAPATH__abc_16259_n5353;
  wire AES_CORE_DATAPATH__abc_16259_n5354;
  wire AES_CORE_DATAPATH__abc_16259_n5355_1;
  wire AES_CORE_DATAPATH__abc_16259_n5357;
  wire AES_CORE_DATAPATH__abc_16259_n5358_1;
  wire AES_CORE_DATAPATH__abc_16259_n5359;
  wire AES_CORE_DATAPATH__abc_16259_n5360;
  wire AES_CORE_DATAPATH__abc_16259_n5361_1;
  wire AES_CORE_DATAPATH__abc_16259_n5362;
  wire AES_CORE_DATAPATH__abc_16259_n5363;
  wire AES_CORE_DATAPATH__abc_16259_n5364_1;
  wire AES_CORE_DATAPATH__abc_16259_n5366;
  wire AES_CORE_DATAPATH__abc_16259_n5367_1;
  wire AES_CORE_DATAPATH__abc_16259_n5368_1;
  wire AES_CORE_DATAPATH__abc_16259_n5369_1;
  wire AES_CORE_DATAPATH__abc_16259_n5370_1;
  wire AES_CORE_DATAPATH__abc_16259_n5371_1;
  wire AES_CORE_DATAPATH__abc_16259_n5372_1;
  wire AES_CORE_DATAPATH__abc_16259_n5373_1;
  wire AES_CORE_DATAPATH__abc_16259_n5375_1;
  wire AES_CORE_DATAPATH__abc_16259_n5376_1;
  wire AES_CORE_DATAPATH__abc_16259_n5377_1;
  wire AES_CORE_DATAPATH__abc_16259_n5378_1;
  wire AES_CORE_DATAPATH__abc_16259_n5379_1;
  wire AES_CORE_DATAPATH__abc_16259_n5380_1;
  wire AES_CORE_DATAPATH__abc_16259_n5381_1;
  wire AES_CORE_DATAPATH__abc_16259_n5382_1;
  wire AES_CORE_DATAPATH__abc_16259_n5384_1;
  wire AES_CORE_DATAPATH__abc_16259_n5385_1;
  wire AES_CORE_DATAPATH__abc_16259_n5386_1;
  wire AES_CORE_DATAPATH__abc_16259_n5387_1;
  wire AES_CORE_DATAPATH__abc_16259_n5388_1;
  wire AES_CORE_DATAPATH__abc_16259_n5389_1;
  wire AES_CORE_DATAPATH__abc_16259_n5390_1;
  wire AES_CORE_DATAPATH__abc_16259_n5391_1;
  wire AES_CORE_DATAPATH__abc_16259_n5393_1;
  wire AES_CORE_DATAPATH__abc_16259_n5394_1;
  wire AES_CORE_DATAPATH__abc_16259_n5395_1;
  wire AES_CORE_DATAPATH__abc_16259_n5396_1;
  wire AES_CORE_DATAPATH__abc_16259_n5397_1;
  wire AES_CORE_DATAPATH__abc_16259_n5398_1;
  wire AES_CORE_DATAPATH__abc_16259_n5399_1;
  wire AES_CORE_DATAPATH__abc_16259_n5400_1;
  wire AES_CORE_DATAPATH__abc_16259_n5402_1;
  wire AES_CORE_DATAPATH__abc_16259_n5403_1;
  wire AES_CORE_DATAPATH__abc_16259_n5404_1;
  wire AES_CORE_DATAPATH__abc_16259_n5405_1;
  wire AES_CORE_DATAPATH__abc_16259_n5406_1;
  wire AES_CORE_DATAPATH__abc_16259_n5407_1;
  wire AES_CORE_DATAPATH__abc_16259_n5408_1;
  wire AES_CORE_DATAPATH__abc_16259_n5409_1;
  wire AES_CORE_DATAPATH__abc_16259_n5411_1;
  wire AES_CORE_DATAPATH__abc_16259_n5412_1;
  wire AES_CORE_DATAPATH__abc_16259_n5413_1;
  wire AES_CORE_DATAPATH__abc_16259_n5414_1;
  wire AES_CORE_DATAPATH__abc_16259_n5415_1;
  wire AES_CORE_DATAPATH__abc_16259_n5416_1;
  wire AES_CORE_DATAPATH__abc_16259_n5417_1;
  wire AES_CORE_DATAPATH__abc_16259_n5418_1;
  wire AES_CORE_DATAPATH__abc_16259_n5420_1;
  wire AES_CORE_DATAPATH__abc_16259_n5421_1;
  wire AES_CORE_DATAPATH__abc_16259_n5422_1;
  wire AES_CORE_DATAPATH__abc_16259_n5423_1;
  wire AES_CORE_DATAPATH__abc_16259_n5424_1;
  wire AES_CORE_DATAPATH__abc_16259_n5425_1;
  wire AES_CORE_DATAPATH__abc_16259_n5426_1;
  wire AES_CORE_DATAPATH__abc_16259_n5427_1;
  wire AES_CORE_DATAPATH__abc_16259_n5429_1;
  wire AES_CORE_DATAPATH__abc_16259_n5430_1;
  wire AES_CORE_DATAPATH__abc_16259_n5431_1;
  wire AES_CORE_DATAPATH__abc_16259_n5432_1;
  wire AES_CORE_DATAPATH__abc_16259_n5433_1;
  wire AES_CORE_DATAPATH__abc_16259_n5434_1;
  wire AES_CORE_DATAPATH__abc_16259_n5435_1;
  wire AES_CORE_DATAPATH__abc_16259_n5436_1;
  wire AES_CORE_DATAPATH__abc_16259_n5438_1;
  wire AES_CORE_DATAPATH__abc_16259_n5439_1;
  wire AES_CORE_DATAPATH__abc_16259_n5440_1;
  wire AES_CORE_DATAPATH__abc_16259_n5441_1;
  wire AES_CORE_DATAPATH__abc_16259_n5442_1;
  wire AES_CORE_DATAPATH__abc_16259_n5443_1;
  wire AES_CORE_DATAPATH__abc_16259_n5444_1;
  wire AES_CORE_DATAPATH__abc_16259_n5445_1;
  wire AES_CORE_DATAPATH__abc_16259_n5447_1;
  wire AES_CORE_DATAPATH__abc_16259_n5448_1;
  wire AES_CORE_DATAPATH__abc_16259_n5449_1;
  wire AES_CORE_DATAPATH__abc_16259_n5450_1;
  wire AES_CORE_DATAPATH__abc_16259_n5451_1;
  wire AES_CORE_DATAPATH__abc_16259_n5452;
  wire AES_CORE_DATAPATH__abc_16259_n5453;
  wire AES_CORE_DATAPATH__abc_16259_n5454;
  wire AES_CORE_DATAPATH__abc_16259_n5456;
  wire AES_CORE_DATAPATH__abc_16259_n5457;
  wire AES_CORE_DATAPATH__abc_16259_n5458;
  wire AES_CORE_DATAPATH__abc_16259_n5459;
  wire AES_CORE_DATAPATH__abc_16259_n5460;
  wire AES_CORE_DATAPATH__abc_16259_n5461;
  wire AES_CORE_DATAPATH__abc_16259_n5462;
  wire AES_CORE_DATAPATH__abc_16259_n5463;
  wire AES_CORE_DATAPATH__abc_16259_n5465;
  wire AES_CORE_DATAPATH__abc_16259_n5466;
  wire AES_CORE_DATAPATH__abc_16259_n5467;
  wire AES_CORE_DATAPATH__abc_16259_n5468;
  wire AES_CORE_DATAPATH__abc_16259_n5469;
  wire AES_CORE_DATAPATH__abc_16259_n5470;
  wire AES_CORE_DATAPATH__abc_16259_n5471;
  wire AES_CORE_DATAPATH__abc_16259_n5472;
  wire AES_CORE_DATAPATH__abc_16259_n5474;
  wire AES_CORE_DATAPATH__abc_16259_n5475;
  wire AES_CORE_DATAPATH__abc_16259_n5476;
  wire AES_CORE_DATAPATH__abc_16259_n5477;
  wire AES_CORE_DATAPATH__abc_16259_n5478;
  wire AES_CORE_DATAPATH__abc_16259_n5479;
  wire AES_CORE_DATAPATH__abc_16259_n5480;
  wire AES_CORE_DATAPATH__abc_16259_n5481;
  wire AES_CORE_DATAPATH__abc_16259_n5483;
  wire AES_CORE_DATAPATH__abc_16259_n5484;
  wire AES_CORE_DATAPATH__abc_16259_n5485;
  wire AES_CORE_DATAPATH__abc_16259_n5486;
  wire AES_CORE_DATAPATH__abc_16259_n5487;
  wire AES_CORE_DATAPATH__abc_16259_n5488;
  wire AES_CORE_DATAPATH__abc_16259_n5489;
  wire AES_CORE_DATAPATH__abc_16259_n5490;
  wire AES_CORE_DATAPATH__abc_16259_n5492;
  wire AES_CORE_DATAPATH__abc_16259_n5493;
  wire AES_CORE_DATAPATH__abc_16259_n5494;
  wire AES_CORE_DATAPATH__abc_16259_n5495;
  wire AES_CORE_DATAPATH__abc_16259_n5496;
  wire AES_CORE_DATAPATH__abc_16259_n5497;
  wire AES_CORE_DATAPATH__abc_16259_n5498;
  wire AES_CORE_DATAPATH__abc_16259_n5499;
  wire AES_CORE_DATAPATH__abc_16259_n5501;
  wire AES_CORE_DATAPATH__abc_16259_n5502;
  wire AES_CORE_DATAPATH__abc_16259_n5503;
  wire AES_CORE_DATAPATH__abc_16259_n5504;
  wire AES_CORE_DATAPATH__abc_16259_n5505;
  wire AES_CORE_DATAPATH__abc_16259_n5506;
  wire AES_CORE_DATAPATH__abc_16259_n5507;
  wire AES_CORE_DATAPATH__abc_16259_n5508;
  wire AES_CORE_DATAPATH__abc_16259_n5510;
  wire AES_CORE_DATAPATH__abc_16259_n5511;
  wire AES_CORE_DATAPATH__abc_16259_n5512;
  wire AES_CORE_DATAPATH__abc_16259_n5513;
  wire AES_CORE_DATAPATH__abc_16259_n5514;
  wire AES_CORE_DATAPATH__abc_16259_n5515;
  wire AES_CORE_DATAPATH__abc_16259_n5516;
  wire AES_CORE_DATAPATH__abc_16259_n5517;
  wire AES_CORE_DATAPATH__abc_16259_n5519;
  wire AES_CORE_DATAPATH__abc_16259_n5520;
  wire AES_CORE_DATAPATH__abc_16259_n5521;
  wire AES_CORE_DATAPATH__abc_16259_n5522;
  wire AES_CORE_DATAPATH__abc_16259_n5523;
  wire AES_CORE_DATAPATH__abc_16259_n5524;
  wire AES_CORE_DATAPATH__abc_16259_n5525;
  wire AES_CORE_DATAPATH__abc_16259_n5526;
  wire AES_CORE_DATAPATH__abc_16259_n5528;
  wire AES_CORE_DATAPATH__abc_16259_n5529;
  wire AES_CORE_DATAPATH__abc_16259_n5530;
  wire AES_CORE_DATAPATH__abc_16259_n5531;
  wire AES_CORE_DATAPATH__abc_16259_n5532;
  wire AES_CORE_DATAPATH__abc_16259_n5533;
  wire AES_CORE_DATAPATH__abc_16259_n5534;
  wire AES_CORE_DATAPATH__abc_16259_n5535;
  wire AES_CORE_DATAPATH__abc_16259_n5537;
  wire AES_CORE_DATAPATH__abc_16259_n5538;
  wire AES_CORE_DATAPATH__abc_16259_n5539;
  wire AES_CORE_DATAPATH__abc_16259_n5540;
  wire AES_CORE_DATAPATH__abc_16259_n5541;
  wire AES_CORE_DATAPATH__abc_16259_n5542;
  wire AES_CORE_DATAPATH__abc_16259_n5543;
  wire AES_CORE_DATAPATH__abc_16259_n5544;
  wire AES_CORE_DATAPATH__abc_16259_n5546;
  wire AES_CORE_DATAPATH__abc_16259_n5547;
  wire AES_CORE_DATAPATH__abc_16259_n5548;
  wire AES_CORE_DATAPATH__abc_16259_n5549;
  wire AES_CORE_DATAPATH__abc_16259_n5550;
  wire AES_CORE_DATAPATH__abc_16259_n5551;
  wire AES_CORE_DATAPATH__abc_16259_n5552;
  wire AES_CORE_DATAPATH__abc_16259_n5553;
  wire AES_CORE_DATAPATH__abc_16259_n5555;
  wire AES_CORE_DATAPATH__abc_16259_n5556;
  wire AES_CORE_DATAPATH__abc_16259_n5558;
  wire AES_CORE_DATAPATH__abc_16259_n5559;
  wire AES_CORE_DATAPATH__abc_16259_n5561;
  wire AES_CORE_DATAPATH__abc_16259_n5562;
  wire AES_CORE_DATAPATH__abc_16259_n5564;
  wire AES_CORE_DATAPATH__abc_16259_n5565;
  wire AES_CORE_DATAPATH__abc_16259_n5567;
  wire AES_CORE_DATAPATH__abc_16259_n5568;
  wire AES_CORE_DATAPATH__abc_16259_n5570;
  wire AES_CORE_DATAPATH__abc_16259_n5571;
  wire AES_CORE_DATAPATH__abc_16259_n5573;
  wire AES_CORE_DATAPATH__abc_16259_n5574;
  wire AES_CORE_DATAPATH__abc_16259_n5576;
  wire AES_CORE_DATAPATH__abc_16259_n5577;
  wire AES_CORE_DATAPATH__abc_16259_n5579;
  wire AES_CORE_DATAPATH__abc_16259_n5580;
  wire AES_CORE_DATAPATH__abc_16259_n5582;
  wire AES_CORE_DATAPATH__abc_16259_n5583;
  wire AES_CORE_DATAPATH__abc_16259_n5585;
  wire AES_CORE_DATAPATH__abc_16259_n5586;
  wire AES_CORE_DATAPATH__abc_16259_n5588;
  wire AES_CORE_DATAPATH__abc_16259_n5589;
  wire AES_CORE_DATAPATH__abc_16259_n5591;
  wire AES_CORE_DATAPATH__abc_16259_n5592;
  wire AES_CORE_DATAPATH__abc_16259_n5594;
  wire AES_CORE_DATAPATH__abc_16259_n5595;
  wire AES_CORE_DATAPATH__abc_16259_n5597;
  wire AES_CORE_DATAPATH__abc_16259_n5598;
  wire AES_CORE_DATAPATH__abc_16259_n5600;
  wire AES_CORE_DATAPATH__abc_16259_n5601;
  wire AES_CORE_DATAPATH__abc_16259_n5603;
  wire AES_CORE_DATAPATH__abc_16259_n5604;
  wire AES_CORE_DATAPATH__abc_16259_n5606;
  wire AES_CORE_DATAPATH__abc_16259_n5607;
  wire AES_CORE_DATAPATH__abc_16259_n5609;
  wire AES_CORE_DATAPATH__abc_16259_n5610;
  wire AES_CORE_DATAPATH__abc_16259_n5612;
  wire AES_CORE_DATAPATH__abc_16259_n5613;
  wire AES_CORE_DATAPATH__abc_16259_n5615;
  wire AES_CORE_DATAPATH__abc_16259_n5616;
  wire AES_CORE_DATAPATH__abc_16259_n5618;
  wire AES_CORE_DATAPATH__abc_16259_n5619;
  wire AES_CORE_DATAPATH__abc_16259_n5621;
  wire AES_CORE_DATAPATH__abc_16259_n5622;
  wire AES_CORE_DATAPATH__abc_16259_n5624;
  wire AES_CORE_DATAPATH__abc_16259_n5625;
  wire AES_CORE_DATAPATH__abc_16259_n5627;
  wire AES_CORE_DATAPATH__abc_16259_n5628;
  wire AES_CORE_DATAPATH__abc_16259_n5630;
  wire AES_CORE_DATAPATH__abc_16259_n5631;
  wire AES_CORE_DATAPATH__abc_16259_n5633;
  wire AES_CORE_DATAPATH__abc_16259_n5634;
  wire AES_CORE_DATAPATH__abc_16259_n5636;
  wire AES_CORE_DATAPATH__abc_16259_n5637;
  wire AES_CORE_DATAPATH__abc_16259_n5639;
  wire AES_CORE_DATAPATH__abc_16259_n5640;
  wire AES_CORE_DATAPATH__abc_16259_n5642;
  wire AES_CORE_DATAPATH__abc_16259_n5643;
  wire AES_CORE_DATAPATH__abc_16259_n5645;
  wire AES_CORE_DATAPATH__abc_16259_n5646;
  wire AES_CORE_DATAPATH__abc_16259_n5648;
  wire AES_CORE_DATAPATH__abc_16259_n5649;
  wire AES_CORE_DATAPATH__abc_16259_n5651;
  wire AES_CORE_DATAPATH__abc_16259_n5652;
  wire AES_CORE_DATAPATH__abc_16259_n5653;
  wire AES_CORE_DATAPATH__abc_16259_n5653_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n5653_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n5653_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n5653_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n5653_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n5654;
  wire AES_CORE_DATAPATH__abc_16259_n5655;
  wire AES_CORE_DATAPATH__abc_16259_n5656;
  wire AES_CORE_DATAPATH__abc_16259_n5657;
  wire AES_CORE_DATAPATH__abc_16259_n5658;
  wire AES_CORE_DATAPATH__abc_16259_n5658_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n5658_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n5658_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n5658_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n5658_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n5659;
  wire AES_CORE_DATAPATH__abc_16259_n5659_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n5659_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n5659_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n5659_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n5659_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n5660;
  wire AES_CORE_DATAPATH__abc_16259_n5661;
  wire AES_CORE_DATAPATH__abc_16259_n5662;
  wire AES_CORE_DATAPATH__abc_16259_n5663;
  wire AES_CORE_DATAPATH__abc_16259_n5664;
  wire AES_CORE_DATAPATH__abc_16259_n5665;
  wire AES_CORE_DATAPATH__abc_16259_n5666;
  wire AES_CORE_DATAPATH__abc_16259_n5667;
  wire AES_CORE_DATAPATH__abc_16259_n5669;
  wire AES_CORE_DATAPATH__abc_16259_n5670;
  wire AES_CORE_DATAPATH__abc_16259_n5671;
  wire AES_CORE_DATAPATH__abc_16259_n5672;
  wire AES_CORE_DATAPATH__abc_16259_n5673;
  wire AES_CORE_DATAPATH__abc_16259_n5674;
  wire AES_CORE_DATAPATH__abc_16259_n5675;
  wire AES_CORE_DATAPATH__abc_16259_n5676;
  wire AES_CORE_DATAPATH__abc_16259_n5678;
  wire AES_CORE_DATAPATH__abc_16259_n5679;
  wire AES_CORE_DATAPATH__abc_16259_n5680;
  wire AES_CORE_DATAPATH__abc_16259_n5681;
  wire AES_CORE_DATAPATH__abc_16259_n5682;
  wire AES_CORE_DATAPATH__abc_16259_n5683;
  wire AES_CORE_DATAPATH__abc_16259_n5684;
  wire AES_CORE_DATAPATH__abc_16259_n5685;
  wire AES_CORE_DATAPATH__abc_16259_n5687;
  wire AES_CORE_DATAPATH__abc_16259_n5688;
  wire AES_CORE_DATAPATH__abc_16259_n5689;
  wire AES_CORE_DATAPATH__abc_16259_n5690;
  wire AES_CORE_DATAPATH__abc_16259_n5691;
  wire AES_CORE_DATAPATH__abc_16259_n5692;
  wire AES_CORE_DATAPATH__abc_16259_n5693;
  wire AES_CORE_DATAPATH__abc_16259_n5694;
  wire AES_CORE_DATAPATH__abc_16259_n5696;
  wire AES_CORE_DATAPATH__abc_16259_n5697;
  wire AES_CORE_DATAPATH__abc_16259_n5698;
  wire AES_CORE_DATAPATH__abc_16259_n5699;
  wire AES_CORE_DATAPATH__abc_16259_n5700;
  wire AES_CORE_DATAPATH__abc_16259_n5701;
  wire AES_CORE_DATAPATH__abc_16259_n5702;
  wire AES_CORE_DATAPATH__abc_16259_n5703;
  wire AES_CORE_DATAPATH__abc_16259_n5705;
  wire AES_CORE_DATAPATH__abc_16259_n5706;
  wire AES_CORE_DATAPATH__abc_16259_n5707;
  wire AES_CORE_DATAPATH__abc_16259_n5708;
  wire AES_CORE_DATAPATH__abc_16259_n5709;
  wire AES_CORE_DATAPATH__abc_16259_n5710;
  wire AES_CORE_DATAPATH__abc_16259_n5711;
  wire AES_CORE_DATAPATH__abc_16259_n5712;
  wire AES_CORE_DATAPATH__abc_16259_n5714;
  wire AES_CORE_DATAPATH__abc_16259_n5715;
  wire AES_CORE_DATAPATH__abc_16259_n5716;
  wire AES_CORE_DATAPATH__abc_16259_n5717;
  wire AES_CORE_DATAPATH__abc_16259_n5718;
  wire AES_CORE_DATAPATH__abc_16259_n5719;
  wire AES_CORE_DATAPATH__abc_16259_n5720;
  wire AES_CORE_DATAPATH__abc_16259_n5721;
  wire AES_CORE_DATAPATH__abc_16259_n5723;
  wire AES_CORE_DATAPATH__abc_16259_n5724;
  wire AES_CORE_DATAPATH__abc_16259_n5725;
  wire AES_CORE_DATAPATH__abc_16259_n5726;
  wire AES_CORE_DATAPATH__abc_16259_n5727;
  wire AES_CORE_DATAPATH__abc_16259_n5728;
  wire AES_CORE_DATAPATH__abc_16259_n5729;
  wire AES_CORE_DATAPATH__abc_16259_n5730;
  wire AES_CORE_DATAPATH__abc_16259_n5732;
  wire AES_CORE_DATAPATH__abc_16259_n5733;
  wire AES_CORE_DATAPATH__abc_16259_n5734;
  wire AES_CORE_DATAPATH__abc_16259_n5735;
  wire AES_CORE_DATAPATH__abc_16259_n5736;
  wire AES_CORE_DATAPATH__abc_16259_n5737;
  wire AES_CORE_DATAPATH__abc_16259_n5738;
  wire AES_CORE_DATAPATH__abc_16259_n5739;
  wire AES_CORE_DATAPATH__abc_16259_n5741;
  wire AES_CORE_DATAPATH__abc_16259_n5742;
  wire AES_CORE_DATAPATH__abc_16259_n5743;
  wire AES_CORE_DATAPATH__abc_16259_n5744;
  wire AES_CORE_DATAPATH__abc_16259_n5745;
  wire AES_CORE_DATAPATH__abc_16259_n5746;
  wire AES_CORE_DATAPATH__abc_16259_n5747;
  wire AES_CORE_DATAPATH__abc_16259_n5748;
  wire AES_CORE_DATAPATH__abc_16259_n5750;
  wire AES_CORE_DATAPATH__abc_16259_n5751;
  wire AES_CORE_DATAPATH__abc_16259_n5752;
  wire AES_CORE_DATAPATH__abc_16259_n5753;
  wire AES_CORE_DATAPATH__abc_16259_n5754;
  wire AES_CORE_DATAPATH__abc_16259_n5755;
  wire AES_CORE_DATAPATH__abc_16259_n5756;
  wire AES_CORE_DATAPATH__abc_16259_n5757;
  wire AES_CORE_DATAPATH__abc_16259_n5759;
  wire AES_CORE_DATAPATH__abc_16259_n5760;
  wire AES_CORE_DATAPATH__abc_16259_n5761;
  wire AES_CORE_DATAPATH__abc_16259_n5762;
  wire AES_CORE_DATAPATH__abc_16259_n5763;
  wire AES_CORE_DATAPATH__abc_16259_n5764;
  wire AES_CORE_DATAPATH__abc_16259_n5765;
  wire AES_CORE_DATAPATH__abc_16259_n5766;
  wire AES_CORE_DATAPATH__abc_16259_n5768;
  wire AES_CORE_DATAPATH__abc_16259_n5769;
  wire AES_CORE_DATAPATH__abc_16259_n5770;
  wire AES_CORE_DATAPATH__abc_16259_n5771;
  wire AES_CORE_DATAPATH__abc_16259_n5772;
  wire AES_CORE_DATAPATH__abc_16259_n5773;
  wire AES_CORE_DATAPATH__abc_16259_n5774;
  wire AES_CORE_DATAPATH__abc_16259_n5775;
  wire AES_CORE_DATAPATH__abc_16259_n5777;
  wire AES_CORE_DATAPATH__abc_16259_n5778;
  wire AES_CORE_DATAPATH__abc_16259_n5779;
  wire AES_CORE_DATAPATH__abc_16259_n5780;
  wire AES_CORE_DATAPATH__abc_16259_n5781;
  wire AES_CORE_DATAPATH__abc_16259_n5782;
  wire AES_CORE_DATAPATH__abc_16259_n5783;
  wire AES_CORE_DATAPATH__abc_16259_n5784;
  wire AES_CORE_DATAPATH__abc_16259_n5786;
  wire AES_CORE_DATAPATH__abc_16259_n5787;
  wire AES_CORE_DATAPATH__abc_16259_n5788;
  wire AES_CORE_DATAPATH__abc_16259_n5789;
  wire AES_CORE_DATAPATH__abc_16259_n5790;
  wire AES_CORE_DATAPATH__abc_16259_n5791;
  wire AES_CORE_DATAPATH__abc_16259_n5792;
  wire AES_CORE_DATAPATH__abc_16259_n5793;
  wire AES_CORE_DATAPATH__abc_16259_n5795;
  wire AES_CORE_DATAPATH__abc_16259_n5796;
  wire AES_CORE_DATAPATH__abc_16259_n5797;
  wire AES_CORE_DATAPATH__abc_16259_n5798;
  wire AES_CORE_DATAPATH__abc_16259_n5799;
  wire AES_CORE_DATAPATH__abc_16259_n5800;
  wire AES_CORE_DATAPATH__abc_16259_n5801;
  wire AES_CORE_DATAPATH__abc_16259_n5802;
  wire AES_CORE_DATAPATH__abc_16259_n5804;
  wire AES_CORE_DATAPATH__abc_16259_n5805;
  wire AES_CORE_DATAPATH__abc_16259_n5806;
  wire AES_CORE_DATAPATH__abc_16259_n5807;
  wire AES_CORE_DATAPATH__abc_16259_n5808;
  wire AES_CORE_DATAPATH__abc_16259_n5809;
  wire AES_CORE_DATAPATH__abc_16259_n5810;
  wire AES_CORE_DATAPATH__abc_16259_n5811;
  wire AES_CORE_DATAPATH__abc_16259_n5813;
  wire AES_CORE_DATAPATH__abc_16259_n5814;
  wire AES_CORE_DATAPATH__abc_16259_n5815;
  wire AES_CORE_DATAPATH__abc_16259_n5816;
  wire AES_CORE_DATAPATH__abc_16259_n5817;
  wire AES_CORE_DATAPATH__abc_16259_n5818;
  wire AES_CORE_DATAPATH__abc_16259_n5819;
  wire AES_CORE_DATAPATH__abc_16259_n5820;
  wire AES_CORE_DATAPATH__abc_16259_n5822;
  wire AES_CORE_DATAPATH__abc_16259_n5823;
  wire AES_CORE_DATAPATH__abc_16259_n5824;
  wire AES_CORE_DATAPATH__abc_16259_n5825;
  wire AES_CORE_DATAPATH__abc_16259_n5826;
  wire AES_CORE_DATAPATH__abc_16259_n5827;
  wire AES_CORE_DATAPATH__abc_16259_n5828;
  wire AES_CORE_DATAPATH__abc_16259_n5829;
  wire AES_CORE_DATAPATH__abc_16259_n5831;
  wire AES_CORE_DATAPATH__abc_16259_n5832;
  wire AES_CORE_DATAPATH__abc_16259_n5833;
  wire AES_CORE_DATAPATH__abc_16259_n5834;
  wire AES_CORE_DATAPATH__abc_16259_n5835;
  wire AES_CORE_DATAPATH__abc_16259_n5836;
  wire AES_CORE_DATAPATH__abc_16259_n5837;
  wire AES_CORE_DATAPATH__abc_16259_n5838;
  wire AES_CORE_DATAPATH__abc_16259_n5840;
  wire AES_CORE_DATAPATH__abc_16259_n5841;
  wire AES_CORE_DATAPATH__abc_16259_n5842;
  wire AES_CORE_DATAPATH__abc_16259_n5843;
  wire AES_CORE_DATAPATH__abc_16259_n5844;
  wire AES_CORE_DATAPATH__abc_16259_n5845;
  wire AES_CORE_DATAPATH__abc_16259_n5846;
  wire AES_CORE_DATAPATH__abc_16259_n5847;
  wire AES_CORE_DATAPATH__abc_16259_n5849;
  wire AES_CORE_DATAPATH__abc_16259_n5850;
  wire AES_CORE_DATAPATH__abc_16259_n5851;
  wire AES_CORE_DATAPATH__abc_16259_n5852;
  wire AES_CORE_DATAPATH__abc_16259_n5853;
  wire AES_CORE_DATAPATH__abc_16259_n5854;
  wire AES_CORE_DATAPATH__abc_16259_n5855;
  wire AES_CORE_DATAPATH__abc_16259_n5856;
  wire AES_CORE_DATAPATH__abc_16259_n5858;
  wire AES_CORE_DATAPATH__abc_16259_n5859;
  wire AES_CORE_DATAPATH__abc_16259_n5860;
  wire AES_CORE_DATAPATH__abc_16259_n5861;
  wire AES_CORE_DATAPATH__abc_16259_n5862;
  wire AES_CORE_DATAPATH__abc_16259_n5863;
  wire AES_CORE_DATAPATH__abc_16259_n5864;
  wire AES_CORE_DATAPATH__abc_16259_n5865;
  wire AES_CORE_DATAPATH__abc_16259_n5867;
  wire AES_CORE_DATAPATH__abc_16259_n5868;
  wire AES_CORE_DATAPATH__abc_16259_n5869;
  wire AES_CORE_DATAPATH__abc_16259_n5870;
  wire AES_CORE_DATAPATH__abc_16259_n5871;
  wire AES_CORE_DATAPATH__abc_16259_n5872;
  wire AES_CORE_DATAPATH__abc_16259_n5873;
  wire AES_CORE_DATAPATH__abc_16259_n5874;
  wire AES_CORE_DATAPATH__abc_16259_n5876;
  wire AES_CORE_DATAPATH__abc_16259_n5877;
  wire AES_CORE_DATAPATH__abc_16259_n5878;
  wire AES_CORE_DATAPATH__abc_16259_n5879;
  wire AES_CORE_DATAPATH__abc_16259_n5880;
  wire AES_CORE_DATAPATH__abc_16259_n5881;
  wire AES_CORE_DATAPATH__abc_16259_n5882;
  wire AES_CORE_DATAPATH__abc_16259_n5883;
  wire AES_CORE_DATAPATH__abc_16259_n5885;
  wire AES_CORE_DATAPATH__abc_16259_n5886;
  wire AES_CORE_DATAPATH__abc_16259_n5887;
  wire AES_CORE_DATAPATH__abc_16259_n5888;
  wire AES_CORE_DATAPATH__abc_16259_n5889;
  wire AES_CORE_DATAPATH__abc_16259_n5890;
  wire AES_CORE_DATAPATH__abc_16259_n5891;
  wire AES_CORE_DATAPATH__abc_16259_n5892;
  wire AES_CORE_DATAPATH__abc_16259_n5894;
  wire AES_CORE_DATAPATH__abc_16259_n5895;
  wire AES_CORE_DATAPATH__abc_16259_n5896;
  wire AES_CORE_DATAPATH__abc_16259_n5897;
  wire AES_CORE_DATAPATH__abc_16259_n5898;
  wire AES_CORE_DATAPATH__abc_16259_n5899;
  wire AES_CORE_DATAPATH__abc_16259_n5900;
  wire AES_CORE_DATAPATH__abc_16259_n5901;
  wire AES_CORE_DATAPATH__abc_16259_n5903;
  wire AES_CORE_DATAPATH__abc_16259_n5904;
  wire AES_CORE_DATAPATH__abc_16259_n5905;
  wire AES_CORE_DATAPATH__abc_16259_n5906;
  wire AES_CORE_DATAPATH__abc_16259_n5907;
  wire AES_CORE_DATAPATH__abc_16259_n5908;
  wire AES_CORE_DATAPATH__abc_16259_n5909;
  wire AES_CORE_DATAPATH__abc_16259_n5910;
  wire AES_CORE_DATAPATH__abc_16259_n5912;
  wire AES_CORE_DATAPATH__abc_16259_n5913;
  wire AES_CORE_DATAPATH__abc_16259_n5914;
  wire AES_CORE_DATAPATH__abc_16259_n5915;
  wire AES_CORE_DATAPATH__abc_16259_n5916;
  wire AES_CORE_DATAPATH__abc_16259_n5917;
  wire AES_CORE_DATAPATH__abc_16259_n5918;
  wire AES_CORE_DATAPATH__abc_16259_n5919;
  wire AES_CORE_DATAPATH__abc_16259_n5921;
  wire AES_CORE_DATAPATH__abc_16259_n5922;
  wire AES_CORE_DATAPATH__abc_16259_n5923;
  wire AES_CORE_DATAPATH__abc_16259_n5924;
  wire AES_CORE_DATAPATH__abc_16259_n5925;
  wire AES_CORE_DATAPATH__abc_16259_n5926;
  wire AES_CORE_DATAPATH__abc_16259_n5927;
  wire AES_CORE_DATAPATH__abc_16259_n5928;
  wire AES_CORE_DATAPATH__abc_16259_n5930;
  wire AES_CORE_DATAPATH__abc_16259_n5931;
  wire AES_CORE_DATAPATH__abc_16259_n5932;
  wire AES_CORE_DATAPATH__abc_16259_n5933;
  wire AES_CORE_DATAPATH__abc_16259_n5934;
  wire AES_CORE_DATAPATH__abc_16259_n5935;
  wire AES_CORE_DATAPATH__abc_16259_n5936;
  wire AES_CORE_DATAPATH__abc_16259_n5937;
  wire AES_CORE_DATAPATH__abc_16259_n5939;
  wire AES_CORE_DATAPATH__abc_16259_n5940;
  wire AES_CORE_DATAPATH__abc_16259_n5941;
  wire AES_CORE_DATAPATH__abc_16259_n5942;
  wire AES_CORE_DATAPATH__abc_16259_n5943;
  wire AES_CORE_DATAPATH__abc_16259_n5944;
  wire AES_CORE_DATAPATH__abc_16259_n5945;
  wire AES_CORE_DATAPATH__abc_16259_n5946;
  wire AES_CORE_DATAPATH__abc_16259_n5948;
  wire AES_CORE_DATAPATH__abc_16259_n5949;
  wire AES_CORE_DATAPATH__abc_16259_n5951;
  wire AES_CORE_DATAPATH__abc_16259_n5952;
  wire AES_CORE_DATAPATH__abc_16259_n5954;
  wire AES_CORE_DATAPATH__abc_16259_n5955;
  wire AES_CORE_DATAPATH__abc_16259_n5957;
  wire AES_CORE_DATAPATH__abc_16259_n5958;
  wire AES_CORE_DATAPATH__abc_16259_n5960;
  wire AES_CORE_DATAPATH__abc_16259_n5961;
  wire AES_CORE_DATAPATH__abc_16259_n5963;
  wire AES_CORE_DATAPATH__abc_16259_n5964;
  wire AES_CORE_DATAPATH__abc_16259_n5966;
  wire AES_CORE_DATAPATH__abc_16259_n5967;
  wire AES_CORE_DATAPATH__abc_16259_n5969;
  wire AES_CORE_DATAPATH__abc_16259_n5970;
  wire AES_CORE_DATAPATH__abc_16259_n5972;
  wire AES_CORE_DATAPATH__abc_16259_n5973;
  wire AES_CORE_DATAPATH__abc_16259_n5975;
  wire AES_CORE_DATAPATH__abc_16259_n5976;
  wire AES_CORE_DATAPATH__abc_16259_n5978;
  wire AES_CORE_DATAPATH__abc_16259_n5979;
  wire AES_CORE_DATAPATH__abc_16259_n5981;
  wire AES_CORE_DATAPATH__abc_16259_n5982;
  wire AES_CORE_DATAPATH__abc_16259_n5984;
  wire AES_CORE_DATAPATH__abc_16259_n5985;
  wire AES_CORE_DATAPATH__abc_16259_n5987;
  wire AES_CORE_DATAPATH__abc_16259_n5988;
  wire AES_CORE_DATAPATH__abc_16259_n5990;
  wire AES_CORE_DATAPATH__abc_16259_n5991;
  wire AES_CORE_DATAPATH__abc_16259_n5993;
  wire AES_CORE_DATAPATH__abc_16259_n5994;
  wire AES_CORE_DATAPATH__abc_16259_n5996;
  wire AES_CORE_DATAPATH__abc_16259_n5997;
  wire AES_CORE_DATAPATH__abc_16259_n5999;
  wire AES_CORE_DATAPATH__abc_16259_n6000;
  wire AES_CORE_DATAPATH__abc_16259_n6002;
  wire AES_CORE_DATAPATH__abc_16259_n6003;
  wire AES_CORE_DATAPATH__abc_16259_n6005;
  wire AES_CORE_DATAPATH__abc_16259_n6006;
  wire AES_CORE_DATAPATH__abc_16259_n6008;
  wire AES_CORE_DATAPATH__abc_16259_n6009;
  wire AES_CORE_DATAPATH__abc_16259_n6011;
  wire AES_CORE_DATAPATH__abc_16259_n6012;
  wire AES_CORE_DATAPATH__abc_16259_n6014;
  wire AES_CORE_DATAPATH__abc_16259_n6015;
  wire AES_CORE_DATAPATH__abc_16259_n6017;
  wire AES_CORE_DATAPATH__abc_16259_n6018;
  wire AES_CORE_DATAPATH__abc_16259_n6020;
  wire AES_CORE_DATAPATH__abc_16259_n6021;
  wire AES_CORE_DATAPATH__abc_16259_n6023;
  wire AES_CORE_DATAPATH__abc_16259_n6024;
  wire AES_CORE_DATAPATH__abc_16259_n6026;
  wire AES_CORE_DATAPATH__abc_16259_n6027;
  wire AES_CORE_DATAPATH__abc_16259_n6029;
  wire AES_CORE_DATAPATH__abc_16259_n6030;
  wire AES_CORE_DATAPATH__abc_16259_n6032;
  wire AES_CORE_DATAPATH__abc_16259_n6033;
  wire AES_CORE_DATAPATH__abc_16259_n6035;
  wire AES_CORE_DATAPATH__abc_16259_n6036;
  wire AES_CORE_DATAPATH__abc_16259_n6038;
  wire AES_CORE_DATAPATH__abc_16259_n6039;
  wire AES_CORE_DATAPATH__abc_16259_n6041;
  wire AES_CORE_DATAPATH__abc_16259_n6042;
  wire AES_CORE_DATAPATH__abc_16259_n6044;
  wire AES_CORE_DATAPATH__abc_16259_n6044_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n6044_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n6044_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n6044_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n6044_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n6045;
  wire AES_CORE_DATAPATH__abc_16259_n6046;
  wire AES_CORE_DATAPATH__abc_16259_n6047;
  wire AES_CORE_DATAPATH__abc_16259_n6048;
  wire AES_CORE_DATAPATH__abc_16259_n6049;
  wire AES_CORE_DATAPATH__abc_16259_n6050;
  wire AES_CORE_DATAPATH__abc_16259_n6051;
  wire AES_CORE_DATAPATH__abc_16259_n6052;
  wire AES_CORE_DATAPATH__abc_16259_n6053;
  wire AES_CORE_DATAPATH__abc_16259_n6053_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n6053_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n6053_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n6053_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n6053_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n6054;
  wire AES_CORE_DATAPATH__abc_16259_n6055;
  wire AES_CORE_DATAPATH__abc_16259_n6056;
  wire AES_CORE_DATAPATH__abc_16259_n6056_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n6056_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n6056_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n6056_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n6056_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n6057;
  wire AES_CORE_DATAPATH__abc_16259_n6057_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n6057_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n6057_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n6057_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n6057_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n6058;
  wire AES_CORE_DATAPATH__abc_16259_n6058_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n6058_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n6058_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n6058_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n6058_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n6058_bF_buf5;
  wire AES_CORE_DATAPATH__abc_16259_n6058_bF_buf6;
  wire AES_CORE_DATAPATH__abc_16259_n6059;
  wire AES_CORE_DATAPATH__abc_16259_n6059_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n6059_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n6059_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n6059_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n6059_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n6059_bF_buf5;
  wire AES_CORE_DATAPATH__abc_16259_n6060;
  wire AES_CORE_DATAPATH__abc_16259_n6061;
  wire AES_CORE_DATAPATH__abc_16259_n6062;
  wire AES_CORE_DATAPATH__abc_16259_n6063;
  wire AES_CORE_DATAPATH__abc_16259_n6063_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n6063_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n6063_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n6063_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n6063_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n6064;
  wire AES_CORE_DATAPATH__abc_16259_n6065;
  wire AES_CORE_DATAPATH__abc_16259_n6066;
  wire AES_CORE_DATAPATH__abc_16259_n6067;
  wire AES_CORE_DATAPATH__abc_16259_n6068;
  wire AES_CORE_DATAPATH__abc_16259_n6069;
  wire AES_CORE_DATAPATH__abc_16259_n6070;
  wire AES_CORE_DATAPATH__abc_16259_n6071;
  wire AES_CORE_DATAPATH__abc_16259_n6072;
  wire AES_CORE_DATAPATH__abc_16259_n6073;
  wire AES_CORE_DATAPATH__abc_16259_n6074;
  wire AES_CORE_DATAPATH__abc_16259_n6074_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n6074_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n6074_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n6074_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n6074_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n6075;
  wire AES_CORE_DATAPATH__abc_16259_n6076;
  wire AES_CORE_DATAPATH__abc_16259_n6077;
  wire AES_CORE_DATAPATH__abc_16259_n6078;
  wire AES_CORE_DATAPATH__abc_16259_n6079;
  wire AES_CORE_DATAPATH__abc_16259_n6080;
  wire AES_CORE_DATAPATH__abc_16259_n6081;
  wire AES_CORE_DATAPATH__abc_16259_n6082;
  wire AES_CORE_DATAPATH__abc_16259_n6083;
  wire AES_CORE_DATAPATH__abc_16259_n6084;
  wire AES_CORE_DATAPATH__abc_16259_n6085;
  wire AES_CORE_DATAPATH__abc_16259_n6086;
  wire AES_CORE_DATAPATH__abc_16259_n6087;
  wire AES_CORE_DATAPATH__abc_16259_n6088;
  wire AES_CORE_DATAPATH__abc_16259_n6089;
  wire AES_CORE_DATAPATH__abc_16259_n6090;
  wire AES_CORE_DATAPATH__abc_16259_n6091;
  wire AES_CORE_DATAPATH__abc_16259_n6092;
  wire AES_CORE_DATAPATH__abc_16259_n6092_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n6092_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n6092_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n6092_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n6092_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n6093;
  wire AES_CORE_DATAPATH__abc_16259_n6094;
  wire AES_CORE_DATAPATH__abc_16259_n6095;
  wire AES_CORE_DATAPATH__abc_16259_n6095_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n6095_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n6095_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n6095_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n6095_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n6096;
  wire AES_CORE_DATAPATH__abc_16259_n6097;
  wire AES_CORE_DATAPATH__abc_16259_n6097_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n6097_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n6097_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n6097_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n6097_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n6098;
  wire AES_CORE_DATAPATH__abc_16259_n6099;
  wire AES_CORE_DATAPATH__abc_16259_n6100;
  wire AES_CORE_DATAPATH__abc_16259_n6101;
  wire AES_CORE_DATAPATH__abc_16259_n6101_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n6101_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n6101_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n6101_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n6101_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n6102;
  wire AES_CORE_DATAPATH__abc_16259_n6103;
  wire AES_CORE_DATAPATH__abc_16259_n6104;
  wire AES_CORE_DATAPATH__abc_16259_n6105;
  wire AES_CORE_DATAPATH__abc_16259_n6106;
  wire AES_CORE_DATAPATH__abc_16259_n6107;
  wire AES_CORE_DATAPATH__abc_16259_n6107_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n6107_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n6107_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n6107_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n6107_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n6107_bF_buf5;
  wire AES_CORE_DATAPATH__abc_16259_n6107_bF_buf6;
  wire AES_CORE_DATAPATH__abc_16259_n6107_bF_buf7;
  wire AES_CORE_DATAPATH__abc_16259_n6107_bF_buf8;
  wire AES_CORE_DATAPATH__abc_16259_n6107_bF_buf9;
  wire AES_CORE_DATAPATH__abc_16259_n6108;
  wire AES_CORE_DATAPATH__abc_16259_n6109;
  wire AES_CORE_DATAPATH__abc_16259_n6110;
  wire AES_CORE_DATAPATH__abc_16259_n6111;
  wire AES_CORE_DATAPATH__abc_16259_n6112;
  wire AES_CORE_DATAPATH__abc_16259_n6113;
  wire AES_CORE_DATAPATH__abc_16259_n6115;
  wire AES_CORE_DATAPATH__abc_16259_n6116;
  wire AES_CORE_DATAPATH__abc_16259_n6117;
  wire AES_CORE_DATAPATH__abc_16259_n6118;
  wire AES_CORE_DATAPATH__abc_16259_n6119;
  wire AES_CORE_DATAPATH__abc_16259_n6120;
  wire AES_CORE_DATAPATH__abc_16259_n6121;
  wire AES_CORE_DATAPATH__abc_16259_n6122;
  wire AES_CORE_DATAPATH__abc_16259_n6123;
  wire AES_CORE_DATAPATH__abc_16259_n6124;
  wire AES_CORE_DATAPATH__abc_16259_n6125;
  wire AES_CORE_DATAPATH__abc_16259_n6126;
  wire AES_CORE_DATAPATH__abc_16259_n6127;
  wire AES_CORE_DATAPATH__abc_16259_n6128;
  wire AES_CORE_DATAPATH__abc_16259_n6129;
  wire AES_CORE_DATAPATH__abc_16259_n6130;
  wire AES_CORE_DATAPATH__abc_16259_n6131;
  wire AES_CORE_DATAPATH__abc_16259_n6132;
  wire AES_CORE_DATAPATH__abc_16259_n6133;
  wire AES_CORE_DATAPATH__abc_16259_n6134;
  wire AES_CORE_DATAPATH__abc_16259_n6135;
  wire AES_CORE_DATAPATH__abc_16259_n6136;
  wire AES_CORE_DATAPATH__abc_16259_n6137;
  wire AES_CORE_DATAPATH__abc_16259_n6138;
  wire AES_CORE_DATAPATH__abc_16259_n6139;
  wire AES_CORE_DATAPATH__abc_16259_n6140;
  wire AES_CORE_DATAPATH__abc_16259_n6141;
  wire AES_CORE_DATAPATH__abc_16259_n6142;
  wire AES_CORE_DATAPATH__abc_16259_n6143;
  wire AES_CORE_DATAPATH__abc_16259_n6144;
  wire AES_CORE_DATAPATH__abc_16259_n6145;
  wire AES_CORE_DATAPATH__abc_16259_n6146;
  wire AES_CORE_DATAPATH__abc_16259_n6147;
  wire AES_CORE_DATAPATH__abc_16259_n6148;
  wire AES_CORE_DATAPATH__abc_16259_n6149;
  wire AES_CORE_DATAPATH__abc_16259_n6150;
  wire AES_CORE_DATAPATH__abc_16259_n6151;
  wire AES_CORE_DATAPATH__abc_16259_n6152;
  wire AES_CORE_DATAPATH__abc_16259_n6153;
  wire AES_CORE_DATAPATH__abc_16259_n6154;
  wire AES_CORE_DATAPATH__abc_16259_n6155;
  wire AES_CORE_DATAPATH__abc_16259_n6156;
  wire AES_CORE_DATAPATH__abc_16259_n6157;
  wire AES_CORE_DATAPATH__abc_16259_n6158;
  wire AES_CORE_DATAPATH__abc_16259_n6159;
  wire AES_CORE_DATAPATH__abc_16259_n6160;
  wire AES_CORE_DATAPATH__abc_16259_n6161;
  wire AES_CORE_DATAPATH__abc_16259_n6162;
  wire AES_CORE_DATAPATH__abc_16259_n6164;
  wire AES_CORE_DATAPATH__abc_16259_n6165;
  wire AES_CORE_DATAPATH__abc_16259_n6166;
  wire AES_CORE_DATAPATH__abc_16259_n6167;
  wire AES_CORE_DATAPATH__abc_16259_n6168;
  wire AES_CORE_DATAPATH__abc_16259_n6169;
  wire AES_CORE_DATAPATH__abc_16259_n6170;
  wire AES_CORE_DATAPATH__abc_16259_n6171;
  wire AES_CORE_DATAPATH__abc_16259_n6172;
  wire AES_CORE_DATAPATH__abc_16259_n6173;
  wire AES_CORE_DATAPATH__abc_16259_n6174;
  wire AES_CORE_DATAPATH__abc_16259_n6175;
  wire AES_CORE_DATAPATH__abc_16259_n6176;
  wire AES_CORE_DATAPATH__abc_16259_n6177;
  wire AES_CORE_DATAPATH__abc_16259_n6178;
  wire AES_CORE_DATAPATH__abc_16259_n6179;
  wire AES_CORE_DATAPATH__abc_16259_n6180;
  wire AES_CORE_DATAPATH__abc_16259_n6181;
  wire AES_CORE_DATAPATH__abc_16259_n6182;
  wire AES_CORE_DATAPATH__abc_16259_n6183;
  wire AES_CORE_DATAPATH__abc_16259_n6184;
  wire AES_CORE_DATAPATH__abc_16259_n6185;
  wire AES_CORE_DATAPATH__abc_16259_n6186;
  wire AES_CORE_DATAPATH__abc_16259_n6187;
  wire AES_CORE_DATAPATH__abc_16259_n6188;
  wire AES_CORE_DATAPATH__abc_16259_n6189;
  wire AES_CORE_DATAPATH__abc_16259_n6190;
  wire AES_CORE_DATAPATH__abc_16259_n6191;
  wire AES_CORE_DATAPATH__abc_16259_n6192;
  wire AES_CORE_DATAPATH__abc_16259_n6193;
  wire AES_CORE_DATAPATH__abc_16259_n6194;
  wire AES_CORE_DATAPATH__abc_16259_n6195;
  wire AES_CORE_DATAPATH__abc_16259_n6196;
  wire AES_CORE_DATAPATH__abc_16259_n6197;
  wire AES_CORE_DATAPATH__abc_16259_n6198;
  wire AES_CORE_DATAPATH__abc_16259_n6199;
  wire AES_CORE_DATAPATH__abc_16259_n6200;
  wire AES_CORE_DATAPATH__abc_16259_n6201;
  wire AES_CORE_DATAPATH__abc_16259_n6202;
  wire AES_CORE_DATAPATH__abc_16259_n6203;
  wire AES_CORE_DATAPATH__abc_16259_n6204;
  wire AES_CORE_DATAPATH__abc_16259_n6205;
  wire AES_CORE_DATAPATH__abc_16259_n6206;
  wire AES_CORE_DATAPATH__abc_16259_n6207;
  wire AES_CORE_DATAPATH__abc_16259_n6208;
  wire AES_CORE_DATAPATH__abc_16259_n6209;
  wire AES_CORE_DATAPATH__abc_16259_n6210;
  wire AES_CORE_DATAPATH__abc_16259_n6211;
  wire AES_CORE_DATAPATH__abc_16259_n6213;
  wire AES_CORE_DATAPATH__abc_16259_n6214;
  wire AES_CORE_DATAPATH__abc_16259_n6215;
  wire AES_CORE_DATAPATH__abc_16259_n6216;
  wire AES_CORE_DATAPATH__abc_16259_n6217;
  wire AES_CORE_DATAPATH__abc_16259_n6218;
  wire AES_CORE_DATAPATH__abc_16259_n6219;
  wire AES_CORE_DATAPATH__abc_16259_n6220;
  wire AES_CORE_DATAPATH__abc_16259_n6221;
  wire AES_CORE_DATAPATH__abc_16259_n6222;
  wire AES_CORE_DATAPATH__abc_16259_n6223;
  wire AES_CORE_DATAPATH__abc_16259_n6224;
  wire AES_CORE_DATAPATH__abc_16259_n6225;
  wire AES_CORE_DATAPATH__abc_16259_n6226;
  wire AES_CORE_DATAPATH__abc_16259_n6227;
  wire AES_CORE_DATAPATH__abc_16259_n6228;
  wire AES_CORE_DATAPATH__abc_16259_n6229;
  wire AES_CORE_DATAPATH__abc_16259_n6230;
  wire AES_CORE_DATAPATH__abc_16259_n6231;
  wire AES_CORE_DATAPATH__abc_16259_n6232;
  wire AES_CORE_DATAPATH__abc_16259_n6233;
  wire AES_CORE_DATAPATH__abc_16259_n6234;
  wire AES_CORE_DATAPATH__abc_16259_n6235;
  wire AES_CORE_DATAPATH__abc_16259_n6236;
  wire AES_CORE_DATAPATH__abc_16259_n6237;
  wire AES_CORE_DATAPATH__abc_16259_n6238;
  wire AES_CORE_DATAPATH__abc_16259_n6239;
  wire AES_CORE_DATAPATH__abc_16259_n6240;
  wire AES_CORE_DATAPATH__abc_16259_n6241;
  wire AES_CORE_DATAPATH__abc_16259_n6242;
  wire AES_CORE_DATAPATH__abc_16259_n6243;
  wire AES_CORE_DATAPATH__abc_16259_n6244;
  wire AES_CORE_DATAPATH__abc_16259_n6245;
  wire AES_CORE_DATAPATH__abc_16259_n6246;
  wire AES_CORE_DATAPATH__abc_16259_n6247;
  wire AES_CORE_DATAPATH__abc_16259_n6248;
  wire AES_CORE_DATAPATH__abc_16259_n6249;
  wire AES_CORE_DATAPATH__abc_16259_n6250;
  wire AES_CORE_DATAPATH__abc_16259_n6251;
  wire AES_CORE_DATAPATH__abc_16259_n6252;
  wire AES_CORE_DATAPATH__abc_16259_n6253;
  wire AES_CORE_DATAPATH__abc_16259_n6254;
  wire AES_CORE_DATAPATH__abc_16259_n6255;
  wire AES_CORE_DATAPATH__abc_16259_n6256;
  wire AES_CORE_DATAPATH__abc_16259_n6257;
  wire AES_CORE_DATAPATH__abc_16259_n6258;
  wire AES_CORE_DATAPATH__abc_16259_n6259;
  wire AES_CORE_DATAPATH__abc_16259_n6260;
  wire AES_CORE_DATAPATH__abc_16259_n6262;
  wire AES_CORE_DATAPATH__abc_16259_n6263;
  wire AES_CORE_DATAPATH__abc_16259_n6264;
  wire AES_CORE_DATAPATH__abc_16259_n6265;
  wire AES_CORE_DATAPATH__abc_16259_n6266;
  wire AES_CORE_DATAPATH__abc_16259_n6267;
  wire AES_CORE_DATAPATH__abc_16259_n6268;
  wire AES_CORE_DATAPATH__abc_16259_n6269;
  wire AES_CORE_DATAPATH__abc_16259_n6270;
  wire AES_CORE_DATAPATH__abc_16259_n6271;
  wire AES_CORE_DATAPATH__abc_16259_n6272;
  wire AES_CORE_DATAPATH__abc_16259_n6273;
  wire AES_CORE_DATAPATH__abc_16259_n6274;
  wire AES_CORE_DATAPATH__abc_16259_n6275;
  wire AES_CORE_DATAPATH__abc_16259_n6276;
  wire AES_CORE_DATAPATH__abc_16259_n6277;
  wire AES_CORE_DATAPATH__abc_16259_n6278;
  wire AES_CORE_DATAPATH__abc_16259_n6279;
  wire AES_CORE_DATAPATH__abc_16259_n6280;
  wire AES_CORE_DATAPATH__abc_16259_n6281;
  wire AES_CORE_DATAPATH__abc_16259_n6282;
  wire AES_CORE_DATAPATH__abc_16259_n6283;
  wire AES_CORE_DATAPATH__abc_16259_n6284;
  wire AES_CORE_DATAPATH__abc_16259_n6285;
  wire AES_CORE_DATAPATH__abc_16259_n6286;
  wire AES_CORE_DATAPATH__abc_16259_n6287;
  wire AES_CORE_DATAPATH__abc_16259_n6288;
  wire AES_CORE_DATAPATH__abc_16259_n6289;
  wire AES_CORE_DATAPATH__abc_16259_n6290;
  wire AES_CORE_DATAPATH__abc_16259_n6291;
  wire AES_CORE_DATAPATH__abc_16259_n6292;
  wire AES_CORE_DATAPATH__abc_16259_n6293;
  wire AES_CORE_DATAPATH__abc_16259_n6294;
  wire AES_CORE_DATAPATH__abc_16259_n6295;
  wire AES_CORE_DATAPATH__abc_16259_n6296;
  wire AES_CORE_DATAPATH__abc_16259_n6297;
  wire AES_CORE_DATAPATH__abc_16259_n6298;
  wire AES_CORE_DATAPATH__abc_16259_n6299;
  wire AES_CORE_DATAPATH__abc_16259_n6300;
  wire AES_CORE_DATAPATH__abc_16259_n6301;
  wire AES_CORE_DATAPATH__abc_16259_n6302;
  wire AES_CORE_DATAPATH__abc_16259_n6303;
  wire AES_CORE_DATAPATH__abc_16259_n6304;
  wire AES_CORE_DATAPATH__abc_16259_n6305;
  wire AES_CORE_DATAPATH__abc_16259_n6306;
  wire AES_CORE_DATAPATH__abc_16259_n6307;
  wire AES_CORE_DATAPATH__abc_16259_n6308;
  wire AES_CORE_DATAPATH__abc_16259_n6309;
  wire AES_CORE_DATAPATH__abc_16259_n6311;
  wire AES_CORE_DATAPATH__abc_16259_n6312;
  wire AES_CORE_DATAPATH__abc_16259_n6313;
  wire AES_CORE_DATAPATH__abc_16259_n6314;
  wire AES_CORE_DATAPATH__abc_16259_n6315;
  wire AES_CORE_DATAPATH__abc_16259_n6316;
  wire AES_CORE_DATAPATH__abc_16259_n6317;
  wire AES_CORE_DATAPATH__abc_16259_n6318;
  wire AES_CORE_DATAPATH__abc_16259_n6319;
  wire AES_CORE_DATAPATH__abc_16259_n6320;
  wire AES_CORE_DATAPATH__abc_16259_n6321;
  wire AES_CORE_DATAPATH__abc_16259_n6322;
  wire AES_CORE_DATAPATH__abc_16259_n6323;
  wire AES_CORE_DATAPATH__abc_16259_n6324;
  wire AES_CORE_DATAPATH__abc_16259_n6325;
  wire AES_CORE_DATAPATH__abc_16259_n6326;
  wire AES_CORE_DATAPATH__abc_16259_n6327;
  wire AES_CORE_DATAPATH__abc_16259_n6328;
  wire AES_CORE_DATAPATH__abc_16259_n6329;
  wire AES_CORE_DATAPATH__abc_16259_n6330;
  wire AES_CORE_DATAPATH__abc_16259_n6331;
  wire AES_CORE_DATAPATH__abc_16259_n6332;
  wire AES_CORE_DATAPATH__abc_16259_n6333;
  wire AES_CORE_DATAPATH__abc_16259_n6334;
  wire AES_CORE_DATAPATH__abc_16259_n6335;
  wire AES_CORE_DATAPATH__abc_16259_n6336;
  wire AES_CORE_DATAPATH__abc_16259_n6337;
  wire AES_CORE_DATAPATH__abc_16259_n6338;
  wire AES_CORE_DATAPATH__abc_16259_n6339;
  wire AES_CORE_DATAPATH__abc_16259_n6340;
  wire AES_CORE_DATAPATH__abc_16259_n6341;
  wire AES_CORE_DATAPATH__abc_16259_n6342;
  wire AES_CORE_DATAPATH__abc_16259_n6343;
  wire AES_CORE_DATAPATH__abc_16259_n6344;
  wire AES_CORE_DATAPATH__abc_16259_n6345;
  wire AES_CORE_DATAPATH__abc_16259_n6346;
  wire AES_CORE_DATAPATH__abc_16259_n6347;
  wire AES_CORE_DATAPATH__abc_16259_n6348;
  wire AES_CORE_DATAPATH__abc_16259_n6349;
  wire AES_CORE_DATAPATH__abc_16259_n6350;
  wire AES_CORE_DATAPATH__abc_16259_n6351;
  wire AES_CORE_DATAPATH__abc_16259_n6352;
  wire AES_CORE_DATAPATH__abc_16259_n6353;
  wire AES_CORE_DATAPATH__abc_16259_n6354;
  wire AES_CORE_DATAPATH__abc_16259_n6355;
  wire AES_CORE_DATAPATH__abc_16259_n6356;
  wire AES_CORE_DATAPATH__abc_16259_n6357;
  wire AES_CORE_DATAPATH__abc_16259_n6358;
  wire AES_CORE_DATAPATH__abc_16259_n6360;
  wire AES_CORE_DATAPATH__abc_16259_n6361;
  wire AES_CORE_DATAPATH__abc_16259_n6362;
  wire AES_CORE_DATAPATH__abc_16259_n6363;
  wire AES_CORE_DATAPATH__abc_16259_n6364;
  wire AES_CORE_DATAPATH__abc_16259_n6365;
  wire AES_CORE_DATAPATH__abc_16259_n6366;
  wire AES_CORE_DATAPATH__abc_16259_n6367;
  wire AES_CORE_DATAPATH__abc_16259_n6368;
  wire AES_CORE_DATAPATH__abc_16259_n6369;
  wire AES_CORE_DATAPATH__abc_16259_n6370;
  wire AES_CORE_DATAPATH__abc_16259_n6371;
  wire AES_CORE_DATAPATH__abc_16259_n6372;
  wire AES_CORE_DATAPATH__abc_16259_n6373;
  wire AES_CORE_DATAPATH__abc_16259_n6374;
  wire AES_CORE_DATAPATH__abc_16259_n6375;
  wire AES_CORE_DATAPATH__abc_16259_n6376;
  wire AES_CORE_DATAPATH__abc_16259_n6377;
  wire AES_CORE_DATAPATH__abc_16259_n6378;
  wire AES_CORE_DATAPATH__abc_16259_n6379;
  wire AES_CORE_DATAPATH__abc_16259_n6380;
  wire AES_CORE_DATAPATH__abc_16259_n6381;
  wire AES_CORE_DATAPATH__abc_16259_n6382;
  wire AES_CORE_DATAPATH__abc_16259_n6383;
  wire AES_CORE_DATAPATH__abc_16259_n6384;
  wire AES_CORE_DATAPATH__abc_16259_n6385;
  wire AES_CORE_DATAPATH__abc_16259_n6386;
  wire AES_CORE_DATAPATH__abc_16259_n6387;
  wire AES_CORE_DATAPATH__abc_16259_n6388;
  wire AES_CORE_DATAPATH__abc_16259_n6389;
  wire AES_CORE_DATAPATH__abc_16259_n6390;
  wire AES_CORE_DATAPATH__abc_16259_n6391;
  wire AES_CORE_DATAPATH__abc_16259_n6392;
  wire AES_CORE_DATAPATH__abc_16259_n6393;
  wire AES_CORE_DATAPATH__abc_16259_n6394;
  wire AES_CORE_DATAPATH__abc_16259_n6395;
  wire AES_CORE_DATAPATH__abc_16259_n6396;
  wire AES_CORE_DATAPATH__abc_16259_n6397;
  wire AES_CORE_DATAPATH__abc_16259_n6398;
  wire AES_CORE_DATAPATH__abc_16259_n6399;
  wire AES_CORE_DATAPATH__abc_16259_n6400;
  wire AES_CORE_DATAPATH__abc_16259_n6401;
  wire AES_CORE_DATAPATH__abc_16259_n6402;
  wire AES_CORE_DATAPATH__abc_16259_n6403;
  wire AES_CORE_DATAPATH__abc_16259_n6404;
  wire AES_CORE_DATAPATH__abc_16259_n6405;
  wire AES_CORE_DATAPATH__abc_16259_n6406;
  wire AES_CORE_DATAPATH__abc_16259_n6407;
  wire AES_CORE_DATAPATH__abc_16259_n6409;
  wire AES_CORE_DATAPATH__abc_16259_n6410;
  wire AES_CORE_DATAPATH__abc_16259_n6411;
  wire AES_CORE_DATAPATH__abc_16259_n6412;
  wire AES_CORE_DATAPATH__abc_16259_n6413;
  wire AES_CORE_DATAPATH__abc_16259_n6414;
  wire AES_CORE_DATAPATH__abc_16259_n6415;
  wire AES_CORE_DATAPATH__abc_16259_n6416;
  wire AES_CORE_DATAPATH__abc_16259_n6417;
  wire AES_CORE_DATAPATH__abc_16259_n6418;
  wire AES_CORE_DATAPATH__abc_16259_n6419;
  wire AES_CORE_DATAPATH__abc_16259_n6420;
  wire AES_CORE_DATAPATH__abc_16259_n6421;
  wire AES_CORE_DATAPATH__abc_16259_n6422;
  wire AES_CORE_DATAPATH__abc_16259_n6423;
  wire AES_CORE_DATAPATH__abc_16259_n6424;
  wire AES_CORE_DATAPATH__abc_16259_n6425;
  wire AES_CORE_DATAPATH__abc_16259_n6426;
  wire AES_CORE_DATAPATH__abc_16259_n6427;
  wire AES_CORE_DATAPATH__abc_16259_n6428;
  wire AES_CORE_DATAPATH__abc_16259_n6429;
  wire AES_CORE_DATAPATH__abc_16259_n6430;
  wire AES_CORE_DATAPATH__abc_16259_n6431;
  wire AES_CORE_DATAPATH__abc_16259_n6432;
  wire AES_CORE_DATAPATH__abc_16259_n6433;
  wire AES_CORE_DATAPATH__abc_16259_n6434;
  wire AES_CORE_DATAPATH__abc_16259_n6435;
  wire AES_CORE_DATAPATH__abc_16259_n6436;
  wire AES_CORE_DATAPATH__abc_16259_n6437;
  wire AES_CORE_DATAPATH__abc_16259_n6438;
  wire AES_CORE_DATAPATH__abc_16259_n6439;
  wire AES_CORE_DATAPATH__abc_16259_n6440;
  wire AES_CORE_DATAPATH__abc_16259_n6441;
  wire AES_CORE_DATAPATH__abc_16259_n6442;
  wire AES_CORE_DATAPATH__abc_16259_n6443;
  wire AES_CORE_DATAPATH__abc_16259_n6444;
  wire AES_CORE_DATAPATH__abc_16259_n6445;
  wire AES_CORE_DATAPATH__abc_16259_n6446;
  wire AES_CORE_DATAPATH__abc_16259_n6447;
  wire AES_CORE_DATAPATH__abc_16259_n6448;
  wire AES_CORE_DATAPATH__abc_16259_n6449;
  wire AES_CORE_DATAPATH__abc_16259_n6450;
  wire AES_CORE_DATAPATH__abc_16259_n6451;
  wire AES_CORE_DATAPATH__abc_16259_n6452;
  wire AES_CORE_DATAPATH__abc_16259_n6453;
  wire AES_CORE_DATAPATH__abc_16259_n6454;
  wire AES_CORE_DATAPATH__abc_16259_n6455;
  wire AES_CORE_DATAPATH__abc_16259_n6456;
  wire AES_CORE_DATAPATH__abc_16259_n6458;
  wire AES_CORE_DATAPATH__abc_16259_n6459;
  wire AES_CORE_DATAPATH__abc_16259_n6460;
  wire AES_CORE_DATAPATH__abc_16259_n6461;
  wire AES_CORE_DATAPATH__abc_16259_n6462;
  wire AES_CORE_DATAPATH__abc_16259_n6463;
  wire AES_CORE_DATAPATH__abc_16259_n6464;
  wire AES_CORE_DATAPATH__abc_16259_n6465;
  wire AES_CORE_DATAPATH__abc_16259_n6466;
  wire AES_CORE_DATAPATH__abc_16259_n6467;
  wire AES_CORE_DATAPATH__abc_16259_n6468;
  wire AES_CORE_DATAPATH__abc_16259_n6469;
  wire AES_CORE_DATAPATH__abc_16259_n6470;
  wire AES_CORE_DATAPATH__abc_16259_n6471;
  wire AES_CORE_DATAPATH__abc_16259_n6472;
  wire AES_CORE_DATAPATH__abc_16259_n6473;
  wire AES_CORE_DATAPATH__abc_16259_n6474;
  wire AES_CORE_DATAPATH__abc_16259_n6475;
  wire AES_CORE_DATAPATH__abc_16259_n6476;
  wire AES_CORE_DATAPATH__abc_16259_n6477;
  wire AES_CORE_DATAPATH__abc_16259_n6478;
  wire AES_CORE_DATAPATH__abc_16259_n6479;
  wire AES_CORE_DATAPATH__abc_16259_n6480;
  wire AES_CORE_DATAPATH__abc_16259_n6481;
  wire AES_CORE_DATAPATH__abc_16259_n6482;
  wire AES_CORE_DATAPATH__abc_16259_n6483;
  wire AES_CORE_DATAPATH__abc_16259_n6484;
  wire AES_CORE_DATAPATH__abc_16259_n6485;
  wire AES_CORE_DATAPATH__abc_16259_n6486;
  wire AES_CORE_DATAPATH__abc_16259_n6487;
  wire AES_CORE_DATAPATH__abc_16259_n6488;
  wire AES_CORE_DATAPATH__abc_16259_n6489;
  wire AES_CORE_DATAPATH__abc_16259_n6490;
  wire AES_CORE_DATAPATH__abc_16259_n6491;
  wire AES_CORE_DATAPATH__abc_16259_n6492;
  wire AES_CORE_DATAPATH__abc_16259_n6493;
  wire AES_CORE_DATAPATH__abc_16259_n6494;
  wire AES_CORE_DATAPATH__abc_16259_n6495;
  wire AES_CORE_DATAPATH__abc_16259_n6496;
  wire AES_CORE_DATAPATH__abc_16259_n6497;
  wire AES_CORE_DATAPATH__abc_16259_n6498;
  wire AES_CORE_DATAPATH__abc_16259_n6499;
  wire AES_CORE_DATAPATH__abc_16259_n6500;
  wire AES_CORE_DATAPATH__abc_16259_n6501;
  wire AES_CORE_DATAPATH__abc_16259_n6502;
  wire AES_CORE_DATAPATH__abc_16259_n6503;
  wire AES_CORE_DATAPATH__abc_16259_n6504;
  wire AES_CORE_DATAPATH__abc_16259_n6505;
  wire AES_CORE_DATAPATH__abc_16259_n6507;
  wire AES_CORE_DATAPATH__abc_16259_n6508;
  wire AES_CORE_DATAPATH__abc_16259_n6509;
  wire AES_CORE_DATAPATH__abc_16259_n6510;
  wire AES_CORE_DATAPATH__abc_16259_n6511;
  wire AES_CORE_DATAPATH__abc_16259_n6512;
  wire AES_CORE_DATAPATH__abc_16259_n6513;
  wire AES_CORE_DATAPATH__abc_16259_n6514;
  wire AES_CORE_DATAPATH__abc_16259_n6515;
  wire AES_CORE_DATAPATH__abc_16259_n6516;
  wire AES_CORE_DATAPATH__abc_16259_n6517;
  wire AES_CORE_DATAPATH__abc_16259_n6518;
  wire AES_CORE_DATAPATH__abc_16259_n6519;
  wire AES_CORE_DATAPATH__abc_16259_n6520;
  wire AES_CORE_DATAPATH__abc_16259_n6521;
  wire AES_CORE_DATAPATH__abc_16259_n6522;
  wire AES_CORE_DATAPATH__abc_16259_n6523;
  wire AES_CORE_DATAPATH__abc_16259_n6524;
  wire AES_CORE_DATAPATH__abc_16259_n6525;
  wire AES_CORE_DATAPATH__abc_16259_n6526;
  wire AES_CORE_DATAPATH__abc_16259_n6527;
  wire AES_CORE_DATAPATH__abc_16259_n6528;
  wire AES_CORE_DATAPATH__abc_16259_n6529;
  wire AES_CORE_DATAPATH__abc_16259_n6530;
  wire AES_CORE_DATAPATH__abc_16259_n6531;
  wire AES_CORE_DATAPATH__abc_16259_n6532;
  wire AES_CORE_DATAPATH__abc_16259_n6533;
  wire AES_CORE_DATAPATH__abc_16259_n6534;
  wire AES_CORE_DATAPATH__abc_16259_n6535;
  wire AES_CORE_DATAPATH__abc_16259_n6536;
  wire AES_CORE_DATAPATH__abc_16259_n6537;
  wire AES_CORE_DATAPATH__abc_16259_n6538;
  wire AES_CORE_DATAPATH__abc_16259_n6539;
  wire AES_CORE_DATAPATH__abc_16259_n6540;
  wire AES_CORE_DATAPATH__abc_16259_n6541;
  wire AES_CORE_DATAPATH__abc_16259_n6542;
  wire AES_CORE_DATAPATH__abc_16259_n6543;
  wire AES_CORE_DATAPATH__abc_16259_n6544;
  wire AES_CORE_DATAPATH__abc_16259_n6545;
  wire AES_CORE_DATAPATH__abc_16259_n6546;
  wire AES_CORE_DATAPATH__abc_16259_n6547;
  wire AES_CORE_DATAPATH__abc_16259_n6548;
  wire AES_CORE_DATAPATH__abc_16259_n6549;
  wire AES_CORE_DATAPATH__abc_16259_n6550;
  wire AES_CORE_DATAPATH__abc_16259_n6551;
  wire AES_CORE_DATAPATH__abc_16259_n6552;
  wire AES_CORE_DATAPATH__abc_16259_n6553;
  wire AES_CORE_DATAPATH__abc_16259_n6554;
  wire AES_CORE_DATAPATH__abc_16259_n6556;
  wire AES_CORE_DATAPATH__abc_16259_n6557;
  wire AES_CORE_DATAPATH__abc_16259_n6558;
  wire AES_CORE_DATAPATH__abc_16259_n6559;
  wire AES_CORE_DATAPATH__abc_16259_n6560;
  wire AES_CORE_DATAPATH__abc_16259_n6561;
  wire AES_CORE_DATAPATH__abc_16259_n6562;
  wire AES_CORE_DATAPATH__abc_16259_n6563;
  wire AES_CORE_DATAPATH__abc_16259_n6564;
  wire AES_CORE_DATAPATH__abc_16259_n6565;
  wire AES_CORE_DATAPATH__abc_16259_n6566;
  wire AES_CORE_DATAPATH__abc_16259_n6567;
  wire AES_CORE_DATAPATH__abc_16259_n6568;
  wire AES_CORE_DATAPATH__abc_16259_n6569;
  wire AES_CORE_DATAPATH__abc_16259_n6570;
  wire AES_CORE_DATAPATH__abc_16259_n6571;
  wire AES_CORE_DATAPATH__abc_16259_n6572;
  wire AES_CORE_DATAPATH__abc_16259_n6573;
  wire AES_CORE_DATAPATH__abc_16259_n6574;
  wire AES_CORE_DATAPATH__abc_16259_n6575;
  wire AES_CORE_DATAPATH__abc_16259_n6576;
  wire AES_CORE_DATAPATH__abc_16259_n6577;
  wire AES_CORE_DATAPATH__abc_16259_n6578;
  wire AES_CORE_DATAPATH__abc_16259_n6579;
  wire AES_CORE_DATAPATH__abc_16259_n6580;
  wire AES_CORE_DATAPATH__abc_16259_n6581;
  wire AES_CORE_DATAPATH__abc_16259_n6582;
  wire AES_CORE_DATAPATH__abc_16259_n6583;
  wire AES_CORE_DATAPATH__abc_16259_n6584;
  wire AES_CORE_DATAPATH__abc_16259_n6585;
  wire AES_CORE_DATAPATH__abc_16259_n6586;
  wire AES_CORE_DATAPATH__abc_16259_n6587;
  wire AES_CORE_DATAPATH__abc_16259_n6588;
  wire AES_CORE_DATAPATH__abc_16259_n6589;
  wire AES_CORE_DATAPATH__abc_16259_n6590;
  wire AES_CORE_DATAPATH__abc_16259_n6591;
  wire AES_CORE_DATAPATH__abc_16259_n6592;
  wire AES_CORE_DATAPATH__abc_16259_n6593;
  wire AES_CORE_DATAPATH__abc_16259_n6594;
  wire AES_CORE_DATAPATH__abc_16259_n6595;
  wire AES_CORE_DATAPATH__abc_16259_n6596;
  wire AES_CORE_DATAPATH__abc_16259_n6597;
  wire AES_CORE_DATAPATH__abc_16259_n6598;
  wire AES_CORE_DATAPATH__abc_16259_n6599;
  wire AES_CORE_DATAPATH__abc_16259_n6600;
  wire AES_CORE_DATAPATH__abc_16259_n6601;
  wire AES_CORE_DATAPATH__abc_16259_n6602;
  wire AES_CORE_DATAPATH__abc_16259_n6603;
  wire AES_CORE_DATAPATH__abc_16259_n6603_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n6603_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n6603_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n6603_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n6604;
  wire AES_CORE_DATAPATH__abc_16259_n6605;
  wire AES_CORE_DATAPATH__abc_16259_n6606;
  wire AES_CORE_DATAPATH__abc_16259_n6607;
  wire AES_CORE_DATAPATH__abc_16259_n6608;
  wire AES_CORE_DATAPATH__abc_16259_n6609;
  wire AES_CORE_DATAPATH__abc_16259_n6610;
  wire AES_CORE_DATAPATH__abc_16259_n6611;
  wire AES_CORE_DATAPATH__abc_16259_n6612;
  wire AES_CORE_DATAPATH__abc_16259_n6613;
  wire AES_CORE_DATAPATH__abc_16259_n6615;
  wire AES_CORE_DATAPATH__abc_16259_n6616;
  wire AES_CORE_DATAPATH__abc_16259_n6617;
  wire AES_CORE_DATAPATH__abc_16259_n6618;
  wire AES_CORE_DATAPATH__abc_16259_n6619;
  wire AES_CORE_DATAPATH__abc_16259_n6620;
  wire AES_CORE_DATAPATH__abc_16259_n6621;
  wire AES_CORE_DATAPATH__abc_16259_n6622;
  wire AES_CORE_DATAPATH__abc_16259_n6623;
  wire AES_CORE_DATAPATH__abc_16259_n6624;
  wire AES_CORE_DATAPATH__abc_16259_n6625;
  wire AES_CORE_DATAPATH__abc_16259_n6626;
  wire AES_CORE_DATAPATH__abc_16259_n6627;
  wire AES_CORE_DATAPATH__abc_16259_n6628;
  wire AES_CORE_DATAPATH__abc_16259_n6629;
  wire AES_CORE_DATAPATH__abc_16259_n6630;
  wire AES_CORE_DATAPATH__abc_16259_n6631;
  wire AES_CORE_DATAPATH__abc_16259_n6632;
  wire AES_CORE_DATAPATH__abc_16259_n6633;
  wire AES_CORE_DATAPATH__abc_16259_n6634;
  wire AES_CORE_DATAPATH__abc_16259_n6635;
  wire AES_CORE_DATAPATH__abc_16259_n6636;
  wire AES_CORE_DATAPATH__abc_16259_n6637;
  wire AES_CORE_DATAPATH__abc_16259_n6638;
  wire AES_CORE_DATAPATH__abc_16259_n6639;
  wire AES_CORE_DATAPATH__abc_16259_n6640;
  wire AES_CORE_DATAPATH__abc_16259_n6641;
  wire AES_CORE_DATAPATH__abc_16259_n6642;
  wire AES_CORE_DATAPATH__abc_16259_n6643;
  wire AES_CORE_DATAPATH__abc_16259_n6644;
  wire AES_CORE_DATAPATH__abc_16259_n6645;
  wire AES_CORE_DATAPATH__abc_16259_n6646;
  wire AES_CORE_DATAPATH__abc_16259_n6647;
  wire AES_CORE_DATAPATH__abc_16259_n6648;
  wire AES_CORE_DATAPATH__abc_16259_n6649;
  wire AES_CORE_DATAPATH__abc_16259_n6650;
  wire AES_CORE_DATAPATH__abc_16259_n6651;
  wire AES_CORE_DATAPATH__abc_16259_n6652;
  wire AES_CORE_DATAPATH__abc_16259_n6653;
  wire AES_CORE_DATAPATH__abc_16259_n6654;
  wire AES_CORE_DATAPATH__abc_16259_n6655;
  wire AES_CORE_DATAPATH__abc_16259_n6656;
  wire AES_CORE_DATAPATH__abc_16259_n6657;
  wire AES_CORE_DATAPATH__abc_16259_n6658;
  wire AES_CORE_DATAPATH__abc_16259_n6659;
  wire AES_CORE_DATAPATH__abc_16259_n6660;
  wire AES_CORE_DATAPATH__abc_16259_n6661;
  wire AES_CORE_DATAPATH__abc_16259_n6662;
  wire AES_CORE_DATAPATH__abc_16259_n6663;
  wire AES_CORE_DATAPATH__abc_16259_n6664;
  wire AES_CORE_DATAPATH__abc_16259_n6665;
  wire AES_CORE_DATAPATH__abc_16259_n6666;
  wire AES_CORE_DATAPATH__abc_16259_n6667;
  wire AES_CORE_DATAPATH__abc_16259_n6669;
  wire AES_CORE_DATAPATH__abc_16259_n6670;
  wire AES_CORE_DATAPATH__abc_16259_n6671;
  wire AES_CORE_DATAPATH__abc_16259_n6672;
  wire AES_CORE_DATAPATH__abc_16259_n6673;
  wire AES_CORE_DATAPATH__abc_16259_n6674;
  wire AES_CORE_DATAPATH__abc_16259_n6675;
  wire AES_CORE_DATAPATH__abc_16259_n6676;
  wire AES_CORE_DATAPATH__abc_16259_n6677;
  wire AES_CORE_DATAPATH__abc_16259_n6678;
  wire AES_CORE_DATAPATH__abc_16259_n6679;
  wire AES_CORE_DATAPATH__abc_16259_n6680;
  wire AES_CORE_DATAPATH__abc_16259_n6681;
  wire AES_CORE_DATAPATH__abc_16259_n6682;
  wire AES_CORE_DATAPATH__abc_16259_n6683;
  wire AES_CORE_DATAPATH__abc_16259_n6684;
  wire AES_CORE_DATAPATH__abc_16259_n6685;
  wire AES_CORE_DATAPATH__abc_16259_n6686;
  wire AES_CORE_DATAPATH__abc_16259_n6687;
  wire AES_CORE_DATAPATH__abc_16259_n6688;
  wire AES_CORE_DATAPATH__abc_16259_n6689;
  wire AES_CORE_DATAPATH__abc_16259_n6690;
  wire AES_CORE_DATAPATH__abc_16259_n6691;
  wire AES_CORE_DATAPATH__abc_16259_n6692;
  wire AES_CORE_DATAPATH__abc_16259_n6693;
  wire AES_CORE_DATAPATH__abc_16259_n6694;
  wire AES_CORE_DATAPATH__abc_16259_n6695;
  wire AES_CORE_DATAPATH__abc_16259_n6696;
  wire AES_CORE_DATAPATH__abc_16259_n6697;
  wire AES_CORE_DATAPATH__abc_16259_n6698;
  wire AES_CORE_DATAPATH__abc_16259_n6699;
  wire AES_CORE_DATAPATH__abc_16259_n6700;
  wire AES_CORE_DATAPATH__abc_16259_n6701;
  wire AES_CORE_DATAPATH__abc_16259_n6702;
  wire AES_CORE_DATAPATH__abc_16259_n6703;
  wire AES_CORE_DATAPATH__abc_16259_n6704;
  wire AES_CORE_DATAPATH__abc_16259_n6705;
  wire AES_CORE_DATAPATH__abc_16259_n6706;
  wire AES_CORE_DATAPATH__abc_16259_n6707;
  wire AES_CORE_DATAPATH__abc_16259_n6708;
  wire AES_CORE_DATAPATH__abc_16259_n6709;
  wire AES_CORE_DATAPATH__abc_16259_n6710;
  wire AES_CORE_DATAPATH__abc_16259_n6711;
  wire AES_CORE_DATAPATH__abc_16259_n6712;
  wire AES_CORE_DATAPATH__abc_16259_n6713;
  wire AES_CORE_DATAPATH__abc_16259_n6714;
  wire AES_CORE_DATAPATH__abc_16259_n6715;
  wire AES_CORE_DATAPATH__abc_16259_n6716;
  wire AES_CORE_DATAPATH__abc_16259_n6718;
  wire AES_CORE_DATAPATH__abc_16259_n6719;
  wire AES_CORE_DATAPATH__abc_16259_n6720;
  wire AES_CORE_DATAPATH__abc_16259_n6721;
  wire AES_CORE_DATAPATH__abc_16259_n6722;
  wire AES_CORE_DATAPATH__abc_16259_n6723;
  wire AES_CORE_DATAPATH__abc_16259_n6724;
  wire AES_CORE_DATAPATH__abc_16259_n6725;
  wire AES_CORE_DATAPATH__abc_16259_n6726;
  wire AES_CORE_DATAPATH__abc_16259_n6727;
  wire AES_CORE_DATAPATH__abc_16259_n6728;
  wire AES_CORE_DATAPATH__abc_16259_n6729;
  wire AES_CORE_DATAPATH__abc_16259_n6730;
  wire AES_CORE_DATAPATH__abc_16259_n6731;
  wire AES_CORE_DATAPATH__abc_16259_n6732;
  wire AES_CORE_DATAPATH__abc_16259_n6733;
  wire AES_CORE_DATAPATH__abc_16259_n6734;
  wire AES_CORE_DATAPATH__abc_16259_n6735;
  wire AES_CORE_DATAPATH__abc_16259_n6736;
  wire AES_CORE_DATAPATH__abc_16259_n6737;
  wire AES_CORE_DATAPATH__abc_16259_n6738;
  wire AES_CORE_DATAPATH__abc_16259_n6739;
  wire AES_CORE_DATAPATH__abc_16259_n6740;
  wire AES_CORE_DATAPATH__abc_16259_n6741;
  wire AES_CORE_DATAPATH__abc_16259_n6742;
  wire AES_CORE_DATAPATH__abc_16259_n6743;
  wire AES_CORE_DATAPATH__abc_16259_n6744;
  wire AES_CORE_DATAPATH__abc_16259_n6745;
  wire AES_CORE_DATAPATH__abc_16259_n6746;
  wire AES_CORE_DATAPATH__abc_16259_n6747;
  wire AES_CORE_DATAPATH__abc_16259_n6748;
  wire AES_CORE_DATAPATH__abc_16259_n6749;
  wire AES_CORE_DATAPATH__abc_16259_n6750;
  wire AES_CORE_DATAPATH__abc_16259_n6751;
  wire AES_CORE_DATAPATH__abc_16259_n6752;
  wire AES_CORE_DATAPATH__abc_16259_n6753;
  wire AES_CORE_DATAPATH__abc_16259_n6754;
  wire AES_CORE_DATAPATH__abc_16259_n6755;
  wire AES_CORE_DATAPATH__abc_16259_n6756;
  wire AES_CORE_DATAPATH__abc_16259_n6757;
  wire AES_CORE_DATAPATH__abc_16259_n6758;
  wire AES_CORE_DATAPATH__abc_16259_n6759;
  wire AES_CORE_DATAPATH__abc_16259_n6760;
  wire AES_CORE_DATAPATH__abc_16259_n6761;
  wire AES_CORE_DATAPATH__abc_16259_n6762;
  wire AES_CORE_DATAPATH__abc_16259_n6763;
  wire AES_CORE_DATAPATH__abc_16259_n6764;
  wire AES_CORE_DATAPATH__abc_16259_n6765;
  wire AES_CORE_DATAPATH__abc_16259_n6766;
  wire AES_CORE_DATAPATH__abc_16259_n6767;
  wire AES_CORE_DATAPATH__abc_16259_n6768;
  wire AES_CORE_DATAPATH__abc_16259_n6769;
  wire AES_CORE_DATAPATH__abc_16259_n6770;
  wire AES_CORE_DATAPATH__abc_16259_n6772;
  wire AES_CORE_DATAPATH__abc_16259_n6773;
  wire AES_CORE_DATAPATH__abc_16259_n6774;
  wire AES_CORE_DATAPATH__abc_16259_n6775;
  wire AES_CORE_DATAPATH__abc_16259_n6776;
  wire AES_CORE_DATAPATH__abc_16259_n6777;
  wire AES_CORE_DATAPATH__abc_16259_n6778;
  wire AES_CORE_DATAPATH__abc_16259_n6779;
  wire AES_CORE_DATAPATH__abc_16259_n6780;
  wire AES_CORE_DATAPATH__abc_16259_n6781;
  wire AES_CORE_DATAPATH__abc_16259_n6782;
  wire AES_CORE_DATAPATH__abc_16259_n6783;
  wire AES_CORE_DATAPATH__abc_16259_n6784;
  wire AES_CORE_DATAPATH__abc_16259_n6785;
  wire AES_CORE_DATAPATH__abc_16259_n6786;
  wire AES_CORE_DATAPATH__abc_16259_n6787;
  wire AES_CORE_DATAPATH__abc_16259_n6788;
  wire AES_CORE_DATAPATH__abc_16259_n6789;
  wire AES_CORE_DATAPATH__abc_16259_n6790;
  wire AES_CORE_DATAPATH__abc_16259_n6791;
  wire AES_CORE_DATAPATH__abc_16259_n6792;
  wire AES_CORE_DATAPATH__abc_16259_n6793;
  wire AES_CORE_DATAPATH__abc_16259_n6794;
  wire AES_CORE_DATAPATH__abc_16259_n6795;
  wire AES_CORE_DATAPATH__abc_16259_n6796;
  wire AES_CORE_DATAPATH__abc_16259_n6797;
  wire AES_CORE_DATAPATH__abc_16259_n6798;
  wire AES_CORE_DATAPATH__abc_16259_n6799;
  wire AES_CORE_DATAPATH__abc_16259_n6800;
  wire AES_CORE_DATAPATH__abc_16259_n6801;
  wire AES_CORE_DATAPATH__abc_16259_n6802;
  wire AES_CORE_DATAPATH__abc_16259_n6803;
  wire AES_CORE_DATAPATH__abc_16259_n6804;
  wire AES_CORE_DATAPATH__abc_16259_n6805;
  wire AES_CORE_DATAPATH__abc_16259_n6806;
  wire AES_CORE_DATAPATH__abc_16259_n6807;
  wire AES_CORE_DATAPATH__abc_16259_n6808;
  wire AES_CORE_DATAPATH__abc_16259_n6809;
  wire AES_CORE_DATAPATH__abc_16259_n6810;
  wire AES_CORE_DATAPATH__abc_16259_n6811;
  wire AES_CORE_DATAPATH__abc_16259_n6812;
  wire AES_CORE_DATAPATH__abc_16259_n6813;
  wire AES_CORE_DATAPATH__abc_16259_n6814;
  wire AES_CORE_DATAPATH__abc_16259_n6815;
  wire AES_CORE_DATAPATH__abc_16259_n6816;
  wire AES_CORE_DATAPATH__abc_16259_n6817;
  wire AES_CORE_DATAPATH__abc_16259_n6818;
  wire AES_CORE_DATAPATH__abc_16259_n6819;
  wire AES_CORE_DATAPATH__abc_16259_n6821;
  wire AES_CORE_DATAPATH__abc_16259_n6822;
  wire AES_CORE_DATAPATH__abc_16259_n6823;
  wire AES_CORE_DATAPATH__abc_16259_n6824;
  wire AES_CORE_DATAPATH__abc_16259_n6825;
  wire AES_CORE_DATAPATH__abc_16259_n6826;
  wire AES_CORE_DATAPATH__abc_16259_n6827;
  wire AES_CORE_DATAPATH__abc_16259_n6828;
  wire AES_CORE_DATAPATH__abc_16259_n6829;
  wire AES_CORE_DATAPATH__abc_16259_n6830;
  wire AES_CORE_DATAPATH__abc_16259_n6831;
  wire AES_CORE_DATAPATH__abc_16259_n6832;
  wire AES_CORE_DATAPATH__abc_16259_n6833;
  wire AES_CORE_DATAPATH__abc_16259_n6834;
  wire AES_CORE_DATAPATH__abc_16259_n6835;
  wire AES_CORE_DATAPATH__abc_16259_n6836;
  wire AES_CORE_DATAPATH__abc_16259_n6837;
  wire AES_CORE_DATAPATH__abc_16259_n6838;
  wire AES_CORE_DATAPATH__abc_16259_n6839;
  wire AES_CORE_DATAPATH__abc_16259_n6840;
  wire AES_CORE_DATAPATH__abc_16259_n6841;
  wire AES_CORE_DATAPATH__abc_16259_n6842;
  wire AES_CORE_DATAPATH__abc_16259_n6843;
  wire AES_CORE_DATAPATH__abc_16259_n6844;
  wire AES_CORE_DATAPATH__abc_16259_n6845;
  wire AES_CORE_DATAPATH__abc_16259_n6846;
  wire AES_CORE_DATAPATH__abc_16259_n6847;
  wire AES_CORE_DATAPATH__abc_16259_n6848;
  wire AES_CORE_DATAPATH__abc_16259_n6849;
  wire AES_CORE_DATAPATH__abc_16259_n6850;
  wire AES_CORE_DATAPATH__abc_16259_n6851;
  wire AES_CORE_DATAPATH__abc_16259_n6852;
  wire AES_CORE_DATAPATH__abc_16259_n6853;
  wire AES_CORE_DATAPATH__abc_16259_n6854;
  wire AES_CORE_DATAPATH__abc_16259_n6855;
  wire AES_CORE_DATAPATH__abc_16259_n6856;
  wire AES_CORE_DATAPATH__abc_16259_n6857;
  wire AES_CORE_DATAPATH__abc_16259_n6858;
  wire AES_CORE_DATAPATH__abc_16259_n6859;
  wire AES_CORE_DATAPATH__abc_16259_n6860;
  wire AES_CORE_DATAPATH__abc_16259_n6861;
  wire AES_CORE_DATAPATH__abc_16259_n6862;
  wire AES_CORE_DATAPATH__abc_16259_n6863;
  wire AES_CORE_DATAPATH__abc_16259_n6864;
  wire AES_CORE_DATAPATH__abc_16259_n6865;
  wire AES_CORE_DATAPATH__abc_16259_n6866;
  wire AES_CORE_DATAPATH__abc_16259_n6867;
  wire AES_CORE_DATAPATH__abc_16259_n6868;
  wire AES_CORE_DATAPATH__abc_16259_n6869;
  wire AES_CORE_DATAPATH__abc_16259_n6870;
  wire AES_CORE_DATAPATH__abc_16259_n6871;
  wire AES_CORE_DATAPATH__abc_16259_n6872;
  wire AES_CORE_DATAPATH__abc_16259_n6873;
  wire AES_CORE_DATAPATH__abc_16259_n6875;
  wire AES_CORE_DATAPATH__abc_16259_n6876;
  wire AES_CORE_DATAPATH__abc_16259_n6877;
  wire AES_CORE_DATAPATH__abc_16259_n6878;
  wire AES_CORE_DATAPATH__abc_16259_n6879;
  wire AES_CORE_DATAPATH__abc_16259_n6880;
  wire AES_CORE_DATAPATH__abc_16259_n6881;
  wire AES_CORE_DATAPATH__abc_16259_n6882;
  wire AES_CORE_DATAPATH__abc_16259_n6883;
  wire AES_CORE_DATAPATH__abc_16259_n6884;
  wire AES_CORE_DATAPATH__abc_16259_n6885;
  wire AES_CORE_DATAPATH__abc_16259_n6886;
  wire AES_CORE_DATAPATH__abc_16259_n6887;
  wire AES_CORE_DATAPATH__abc_16259_n6888;
  wire AES_CORE_DATAPATH__abc_16259_n6889;
  wire AES_CORE_DATAPATH__abc_16259_n6890;
  wire AES_CORE_DATAPATH__abc_16259_n6891;
  wire AES_CORE_DATAPATH__abc_16259_n6892;
  wire AES_CORE_DATAPATH__abc_16259_n6893;
  wire AES_CORE_DATAPATH__abc_16259_n6894;
  wire AES_CORE_DATAPATH__abc_16259_n6895;
  wire AES_CORE_DATAPATH__abc_16259_n6896;
  wire AES_CORE_DATAPATH__abc_16259_n6897;
  wire AES_CORE_DATAPATH__abc_16259_n6898;
  wire AES_CORE_DATAPATH__abc_16259_n6899;
  wire AES_CORE_DATAPATH__abc_16259_n6900;
  wire AES_CORE_DATAPATH__abc_16259_n6901;
  wire AES_CORE_DATAPATH__abc_16259_n6902;
  wire AES_CORE_DATAPATH__abc_16259_n6903;
  wire AES_CORE_DATAPATH__abc_16259_n6904;
  wire AES_CORE_DATAPATH__abc_16259_n6905;
  wire AES_CORE_DATAPATH__abc_16259_n6906;
  wire AES_CORE_DATAPATH__abc_16259_n6907;
  wire AES_CORE_DATAPATH__abc_16259_n6908;
  wire AES_CORE_DATAPATH__abc_16259_n6909;
  wire AES_CORE_DATAPATH__abc_16259_n6910;
  wire AES_CORE_DATAPATH__abc_16259_n6911;
  wire AES_CORE_DATAPATH__abc_16259_n6912;
  wire AES_CORE_DATAPATH__abc_16259_n6913;
  wire AES_CORE_DATAPATH__abc_16259_n6914;
  wire AES_CORE_DATAPATH__abc_16259_n6915;
  wire AES_CORE_DATAPATH__abc_16259_n6916;
  wire AES_CORE_DATAPATH__abc_16259_n6917;
  wire AES_CORE_DATAPATH__abc_16259_n6918;
  wire AES_CORE_DATAPATH__abc_16259_n6919;
  wire AES_CORE_DATAPATH__abc_16259_n6920;
  wire AES_CORE_DATAPATH__abc_16259_n6921;
  wire AES_CORE_DATAPATH__abc_16259_n6922;
  wire AES_CORE_DATAPATH__abc_16259_n6924;
  wire AES_CORE_DATAPATH__abc_16259_n6925;
  wire AES_CORE_DATAPATH__abc_16259_n6926;
  wire AES_CORE_DATAPATH__abc_16259_n6927;
  wire AES_CORE_DATAPATH__abc_16259_n6928;
  wire AES_CORE_DATAPATH__abc_16259_n6929;
  wire AES_CORE_DATAPATH__abc_16259_n6930;
  wire AES_CORE_DATAPATH__abc_16259_n6931;
  wire AES_CORE_DATAPATH__abc_16259_n6932;
  wire AES_CORE_DATAPATH__abc_16259_n6933;
  wire AES_CORE_DATAPATH__abc_16259_n6934;
  wire AES_CORE_DATAPATH__abc_16259_n6935;
  wire AES_CORE_DATAPATH__abc_16259_n6936;
  wire AES_CORE_DATAPATH__abc_16259_n6937;
  wire AES_CORE_DATAPATH__abc_16259_n6938;
  wire AES_CORE_DATAPATH__abc_16259_n6939;
  wire AES_CORE_DATAPATH__abc_16259_n6940;
  wire AES_CORE_DATAPATH__abc_16259_n6941;
  wire AES_CORE_DATAPATH__abc_16259_n6942;
  wire AES_CORE_DATAPATH__abc_16259_n6943;
  wire AES_CORE_DATAPATH__abc_16259_n6944;
  wire AES_CORE_DATAPATH__abc_16259_n6945;
  wire AES_CORE_DATAPATH__abc_16259_n6946;
  wire AES_CORE_DATAPATH__abc_16259_n6947;
  wire AES_CORE_DATAPATH__abc_16259_n6948;
  wire AES_CORE_DATAPATH__abc_16259_n6949;
  wire AES_CORE_DATAPATH__abc_16259_n6950;
  wire AES_CORE_DATAPATH__abc_16259_n6951;
  wire AES_CORE_DATAPATH__abc_16259_n6952;
  wire AES_CORE_DATAPATH__abc_16259_n6953;
  wire AES_CORE_DATAPATH__abc_16259_n6954;
  wire AES_CORE_DATAPATH__abc_16259_n6955;
  wire AES_CORE_DATAPATH__abc_16259_n6956;
  wire AES_CORE_DATAPATH__abc_16259_n6957;
  wire AES_CORE_DATAPATH__abc_16259_n6958;
  wire AES_CORE_DATAPATH__abc_16259_n6959;
  wire AES_CORE_DATAPATH__abc_16259_n6960;
  wire AES_CORE_DATAPATH__abc_16259_n6961;
  wire AES_CORE_DATAPATH__abc_16259_n6962;
  wire AES_CORE_DATAPATH__abc_16259_n6963;
  wire AES_CORE_DATAPATH__abc_16259_n6964;
  wire AES_CORE_DATAPATH__abc_16259_n6965;
  wire AES_CORE_DATAPATH__abc_16259_n6966;
  wire AES_CORE_DATAPATH__abc_16259_n6967;
  wire AES_CORE_DATAPATH__abc_16259_n6968;
  wire AES_CORE_DATAPATH__abc_16259_n6969;
  wire AES_CORE_DATAPATH__abc_16259_n6970;
  wire AES_CORE_DATAPATH__abc_16259_n6971;
  wire AES_CORE_DATAPATH__abc_16259_n6972;
  wire AES_CORE_DATAPATH__abc_16259_n6973;
  wire AES_CORE_DATAPATH__abc_16259_n6974;
  wire AES_CORE_DATAPATH__abc_16259_n6975;
  wire AES_CORE_DATAPATH__abc_16259_n6976;
  wire AES_CORE_DATAPATH__abc_16259_n6978;
  wire AES_CORE_DATAPATH__abc_16259_n6979;
  wire AES_CORE_DATAPATH__abc_16259_n6980;
  wire AES_CORE_DATAPATH__abc_16259_n6981;
  wire AES_CORE_DATAPATH__abc_16259_n6982;
  wire AES_CORE_DATAPATH__abc_16259_n6983;
  wire AES_CORE_DATAPATH__abc_16259_n6984;
  wire AES_CORE_DATAPATH__abc_16259_n6985;
  wire AES_CORE_DATAPATH__abc_16259_n6986;
  wire AES_CORE_DATAPATH__abc_16259_n6987;
  wire AES_CORE_DATAPATH__abc_16259_n6988;
  wire AES_CORE_DATAPATH__abc_16259_n6989;
  wire AES_CORE_DATAPATH__abc_16259_n6990;
  wire AES_CORE_DATAPATH__abc_16259_n6991;
  wire AES_CORE_DATAPATH__abc_16259_n6992;
  wire AES_CORE_DATAPATH__abc_16259_n6993;
  wire AES_CORE_DATAPATH__abc_16259_n6994;
  wire AES_CORE_DATAPATH__abc_16259_n6995;
  wire AES_CORE_DATAPATH__abc_16259_n6996;
  wire AES_CORE_DATAPATH__abc_16259_n6997;
  wire AES_CORE_DATAPATH__abc_16259_n6998;
  wire AES_CORE_DATAPATH__abc_16259_n6999;
  wire AES_CORE_DATAPATH__abc_16259_n7000;
  wire AES_CORE_DATAPATH__abc_16259_n7001;
  wire AES_CORE_DATAPATH__abc_16259_n7002;
  wire AES_CORE_DATAPATH__abc_16259_n7003;
  wire AES_CORE_DATAPATH__abc_16259_n7004;
  wire AES_CORE_DATAPATH__abc_16259_n7005;
  wire AES_CORE_DATAPATH__abc_16259_n7006;
  wire AES_CORE_DATAPATH__abc_16259_n7007;
  wire AES_CORE_DATAPATH__abc_16259_n7008;
  wire AES_CORE_DATAPATH__abc_16259_n7009;
  wire AES_CORE_DATAPATH__abc_16259_n7010;
  wire AES_CORE_DATAPATH__abc_16259_n7011;
  wire AES_CORE_DATAPATH__abc_16259_n7012;
  wire AES_CORE_DATAPATH__abc_16259_n7013;
  wire AES_CORE_DATAPATH__abc_16259_n7014;
  wire AES_CORE_DATAPATH__abc_16259_n7015;
  wire AES_CORE_DATAPATH__abc_16259_n7016;
  wire AES_CORE_DATAPATH__abc_16259_n7017;
  wire AES_CORE_DATAPATH__abc_16259_n7018;
  wire AES_CORE_DATAPATH__abc_16259_n7019;
  wire AES_CORE_DATAPATH__abc_16259_n7020;
  wire AES_CORE_DATAPATH__abc_16259_n7021;
  wire AES_CORE_DATAPATH__abc_16259_n7022;
  wire AES_CORE_DATAPATH__abc_16259_n7023;
  wire AES_CORE_DATAPATH__abc_16259_n7024;
  wire AES_CORE_DATAPATH__abc_16259_n7025;
  wire AES_CORE_DATAPATH__abc_16259_n7027;
  wire AES_CORE_DATAPATH__abc_16259_n7028;
  wire AES_CORE_DATAPATH__abc_16259_n7029;
  wire AES_CORE_DATAPATH__abc_16259_n7030;
  wire AES_CORE_DATAPATH__abc_16259_n7031;
  wire AES_CORE_DATAPATH__abc_16259_n7032;
  wire AES_CORE_DATAPATH__abc_16259_n7033;
  wire AES_CORE_DATAPATH__abc_16259_n7034;
  wire AES_CORE_DATAPATH__abc_16259_n7035;
  wire AES_CORE_DATAPATH__abc_16259_n7036;
  wire AES_CORE_DATAPATH__abc_16259_n7037;
  wire AES_CORE_DATAPATH__abc_16259_n7038;
  wire AES_CORE_DATAPATH__abc_16259_n7039;
  wire AES_CORE_DATAPATH__abc_16259_n7040;
  wire AES_CORE_DATAPATH__abc_16259_n7041;
  wire AES_CORE_DATAPATH__abc_16259_n7042;
  wire AES_CORE_DATAPATH__abc_16259_n7043;
  wire AES_CORE_DATAPATH__abc_16259_n7044;
  wire AES_CORE_DATAPATH__abc_16259_n7045;
  wire AES_CORE_DATAPATH__abc_16259_n7046;
  wire AES_CORE_DATAPATH__abc_16259_n7047;
  wire AES_CORE_DATAPATH__abc_16259_n7048;
  wire AES_CORE_DATAPATH__abc_16259_n7049;
  wire AES_CORE_DATAPATH__abc_16259_n7050;
  wire AES_CORE_DATAPATH__abc_16259_n7051;
  wire AES_CORE_DATAPATH__abc_16259_n7052;
  wire AES_CORE_DATAPATH__abc_16259_n7053;
  wire AES_CORE_DATAPATH__abc_16259_n7054;
  wire AES_CORE_DATAPATH__abc_16259_n7055;
  wire AES_CORE_DATAPATH__abc_16259_n7056;
  wire AES_CORE_DATAPATH__abc_16259_n7057;
  wire AES_CORE_DATAPATH__abc_16259_n7058;
  wire AES_CORE_DATAPATH__abc_16259_n7059;
  wire AES_CORE_DATAPATH__abc_16259_n7060;
  wire AES_CORE_DATAPATH__abc_16259_n7061;
  wire AES_CORE_DATAPATH__abc_16259_n7062;
  wire AES_CORE_DATAPATH__abc_16259_n7063;
  wire AES_CORE_DATAPATH__abc_16259_n7064;
  wire AES_CORE_DATAPATH__abc_16259_n7065;
  wire AES_CORE_DATAPATH__abc_16259_n7066;
  wire AES_CORE_DATAPATH__abc_16259_n7067;
  wire AES_CORE_DATAPATH__abc_16259_n7068;
  wire AES_CORE_DATAPATH__abc_16259_n7069;
  wire AES_CORE_DATAPATH__abc_16259_n7070;
  wire AES_CORE_DATAPATH__abc_16259_n7071;
  wire AES_CORE_DATAPATH__abc_16259_n7072;
  wire AES_CORE_DATAPATH__abc_16259_n7073;
  wire AES_CORE_DATAPATH__abc_16259_n7074;
  wire AES_CORE_DATAPATH__abc_16259_n7076;
  wire AES_CORE_DATAPATH__abc_16259_n7077;
  wire AES_CORE_DATAPATH__abc_16259_n7078;
  wire AES_CORE_DATAPATH__abc_16259_n7079;
  wire AES_CORE_DATAPATH__abc_16259_n7080;
  wire AES_CORE_DATAPATH__abc_16259_n7081;
  wire AES_CORE_DATAPATH__abc_16259_n7082;
  wire AES_CORE_DATAPATH__abc_16259_n7083;
  wire AES_CORE_DATAPATH__abc_16259_n7084;
  wire AES_CORE_DATAPATH__abc_16259_n7085;
  wire AES_CORE_DATAPATH__abc_16259_n7086;
  wire AES_CORE_DATAPATH__abc_16259_n7087;
  wire AES_CORE_DATAPATH__abc_16259_n7088;
  wire AES_CORE_DATAPATH__abc_16259_n7089;
  wire AES_CORE_DATAPATH__abc_16259_n7090;
  wire AES_CORE_DATAPATH__abc_16259_n7091;
  wire AES_CORE_DATAPATH__abc_16259_n7092;
  wire AES_CORE_DATAPATH__abc_16259_n7093;
  wire AES_CORE_DATAPATH__abc_16259_n7094;
  wire AES_CORE_DATAPATH__abc_16259_n7095;
  wire AES_CORE_DATAPATH__abc_16259_n7096;
  wire AES_CORE_DATAPATH__abc_16259_n7097;
  wire AES_CORE_DATAPATH__abc_16259_n7098;
  wire AES_CORE_DATAPATH__abc_16259_n7099;
  wire AES_CORE_DATAPATH__abc_16259_n7100;
  wire AES_CORE_DATAPATH__abc_16259_n7101;
  wire AES_CORE_DATAPATH__abc_16259_n7102;
  wire AES_CORE_DATAPATH__abc_16259_n7103;
  wire AES_CORE_DATAPATH__abc_16259_n7104;
  wire AES_CORE_DATAPATH__abc_16259_n7105;
  wire AES_CORE_DATAPATH__abc_16259_n7106;
  wire AES_CORE_DATAPATH__abc_16259_n7107;
  wire AES_CORE_DATAPATH__abc_16259_n7108;
  wire AES_CORE_DATAPATH__abc_16259_n7109;
  wire AES_CORE_DATAPATH__abc_16259_n7110;
  wire AES_CORE_DATAPATH__abc_16259_n7111;
  wire AES_CORE_DATAPATH__abc_16259_n7112;
  wire AES_CORE_DATAPATH__abc_16259_n7113;
  wire AES_CORE_DATAPATH__abc_16259_n7114;
  wire AES_CORE_DATAPATH__abc_16259_n7115;
  wire AES_CORE_DATAPATH__abc_16259_n7116;
  wire AES_CORE_DATAPATH__abc_16259_n7117;
  wire AES_CORE_DATAPATH__abc_16259_n7118;
  wire AES_CORE_DATAPATH__abc_16259_n7119;
  wire AES_CORE_DATAPATH__abc_16259_n7120;
  wire AES_CORE_DATAPATH__abc_16259_n7121;
  wire AES_CORE_DATAPATH__abc_16259_n7122;
  wire AES_CORE_DATAPATH__abc_16259_n7123;
  wire AES_CORE_DATAPATH__abc_16259_n7125;
  wire AES_CORE_DATAPATH__abc_16259_n7126;
  wire AES_CORE_DATAPATH__abc_16259_n7127;
  wire AES_CORE_DATAPATH__abc_16259_n7128;
  wire AES_CORE_DATAPATH__abc_16259_n7129;
  wire AES_CORE_DATAPATH__abc_16259_n7130;
  wire AES_CORE_DATAPATH__abc_16259_n7131;
  wire AES_CORE_DATAPATH__abc_16259_n7132;
  wire AES_CORE_DATAPATH__abc_16259_n7133;
  wire AES_CORE_DATAPATH__abc_16259_n7134;
  wire AES_CORE_DATAPATH__abc_16259_n7135;
  wire AES_CORE_DATAPATH__abc_16259_n7136;
  wire AES_CORE_DATAPATH__abc_16259_n7137;
  wire AES_CORE_DATAPATH__abc_16259_n7138;
  wire AES_CORE_DATAPATH__abc_16259_n7139;
  wire AES_CORE_DATAPATH__abc_16259_n7140;
  wire AES_CORE_DATAPATH__abc_16259_n7141;
  wire AES_CORE_DATAPATH__abc_16259_n7142;
  wire AES_CORE_DATAPATH__abc_16259_n7143;
  wire AES_CORE_DATAPATH__abc_16259_n7144;
  wire AES_CORE_DATAPATH__abc_16259_n7145;
  wire AES_CORE_DATAPATH__abc_16259_n7146;
  wire AES_CORE_DATAPATH__abc_16259_n7147;
  wire AES_CORE_DATAPATH__abc_16259_n7148;
  wire AES_CORE_DATAPATH__abc_16259_n7149;
  wire AES_CORE_DATAPATH__abc_16259_n7150;
  wire AES_CORE_DATAPATH__abc_16259_n7151;
  wire AES_CORE_DATAPATH__abc_16259_n7152;
  wire AES_CORE_DATAPATH__abc_16259_n7153;
  wire AES_CORE_DATAPATH__abc_16259_n7154;
  wire AES_CORE_DATAPATH__abc_16259_n7155;
  wire AES_CORE_DATAPATH__abc_16259_n7156;
  wire AES_CORE_DATAPATH__abc_16259_n7157;
  wire AES_CORE_DATAPATH__abc_16259_n7158;
  wire AES_CORE_DATAPATH__abc_16259_n7159;
  wire AES_CORE_DATAPATH__abc_16259_n7160;
  wire AES_CORE_DATAPATH__abc_16259_n7161;
  wire AES_CORE_DATAPATH__abc_16259_n7162;
  wire AES_CORE_DATAPATH__abc_16259_n7163;
  wire AES_CORE_DATAPATH__abc_16259_n7164;
  wire AES_CORE_DATAPATH__abc_16259_n7165;
  wire AES_CORE_DATAPATH__abc_16259_n7166;
  wire AES_CORE_DATAPATH__abc_16259_n7167;
  wire AES_CORE_DATAPATH__abc_16259_n7168;
  wire AES_CORE_DATAPATH__abc_16259_n7169;
  wire AES_CORE_DATAPATH__abc_16259_n7170;
  wire AES_CORE_DATAPATH__abc_16259_n7171;
  wire AES_CORE_DATAPATH__abc_16259_n7172;
  wire AES_CORE_DATAPATH__abc_16259_n7173;
  wire AES_CORE_DATAPATH__abc_16259_n7174;
  wire AES_CORE_DATAPATH__abc_16259_n7175;
  wire AES_CORE_DATAPATH__abc_16259_n7176;
  wire AES_CORE_DATAPATH__abc_16259_n7177;
  wire AES_CORE_DATAPATH__abc_16259_n7179;
  wire AES_CORE_DATAPATH__abc_16259_n7180;
  wire AES_CORE_DATAPATH__abc_16259_n7181;
  wire AES_CORE_DATAPATH__abc_16259_n7182;
  wire AES_CORE_DATAPATH__abc_16259_n7183;
  wire AES_CORE_DATAPATH__abc_16259_n7184;
  wire AES_CORE_DATAPATH__abc_16259_n7185;
  wire AES_CORE_DATAPATH__abc_16259_n7186;
  wire AES_CORE_DATAPATH__abc_16259_n7187;
  wire AES_CORE_DATAPATH__abc_16259_n7188;
  wire AES_CORE_DATAPATH__abc_16259_n7189;
  wire AES_CORE_DATAPATH__abc_16259_n7190;
  wire AES_CORE_DATAPATH__abc_16259_n7191;
  wire AES_CORE_DATAPATH__abc_16259_n7192;
  wire AES_CORE_DATAPATH__abc_16259_n7193;
  wire AES_CORE_DATAPATH__abc_16259_n7194;
  wire AES_CORE_DATAPATH__abc_16259_n7195;
  wire AES_CORE_DATAPATH__abc_16259_n7196;
  wire AES_CORE_DATAPATH__abc_16259_n7197;
  wire AES_CORE_DATAPATH__abc_16259_n7198;
  wire AES_CORE_DATAPATH__abc_16259_n7199;
  wire AES_CORE_DATAPATH__abc_16259_n7200;
  wire AES_CORE_DATAPATH__abc_16259_n7201;
  wire AES_CORE_DATAPATH__abc_16259_n7202;
  wire AES_CORE_DATAPATH__abc_16259_n7203;
  wire AES_CORE_DATAPATH__abc_16259_n7204;
  wire AES_CORE_DATAPATH__abc_16259_n7205;
  wire AES_CORE_DATAPATH__abc_16259_n7206;
  wire AES_CORE_DATAPATH__abc_16259_n7207;
  wire AES_CORE_DATAPATH__abc_16259_n7208;
  wire AES_CORE_DATAPATH__abc_16259_n7209;
  wire AES_CORE_DATAPATH__abc_16259_n7210;
  wire AES_CORE_DATAPATH__abc_16259_n7211;
  wire AES_CORE_DATAPATH__abc_16259_n7212;
  wire AES_CORE_DATAPATH__abc_16259_n7213;
  wire AES_CORE_DATAPATH__abc_16259_n7214;
  wire AES_CORE_DATAPATH__abc_16259_n7215;
  wire AES_CORE_DATAPATH__abc_16259_n7216;
  wire AES_CORE_DATAPATH__abc_16259_n7217;
  wire AES_CORE_DATAPATH__abc_16259_n7218;
  wire AES_CORE_DATAPATH__abc_16259_n7219;
  wire AES_CORE_DATAPATH__abc_16259_n7220;
  wire AES_CORE_DATAPATH__abc_16259_n7221;
  wire AES_CORE_DATAPATH__abc_16259_n7222;
  wire AES_CORE_DATAPATH__abc_16259_n7223;
  wire AES_CORE_DATAPATH__abc_16259_n7224;
  wire AES_CORE_DATAPATH__abc_16259_n7225;
  wire AES_CORE_DATAPATH__abc_16259_n7226;
  wire AES_CORE_DATAPATH__abc_16259_n7228;
  wire AES_CORE_DATAPATH__abc_16259_n7229;
  wire AES_CORE_DATAPATH__abc_16259_n7230;
  wire AES_CORE_DATAPATH__abc_16259_n7231;
  wire AES_CORE_DATAPATH__abc_16259_n7232;
  wire AES_CORE_DATAPATH__abc_16259_n7233;
  wire AES_CORE_DATAPATH__abc_16259_n7234;
  wire AES_CORE_DATAPATH__abc_16259_n7235;
  wire AES_CORE_DATAPATH__abc_16259_n7236;
  wire AES_CORE_DATAPATH__abc_16259_n7237;
  wire AES_CORE_DATAPATH__abc_16259_n7238;
  wire AES_CORE_DATAPATH__abc_16259_n7239;
  wire AES_CORE_DATAPATH__abc_16259_n7240;
  wire AES_CORE_DATAPATH__abc_16259_n7241;
  wire AES_CORE_DATAPATH__abc_16259_n7242;
  wire AES_CORE_DATAPATH__abc_16259_n7243;
  wire AES_CORE_DATAPATH__abc_16259_n7244;
  wire AES_CORE_DATAPATH__abc_16259_n7245;
  wire AES_CORE_DATAPATH__abc_16259_n7246;
  wire AES_CORE_DATAPATH__abc_16259_n7247;
  wire AES_CORE_DATAPATH__abc_16259_n7248;
  wire AES_CORE_DATAPATH__abc_16259_n7249;
  wire AES_CORE_DATAPATH__abc_16259_n7250;
  wire AES_CORE_DATAPATH__abc_16259_n7251;
  wire AES_CORE_DATAPATH__abc_16259_n7252;
  wire AES_CORE_DATAPATH__abc_16259_n7253;
  wire AES_CORE_DATAPATH__abc_16259_n7254;
  wire AES_CORE_DATAPATH__abc_16259_n7255;
  wire AES_CORE_DATAPATH__abc_16259_n7256;
  wire AES_CORE_DATAPATH__abc_16259_n7257;
  wire AES_CORE_DATAPATH__abc_16259_n7258;
  wire AES_CORE_DATAPATH__abc_16259_n7259;
  wire AES_CORE_DATAPATH__abc_16259_n7260;
  wire AES_CORE_DATAPATH__abc_16259_n7261;
  wire AES_CORE_DATAPATH__abc_16259_n7262;
  wire AES_CORE_DATAPATH__abc_16259_n7263;
  wire AES_CORE_DATAPATH__abc_16259_n7264;
  wire AES_CORE_DATAPATH__abc_16259_n7265;
  wire AES_CORE_DATAPATH__abc_16259_n7266;
  wire AES_CORE_DATAPATH__abc_16259_n7267;
  wire AES_CORE_DATAPATH__abc_16259_n7268;
  wire AES_CORE_DATAPATH__abc_16259_n7269;
  wire AES_CORE_DATAPATH__abc_16259_n7270;
  wire AES_CORE_DATAPATH__abc_16259_n7271;
  wire AES_CORE_DATAPATH__abc_16259_n7272;
  wire AES_CORE_DATAPATH__abc_16259_n7273;
  wire AES_CORE_DATAPATH__abc_16259_n7274;
  wire AES_CORE_DATAPATH__abc_16259_n7275;
  wire AES_CORE_DATAPATH__abc_16259_n7277;
  wire AES_CORE_DATAPATH__abc_16259_n7278;
  wire AES_CORE_DATAPATH__abc_16259_n7279;
  wire AES_CORE_DATAPATH__abc_16259_n7280;
  wire AES_CORE_DATAPATH__abc_16259_n7281;
  wire AES_CORE_DATAPATH__abc_16259_n7282;
  wire AES_CORE_DATAPATH__abc_16259_n7283;
  wire AES_CORE_DATAPATH__abc_16259_n7284;
  wire AES_CORE_DATAPATH__abc_16259_n7285;
  wire AES_CORE_DATAPATH__abc_16259_n7286;
  wire AES_CORE_DATAPATH__abc_16259_n7287;
  wire AES_CORE_DATAPATH__abc_16259_n7288;
  wire AES_CORE_DATAPATH__abc_16259_n7289;
  wire AES_CORE_DATAPATH__abc_16259_n7290;
  wire AES_CORE_DATAPATH__abc_16259_n7291;
  wire AES_CORE_DATAPATH__abc_16259_n7292;
  wire AES_CORE_DATAPATH__abc_16259_n7293;
  wire AES_CORE_DATAPATH__abc_16259_n7294;
  wire AES_CORE_DATAPATH__abc_16259_n7295;
  wire AES_CORE_DATAPATH__abc_16259_n7296;
  wire AES_CORE_DATAPATH__abc_16259_n7297;
  wire AES_CORE_DATAPATH__abc_16259_n7298;
  wire AES_CORE_DATAPATH__abc_16259_n7299;
  wire AES_CORE_DATAPATH__abc_16259_n7300;
  wire AES_CORE_DATAPATH__abc_16259_n7301;
  wire AES_CORE_DATAPATH__abc_16259_n7302;
  wire AES_CORE_DATAPATH__abc_16259_n7303;
  wire AES_CORE_DATAPATH__abc_16259_n7304;
  wire AES_CORE_DATAPATH__abc_16259_n7305;
  wire AES_CORE_DATAPATH__abc_16259_n7306;
  wire AES_CORE_DATAPATH__abc_16259_n7307;
  wire AES_CORE_DATAPATH__abc_16259_n7308;
  wire AES_CORE_DATAPATH__abc_16259_n7309;
  wire AES_CORE_DATAPATH__abc_16259_n7310;
  wire AES_CORE_DATAPATH__abc_16259_n7311;
  wire AES_CORE_DATAPATH__abc_16259_n7312;
  wire AES_CORE_DATAPATH__abc_16259_n7313;
  wire AES_CORE_DATAPATH__abc_16259_n7314;
  wire AES_CORE_DATAPATH__abc_16259_n7315;
  wire AES_CORE_DATAPATH__abc_16259_n7316;
  wire AES_CORE_DATAPATH__abc_16259_n7317;
  wire AES_CORE_DATAPATH__abc_16259_n7318;
  wire AES_CORE_DATAPATH__abc_16259_n7319;
  wire AES_CORE_DATAPATH__abc_16259_n7320;
  wire AES_CORE_DATAPATH__abc_16259_n7321;
  wire AES_CORE_DATAPATH__abc_16259_n7322;
  wire AES_CORE_DATAPATH__abc_16259_n7323;
  wire AES_CORE_DATAPATH__abc_16259_n7324;
  wire AES_CORE_DATAPATH__abc_16259_n7326;
  wire AES_CORE_DATAPATH__abc_16259_n7327;
  wire AES_CORE_DATAPATH__abc_16259_n7328;
  wire AES_CORE_DATAPATH__abc_16259_n7329;
  wire AES_CORE_DATAPATH__abc_16259_n7330;
  wire AES_CORE_DATAPATH__abc_16259_n7331;
  wire AES_CORE_DATAPATH__abc_16259_n7332;
  wire AES_CORE_DATAPATH__abc_16259_n7333;
  wire AES_CORE_DATAPATH__abc_16259_n7334;
  wire AES_CORE_DATAPATH__abc_16259_n7335;
  wire AES_CORE_DATAPATH__abc_16259_n7336;
  wire AES_CORE_DATAPATH__abc_16259_n7337;
  wire AES_CORE_DATAPATH__abc_16259_n7338;
  wire AES_CORE_DATAPATH__abc_16259_n7339;
  wire AES_CORE_DATAPATH__abc_16259_n7340;
  wire AES_CORE_DATAPATH__abc_16259_n7341;
  wire AES_CORE_DATAPATH__abc_16259_n7342;
  wire AES_CORE_DATAPATH__abc_16259_n7343;
  wire AES_CORE_DATAPATH__abc_16259_n7344;
  wire AES_CORE_DATAPATH__abc_16259_n7345;
  wire AES_CORE_DATAPATH__abc_16259_n7346;
  wire AES_CORE_DATAPATH__abc_16259_n7347;
  wire AES_CORE_DATAPATH__abc_16259_n7348;
  wire AES_CORE_DATAPATH__abc_16259_n7349;
  wire AES_CORE_DATAPATH__abc_16259_n7350;
  wire AES_CORE_DATAPATH__abc_16259_n7351;
  wire AES_CORE_DATAPATH__abc_16259_n7352;
  wire AES_CORE_DATAPATH__abc_16259_n7353;
  wire AES_CORE_DATAPATH__abc_16259_n7354;
  wire AES_CORE_DATAPATH__abc_16259_n7355;
  wire AES_CORE_DATAPATH__abc_16259_n7356;
  wire AES_CORE_DATAPATH__abc_16259_n7357;
  wire AES_CORE_DATAPATH__abc_16259_n7358;
  wire AES_CORE_DATAPATH__abc_16259_n7359;
  wire AES_CORE_DATAPATH__abc_16259_n7360;
  wire AES_CORE_DATAPATH__abc_16259_n7361;
  wire AES_CORE_DATAPATH__abc_16259_n7362;
  wire AES_CORE_DATAPATH__abc_16259_n7363;
  wire AES_CORE_DATAPATH__abc_16259_n7364;
  wire AES_CORE_DATAPATH__abc_16259_n7365;
  wire AES_CORE_DATAPATH__abc_16259_n7366;
  wire AES_CORE_DATAPATH__abc_16259_n7367;
  wire AES_CORE_DATAPATH__abc_16259_n7368;
  wire AES_CORE_DATAPATH__abc_16259_n7369;
  wire AES_CORE_DATAPATH__abc_16259_n7370;
  wire AES_CORE_DATAPATH__abc_16259_n7371;
  wire AES_CORE_DATAPATH__abc_16259_n7372;
  wire AES_CORE_DATAPATH__abc_16259_n7373;
  wire AES_CORE_DATAPATH__abc_16259_n7375;
  wire AES_CORE_DATAPATH__abc_16259_n7376;
  wire AES_CORE_DATAPATH__abc_16259_n7377;
  wire AES_CORE_DATAPATH__abc_16259_n7378;
  wire AES_CORE_DATAPATH__abc_16259_n7379;
  wire AES_CORE_DATAPATH__abc_16259_n7380;
  wire AES_CORE_DATAPATH__abc_16259_n7381;
  wire AES_CORE_DATAPATH__abc_16259_n7382;
  wire AES_CORE_DATAPATH__abc_16259_n7383;
  wire AES_CORE_DATAPATH__abc_16259_n7384;
  wire AES_CORE_DATAPATH__abc_16259_n7385;
  wire AES_CORE_DATAPATH__abc_16259_n7386;
  wire AES_CORE_DATAPATH__abc_16259_n7387;
  wire AES_CORE_DATAPATH__abc_16259_n7388;
  wire AES_CORE_DATAPATH__abc_16259_n7389;
  wire AES_CORE_DATAPATH__abc_16259_n7390;
  wire AES_CORE_DATAPATH__abc_16259_n7391;
  wire AES_CORE_DATAPATH__abc_16259_n7392;
  wire AES_CORE_DATAPATH__abc_16259_n7393;
  wire AES_CORE_DATAPATH__abc_16259_n7394;
  wire AES_CORE_DATAPATH__abc_16259_n7395;
  wire AES_CORE_DATAPATH__abc_16259_n7396;
  wire AES_CORE_DATAPATH__abc_16259_n7397;
  wire AES_CORE_DATAPATH__abc_16259_n7398;
  wire AES_CORE_DATAPATH__abc_16259_n7399;
  wire AES_CORE_DATAPATH__abc_16259_n7400;
  wire AES_CORE_DATAPATH__abc_16259_n7401;
  wire AES_CORE_DATAPATH__abc_16259_n7402;
  wire AES_CORE_DATAPATH__abc_16259_n7403;
  wire AES_CORE_DATAPATH__abc_16259_n7404;
  wire AES_CORE_DATAPATH__abc_16259_n7405;
  wire AES_CORE_DATAPATH__abc_16259_n7406;
  wire AES_CORE_DATAPATH__abc_16259_n7407;
  wire AES_CORE_DATAPATH__abc_16259_n7408;
  wire AES_CORE_DATAPATH__abc_16259_n7409;
  wire AES_CORE_DATAPATH__abc_16259_n7410;
  wire AES_CORE_DATAPATH__abc_16259_n7411;
  wire AES_CORE_DATAPATH__abc_16259_n7412;
  wire AES_CORE_DATAPATH__abc_16259_n7413;
  wire AES_CORE_DATAPATH__abc_16259_n7414;
  wire AES_CORE_DATAPATH__abc_16259_n7415;
  wire AES_CORE_DATAPATH__abc_16259_n7416;
  wire AES_CORE_DATAPATH__abc_16259_n7417;
  wire AES_CORE_DATAPATH__abc_16259_n7418;
  wire AES_CORE_DATAPATH__abc_16259_n7419;
  wire AES_CORE_DATAPATH__abc_16259_n7420;
  wire AES_CORE_DATAPATH__abc_16259_n7421;
  wire AES_CORE_DATAPATH__abc_16259_n7422;
  wire AES_CORE_DATAPATH__abc_16259_n7424;
  wire AES_CORE_DATAPATH__abc_16259_n7425;
  wire AES_CORE_DATAPATH__abc_16259_n7426;
  wire AES_CORE_DATAPATH__abc_16259_n7427;
  wire AES_CORE_DATAPATH__abc_16259_n7428;
  wire AES_CORE_DATAPATH__abc_16259_n7429;
  wire AES_CORE_DATAPATH__abc_16259_n7430;
  wire AES_CORE_DATAPATH__abc_16259_n7431;
  wire AES_CORE_DATAPATH__abc_16259_n7432;
  wire AES_CORE_DATAPATH__abc_16259_n7433;
  wire AES_CORE_DATAPATH__abc_16259_n7434;
  wire AES_CORE_DATAPATH__abc_16259_n7435;
  wire AES_CORE_DATAPATH__abc_16259_n7436;
  wire AES_CORE_DATAPATH__abc_16259_n7437;
  wire AES_CORE_DATAPATH__abc_16259_n7438;
  wire AES_CORE_DATAPATH__abc_16259_n7439;
  wire AES_CORE_DATAPATH__abc_16259_n7440;
  wire AES_CORE_DATAPATH__abc_16259_n7441;
  wire AES_CORE_DATAPATH__abc_16259_n7442;
  wire AES_CORE_DATAPATH__abc_16259_n7443;
  wire AES_CORE_DATAPATH__abc_16259_n7444;
  wire AES_CORE_DATAPATH__abc_16259_n7445;
  wire AES_CORE_DATAPATH__abc_16259_n7446;
  wire AES_CORE_DATAPATH__abc_16259_n7447;
  wire AES_CORE_DATAPATH__abc_16259_n7448;
  wire AES_CORE_DATAPATH__abc_16259_n7449;
  wire AES_CORE_DATAPATH__abc_16259_n7450;
  wire AES_CORE_DATAPATH__abc_16259_n7451;
  wire AES_CORE_DATAPATH__abc_16259_n7452;
  wire AES_CORE_DATAPATH__abc_16259_n7453;
  wire AES_CORE_DATAPATH__abc_16259_n7454;
  wire AES_CORE_DATAPATH__abc_16259_n7455;
  wire AES_CORE_DATAPATH__abc_16259_n7456;
  wire AES_CORE_DATAPATH__abc_16259_n7457;
  wire AES_CORE_DATAPATH__abc_16259_n7458;
  wire AES_CORE_DATAPATH__abc_16259_n7459;
  wire AES_CORE_DATAPATH__abc_16259_n7460;
  wire AES_CORE_DATAPATH__abc_16259_n7461;
  wire AES_CORE_DATAPATH__abc_16259_n7462;
  wire AES_CORE_DATAPATH__abc_16259_n7463;
  wire AES_CORE_DATAPATH__abc_16259_n7464;
  wire AES_CORE_DATAPATH__abc_16259_n7465;
  wire AES_CORE_DATAPATH__abc_16259_n7466;
  wire AES_CORE_DATAPATH__abc_16259_n7467;
  wire AES_CORE_DATAPATH__abc_16259_n7468;
  wire AES_CORE_DATAPATH__abc_16259_n7469;
  wire AES_CORE_DATAPATH__abc_16259_n7470;
  wire AES_CORE_DATAPATH__abc_16259_n7471;
  wire AES_CORE_DATAPATH__abc_16259_n7473;
  wire AES_CORE_DATAPATH__abc_16259_n7474;
  wire AES_CORE_DATAPATH__abc_16259_n7475;
  wire AES_CORE_DATAPATH__abc_16259_n7476;
  wire AES_CORE_DATAPATH__abc_16259_n7477;
  wire AES_CORE_DATAPATH__abc_16259_n7478;
  wire AES_CORE_DATAPATH__abc_16259_n7479;
  wire AES_CORE_DATAPATH__abc_16259_n7480;
  wire AES_CORE_DATAPATH__abc_16259_n7481;
  wire AES_CORE_DATAPATH__abc_16259_n7482;
  wire AES_CORE_DATAPATH__abc_16259_n7483;
  wire AES_CORE_DATAPATH__abc_16259_n7484;
  wire AES_CORE_DATAPATH__abc_16259_n7485;
  wire AES_CORE_DATAPATH__abc_16259_n7486;
  wire AES_CORE_DATAPATH__abc_16259_n7487;
  wire AES_CORE_DATAPATH__abc_16259_n7488;
  wire AES_CORE_DATAPATH__abc_16259_n7489;
  wire AES_CORE_DATAPATH__abc_16259_n7490;
  wire AES_CORE_DATAPATH__abc_16259_n7491;
  wire AES_CORE_DATAPATH__abc_16259_n7492;
  wire AES_CORE_DATAPATH__abc_16259_n7493;
  wire AES_CORE_DATAPATH__abc_16259_n7494;
  wire AES_CORE_DATAPATH__abc_16259_n7495;
  wire AES_CORE_DATAPATH__abc_16259_n7496;
  wire AES_CORE_DATAPATH__abc_16259_n7497;
  wire AES_CORE_DATAPATH__abc_16259_n7498;
  wire AES_CORE_DATAPATH__abc_16259_n7499;
  wire AES_CORE_DATAPATH__abc_16259_n7500;
  wire AES_CORE_DATAPATH__abc_16259_n7501;
  wire AES_CORE_DATAPATH__abc_16259_n7502;
  wire AES_CORE_DATAPATH__abc_16259_n7503;
  wire AES_CORE_DATAPATH__abc_16259_n7504;
  wire AES_CORE_DATAPATH__abc_16259_n7505;
  wire AES_CORE_DATAPATH__abc_16259_n7506;
  wire AES_CORE_DATAPATH__abc_16259_n7507;
  wire AES_CORE_DATAPATH__abc_16259_n7508;
  wire AES_CORE_DATAPATH__abc_16259_n7509;
  wire AES_CORE_DATAPATH__abc_16259_n7510;
  wire AES_CORE_DATAPATH__abc_16259_n7511;
  wire AES_CORE_DATAPATH__abc_16259_n7512;
  wire AES_CORE_DATAPATH__abc_16259_n7513;
  wire AES_CORE_DATAPATH__abc_16259_n7514;
  wire AES_CORE_DATAPATH__abc_16259_n7515;
  wire AES_CORE_DATAPATH__abc_16259_n7516;
  wire AES_CORE_DATAPATH__abc_16259_n7517;
  wire AES_CORE_DATAPATH__abc_16259_n7518;
  wire AES_CORE_DATAPATH__abc_16259_n7519;
  wire AES_CORE_DATAPATH__abc_16259_n7520;
  wire AES_CORE_DATAPATH__abc_16259_n7522;
  wire AES_CORE_DATAPATH__abc_16259_n7523;
  wire AES_CORE_DATAPATH__abc_16259_n7524;
  wire AES_CORE_DATAPATH__abc_16259_n7525;
  wire AES_CORE_DATAPATH__abc_16259_n7526;
  wire AES_CORE_DATAPATH__abc_16259_n7527;
  wire AES_CORE_DATAPATH__abc_16259_n7528;
  wire AES_CORE_DATAPATH__abc_16259_n7529;
  wire AES_CORE_DATAPATH__abc_16259_n7530;
  wire AES_CORE_DATAPATH__abc_16259_n7531;
  wire AES_CORE_DATAPATH__abc_16259_n7532;
  wire AES_CORE_DATAPATH__abc_16259_n7533;
  wire AES_CORE_DATAPATH__abc_16259_n7534;
  wire AES_CORE_DATAPATH__abc_16259_n7535;
  wire AES_CORE_DATAPATH__abc_16259_n7536;
  wire AES_CORE_DATAPATH__abc_16259_n7537;
  wire AES_CORE_DATAPATH__abc_16259_n7538;
  wire AES_CORE_DATAPATH__abc_16259_n7539;
  wire AES_CORE_DATAPATH__abc_16259_n7540;
  wire AES_CORE_DATAPATH__abc_16259_n7541;
  wire AES_CORE_DATAPATH__abc_16259_n7542;
  wire AES_CORE_DATAPATH__abc_16259_n7543;
  wire AES_CORE_DATAPATH__abc_16259_n7544;
  wire AES_CORE_DATAPATH__abc_16259_n7545;
  wire AES_CORE_DATAPATH__abc_16259_n7546;
  wire AES_CORE_DATAPATH__abc_16259_n7547;
  wire AES_CORE_DATAPATH__abc_16259_n7548;
  wire AES_CORE_DATAPATH__abc_16259_n7549;
  wire AES_CORE_DATAPATH__abc_16259_n7550;
  wire AES_CORE_DATAPATH__abc_16259_n7551;
  wire AES_CORE_DATAPATH__abc_16259_n7552;
  wire AES_CORE_DATAPATH__abc_16259_n7553;
  wire AES_CORE_DATAPATH__abc_16259_n7554;
  wire AES_CORE_DATAPATH__abc_16259_n7555;
  wire AES_CORE_DATAPATH__abc_16259_n7556;
  wire AES_CORE_DATAPATH__abc_16259_n7557;
  wire AES_CORE_DATAPATH__abc_16259_n7558;
  wire AES_CORE_DATAPATH__abc_16259_n7559;
  wire AES_CORE_DATAPATH__abc_16259_n7560;
  wire AES_CORE_DATAPATH__abc_16259_n7561;
  wire AES_CORE_DATAPATH__abc_16259_n7562;
  wire AES_CORE_DATAPATH__abc_16259_n7563;
  wire AES_CORE_DATAPATH__abc_16259_n7564;
  wire AES_CORE_DATAPATH__abc_16259_n7565;
  wire AES_CORE_DATAPATH__abc_16259_n7566;
  wire AES_CORE_DATAPATH__abc_16259_n7567;
  wire AES_CORE_DATAPATH__abc_16259_n7568;
  wire AES_CORE_DATAPATH__abc_16259_n7569;
  wire AES_CORE_DATAPATH__abc_16259_n7571;
  wire AES_CORE_DATAPATH__abc_16259_n7572;
  wire AES_CORE_DATAPATH__abc_16259_n7573;
  wire AES_CORE_DATAPATH__abc_16259_n7574;
  wire AES_CORE_DATAPATH__abc_16259_n7575;
  wire AES_CORE_DATAPATH__abc_16259_n7576;
  wire AES_CORE_DATAPATH__abc_16259_n7577;
  wire AES_CORE_DATAPATH__abc_16259_n7578;
  wire AES_CORE_DATAPATH__abc_16259_n7579;
  wire AES_CORE_DATAPATH__abc_16259_n7580;
  wire AES_CORE_DATAPATH__abc_16259_n7581;
  wire AES_CORE_DATAPATH__abc_16259_n7582;
  wire AES_CORE_DATAPATH__abc_16259_n7583;
  wire AES_CORE_DATAPATH__abc_16259_n7584;
  wire AES_CORE_DATAPATH__abc_16259_n7585;
  wire AES_CORE_DATAPATH__abc_16259_n7586;
  wire AES_CORE_DATAPATH__abc_16259_n7587;
  wire AES_CORE_DATAPATH__abc_16259_n7588;
  wire AES_CORE_DATAPATH__abc_16259_n7589;
  wire AES_CORE_DATAPATH__abc_16259_n7590;
  wire AES_CORE_DATAPATH__abc_16259_n7591;
  wire AES_CORE_DATAPATH__abc_16259_n7592;
  wire AES_CORE_DATAPATH__abc_16259_n7593;
  wire AES_CORE_DATAPATH__abc_16259_n7594;
  wire AES_CORE_DATAPATH__abc_16259_n7595;
  wire AES_CORE_DATAPATH__abc_16259_n7596;
  wire AES_CORE_DATAPATH__abc_16259_n7597;
  wire AES_CORE_DATAPATH__abc_16259_n7598;
  wire AES_CORE_DATAPATH__abc_16259_n7599;
  wire AES_CORE_DATAPATH__abc_16259_n7600;
  wire AES_CORE_DATAPATH__abc_16259_n7601;
  wire AES_CORE_DATAPATH__abc_16259_n7602;
  wire AES_CORE_DATAPATH__abc_16259_n7603;
  wire AES_CORE_DATAPATH__abc_16259_n7604;
  wire AES_CORE_DATAPATH__abc_16259_n7605;
  wire AES_CORE_DATAPATH__abc_16259_n7606;
  wire AES_CORE_DATAPATH__abc_16259_n7607;
  wire AES_CORE_DATAPATH__abc_16259_n7608;
  wire AES_CORE_DATAPATH__abc_16259_n7609;
  wire AES_CORE_DATAPATH__abc_16259_n7610;
  wire AES_CORE_DATAPATH__abc_16259_n7611;
  wire AES_CORE_DATAPATH__abc_16259_n7612;
  wire AES_CORE_DATAPATH__abc_16259_n7613;
  wire AES_CORE_DATAPATH__abc_16259_n7614;
  wire AES_CORE_DATAPATH__abc_16259_n7615;
  wire AES_CORE_DATAPATH__abc_16259_n7616;
  wire AES_CORE_DATAPATH__abc_16259_n7617;
  wire AES_CORE_DATAPATH__abc_16259_n7618;
  wire AES_CORE_DATAPATH__abc_16259_n7620;
  wire AES_CORE_DATAPATH__abc_16259_n7621;
  wire AES_CORE_DATAPATH__abc_16259_n7622;
  wire AES_CORE_DATAPATH__abc_16259_n7623;
  wire AES_CORE_DATAPATH__abc_16259_n7624;
  wire AES_CORE_DATAPATH__abc_16259_n7625;
  wire AES_CORE_DATAPATH__abc_16259_n7626;
  wire AES_CORE_DATAPATH__abc_16259_n7627;
  wire AES_CORE_DATAPATH__abc_16259_n7628;
  wire AES_CORE_DATAPATH__abc_16259_n7629;
  wire AES_CORE_DATAPATH__abc_16259_n7630;
  wire AES_CORE_DATAPATH__abc_16259_n7631;
  wire AES_CORE_DATAPATH__abc_16259_n7632;
  wire AES_CORE_DATAPATH__abc_16259_n7633;
  wire AES_CORE_DATAPATH__abc_16259_n7634;
  wire AES_CORE_DATAPATH__abc_16259_n7635;
  wire AES_CORE_DATAPATH__abc_16259_n7636;
  wire AES_CORE_DATAPATH__abc_16259_n7637;
  wire AES_CORE_DATAPATH__abc_16259_n7638;
  wire AES_CORE_DATAPATH__abc_16259_n7639;
  wire AES_CORE_DATAPATH__abc_16259_n7640;
  wire AES_CORE_DATAPATH__abc_16259_n7641;
  wire AES_CORE_DATAPATH__abc_16259_n7642;
  wire AES_CORE_DATAPATH__abc_16259_n7643;
  wire AES_CORE_DATAPATH__abc_16259_n7644;
  wire AES_CORE_DATAPATH__abc_16259_n7645;
  wire AES_CORE_DATAPATH__abc_16259_n7646;
  wire AES_CORE_DATAPATH__abc_16259_n7647;
  wire AES_CORE_DATAPATH__abc_16259_n7648;
  wire AES_CORE_DATAPATH__abc_16259_n7649;
  wire AES_CORE_DATAPATH__abc_16259_n7650;
  wire AES_CORE_DATAPATH__abc_16259_n7651;
  wire AES_CORE_DATAPATH__abc_16259_n7652;
  wire AES_CORE_DATAPATH__abc_16259_n7653;
  wire AES_CORE_DATAPATH__abc_16259_n7654;
  wire AES_CORE_DATAPATH__abc_16259_n7655;
  wire AES_CORE_DATAPATH__abc_16259_n7656;
  wire AES_CORE_DATAPATH__abc_16259_n7657;
  wire AES_CORE_DATAPATH__abc_16259_n7658;
  wire AES_CORE_DATAPATH__abc_16259_n7659;
  wire AES_CORE_DATAPATH__abc_16259_n7660;
  wire AES_CORE_DATAPATH__abc_16259_n7661;
  wire AES_CORE_DATAPATH__abc_16259_n7662;
  wire AES_CORE_DATAPATH__abc_16259_n7663;
  wire AES_CORE_DATAPATH__abc_16259_n7664;
  wire AES_CORE_DATAPATH__abc_16259_n7665;
  wire AES_CORE_DATAPATH__abc_16259_n7666;
  wire AES_CORE_DATAPATH__abc_16259_n7667;
  wire AES_CORE_DATAPATH__abc_16259_n7669;
  wire AES_CORE_DATAPATH__abc_16259_n7669_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n7669_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n7669_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n7669_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n7669_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n7670;
  wire AES_CORE_DATAPATH__abc_16259_n7671;
  wire AES_CORE_DATAPATH__abc_16259_n7672;
  wire AES_CORE_DATAPATH__abc_16259_n7673;
  wire AES_CORE_DATAPATH__abc_16259_n7674;
  wire AES_CORE_DATAPATH__abc_16259_n7675;
  wire AES_CORE_DATAPATH__abc_16259_n7676;
  wire AES_CORE_DATAPATH__abc_16259_n7678;
  wire AES_CORE_DATAPATH__abc_16259_n7679;
  wire AES_CORE_DATAPATH__abc_16259_n7680;
  wire AES_CORE_DATAPATH__abc_16259_n7681;
  wire AES_CORE_DATAPATH__abc_16259_n7682;
  wire AES_CORE_DATAPATH__abc_16259_n7683;
  wire AES_CORE_DATAPATH__abc_16259_n7684;
  wire AES_CORE_DATAPATH__abc_16259_n7686;
  wire AES_CORE_DATAPATH__abc_16259_n7687;
  wire AES_CORE_DATAPATH__abc_16259_n7688;
  wire AES_CORE_DATAPATH__abc_16259_n7689;
  wire AES_CORE_DATAPATH__abc_16259_n7690;
  wire AES_CORE_DATAPATH__abc_16259_n7691;
  wire AES_CORE_DATAPATH__abc_16259_n7692;
  wire AES_CORE_DATAPATH__abc_16259_n7694;
  wire AES_CORE_DATAPATH__abc_16259_n7695;
  wire AES_CORE_DATAPATH__abc_16259_n7696;
  wire AES_CORE_DATAPATH__abc_16259_n7697;
  wire AES_CORE_DATAPATH__abc_16259_n7698;
  wire AES_CORE_DATAPATH__abc_16259_n7699;
  wire AES_CORE_DATAPATH__abc_16259_n7700;
  wire AES_CORE_DATAPATH__abc_16259_n7702;
  wire AES_CORE_DATAPATH__abc_16259_n7703;
  wire AES_CORE_DATAPATH__abc_16259_n7704;
  wire AES_CORE_DATAPATH__abc_16259_n7705;
  wire AES_CORE_DATAPATH__abc_16259_n7706;
  wire AES_CORE_DATAPATH__abc_16259_n7707;
  wire AES_CORE_DATAPATH__abc_16259_n7708;
  wire AES_CORE_DATAPATH__abc_16259_n7710;
  wire AES_CORE_DATAPATH__abc_16259_n7711;
  wire AES_CORE_DATAPATH__abc_16259_n7712;
  wire AES_CORE_DATAPATH__abc_16259_n7713;
  wire AES_CORE_DATAPATH__abc_16259_n7714;
  wire AES_CORE_DATAPATH__abc_16259_n7715;
  wire AES_CORE_DATAPATH__abc_16259_n7716;
  wire AES_CORE_DATAPATH__abc_16259_n7718;
  wire AES_CORE_DATAPATH__abc_16259_n7719;
  wire AES_CORE_DATAPATH__abc_16259_n7720;
  wire AES_CORE_DATAPATH__abc_16259_n7721;
  wire AES_CORE_DATAPATH__abc_16259_n7722;
  wire AES_CORE_DATAPATH__abc_16259_n7723;
  wire AES_CORE_DATAPATH__abc_16259_n7724;
  wire AES_CORE_DATAPATH__abc_16259_n7726;
  wire AES_CORE_DATAPATH__abc_16259_n7727;
  wire AES_CORE_DATAPATH__abc_16259_n7728;
  wire AES_CORE_DATAPATH__abc_16259_n7729;
  wire AES_CORE_DATAPATH__abc_16259_n7730;
  wire AES_CORE_DATAPATH__abc_16259_n7731;
  wire AES_CORE_DATAPATH__abc_16259_n7732;
  wire AES_CORE_DATAPATH__abc_16259_n7734;
  wire AES_CORE_DATAPATH__abc_16259_n7735;
  wire AES_CORE_DATAPATH__abc_16259_n7736;
  wire AES_CORE_DATAPATH__abc_16259_n7737;
  wire AES_CORE_DATAPATH__abc_16259_n7738;
  wire AES_CORE_DATAPATH__abc_16259_n7739;
  wire AES_CORE_DATAPATH__abc_16259_n7740;
  wire AES_CORE_DATAPATH__abc_16259_n7742;
  wire AES_CORE_DATAPATH__abc_16259_n7743;
  wire AES_CORE_DATAPATH__abc_16259_n7744;
  wire AES_CORE_DATAPATH__abc_16259_n7745;
  wire AES_CORE_DATAPATH__abc_16259_n7746;
  wire AES_CORE_DATAPATH__abc_16259_n7747;
  wire AES_CORE_DATAPATH__abc_16259_n7748;
  wire AES_CORE_DATAPATH__abc_16259_n7750;
  wire AES_CORE_DATAPATH__abc_16259_n7751;
  wire AES_CORE_DATAPATH__abc_16259_n7752;
  wire AES_CORE_DATAPATH__abc_16259_n7753;
  wire AES_CORE_DATAPATH__abc_16259_n7754;
  wire AES_CORE_DATAPATH__abc_16259_n7755;
  wire AES_CORE_DATAPATH__abc_16259_n7756;
  wire AES_CORE_DATAPATH__abc_16259_n7757;
  wire AES_CORE_DATAPATH__abc_16259_n7758;
  wire AES_CORE_DATAPATH__abc_16259_n7759;
  wire AES_CORE_DATAPATH__abc_16259_n7761;
  wire AES_CORE_DATAPATH__abc_16259_n7762;
  wire AES_CORE_DATAPATH__abc_16259_n7763;
  wire AES_CORE_DATAPATH__abc_16259_n7764;
  wire AES_CORE_DATAPATH__abc_16259_n7765;
  wire AES_CORE_DATAPATH__abc_16259_n7766;
  wire AES_CORE_DATAPATH__abc_16259_n7767;
  wire AES_CORE_DATAPATH__abc_16259_n7768;
  wire AES_CORE_DATAPATH__abc_16259_n7769;
  wire AES_CORE_DATAPATH__abc_16259_n7770;
  wire AES_CORE_DATAPATH__abc_16259_n7772;
  wire AES_CORE_DATAPATH__abc_16259_n7773;
  wire AES_CORE_DATAPATH__abc_16259_n7774;
  wire AES_CORE_DATAPATH__abc_16259_n7775;
  wire AES_CORE_DATAPATH__abc_16259_n7776;
  wire AES_CORE_DATAPATH__abc_16259_n7777;
  wire AES_CORE_DATAPATH__abc_16259_n7778;
  wire AES_CORE_DATAPATH__abc_16259_n7780;
  wire AES_CORE_DATAPATH__abc_16259_n7781;
  wire AES_CORE_DATAPATH__abc_16259_n7782;
  wire AES_CORE_DATAPATH__abc_16259_n7783;
  wire AES_CORE_DATAPATH__abc_16259_n7784;
  wire AES_CORE_DATAPATH__abc_16259_n7785;
  wire AES_CORE_DATAPATH__abc_16259_n7786;
  wire AES_CORE_DATAPATH__abc_16259_n7787;
  wire AES_CORE_DATAPATH__abc_16259_n7788;
  wire AES_CORE_DATAPATH__abc_16259_n7789;
  wire AES_CORE_DATAPATH__abc_16259_n7791;
  wire AES_CORE_DATAPATH__abc_16259_n7792;
  wire AES_CORE_DATAPATH__abc_16259_n7793;
  wire AES_CORE_DATAPATH__abc_16259_n7794;
  wire AES_CORE_DATAPATH__abc_16259_n7795;
  wire AES_CORE_DATAPATH__abc_16259_n7796;
  wire AES_CORE_DATAPATH__abc_16259_n7797;
  wire AES_CORE_DATAPATH__abc_16259_n7799;
  wire AES_CORE_DATAPATH__abc_16259_n7800;
  wire AES_CORE_DATAPATH__abc_16259_n7801;
  wire AES_CORE_DATAPATH__abc_16259_n7802;
  wire AES_CORE_DATAPATH__abc_16259_n7803;
  wire AES_CORE_DATAPATH__abc_16259_n7804;
  wire AES_CORE_DATAPATH__abc_16259_n7805;
  wire AES_CORE_DATAPATH__abc_16259_n7806;
  wire AES_CORE_DATAPATH__abc_16259_n7807;
  wire AES_CORE_DATAPATH__abc_16259_n7808;
  wire AES_CORE_DATAPATH__abc_16259_n7810;
  wire AES_CORE_DATAPATH__abc_16259_n7811;
  wire AES_CORE_DATAPATH__abc_16259_n7812;
  wire AES_CORE_DATAPATH__abc_16259_n7813;
  wire AES_CORE_DATAPATH__abc_16259_n7814;
  wire AES_CORE_DATAPATH__abc_16259_n7815;
  wire AES_CORE_DATAPATH__abc_16259_n7816;
  wire AES_CORE_DATAPATH__abc_16259_n7818;
  wire AES_CORE_DATAPATH__abc_16259_n7819;
  wire AES_CORE_DATAPATH__abc_16259_n7820;
  wire AES_CORE_DATAPATH__abc_16259_n7821;
  wire AES_CORE_DATAPATH__abc_16259_n7822;
  wire AES_CORE_DATAPATH__abc_16259_n7823;
  wire AES_CORE_DATAPATH__abc_16259_n7824;
  wire AES_CORE_DATAPATH__abc_16259_n7825;
  wire AES_CORE_DATAPATH__abc_16259_n7826;
  wire AES_CORE_DATAPATH__abc_16259_n7827;
  wire AES_CORE_DATAPATH__abc_16259_n7829;
  wire AES_CORE_DATAPATH__abc_16259_n7830;
  wire AES_CORE_DATAPATH__abc_16259_n7831;
  wire AES_CORE_DATAPATH__abc_16259_n7832;
  wire AES_CORE_DATAPATH__abc_16259_n7833;
  wire AES_CORE_DATAPATH__abc_16259_n7834;
  wire AES_CORE_DATAPATH__abc_16259_n7835;
  wire AES_CORE_DATAPATH__abc_16259_n7837;
  wire AES_CORE_DATAPATH__abc_16259_n7838;
  wire AES_CORE_DATAPATH__abc_16259_n7839;
  wire AES_CORE_DATAPATH__abc_16259_n7840;
  wire AES_CORE_DATAPATH__abc_16259_n7841;
  wire AES_CORE_DATAPATH__abc_16259_n7842;
  wire AES_CORE_DATAPATH__abc_16259_n7843;
  wire AES_CORE_DATAPATH__abc_16259_n7845;
  wire AES_CORE_DATAPATH__abc_16259_n7846;
  wire AES_CORE_DATAPATH__abc_16259_n7847;
  wire AES_CORE_DATAPATH__abc_16259_n7848;
  wire AES_CORE_DATAPATH__abc_16259_n7849;
  wire AES_CORE_DATAPATH__abc_16259_n7850;
  wire AES_CORE_DATAPATH__abc_16259_n7851;
  wire AES_CORE_DATAPATH__abc_16259_n7853;
  wire AES_CORE_DATAPATH__abc_16259_n7854;
  wire AES_CORE_DATAPATH__abc_16259_n7855;
  wire AES_CORE_DATAPATH__abc_16259_n7856;
  wire AES_CORE_DATAPATH__abc_16259_n7857;
  wire AES_CORE_DATAPATH__abc_16259_n7858;
  wire AES_CORE_DATAPATH__abc_16259_n7859;
  wire AES_CORE_DATAPATH__abc_16259_n7860;
  wire AES_CORE_DATAPATH__abc_16259_n7861;
  wire AES_CORE_DATAPATH__abc_16259_n7862;
  wire AES_CORE_DATAPATH__abc_16259_n7864;
  wire AES_CORE_DATAPATH__abc_16259_n7865;
  wire AES_CORE_DATAPATH__abc_16259_n7866;
  wire AES_CORE_DATAPATH__abc_16259_n7867;
  wire AES_CORE_DATAPATH__abc_16259_n7868;
  wire AES_CORE_DATAPATH__abc_16259_n7869;
  wire AES_CORE_DATAPATH__abc_16259_n7870;
  wire AES_CORE_DATAPATH__abc_16259_n7872;
  wire AES_CORE_DATAPATH__abc_16259_n7873;
  wire AES_CORE_DATAPATH__abc_16259_n7874;
  wire AES_CORE_DATAPATH__abc_16259_n7875;
  wire AES_CORE_DATAPATH__abc_16259_n7876;
  wire AES_CORE_DATAPATH__abc_16259_n7877;
  wire AES_CORE_DATAPATH__abc_16259_n7878;
  wire AES_CORE_DATAPATH__abc_16259_n7880;
  wire AES_CORE_DATAPATH__abc_16259_n7881;
  wire AES_CORE_DATAPATH__abc_16259_n7882;
  wire AES_CORE_DATAPATH__abc_16259_n7883;
  wire AES_CORE_DATAPATH__abc_16259_n7884;
  wire AES_CORE_DATAPATH__abc_16259_n7885;
  wire AES_CORE_DATAPATH__abc_16259_n7886;
  wire AES_CORE_DATAPATH__abc_16259_n7888;
  wire AES_CORE_DATAPATH__abc_16259_n7889;
  wire AES_CORE_DATAPATH__abc_16259_n7890;
  wire AES_CORE_DATAPATH__abc_16259_n7891;
  wire AES_CORE_DATAPATH__abc_16259_n7892;
  wire AES_CORE_DATAPATH__abc_16259_n7893;
  wire AES_CORE_DATAPATH__abc_16259_n7894;
  wire AES_CORE_DATAPATH__abc_16259_n7896;
  wire AES_CORE_DATAPATH__abc_16259_n7897;
  wire AES_CORE_DATAPATH__abc_16259_n7898;
  wire AES_CORE_DATAPATH__abc_16259_n7899;
  wire AES_CORE_DATAPATH__abc_16259_n7900;
  wire AES_CORE_DATAPATH__abc_16259_n7901;
  wire AES_CORE_DATAPATH__abc_16259_n7902;
  wire AES_CORE_DATAPATH__abc_16259_n7904;
  wire AES_CORE_DATAPATH__abc_16259_n7905;
  wire AES_CORE_DATAPATH__abc_16259_n7906;
  wire AES_CORE_DATAPATH__abc_16259_n7907;
  wire AES_CORE_DATAPATH__abc_16259_n7908;
  wire AES_CORE_DATAPATH__abc_16259_n7909;
  wire AES_CORE_DATAPATH__abc_16259_n7910;
  wire AES_CORE_DATAPATH__abc_16259_n7912;
  wire AES_CORE_DATAPATH__abc_16259_n7913;
  wire AES_CORE_DATAPATH__abc_16259_n7914;
  wire AES_CORE_DATAPATH__abc_16259_n7915;
  wire AES_CORE_DATAPATH__abc_16259_n7916;
  wire AES_CORE_DATAPATH__abc_16259_n7917;
  wire AES_CORE_DATAPATH__abc_16259_n7918;
  wire AES_CORE_DATAPATH__abc_16259_n7920;
  wire AES_CORE_DATAPATH__abc_16259_n7921;
  wire AES_CORE_DATAPATH__abc_16259_n7922;
  wire AES_CORE_DATAPATH__abc_16259_n7923;
  wire AES_CORE_DATAPATH__abc_16259_n7924;
  wire AES_CORE_DATAPATH__abc_16259_n7925;
  wire AES_CORE_DATAPATH__abc_16259_n7926;
  wire AES_CORE_DATAPATH__abc_16259_n7928;
  wire AES_CORE_DATAPATH__abc_16259_n7929;
  wire AES_CORE_DATAPATH__abc_16259_n7930;
  wire AES_CORE_DATAPATH__abc_16259_n7931;
  wire AES_CORE_DATAPATH__abc_16259_n7932;
  wire AES_CORE_DATAPATH__abc_16259_n7933;
  wire AES_CORE_DATAPATH__abc_16259_n7934;
  wire AES_CORE_DATAPATH__abc_16259_n7936;
  wire AES_CORE_DATAPATH__abc_16259_n7937;
  wire AES_CORE_DATAPATH__abc_16259_n7938;
  wire AES_CORE_DATAPATH__abc_16259_n7939;
  wire AES_CORE_DATAPATH__abc_16259_n7940;
  wire AES_CORE_DATAPATH__abc_16259_n7941;
  wire AES_CORE_DATAPATH__abc_16259_n7942;
  wire AES_CORE_DATAPATH__abc_16259_n7944;
  wire AES_CORE_DATAPATH__abc_16259_n7944_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n7944_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n7944_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n7944_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n7944_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n7945;
  wire AES_CORE_DATAPATH__abc_16259_n7946;
  wire AES_CORE_DATAPATH__abc_16259_n7947;
  wire AES_CORE_DATAPATH__abc_16259_n7948;
  wire AES_CORE_DATAPATH__abc_16259_n7949;
  wire AES_CORE_DATAPATH__abc_16259_n7950;
  wire AES_CORE_DATAPATH__abc_16259_n7951;
  wire AES_CORE_DATAPATH__abc_16259_n7953;
  wire AES_CORE_DATAPATH__abc_16259_n7954;
  wire AES_CORE_DATAPATH__abc_16259_n7955;
  wire AES_CORE_DATAPATH__abc_16259_n7956;
  wire AES_CORE_DATAPATH__abc_16259_n7957;
  wire AES_CORE_DATAPATH__abc_16259_n7958;
  wire AES_CORE_DATAPATH__abc_16259_n7959;
  wire AES_CORE_DATAPATH__abc_16259_n7961;
  wire AES_CORE_DATAPATH__abc_16259_n7962;
  wire AES_CORE_DATAPATH__abc_16259_n7963;
  wire AES_CORE_DATAPATH__abc_16259_n7964;
  wire AES_CORE_DATAPATH__abc_16259_n7965;
  wire AES_CORE_DATAPATH__abc_16259_n7966;
  wire AES_CORE_DATAPATH__abc_16259_n7967;
  wire AES_CORE_DATAPATH__abc_16259_n7969;
  wire AES_CORE_DATAPATH__abc_16259_n7970;
  wire AES_CORE_DATAPATH__abc_16259_n7971;
  wire AES_CORE_DATAPATH__abc_16259_n7972;
  wire AES_CORE_DATAPATH__abc_16259_n7973;
  wire AES_CORE_DATAPATH__abc_16259_n7974;
  wire AES_CORE_DATAPATH__abc_16259_n7975;
  wire AES_CORE_DATAPATH__abc_16259_n7977;
  wire AES_CORE_DATAPATH__abc_16259_n7978;
  wire AES_CORE_DATAPATH__abc_16259_n7979;
  wire AES_CORE_DATAPATH__abc_16259_n7980;
  wire AES_CORE_DATAPATH__abc_16259_n7981;
  wire AES_CORE_DATAPATH__abc_16259_n7982;
  wire AES_CORE_DATAPATH__abc_16259_n7983;
  wire AES_CORE_DATAPATH__abc_16259_n7985;
  wire AES_CORE_DATAPATH__abc_16259_n7986;
  wire AES_CORE_DATAPATH__abc_16259_n7987;
  wire AES_CORE_DATAPATH__abc_16259_n7988;
  wire AES_CORE_DATAPATH__abc_16259_n7989;
  wire AES_CORE_DATAPATH__abc_16259_n7990;
  wire AES_CORE_DATAPATH__abc_16259_n7991;
  wire AES_CORE_DATAPATH__abc_16259_n7993;
  wire AES_CORE_DATAPATH__abc_16259_n7994;
  wire AES_CORE_DATAPATH__abc_16259_n7995;
  wire AES_CORE_DATAPATH__abc_16259_n7996;
  wire AES_CORE_DATAPATH__abc_16259_n7997;
  wire AES_CORE_DATAPATH__abc_16259_n7998;
  wire AES_CORE_DATAPATH__abc_16259_n7999;
  wire AES_CORE_DATAPATH__abc_16259_n8001;
  wire AES_CORE_DATAPATH__abc_16259_n8002;
  wire AES_CORE_DATAPATH__abc_16259_n8003;
  wire AES_CORE_DATAPATH__abc_16259_n8004;
  wire AES_CORE_DATAPATH__abc_16259_n8005;
  wire AES_CORE_DATAPATH__abc_16259_n8006;
  wire AES_CORE_DATAPATH__abc_16259_n8007;
  wire AES_CORE_DATAPATH__abc_16259_n8009;
  wire AES_CORE_DATAPATH__abc_16259_n8010;
  wire AES_CORE_DATAPATH__abc_16259_n8011;
  wire AES_CORE_DATAPATH__abc_16259_n8012;
  wire AES_CORE_DATAPATH__abc_16259_n8013;
  wire AES_CORE_DATAPATH__abc_16259_n8014;
  wire AES_CORE_DATAPATH__abc_16259_n8015;
  wire AES_CORE_DATAPATH__abc_16259_n8017;
  wire AES_CORE_DATAPATH__abc_16259_n8018;
  wire AES_CORE_DATAPATH__abc_16259_n8019;
  wire AES_CORE_DATAPATH__abc_16259_n8020;
  wire AES_CORE_DATAPATH__abc_16259_n8021;
  wire AES_CORE_DATAPATH__abc_16259_n8022;
  wire AES_CORE_DATAPATH__abc_16259_n8023;
  wire AES_CORE_DATAPATH__abc_16259_n8025;
  wire AES_CORE_DATAPATH__abc_16259_n8026;
  wire AES_CORE_DATAPATH__abc_16259_n8027;
  wire AES_CORE_DATAPATH__abc_16259_n8028;
  wire AES_CORE_DATAPATH__abc_16259_n8029;
  wire AES_CORE_DATAPATH__abc_16259_n8030;
  wire AES_CORE_DATAPATH__abc_16259_n8031;
  wire AES_CORE_DATAPATH__abc_16259_n8032;
  wire AES_CORE_DATAPATH__abc_16259_n8033;
  wire AES_CORE_DATAPATH__abc_16259_n8034;
  wire AES_CORE_DATAPATH__abc_16259_n8036;
  wire AES_CORE_DATAPATH__abc_16259_n8037;
  wire AES_CORE_DATAPATH__abc_16259_n8038;
  wire AES_CORE_DATAPATH__abc_16259_n8039;
  wire AES_CORE_DATAPATH__abc_16259_n8040;
  wire AES_CORE_DATAPATH__abc_16259_n8041;
  wire AES_CORE_DATAPATH__abc_16259_n8042;
  wire AES_CORE_DATAPATH__abc_16259_n8043;
  wire AES_CORE_DATAPATH__abc_16259_n8044;
  wire AES_CORE_DATAPATH__abc_16259_n8045;
  wire AES_CORE_DATAPATH__abc_16259_n8047;
  wire AES_CORE_DATAPATH__abc_16259_n8048;
  wire AES_CORE_DATAPATH__abc_16259_n8049;
  wire AES_CORE_DATAPATH__abc_16259_n8050;
  wire AES_CORE_DATAPATH__abc_16259_n8051;
  wire AES_CORE_DATAPATH__abc_16259_n8052;
  wire AES_CORE_DATAPATH__abc_16259_n8053;
  wire AES_CORE_DATAPATH__abc_16259_n8055;
  wire AES_CORE_DATAPATH__abc_16259_n8056;
  wire AES_CORE_DATAPATH__abc_16259_n8057;
  wire AES_CORE_DATAPATH__abc_16259_n8058;
  wire AES_CORE_DATAPATH__abc_16259_n8059;
  wire AES_CORE_DATAPATH__abc_16259_n8060;
  wire AES_CORE_DATAPATH__abc_16259_n8061;
  wire AES_CORE_DATAPATH__abc_16259_n8062;
  wire AES_CORE_DATAPATH__abc_16259_n8063;
  wire AES_CORE_DATAPATH__abc_16259_n8064;
  wire AES_CORE_DATAPATH__abc_16259_n8066;
  wire AES_CORE_DATAPATH__abc_16259_n8067;
  wire AES_CORE_DATAPATH__abc_16259_n8068;
  wire AES_CORE_DATAPATH__abc_16259_n8069;
  wire AES_CORE_DATAPATH__abc_16259_n8070;
  wire AES_CORE_DATAPATH__abc_16259_n8071;
  wire AES_CORE_DATAPATH__abc_16259_n8072;
  wire AES_CORE_DATAPATH__abc_16259_n8074;
  wire AES_CORE_DATAPATH__abc_16259_n8075;
  wire AES_CORE_DATAPATH__abc_16259_n8076;
  wire AES_CORE_DATAPATH__abc_16259_n8077;
  wire AES_CORE_DATAPATH__abc_16259_n8078;
  wire AES_CORE_DATAPATH__abc_16259_n8079;
  wire AES_CORE_DATAPATH__abc_16259_n8080;
  wire AES_CORE_DATAPATH__abc_16259_n8081;
  wire AES_CORE_DATAPATH__abc_16259_n8082;
  wire AES_CORE_DATAPATH__abc_16259_n8083;
  wire AES_CORE_DATAPATH__abc_16259_n8085;
  wire AES_CORE_DATAPATH__abc_16259_n8086;
  wire AES_CORE_DATAPATH__abc_16259_n8087;
  wire AES_CORE_DATAPATH__abc_16259_n8088;
  wire AES_CORE_DATAPATH__abc_16259_n8089;
  wire AES_CORE_DATAPATH__abc_16259_n8090;
  wire AES_CORE_DATAPATH__abc_16259_n8091;
  wire AES_CORE_DATAPATH__abc_16259_n8093;
  wire AES_CORE_DATAPATH__abc_16259_n8094;
  wire AES_CORE_DATAPATH__abc_16259_n8095;
  wire AES_CORE_DATAPATH__abc_16259_n8096;
  wire AES_CORE_DATAPATH__abc_16259_n8097;
  wire AES_CORE_DATAPATH__abc_16259_n8098;
  wire AES_CORE_DATAPATH__abc_16259_n8099;
  wire AES_CORE_DATAPATH__abc_16259_n8100;
  wire AES_CORE_DATAPATH__abc_16259_n8101;
  wire AES_CORE_DATAPATH__abc_16259_n8102;
  wire AES_CORE_DATAPATH__abc_16259_n8104;
  wire AES_CORE_DATAPATH__abc_16259_n8105;
  wire AES_CORE_DATAPATH__abc_16259_n8106;
  wire AES_CORE_DATAPATH__abc_16259_n8107;
  wire AES_CORE_DATAPATH__abc_16259_n8108;
  wire AES_CORE_DATAPATH__abc_16259_n8109;
  wire AES_CORE_DATAPATH__abc_16259_n8110;
  wire AES_CORE_DATAPATH__abc_16259_n8112;
  wire AES_CORE_DATAPATH__abc_16259_n8113;
  wire AES_CORE_DATAPATH__abc_16259_n8114;
  wire AES_CORE_DATAPATH__abc_16259_n8115;
  wire AES_CORE_DATAPATH__abc_16259_n8116;
  wire AES_CORE_DATAPATH__abc_16259_n8117;
  wire AES_CORE_DATAPATH__abc_16259_n8118;
  wire AES_CORE_DATAPATH__abc_16259_n8120;
  wire AES_CORE_DATAPATH__abc_16259_n8121;
  wire AES_CORE_DATAPATH__abc_16259_n8122;
  wire AES_CORE_DATAPATH__abc_16259_n8123;
  wire AES_CORE_DATAPATH__abc_16259_n8124;
  wire AES_CORE_DATAPATH__abc_16259_n8125;
  wire AES_CORE_DATAPATH__abc_16259_n8126;
  wire AES_CORE_DATAPATH__abc_16259_n8128;
  wire AES_CORE_DATAPATH__abc_16259_n8129;
  wire AES_CORE_DATAPATH__abc_16259_n8130;
  wire AES_CORE_DATAPATH__abc_16259_n8131;
  wire AES_CORE_DATAPATH__abc_16259_n8132;
  wire AES_CORE_DATAPATH__abc_16259_n8133;
  wire AES_CORE_DATAPATH__abc_16259_n8134;
  wire AES_CORE_DATAPATH__abc_16259_n8135;
  wire AES_CORE_DATAPATH__abc_16259_n8136;
  wire AES_CORE_DATAPATH__abc_16259_n8137;
  wire AES_CORE_DATAPATH__abc_16259_n8139;
  wire AES_CORE_DATAPATH__abc_16259_n8140;
  wire AES_CORE_DATAPATH__abc_16259_n8141;
  wire AES_CORE_DATAPATH__abc_16259_n8142;
  wire AES_CORE_DATAPATH__abc_16259_n8143;
  wire AES_CORE_DATAPATH__abc_16259_n8144;
  wire AES_CORE_DATAPATH__abc_16259_n8145;
  wire AES_CORE_DATAPATH__abc_16259_n8147;
  wire AES_CORE_DATAPATH__abc_16259_n8148;
  wire AES_CORE_DATAPATH__abc_16259_n8149;
  wire AES_CORE_DATAPATH__abc_16259_n8150;
  wire AES_CORE_DATAPATH__abc_16259_n8151;
  wire AES_CORE_DATAPATH__abc_16259_n8152;
  wire AES_CORE_DATAPATH__abc_16259_n8153;
  wire AES_CORE_DATAPATH__abc_16259_n8155;
  wire AES_CORE_DATAPATH__abc_16259_n8156;
  wire AES_CORE_DATAPATH__abc_16259_n8157;
  wire AES_CORE_DATAPATH__abc_16259_n8158;
  wire AES_CORE_DATAPATH__abc_16259_n8159;
  wire AES_CORE_DATAPATH__abc_16259_n8160;
  wire AES_CORE_DATAPATH__abc_16259_n8161;
  wire AES_CORE_DATAPATH__abc_16259_n8163;
  wire AES_CORE_DATAPATH__abc_16259_n8164;
  wire AES_CORE_DATAPATH__abc_16259_n8165;
  wire AES_CORE_DATAPATH__abc_16259_n8166;
  wire AES_CORE_DATAPATH__abc_16259_n8167;
  wire AES_CORE_DATAPATH__abc_16259_n8168;
  wire AES_CORE_DATAPATH__abc_16259_n8169;
  wire AES_CORE_DATAPATH__abc_16259_n8171;
  wire AES_CORE_DATAPATH__abc_16259_n8172;
  wire AES_CORE_DATAPATH__abc_16259_n8173;
  wire AES_CORE_DATAPATH__abc_16259_n8174;
  wire AES_CORE_DATAPATH__abc_16259_n8175;
  wire AES_CORE_DATAPATH__abc_16259_n8176;
  wire AES_CORE_DATAPATH__abc_16259_n8177;
  wire AES_CORE_DATAPATH__abc_16259_n8179;
  wire AES_CORE_DATAPATH__abc_16259_n8180;
  wire AES_CORE_DATAPATH__abc_16259_n8181;
  wire AES_CORE_DATAPATH__abc_16259_n8182;
  wire AES_CORE_DATAPATH__abc_16259_n8183;
  wire AES_CORE_DATAPATH__abc_16259_n8184;
  wire AES_CORE_DATAPATH__abc_16259_n8185;
  wire AES_CORE_DATAPATH__abc_16259_n8187;
  wire AES_CORE_DATAPATH__abc_16259_n8188;
  wire AES_CORE_DATAPATH__abc_16259_n8189;
  wire AES_CORE_DATAPATH__abc_16259_n8190;
  wire AES_CORE_DATAPATH__abc_16259_n8191;
  wire AES_CORE_DATAPATH__abc_16259_n8192;
  wire AES_CORE_DATAPATH__abc_16259_n8193;
  wire AES_CORE_DATAPATH__abc_16259_n8195;
  wire AES_CORE_DATAPATH__abc_16259_n8196;
  wire AES_CORE_DATAPATH__abc_16259_n8197;
  wire AES_CORE_DATAPATH__abc_16259_n8198;
  wire AES_CORE_DATAPATH__abc_16259_n8199;
  wire AES_CORE_DATAPATH__abc_16259_n8200;
  wire AES_CORE_DATAPATH__abc_16259_n8201;
  wire AES_CORE_DATAPATH__abc_16259_n8203;
  wire AES_CORE_DATAPATH__abc_16259_n8204;
  wire AES_CORE_DATAPATH__abc_16259_n8205;
  wire AES_CORE_DATAPATH__abc_16259_n8206;
  wire AES_CORE_DATAPATH__abc_16259_n8207;
  wire AES_CORE_DATAPATH__abc_16259_n8208;
  wire AES_CORE_DATAPATH__abc_16259_n8209;
  wire AES_CORE_DATAPATH__abc_16259_n8211;
  wire AES_CORE_DATAPATH__abc_16259_n8212;
  wire AES_CORE_DATAPATH__abc_16259_n8213;
  wire AES_CORE_DATAPATH__abc_16259_n8214;
  wire AES_CORE_DATAPATH__abc_16259_n8215;
  wire AES_CORE_DATAPATH__abc_16259_n8216;
  wire AES_CORE_DATAPATH__abc_16259_n8217;
  wire AES_CORE_DATAPATH__abc_16259_n8219;
  wire AES_CORE_DATAPATH__abc_16259_n8219_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n8219_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n8219_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n8219_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n8219_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n8220;
  wire AES_CORE_DATAPATH__abc_16259_n8221;
  wire AES_CORE_DATAPATH__abc_16259_n8222;
  wire AES_CORE_DATAPATH__abc_16259_n8223;
  wire AES_CORE_DATAPATH__abc_16259_n8224;
  wire AES_CORE_DATAPATH__abc_16259_n8225;
  wire AES_CORE_DATAPATH__abc_16259_n8226;
  wire AES_CORE_DATAPATH__abc_16259_n8228;
  wire AES_CORE_DATAPATH__abc_16259_n8229;
  wire AES_CORE_DATAPATH__abc_16259_n8230;
  wire AES_CORE_DATAPATH__abc_16259_n8231;
  wire AES_CORE_DATAPATH__abc_16259_n8232;
  wire AES_CORE_DATAPATH__abc_16259_n8233;
  wire AES_CORE_DATAPATH__abc_16259_n8234;
  wire AES_CORE_DATAPATH__abc_16259_n8236;
  wire AES_CORE_DATAPATH__abc_16259_n8237;
  wire AES_CORE_DATAPATH__abc_16259_n8238;
  wire AES_CORE_DATAPATH__abc_16259_n8239;
  wire AES_CORE_DATAPATH__abc_16259_n8240;
  wire AES_CORE_DATAPATH__abc_16259_n8241;
  wire AES_CORE_DATAPATH__abc_16259_n8242;
  wire AES_CORE_DATAPATH__abc_16259_n8244;
  wire AES_CORE_DATAPATH__abc_16259_n8245;
  wire AES_CORE_DATAPATH__abc_16259_n8246;
  wire AES_CORE_DATAPATH__abc_16259_n8247;
  wire AES_CORE_DATAPATH__abc_16259_n8248;
  wire AES_CORE_DATAPATH__abc_16259_n8249;
  wire AES_CORE_DATAPATH__abc_16259_n8250;
  wire AES_CORE_DATAPATH__abc_16259_n8252;
  wire AES_CORE_DATAPATH__abc_16259_n8253;
  wire AES_CORE_DATAPATH__abc_16259_n8254;
  wire AES_CORE_DATAPATH__abc_16259_n8255;
  wire AES_CORE_DATAPATH__abc_16259_n8256;
  wire AES_CORE_DATAPATH__abc_16259_n8257;
  wire AES_CORE_DATAPATH__abc_16259_n8258;
  wire AES_CORE_DATAPATH__abc_16259_n8260;
  wire AES_CORE_DATAPATH__abc_16259_n8261;
  wire AES_CORE_DATAPATH__abc_16259_n8262;
  wire AES_CORE_DATAPATH__abc_16259_n8263;
  wire AES_CORE_DATAPATH__abc_16259_n8264;
  wire AES_CORE_DATAPATH__abc_16259_n8265;
  wire AES_CORE_DATAPATH__abc_16259_n8266;
  wire AES_CORE_DATAPATH__abc_16259_n8268;
  wire AES_CORE_DATAPATH__abc_16259_n8269;
  wire AES_CORE_DATAPATH__abc_16259_n8270;
  wire AES_CORE_DATAPATH__abc_16259_n8271;
  wire AES_CORE_DATAPATH__abc_16259_n8272;
  wire AES_CORE_DATAPATH__abc_16259_n8273;
  wire AES_CORE_DATAPATH__abc_16259_n8274;
  wire AES_CORE_DATAPATH__abc_16259_n8276;
  wire AES_CORE_DATAPATH__abc_16259_n8277;
  wire AES_CORE_DATAPATH__abc_16259_n8278;
  wire AES_CORE_DATAPATH__abc_16259_n8279;
  wire AES_CORE_DATAPATH__abc_16259_n8280;
  wire AES_CORE_DATAPATH__abc_16259_n8281;
  wire AES_CORE_DATAPATH__abc_16259_n8282;
  wire AES_CORE_DATAPATH__abc_16259_n8284;
  wire AES_CORE_DATAPATH__abc_16259_n8285;
  wire AES_CORE_DATAPATH__abc_16259_n8286;
  wire AES_CORE_DATAPATH__abc_16259_n8287;
  wire AES_CORE_DATAPATH__abc_16259_n8288;
  wire AES_CORE_DATAPATH__abc_16259_n8289;
  wire AES_CORE_DATAPATH__abc_16259_n8290;
  wire AES_CORE_DATAPATH__abc_16259_n8292;
  wire AES_CORE_DATAPATH__abc_16259_n8293;
  wire AES_CORE_DATAPATH__abc_16259_n8294;
  wire AES_CORE_DATAPATH__abc_16259_n8295;
  wire AES_CORE_DATAPATH__abc_16259_n8296;
  wire AES_CORE_DATAPATH__abc_16259_n8297;
  wire AES_CORE_DATAPATH__abc_16259_n8298;
  wire AES_CORE_DATAPATH__abc_16259_n8300;
  wire AES_CORE_DATAPATH__abc_16259_n8301;
  wire AES_CORE_DATAPATH__abc_16259_n8302;
  wire AES_CORE_DATAPATH__abc_16259_n8303;
  wire AES_CORE_DATAPATH__abc_16259_n8304;
  wire AES_CORE_DATAPATH__abc_16259_n8305;
  wire AES_CORE_DATAPATH__abc_16259_n8306;
  wire AES_CORE_DATAPATH__abc_16259_n8307;
  wire AES_CORE_DATAPATH__abc_16259_n8308;
  wire AES_CORE_DATAPATH__abc_16259_n8309;
  wire AES_CORE_DATAPATH__abc_16259_n8311;
  wire AES_CORE_DATAPATH__abc_16259_n8312;
  wire AES_CORE_DATAPATH__abc_16259_n8313;
  wire AES_CORE_DATAPATH__abc_16259_n8314;
  wire AES_CORE_DATAPATH__abc_16259_n8315;
  wire AES_CORE_DATAPATH__abc_16259_n8316;
  wire AES_CORE_DATAPATH__abc_16259_n8317;
  wire AES_CORE_DATAPATH__abc_16259_n8318;
  wire AES_CORE_DATAPATH__abc_16259_n8319;
  wire AES_CORE_DATAPATH__abc_16259_n8320;
  wire AES_CORE_DATAPATH__abc_16259_n8322;
  wire AES_CORE_DATAPATH__abc_16259_n8323;
  wire AES_CORE_DATAPATH__abc_16259_n8324;
  wire AES_CORE_DATAPATH__abc_16259_n8325;
  wire AES_CORE_DATAPATH__abc_16259_n8326;
  wire AES_CORE_DATAPATH__abc_16259_n8327;
  wire AES_CORE_DATAPATH__abc_16259_n8328;
  wire AES_CORE_DATAPATH__abc_16259_n8330;
  wire AES_CORE_DATAPATH__abc_16259_n8331;
  wire AES_CORE_DATAPATH__abc_16259_n8332;
  wire AES_CORE_DATAPATH__abc_16259_n8333;
  wire AES_CORE_DATAPATH__abc_16259_n8334;
  wire AES_CORE_DATAPATH__abc_16259_n8335;
  wire AES_CORE_DATAPATH__abc_16259_n8336;
  wire AES_CORE_DATAPATH__abc_16259_n8337;
  wire AES_CORE_DATAPATH__abc_16259_n8338;
  wire AES_CORE_DATAPATH__abc_16259_n8339;
  wire AES_CORE_DATAPATH__abc_16259_n8341;
  wire AES_CORE_DATAPATH__abc_16259_n8342;
  wire AES_CORE_DATAPATH__abc_16259_n8343;
  wire AES_CORE_DATAPATH__abc_16259_n8344;
  wire AES_CORE_DATAPATH__abc_16259_n8345;
  wire AES_CORE_DATAPATH__abc_16259_n8346;
  wire AES_CORE_DATAPATH__abc_16259_n8347;
  wire AES_CORE_DATAPATH__abc_16259_n8349;
  wire AES_CORE_DATAPATH__abc_16259_n8350;
  wire AES_CORE_DATAPATH__abc_16259_n8351;
  wire AES_CORE_DATAPATH__abc_16259_n8352;
  wire AES_CORE_DATAPATH__abc_16259_n8353;
  wire AES_CORE_DATAPATH__abc_16259_n8354;
  wire AES_CORE_DATAPATH__abc_16259_n8355;
  wire AES_CORE_DATAPATH__abc_16259_n8356;
  wire AES_CORE_DATAPATH__abc_16259_n8357;
  wire AES_CORE_DATAPATH__abc_16259_n8358;
  wire AES_CORE_DATAPATH__abc_16259_n8360;
  wire AES_CORE_DATAPATH__abc_16259_n8361;
  wire AES_CORE_DATAPATH__abc_16259_n8362;
  wire AES_CORE_DATAPATH__abc_16259_n8363;
  wire AES_CORE_DATAPATH__abc_16259_n8364;
  wire AES_CORE_DATAPATH__abc_16259_n8365;
  wire AES_CORE_DATAPATH__abc_16259_n8366;
  wire AES_CORE_DATAPATH__abc_16259_n8368;
  wire AES_CORE_DATAPATH__abc_16259_n8369;
  wire AES_CORE_DATAPATH__abc_16259_n8370;
  wire AES_CORE_DATAPATH__abc_16259_n8371;
  wire AES_CORE_DATAPATH__abc_16259_n8372;
  wire AES_CORE_DATAPATH__abc_16259_n8373;
  wire AES_CORE_DATAPATH__abc_16259_n8374;
  wire AES_CORE_DATAPATH__abc_16259_n8375;
  wire AES_CORE_DATAPATH__abc_16259_n8376;
  wire AES_CORE_DATAPATH__abc_16259_n8377;
  wire AES_CORE_DATAPATH__abc_16259_n8379;
  wire AES_CORE_DATAPATH__abc_16259_n8380;
  wire AES_CORE_DATAPATH__abc_16259_n8381;
  wire AES_CORE_DATAPATH__abc_16259_n8382;
  wire AES_CORE_DATAPATH__abc_16259_n8383;
  wire AES_CORE_DATAPATH__abc_16259_n8384;
  wire AES_CORE_DATAPATH__abc_16259_n8385;
  wire AES_CORE_DATAPATH__abc_16259_n8387;
  wire AES_CORE_DATAPATH__abc_16259_n8388;
  wire AES_CORE_DATAPATH__abc_16259_n8389;
  wire AES_CORE_DATAPATH__abc_16259_n8390;
  wire AES_CORE_DATAPATH__abc_16259_n8391;
  wire AES_CORE_DATAPATH__abc_16259_n8392;
  wire AES_CORE_DATAPATH__abc_16259_n8393;
  wire AES_CORE_DATAPATH__abc_16259_n8395;
  wire AES_CORE_DATAPATH__abc_16259_n8396;
  wire AES_CORE_DATAPATH__abc_16259_n8397;
  wire AES_CORE_DATAPATH__abc_16259_n8398;
  wire AES_CORE_DATAPATH__abc_16259_n8399;
  wire AES_CORE_DATAPATH__abc_16259_n8400;
  wire AES_CORE_DATAPATH__abc_16259_n8401;
  wire AES_CORE_DATAPATH__abc_16259_n8403;
  wire AES_CORE_DATAPATH__abc_16259_n8404;
  wire AES_CORE_DATAPATH__abc_16259_n8405;
  wire AES_CORE_DATAPATH__abc_16259_n8406;
  wire AES_CORE_DATAPATH__abc_16259_n8407;
  wire AES_CORE_DATAPATH__abc_16259_n8408;
  wire AES_CORE_DATAPATH__abc_16259_n8409;
  wire AES_CORE_DATAPATH__abc_16259_n8410;
  wire AES_CORE_DATAPATH__abc_16259_n8411;
  wire AES_CORE_DATAPATH__abc_16259_n8412;
  wire AES_CORE_DATAPATH__abc_16259_n8414;
  wire AES_CORE_DATAPATH__abc_16259_n8415;
  wire AES_CORE_DATAPATH__abc_16259_n8416;
  wire AES_CORE_DATAPATH__abc_16259_n8417;
  wire AES_CORE_DATAPATH__abc_16259_n8418;
  wire AES_CORE_DATAPATH__abc_16259_n8419;
  wire AES_CORE_DATAPATH__abc_16259_n8420;
  wire AES_CORE_DATAPATH__abc_16259_n8422;
  wire AES_CORE_DATAPATH__abc_16259_n8423;
  wire AES_CORE_DATAPATH__abc_16259_n8424;
  wire AES_CORE_DATAPATH__abc_16259_n8425;
  wire AES_CORE_DATAPATH__abc_16259_n8426;
  wire AES_CORE_DATAPATH__abc_16259_n8427;
  wire AES_CORE_DATAPATH__abc_16259_n8428;
  wire AES_CORE_DATAPATH__abc_16259_n8430;
  wire AES_CORE_DATAPATH__abc_16259_n8431;
  wire AES_CORE_DATAPATH__abc_16259_n8432;
  wire AES_CORE_DATAPATH__abc_16259_n8433;
  wire AES_CORE_DATAPATH__abc_16259_n8434;
  wire AES_CORE_DATAPATH__abc_16259_n8435;
  wire AES_CORE_DATAPATH__abc_16259_n8436;
  wire AES_CORE_DATAPATH__abc_16259_n8438;
  wire AES_CORE_DATAPATH__abc_16259_n8439;
  wire AES_CORE_DATAPATH__abc_16259_n8440;
  wire AES_CORE_DATAPATH__abc_16259_n8441;
  wire AES_CORE_DATAPATH__abc_16259_n8442;
  wire AES_CORE_DATAPATH__abc_16259_n8443;
  wire AES_CORE_DATAPATH__abc_16259_n8444;
  wire AES_CORE_DATAPATH__abc_16259_n8446;
  wire AES_CORE_DATAPATH__abc_16259_n8447;
  wire AES_CORE_DATAPATH__abc_16259_n8448;
  wire AES_CORE_DATAPATH__abc_16259_n8449;
  wire AES_CORE_DATAPATH__abc_16259_n8450;
  wire AES_CORE_DATAPATH__abc_16259_n8451;
  wire AES_CORE_DATAPATH__abc_16259_n8452;
  wire AES_CORE_DATAPATH__abc_16259_n8454;
  wire AES_CORE_DATAPATH__abc_16259_n8455;
  wire AES_CORE_DATAPATH__abc_16259_n8456;
  wire AES_CORE_DATAPATH__abc_16259_n8457;
  wire AES_CORE_DATAPATH__abc_16259_n8458;
  wire AES_CORE_DATAPATH__abc_16259_n8459;
  wire AES_CORE_DATAPATH__abc_16259_n8460;
  wire AES_CORE_DATAPATH__abc_16259_n8462;
  wire AES_CORE_DATAPATH__abc_16259_n8463;
  wire AES_CORE_DATAPATH__abc_16259_n8464;
  wire AES_CORE_DATAPATH__abc_16259_n8465;
  wire AES_CORE_DATAPATH__abc_16259_n8466;
  wire AES_CORE_DATAPATH__abc_16259_n8467;
  wire AES_CORE_DATAPATH__abc_16259_n8468;
  wire AES_CORE_DATAPATH__abc_16259_n8470;
  wire AES_CORE_DATAPATH__abc_16259_n8471;
  wire AES_CORE_DATAPATH__abc_16259_n8472;
  wire AES_CORE_DATAPATH__abc_16259_n8473;
  wire AES_CORE_DATAPATH__abc_16259_n8474;
  wire AES_CORE_DATAPATH__abc_16259_n8475;
  wire AES_CORE_DATAPATH__abc_16259_n8476;
  wire AES_CORE_DATAPATH__abc_16259_n8478;
  wire AES_CORE_DATAPATH__abc_16259_n8479;
  wire AES_CORE_DATAPATH__abc_16259_n8480;
  wire AES_CORE_DATAPATH__abc_16259_n8481;
  wire AES_CORE_DATAPATH__abc_16259_n8482;
  wire AES_CORE_DATAPATH__abc_16259_n8483;
  wire AES_CORE_DATAPATH__abc_16259_n8484;
  wire AES_CORE_DATAPATH__abc_16259_n8486;
  wire AES_CORE_DATAPATH__abc_16259_n8487;
  wire AES_CORE_DATAPATH__abc_16259_n8488;
  wire AES_CORE_DATAPATH__abc_16259_n8489;
  wire AES_CORE_DATAPATH__abc_16259_n8490;
  wire AES_CORE_DATAPATH__abc_16259_n8491;
  wire AES_CORE_DATAPATH__abc_16259_n8492;
  wire AES_CORE_DATAPATH__abc_16259_n8494;
  wire AES_CORE_DATAPATH__abc_16259_n8495;
  wire AES_CORE_DATAPATH__abc_16259_n8496;
  wire AES_CORE_DATAPATH__abc_16259_n8496_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n8496_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n8496_bF_buf10;
  wire AES_CORE_DATAPATH__abc_16259_n8496_bF_buf11;
  wire AES_CORE_DATAPATH__abc_16259_n8496_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n8496_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n8496_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n8496_bF_buf5;
  wire AES_CORE_DATAPATH__abc_16259_n8496_bF_buf6;
  wire AES_CORE_DATAPATH__abc_16259_n8496_bF_buf7;
  wire AES_CORE_DATAPATH__abc_16259_n8496_bF_buf8;
  wire AES_CORE_DATAPATH__abc_16259_n8496_bF_buf9;
  wire AES_CORE_DATAPATH__abc_16259_n8497;
  wire AES_CORE_DATAPATH__abc_16259_n8498;
  wire AES_CORE_DATAPATH__abc_16259_n8499;
  wire AES_CORE_DATAPATH__abc_16259_n8499_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n8499_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n8499_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n8499_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n8499_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n8499_bF_buf5;
  wire AES_CORE_DATAPATH__abc_16259_n8499_bF_buf6;
  wire AES_CORE_DATAPATH__abc_16259_n8499_bF_buf7;
  wire AES_CORE_DATAPATH__abc_16259_n8500;
  wire AES_CORE_DATAPATH__abc_16259_n8500_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n8500_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n8500_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n8500_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n8500_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n8500_bF_buf5;
  wire AES_CORE_DATAPATH__abc_16259_n8500_bF_buf6;
  wire AES_CORE_DATAPATH__abc_16259_n8501;
  wire AES_CORE_DATAPATH__abc_16259_n8502;
  wire AES_CORE_DATAPATH__abc_16259_n8504;
  wire AES_CORE_DATAPATH__abc_16259_n8505;
  wire AES_CORE_DATAPATH__abc_16259_n8507;
  wire AES_CORE_DATAPATH__abc_16259_n8508;
  wire AES_CORE_DATAPATH__abc_16259_n8510;
  wire AES_CORE_DATAPATH__abc_16259_n8511;
  wire AES_CORE_DATAPATH__abc_16259_n8513;
  wire AES_CORE_DATAPATH__abc_16259_n8514;
  wire AES_CORE_DATAPATH__abc_16259_n8516;
  wire AES_CORE_DATAPATH__abc_16259_n8517;
  wire AES_CORE_DATAPATH__abc_16259_n8519;
  wire AES_CORE_DATAPATH__abc_16259_n8520;
  wire AES_CORE_DATAPATH__abc_16259_n8522;
  wire AES_CORE_DATAPATH__abc_16259_n8523;
  wire AES_CORE_DATAPATH__abc_16259_n8525;
  wire AES_CORE_DATAPATH__abc_16259_n8526;
  wire AES_CORE_DATAPATH__abc_16259_n8528;
  wire AES_CORE_DATAPATH__abc_16259_n8529;
  wire AES_CORE_DATAPATH__abc_16259_n8531;
  wire AES_CORE_DATAPATH__abc_16259_n8532;
  wire AES_CORE_DATAPATH__abc_16259_n8533;
  wire AES_CORE_DATAPATH__abc_16259_n8535;
  wire AES_CORE_DATAPATH__abc_16259_n8536;
  wire AES_CORE_DATAPATH__abc_16259_n8537;
  wire AES_CORE_DATAPATH__abc_16259_n8539;
  wire AES_CORE_DATAPATH__abc_16259_n8540;
  wire AES_CORE_DATAPATH__abc_16259_n8542;
  wire AES_CORE_DATAPATH__abc_16259_n8543;
  wire AES_CORE_DATAPATH__abc_16259_n8544;
  wire AES_CORE_DATAPATH__abc_16259_n8546;
  wire AES_CORE_DATAPATH__abc_16259_n8547;
  wire AES_CORE_DATAPATH__abc_16259_n8549;
  wire AES_CORE_DATAPATH__abc_16259_n8550;
  wire AES_CORE_DATAPATH__abc_16259_n8551;
  wire AES_CORE_DATAPATH__abc_16259_n8553;
  wire AES_CORE_DATAPATH__abc_16259_n8554;
  wire AES_CORE_DATAPATH__abc_16259_n8556;
  wire AES_CORE_DATAPATH__abc_16259_n8557;
  wire AES_CORE_DATAPATH__abc_16259_n8558;
  wire AES_CORE_DATAPATH__abc_16259_n8560;
  wire AES_CORE_DATAPATH__abc_16259_n8561;
  wire AES_CORE_DATAPATH__abc_16259_n8563;
  wire AES_CORE_DATAPATH__abc_16259_n8564;
  wire AES_CORE_DATAPATH__abc_16259_n8566;
  wire AES_CORE_DATAPATH__abc_16259_n8567;
  wire AES_CORE_DATAPATH__abc_16259_n8569;
  wire AES_CORE_DATAPATH__abc_16259_n8570;
  wire AES_CORE_DATAPATH__abc_16259_n8571;
  wire AES_CORE_DATAPATH__abc_16259_n8573;
  wire AES_CORE_DATAPATH__abc_16259_n8574;
  wire AES_CORE_DATAPATH__abc_16259_n8576;
  wire AES_CORE_DATAPATH__abc_16259_n8577;
  wire AES_CORE_DATAPATH__abc_16259_n8579;
  wire AES_CORE_DATAPATH__abc_16259_n8580;
  wire AES_CORE_DATAPATH__abc_16259_n8582;
  wire AES_CORE_DATAPATH__abc_16259_n8583;
  wire AES_CORE_DATAPATH__abc_16259_n8585;
  wire AES_CORE_DATAPATH__abc_16259_n8586;
  wire AES_CORE_DATAPATH__abc_16259_n8588;
  wire AES_CORE_DATAPATH__abc_16259_n8589;
  wire AES_CORE_DATAPATH__abc_16259_n8591;
  wire AES_CORE_DATAPATH__abc_16259_n8592;
  wire AES_CORE_DATAPATH__abc_16259_n8594;
  wire AES_CORE_DATAPATH__abc_16259_n8595;
  wire AES_CORE_DATAPATH__abc_16259_n8597;
  wire AES_CORE_DATAPATH__abc_16259_n8598;
  wire AES_CORE_DATAPATH__abc_16259_n8600;
  wire AES_CORE_DATAPATH__abc_16259_n8601;
  wire AES_CORE_DATAPATH__abc_16259_n8603;
  wire AES_CORE_DATAPATH__abc_16259_n8603_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n8603_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n8603_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n8603_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n8603_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n8603_bF_buf5;
  wire AES_CORE_DATAPATH__abc_16259_n8603_bF_buf6;
  wire AES_CORE_DATAPATH__abc_16259_n8603_bF_buf7;
  wire AES_CORE_DATAPATH__abc_16259_n8603_bF_buf8;
  wire AES_CORE_DATAPATH__abc_16259_n8603_bF_buf9;
  wire AES_CORE_DATAPATH__abc_16259_n8604;
  wire AES_CORE_DATAPATH__abc_16259_n8605;
  wire AES_CORE_DATAPATH__abc_16259_n8606;
  wire AES_CORE_DATAPATH__abc_16259_n8607;
  wire AES_CORE_DATAPATH__abc_16259_n8608;
  wire AES_CORE_DATAPATH__abc_16259_n8609;
  wire AES_CORE_DATAPATH__abc_16259_n8610;
  wire AES_CORE_DATAPATH__abc_16259_n8611;
  wire AES_CORE_DATAPATH__abc_16259_n8613;
  wire AES_CORE_DATAPATH__abc_16259_n8614;
  wire AES_CORE_DATAPATH__abc_16259_n8615;
  wire AES_CORE_DATAPATH__abc_16259_n8616;
  wire AES_CORE_DATAPATH__abc_16259_n8617;
  wire AES_CORE_DATAPATH__abc_16259_n8618;
  wire AES_CORE_DATAPATH__abc_16259_n8619;
  wire AES_CORE_DATAPATH__abc_16259_n8620;
  wire AES_CORE_DATAPATH__abc_16259_n8622;
  wire AES_CORE_DATAPATH__abc_16259_n8623;
  wire AES_CORE_DATAPATH__abc_16259_n8624;
  wire AES_CORE_DATAPATH__abc_16259_n8625;
  wire AES_CORE_DATAPATH__abc_16259_n8626;
  wire AES_CORE_DATAPATH__abc_16259_n8627;
  wire AES_CORE_DATAPATH__abc_16259_n8628;
  wire AES_CORE_DATAPATH__abc_16259_n8629;
  wire AES_CORE_DATAPATH__abc_16259_n8631;
  wire AES_CORE_DATAPATH__abc_16259_n8632;
  wire AES_CORE_DATAPATH__abc_16259_n8633;
  wire AES_CORE_DATAPATH__abc_16259_n8634;
  wire AES_CORE_DATAPATH__abc_16259_n8635;
  wire AES_CORE_DATAPATH__abc_16259_n8636;
  wire AES_CORE_DATAPATH__abc_16259_n8637;
  wire AES_CORE_DATAPATH__abc_16259_n8638;
  wire AES_CORE_DATAPATH__abc_16259_n8640;
  wire AES_CORE_DATAPATH__abc_16259_n8641;
  wire AES_CORE_DATAPATH__abc_16259_n8642;
  wire AES_CORE_DATAPATH__abc_16259_n8643;
  wire AES_CORE_DATAPATH__abc_16259_n8644;
  wire AES_CORE_DATAPATH__abc_16259_n8645;
  wire AES_CORE_DATAPATH__abc_16259_n8646;
  wire AES_CORE_DATAPATH__abc_16259_n8647;
  wire AES_CORE_DATAPATH__abc_16259_n8649;
  wire AES_CORE_DATAPATH__abc_16259_n8650;
  wire AES_CORE_DATAPATH__abc_16259_n8651;
  wire AES_CORE_DATAPATH__abc_16259_n8652;
  wire AES_CORE_DATAPATH__abc_16259_n8653;
  wire AES_CORE_DATAPATH__abc_16259_n8654;
  wire AES_CORE_DATAPATH__abc_16259_n8655;
  wire AES_CORE_DATAPATH__abc_16259_n8656;
  wire AES_CORE_DATAPATH__abc_16259_n8658;
  wire AES_CORE_DATAPATH__abc_16259_n8659;
  wire AES_CORE_DATAPATH__abc_16259_n8660;
  wire AES_CORE_DATAPATH__abc_16259_n8661;
  wire AES_CORE_DATAPATH__abc_16259_n8662;
  wire AES_CORE_DATAPATH__abc_16259_n8663;
  wire AES_CORE_DATAPATH__abc_16259_n8664;
  wire AES_CORE_DATAPATH__abc_16259_n8665;
  wire AES_CORE_DATAPATH__abc_16259_n8667;
  wire AES_CORE_DATAPATH__abc_16259_n8668;
  wire AES_CORE_DATAPATH__abc_16259_n8669;
  wire AES_CORE_DATAPATH__abc_16259_n8670;
  wire AES_CORE_DATAPATH__abc_16259_n8671;
  wire AES_CORE_DATAPATH__abc_16259_n8672;
  wire AES_CORE_DATAPATH__abc_16259_n8673;
  wire AES_CORE_DATAPATH__abc_16259_n8674;
  wire AES_CORE_DATAPATH__abc_16259_n8676;
  wire AES_CORE_DATAPATH__abc_16259_n8677;
  wire AES_CORE_DATAPATH__abc_16259_n8678;
  wire AES_CORE_DATAPATH__abc_16259_n8679;
  wire AES_CORE_DATAPATH__abc_16259_n8680;
  wire AES_CORE_DATAPATH__abc_16259_n8681;
  wire AES_CORE_DATAPATH__abc_16259_n8682;
  wire AES_CORE_DATAPATH__abc_16259_n8683;
  wire AES_CORE_DATAPATH__abc_16259_n8685;
  wire AES_CORE_DATAPATH__abc_16259_n8686;
  wire AES_CORE_DATAPATH__abc_16259_n8687;
  wire AES_CORE_DATAPATH__abc_16259_n8688;
  wire AES_CORE_DATAPATH__abc_16259_n8689;
  wire AES_CORE_DATAPATH__abc_16259_n8690;
  wire AES_CORE_DATAPATH__abc_16259_n8691;
  wire AES_CORE_DATAPATH__abc_16259_n8692;
  wire AES_CORE_DATAPATH__abc_16259_n8694;
  wire AES_CORE_DATAPATH__abc_16259_n8695;
  wire AES_CORE_DATAPATH__abc_16259_n8696;
  wire AES_CORE_DATAPATH__abc_16259_n8697;
  wire AES_CORE_DATAPATH__abc_16259_n8698;
  wire AES_CORE_DATAPATH__abc_16259_n8699;
  wire AES_CORE_DATAPATH__abc_16259_n8700;
  wire AES_CORE_DATAPATH__abc_16259_n8701;
  wire AES_CORE_DATAPATH__abc_16259_n8702;
  wire AES_CORE_DATAPATH__abc_16259_n8704;
  wire AES_CORE_DATAPATH__abc_16259_n8705;
  wire AES_CORE_DATAPATH__abc_16259_n8706;
  wire AES_CORE_DATAPATH__abc_16259_n8707;
  wire AES_CORE_DATAPATH__abc_16259_n8708;
  wire AES_CORE_DATAPATH__abc_16259_n8709;
  wire AES_CORE_DATAPATH__abc_16259_n8710;
  wire AES_CORE_DATAPATH__abc_16259_n8711;
  wire AES_CORE_DATAPATH__abc_16259_n8712;
  wire AES_CORE_DATAPATH__abc_16259_n8714;
  wire AES_CORE_DATAPATH__abc_16259_n8715;
  wire AES_CORE_DATAPATH__abc_16259_n8716;
  wire AES_CORE_DATAPATH__abc_16259_n8717;
  wire AES_CORE_DATAPATH__abc_16259_n8718;
  wire AES_CORE_DATAPATH__abc_16259_n8719;
  wire AES_CORE_DATAPATH__abc_16259_n8720;
  wire AES_CORE_DATAPATH__abc_16259_n8721;
  wire AES_CORE_DATAPATH__abc_16259_n8723;
  wire AES_CORE_DATAPATH__abc_16259_n8724;
  wire AES_CORE_DATAPATH__abc_16259_n8725;
  wire AES_CORE_DATAPATH__abc_16259_n8726;
  wire AES_CORE_DATAPATH__abc_16259_n8727;
  wire AES_CORE_DATAPATH__abc_16259_n8728;
  wire AES_CORE_DATAPATH__abc_16259_n8729;
  wire AES_CORE_DATAPATH__abc_16259_n8730;
  wire AES_CORE_DATAPATH__abc_16259_n8731;
  wire AES_CORE_DATAPATH__abc_16259_n8733;
  wire AES_CORE_DATAPATH__abc_16259_n8734;
  wire AES_CORE_DATAPATH__abc_16259_n8735;
  wire AES_CORE_DATAPATH__abc_16259_n8736;
  wire AES_CORE_DATAPATH__abc_16259_n8737;
  wire AES_CORE_DATAPATH__abc_16259_n8738;
  wire AES_CORE_DATAPATH__abc_16259_n8739;
  wire AES_CORE_DATAPATH__abc_16259_n8740;
  wire AES_CORE_DATAPATH__abc_16259_n8742;
  wire AES_CORE_DATAPATH__abc_16259_n8743;
  wire AES_CORE_DATAPATH__abc_16259_n8744;
  wire AES_CORE_DATAPATH__abc_16259_n8745;
  wire AES_CORE_DATAPATH__abc_16259_n8746;
  wire AES_CORE_DATAPATH__abc_16259_n8747;
  wire AES_CORE_DATAPATH__abc_16259_n8748;
  wire AES_CORE_DATAPATH__abc_16259_n8749;
  wire AES_CORE_DATAPATH__abc_16259_n8750;
  wire AES_CORE_DATAPATH__abc_16259_n8752;
  wire AES_CORE_DATAPATH__abc_16259_n8753;
  wire AES_CORE_DATAPATH__abc_16259_n8754;
  wire AES_CORE_DATAPATH__abc_16259_n8755;
  wire AES_CORE_DATAPATH__abc_16259_n8756;
  wire AES_CORE_DATAPATH__abc_16259_n8757;
  wire AES_CORE_DATAPATH__abc_16259_n8758;
  wire AES_CORE_DATAPATH__abc_16259_n8759;
  wire AES_CORE_DATAPATH__abc_16259_n8761;
  wire AES_CORE_DATAPATH__abc_16259_n8762;
  wire AES_CORE_DATAPATH__abc_16259_n8763;
  wire AES_CORE_DATAPATH__abc_16259_n8764;
  wire AES_CORE_DATAPATH__abc_16259_n8765;
  wire AES_CORE_DATAPATH__abc_16259_n8766;
  wire AES_CORE_DATAPATH__abc_16259_n8767;
  wire AES_CORE_DATAPATH__abc_16259_n8768;
  wire AES_CORE_DATAPATH__abc_16259_n8769;
  wire AES_CORE_DATAPATH__abc_16259_n8771;
  wire AES_CORE_DATAPATH__abc_16259_n8772;
  wire AES_CORE_DATAPATH__abc_16259_n8773;
  wire AES_CORE_DATAPATH__abc_16259_n8774;
  wire AES_CORE_DATAPATH__abc_16259_n8775;
  wire AES_CORE_DATAPATH__abc_16259_n8776;
  wire AES_CORE_DATAPATH__abc_16259_n8777;
  wire AES_CORE_DATAPATH__abc_16259_n8778;
  wire AES_CORE_DATAPATH__abc_16259_n8780;
  wire AES_CORE_DATAPATH__abc_16259_n8781;
  wire AES_CORE_DATAPATH__abc_16259_n8782;
  wire AES_CORE_DATAPATH__abc_16259_n8783;
  wire AES_CORE_DATAPATH__abc_16259_n8784;
  wire AES_CORE_DATAPATH__abc_16259_n8785;
  wire AES_CORE_DATAPATH__abc_16259_n8786;
  wire AES_CORE_DATAPATH__abc_16259_n8787;
  wire AES_CORE_DATAPATH__abc_16259_n8789;
  wire AES_CORE_DATAPATH__abc_16259_n8790;
  wire AES_CORE_DATAPATH__abc_16259_n8791;
  wire AES_CORE_DATAPATH__abc_16259_n8792;
  wire AES_CORE_DATAPATH__abc_16259_n8793;
  wire AES_CORE_DATAPATH__abc_16259_n8794;
  wire AES_CORE_DATAPATH__abc_16259_n8795;
  wire AES_CORE_DATAPATH__abc_16259_n8796;
  wire AES_CORE_DATAPATH__abc_16259_n8798;
  wire AES_CORE_DATAPATH__abc_16259_n8799;
  wire AES_CORE_DATAPATH__abc_16259_n8800;
  wire AES_CORE_DATAPATH__abc_16259_n8801;
  wire AES_CORE_DATAPATH__abc_16259_n8802;
  wire AES_CORE_DATAPATH__abc_16259_n8803;
  wire AES_CORE_DATAPATH__abc_16259_n8804;
  wire AES_CORE_DATAPATH__abc_16259_n8805;
  wire AES_CORE_DATAPATH__abc_16259_n8806;
  wire AES_CORE_DATAPATH__abc_16259_n8808;
  wire AES_CORE_DATAPATH__abc_16259_n8809;
  wire AES_CORE_DATAPATH__abc_16259_n8810;
  wire AES_CORE_DATAPATH__abc_16259_n8811;
  wire AES_CORE_DATAPATH__abc_16259_n8812;
  wire AES_CORE_DATAPATH__abc_16259_n8813;
  wire AES_CORE_DATAPATH__abc_16259_n8814;
  wire AES_CORE_DATAPATH__abc_16259_n8815;
  wire AES_CORE_DATAPATH__abc_16259_n8817;
  wire AES_CORE_DATAPATH__abc_16259_n8818;
  wire AES_CORE_DATAPATH__abc_16259_n8819;
  wire AES_CORE_DATAPATH__abc_16259_n8820;
  wire AES_CORE_DATAPATH__abc_16259_n8821;
  wire AES_CORE_DATAPATH__abc_16259_n8822;
  wire AES_CORE_DATAPATH__abc_16259_n8823;
  wire AES_CORE_DATAPATH__abc_16259_n8824;
  wire AES_CORE_DATAPATH__abc_16259_n8826;
  wire AES_CORE_DATAPATH__abc_16259_n8827;
  wire AES_CORE_DATAPATH__abc_16259_n8828;
  wire AES_CORE_DATAPATH__abc_16259_n8829;
  wire AES_CORE_DATAPATH__abc_16259_n8830;
  wire AES_CORE_DATAPATH__abc_16259_n8831;
  wire AES_CORE_DATAPATH__abc_16259_n8832;
  wire AES_CORE_DATAPATH__abc_16259_n8833;
  wire AES_CORE_DATAPATH__abc_16259_n8835;
  wire AES_CORE_DATAPATH__abc_16259_n8836;
  wire AES_CORE_DATAPATH__abc_16259_n8837;
  wire AES_CORE_DATAPATH__abc_16259_n8838;
  wire AES_CORE_DATAPATH__abc_16259_n8839;
  wire AES_CORE_DATAPATH__abc_16259_n8840;
  wire AES_CORE_DATAPATH__abc_16259_n8841;
  wire AES_CORE_DATAPATH__abc_16259_n8842;
  wire AES_CORE_DATAPATH__abc_16259_n8844;
  wire AES_CORE_DATAPATH__abc_16259_n8845;
  wire AES_CORE_DATAPATH__abc_16259_n8846;
  wire AES_CORE_DATAPATH__abc_16259_n8847;
  wire AES_CORE_DATAPATH__abc_16259_n8848;
  wire AES_CORE_DATAPATH__abc_16259_n8849;
  wire AES_CORE_DATAPATH__abc_16259_n8850;
  wire AES_CORE_DATAPATH__abc_16259_n8851;
  wire AES_CORE_DATAPATH__abc_16259_n8853;
  wire AES_CORE_DATAPATH__abc_16259_n8854;
  wire AES_CORE_DATAPATH__abc_16259_n8855;
  wire AES_CORE_DATAPATH__abc_16259_n8856;
  wire AES_CORE_DATAPATH__abc_16259_n8857;
  wire AES_CORE_DATAPATH__abc_16259_n8858;
  wire AES_CORE_DATAPATH__abc_16259_n8859;
  wire AES_CORE_DATAPATH__abc_16259_n8860;
  wire AES_CORE_DATAPATH__abc_16259_n8862;
  wire AES_CORE_DATAPATH__abc_16259_n8863;
  wire AES_CORE_DATAPATH__abc_16259_n8864;
  wire AES_CORE_DATAPATH__abc_16259_n8865;
  wire AES_CORE_DATAPATH__abc_16259_n8866;
  wire AES_CORE_DATAPATH__abc_16259_n8867;
  wire AES_CORE_DATAPATH__abc_16259_n8868;
  wire AES_CORE_DATAPATH__abc_16259_n8869;
  wire AES_CORE_DATAPATH__abc_16259_n8871;
  wire AES_CORE_DATAPATH__abc_16259_n8872;
  wire AES_CORE_DATAPATH__abc_16259_n8873;
  wire AES_CORE_DATAPATH__abc_16259_n8874;
  wire AES_CORE_DATAPATH__abc_16259_n8875;
  wire AES_CORE_DATAPATH__abc_16259_n8876;
  wire AES_CORE_DATAPATH__abc_16259_n8877;
  wire AES_CORE_DATAPATH__abc_16259_n8878;
  wire AES_CORE_DATAPATH__abc_16259_n8880;
  wire AES_CORE_DATAPATH__abc_16259_n8881;
  wire AES_CORE_DATAPATH__abc_16259_n8882;
  wire AES_CORE_DATAPATH__abc_16259_n8883;
  wire AES_CORE_DATAPATH__abc_16259_n8884;
  wire AES_CORE_DATAPATH__abc_16259_n8885;
  wire AES_CORE_DATAPATH__abc_16259_n8886;
  wire AES_CORE_DATAPATH__abc_16259_n8887;
  wire AES_CORE_DATAPATH__abc_16259_n8889;
  wire AES_CORE_DATAPATH__abc_16259_n8890;
  wire AES_CORE_DATAPATH__abc_16259_n8891;
  wire AES_CORE_DATAPATH__abc_16259_n8892;
  wire AES_CORE_DATAPATH__abc_16259_n8893;
  wire AES_CORE_DATAPATH__abc_16259_n8894;
  wire AES_CORE_DATAPATH__abc_16259_n8895;
  wire AES_CORE_DATAPATH__abc_16259_n8896;
  wire AES_CORE_DATAPATH__abc_16259_n8898;
  wire AES_CORE_DATAPATH__abc_16259_n8898_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n8898_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n8898_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n8898_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n8898_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n8899;
  wire AES_CORE_DATAPATH__abc_16259_n8899_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n8899_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n8899_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n8899_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n8899_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n8900;
  wire AES_CORE_DATAPATH__abc_16259_n8900_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n8900_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n8900_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n8900_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n8901;
  wire AES_CORE_DATAPATH__abc_16259_n8902;
  wire AES_CORE_DATAPATH__abc_16259_n8903;
  wire AES_CORE_DATAPATH__abc_16259_n8904;
  wire AES_CORE_DATAPATH__abc_16259_n8905;
  wire AES_CORE_DATAPATH__abc_16259_n8905_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n8905_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n8905_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n8905_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n8905_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n8906;
  wire AES_CORE_DATAPATH__abc_16259_n8907;
  wire AES_CORE_DATAPATH__abc_16259_n8908;
  wire AES_CORE_DATAPATH__abc_16259_n8909;
  wire AES_CORE_DATAPATH__abc_16259_n8911;
  wire AES_CORE_DATAPATH__abc_16259_n8912;
  wire AES_CORE_DATAPATH__abc_16259_n8913;
  wire AES_CORE_DATAPATH__abc_16259_n8914;
  wire AES_CORE_DATAPATH__abc_16259_n8915;
  wire AES_CORE_DATAPATH__abc_16259_n8916;
  wire AES_CORE_DATAPATH__abc_16259_n8917;
  wire AES_CORE_DATAPATH__abc_16259_n8918;
  wire AES_CORE_DATAPATH__abc_16259_n8918_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n8918_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n8918_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n8918_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n8918_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n8919;
  wire AES_CORE_DATAPATH__abc_16259_n8920;
  wire AES_CORE_DATAPATH__abc_16259_n8921;
  wire AES_CORE_DATAPATH__abc_16259_n8922;
  wire AES_CORE_DATAPATH__abc_16259_n8924;
  wire AES_CORE_DATAPATH__abc_16259_n8925;
  wire AES_CORE_DATAPATH__abc_16259_n8926;
  wire AES_CORE_DATAPATH__abc_16259_n8927;
  wire AES_CORE_DATAPATH__abc_16259_n8928;
  wire AES_CORE_DATAPATH__abc_16259_n8929;
  wire AES_CORE_DATAPATH__abc_16259_n8930;
  wire AES_CORE_DATAPATH__abc_16259_n8931;
  wire AES_CORE_DATAPATH__abc_16259_n8932;
  wire AES_CORE_DATAPATH__abc_16259_n8934;
  wire AES_CORE_DATAPATH__abc_16259_n8935;
  wire AES_CORE_DATAPATH__abc_16259_n8936;
  wire AES_CORE_DATAPATH__abc_16259_n8937;
  wire AES_CORE_DATAPATH__abc_16259_n8938;
  wire AES_CORE_DATAPATH__abc_16259_n8939;
  wire AES_CORE_DATAPATH__abc_16259_n8940;
  wire AES_CORE_DATAPATH__abc_16259_n8941;
  wire AES_CORE_DATAPATH__abc_16259_n8942;
  wire AES_CORE_DATAPATH__abc_16259_n8943;
  wire AES_CORE_DATAPATH__abc_16259_n8944;
  wire AES_CORE_DATAPATH__abc_16259_n8946;
  wire AES_CORE_DATAPATH__abc_16259_n8947;
  wire AES_CORE_DATAPATH__abc_16259_n8948;
  wire AES_CORE_DATAPATH__abc_16259_n8949;
  wire AES_CORE_DATAPATH__abc_16259_n8950;
  wire AES_CORE_DATAPATH__abc_16259_n8951;
  wire AES_CORE_DATAPATH__abc_16259_n8952;
  wire AES_CORE_DATAPATH__abc_16259_n8953;
  wire AES_CORE_DATAPATH__abc_16259_n8954;
  wire AES_CORE_DATAPATH__abc_16259_n8956;
  wire AES_CORE_DATAPATH__abc_16259_n8957;
  wire AES_CORE_DATAPATH__abc_16259_n8958;
  wire AES_CORE_DATAPATH__abc_16259_n8959;
  wire AES_CORE_DATAPATH__abc_16259_n8960;
  wire AES_CORE_DATAPATH__abc_16259_n8961;
  wire AES_CORE_DATAPATH__abc_16259_n8962;
  wire AES_CORE_DATAPATH__abc_16259_n8963;
  wire AES_CORE_DATAPATH__abc_16259_n8964;
  wire AES_CORE_DATAPATH__abc_16259_n8965;
  wire AES_CORE_DATAPATH__abc_16259_n8967;
  wire AES_CORE_DATAPATH__abc_16259_n8968;
  wire AES_CORE_DATAPATH__abc_16259_n8969;
  wire AES_CORE_DATAPATH__abc_16259_n8970;
  wire AES_CORE_DATAPATH__abc_16259_n8971;
  wire AES_CORE_DATAPATH__abc_16259_n8972;
  wire AES_CORE_DATAPATH__abc_16259_n8973;
  wire AES_CORE_DATAPATH__abc_16259_n8974;
  wire AES_CORE_DATAPATH__abc_16259_n8975;
  wire AES_CORE_DATAPATH__abc_16259_n8977;
  wire AES_CORE_DATAPATH__abc_16259_n8978;
  wire AES_CORE_DATAPATH__abc_16259_n8979;
  wire AES_CORE_DATAPATH__abc_16259_n8980;
  wire AES_CORE_DATAPATH__abc_16259_n8981;
  wire AES_CORE_DATAPATH__abc_16259_n8982;
  wire AES_CORE_DATAPATH__abc_16259_n8983;
  wire AES_CORE_DATAPATH__abc_16259_n8984;
  wire AES_CORE_DATAPATH__abc_16259_n8985;
  wire AES_CORE_DATAPATH__abc_16259_n8986;
  wire AES_CORE_DATAPATH__abc_16259_n8987;
  wire AES_CORE_DATAPATH__abc_16259_n8989;
  wire AES_CORE_DATAPATH__abc_16259_n8990;
  wire AES_CORE_DATAPATH__abc_16259_n8991;
  wire AES_CORE_DATAPATH__abc_16259_n8992;
  wire AES_CORE_DATAPATH__abc_16259_n8993;
  wire AES_CORE_DATAPATH__abc_16259_n8994;
  wire AES_CORE_DATAPATH__abc_16259_n8995;
  wire AES_CORE_DATAPATH__abc_16259_n8996;
  wire AES_CORE_DATAPATH__abc_16259_n8997;
  wire AES_CORE_DATAPATH__abc_16259_n8999;
  wire AES_CORE_DATAPATH__abc_16259_n9000;
  wire AES_CORE_DATAPATH__abc_16259_n9001;
  wire AES_CORE_DATAPATH__abc_16259_n9002;
  wire AES_CORE_DATAPATH__abc_16259_n9003;
  wire AES_CORE_DATAPATH__abc_16259_n9004;
  wire AES_CORE_DATAPATH__abc_16259_n9005;
  wire AES_CORE_DATAPATH__abc_16259_n9006;
  wire AES_CORE_DATAPATH__abc_16259_n9007;
  wire AES_CORE_DATAPATH__abc_16259_n9008;
  wire AES_CORE_DATAPATH__abc_16259_n9009;
  wire AES_CORE_DATAPATH__abc_16259_n9010;
  wire AES_CORE_DATAPATH__abc_16259_n9012;
  wire AES_CORE_DATAPATH__abc_16259_n9013;
  wire AES_CORE_DATAPATH__abc_16259_n9014;
  wire AES_CORE_DATAPATH__abc_16259_n9015;
  wire AES_CORE_DATAPATH__abc_16259_n9016;
  wire AES_CORE_DATAPATH__abc_16259_n9017;
  wire AES_CORE_DATAPATH__abc_16259_n9018;
  wire AES_CORE_DATAPATH__abc_16259_n9019;
  wire AES_CORE_DATAPATH__abc_16259_n9020;
  wire AES_CORE_DATAPATH__abc_16259_n9021;
  wire AES_CORE_DATAPATH__abc_16259_n9022;
  wire AES_CORE_DATAPATH__abc_16259_n9024;
  wire AES_CORE_DATAPATH__abc_16259_n9025;
  wire AES_CORE_DATAPATH__abc_16259_n9026;
  wire AES_CORE_DATAPATH__abc_16259_n9027;
  wire AES_CORE_DATAPATH__abc_16259_n9028;
  wire AES_CORE_DATAPATH__abc_16259_n9029;
  wire AES_CORE_DATAPATH__abc_16259_n9030;
  wire AES_CORE_DATAPATH__abc_16259_n9031;
  wire AES_CORE_DATAPATH__abc_16259_n9032;
  wire AES_CORE_DATAPATH__abc_16259_n9033;
  wire AES_CORE_DATAPATH__abc_16259_n9034;
  wire AES_CORE_DATAPATH__abc_16259_n9036;
  wire AES_CORE_DATAPATH__abc_16259_n9037;
  wire AES_CORE_DATAPATH__abc_16259_n9038;
  wire AES_CORE_DATAPATH__abc_16259_n9039;
  wire AES_CORE_DATAPATH__abc_16259_n9040;
  wire AES_CORE_DATAPATH__abc_16259_n9041;
  wire AES_CORE_DATAPATH__abc_16259_n9042;
  wire AES_CORE_DATAPATH__abc_16259_n9043;
  wire AES_CORE_DATAPATH__abc_16259_n9044;
  wire AES_CORE_DATAPATH__abc_16259_n9045;
  wire AES_CORE_DATAPATH__abc_16259_n9046;
  wire AES_CORE_DATAPATH__abc_16259_n9048;
  wire AES_CORE_DATAPATH__abc_16259_n9049;
  wire AES_CORE_DATAPATH__abc_16259_n9050;
  wire AES_CORE_DATAPATH__abc_16259_n9051;
  wire AES_CORE_DATAPATH__abc_16259_n9052;
  wire AES_CORE_DATAPATH__abc_16259_n9053;
  wire AES_CORE_DATAPATH__abc_16259_n9054;
  wire AES_CORE_DATAPATH__abc_16259_n9055;
  wire AES_CORE_DATAPATH__abc_16259_n9056;
  wire AES_CORE_DATAPATH__abc_16259_n9057;
  wire AES_CORE_DATAPATH__abc_16259_n9058;
  wire AES_CORE_DATAPATH__abc_16259_n9060;
  wire AES_CORE_DATAPATH__abc_16259_n9061;
  wire AES_CORE_DATAPATH__abc_16259_n9062;
  wire AES_CORE_DATAPATH__abc_16259_n9063;
  wire AES_CORE_DATAPATH__abc_16259_n9064;
  wire AES_CORE_DATAPATH__abc_16259_n9065;
  wire AES_CORE_DATAPATH__abc_16259_n9066;
  wire AES_CORE_DATAPATH__abc_16259_n9067;
  wire AES_CORE_DATAPATH__abc_16259_n9068;
  wire AES_CORE_DATAPATH__abc_16259_n9069;
  wire AES_CORE_DATAPATH__abc_16259_n9070;
  wire AES_CORE_DATAPATH__abc_16259_n9072;
  wire AES_CORE_DATAPATH__abc_16259_n9073;
  wire AES_CORE_DATAPATH__abc_16259_n9074;
  wire AES_CORE_DATAPATH__abc_16259_n9075;
  wire AES_CORE_DATAPATH__abc_16259_n9076;
  wire AES_CORE_DATAPATH__abc_16259_n9077;
  wire AES_CORE_DATAPATH__abc_16259_n9078;
  wire AES_CORE_DATAPATH__abc_16259_n9079;
  wire AES_CORE_DATAPATH__abc_16259_n9080;
  wire AES_CORE_DATAPATH__abc_16259_n9081;
  wire AES_CORE_DATAPATH__abc_16259_n9082;
  wire AES_CORE_DATAPATH__abc_16259_n9084;
  wire AES_CORE_DATAPATH__abc_16259_n9085;
  wire AES_CORE_DATAPATH__abc_16259_n9086;
  wire AES_CORE_DATAPATH__abc_16259_n9087;
  wire AES_CORE_DATAPATH__abc_16259_n9088;
  wire AES_CORE_DATAPATH__abc_16259_n9089;
  wire AES_CORE_DATAPATH__abc_16259_n9090;
  wire AES_CORE_DATAPATH__abc_16259_n9091;
  wire AES_CORE_DATAPATH__abc_16259_n9092;
  wire AES_CORE_DATAPATH__abc_16259_n9093;
  wire AES_CORE_DATAPATH__abc_16259_n9094;
  wire AES_CORE_DATAPATH__abc_16259_n9096;
  wire AES_CORE_DATAPATH__abc_16259_n9097;
  wire AES_CORE_DATAPATH__abc_16259_n9098;
  wire AES_CORE_DATAPATH__abc_16259_n9099;
  wire AES_CORE_DATAPATH__abc_16259_n9100;
  wire AES_CORE_DATAPATH__abc_16259_n9101;
  wire AES_CORE_DATAPATH__abc_16259_n9102;
  wire AES_CORE_DATAPATH__abc_16259_n9103;
  wire AES_CORE_DATAPATH__abc_16259_n9104;
  wire AES_CORE_DATAPATH__abc_16259_n9105;
  wire AES_CORE_DATAPATH__abc_16259_n9106;
  wire AES_CORE_DATAPATH__abc_16259_n9108;
  wire AES_CORE_DATAPATH__abc_16259_n9109;
  wire AES_CORE_DATAPATH__abc_16259_n9110;
  wire AES_CORE_DATAPATH__abc_16259_n9111;
  wire AES_CORE_DATAPATH__abc_16259_n9112;
  wire AES_CORE_DATAPATH__abc_16259_n9113;
  wire AES_CORE_DATAPATH__abc_16259_n9114;
  wire AES_CORE_DATAPATH__abc_16259_n9115;
  wire AES_CORE_DATAPATH__abc_16259_n9116;
  wire AES_CORE_DATAPATH__abc_16259_n9117;
  wire AES_CORE_DATAPATH__abc_16259_n9118;
  wire AES_CORE_DATAPATH__abc_16259_n9119;
  wire AES_CORE_DATAPATH__abc_16259_n9121;
  wire AES_CORE_DATAPATH__abc_16259_n9122;
  wire AES_CORE_DATAPATH__abc_16259_n9123;
  wire AES_CORE_DATAPATH__abc_16259_n9124;
  wire AES_CORE_DATAPATH__abc_16259_n9125;
  wire AES_CORE_DATAPATH__abc_16259_n9126;
  wire AES_CORE_DATAPATH__abc_16259_n9127;
  wire AES_CORE_DATAPATH__abc_16259_n9128;
  wire AES_CORE_DATAPATH__abc_16259_n9129;
  wire AES_CORE_DATAPATH__abc_16259_n9130;
  wire AES_CORE_DATAPATH__abc_16259_n9131;
  wire AES_CORE_DATAPATH__abc_16259_n9133;
  wire AES_CORE_DATAPATH__abc_16259_n9134;
  wire AES_CORE_DATAPATH__abc_16259_n9135;
  wire AES_CORE_DATAPATH__abc_16259_n9136;
  wire AES_CORE_DATAPATH__abc_16259_n9137;
  wire AES_CORE_DATAPATH__abc_16259_n9138;
  wire AES_CORE_DATAPATH__abc_16259_n9139;
  wire AES_CORE_DATAPATH__abc_16259_n9140;
  wire AES_CORE_DATAPATH__abc_16259_n9141;
  wire AES_CORE_DATAPATH__abc_16259_n9142;
  wire AES_CORE_DATAPATH__abc_16259_n9143;
  wire AES_CORE_DATAPATH__abc_16259_n9144;
  wire AES_CORE_DATAPATH__abc_16259_n9145;
  wire AES_CORE_DATAPATH__abc_16259_n9147;
  wire AES_CORE_DATAPATH__abc_16259_n9148;
  wire AES_CORE_DATAPATH__abc_16259_n9149;
  wire AES_CORE_DATAPATH__abc_16259_n9150;
  wire AES_CORE_DATAPATH__abc_16259_n9151;
  wire AES_CORE_DATAPATH__abc_16259_n9152;
  wire AES_CORE_DATAPATH__abc_16259_n9153;
  wire AES_CORE_DATAPATH__abc_16259_n9154;
  wire AES_CORE_DATAPATH__abc_16259_n9155;
  wire AES_CORE_DATAPATH__abc_16259_n9156;
  wire AES_CORE_DATAPATH__abc_16259_n9157;
  wire AES_CORE_DATAPATH__abc_16259_n9159;
  wire AES_CORE_DATAPATH__abc_16259_n9160;
  wire AES_CORE_DATAPATH__abc_16259_n9161;
  wire AES_CORE_DATAPATH__abc_16259_n9162;
  wire AES_CORE_DATAPATH__abc_16259_n9163;
  wire AES_CORE_DATAPATH__abc_16259_n9164;
  wire AES_CORE_DATAPATH__abc_16259_n9165;
  wire AES_CORE_DATAPATH__abc_16259_n9166;
  wire AES_CORE_DATAPATH__abc_16259_n9167;
  wire AES_CORE_DATAPATH__abc_16259_n9168;
  wire AES_CORE_DATAPATH__abc_16259_n9169;
  wire AES_CORE_DATAPATH__abc_16259_n9170;
  wire AES_CORE_DATAPATH__abc_16259_n9171;
  wire AES_CORE_DATAPATH__abc_16259_n9172;
  wire AES_CORE_DATAPATH__abc_16259_n9174;
  wire AES_CORE_DATAPATH__abc_16259_n9175;
  wire AES_CORE_DATAPATH__abc_16259_n9176;
  wire AES_CORE_DATAPATH__abc_16259_n9177;
  wire AES_CORE_DATAPATH__abc_16259_n9178;
  wire AES_CORE_DATAPATH__abc_16259_n9179;
  wire AES_CORE_DATAPATH__abc_16259_n9180;
  wire AES_CORE_DATAPATH__abc_16259_n9181;
  wire AES_CORE_DATAPATH__abc_16259_n9182;
  wire AES_CORE_DATAPATH__abc_16259_n9183;
  wire AES_CORE_DATAPATH__abc_16259_n9184;
  wire AES_CORE_DATAPATH__abc_16259_n9186;
  wire AES_CORE_DATAPATH__abc_16259_n9187;
  wire AES_CORE_DATAPATH__abc_16259_n9188;
  wire AES_CORE_DATAPATH__abc_16259_n9189;
  wire AES_CORE_DATAPATH__abc_16259_n9190;
  wire AES_CORE_DATAPATH__abc_16259_n9191;
  wire AES_CORE_DATAPATH__abc_16259_n9192;
  wire AES_CORE_DATAPATH__abc_16259_n9193;
  wire AES_CORE_DATAPATH__abc_16259_n9194;
  wire AES_CORE_DATAPATH__abc_16259_n9195;
  wire AES_CORE_DATAPATH__abc_16259_n9196;
  wire AES_CORE_DATAPATH__abc_16259_n9197;
  wire AES_CORE_DATAPATH__abc_16259_n9198;
  wire AES_CORE_DATAPATH__abc_16259_n9200;
  wire AES_CORE_DATAPATH__abc_16259_n9201;
  wire AES_CORE_DATAPATH__abc_16259_n9202;
  wire AES_CORE_DATAPATH__abc_16259_n9203;
  wire AES_CORE_DATAPATH__abc_16259_n9204;
  wire AES_CORE_DATAPATH__abc_16259_n9205;
  wire AES_CORE_DATAPATH__abc_16259_n9206;
  wire AES_CORE_DATAPATH__abc_16259_n9207;
  wire AES_CORE_DATAPATH__abc_16259_n9208;
  wire AES_CORE_DATAPATH__abc_16259_n9209;
  wire AES_CORE_DATAPATH__abc_16259_n9210;
  wire AES_CORE_DATAPATH__abc_16259_n9212;
  wire AES_CORE_DATAPATH__abc_16259_n9213;
  wire AES_CORE_DATAPATH__abc_16259_n9214;
  wire AES_CORE_DATAPATH__abc_16259_n9215;
  wire AES_CORE_DATAPATH__abc_16259_n9216;
  wire AES_CORE_DATAPATH__abc_16259_n9217;
  wire AES_CORE_DATAPATH__abc_16259_n9218;
  wire AES_CORE_DATAPATH__abc_16259_n9219;
  wire AES_CORE_DATAPATH__abc_16259_n9220;
  wire AES_CORE_DATAPATH__abc_16259_n9221;
  wire AES_CORE_DATAPATH__abc_16259_n9222;
  wire AES_CORE_DATAPATH__abc_16259_n9223;
  wire AES_CORE_DATAPATH__abc_16259_n9225;
  wire AES_CORE_DATAPATH__abc_16259_n9226;
  wire AES_CORE_DATAPATH__abc_16259_n9227;
  wire AES_CORE_DATAPATH__abc_16259_n9228;
  wire AES_CORE_DATAPATH__abc_16259_n9229;
  wire AES_CORE_DATAPATH__abc_16259_n9230;
  wire AES_CORE_DATAPATH__abc_16259_n9231;
  wire AES_CORE_DATAPATH__abc_16259_n9232;
  wire AES_CORE_DATAPATH__abc_16259_n9233;
  wire AES_CORE_DATAPATH__abc_16259_n9234;
  wire AES_CORE_DATAPATH__abc_16259_n9235;
  wire AES_CORE_DATAPATH__abc_16259_n9237;
  wire AES_CORE_DATAPATH__abc_16259_n9238;
  wire AES_CORE_DATAPATH__abc_16259_n9239;
  wire AES_CORE_DATAPATH__abc_16259_n9240;
  wire AES_CORE_DATAPATH__abc_16259_n9241;
  wire AES_CORE_DATAPATH__abc_16259_n9242;
  wire AES_CORE_DATAPATH__abc_16259_n9243;
  wire AES_CORE_DATAPATH__abc_16259_n9244;
  wire AES_CORE_DATAPATH__abc_16259_n9245;
  wire AES_CORE_DATAPATH__abc_16259_n9246;
  wire AES_CORE_DATAPATH__abc_16259_n9247;
  wire AES_CORE_DATAPATH__abc_16259_n9249;
  wire AES_CORE_DATAPATH__abc_16259_n9250;
  wire AES_CORE_DATAPATH__abc_16259_n9251;
  wire AES_CORE_DATAPATH__abc_16259_n9252;
  wire AES_CORE_DATAPATH__abc_16259_n9253;
  wire AES_CORE_DATAPATH__abc_16259_n9254;
  wire AES_CORE_DATAPATH__abc_16259_n9255;
  wire AES_CORE_DATAPATH__abc_16259_n9256;
  wire AES_CORE_DATAPATH__abc_16259_n9257;
  wire AES_CORE_DATAPATH__abc_16259_n9258;
  wire AES_CORE_DATAPATH__abc_16259_n9259;
  wire AES_CORE_DATAPATH__abc_16259_n9261;
  wire AES_CORE_DATAPATH__abc_16259_n9262;
  wire AES_CORE_DATAPATH__abc_16259_n9263;
  wire AES_CORE_DATAPATH__abc_16259_n9264;
  wire AES_CORE_DATAPATH__abc_16259_n9265;
  wire AES_CORE_DATAPATH__abc_16259_n9266;
  wire AES_CORE_DATAPATH__abc_16259_n9267;
  wire AES_CORE_DATAPATH__abc_16259_n9268;
  wire AES_CORE_DATAPATH__abc_16259_n9269;
  wire AES_CORE_DATAPATH__abc_16259_n9270;
  wire AES_CORE_DATAPATH__abc_16259_n9271;
  wire AES_CORE_DATAPATH__abc_16259_n9273;
  wire AES_CORE_DATAPATH__abc_16259_n9274;
  wire AES_CORE_DATAPATH__abc_16259_n9275;
  wire AES_CORE_DATAPATH__abc_16259_n9276;
  wire AES_CORE_DATAPATH__abc_16259_n9277;
  wire AES_CORE_DATAPATH__abc_16259_n9278;
  wire AES_CORE_DATAPATH__abc_16259_n9279;
  wire AES_CORE_DATAPATH__abc_16259_n9280;
  wire AES_CORE_DATAPATH__abc_16259_n9281;
  wire AES_CORE_DATAPATH__abc_16259_n9282;
  wire AES_CORE_DATAPATH__abc_16259_n9283;
  wire AES_CORE_DATAPATH__abc_16259_n9285;
  wire AES_CORE_DATAPATH__abc_16259_n9286;
  wire AES_CORE_DATAPATH__abc_16259_n9287;
  wire AES_CORE_DATAPATH__abc_16259_n9287_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n9287_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n9287_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n9287_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n9287_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n9287_bF_buf5;
  wire AES_CORE_DATAPATH__abc_16259_n9287_bF_buf6;
  wire AES_CORE_DATAPATH__abc_16259_n9287_bF_buf7;
  wire AES_CORE_DATAPATH__abc_16259_n9288;
  wire AES_CORE_DATAPATH__abc_16259_n9288_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n9288_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n9288_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n9288_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n9288_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n9288_bF_buf5;
  wire AES_CORE_DATAPATH__abc_16259_n9288_bF_buf6;
  wire AES_CORE_DATAPATH__abc_16259_n9289;
  wire AES_CORE_DATAPATH__abc_16259_n9290;
  wire AES_CORE_DATAPATH__abc_16259_n9292;
  wire AES_CORE_DATAPATH__abc_16259_n9293;
  wire AES_CORE_DATAPATH__abc_16259_n9295;
  wire AES_CORE_DATAPATH__abc_16259_n9296;
  wire AES_CORE_DATAPATH__abc_16259_n9298;
  wire AES_CORE_DATAPATH__abc_16259_n9299;
  wire AES_CORE_DATAPATH__abc_16259_n9301;
  wire AES_CORE_DATAPATH__abc_16259_n9302;
  wire AES_CORE_DATAPATH__abc_16259_n9304;
  wire AES_CORE_DATAPATH__abc_16259_n9305;
  wire AES_CORE_DATAPATH__abc_16259_n9307;
  wire AES_CORE_DATAPATH__abc_16259_n9308;
  wire AES_CORE_DATAPATH__abc_16259_n9310;
  wire AES_CORE_DATAPATH__abc_16259_n9311;
  wire AES_CORE_DATAPATH__abc_16259_n9313;
  wire AES_CORE_DATAPATH__abc_16259_n9314;
  wire AES_CORE_DATAPATH__abc_16259_n9316;
  wire AES_CORE_DATAPATH__abc_16259_n9317;
  wire AES_CORE_DATAPATH__abc_16259_n9319;
  wire AES_CORE_DATAPATH__abc_16259_n9320;
  wire AES_CORE_DATAPATH__abc_16259_n9321;
  wire AES_CORE_DATAPATH__abc_16259_n9323;
  wire AES_CORE_DATAPATH__abc_16259_n9324;
  wire AES_CORE_DATAPATH__abc_16259_n9325;
  wire AES_CORE_DATAPATH__abc_16259_n9327;
  wire AES_CORE_DATAPATH__abc_16259_n9328;
  wire AES_CORE_DATAPATH__abc_16259_n9330;
  wire AES_CORE_DATAPATH__abc_16259_n9331;
  wire AES_CORE_DATAPATH__abc_16259_n9332;
  wire AES_CORE_DATAPATH__abc_16259_n9334;
  wire AES_CORE_DATAPATH__abc_16259_n9335;
  wire AES_CORE_DATAPATH__abc_16259_n9337;
  wire AES_CORE_DATAPATH__abc_16259_n9338;
  wire AES_CORE_DATAPATH__abc_16259_n9339;
  wire AES_CORE_DATAPATH__abc_16259_n9341;
  wire AES_CORE_DATAPATH__abc_16259_n9342;
  wire AES_CORE_DATAPATH__abc_16259_n9344;
  wire AES_CORE_DATAPATH__abc_16259_n9345;
  wire AES_CORE_DATAPATH__abc_16259_n9346;
  wire AES_CORE_DATAPATH__abc_16259_n9348;
  wire AES_CORE_DATAPATH__abc_16259_n9349;
  wire AES_CORE_DATAPATH__abc_16259_n9351;
  wire AES_CORE_DATAPATH__abc_16259_n9352;
  wire AES_CORE_DATAPATH__abc_16259_n9354;
  wire AES_CORE_DATAPATH__abc_16259_n9355;
  wire AES_CORE_DATAPATH__abc_16259_n9357;
  wire AES_CORE_DATAPATH__abc_16259_n9358;
  wire AES_CORE_DATAPATH__abc_16259_n9359;
  wire AES_CORE_DATAPATH__abc_16259_n9361;
  wire AES_CORE_DATAPATH__abc_16259_n9362;
  wire AES_CORE_DATAPATH__abc_16259_n9364;
  wire AES_CORE_DATAPATH__abc_16259_n9365;
  wire AES_CORE_DATAPATH__abc_16259_n9367;
  wire AES_CORE_DATAPATH__abc_16259_n9368;
  wire AES_CORE_DATAPATH__abc_16259_n9370;
  wire AES_CORE_DATAPATH__abc_16259_n9371;
  wire AES_CORE_DATAPATH__abc_16259_n9373;
  wire AES_CORE_DATAPATH__abc_16259_n9374;
  wire AES_CORE_DATAPATH__abc_16259_n9376;
  wire AES_CORE_DATAPATH__abc_16259_n9377;
  wire AES_CORE_DATAPATH__abc_16259_n9379;
  wire AES_CORE_DATAPATH__abc_16259_n9380;
  wire AES_CORE_DATAPATH__abc_16259_n9382;
  wire AES_CORE_DATAPATH__abc_16259_n9383;
  wire AES_CORE_DATAPATH__abc_16259_n9385;
  wire AES_CORE_DATAPATH__abc_16259_n9386;
  wire AES_CORE_DATAPATH__abc_16259_n9388;
  wire AES_CORE_DATAPATH__abc_16259_n9389;
  wire AES_CORE_DATAPATH__abc_16259_n9391;
  wire AES_CORE_DATAPATH__abc_16259_n9392;
  wire AES_CORE_DATAPATH__abc_16259_n9393;
  wire AES_CORE_DATAPATH__abc_16259_n9394;
  wire AES_CORE_DATAPATH__abc_16259_n9395;
  wire AES_CORE_DATAPATH__abc_16259_n9396;
  wire AES_CORE_DATAPATH__abc_16259_n9397;
  wire AES_CORE_DATAPATH__abc_16259_n9399;
  wire AES_CORE_DATAPATH__abc_16259_n9400;
  wire AES_CORE_DATAPATH__abc_16259_n9401;
  wire AES_CORE_DATAPATH__abc_16259_n9402;
  wire AES_CORE_DATAPATH__abc_16259_n9403;
  wire AES_CORE_DATAPATH__abc_16259_n9404;
  wire AES_CORE_DATAPATH__abc_16259_n9405;
  wire AES_CORE_DATAPATH__abc_16259_n9407;
  wire AES_CORE_DATAPATH__abc_16259_n9408;
  wire AES_CORE_DATAPATH__abc_16259_n9409;
  wire AES_CORE_DATAPATH__abc_16259_n9410;
  wire AES_CORE_DATAPATH__abc_16259_n9411;
  wire AES_CORE_DATAPATH__abc_16259_n9412;
  wire AES_CORE_DATAPATH__abc_16259_n9413;
  wire AES_CORE_DATAPATH__abc_16259_n9415;
  wire AES_CORE_DATAPATH__abc_16259_n9416;
  wire AES_CORE_DATAPATH__abc_16259_n9417;
  wire AES_CORE_DATAPATH__abc_16259_n9418;
  wire AES_CORE_DATAPATH__abc_16259_n9419;
  wire AES_CORE_DATAPATH__abc_16259_n9420;
  wire AES_CORE_DATAPATH__abc_16259_n9421;
  wire AES_CORE_DATAPATH__abc_16259_n9423;
  wire AES_CORE_DATAPATH__abc_16259_n9424;
  wire AES_CORE_DATAPATH__abc_16259_n9425;
  wire AES_CORE_DATAPATH__abc_16259_n9426;
  wire AES_CORE_DATAPATH__abc_16259_n9427;
  wire AES_CORE_DATAPATH__abc_16259_n9428;
  wire AES_CORE_DATAPATH__abc_16259_n9429;
  wire AES_CORE_DATAPATH__abc_16259_n9431;
  wire AES_CORE_DATAPATH__abc_16259_n9432;
  wire AES_CORE_DATAPATH__abc_16259_n9433;
  wire AES_CORE_DATAPATH__abc_16259_n9434;
  wire AES_CORE_DATAPATH__abc_16259_n9435;
  wire AES_CORE_DATAPATH__abc_16259_n9436;
  wire AES_CORE_DATAPATH__abc_16259_n9437;
  wire AES_CORE_DATAPATH__abc_16259_n9439;
  wire AES_CORE_DATAPATH__abc_16259_n9440;
  wire AES_CORE_DATAPATH__abc_16259_n9441;
  wire AES_CORE_DATAPATH__abc_16259_n9442;
  wire AES_CORE_DATAPATH__abc_16259_n9443;
  wire AES_CORE_DATAPATH__abc_16259_n9444;
  wire AES_CORE_DATAPATH__abc_16259_n9445;
  wire AES_CORE_DATAPATH__abc_16259_n9447;
  wire AES_CORE_DATAPATH__abc_16259_n9448;
  wire AES_CORE_DATAPATH__abc_16259_n9449;
  wire AES_CORE_DATAPATH__abc_16259_n9450;
  wire AES_CORE_DATAPATH__abc_16259_n9451;
  wire AES_CORE_DATAPATH__abc_16259_n9452;
  wire AES_CORE_DATAPATH__abc_16259_n9453;
  wire AES_CORE_DATAPATH__abc_16259_n9455;
  wire AES_CORE_DATAPATH__abc_16259_n9456;
  wire AES_CORE_DATAPATH__abc_16259_n9457;
  wire AES_CORE_DATAPATH__abc_16259_n9458;
  wire AES_CORE_DATAPATH__abc_16259_n9459;
  wire AES_CORE_DATAPATH__abc_16259_n9460;
  wire AES_CORE_DATAPATH__abc_16259_n9461;
  wire AES_CORE_DATAPATH__abc_16259_n9463;
  wire AES_CORE_DATAPATH__abc_16259_n9464;
  wire AES_CORE_DATAPATH__abc_16259_n9465;
  wire AES_CORE_DATAPATH__abc_16259_n9466;
  wire AES_CORE_DATAPATH__abc_16259_n9467;
  wire AES_CORE_DATAPATH__abc_16259_n9468;
  wire AES_CORE_DATAPATH__abc_16259_n9469;
  wire AES_CORE_DATAPATH__abc_16259_n9471;
  wire AES_CORE_DATAPATH__abc_16259_n9472;
  wire AES_CORE_DATAPATH__abc_16259_n9473;
  wire AES_CORE_DATAPATH__abc_16259_n9474;
  wire AES_CORE_DATAPATH__abc_16259_n9475;
  wire AES_CORE_DATAPATH__abc_16259_n9476;
  wire AES_CORE_DATAPATH__abc_16259_n9477;
  wire AES_CORE_DATAPATH__abc_16259_n9478;
  wire AES_CORE_DATAPATH__abc_16259_n9480;
  wire AES_CORE_DATAPATH__abc_16259_n9481;
  wire AES_CORE_DATAPATH__abc_16259_n9482;
  wire AES_CORE_DATAPATH__abc_16259_n9483;
  wire AES_CORE_DATAPATH__abc_16259_n9484;
  wire AES_CORE_DATAPATH__abc_16259_n9485;
  wire AES_CORE_DATAPATH__abc_16259_n9486;
  wire AES_CORE_DATAPATH__abc_16259_n9487;
  wire AES_CORE_DATAPATH__abc_16259_n9489;
  wire AES_CORE_DATAPATH__abc_16259_n9490;
  wire AES_CORE_DATAPATH__abc_16259_n9491;
  wire AES_CORE_DATAPATH__abc_16259_n9492;
  wire AES_CORE_DATAPATH__abc_16259_n9493;
  wire AES_CORE_DATAPATH__abc_16259_n9494;
  wire AES_CORE_DATAPATH__abc_16259_n9495;
  wire AES_CORE_DATAPATH__abc_16259_n9497;
  wire AES_CORE_DATAPATH__abc_16259_n9498;
  wire AES_CORE_DATAPATH__abc_16259_n9499;
  wire AES_CORE_DATAPATH__abc_16259_n9500;
  wire AES_CORE_DATAPATH__abc_16259_n9501;
  wire AES_CORE_DATAPATH__abc_16259_n9502;
  wire AES_CORE_DATAPATH__abc_16259_n9503;
  wire AES_CORE_DATAPATH__abc_16259_n9504;
  wire AES_CORE_DATAPATH__abc_16259_n9506;
  wire AES_CORE_DATAPATH__abc_16259_n9507;
  wire AES_CORE_DATAPATH__abc_16259_n9508;
  wire AES_CORE_DATAPATH__abc_16259_n9509;
  wire AES_CORE_DATAPATH__abc_16259_n9510;
  wire AES_CORE_DATAPATH__abc_16259_n9511;
  wire AES_CORE_DATAPATH__abc_16259_n9512;
  wire AES_CORE_DATAPATH__abc_16259_n9514;
  wire AES_CORE_DATAPATH__abc_16259_n9515;
  wire AES_CORE_DATAPATH__abc_16259_n9516;
  wire AES_CORE_DATAPATH__abc_16259_n9517;
  wire AES_CORE_DATAPATH__abc_16259_n9518;
  wire AES_CORE_DATAPATH__abc_16259_n9519;
  wire AES_CORE_DATAPATH__abc_16259_n9520;
  wire AES_CORE_DATAPATH__abc_16259_n9521;
  wire AES_CORE_DATAPATH__abc_16259_n9523;
  wire AES_CORE_DATAPATH__abc_16259_n9524;
  wire AES_CORE_DATAPATH__abc_16259_n9525;
  wire AES_CORE_DATAPATH__abc_16259_n9526;
  wire AES_CORE_DATAPATH__abc_16259_n9527;
  wire AES_CORE_DATAPATH__abc_16259_n9528;
  wire AES_CORE_DATAPATH__abc_16259_n9529;
  wire AES_CORE_DATAPATH__abc_16259_n9531;
  wire AES_CORE_DATAPATH__abc_16259_n9532;
  wire AES_CORE_DATAPATH__abc_16259_n9533;
  wire AES_CORE_DATAPATH__abc_16259_n9534;
  wire AES_CORE_DATAPATH__abc_16259_n9535;
  wire AES_CORE_DATAPATH__abc_16259_n9536;
  wire AES_CORE_DATAPATH__abc_16259_n9537;
  wire AES_CORE_DATAPATH__abc_16259_n9538;
  wire AES_CORE_DATAPATH__abc_16259_n9540;
  wire AES_CORE_DATAPATH__abc_16259_n9541;
  wire AES_CORE_DATAPATH__abc_16259_n9542;
  wire AES_CORE_DATAPATH__abc_16259_n9543;
  wire AES_CORE_DATAPATH__abc_16259_n9544;
  wire AES_CORE_DATAPATH__abc_16259_n9545;
  wire AES_CORE_DATAPATH__abc_16259_n9546;
  wire AES_CORE_DATAPATH__abc_16259_n9548;
  wire AES_CORE_DATAPATH__abc_16259_n9549;
  wire AES_CORE_DATAPATH__abc_16259_n9550;
  wire AES_CORE_DATAPATH__abc_16259_n9551;
  wire AES_CORE_DATAPATH__abc_16259_n9552;
  wire AES_CORE_DATAPATH__abc_16259_n9553;
  wire AES_CORE_DATAPATH__abc_16259_n9554;
  wire AES_CORE_DATAPATH__abc_16259_n9556;
  wire AES_CORE_DATAPATH__abc_16259_n9557;
  wire AES_CORE_DATAPATH__abc_16259_n9558;
  wire AES_CORE_DATAPATH__abc_16259_n9559;
  wire AES_CORE_DATAPATH__abc_16259_n9560;
  wire AES_CORE_DATAPATH__abc_16259_n9561;
  wire AES_CORE_DATAPATH__abc_16259_n9562;
  wire AES_CORE_DATAPATH__abc_16259_n9564;
  wire AES_CORE_DATAPATH__abc_16259_n9565;
  wire AES_CORE_DATAPATH__abc_16259_n9566;
  wire AES_CORE_DATAPATH__abc_16259_n9567;
  wire AES_CORE_DATAPATH__abc_16259_n9568;
  wire AES_CORE_DATAPATH__abc_16259_n9569;
  wire AES_CORE_DATAPATH__abc_16259_n9570;
  wire AES_CORE_DATAPATH__abc_16259_n9571;
  wire AES_CORE_DATAPATH__abc_16259_n9573;
  wire AES_CORE_DATAPATH__abc_16259_n9574;
  wire AES_CORE_DATAPATH__abc_16259_n9575;
  wire AES_CORE_DATAPATH__abc_16259_n9576;
  wire AES_CORE_DATAPATH__abc_16259_n9577;
  wire AES_CORE_DATAPATH__abc_16259_n9578;
  wire AES_CORE_DATAPATH__abc_16259_n9579;
  wire AES_CORE_DATAPATH__abc_16259_n9581;
  wire AES_CORE_DATAPATH__abc_16259_n9582;
  wire AES_CORE_DATAPATH__abc_16259_n9583;
  wire AES_CORE_DATAPATH__abc_16259_n9584;
  wire AES_CORE_DATAPATH__abc_16259_n9585;
  wire AES_CORE_DATAPATH__abc_16259_n9586;
  wire AES_CORE_DATAPATH__abc_16259_n9587;
  wire AES_CORE_DATAPATH__abc_16259_n9589;
  wire AES_CORE_DATAPATH__abc_16259_n9590;
  wire AES_CORE_DATAPATH__abc_16259_n9591;
  wire AES_CORE_DATAPATH__abc_16259_n9592;
  wire AES_CORE_DATAPATH__abc_16259_n9593;
  wire AES_CORE_DATAPATH__abc_16259_n9594;
  wire AES_CORE_DATAPATH__abc_16259_n9595;
  wire AES_CORE_DATAPATH__abc_16259_n9597;
  wire AES_CORE_DATAPATH__abc_16259_n9598;
  wire AES_CORE_DATAPATH__abc_16259_n9599;
  wire AES_CORE_DATAPATH__abc_16259_n9600;
  wire AES_CORE_DATAPATH__abc_16259_n9601;
  wire AES_CORE_DATAPATH__abc_16259_n9602;
  wire AES_CORE_DATAPATH__abc_16259_n9603;
  wire AES_CORE_DATAPATH__abc_16259_n9605;
  wire AES_CORE_DATAPATH__abc_16259_n9606;
  wire AES_CORE_DATAPATH__abc_16259_n9607;
  wire AES_CORE_DATAPATH__abc_16259_n9608;
  wire AES_CORE_DATAPATH__abc_16259_n9609;
  wire AES_CORE_DATAPATH__abc_16259_n9610;
  wire AES_CORE_DATAPATH__abc_16259_n9611;
  wire AES_CORE_DATAPATH__abc_16259_n9613;
  wire AES_CORE_DATAPATH__abc_16259_n9614;
  wire AES_CORE_DATAPATH__abc_16259_n9615;
  wire AES_CORE_DATAPATH__abc_16259_n9616;
  wire AES_CORE_DATAPATH__abc_16259_n9617;
  wire AES_CORE_DATAPATH__abc_16259_n9618;
  wire AES_CORE_DATAPATH__abc_16259_n9619;
  wire AES_CORE_DATAPATH__abc_16259_n9621;
  wire AES_CORE_DATAPATH__abc_16259_n9622;
  wire AES_CORE_DATAPATH__abc_16259_n9623;
  wire AES_CORE_DATAPATH__abc_16259_n9624;
  wire AES_CORE_DATAPATH__abc_16259_n9625;
  wire AES_CORE_DATAPATH__abc_16259_n9626;
  wire AES_CORE_DATAPATH__abc_16259_n9627;
  wire AES_CORE_DATAPATH__abc_16259_n9629;
  wire AES_CORE_DATAPATH__abc_16259_n9630;
  wire AES_CORE_DATAPATH__abc_16259_n9631;
  wire AES_CORE_DATAPATH__abc_16259_n9632;
  wire AES_CORE_DATAPATH__abc_16259_n9633;
  wire AES_CORE_DATAPATH__abc_16259_n9634;
  wire AES_CORE_DATAPATH__abc_16259_n9635;
  wire AES_CORE_DATAPATH__abc_16259_n9637;
  wire AES_CORE_DATAPATH__abc_16259_n9638;
  wire AES_CORE_DATAPATH__abc_16259_n9639;
  wire AES_CORE_DATAPATH__abc_16259_n9640;
  wire AES_CORE_DATAPATH__abc_16259_n9641;
  wire AES_CORE_DATAPATH__abc_16259_n9642;
  wire AES_CORE_DATAPATH__abc_16259_n9643;
  wire AES_CORE_DATAPATH__abc_16259_n9645;
  wire AES_CORE_DATAPATH__abc_16259_n9646;
  wire AES_CORE_DATAPATH__abc_16259_n9647;
  wire AES_CORE_DATAPATH__abc_16259_n9648;
  wire AES_CORE_DATAPATH__abc_16259_n9649;
  wire AES_CORE_DATAPATH__abc_16259_n9650;
  wire AES_CORE_DATAPATH__abc_16259_n9651;
  wire AES_CORE_DATAPATH__abc_16259_n9653;
  wire AES_CORE_DATAPATH__abc_16259_n9654;
  wire AES_CORE_DATAPATH__abc_16259_n9654_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n9654_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n9654_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n9654_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n9654_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n9655;
  wire AES_CORE_DATAPATH__abc_16259_n9657;
  wire AES_CORE_DATAPATH__abc_16259_n9658;
  wire AES_CORE_DATAPATH__abc_16259_n9660;
  wire AES_CORE_DATAPATH__abc_16259_n9661;
  wire AES_CORE_DATAPATH__abc_16259_n9663;
  wire AES_CORE_DATAPATH__abc_16259_n9664;
  wire AES_CORE_DATAPATH__abc_16259_n9666;
  wire AES_CORE_DATAPATH__abc_16259_n9667;
  wire AES_CORE_DATAPATH__abc_16259_n9669;
  wire AES_CORE_DATAPATH__abc_16259_n9670;
  wire AES_CORE_DATAPATH__abc_16259_n9672;
  wire AES_CORE_DATAPATH__abc_16259_n9673;
  wire AES_CORE_DATAPATH__abc_16259_n9675;
  wire AES_CORE_DATAPATH__abc_16259_n9676;
  wire AES_CORE_DATAPATH__abc_16259_n9678;
  wire AES_CORE_DATAPATH__abc_16259_n9679;
  wire AES_CORE_DATAPATH__abc_16259_n9681;
  wire AES_CORE_DATAPATH__abc_16259_n9682;
  wire AES_CORE_DATAPATH__abc_16259_n9684;
  wire AES_CORE_DATAPATH__abc_16259_n9685;
  wire AES_CORE_DATAPATH__abc_16259_n9687;
  wire AES_CORE_DATAPATH__abc_16259_n9688;
  wire AES_CORE_DATAPATH__abc_16259_n9690;
  wire AES_CORE_DATAPATH__abc_16259_n9691;
  wire AES_CORE_DATAPATH__abc_16259_n9693;
  wire AES_CORE_DATAPATH__abc_16259_n9694;
  wire AES_CORE_DATAPATH__abc_16259_n9696;
  wire AES_CORE_DATAPATH__abc_16259_n9697;
  wire AES_CORE_DATAPATH__abc_16259_n9699;
  wire AES_CORE_DATAPATH__abc_16259_n9700;
  wire AES_CORE_DATAPATH__abc_16259_n9702;
  wire AES_CORE_DATAPATH__abc_16259_n9703;
  wire AES_CORE_DATAPATH__abc_16259_n9705;
  wire AES_CORE_DATAPATH__abc_16259_n9706;
  wire AES_CORE_DATAPATH__abc_16259_n9708;
  wire AES_CORE_DATAPATH__abc_16259_n9709;
  wire AES_CORE_DATAPATH__abc_16259_n9711;
  wire AES_CORE_DATAPATH__abc_16259_n9712;
  wire AES_CORE_DATAPATH__abc_16259_n9714;
  wire AES_CORE_DATAPATH__abc_16259_n9715;
  wire AES_CORE_DATAPATH__abc_16259_n9717;
  wire AES_CORE_DATAPATH__abc_16259_n9718;
  wire AES_CORE_DATAPATH__abc_16259_n9720;
  wire AES_CORE_DATAPATH__abc_16259_n9721;
  wire AES_CORE_DATAPATH__abc_16259_n9723;
  wire AES_CORE_DATAPATH__abc_16259_n9724;
  wire AES_CORE_DATAPATH__abc_16259_n9726;
  wire AES_CORE_DATAPATH__abc_16259_n9727;
  wire AES_CORE_DATAPATH__abc_16259_n9729;
  wire AES_CORE_DATAPATH__abc_16259_n9730;
  wire AES_CORE_DATAPATH__abc_16259_n9732;
  wire AES_CORE_DATAPATH__abc_16259_n9733;
  wire AES_CORE_DATAPATH__abc_16259_n9735;
  wire AES_CORE_DATAPATH__abc_16259_n9736;
  wire AES_CORE_DATAPATH__abc_16259_n9738;
  wire AES_CORE_DATAPATH__abc_16259_n9739;
  wire AES_CORE_DATAPATH__abc_16259_n9741;
  wire AES_CORE_DATAPATH__abc_16259_n9742;
  wire AES_CORE_DATAPATH__abc_16259_n9744;
  wire AES_CORE_DATAPATH__abc_16259_n9745;
  wire AES_CORE_DATAPATH__abc_16259_n9747;
  wire AES_CORE_DATAPATH__abc_16259_n9748;
  wire AES_CORE_DATAPATH__abc_16259_n9750;
  wire AES_CORE_DATAPATH__abc_16259_n9751;
  wire AES_CORE_DATAPATH__abc_16259_n9752;
  wire AES_CORE_DATAPATH__abc_16259_n9752_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n9752_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n9752_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n9752_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n9752_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n9752_bF_buf5;
  wire AES_CORE_DATAPATH__abc_16259_n9752_bF_buf6;
  wire AES_CORE_DATAPATH__abc_16259_n9752_bF_buf7;
  wire AES_CORE_DATAPATH__abc_16259_n9753;
  wire AES_CORE_DATAPATH__abc_16259_n9753_bF_buf0;
  wire AES_CORE_DATAPATH__abc_16259_n9753_bF_buf1;
  wire AES_CORE_DATAPATH__abc_16259_n9753_bF_buf2;
  wire AES_CORE_DATAPATH__abc_16259_n9753_bF_buf3;
  wire AES_CORE_DATAPATH__abc_16259_n9753_bF_buf4;
  wire AES_CORE_DATAPATH__abc_16259_n9753_bF_buf5;
  wire AES_CORE_DATAPATH__abc_16259_n9753_bF_buf6;
  wire AES_CORE_DATAPATH__abc_16259_n9754;
  wire AES_CORE_DATAPATH__abc_16259_n9755;
  wire AES_CORE_DATAPATH__abc_16259_n9757;
  wire AES_CORE_DATAPATH__abc_16259_n9758;
  wire AES_CORE_DATAPATH__abc_16259_n9760;
  wire AES_CORE_DATAPATH__abc_16259_n9761;
  wire AES_CORE_DATAPATH__abc_16259_n9763;
  wire AES_CORE_DATAPATH__abc_16259_n9764;
  wire AES_CORE_DATAPATH__abc_16259_n9766;
  wire AES_CORE_DATAPATH__abc_16259_n9767;
  wire AES_CORE_DATAPATH__abc_16259_n9769;
  wire AES_CORE_DATAPATH__abc_16259_n9770;
  wire AES_CORE_DATAPATH__abc_16259_n9772;
  wire AES_CORE_DATAPATH__abc_16259_n9773;
  wire AES_CORE_DATAPATH__abc_16259_n9775;
  wire AES_CORE_DATAPATH__abc_16259_n9776;
  wire AES_CORE_DATAPATH__abc_16259_n9778;
  wire AES_CORE_DATAPATH__abc_16259_n9779;
  wire AES_CORE_DATAPATH__abc_16259_n9781;
  wire AES_CORE_DATAPATH__abc_16259_n9782;
  wire AES_CORE_DATAPATH__abc_16259_n9784;
  wire AES_CORE_DATAPATH__abc_16259_n9785;
  wire AES_CORE_DATAPATH__abc_16259_n9786;
  wire AES_CORE_DATAPATH__abc_16259_n9788;
  wire AES_CORE_DATAPATH__abc_16259_n9789;
  wire AES_CORE_DATAPATH__abc_16259_n9790;
  wire AES_CORE_DATAPATH__abc_16259_n9792;
  wire AES_CORE_DATAPATH__abc_16259_n9793;
  wire AES_CORE_DATAPATH__abc_16259_n9795;
  wire AES_CORE_DATAPATH__abc_16259_n9796;
  wire AES_CORE_DATAPATH__abc_16259_n9797;
  wire AES_CORE_DATAPATH__abc_16259_n9799;
  wire AES_CORE_DATAPATH__abc_16259_n9800;
  wire AES_CORE_DATAPATH__abc_16259_n9802;
  wire AES_CORE_DATAPATH__abc_16259_n9803;
  wire AES_CORE_DATAPATH__abc_16259_n9804;
  wire AES_CORE_DATAPATH__abc_16259_n9806;
  wire AES_CORE_DATAPATH__abc_16259_n9807;
  wire AES_CORE_DATAPATH__abc_16259_n9809;
  wire AES_CORE_DATAPATH__abc_16259_n9810;
  wire AES_CORE_DATAPATH__abc_16259_n9811;
  wire AES_CORE_DATAPATH__abc_16259_n9813;
  wire AES_CORE_DATAPATH__abc_16259_n9814;
  wire AES_CORE_DATAPATH__abc_16259_n9816;
  wire AES_CORE_DATAPATH__abc_16259_n9817;
  wire AES_CORE_DATAPATH__abc_16259_n9819;
  wire AES_CORE_DATAPATH__abc_16259_n9820;
  wire AES_CORE_DATAPATH__abc_16259_n9822;
  wire AES_CORE_DATAPATH__abc_16259_n9823;
  wire AES_CORE_DATAPATH__abc_16259_n9824;
  wire AES_CORE_DATAPATH__abc_16259_n9826;
  wire AES_CORE_DATAPATH__abc_16259_n9827;
  wire AES_CORE_DATAPATH__abc_16259_n9829;
  wire AES_CORE_DATAPATH__abc_16259_n9830;
  wire AES_CORE_DATAPATH__abc_16259_n9832;
  wire AES_CORE_DATAPATH__abc_16259_n9833;
  wire AES_CORE_DATAPATH__abc_16259_n9835;
  wire AES_CORE_DATAPATH__abc_16259_n9836;
  wire AES_CORE_DATAPATH__abc_16259_n9838;
  wire AES_CORE_DATAPATH__abc_16259_n9839;
  wire AES_CORE_DATAPATH__abc_16259_n9841;
  wire AES_CORE_DATAPATH__abc_16259_n9842;
  wire AES_CORE_DATAPATH__abc_16259_n9844;
  wire AES_CORE_DATAPATH__abc_16259_n9845;
  wire AES_CORE_DATAPATH__abc_16259_n9847;
  wire AES_CORE_DATAPATH__abc_16259_n9848;
  wire AES_CORE_DATAPATH__abc_16259_n9850;
  wire AES_CORE_DATAPATH__abc_16259_n9851;
  wire AES_CORE_DATAPATH__abc_16259_n9853;
  wire AES_CORE_DATAPATH__abc_16259_n9854;
  wire AES_CORE_DATAPATH__abc_16259_n9856;
  wire AES_CORE_DATAPATH__abc_16259_n9857;
  wire AES_CORE_DATAPATH__abc_16259_n9858;
  wire AES_CORE_DATAPATH__abc_16259_n9859;
  wire AES_CORE_DATAPATH__abc_16259_n9860;
  wire AES_CORE_DATAPATH__abc_16259_n9861;
  wire AES_CORE_DATAPATH__abc_16259_n9862;
  wire AES_CORE_DATAPATH__abc_16259_n9864;
  wire AES_CORE_DATAPATH__abc_16259_n9865;
  wire AES_CORE_DATAPATH__abc_16259_n9866;
  wire AES_CORE_DATAPATH__abc_16259_n9867;
  wire AES_CORE_DATAPATH__abc_16259_n9868;
  wire AES_CORE_DATAPATH__abc_16259_n9869;
  wire AES_CORE_DATAPATH__abc_16259_n9870;
  wire AES_CORE_DATAPATH__abc_16259_n9872;
  wire AES_CORE_DATAPATH__abc_16259_n9873;
  wire AES_CORE_DATAPATH__abc_16259_n9874;
  wire AES_CORE_DATAPATH__abc_16259_n9875;
  wire AES_CORE_DATAPATH__abc_16259_n9876;
  wire AES_CORE_DATAPATH__abc_16259_n9877;
  wire AES_CORE_DATAPATH__abc_16259_n9878;
  wire AES_CORE_DATAPATH__abc_16259_n9880;
  wire AES_CORE_DATAPATH__abc_16259_n9881;
  wire AES_CORE_DATAPATH__abc_16259_n9882;
  wire AES_CORE_DATAPATH__abc_16259_n9883;
  wire AES_CORE_DATAPATH__abc_16259_n9884;
  wire AES_CORE_DATAPATH__abc_16259_n9885;
  wire AES_CORE_DATAPATH__abc_16259_n9886;
  wire AES_CORE_DATAPATH__abc_16259_n9888;
  wire AES_CORE_DATAPATH__abc_16259_n9889;
  wire AES_CORE_DATAPATH__abc_16259_n9890;
  wire AES_CORE_DATAPATH__abc_16259_n9891;
  wire AES_CORE_DATAPATH__abc_16259_n9892;
  wire AES_CORE_DATAPATH__abc_16259_n9893;
  wire AES_CORE_DATAPATH__abc_16259_n9894;
  wire AES_CORE_DATAPATH__abc_16259_n9896;
  wire AES_CORE_DATAPATH__abc_16259_n9897;
  wire AES_CORE_DATAPATH__abc_16259_n9898;
  wire AES_CORE_DATAPATH__abc_16259_n9899;
  wire AES_CORE_DATAPATH__abc_16259_n9900;
  wire AES_CORE_DATAPATH__abc_16259_n9901;
  wire AES_CORE_DATAPATH__abc_16259_n9902;
  wire AES_CORE_DATAPATH__abc_16259_n9904;
  wire AES_CORE_DATAPATH__abc_16259_n9905;
  wire AES_CORE_DATAPATH__abc_16259_n9906;
  wire AES_CORE_DATAPATH__abc_16259_n9907;
  wire AES_CORE_DATAPATH__abc_16259_n9908;
  wire AES_CORE_DATAPATH__abc_16259_n9909;
  wire AES_CORE_DATAPATH__abc_16259_n9910;
  wire AES_CORE_DATAPATH__abc_16259_n9912;
  wire AES_CORE_DATAPATH__abc_16259_n9913;
  wire AES_CORE_DATAPATH__abc_16259_n9914;
  wire AES_CORE_DATAPATH__abc_16259_n9915;
  wire AES_CORE_DATAPATH__abc_16259_n9916;
  wire AES_CORE_DATAPATH__abc_16259_n9917;
  wire AES_CORE_DATAPATH__abc_16259_n9918;
  wire AES_CORE_DATAPATH__abc_16259_n9920;
  wire AES_CORE_DATAPATH__abc_16259_n9921;
  wire AES_CORE_DATAPATH__abc_16259_n9922;
  wire AES_CORE_DATAPATH__abc_16259_n9923;
  wire AES_CORE_DATAPATH__abc_16259_n9924;
  wire AES_CORE_DATAPATH__abc_16259_n9925;
  wire AES_CORE_DATAPATH__abc_16259_n9926;
  wire AES_CORE_DATAPATH__abc_16259_n9928;
  wire AES_CORE_DATAPATH__abc_16259_n9929;
  wire AES_CORE_DATAPATH__abc_16259_n9930;
  wire AES_CORE_DATAPATH__abc_16259_n9931;
  wire AES_CORE_DATAPATH__abc_16259_n9932;
  wire AES_CORE_DATAPATH__abc_16259_n9933;
  wire AES_CORE_DATAPATH__abc_16259_n9934;
  wire AES_CORE_DATAPATH__abc_16259_n9936;
  wire AES_CORE_DATAPATH__abc_16259_n9937;
  wire AES_CORE_DATAPATH__abc_16259_n9938;
  wire AES_CORE_DATAPATH__abc_16259_n9939;
  wire AES_CORE_DATAPATH__abc_16259_n9940;
  wire AES_CORE_DATAPATH__abc_16259_n9941;
  wire AES_CORE_DATAPATH__abc_16259_n9942;
  wire AES_CORE_DATAPATH__abc_16259_n9943;
  wire AES_CORE_DATAPATH__abc_16259_n9945;
  wire AES_CORE_DATAPATH__abc_16259_n9946;
  wire AES_CORE_DATAPATH__abc_16259_n9947;
  wire AES_CORE_DATAPATH__abc_16259_n9948;
  wire AES_CORE_DATAPATH__abc_16259_n9949;
  wire AES_CORE_DATAPATH__abc_16259_n9950;
  wire AES_CORE_DATAPATH__abc_16259_n9951;
  wire AES_CORE_DATAPATH__abc_16259_n9952;
  wire AES_CORE_DATAPATH__abc_16259_n9954;
  wire AES_CORE_DATAPATH__abc_16259_n9955;
  wire AES_CORE_DATAPATH__abc_16259_n9956;
  wire AES_CORE_DATAPATH__abc_16259_n9957;
  wire AES_CORE_DATAPATH__abc_16259_n9958;
  wire AES_CORE_DATAPATH__abc_16259_n9959;
  wire AES_CORE_DATAPATH__abc_16259_n9960;
  wire AES_CORE_DATAPATH__abc_16259_n9962;
  wire AES_CORE_DATAPATH__abc_16259_n9963;
  wire AES_CORE_DATAPATH__abc_16259_n9964;
  wire AES_CORE_DATAPATH__abc_16259_n9965;
  wire AES_CORE_DATAPATH__abc_16259_n9966;
  wire AES_CORE_DATAPATH__abc_16259_n9967;
  wire AES_CORE_DATAPATH__abc_16259_n9968;
  wire AES_CORE_DATAPATH__abc_16259_n9969;
  wire AES_CORE_DATAPATH__abc_16259_n9971;
  wire AES_CORE_DATAPATH__abc_16259_n9972;
  wire AES_CORE_DATAPATH__abc_16259_n9973;
  wire AES_CORE_DATAPATH__abc_16259_n9974;
  wire AES_CORE_DATAPATH__abc_16259_n9975;
  wire AES_CORE_DATAPATH__abc_16259_n9976;
  wire AES_CORE_DATAPATH__abc_16259_n9977;
  wire AES_CORE_DATAPATH__abc_16259_n9979;
  wire AES_CORE_DATAPATH__abc_16259_n9980;
  wire AES_CORE_DATAPATH__abc_16259_n9981;
  wire AES_CORE_DATAPATH__abc_16259_n9982;
  wire AES_CORE_DATAPATH__abc_16259_n9983;
  wire AES_CORE_DATAPATH__abc_16259_n9984;
  wire AES_CORE_DATAPATH__abc_16259_n9985;
  wire AES_CORE_DATAPATH__abc_16259_n9986;
  wire AES_CORE_DATAPATH__abc_16259_n9988;
  wire AES_CORE_DATAPATH__abc_16259_n9989;
  wire AES_CORE_DATAPATH__abc_16259_n9990;
  wire AES_CORE_DATAPATH__abc_16259_n9991;
  wire AES_CORE_DATAPATH__abc_16259_n9992;
  wire AES_CORE_DATAPATH__abc_16259_n9993;
  wire AES_CORE_DATAPATH__abc_16259_n9994;
  wire AES_CORE_DATAPATH__abc_16259_n9996;
  wire AES_CORE_DATAPATH__abc_16259_n9997;
  wire AES_CORE_DATAPATH__abc_16259_n9998;
  wire AES_CORE_DATAPATH__abc_16259_n9999;
  wire AES_CORE_DATAPATH_bkp_0__0_;
  wire AES_CORE_DATAPATH_bkp_0__10_;
  wire AES_CORE_DATAPATH_bkp_0__11_;
  wire AES_CORE_DATAPATH_bkp_0__12_;
  wire AES_CORE_DATAPATH_bkp_0__13_;
  wire AES_CORE_DATAPATH_bkp_0__14_;
  wire AES_CORE_DATAPATH_bkp_0__15_;
  wire AES_CORE_DATAPATH_bkp_0__16_;
  wire AES_CORE_DATAPATH_bkp_0__17_;
  wire AES_CORE_DATAPATH_bkp_0__18_;
  wire AES_CORE_DATAPATH_bkp_0__19_;
  wire AES_CORE_DATAPATH_bkp_0__1_;
  wire AES_CORE_DATAPATH_bkp_0__20_;
  wire AES_CORE_DATAPATH_bkp_0__21_;
  wire AES_CORE_DATAPATH_bkp_0__22_;
  wire AES_CORE_DATAPATH_bkp_0__23_;
  wire AES_CORE_DATAPATH_bkp_0__24_;
  wire AES_CORE_DATAPATH_bkp_0__25_;
  wire AES_CORE_DATAPATH_bkp_0__26_;
  wire AES_CORE_DATAPATH_bkp_0__27_;
  wire AES_CORE_DATAPATH_bkp_0__28_;
  wire AES_CORE_DATAPATH_bkp_0__29_;
  wire AES_CORE_DATAPATH_bkp_0__2_;
  wire AES_CORE_DATAPATH_bkp_0__30_;
  wire AES_CORE_DATAPATH_bkp_0__31_;
  wire AES_CORE_DATAPATH_bkp_0__3_;
  wire AES_CORE_DATAPATH_bkp_0__4_;
  wire AES_CORE_DATAPATH_bkp_0__5_;
  wire AES_CORE_DATAPATH_bkp_0__6_;
  wire AES_CORE_DATAPATH_bkp_0__7_;
  wire AES_CORE_DATAPATH_bkp_0__8_;
  wire AES_CORE_DATAPATH_bkp_0__9_;
  wire AES_CORE_DATAPATH_bkp_1_0__0_;
  wire AES_CORE_DATAPATH_bkp_1_0__10_;
  wire AES_CORE_DATAPATH_bkp_1_0__11_;
  wire AES_CORE_DATAPATH_bkp_1_0__12_;
  wire AES_CORE_DATAPATH_bkp_1_0__13_;
  wire AES_CORE_DATAPATH_bkp_1_0__14_;
  wire AES_CORE_DATAPATH_bkp_1_0__15_;
  wire AES_CORE_DATAPATH_bkp_1_0__16_;
  wire AES_CORE_DATAPATH_bkp_1_0__17_;
  wire AES_CORE_DATAPATH_bkp_1_0__18_;
  wire AES_CORE_DATAPATH_bkp_1_0__19_;
  wire AES_CORE_DATAPATH_bkp_1_0__1_;
  wire AES_CORE_DATAPATH_bkp_1_0__20_;
  wire AES_CORE_DATAPATH_bkp_1_0__21_;
  wire AES_CORE_DATAPATH_bkp_1_0__22_;
  wire AES_CORE_DATAPATH_bkp_1_0__23_;
  wire AES_CORE_DATAPATH_bkp_1_0__24_;
  wire AES_CORE_DATAPATH_bkp_1_0__25_;
  wire AES_CORE_DATAPATH_bkp_1_0__26_;
  wire AES_CORE_DATAPATH_bkp_1_0__27_;
  wire AES_CORE_DATAPATH_bkp_1_0__28_;
  wire AES_CORE_DATAPATH_bkp_1_0__29_;
  wire AES_CORE_DATAPATH_bkp_1_0__2_;
  wire AES_CORE_DATAPATH_bkp_1_0__30_;
  wire AES_CORE_DATAPATH_bkp_1_0__31_;
  wire AES_CORE_DATAPATH_bkp_1_0__3_;
  wire AES_CORE_DATAPATH_bkp_1_0__4_;
  wire AES_CORE_DATAPATH_bkp_1_0__5_;
  wire AES_CORE_DATAPATH_bkp_1_0__6_;
  wire AES_CORE_DATAPATH_bkp_1_0__7_;
  wire AES_CORE_DATAPATH_bkp_1_0__8_;
  wire AES_CORE_DATAPATH_bkp_1_0__9_;
  wire AES_CORE_DATAPATH_bkp_1_1__0_;
  wire AES_CORE_DATAPATH_bkp_1_1__10_;
  wire AES_CORE_DATAPATH_bkp_1_1__11_;
  wire AES_CORE_DATAPATH_bkp_1_1__12_;
  wire AES_CORE_DATAPATH_bkp_1_1__13_;
  wire AES_CORE_DATAPATH_bkp_1_1__14_;
  wire AES_CORE_DATAPATH_bkp_1_1__15_;
  wire AES_CORE_DATAPATH_bkp_1_1__16_;
  wire AES_CORE_DATAPATH_bkp_1_1__17_;
  wire AES_CORE_DATAPATH_bkp_1_1__18_;
  wire AES_CORE_DATAPATH_bkp_1_1__19_;
  wire AES_CORE_DATAPATH_bkp_1_1__1_;
  wire AES_CORE_DATAPATH_bkp_1_1__20_;
  wire AES_CORE_DATAPATH_bkp_1_1__21_;
  wire AES_CORE_DATAPATH_bkp_1_1__22_;
  wire AES_CORE_DATAPATH_bkp_1_1__23_;
  wire AES_CORE_DATAPATH_bkp_1_1__24_;
  wire AES_CORE_DATAPATH_bkp_1_1__25_;
  wire AES_CORE_DATAPATH_bkp_1_1__26_;
  wire AES_CORE_DATAPATH_bkp_1_1__27_;
  wire AES_CORE_DATAPATH_bkp_1_1__28_;
  wire AES_CORE_DATAPATH_bkp_1_1__29_;
  wire AES_CORE_DATAPATH_bkp_1_1__2_;
  wire AES_CORE_DATAPATH_bkp_1_1__30_;
  wire AES_CORE_DATAPATH_bkp_1_1__31_;
  wire AES_CORE_DATAPATH_bkp_1_1__3_;
  wire AES_CORE_DATAPATH_bkp_1_1__4_;
  wire AES_CORE_DATAPATH_bkp_1_1__5_;
  wire AES_CORE_DATAPATH_bkp_1_1__6_;
  wire AES_CORE_DATAPATH_bkp_1_1__7_;
  wire AES_CORE_DATAPATH_bkp_1_1__8_;
  wire AES_CORE_DATAPATH_bkp_1_1__9_;
  wire AES_CORE_DATAPATH_bkp_1_2__0_;
  wire AES_CORE_DATAPATH_bkp_1_2__10_;
  wire AES_CORE_DATAPATH_bkp_1_2__11_;
  wire AES_CORE_DATAPATH_bkp_1_2__12_;
  wire AES_CORE_DATAPATH_bkp_1_2__13_;
  wire AES_CORE_DATAPATH_bkp_1_2__14_;
  wire AES_CORE_DATAPATH_bkp_1_2__15_;
  wire AES_CORE_DATAPATH_bkp_1_2__16_;
  wire AES_CORE_DATAPATH_bkp_1_2__17_;
  wire AES_CORE_DATAPATH_bkp_1_2__18_;
  wire AES_CORE_DATAPATH_bkp_1_2__19_;
  wire AES_CORE_DATAPATH_bkp_1_2__1_;
  wire AES_CORE_DATAPATH_bkp_1_2__20_;
  wire AES_CORE_DATAPATH_bkp_1_2__21_;
  wire AES_CORE_DATAPATH_bkp_1_2__22_;
  wire AES_CORE_DATAPATH_bkp_1_2__23_;
  wire AES_CORE_DATAPATH_bkp_1_2__24_;
  wire AES_CORE_DATAPATH_bkp_1_2__25_;
  wire AES_CORE_DATAPATH_bkp_1_2__26_;
  wire AES_CORE_DATAPATH_bkp_1_2__27_;
  wire AES_CORE_DATAPATH_bkp_1_2__28_;
  wire AES_CORE_DATAPATH_bkp_1_2__29_;
  wire AES_CORE_DATAPATH_bkp_1_2__2_;
  wire AES_CORE_DATAPATH_bkp_1_2__30_;
  wire AES_CORE_DATAPATH_bkp_1_2__31_;
  wire AES_CORE_DATAPATH_bkp_1_2__3_;
  wire AES_CORE_DATAPATH_bkp_1_2__4_;
  wire AES_CORE_DATAPATH_bkp_1_2__5_;
  wire AES_CORE_DATAPATH_bkp_1_2__6_;
  wire AES_CORE_DATAPATH_bkp_1_2__7_;
  wire AES_CORE_DATAPATH_bkp_1_2__8_;
  wire AES_CORE_DATAPATH_bkp_1_2__9_;
  wire AES_CORE_DATAPATH_bkp_1_3__0_;
  wire AES_CORE_DATAPATH_bkp_1_3__10_;
  wire AES_CORE_DATAPATH_bkp_1_3__11_;
  wire AES_CORE_DATAPATH_bkp_1_3__12_;
  wire AES_CORE_DATAPATH_bkp_1_3__13_;
  wire AES_CORE_DATAPATH_bkp_1_3__14_;
  wire AES_CORE_DATAPATH_bkp_1_3__15_;
  wire AES_CORE_DATAPATH_bkp_1_3__16_;
  wire AES_CORE_DATAPATH_bkp_1_3__17_;
  wire AES_CORE_DATAPATH_bkp_1_3__18_;
  wire AES_CORE_DATAPATH_bkp_1_3__19_;
  wire AES_CORE_DATAPATH_bkp_1_3__1_;
  wire AES_CORE_DATAPATH_bkp_1_3__20_;
  wire AES_CORE_DATAPATH_bkp_1_3__21_;
  wire AES_CORE_DATAPATH_bkp_1_3__22_;
  wire AES_CORE_DATAPATH_bkp_1_3__23_;
  wire AES_CORE_DATAPATH_bkp_1_3__24_;
  wire AES_CORE_DATAPATH_bkp_1_3__25_;
  wire AES_CORE_DATAPATH_bkp_1_3__26_;
  wire AES_CORE_DATAPATH_bkp_1_3__27_;
  wire AES_CORE_DATAPATH_bkp_1_3__28_;
  wire AES_CORE_DATAPATH_bkp_1_3__29_;
  wire AES_CORE_DATAPATH_bkp_1_3__2_;
  wire AES_CORE_DATAPATH_bkp_1_3__30_;
  wire AES_CORE_DATAPATH_bkp_1_3__31_;
  wire AES_CORE_DATAPATH_bkp_1_3__3_;
  wire AES_CORE_DATAPATH_bkp_1_3__4_;
  wire AES_CORE_DATAPATH_bkp_1_3__5_;
  wire AES_CORE_DATAPATH_bkp_1_3__6_;
  wire AES_CORE_DATAPATH_bkp_1_3__7_;
  wire AES_CORE_DATAPATH_bkp_1_3__8_;
  wire AES_CORE_DATAPATH_bkp_1_3__9_;
  wire AES_CORE_DATAPATH_bkp_1__0_;
  wire AES_CORE_DATAPATH_bkp_1__10_;
  wire AES_CORE_DATAPATH_bkp_1__11_;
  wire AES_CORE_DATAPATH_bkp_1__12_;
  wire AES_CORE_DATAPATH_bkp_1__13_;
  wire AES_CORE_DATAPATH_bkp_1__14_;
  wire AES_CORE_DATAPATH_bkp_1__15_;
  wire AES_CORE_DATAPATH_bkp_1__16_;
  wire AES_CORE_DATAPATH_bkp_1__17_;
  wire AES_CORE_DATAPATH_bkp_1__18_;
  wire AES_CORE_DATAPATH_bkp_1__19_;
  wire AES_CORE_DATAPATH_bkp_1__1_;
  wire AES_CORE_DATAPATH_bkp_1__20_;
  wire AES_CORE_DATAPATH_bkp_1__21_;
  wire AES_CORE_DATAPATH_bkp_1__22_;
  wire AES_CORE_DATAPATH_bkp_1__23_;
  wire AES_CORE_DATAPATH_bkp_1__24_;
  wire AES_CORE_DATAPATH_bkp_1__25_;
  wire AES_CORE_DATAPATH_bkp_1__26_;
  wire AES_CORE_DATAPATH_bkp_1__27_;
  wire AES_CORE_DATAPATH_bkp_1__28_;
  wire AES_CORE_DATAPATH_bkp_1__29_;
  wire AES_CORE_DATAPATH_bkp_1__2_;
  wire AES_CORE_DATAPATH_bkp_1__30_;
  wire AES_CORE_DATAPATH_bkp_1__31_;
  wire AES_CORE_DATAPATH_bkp_1__3_;
  wire AES_CORE_DATAPATH_bkp_1__4_;
  wire AES_CORE_DATAPATH_bkp_1__5_;
  wire AES_CORE_DATAPATH_bkp_1__6_;
  wire AES_CORE_DATAPATH_bkp_1__7_;
  wire AES_CORE_DATAPATH_bkp_1__8_;
  wire AES_CORE_DATAPATH_bkp_1__9_;
  wire AES_CORE_DATAPATH_bkp_2__0_;
  wire AES_CORE_DATAPATH_bkp_2__10_;
  wire AES_CORE_DATAPATH_bkp_2__11_;
  wire AES_CORE_DATAPATH_bkp_2__12_;
  wire AES_CORE_DATAPATH_bkp_2__13_;
  wire AES_CORE_DATAPATH_bkp_2__14_;
  wire AES_CORE_DATAPATH_bkp_2__15_;
  wire AES_CORE_DATAPATH_bkp_2__16_;
  wire AES_CORE_DATAPATH_bkp_2__17_;
  wire AES_CORE_DATAPATH_bkp_2__18_;
  wire AES_CORE_DATAPATH_bkp_2__19_;
  wire AES_CORE_DATAPATH_bkp_2__1_;
  wire AES_CORE_DATAPATH_bkp_2__20_;
  wire AES_CORE_DATAPATH_bkp_2__21_;
  wire AES_CORE_DATAPATH_bkp_2__22_;
  wire AES_CORE_DATAPATH_bkp_2__23_;
  wire AES_CORE_DATAPATH_bkp_2__24_;
  wire AES_CORE_DATAPATH_bkp_2__25_;
  wire AES_CORE_DATAPATH_bkp_2__26_;
  wire AES_CORE_DATAPATH_bkp_2__27_;
  wire AES_CORE_DATAPATH_bkp_2__28_;
  wire AES_CORE_DATAPATH_bkp_2__29_;
  wire AES_CORE_DATAPATH_bkp_2__2_;
  wire AES_CORE_DATAPATH_bkp_2__30_;
  wire AES_CORE_DATAPATH_bkp_2__31_;
  wire AES_CORE_DATAPATH_bkp_2__3_;
  wire AES_CORE_DATAPATH_bkp_2__4_;
  wire AES_CORE_DATAPATH_bkp_2__5_;
  wire AES_CORE_DATAPATH_bkp_2__6_;
  wire AES_CORE_DATAPATH_bkp_2__7_;
  wire AES_CORE_DATAPATH_bkp_2__8_;
  wire AES_CORE_DATAPATH_bkp_2__9_;
  wire AES_CORE_DATAPATH_bkp_3__0_;
  wire AES_CORE_DATAPATH_bkp_3__10_;
  wire AES_CORE_DATAPATH_bkp_3__11_;
  wire AES_CORE_DATAPATH_bkp_3__12_;
  wire AES_CORE_DATAPATH_bkp_3__13_;
  wire AES_CORE_DATAPATH_bkp_3__14_;
  wire AES_CORE_DATAPATH_bkp_3__15_;
  wire AES_CORE_DATAPATH_bkp_3__16_;
  wire AES_CORE_DATAPATH_bkp_3__17_;
  wire AES_CORE_DATAPATH_bkp_3__18_;
  wire AES_CORE_DATAPATH_bkp_3__19_;
  wire AES_CORE_DATAPATH_bkp_3__1_;
  wire AES_CORE_DATAPATH_bkp_3__20_;
  wire AES_CORE_DATAPATH_bkp_3__21_;
  wire AES_CORE_DATAPATH_bkp_3__22_;
  wire AES_CORE_DATAPATH_bkp_3__23_;
  wire AES_CORE_DATAPATH_bkp_3__24_;
  wire AES_CORE_DATAPATH_bkp_3__25_;
  wire AES_CORE_DATAPATH_bkp_3__26_;
  wire AES_CORE_DATAPATH_bkp_3__27_;
  wire AES_CORE_DATAPATH_bkp_3__28_;
  wire AES_CORE_DATAPATH_bkp_3__29_;
  wire AES_CORE_DATAPATH_bkp_3__2_;
  wire AES_CORE_DATAPATH_bkp_3__30_;
  wire AES_CORE_DATAPATH_bkp_3__31_;
  wire AES_CORE_DATAPATH_bkp_3__3_;
  wire AES_CORE_DATAPATH_bkp_3__4_;
  wire AES_CORE_DATAPATH_bkp_3__5_;
  wire AES_CORE_DATAPATH_bkp_3__6_;
  wire AES_CORE_DATAPATH_bkp_3__7_;
  wire AES_CORE_DATAPATH_bkp_3__8_;
  wire AES_CORE_DATAPATH_bkp_3__9_;
  wire AES_CORE_DATAPATH_col_0__0_;
  wire AES_CORE_DATAPATH_col_0__10_;
  wire AES_CORE_DATAPATH_col_0__11_;
  wire AES_CORE_DATAPATH_col_0__12_;
  wire AES_CORE_DATAPATH_col_0__13_;
  wire AES_CORE_DATAPATH_col_0__14_;
  wire AES_CORE_DATAPATH_col_0__15_;
  wire AES_CORE_DATAPATH_col_0__16_;
  wire AES_CORE_DATAPATH_col_0__17_;
  wire AES_CORE_DATAPATH_col_0__18_;
  wire AES_CORE_DATAPATH_col_0__19_;
  wire AES_CORE_DATAPATH_col_0__1_;
  wire AES_CORE_DATAPATH_col_0__20_;
  wire AES_CORE_DATAPATH_col_0__21_;
  wire AES_CORE_DATAPATH_col_0__22_;
  wire AES_CORE_DATAPATH_col_0__23_;
  wire AES_CORE_DATAPATH_col_0__24_;
  wire AES_CORE_DATAPATH_col_0__25_;
  wire AES_CORE_DATAPATH_col_0__26_;
  wire AES_CORE_DATAPATH_col_0__27_;
  wire AES_CORE_DATAPATH_col_0__28_;
  wire AES_CORE_DATAPATH_col_0__29_;
  wire AES_CORE_DATAPATH_col_0__2_;
  wire AES_CORE_DATAPATH_col_0__30_;
  wire AES_CORE_DATAPATH_col_0__31_;
  wire AES_CORE_DATAPATH_col_0__3_;
  wire AES_CORE_DATAPATH_col_0__4_;
  wire AES_CORE_DATAPATH_col_0__5_;
  wire AES_CORE_DATAPATH_col_0__6_;
  wire AES_CORE_DATAPATH_col_0__7_;
  wire AES_CORE_DATAPATH_col_0__8_;
  wire AES_CORE_DATAPATH_col_0__9_;
  wire AES_CORE_DATAPATH_col_3__0_;
  wire AES_CORE_DATAPATH_col_3__10_;
  wire AES_CORE_DATAPATH_col_3__11_;
  wire AES_CORE_DATAPATH_col_3__12_;
  wire AES_CORE_DATAPATH_col_3__13_;
  wire AES_CORE_DATAPATH_col_3__14_;
  wire AES_CORE_DATAPATH_col_3__15_;
  wire AES_CORE_DATAPATH_col_3__16_;
  wire AES_CORE_DATAPATH_col_3__17_;
  wire AES_CORE_DATAPATH_col_3__18_;
  wire AES_CORE_DATAPATH_col_3__19_;
  wire AES_CORE_DATAPATH_col_3__1_;
  wire AES_CORE_DATAPATH_col_3__20_;
  wire AES_CORE_DATAPATH_col_3__21_;
  wire AES_CORE_DATAPATH_col_3__22_;
  wire AES_CORE_DATAPATH_col_3__23_;
  wire AES_CORE_DATAPATH_col_3__24_;
  wire AES_CORE_DATAPATH_col_3__25_;
  wire AES_CORE_DATAPATH_col_3__26_;
  wire AES_CORE_DATAPATH_col_3__27_;
  wire AES_CORE_DATAPATH_col_3__28_;
  wire AES_CORE_DATAPATH_col_3__29_;
  wire AES_CORE_DATAPATH_col_3__2_;
  wire AES_CORE_DATAPATH_col_3__30_;
  wire AES_CORE_DATAPATH_col_3__31_;
  wire AES_CORE_DATAPATH_col_3__3_;
  wire AES_CORE_DATAPATH_col_3__4_;
  wire AES_CORE_DATAPATH_col_3__5_;
  wire AES_CORE_DATAPATH_col_3__6_;
  wire AES_CORE_DATAPATH_col_3__7_;
  wire AES_CORE_DATAPATH_col_3__8_;
  wire AES_CORE_DATAPATH_col_3__9_;
  wire AES_CORE_DATAPATH_col_en_cnt_unit_pp1_0_;
  wire AES_CORE_DATAPATH_col_en_cnt_unit_pp1_0__FF_INPUT;
  wire AES_CORE_DATAPATH_col_en_cnt_unit_pp1_1_;
  wire AES_CORE_DATAPATH_col_en_cnt_unit_pp1_1__FF_INPUT;
  wire AES_CORE_DATAPATH_col_en_cnt_unit_pp1_2_;
  wire AES_CORE_DATAPATH_col_en_cnt_unit_pp1_2__FF_INPUT;
  wire AES_CORE_DATAPATH_col_en_cnt_unit_pp1_3_;
  wire AES_CORE_DATAPATH_col_en_cnt_unit_pp1_3__FF_INPUT;
  wire AES_CORE_DATAPATH_col_en_cnt_unit_pp2_0_;
  wire AES_CORE_DATAPATH_col_en_cnt_unit_pp2_0__FF_INPUT;
  wire AES_CORE_DATAPATH_col_en_cnt_unit_pp2_1_;
  wire AES_CORE_DATAPATH_col_en_cnt_unit_pp2_1__FF_INPUT;
  wire AES_CORE_DATAPATH_col_en_cnt_unit_pp2_2_;
  wire AES_CORE_DATAPATH_col_en_cnt_unit_pp2_2__FF_INPUT;
  wire AES_CORE_DATAPATH_col_en_cnt_unit_pp2_3_;
  wire AES_CORE_DATAPATH_col_en_cnt_unit_pp2_3__FF_INPUT;
  wire AES_CORE_DATAPATH_col_en_host_0_;
  wire AES_CORE_DATAPATH_col_en_host_1_;
  wire AES_CORE_DATAPATH_col_en_host_2_;
  wire AES_CORE_DATAPATH_col_en_host_3_;
  wire AES_CORE_DATAPATH_col_sel_host_0_;
  wire AES_CORE_DATAPATH_col_sel_host_1_;
  wire AES_CORE_DATAPATH_col_sel_pp1_0_;
  wire AES_CORE_DATAPATH_col_sel_pp1_1_;
  wire AES_CORE_DATAPATH_col_sel_pp2_0_;
  wire AES_CORE_DATAPATH_col_sel_pp2_1_;
  wire AES_CORE_DATAPATH_iv_0__0_;
  wire AES_CORE_DATAPATH_iv_0__10_;
  wire AES_CORE_DATAPATH_iv_0__11_;
  wire AES_CORE_DATAPATH_iv_0__12_;
  wire AES_CORE_DATAPATH_iv_0__13_;
  wire AES_CORE_DATAPATH_iv_0__14_;
  wire AES_CORE_DATAPATH_iv_0__15_;
  wire AES_CORE_DATAPATH_iv_0__16_;
  wire AES_CORE_DATAPATH_iv_0__17_;
  wire AES_CORE_DATAPATH_iv_0__18_;
  wire AES_CORE_DATAPATH_iv_0__19_;
  wire AES_CORE_DATAPATH_iv_0__1_;
  wire AES_CORE_DATAPATH_iv_0__20_;
  wire AES_CORE_DATAPATH_iv_0__21_;
  wire AES_CORE_DATAPATH_iv_0__22_;
  wire AES_CORE_DATAPATH_iv_0__23_;
  wire AES_CORE_DATAPATH_iv_0__24_;
  wire AES_CORE_DATAPATH_iv_0__25_;
  wire AES_CORE_DATAPATH_iv_0__26_;
  wire AES_CORE_DATAPATH_iv_0__27_;
  wire AES_CORE_DATAPATH_iv_0__28_;
  wire AES_CORE_DATAPATH_iv_0__29_;
  wire AES_CORE_DATAPATH_iv_0__2_;
  wire AES_CORE_DATAPATH_iv_0__30_;
  wire AES_CORE_DATAPATH_iv_0__31_;
  wire AES_CORE_DATAPATH_iv_0__3_;
  wire AES_CORE_DATAPATH_iv_0__4_;
  wire AES_CORE_DATAPATH_iv_0__5_;
  wire AES_CORE_DATAPATH_iv_0__6_;
  wire AES_CORE_DATAPATH_iv_0__7_;
  wire AES_CORE_DATAPATH_iv_0__8_;
  wire AES_CORE_DATAPATH_iv_0__9_;
  wire AES_CORE_DATAPATH_iv_1__0_;
  wire AES_CORE_DATAPATH_iv_1__10_;
  wire AES_CORE_DATAPATH_iv_1__11_;
  wire AES_CORE_DATAPATH_iv_1__12_;
  wire AES_CORE_DATAPATH_iv_1__13_;
  wire AES_CORE_DATAPATH_iv_1__14_;
  wire AES_CORE_DATAPATH_iv_1__15_;
  wire AES_CORE_DATAPATH_iv_1__16_;
  wire AES_CORE_DATAPATH_iv_1__17_;
  wire AES_CORE_DATAPATH_iv_1__18_;
  wire AES_CORE_DATAPATH_iv_1__19_;
  wire AES_CORE_DATAPATH_iv_1__1_;
  wire AES_CORE_DATAPATH_iv_1__20_;
  wire AES_CORE_DATAPATH_iv_1__21_;
  wire AES_CORE_DATAPATH_iv_1__22_;
  wire AES_CORE_DATAPATH_iv_1__23_;
  wire AES_CORE_DATAPATH_iv_1__24_;
  wire AES_CORE_DATAPATH_iv_1__25_;
  wire AES_CORE_DATAPATH_iv_1__26_;
  wire AES_CORE_DATAPATH_iv_1__27_;
  wire AES_CORE_DATAPATH_iv_1__28_;
  wire AES_CORE_DATAPATH_iv_1__29_;
  wire AES_CORE_DATAPATH_iv_1__2_;
  wire AES_CORE_DATAPATH_iv_1__30_;
  wire AES_CORE_DATAPATH_iv_1__31_;
  wire AES_CORE_DATAPATH_iv_1__3_;
  wire AES_CORE_DATAPATH_iv_1__4_;
  wire AES_CORE_DATAPATH_iv_1__5_;
  wire AES_CORE_DATAPATH_iv_1__6_;
  wire AES_CORE_DATAPATH_iv_1__7_;
  wire AES_CORE_DATAPATH_iv_1__8_;
  wire AES_CORE_DATAPATH_iv_1__9_;
  wire AES_CORE_DATAPATH_iv_2__0_;
  wire AES_CORE_DATAPATH_iv_2__10_;
  wire AES_CORE_DATAPATH_iv_2__11_;
  wire AES_CORE_DATAPATH_iv_2__12_;
  wire AES_CORE_DATAPATH_iv_2__13_;
  wire AES_CORE_DATAPATH_iv_2__14_;
  wire AES_CORE_DATAPATH_iv_2__15_;
  wire AES_CORE_DATAPATH_iv_2__16_;
  wire AES_CORE_DATAPATH_iv_2__17_;
  wire AES_CORE_DATAPATH_iv_2__18_;
  wire AES_CORE_DATAPATH_iv_2__19_;
  wire AES_CORE_DATAPATH_iv_2__1_;
  wire AES_CORE_DATAPATH_iv_2__20_;
  wire AES_CORE_DATAPATH_iv_2__21_;
  wire AES_CORE_DATAPATH_iv_2__22_;
  wire AES_CORE_DATAPATH_iv_2__23_;
  wire AES_CORE_DATAPATH_iv_2__24_;
  wire AES_CORE_DATAPATH_iv_2__25_;
  wire AES_CORE_DATAPATH_iv_2__26_;
  wire AES_CORE_DATAPATH_iv_2__27_;
  wire AES_CORE_DATAPATH_iv_2__28_;
  wire AES_CORE_DATAPATH_iv_2__29_;
  wire AES_CORE_DATAPATH_iv_2__2_;
  wire AES_CORE_DATAPATH_iv_2__30_;
  wire AES_CORE_DATAPATH_iv_2__31_;
  wire AES_CORE_DATAPATH_iv_2__3_;
  wire AES_CORE_DATAPATH_iv_2__4_;
  wire AES_CORE_DATAPATH_iv_2__5_;
  wire AES_CORE_DATAPATH_iv_2__6_;
  wire AES_CORE_DATAPATH_iv_2__7_;
  wire AES_CORE_DATAPATH_iv_2__8_;
  wire AES_CORE_DATAPATH_iv_2__9_;
  wire AES_CORE_DATAPATH_iv_3__0_;
  wire AES_CORE_DATAPATH_iv_3__10_;
  wire AES_CORE_DATAPATH_iv_3__11_;
  wire AES_CORE_DATAPATH_iv_3__12_;
  wire AES_CORE_DATAPATH_iv_3__13_;
  wire AES_CORE_DATAPATH_iv_3__14_;
  wire AES_CORE_DATAPATH_iv_3__15_;
  wire AES_CORE_DATAPATH_iv_3__16_;
  wire AES_CORE_DATAPATH_iv_3__17_;
  wire AES_CORE_DATAPATH_iv_3__18_;
  wire AES_CORE_DATAPATH_iv_3__19_;
  wire AES_CORE_DATAPATH_iv_3__1_;
  wire AES_CORE_DATAPATH_iv_3__20_;
  wire AES_CORE_DATAPATH_iv_3__21_;
  wire AES_CORE_DATAPATH_iv_3__22_;
  wire AES_CORE_DATAPATH_iv_3__23_;
  wire AES_CORE_DATAPATH_iv_3__24_;
  wire AES_CORE_DATAPATH_iv_3__25_;
  wire AES_CORE_DATAPATH_iv_3__26_;
  wire AES_CORE_DATAPATH_iv_3__27_;
  wire AES_CORE_DATAPATH_iv_3__28_;
  wire AES_CORE_DATAPATH_iv_3__29_;
  wire AES_CORE_DATAPATH_iv_3__2_;
  wire AES_CORE_DATAPATH_iv_3__30_;
  wire AES_CORE_DATAPATH_iv_3__31_;
  wire AES_CORE_DATAPATH_iv_3__3_;
  wire AES_CORE_DATAPATH_iv_3__4_;
  wire AES_CORE_DATAPATH_iv_3__5_;
  wire AES_CORE_DATAPATH_iv_3__6_;
  wire AES_CORE_DATAPATH_iv_3__7_;
  wire AES_CORE_DATAPATH_iv_3__8_;
  wire AES_CORE_DATAPATH_iv_3__9_;
  wire AES_CORE_DATAPATH_key_en_pp1_0_;
  wire AES_CORE_DATAPATH_key_en_pp1_0__FF_INPUT;
  wire AES_CORE_DATAPATH_key_en_pp1_1_;
  wire AES_CORE_DATAPATH_key_en_pp1_1__FF_INPUT;
  wire AES_CORE_DATAPATH_key_en_pp1_2_;
  wire AES_CORE_DATAPATH_key_en_pp1_2__FF_INPUT;
  wire AES_CORE_DATAPATH_key_en_pp1_3_;
  wire AES_CORE_DATAPATH_key_en_pp1_3__FF_INPUT;
  wire AES_CORE_DATAPATH_key_host_0__0_;
  wire AES_CORE_DATAPATH_key_host_0__10_;
  wire AES_CORE_DATAPATH_key_host_0__11_;
  wire AES_CORE_DATAPATH_key_host_0__12_;
  wire AES_CORE_DATAPATH_key_host_0__13_;
  wire AES_CORE_DATAPATH_key_host_0__14_;
  wire AES_CORE_DATAPATH_key_host_0__15_;
  wire AES_CORE_DATAPATH_key_host_0__16_;
  wire AES_CORE_DATAPATH_key_host_0__17_;
  wire AES_CORE_DATAPATH_key_host_0__18_;
  wire AES_CORE_DATAPATH_key_host_0__19_;
  wire AES_CORE_DATAPATH_key_host_0__1_;
  wire AES_CORE_DATAPATH_key_host_0__20_;
  wire AES_CORE_DATAPATH_key_host_0__21_;
  wire AES_CORE_DATAPATH_key_host_0__22_;
  wire AES_CORE_DATAPATH_key_host_0__23_;
  wire AES_CORE_DATAPATH_key_host_0__24_;
  wire AES_CORE_DATAPATH_key_host_0__25_;
  wire AES_CORE_DATAPATH_key_host_0__26_;
  wire AES_CORE_DATAPATH_key_host_0__27_;
  wire AES_CORE_DATAPATH_key_host_0__28_;
  wire AES_CORE_DATAPATH_key_host_0__29_;
  wire AES_CORE_DATAPATH_key_host_0__2_;
  wire AES_CORE_DATAPATH_key_host_0__30_;
  wire AES_CORE_DATAPATH_key_host_0__31_;
  wire AES_CORE_DATAPATH_key_host_0__3_;
  wire AES_CORE_DATAPATH_key_host_0__4_;
  wire AES_CORE_DATAPATH_key_host_0__5_;
  wire AES_CORE_DATAPATH_key_host_0__6_;
  wire AES_CORE_DATAPATH_key_host_0__7_;
  wire AES_CORE_DATAPATH_key_host_0__8_;
  wire AES_CORE_DATAPATH_key_host_0__9_;
  wire AES_CORE_DATAPATH_key_host_1__0_;
  wire AES_CORE_DATAPATH_key_host_1__10_;
  wire AES_CORE_DATAPATH_key_host_1__11_;
  wire AES_CORE_DATAPATH_key_host_1__12_;
  wire AES_CORE_DATAPATH_key_host_1__13_;
  wire AES_CORE_DATAPATH_key_host_1__14_;
  wire AES_CORE_DATAPATH_key_host_1__15_;
  wire AES_CORE_DATAPATH_key_host_1__16_;
  wire AES_CORE_DATAPATH_key_host_1__17_;
  wire AES_CORE_DATAPATH_key_host_1__18_;
  wire AES_CORE_DATAPATH_key_host_1__19_;
  wire AES_CORE_DATAPATH_key_host_1__1_;
  wire AES_CORE_DATAPATH_key_host_1__20_;
  wire AES_CORE_DATAPATH_key_host_1__21_;
  wire AES_CORE_DATAPATH_key_host_1__22_;
  wire AES_CORE_DATAPATH_key_host_1__23_;
  wire AES_CORE_DATAPATH_key_host_1__24_;
  wire AES_CORE_DATAPATH_key_host_1__25_;
  wire AES_CORE_DATAPATH_key_host_1__26_;
  wire AES_CORE_DATAPATH_key_host_1__27_;
  wire AES_CORE_DATAPATH_key_host_1__28_;
  wire AES_CORE_DATAPATH_key_host_1__29_;
  wire AES_CORE_DATAPATH_key_host_1__2_;
  wire AES_CORE_DATAPATH_key_host_1__30_;
  wire AES_CORE_DATAPATH_key_host_1__31_;
  wire AES_CORE_DATAPATH_key_host_1__3_;
  wire AES_CORE_DATAPATH_key_host_1__4_;
  wire AES_CORE_DATAPATH_key_host_1__5_;
  wire AES_CORE_DATAPATH_key_host_1__6_;
  wire AES_CORE_DATAPATH_key_host_1__7_;
  wire AES_CORE_DATAPATH_key_host_1__8_;
  wire AES_CORE_DATAPATH_key_host_1__9_;
  wire AES_CORE_DATAPATH_key_host_2__0_;
  wire AES_CORE_DATAPATH_key_host_2__10_;
  wire AES_CORE_DATAPATH_key_host_2__11_;
  wire AES_CORE_DATAPATH_key_host_2__12_;
  wire AES_CORE_DATAPATH_key_host_2__13_;
  wire AES_CORE_DATAPATH_key_host_2__14_;
  wire AES_CORE_DATAPATH_key_host_2__15_;
  wire AES_CORE_DATAPATH_key_host_2__16_;
  wire AES_CORE_DATAPATH_key_host_2__17_;
  wire AES_CORE_DATAPATH_key_host_2__18_;
  wire AES_CORE_DATAPATH_key_host_2__19_;
  wire AES_CORE_DATAPATH_key_host_2__1_;
  wire AES_CORE_DATAPATH_key_host_2__20_;
  wire AES_CORE_DATAPATH_key_host_2__21_;
  wire AES_CORE_DATAPATH_key_host_2__22_;
  wire AES_CORE_DATAPATH_key_host_2__23_;
  wire AES_CORE_DATAPATH_key_host_2__24_;
  wire AES_CORE_DATAPATH_key_host_2__25_;
  wire AES_CORE_DATAPATH_key_host_2__26_;
  wire AES_CORE_DATAPATH_key_host_2__27_;
  wire AES_CORE_DATAPATH_key_host_2__28_;
  wire AES_CORE_DATAPATH_key_host_2__29_;
  wire AES_CORE_DATAPATH_key_host_2__2_;
  wire AES_CORE_DATAPATH_key_host_2__30_;
  wire AES_CORE_DATAPATH_key_host_2__31_;
  wire AES_CORE_DATAPATH_key_host_2__3_;
  wire AES_CORE_DATAPATH_key_host_2__4_;
  wire AES_CORE_DATAPATH_key_host_2__5_;
  wire AES_CORE_DATAPATH_key_host_2__6_;
  wire AES_CORE_DATAPATH_key_host_2__7_;
  wire AES_CORE_DATAPATH_key_host_2__8_;
  wire AES_CORE_DATAPATH_key_host_2__9_;
  wire AES_CORE_DATAPATH_key_host_3__0_;
  wire AES_CORE_DATAPATH_key_host_3__10_;
  wire AES_CORE_DATAPATH_key_host_3__11_;
  wire AES_CORE_DATAPATH_key_host_3__12_;
  wire AES_CORE_DATAPATH_key_host_3__13_;
  wire AES_CORE_DATAPATH_key_host_3__14_;
  wire AES_CORE_DATAPATH_key_host_3__15_;
  wire AES_CORE_DATAPATH_key_host_3__16_;
  wire AES_CORE_DATAPATH_key_host_3__17_;
  wire AES_CORE_DATAPATH_key_host_3__18_;
  wire AES_CORE_DATAPATH_key_host_3__19_;
  wire AES_CORE_DATAPATH_key_host_3__1_;
  wire AES_CORE_DATAPATH_key_host_3__20_;
  wire AES_CORE_DATAPATH_key_host_3__21_;
  wire AES_CORE_DATAPATH_key_host_3__22_;
  wire AES_CORE_DATAPATH_key_host_3__23_;
  wire AES_CORE_DATAPATH_key_host_3__24_;
  wire AES_CORE_DATAPATH_key_host_3__25_;
  wire AES_CORE_DATAPATH_key_host_3__26_;
  wire AES_CORE_DATAPATH_key_host_3__27_;
  wire AES_CORE_DATAPATH_key_host_3__28_;
  wire AES_CORE_DATAPATH_key_host_3__29_;
  wire AES_CORE_DATAPATH_key_host_3__2_;
  wire AES_CORE_DATAPATH_key_host_3__30_;
  wire AES_CORE_DATAPATH_key_host_3__31_;
  wire AES_CORE_DATAPATH_key_host_3__3_;
  wire AES_CORE_DATAPATH_key_host_3__4_;
  wire AES_CORE_DATAPATH_key_host_3__5_;
  wire AES_CORE_DATAPATH_key_host_3__6_;
  wire AES_CORE_DATAPATH_key_host_3__7_;
  wire AES_CORE_DATAPATH_key_host_3__8_;
  wire AES_CORE_DATAPATH_key_host_3__9_;
  wire AES_CORE_DATAPATH_key_out_sel_pp1_0_;
  wire AES_CORE_DATAPATH_key_out_sel_pp1_1_;
  wire AES_CORE_DATAPATH_key_out_sel_pp2_0_;
  wire AES_CORE_DATAPATH_key_out_sel_pp2_1_;
  wire AES_CORE_DATAPATH_key_sel_pp1;
  wire AES_CORE_DATAPATH_last_round_pp1;
  wire AES_CORE_DATAPATH_last_round_pp2;
  wire AES_CORE_DATAPATH_last_round_pp2_bF_buf0;
  wire AES_CORE_DATAPATH_last_round_pp2_bF_buf1;
  wire AES_CORE_DATAPATH_last_round_pp2_bF_buf2;
  wire AES_CORE_DATAPATH_last_round_pp2_bF_buf3;
  wire AES_CORE_DATAPATH_last_round_pp2_bF_buf4;
  wire AES_CORE_DATAPATH_rk_out_sel;
  wire AES_CORE_DATAPATH_rk_out_sel_pp1;
  wire AES_CORE_DATAPATH_rk_out_sel_pp2;
  wire AES_CORE_DATAPATH_rk_sel_pp1_0_;
  wire AES_CORE_DATAPATH_rk_sel_pp1_1_;
  wire AES_CORE_DATAPATH_rk_sel_pp2_0_;
  wire AES_CORE_DATAPATH_rk_sel_pp2_1_;
  wire AES_CORE_DATAPATH_sbox_pp2_0__FF_INPUT;
  wire AES_CORE_DATAPATH_sbox_pp2_10__FF_INPUT;
  wire AES_CORE_DATAPATH_sbox_pp2_11__FF_INPUT;
  wire AES_CORE_DATAPATH_sbox_pp2_12__FF_INPUT;
  wire AES_CORE_DATAPATH_sbox_pp2_13__FF_INPUT;
  wire AES_CORE_DATAPATH_sbox_pp2_14__FF_INPUT;
  wire AES_CORE_DATAPATH_sbox_pp2_15__FF_INPUT;
  wire AES_CORE_DATAPATH_sbox_pp2_16__FF_INPUT;
  wire AES_CORE_DATAPATH_sbox_pp2_17__FF_INPUT;
  wire AES_CORE_DATAPATH_sbox_pp2_18__FF_INPUT;
  wire AES_CORE_DATAPATH_sbox_pp2_19__FF_INPUT;
  wire AES_CORE_DATAPATH_sbox_pp2_1__FF_INPUT;
  wire AES_CORE_DATAPATH_sbox_pp2_20__FF_INPUT;
  wire AES_CORE_DATAPATH_sbox_pp2_21__FF_INPUT;
  wire AES_CORE_DATAPATH_sbox_pp2_22__FF_INPUT;
  wire AES_CORE_DATAPATH_sbox_pp2_23__FF_INPUT;
  wire AES_CORE_DATAPATH_sbox_pp2_24__FF_INPUT;
  wire AES_CORE_DATAPATH_sbox_pp2_25__FF_INPUT;
  wire AES_CORE_DATAPATH_sbox_pp2_26__FF_INPUT;
  wire AES_CORE_DATAPATH_sbox_pp2_27__FF_INPUT;
  wire AES_CORE_DATAPATH_sbox_pp2_28__FF_INPUT;
  wire AES_CORE_DATAPATH_sbox_pp2_29__FF_INPUT;
  wire AES_CORE_DATAPATH_sbox_pp2_2__FF_INPUT;
  wire AES_CORE_DATAPATH_sbox_pp2_30__FF_INPUT;
  wire AES_CORE_DATAPATH_sbox_pp2_31__FF_INPUT;
  wire AES_CORE_DATAPATH_sbox_pp2_3__FF_INPUT;
  wire AES_CORE_DATAPATH_sbox_pp2_4__FF_INPUT;
  wire AES_CORE_DATAPATH_sbox_pp2_5__FF_INPUT;
  wire AES_CORE_DATAPATH_sbox_pp2_6__FF_INPUT;
  wire AES_CORE_DATAPATH_sbox_pp2_7__FF_INPUT;
  wire AES_CORE_DATAPATH_sbox_pp2_8__FF_INPUT;
  wire AES_CORE_DATAPATH_sbox_pp2_9__FF_INPUT;
  wire _abc_15830_n11_1;
  wire _abc_15830_n12_1;
  wire _abc_15830_n13_1;
  wire _abc_15830_n15;
  wire _auto_iopadmap_cc_313_execute_26881_0_;
  wire _auto_iopadmap_cc_313_execute_26881_10_;
  wire _auto_iopadmap_cc_313_execute_26881_11_;
  wire _auto_iopadmap_cc_313_execute_26881_12_;
  wire _auto_iopadmap_cc_313_execute_26881_13_;
  wire _auto_iopadmap_cc_313_execute_26881_14_;
  wire _auto_iopadmap_cc_313_execute_26881_15_;
  wire _auto_iopadmap_cc_313_execute_26881_16_;
  wire _auto_iopadmap_cc_313_execute_26881_17_;
  wire _auto_iopadmap_cc_313_execute_26881_18_;
  wire _auto_iopadmap_cc_313_execute_26881_19_;
  wire _auto_iopadmap_cc_313_execute_26881_1_;
  wire _auto_iopadmap_cc_313_execute_26881_20_;
  wire _auto_iopadmap_cc_313_execute_26881_21_;
  wire _auto_iopadmap_cc_313_execute_26881_22_;
  wire _auto_iopadmap_cc_313_execute_26881_23_;
  wire _auto_iopadmap_cc_313_execute_26881_24_;
  wire _auto_iopadmap_cc_313_execute_26881_25_;
  wire _auto_iopadmap_cc_313_execute_26881_26_;
  wire _auto_iopadmap_cc_313_execute_26881_27_;
  wire _auto_iopadmap_cc_313_execute_26881_28_;
  wire _auto_iopadmap_cc_313_execute_26881_29_;
  wire _auto_iopadmap_cc_313_execute_26881_2_;
  wire _auto_iopadmap_cc_313_execute_26881_30_;
  wire _auto_iopadmap_cc_313_execute_26881_31_;
  wire _auto_iopadmap_cc_313_execute_26881_3_;
  wire _auto_iopadmap_cc_313_execute_26881_4_;
  wire _auto_iopadmap_cc_313_execute_26881_5_;
  wire _auto_iopadmap_cc_313_execute_26881_6_;
  wire _auto_iopadmap_cc_313_execute_26881_7_;
  wire _auto_iopadmap_cc_313_execute_26881_8_;
  wire _auto_iopadmap_cc_313_execute_26881_9_;
  wire _auto_iopadmap_cc_313_execute_26914;
  wire _auto_iopadmap_cc_313_execute_26916_0_;
  wire _auto_iopadmap_cc_313_execute_26916_10_;
  wire _auto_iopadmap_cc_313_execute_26916_11_;
  wire _auto_iopadmap_cc_313_execute_26916_12_;
  wire _auto_iopadmap_cc_313_execute_26916_13_;
  wire _auto_iopadmap_cc_313_execute_26916_14_;
  wire _auto_iopadmap_cc_313_execute_26916_15_;
  wire _auto_iopadmap_cc_313_execute_26916_16_;
  wire _auto_iopadmap_cc_313_execute_26916_17_;
  wire _auto_iopadmap_cc_313_execute_26916_18_;
  wire _auto_iopadmap_cc_313_execute_26916_19_;
  wire _auto_iopadmap_cc_313_execute_26916_1_;
  wire _auto_iopadmap_cc_313_execute_26916_20_;
  wire _auto_iopadmap_cc_313_execute_26916_21_;
  wire _auto_iopadmap_cc_313_execute_26916_22_;
  wire _auto_iopadmap_cc_313_execute_26916_23_;
  wire _auto_iopadmap_cc_313_execute_26916_24_;
  wire _auto_iopadmap_cc_313_execute_26916_25_;
  wire _auto_iopadmap_cc_313_execute_26916_26_;
  wire _auto_iopadmap_cc_313_execute_26916_27_;
  wire _auto_iopadmap_cc_313_execute_26916_28_;
  wire _auto_iopadmap_cc_313_execute_26916_29_;
  wire _auto_iopadmap_cc_313_execute_26916_2_;
  wire _auto_iopadmap_cc_313_execute_26916_30_;
  wire _auto_iopadmap_cc_313_execute_26916_31_;
  wire _auto_iopadmap_cc_313_execute_26916_3_;
  wire _auto_iopadmap_cc_313_execute_26916_4_;
  wire _auto_iopadmap_cc_313_execute_26916_5_;
  wire _auto_iopadmap_cc_313_execute_26916_6_;
  wire _auto_iopadmap_cc_313_execute_26916_7_;
  wire _auto_iopadmap_cc_313_execute_26916_8_;
  wire _auto_iopadmap_cc_313_execute_26916_9_;
  wire _auto_iopadmap_cc_313_execute_26949_0_;
  wire _auto_iopadmap_cc_313_execute_26949_10_;
  wire _auto_iopadmap_cc_313_execute_26949_11_;
  wire _auto_iopadmap_cc_313_execute_26949_12_;
  wire _auto_iopadmap_cc_313_execute_26949_13_;
  wire _auto_iopadmap_cc_313_execute_26949_14_;
  wire _auto_iopadmap_cc_313_execute_26949_15_;
  wire _auto_iopadmap_cc_313_execute_26949_16_;
  wire _auto_iopadmap_cc_313_execute_26949_17_;
  wire _auto_iopadmap_cc_313_execute_26949_18_;
  wire _auto_iopadmap_cc_313_execute_26949_19_;
  wire _auto_iopadmap_cc_313_execute_26949_1_;
  wire _auto_iopadmap_cc_313_execute_26949_20_;
  wire _auto_iopadmap_cc_313_execute_26949_21_;
  wire _auto_iopadmap_cc_313_execute_26949_22_;
  wire _auto_iopadmap_cc_313_execute_26949_23_;
  wire _auto_iopadmap_cc_313_execute_26949_24_;
  wire _auto_iopadmap_cc_313_execute_26949_25_;
  wire _auto_iopadmap_cc_313_execute_26949_26_;
  wire _auto_iopadmap_cc_313_execute_26949_27_;
  wire _auto_iopadmap_cc_313_execute_26949_28_;
  wire _auto_iopadmap_cc_313_execute_26949_29_;
  wire _auto_iopadmap_cc_313_execute_26949_2_;
  wire _auto_iopadmap_cc_313_execute_26949_30_;
  wire _auto_iopadmap_cc_313_execute_26949_31_;
  wire _auto_iopadmap_cc_313_execute_26949_3_;
  wire _auto_iopadmap_cc_313_execute_26949_4_;
  wire _auto_iopadmap_cc_313_execute_26949_5_;
  wire _auto_iopadmap_cc_313_execute_26949_6_;
  wire _auto_iopadmap_cc_313_execute_26949_7_;
  wire _auto_iopadmap_cc_313_execute_26949_8_;
  wire _auto_iopadmap_cc_313_execute_26949_9_;
  input \addr[0] ;
  input \addr[1] ;
  input \aes_mode[0] ;
  input \aes_mode[1] ;
  input \bus_in[0] ;
  input \bus_in[10] ;
  input \bus_in[11] ;
  input \bus_in[12] ;
  input \bus_in[13] ;
  input \bus_in[14] ;
  input \bus_in[15] ;
  input \bus_in[16] ;
  input \bus_in[17] ;
  input \bus_in[18] ;
  input \bus_in[19] ;
  input \bus_in[1] ;
  input \bus_in[20] ;
  input \bus_in[21] ;
  input \bus_in[22] ;
  input \bus_in[23] ;
  input \bus_in[24] ;
  input \bus_in[25] ;
  input \bus_in[26] ;
  input \bus_in[27] ;
  input \bus_in[28] ;
  input \bus_in[29] ;
  input \bus_in[2] ;
  input \bus_in[30] ;
  input \bus_in[31] ;
  input \bus_in[3] ;
  input \bus_in[4] ;
  input \bus_in[5] ;
  input \bus_in[6] ;
  input \bus_in[7] ;
  input \bus_in[8] ;
  input \bus_in[9] ;
  input clk;
  wire clk_bF_buf0;
  wire clk_bF_buf1;
  wire clk_bF_buf10;
  wire clk_bF_buf11;
  wire clk_bF_buf12;
  wire clk_bF_buf13;
  wire clk_bF_buf14;
  wire clk_bF_buf15;
  wire clk_bF_buf16;
  wire clk_bF_buf17;
  wire clk_bF_buf18;
  wire clk_bF_buf19;
  wire clk_bF_buf2;
  wire clk_bF_buf20;
  wire clk_bF_buf21;
  wire clk_bF_buf22;
  wire clk_bF_buf23;
  wire clk_bF_buf24;
  wire clk_bF_buf25;
  wire clk_bF_buf26;
  wire clk_bF_buf27;
  wire clk_bF_buf28;
  wire clk_bF_buf29;
  wire clk_bF_buf3;
  wire clk_bF_buf30;
  wire clk_bF_buf31;
  wire clk_bF_buf32;
  wire clk_bF_buf33;
  wire clk_bF_buf34;
  wire clk_bF_buf35;
  wire clk_bF_buf36;
  wire clk_bF_buf37;
  wire clk_bF_buf38;
  wire clk_bF_buf39;
  wire clk_bF_buf4;
  wire clk_bF_buf40;
  wire clk_bF_buf41;
  wire clk_bF_buf42;
  wire clk_bF_buf43;
  wire clk_bF_buf44;
  wire clk_bF_buf45;
  wire clk_bF_buf46;
  wire clk_bF_buf47;
  wire clk_bF_buf48;
  wire clk_bF_buf49;
  wire clk_bF_buf5;
  wire clk_bF_buf50;
  wire clk_bF_buf51;
  wire clk_bF_buf52;
  wire clk_bF_buf53;
  wire clk_bF_buf54;
  wire clk_bF_buf55;
  wire clk_bF_buf56;
  wire clk_bF_buf57;
  wire clk_bF_buf58;
  wire clk_bF_buf59;
  wire clk_bF_buf6;
  wire clk_bF_buf60;
  wire clk_bF_buf61;
  wire clk_bF_buf62;
  wire clk_bF_buf63;
  wire clk_bF_buf64;
  wire clk_bF_buf65;
  wire clk_bF_buf66;
  wire clk_bF_buf67;
  wire clk_bF_buf68;
  wire clk_bF_buf69;
  wire clk_bF_buf7;
  wire clk_bF_buf70;
  wire clk_bF_buf71;
  wire clk_bF_buf72;
  wire clk_bF_buf73;
  wire clk_bF_buf74;
  wire clk_bF_buf75;
  wire clk_bF_buf76;
  wire clk_bF_buf77;
  wire clk_bF_buf78;
  wire clk_bF_buf79;
  wire clk_bF_buf8;
  wire clk_bF_buf80;
  wire clk_bF_buf81;
  wire clk_bF_buf82;
  wire clk_bF_buf83;
  wire clk_bF_buf84;
  wire clk_bF_buf85;
  wire clk_bF_buf86;
  wire clk_bF_buf87;
  wire clk_bF_buf88;
  wire clk_bF_buf89;
  wire clk_bF_buf9;
  wire clk_bF_buf90;
  wire clk_bF_buf91;
  wire clk_bF_buf92;
  wire clk_hier0_bF_buf0;
  wire clk_hier0_bF_buf1;
  wire clk_hier0_bF_buf2;
  wire clk_hier0_bF_buf3;
  wire clk_hier0_bF_buf4;
  wire clk_hier0_bF_buf5;
  wire clk_hier0_bF_buf6;
  wire clk_hier0_bF_buf7;
  wire clk_hier0_bF_buf8;
  output \col_out[0] ;
  output \col_out[10] ;
  output \col_out[11] ;
  output \col_out[12] ;
  output \col_out[13] ;
  output \col_out[14] ;
  output \col_out[15] ;
  output \col_out[16] ;
  output \col_out[17] ;
  output \col_out[18] ;
  output \col_out[19] ;
  output \col_out[1] ;
  output \col_out[20] ;
  output \col_out[21] ;
  output \col_out[22] ;
  output \col_out[23] ;
  output \col_out[24] ;
  output \col_out[25] ;
  output \col_out[26] ;
  output \col_out[27] ;
  output \col_out[28] ;
  output \col_out[29] ;
  output \col_out[2] ;
  output \col_out[30] ;
  output \col_out[31] ;
  output \col_out[3] ;
  output \col_out[4] ;
  output \col_out[5] ;
  output \col_out[6] ;
  output \col_out[7] ;
  output \col_out[8] ;
  output \col_out[9] ;
  input \data_type[0] ;
  input \data_type[1] ;
  input disable_core;
  output end_aes;
  input first_block;
  input \iv_en[0] ;
  input \iv_en[1] ;
  input \iv_en[2] ;
  input \iv_en[3] ;
  wire iv_en_0_bF_buf0;
  wire iv_en_0_bF_buf1;
  wire iv_en_0_bF_buf2;
  wire iv_en_0_bF_buf3;
  wire iv_en_0_bF_buf4;
  wire iv_en_1_bF_buf0;
  wire iv_en_1_bF_buf1;
  wire iv_en_1_bF_buf2;
  wire iv_en_1_bF_buf3;
  wire iv_en_1_bF_buf4;
  wire iv_en_2_bF_buf0;
  wire iv_en_2_bF_buf1;
  wire iv_en_2_bF_buf2;
  wire iv_en_2_bF_buf3;
  wire iv_en_2_bF_buf4;
  output \iv_out[0] ;
  output \iv_out[10] ;
  output \iv_out[11] ;
  output \iv_out[12] ;
  output \iv_out[13] ;
  output \iv_out[14] ;
  output \iv_out[15] ;
  output \iv_out[16] ;
  output \iv_out[17] ;
  output \iv_out[18] ;
  output \iv_out[19] ;
  output \iv_out[1] ;
  output \iv_out[20] ;
  output \iv_out[21] ;
  output \iv_out[22] ;
  output \iv_out[23] ;
  output \iv_out[24] ;
  output \iv_out[25] ;
  output \iv_out[26] ;
  output \iv_out[27] ;
  output \iv_out[28] ;
  output \iv_out[29] ;
  output \iv_out[2] ;
  output \iv_out[30] ;
  output \iv_out[31] ;
  output \iv_out[3] ;
  output \iv_out[4] ;
  output \iv_out[5] ;
  output \iv_out[6] ;
  output \iv_out[7] ;
  output \iv_out[8] ;
  output \iv_out[9] ;
  input \iv_sel_rd[0] ;
  input \iv_sel_rd[1] ;
  input \iv_sel_rd[2] ;
  input \iv_sel_rd[3] ;
  input \key_en[0] ;
  input \key_en[1] ;
  input \key_en[2] ;
  input \key_en[3] ;
  wire key_en_0_bF_buf0;
  wire key_en_0_bF_buf1;
  wire key_en_0_bF_buf2;
  wire key_en_0_bF_buf3;
  wire key_en_0_bF_buf4;
  wire key_en_1_bF_buf0;
  wire key_en_1_bF_buf1;
  wire key_en_1_bF_buf2;
  wire key_en_1_bF_buf3;
  wire key_en_1_bF_buf4;
  wire key_en_2_bF_buf0;
  wire key_en_2_bF_buf1;
  wire key_en_2_bF_buf2;
  wire key_en_2_bF_buf3;
  wire key_en_2_bF_buf4;
  wire key_en_3_bF_buf0;
  wire key_en_3_bF_buf1;
  wire key_en_3_bF_buf2;
  wire key_en_3_bF_buf3;
  wire key_en_3_bF_buf4;
  output \key_out[0] ;
  output \key_out[10] ;
  output \key_out[11] ;
  output \key_out[12] ;
  output \key_out[13] ;
  output \key_out[14] ;
  output \key_out[15] ;
  output \key_out[16] ;
  output \key_out[17] ;
  output \key_out[18] ;
  output \key_out[19] ;
  output \key_out[1] ;
  output \key_out[20] ;
  output \key_out[21] ;
  output \key_out[22] ;
  output \key_out[23] ;
  output \key_out[24] ;
  output \key_out[25] ;
  output \key_out[26] ;
  output \key_out[27] ;
  output \key_out[28] ;
  output \key_out[29] ;
  output \key_out[2] ;
  output \key_out[30] ;
  output \key_out[31] ;
  output \key_out[3] ;
  output \key_out[4] ;
  output \key_out[5] ;
  output \key_out[6] ;
  output \key_out[7] ;
  output \key_out[8] ;
  output \key_out[9] ;
  input \key_sel_rd[0] ;
  input \key_sel_rd[1] ;
  input \op_mode[0] ;
  input \op_mode[1] ;
  input read_en;
  input rst_n;
  wire rst_n_bF_buf0;
  wire rst_n_bF_buf1;
  wire rst_n_bF_buf10;
  wire rst_n_bF_buf11;
  wire rst_n_bF_buf12;
  wire rst_n_bF_buf13;
  wire rst_n_bF_buf14;
  wire rst_n_bF_buf15;
  wire rst_n_bF_buf16;
  wire rst_n_bF_buf17;
  wire rst_n_bF_buf18;
  wire rst_n_bF_buf19;
  wire rst_n_bF_buf2;
  wire rst_n_bF_buf20;
  wire rst_n_bF_buf21;
  wire rst_n_bF_buf22;
  wire rst_n_bF_buf23;
  wire rst_n_bF_buf24;
  wire rst_n_bF_buf25;
  wire rst_n_bF_buf26;
  wire rst_n_bF_buf27;
  wire rst_n_bF_buf28;
  wire rst_n_bF_buf29;
  wire rst_n_bF_buf3;
  wire rst_n_bF_buf30;
  wire rst_n_bF_buf31;
  wire rst_n_bF_buf32;
  wire rst_n_bF_buf33;
  wire rst_n_bF_buf34;
  wire rst_n_bF_buf35;
  wire rst_n_bF_buf36;
  wire rst_n_bF_buf37;
  wire rst_n_bF_buf38;
  wire rst_n_bF_buf39;
  wire rst_n_bF_buf4;
  wire rst_n_bF_buf40;
  wire rst_n_bF_buf41;
  wire rst_n_bF_buf42;
  wire rst_n_bF_buf43;
  wire rst_n_bF_buf44;
  wire rst_n_bF_buf45;
  wire rst_n_bF_buf46;
  wire rst_n_bF_buf47;
  wire rst_n_bF_buf48;
  wire rst_n_bF_buf49;
  wire rst_n_bF_buf5;
  wire rst_n_bF_buf50;
  wire rst_n_bF_buf51;
  wire rst_n_bF_buf52;
  wire rst_n_bF_buf53;
  wire rst_n_bF_buf54;
  wire rst_n_bF_buf55;
  wire rst_n_bF_buf56;
  wire rst_n_bF_buf57;
  wire rst_n_bF_buf58;
  wire rst_n_bF_buf59;
  wire rst_n_bF_buf6;
  wire rst_n_bF_buf60;
  wire rst_n_bF_buf61;
  wire rst_n_bF_buf62;
  wire rst_n_bF_buf63;
  wire rst_n_bF_buf64;
  wire rst_n_bF_buf65;
  wire rst_n_bF_buf66;
  wire rst_n_bF_buf67;
  wire rst_n_bF_buf68;
  wire rst_n_bF_buf69;
  wire rst_n_bF_buf7;
  wire rst_n_bF_buf70;
  wire rst_n_bF_buf71;
  wire rst_n_bF_buf72;
  wire rst_n_bF_buf73;
  wire rst_n_bF_buf74;
  wire rst_n_bF_buf75;
  wire rst_n_bF_buf76;
  wire rst_n_bF_buf77;
  wire rst_n_bF_buf78;
  wire rst_n_bF_buf79;
  wire rst_n_bF_buf8;
  wire rst_n_bF_buf80;
  wire rst_n_bF_buf81;
  wire rst_n_bF_buf82;
  wire rst_n_bF_buf83;
  wire rst_n_bF_buf84;
  wire rst_n_bF_buf85;
  wire rst_n_bF_buf86;
  wire rst_n_bF_buf9;
  wire rst_n_hier0_bF_buf0;
  wire rst_n_hier0_bF_buf1;
  wire rst_n_hier0_bF_buf2;
  wire rst_n_hier0_bF_buf3;
  wire rst_n_hier0_bF_buf4;
  wire rst_n_hier0_bF_buf5;
  wire rst_n_hier0_bF_buf6;
  wire rst_n_hier0_bF_buf7;
  wire rst_n_hier0_bF_buf8;
  input start;
  input write_en;
  AND2X2 AND2X2_1 ( .A(_abc_15830_n12_1), .B(write_en), .Y(_abc_15830_n13_1) );
  AND2X2 AND2X2_10 ( .A(AES_CORE_CONTROL_UNIT_rd_count_1_), .B(AES_CORE_CONTROL_UNIT_rd_count_3_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n82_1) );
  AND2X2 AND2X2_100 ( .A(AES_CORE_DATAPATH__abc_16259_n2457_1), .B(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_0_), .Y(AES_CORE_DATAPATH__abc_16259_n2464) );
  AND2X2 AND2X2_1000 ( .A(_auto_iopadmap_cc_313_execute_26949_22_), .B(AES_CORE_DATAPATH__abc_16259_n4386), .Y(AES_CORE_DATAPATH__abc_16259_n4387) );
  AND2X2 AND2X2_1001 ( .A(AES_CORE_DATAPATH__abc_16259_n4388), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_6_), .Y(AES_CORE_DATAPATH__abc_16259_n4389) );
  AND2X2 AND2X2_1002 ( .A(AES_CORE_DATAPATH__abc_16259_n4391_1), .B(AES_CORE_DATAPATH__abc_16259_n4385_1), .Y(AES_CORE_DATAPATH_sbox_pp2_22__FF_INPUT) );
  AND2X2 AND2X2_1003 ( .A(_auto_iopadmap_cc_313_execute_26949_23_), .B(AES_CORE_DATAPATH__abc_16259_n4394), .Y(AES_CORE_DATAPATH__abc_16259_n4395) );
  AND2X2 AND2X2_1004 ( .A(AES_CORE_DATAPATH__abc_16259_n4396), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_7_), .Y(AES_CORE_DATAPATH__abc_16259_n4397) );
  AND2X2 AND2X2_1005 ( .A(AES_CORE_DATAPATH__abc_16259_n4399_1), .B(AES_CORE_DATAPATH__abc_16259_n4393_1), .Y(AES_CORE_DATAPATH_sbox_pp2_23__FF_INPUT) );
  AND2X2 AND2X2_1006 ( .A(_auto_iopadmap_cc_313_execute_26949_24_), .B(AES_CORE_DATAPATH__abc_16259_n4402), .Y(AES_CORE_DATAPATH__abc_16259_n4403) );
  AND2X2 AND2X2_1007 ( .A(AES_CORE_DATAPATH__abc_16259_n4404), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_1_2_), .Y(AES_CORE_DATAPATH__abc_16259_n4405) );
  AND2X2 AND2X2_1008 ( .A(AES_CORE_DATAPATH__abc_16259_n4407_1), .B(AES_CORE_DATAPATH__abc_16259_n4401_1), .Y(AES_CORE_DATAPATH_sbox_pp2_24__FF_INPUT) );
  AND2X2 AND2X2_1009 ( .A(_auto_iopadmap_cc_313_execute_26949_25_), .B(AES_CORE_DATAPATH__abc_16259_n4410), .Y(AES_CORE_DATAPATH__abc_16259_n4411) );
  AND2X2 AND2X2_101 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk_bF_buf0), .B(AES_CORE_CONTROL_UNIT_col_en_0_), .Y(AES_CORE_DATAPATH__abc_16259_n2465_1) );
  AND2X2 AND2X2_1010 ( .A(AES_CORE_DATAPATH__abc_16259_n4412), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_1_), .Y(AES_CORE_DATAPATH__abc_16259_n4413) );
  AND2X2 AND2X2_1011 ( .A(AES_CORE_DATAPATH__abc_16259_n4415_1), .B(AES_CORE_DATAPATH__abc_16259_n4409_1), .Y(AES_CORE_DATAPATH_sbox_pp2_25__FF_INPUT) );
  AND2X2 AND2X2_1012 ( .A(AES_CORE_DATAPATH__abc_16259_n2807_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_26_), .Y(AES_CORE_DATAPATH__abc_16259_n4417_1) );
  AND2X2 AND2X2_1013 ( .A(AES_CORE_DATAPATH__abc_16259_n4421), .B(AES_CORE_DATAPATH__abc_16259_n2804_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n4422_1) );
  AND2X2 AND2X2_1014 ( .A(AES_CORE_DATAPATH__abc_16259_n4422_1), .B(AES_CORE_DATAPATH__abc_16259_n4420), .Y(AES_CORE_DATAPATH__abc_16259_n4423_1) );
  AND2X2 AND2X2_1015 ( .A(_auto_iopadmap_cc_313_execute_26949_27_), .B(AES_CORE_DATAPATH__abc_16259_n4426), .Y(AES_CORE_DATAPATH__abc_16259_n4427) );
  AND2X2 AND2X2_1016 ( .A(AES_CORE_DATAPATH__abc_16259_n4428), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_3_), .Y(AES_CORE_DATAPATH__abc_16259_n4429) );
  AND2X2 AND2X2_1017 ( .A(AES_CORE_DATAPATH__abc_16259_n4431_1), .B(AES_CORE_DATAPATH__abc_16259_n4425_1), .Y(AES_CORE_DATAPATH_sbox_pp2_27__FF_INPUT) );
  AND2X2 AND2X2_1018 ( .A(_auto_iopadmap_cc_313_execute_26949_28_), .B(AES_CORE_DATAPATH__abc_16259_n4434), .Y(AES_CORE_DATAPATH__abc_16259_n4435) );
  AND2X2 AND2X2_1019 ( .A(AES_CORE_DATAPATH__abc_16259_n4436), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_4_), .Y(AES_CORE_DATAPATH__abc_16259_n4437) );
  AND2X2 AND2X2_102 ( .A(AES_CORE_DATAPATH__abc_16259_n2463_1), .B(AES_CORE_DATAPATH__abc_16259_n2468), .Y(AES_CORE_DATAPATH__abc_16259_n2469_1) );
  AND2X2 AND2X2_1020 ( .A(AES_CORE_DATAPATH__abc_16259_n4439), .B(AES_CORE_DATAPATH__abc_16259_n4433_1), .Y(AES_CORE_DATAPATH_sbox_pp2_28__FF_INPUT) );
  AND2X2 AND2X2_1021 ( .A(_auto_iopadmap_cc_313_execute_26949_29_), .B(AES_CORE_DATAPATH__abc_16259_n4442), .Y(AES_CORE_DATAPATH__abc_16259_n4443_1) );
  AND2X2 AND2X2_1022 ( .A(AES_CORE_DATAPATH__abc_16259_n4444_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_5_), .Y(AES_CORE_DATAPATH__abc_16259_n4445_1) );
  AND2X2 AND2X2_1023 ( .A(AES_CORE_DATAPATH__abc_16259_n4447_1), .B(AES_CORE_DATAPATH__abc_16259_n4441), .Y(AES_CORE_DATAPATH_sbox_pp2_29__FF_INPUT) );
  AND2X2 AND2X2_1024 ( .A(_auto_iopadmap_cc_313_execute_26949_30_), .B(AES_CORE_DATAPATH__abc_16259_n4450_1), .Y(AES_CORE_DATAPATH__abc_16259_n4451_1) );
  AND2X2 AND2X2_1025 ( .A(AES_CORE_DATAPATH__abc_16259_n4452_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_6_), .Y(AES_CORE_DATAPATH__abc_16259_n4453_1) );
  AND2X2 AND2X2_1026 ( .A(AES_CORE_DATAPATH__abc_16259_n4455_1), .B(AES_CORE_DATAPATH__abc_16259_n4449_1), .Y(AES_CORE_DATAPATH_sbox_pp2_30__FF_INPUT) );
  AND2X2 AND2X2_1027 ( .A(_auto_iopadmap_cc_313_execute_26949_31_), .B(AES_CORE_DATAPATH__abc_16259_n4458_1), .Y(AES_CORE_DATAPATH__abc_16259_n4459_1) );
  AND2X2 AND2X2_1028 ( .A(AES_CORE_DATAPATH__abc_16259_n4460_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_7_), .Y(AES_CORE_DATAPATH__abc_16259_n4461_1) );
  AND2X2 AND2X2_1029 ( .A(AES_CORE_DATAPATH__abc_16259_n4463_1), .B(AES_CORE_DATAPATH__abc_16259_n4457_1), .Y(AES_CORE_DATAPATH_sbox_pp2_31__FF_INPUT) );
  AND2X2 AND2X2_103 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf7), .B(AES_CORE_DATAPATH_iv_0__0_), .Y(AES_CORE_DATAPATH__abc_16259_n2470) );
  AND2X2 AND2X2_1030 ( .A(AES_CORE_CONTROL_UNIT_bypass_key_en), .B(AES_CORE_CONTROL_UNIT_key_en_0_), .Y(AES_CORE_DATAPATH__abc_16259_n4466_1) );
  AND2X2 AND2X2_1031 ( .A(AES_CORE_DATAPATH__abc_16259_n4468_1_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n4469_1), .Y(AES_CORE_DATAPATH__abc_16259_n4470_1) );
  AND2X2 AND2X2_1032 ( .A(AES_CORE_DATAPATH__abc_16259_n2806_1), .B(AES_CORE_DATAPATH_key_en_pp1_0_), .Y(AES_CORE_DATAPATH__abc_16259_n4471_1) );
  AND2X2 AND2X2_1033 ( .A(AES_CORE_DATAPATH__abc_16259_n4472_1), .B(AES_CORE_DATAPATH__abc_16259_n4470_1), .Y(AES_CORE_DATAPATH__abc_16259_n4473_1) );
  AND2X2 AND2X2_1034 ( .A(AES_CORE_DATAPATH__abc_16259_n4473_1), .B(AES_CORE_DATAPATH__abc_16259_n4467_1), .Y(AES_CORE_DATAPATH__abc_16259_n4474_1) );
  AND2X2 AND2X2_1035 ( .A(AES_CORE_DATAPATH__abc_16259_n2806_1), .B(AES_CORE_DATAPATH_key_sel_pp1), .Y(AES_CORE_DATAPATH__abc_16259_n4476_1) );
  AND2X2 AND2X2_1036 ( .A(AES_CORE_CONTROL_UNIT_bypass_key_en), .B(AES_CORE_CONTROL_UNIT_key_sel), .Y(AES_CORE_DATAPATH__abc_16259_n4477_1) );
  AND2X2 AND2X2_1037 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf10), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_96_), .Y(AES_CORE_DATAPATH__abc_16259_n4479_1) );
  AND2X2 AND2X2_1038 ( .A(key_en_0_bF_buf3), .B(\bus_in[0] ), .Y(AES_CORE_DATAPATH__abc_16259_n4481_1) );
  AND2X2 AND2X2_1039 ( .A(AES_CORE_DATAPATH__abc_16259_n4468_1_bF_buf3), .B(AES_CORE_DATAPATH_key_host_0__0_), .Y(AES_CORE_DATAPATH__abc_16259_n4482_1) );
  AND2X2 AND2X2_104 ( .A(AES_CORE_DATAPATH__abc_16259_n2457_1), .B(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_2_), .Y(AES_CORE_DATAPATH__abc_16259_n2471_1) );
  AND2X2 AND2X2_1040 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf10), .B(AES_CORE_DATAPATH__abc_16259_n4483_1), .Y(AES_CORE_DATAPATH__abc_16259_n4484_1) );
  AND2X2 AND2X2_1041 ( .A(AES_CORE_DATAPATH__abc_16259_n4485_1), .B(AES_CORE_DATAPATH__abc_16259_n4475_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n4486_1) );
  AND2X2 AND2X2_1042 ( .A(AES_CORE_DATAPATH__abc_16259_n4474_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__0_), .Y(AES_CORE_DATAPATH__abc_16259_n4487_1) );
  AND2X2 AND2X2_1043 ( .A(AES_CORE_DATAPATH__abc_16259_n4468_1_bF_buf2), .B(AES_CORE_DATAPATH_key_host_0__1_), .Y(AES_CORE_DATAPATH__abc_16259_n4490_1) );
  AND2X2 AND2X2_1044 ( .A(key_en_0_bF_buf2), .B(\bus_in[1] ), .Y(AES_CORE_DATAPATH__abc_16259_n4491_1) );
  AND2X2 AND2X2_1045 ( .A(AES_CORE_DATAPATH__abc_16259_n4489_1), .B(AES_CORE_DATAPATH__abc_16259_n4493_1), .Y(AES_CORE_DATAPATH__abc_16259_n4494_1) );
  AND2X2 AND2X2_1046 ( .A(AES_CORE_DATAPATH__abc_16259_n4494_1), .B(AES_CORE_DATAPATH__abc_16259_n4475_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n4495_1) );
  AND2X2 AND2X2_1047 ( .A(AES_CORE_DATAPATH__abc_16259_n4474_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__1_), .Y(AES_CORE_DATAPATH__abc_16259_n4496_1) );
  AND2X2 AND2X2_1048 ( .A(AES_CORE_DATAPATH__abc_16259_n4468_1_bF_buf1), .B(AES_CORE_DATAPATH_key_host_0__2_), .Y(AES_CORE_DATAPATH__abc_16259_n4499_1) );
  AND2X2 AND2X2_1049 ( .A(key_en_0_bF_buf1), .B(\bus_in[2] ), .Y(AES_CORE_DATAPATH__abc_16259_n4500_1) );
  AND2X2 AND2X2_105 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk_bF_buf3), .B(AES_CORE_CONTROL_UNIT_col_en_2_), .Y(AES_CORE_DATAPATH__abc_16259_n2472) );
  AND2X2 AND2X2_1050 ( .A(AES_CORE_DATAPATH__abc_16259_n4498_1), .B(AES_CORE_DATAPATH__abc_16259_n4502_1), .Y(AES_CORE_DATAPATH__abc_16259_n4503_1) );
  AND2X2 AND2X2_1051 ( .A(AES_CORE_DATAPATH__abc_16259_n4503_1), .B(AES_CORE_DATAPATH__abc_16259_n4475_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n4504_1) );
  AND2X2 AND2X2_1052 ( .A(AES_CORE_DATAPATH__abc_16259_n4474_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__2_), .Y(AES_CORE_DATAPATH__abc_16259_n4505_1) );
  AND2X2 AND2X2_1053 ( .A(AES_CORE_DATAPATH__abc_16259_n4468_1_bF_buf0), .B(AES_CORE_DATAPATH_key_host_0__3_), .Y(AES_CORE_DATAPATH__abc_16259_n4508) );
  AND2X2 AND2X2_1054 ( .A(key_en_0_bF_buf0), .B(\bus_in[3] ), .Y(AES_CORE_DATAPATH__abc_16259_n4509) );
  AND2X2 AND2X2_1055 ( .A(AES_CORE_DATAPATH__abc_16259_n4507), .B(AES_CORE_DATAPATH__abc_16259_n4511), .Y(AES_CORE_DATAPATH__abc_16259_n4512) );
  AND2X2 AND2X2_1056 ( .A(AES_CORE_DATAPATH__abc_16259_n4512), .B(AES_CORE_DATAPATH__abc_16259_n4475_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n4513_1) );
  AND2X2 AND2X2_1057 ( .A(AES_CORE_DATAPATH__abc_16259_n4474_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__3_), .Y(AES_CORE_DATAPATH__abc_16259_n4514) );
  AND2X2 AND2X2_1058 ( .A(AES_CORE_DATAPATH__abc_16259_n4468_1_bF_buf4), .B(AES_CORE_DATAPATH_key_host_0__4_), .Y(AES_CORE_DATAPATH__abc_16259_n4517) );
  AND2X2 AND2X2_1059 ( .A(key_en_0_bF_buf4), .B(\bus_in[4] ), .Y(AES_CORE_DATAPATH__abc_16259_n4518) );
  AND2X2 AND2X2_106 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf6), .B(AES_CORE_DATAPATH_iv_1__0_), .Y(AES_CORE_DATAPATH__abc_16259_n2476) );
  AND2X2 AND2X2_1060 ( .A(AES_CORE_DATAPATH__abc_16259_n4516_1), .B(AES_CORE_DATAPATH__abc_16259_n4520), .Y(AES_CORE_DATAPATH__abc_16259_n4521) );
  AND2X2 AND2X2_1061 ( .A(AES_CORE_DATAPATH__abc_16259_n4522_1), .B(AES_CORE_DATAPATH__abc_16259_n4523), .Y(AES_CORE_DATAPATH__0key_0__31_0__4_) );
  AND2X2 AND2X2_1062 ( .A(AES_CORE_DATAPATH__abc_16259_n4468_1_bF_buf3), .B(AES_CORE_DATAPATH_key_host_0__5_), .Y(AES_CORE_DATAPATH__abc_16259_n4526) );
  AND2X2 AND2X2_1063 ( .A(key_en_0_bF_buf3), .B(\bus_in[5] ), .Y(AES_CORE_DATAPATH__abc_16259_n4527) );
  AND2X2 AND2X2_1064 ( .A(AES_CORE_DATAPATH__abc_16259_n4525_1), .B(AES_CORE_DATAPATH__abc_16259_n4529), .Y(AES_CORE_DATAPATH__abc_16259_n4530) );
  AND2X2 AND2X2_1065 ( .A(AES_CORE_DATAPATH__abc_16259_n4531_1), .B(AES_CORE_DATAPATH__abc_16259_n4532), .Y(AES_CORE_DATAPATH__0key_0__31_0__5_) );
  AND2X2 AND2X2_1066 ( .A(AES_CORE_DATAPATH__abc_16259_n4468_1_bF_buf2), .B(AES_CORE_DATAPATH_key_host_0__6_), .Y(AES_CORE_DATAPATH__abc_16259_n4535) );
  AND2X2 AND2X2_1067 ( .A(key_en_0_bF_buf2), .B(\bus_in[6] ), .Y(AES_CORE_DATAPATH__abc_16259_n4536) );
  AND2X2 AND2X2_1068 ( .A(AES_CORE_DATAPATH__abc_16259_n4534_1), .B(AES_CORE_DATAPATH__abc_16259_n4538), .Y(AES_CORE_DATAPATH__abc_16259_n4539) );
  AND2X2 AND2X2_1069 ( .A(AES_CORE_DATAPATH__abc_16259_n4539), .B(AES_CORE_DATAPATH__abc_16259_n4475_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n4540_1) );
  AND2X2 AND2X2_107 ( .A(AES_CORE_DATAPATH__abc_16259_n2457_1), .B(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_3_), .Y(AES_CORE_DATAPATH__abc_16259_n2479_1) );
  AND2X2 AND2X2_1070 ( .A(AES_CORE_DATAPATH__abc_16259_n4474_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__6_), .Y(AES_CORE_DATAPATH__abc_16259_n4541) );
  AND2X2 AND2X2_1071 ( .A(AES_CORE_DATAPATH__abc_16259_n4468_1_bF_buf1), .B(AES_CORE_DATAPATH_key_host_0__7_), .Y(AES_CORE_DATAPATH__abc_16259_n4544) );
  AND2X2 AND2X2_1072 ( .A(key_en_0_bF_buf1), .B(\bus_in[7] ), .Y(AES_CORE_DATAPATH__abc_16259_n4545) );
  AND2X2 AND2X2_1073 ( .A(AES_CORE_DATAPATH__abc_16259_n4543_1), .B(AES_CORE_DATAPATH__abc_16259_n4547), .Y(AES_CORE_DATAPATH__abc_16259_n4548) );
  AND2X2 AND2X2_1074 ( .A(AES_CORE_DATAPATH__abc_16259_n4548), .B(AES_CORE_DATAPATH__abc_16259_n4475_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n4549_1) );
  AND2X2 AND2X2_1075 ( .A(AES_CORE_DATAPATH__abc_16259_n4474_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__7_), .Y(AES_CORE_DATAPATH__abc_16259_n4550) );
  AND2X2 AND2X2_1076 ( .A(AES_CORE_DATAPATH__abc_16259_n4468_1_bF_buf0), .B(AES_CORE_DATAPATH_key_host_0__8_), .Y(AES_CORE_DATAPATH__abc_16259_n4553) );
  AND2X2 AND2X2_1077 ( .A(key_en_0_bF_buf0), .B(\bus_in[8] ), .Y(AES_CORE_DATAPATH__abc_16259_n4554) );
  AND2X2 AND2X2_1078 ( .A(AES_CORE_DATAPATH__abc_16259_n4552_1), .B(AES_CORE_DATAPATH__abc_16259_n4556), .Y(AES_CORE_DATAPATH__abc_16259_n4557) );
  AND2X2 AND2X2_1079 ( .A(AES_CORE_DATAPATH__abc_16259_n4557), .B(AES_CORE_DATAPATH__abc_16259_n4475_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n4558_1) );
  AND2X2 AND2X2_108 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk_bF_buf2), .B(AES_CORE_CONTROL_UNIT_col_en_3_), .Y(AES_CORE_DATAPATH__abc_16259_n2480) );
  AND2X2 AND2X2_1080 ( .A(AES_CORE_DATAPATH__abc_16259_n4474_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__8_), .Y(AES_CORE_DATAPATH__abc_16259_n4559) );
  AND2X2 AND2X2_1081 ( .A(AES_CORE_DATAPATH__abc_16259_n4468_1_bF_buf4), .B(AES_CORE_DATAPATH_key_host_0__9_), .Y(AES_CORE_DATAPATH__abc_16259_n4562) );
  AND2X2 AND2X2_1082 ( .A(key_en_0_bF_buf4), .B(\bus_in[9] ), .Y(AES_CORE_DATAPATH__abc_16259_n4563) );
  AND2X2 AND2X2_1083 ( .A(AES_CORE_DATAPATH__abc_16259_n4561_1), .B(AES_CORE_DATAPATH__abc_16259_n4565), .Y(AES_CORE_DATAPATH__abc_16259_n4566) );
  AND2X2 AND2X2_1084 ( .A(AES_CORE_DATAPATH__abc_16259_n4566), .B(AES_CORE_DATAPATH__abc_16259_n4475_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n4567_1) );
  AND2X2 AND2X2_1085 ( .A(AES_CORE_DATAPATH__abc_16259_n4474_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__9_), .Y(AES_CORE_DATAPATH__abc_16259_n4568) );
  AND2X2 AND2X2_1086 ( .A(AES_CORE_DATAPATH__abc_16259_n4468_1_bF_buf3), .B(AES_CORE_DATAPATH_key_host_0__10_), .Y(AES_CORE_DATAPATH__abc_16259_n4571) );
  AND2X2 AND2X2_1087 ( .A(key_en_0_bF_buf3), .B(\bus_in[10] ), .Y(AES_CORE_DATAPATH__abc_16259_n4572) );
  AND2X2 AND2X2_1088 ( .A(AES_CORE_DATAPATH__abc_16259_n4570_1), .B(AES_CORE_DATAPATH__abc_16259_n4574), .Y(AES_CORE_DATAPATH__abc_16259_n4575) );
  AND2X2 AND2X2_1089 ( .A(AES_CORE_DATAPATH__abc_16259_n4576_1), .B(AES_CORE_DATAPATH__abc_16259_n4577), .Y(AES_CORE_DATAPATH__0key_0__31_0__10_) );
  AND2X2 AND2X2_109 ( .A(AES_CORE_DATAPATH__abc_16259_n2486), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n2487_1) );
  AND2X2 AND2X2_1090 ( .A(AES_CORE_DATAPATH__abc_16259_n4468_1_bF_buf2), .B(AES_CORE_DATAPATH_key_host_0__11_), .Y(AES_CORE_DATAPATH__abc_16259_n4580) );
  AND2X2 AND2X2_1091 ( .A(key_en_0_bF_buf2), .B(\bus_in[11] ), .Y(AES_CORE_DATAPATH__abc_16259_n4581) );
  AND2X2 AND2X2_1092 ( .A(AES_CORE_DATAPATH__abc_16259_n4579_1), .B(AES_CORE_DATAPATH__abc_16259_n4583), .Y(AES_CORE_DATAPATH__abc_16259_n4584) );
  AND2X2 AND2X2_1093 ( .A(AES_CORE_DATAPATH__abc_16259_n4584), .B(AES_CORE_DATAPATH__abc_16259_n4475_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n4585_1) );
  AND2X2 AND2X2_1094 ( .A(AES_CORE_DATAPATH__abc_16259_n4474_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__11_), .Y(AES_CORE_DATAPATH__abc_16259_n4586) );
  AND2X2 AND2X2_1095 ( .A(AES_CORE_DATAPATH__abc_16259_n4468_1_bF_buf1), .B(AES_CORE_DATAPATH_key_host_0__12_), .Y(AES_CORE_DATAPATH__abc_16259_n4589) );
  AND2X2 AND2X2_1096 ( .A(key_en_0_bF_buf1), .B(\bus_in[12] ), .Y(AES_CORE_DATAPATH__abc_16259_n4590) );
  AND2X2 AND2X2_1097 ( .A(AES_CORE_DATAPATH__abc_16259_n4588_1), .B(AES_CORE_DATAPATH__abc_16259_n4592), .Y(AES_CORE_DATAPATH__abc_16259_n4593) );
  AND2X2 AND2X2_1098 ( .A(AES_CORE_DATAPATH__abc_16259_n4593), .B(AES_CORE_DATAPATH__abc_16259_n4475_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n4594_1) );
  AND2X2 AND2X2_1099 ( .A(AES_CORE_DATAPATH__abc_16259_n4474_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__12_), .Y(AES_CORE_DATAPATH__abc_16259_n4595) );
  AND2X2 AND2X2_11 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n82_1), .B(AES_CORE_CONTROL_UNIT__abc_15841_n81_1), .Y(AES_CORE_CONTROL_UNIT_last_round) );
  AND2X2 AND2X2_110 ( .A(AES_CORE_DATAPATH__abc_16259_n2478), .B(AES_CORE_DATAPATH__abc_16259_n2487_1), .Y(AES_CORE_DATAPATH__abc_16259_n2488) );
  AND2X2 AND2X2_1100 ( .A(AES_CORE_DATAPATH__abc_16259_n4468_1_bF_buf0), .B(AES_CORE_DATAPATH_key_host_0__13_), .Y(AES_CORE_DATAPATH__abc_16259_n4598) );
  AND2X2 AND2X2_1101 ( .A(key_en_0_bF_buf0), .B(\bus_in[13] ), .Y(AES_CORE_DATAPATH__abc_16259_n4599) );
  AND2X2 AND2X2_1102 ( .A(AES_CORE_DATAPATH__abc_16259_n4597_1), .B(AES_CORE_DATAPATH__abc_16259_n4601), .Y(AES_CORE_DATAPATH__abc_16259_n4602) );
  AND2X2 AND2X2_1103 ( .A(AES_CORE_DATAPATH__abc_16259_n4603_1), .B(AES_CORE_DATAPATH__abc_16259_n4604_1), .Y(AES_CORE_DATAPATH__0key_0__31_0__13_) );
  AND2X2 AND2X2_1104 ( .A(AES_CORE_DATAPATH__abc_16259_n4468_1_bF_buf4), .B(AES_CORE_DATAPATH_key_host_0__14_), .Y(AES_CORE_DATAPATH__abc_16259_n4607_1) );
  AND2X2 AND2X2_1105 ( .A(key_en_0_bF_buf4), .B(\bus_in[14] ), .Y(AES_CORE_DATAPATH__abc_16259_n4608) );
  AND2X2 AND2X2_1106 ( .A(AES_CORE_DATAPATH__abc_16259_n4606), .B(AES_CORE_DATAPATH__abc_16259_n4610), .Y(AES_CORE_DATAPATH__abc_16259_n4611_1) );
  AND2X2 AND2X2_1107 ( .A(AES_CORE_DATAPATH__abc_16259_n4612), .B(AES_CORE_DATAPATH__abc_16259_n4613), .Y(AES_CORE_DATAPATH__0key_0__31_0__14_) );
  AND2X2 AND2X2_1108 ( .A(AES_CORE_DATAPATH__abc_16259_n4468_1_bF_buf3), .B(AES_CORE_DATAPATH_key_host_0__15_), .Y(AES_CORE_DATAPATH__abc_16259_n4616_1) );
  AND2X2 AND2X2_1109 ( .A(key_en_0_bF_buf3), .B(\bus_in[15] ), .Y(AES_CORE_DATAPATH__abc_16259_n4617) );
  AND2X2 AND2X2_111 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf6), .B(AES_CORE_DATAPATH_iv_3__0_), .Y(AES_CORE_DATAPATH__abc_16259_n2489_1) );
  AND2X2 AND2X2_1110 ( .A(AES_CORE_DATAPATH__abc_16259_n4615), .B(AES_CORE_DATAPATH__abc_16259_n4619), .Y(AES_CORE_DATAPATH__abc_16259_n4620) );
  AND2X2 AND2X2_1111 ( .A(AES_CORE_DATAPATH__abc_16259_n4620), .B(AES_CORE_DATAPATH__abc_16259_n4475_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n4621) );
  AND2X2 AND2X2_1112 ( .A(AES_CORE_DATAPATH__abc_16259_n4474_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__15_), .Y(AES_CORE_DATAPATH__abc_16259_n4622_1) );
  AND2X2 AND2X2_1113 ( .A(AES_CORE_DATAPATH__abc_16259_n4468_1_bF_buf2), .B(AES_CORE_DATAPATH_key_host_0__16_), .Y(AES_CORE_DATAPATH__abc_16259_n4625) );
  AND2X2 AND2X2_1114 ( .A(key_en_0_bF_buf2), .B(\bus_in[16] ), .Y(AES_CORE_DATAPATH__abc_16259_n4626) );
  AND2X2 AND2X2_1115 ( .A(AES_CORE_DATAPATH__abc_16259_n4624), .B(AES_CORE_DATAPATH__abc_16259_n4628_1), .Y(AES_CORE_DATAPATH__abc_16259_n4629) );
  AND2X2 AND2X2_1116 ( .A(AES_CORE_DATAPATH__abc_16259_n4629), .B(AES_CORE_DATAPATH__abc_16259_n4475_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n4630) );
  AND2X2 AND2X2_1117 ( .A(AES_CORE_DATAPATH__abc_16259_n4474_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__16_), .Y(AES_CORE_DATAPATH__abc_16259_n4631) );
  AND2X2 AND2X2_1118 ( .A(AES_CORE_DATAPATH__abc_16259_n4468_1_bF_buf1), .B(AES_CORE_DATAPATH_key_host_0__17_), .Y(AES_CORE_DATAPATH__abc_16259_n4634) );
  AND2X2 AND2X2_1119 ( .A(key_en_0_bF_buf1), .B(\bus_in[17] ), .Y(AES_CORE_DATAPATH__abc_16259_n4635_1) );
  AND2X2 AND2X2_112 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf6), .B(AES_CORE_DATAPATH_iv_0__1_), .Y(AES_CORE_DATAPATH__abc_16259_n2491_1) );
  AND2X2 AND2X2_1120 ( .A(AES_CORE_DATAPATH__abc_16259_n4633), .B(AES_CORE_DATAPATH__abc_16259_n4637), .Y(AES_CORE_DATAPATH__abc_16259_n4638) );
  AND2X2 AND2X2_1121 ( .A(AES_CORE_DATAPATH__abc_16259_n4638), .B(AES_CORE_DATAPATH__abc_16259_n4475_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n4639) );
  AND2X2 AND2X2_1122 ( .A(AES_CORE_DATAPATH__abc_16259_n4474_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__17_), .Y(AES_CORE_DATAPATH__abc_16259_n4640) );
  AND2X2 AND2X2_1123 ( .A(AES_CORE_DATAPATH__abc_16259_n4468_1_bF_buf0), .B(AES_CORE_DATAPATH_key_host_0__18_), .Y(AES_CORE_DATAPATH__abc_16259_n4643) );
  AND2X2 AND2X2_1124 ( .A(key_en_0_bF_buf0), .B(\bus_in[18] ), .Y(AES_CORE_DATAPATH__abc_16259_n4644) );
  AND2X2 AND2X2_1125 ( .A(AES_CORE_DATAPATH__abc_16259_n4642), .B(AES_CORE_DATAPATH__abc_16259_n4646), .Y(AES_CORE_DATAPATH__abc_16259_n4647) );
  AND2X2 AND2X2_1126 ( .A(AES_CORE_DATAPATH__abc_16259_n4648_1), .B(AES_CORE_DATAPATH__abc_16259_n4649), .Y(AES_CORE_DATAPATH__0key_0__31_0__18_) );
  AND2X2 AND2X2_1127 ( .A(AES_CORE_DATAPATH__abc_16259_n4468_1_bF_buf4), .B(AES_CORE_DATAPATH_key_host_0__19_), .Y(AES_CORE_DATAPATH__abc_16259_n4652) );
  AND2X2 AND2X2_1128 ( .A(key_en_0_bF_buf4), .B(\bus_in[19] ), .Y(AES_CORE_DATAPATH__abc_16259_n4653) );
  AND2X2 AND2X2_1129 ( .A(AES_CORE_DATAPATH__abc_16259_n4651), .B(AES_CORE_DATAPATH__abc_16259_n4655), .Y(AES_CORE_DATAPATH__abc_16259_n4656) );
  AND2X2 AND2X2_113 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf5), .B(AES_CORE_DATAPATH_iv_1__1_), .Y(AES_CORE_DATAPATH__abc_16259_n2492_1) );
  AND2X2 AND2X2_1130 ( .A(AES_CORE_DATAPATH__abc_16259_n4656), .B(AES_CORE_DATAPATH__abc_16259_n4475_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n4657) );
  AND2X2 AND2X2_1131 ( .A(AES_CORE_DATAPATH__abc_16259_n4474_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__19_), .Y(AES_CORE_DATAPATH__abc_16259_n4658) );
  AND2X2 AND2X2_1132 ( .A(AES_CORE_DATAPATH__abc_16259_n4468_1_bF_buf3), .B(AES_CORE_DATAPATH_key_host_0__20_), .Y(AES_CORE_DATAPATH__abc_16259_n4661) );
  AND2X2 AND2X2_1133 ( .A(key_en_0_bF_buf3), .B(\bus_in[20] ), .Y(AES_CORE_DATAPATH__abc_16259_n4662_1) );
  AND2X2 AND2X2_1134 ( .A(AES_CORE_DATAPATH__abc_16259_n4660), .B(AES_CORE_DATAPATH__abc_16259_n4664), .Y(AES_CORE_DATAPATH__abc_16259_n4665) );
  AND2X2 AND2X2_1135 ( .A(AES_CORE_DATAPATH__abc_16259_n4665), .B(AES_CORE_DATAPATH__abc_16259_n4475_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n4666) );
  AND2X2 AND2X2_1136 ( .A(AES_CORE_DATAPATH__abc_16259_n4474_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__20_), .Y(AES_CORE_DATAPATH__abc_16259_n4667) );
  AND2X2 AND2X2_1137 ( .A(AES_CORE_DATAPATH__abc_16259_n4468_1_bF_buf2), .B(AES_CORE_DATAPATH_key_host_0__21_), .Y(AES_CORE_DATAPATH__abc_16259_n4670) );
  AND2X2 AND2X2_1138 ( .A(key_en_0_bF_buf2), .B(\bus_in[21] ), .Y(AES_CORE_DATAPATH__abc_16259_n4671) );
  AND2X2 AND2X2_1139 ( .A(AES_CORE_DATAPATH__abc_16259_n4669), .B(AES_CORE_DATAPATH__abc_16259_n4673), .Y(AES_CORE_DATAPATH__abc_16259_n4674) );
  AND2X2 AND2X2_114 ( .A(AES_CORE_DATAPATH__abc_16259_n2495), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n2496) );
  AND2X2 AND2X2_1140 ( .A(AES_CORE_DATAPATH__abc_16259_n4675_1), .B(AES_CORE_DATAPATH__abc_16259_n4676), .Y(AES_CORE_DATAPATH__0key_0__31_0__21_) );
  AND2X2 AND2X2_1141 ( .A(AES_CORE_DATAPATH__abc_16259_n4468_1_bF_buf1), .B(AES_CORE_DATAPATH_key_host_0__22_), .Y(AES_CORE_DATAPATH__abc_16259_n4679) );
  AND2X2 AND2X2_1142 ( .A(key_en_0_bF_buf1), .B(\bus_in[22] ), .Y(AES_CORE_DATAPATH__abc_16259_n4680) );
  AND2X2 AND2X2_1143 ( .A(AES_CORE_DATAPATH__abc_16259_n4678), .B(AES_CORE_DATAPATH__abc_16259_n4682), .Y(AES_CORE_DATAPATH__abc_16259_n4683) );
  AND2X2 AND2X2_1144 ( .A(AES_CORE_DATAPATH__abc_16259_n4684), .B(AES_CORE_DATAPATH__abc_16259_n4685), .Y(AES_CORE_DATAPATH__0key_0__31_0__22_) );
  AND2X2 AND2X2_1145 ( .A(AES_CORE_DATAPATH__abc_16259_n4468_1_bF_buf0), .B(AES_CORE_DATAPATH_key_host_0__23_), .Y(AES_CORE_DATAPATH__abc_16259_n4688) );
  AND2X2 AND2X2_1146 ( .A(key_en_0_bF_buf0), .B(\bus_in[23] ), .Y(AES_CORE_DATAPATH__abc_16259_n4689_1) );
  AND2X2 AND2X2_1147 ( .A(AES_CORE_DATAPATH__abc_16259_n4687), .B(AES_CORE_DATAPATH__abc_16259_n4691), .Y(AES_CORE_DATAPATH__abc_16259_n4692) );
  AND2X2 AND2X2_1148 ( .A(AES_CORE_DATAPATH__abc_16259_n4692), .B(AES_CORE_DATAPATH__abc_16259_n4475_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n4693) );
  AND2X2 AND2X2_1149 ( .A(AES_CORE_DATAPATH__abc_16259_n4474_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__23_), .Y(AES_CORE_DATAPATH__abc_16259_n4694) );
  AND2X2 AND2X2_115 ( .A(AES_CORE_DATAPATH__abc_16259_n2494_1), .B(AES_CORE_DATAPATH__abc_16259_n2496), .Y(AES_CORE_DATAPATH__abc_16259_n2497_1) );
  AND2X2 AND2X2_1150 ( .A(AES_CORE_DATAPATH__abc_16259_n4468_1_bF_buf4), .B(AES_CORE_DATAPATH_key_host_0__24_), .Y(AES_CORE_DATAPATH__abc_16259_n4697) );
  AND2X2 AND2X2_1151 ( .A(key_en_0_bF_buf4), .B(\bus_in[24] ), .Y(AES_CORE_DATAPATH__abc_16259_n4698) );
  AND2X2 AND2X2_1152 ( .A(AES_CORE_DATAPATH__abc_16259_n4696), .B(AES_CORE_DATAPATH__abc_16259_n4700), .Y(AES_CORE_DATAPATH__abc_16259_n4701) );
  AND2X2 AND2X2_1153 ( .A(AES_CORE_DATAPATH__abc_16259_n4701), .B(AES_CORE_DATAPATH__abc_16259_n4475_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n4702_1) );
  AND2X2 AND2X2_1154 ( .A(AES_CORE_DATAPATH__abc_16259_n4474_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__24_), .Y(AES_CORE_DATAPATH__abc_16259_n4703) );
  AND2X2 AND2X2_1155 ( .A(AES_CORE_DATAPATH__abc_16259_n4468_1_bF_buf3), .B(AES_CORE_DATAPATH_key_host_0__25_), .Y(AES_CORE_DATAPATH__abc_16259_n4706) );
  AND2X2 AND2X2_1156 ( .A(key_en_0_bF_buf3), .B(\bus_in[25] ), .Y(AES_CORE_DATAPATH__abc_16259_n4707) );
  AND2X2 AND2X2_1157 ( .A(AES_CORE_DATAPATH__abc_16259_n4705), .B(AES_CORE_DATAPATH__abc_16259_n4709), .Y(AES_CORE_DATAPATH__abc_16259_n4710) );
  AND2X2 AND2X2_1158 ( .A(AES_CORE_DATAPATH__abc_16259_n4710), .B(AES_CORE_DATAPATH__abc_16259_n4475_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n4711) );
  AND2X2 AND2X2_1159 ( .A(AES_CORE_DATAPATH__abc_16259_n4474_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__25_), .Y(AES_CORE_DATAPATH__abc_16259_n4712) );
  AND2X2 AND2X2_116 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf5), .B(AES_CORE_DATAPATH_iv_3__1_), .Y(AES_CORE_DATAPATH__abc_16259_n2498) );
  AND2X2 AND2X2_1160 ( .A(AES_CORE_DATAPATH__abc_16259_n4468_1_bF_buf2), .B(AES_CORE_DATAPATH_key_host_0__26_), .Y(AES_CORE_DATAPATH__abc_16259_n4715) );
  AND2X2 AND2X2_1161 ( .A(key_en_0_bF_buf2), .B(\bus_in[26] ), .Y(AES_CORE_DATAPATH__abc_16259_n4716) );
  AND2X2 AND2X2_1162 ( .A(AES_CORE_DATAPATH__abc_16259_n4714), .B(AES_CORE_DATAPATH__abc_16259_n4718), .Y(AES_CORE_DATAPATH__abc_16259_n4719) );
  AND2X2 AND2X2_1163 ( .A(AES_CORE_DATAPATH__abc_16259_n4719), .B(AES_CORE_DATAPATH__abc_16259_n4475_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n4720) );
  AND2X2 AND2X2_1164 ( .A(AES_CORE_DATAPATH__abc_16259_n4474_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__26_), .Y(AES_CORE_DATAPATH__abc_16259_n4721) );
  AND2X2 AND2X2_1165 ( .A(AES_CORE_DATAPATH__abc_16259_n4468_1_bF_buf1), .B(AES_CORE_DATAPATH_key_host_0__27_), .Y(AES_CORE_DATAPATH__abc_16259_n4724) );
  AND2X2 AND2X2_1166 ( .A(key_en_0_bF_buf1), .B(\bus_in[27] ), .Y(AES_CORE_DATAPATH__abc_16259_n4725) );
  AND2X2 AND2X2_1167 ( .A(AES_CORE_DATAPATH__abc_16259_n4723_1), .B(AES_CORE_DATAPATH__abc_16259_n4727), .Y(AES_CORE_DATAPATH__abc_16259_n4728) );
  AND2X2 AND2X2_1168 ( .A(AES_CORE_DATAPATH__abc_16259_n4728), .B(AES_CORE_DATAPATH__abc_16259_n4475_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n4729) );
  AND2X2 AND2X2_1169 ( .A(AES_CORE_DATAPATH__abc_16259_n4474_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__27_), .Y(AES_CORE_DATAPATH__abc_16259_n4730_1) );
  AND2X2 AND2X2_117 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf5), .B(AES_CORE_DATAPATH_iv_0__2_), .Y(AES_CORE_DATAPATH__abc_16259_n2500) );
  AND2X2 AND2X2_1170 ( .A(AES_CORE_DATAPATH__abc_16259_n4468_1_bF_buf0), .B(AES_CORE_DATAPATH_key_host_0__28_), .Y(AES_CORE_DATAPATH__abc_16259_n4733) );
  AND2X2 AND2X2_1171 ( .A(key_en_0_bF_buf0), .B(\bus_in[28] ), .Y(AES_CORE_DATAPATH__abc_16259_n4734) );
  AND2X2 AND2X2_1172 ( .A(AES_CORE_DATAPATH__abc_16259_n4732), .B(AES_CORE_DATAPATH__abc_16259_n4736_1), .Y(AES_CORE_DATAPATH__abc_16259_n4737) );
  AND2X2 AND2X2_1173 ( .A(AES_CORE_DATAPATH__abc_16259_n4738), .B(AES_CORE_DATAPATH__abc_16259_n4739), .Y(AES_CORE_DATAPATH__0key_0__31_0__28_) );
  AND2X2 AND2X2_1174 ( .A(AES_CORE_DATAPATH__abc_16259_n4468_1_bF_buf4), .B(AES_CORE_DATAPATH_key_host_0__29_), .Y(AES_CORE_DATAPATH__abc_16259_n4742) );
  AND2X2 AND2X2_1175 ( .A(key_en_0_bF_buf4), .B(\bus_in[29] ), .Y(AES_CORE_DATAPATH__abc_16259_n4743) );
  AND2X2 AND2X2_1176 ( .A(AES_CORE_DATAPATH__abc_16259_n4741), .B(AES_CORE_DATAPATH__abc_16259_n4745), .Y(AES_CORE_DATAPATH__abc_16259_n4746) );
  AND2X2 AND2X2_1177 ( .A(AES_CORE_DATAPATH__abc_16259_n4746), .B(AES_CORE_DATAPATH__abc_16259_n4475_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n4747) );
  AND2X2 AND2X2_1178 ( .A(AES_CORE_DATAPATH__abc_16259_n4474_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__29_), .Y(AES_CORE_DATAPATH__abc_16259_n4748) );
  AND2X2 AND2X2_1179 ( .A(AES_CORE_DATAPATH__abc_16259_n4468_1_bF_buf3), .B(AES_CORE_DATAPATH_key_host_0__30_), .Y(AES_CORE_DATAPATH__abc_16259_n4751) );
  AND2X2 AND2X2_118 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf4), .B(AES_CORE_DATAPATH_iv_1__2_), .Y(AES_CORE_DATAPATH__abc_16259_n2501_1) );
  AND2X2 AND2X2_1180 ( .A(key_en_0_bF_buf3), .B(\bus_in[30] ), .Y(AES_CORE_DATAPATH__abc_16259_n4752) );
  AND2X2 AND2X2_1181 ( .A(AES_CORE_DATAPATH__abc_16259_n4750_1), .B(AES_CORE_DATAPATH__abc_16259_n4754), .Y(AES_CORE_DATAPATH__abc_16259_n4755) );
  AND2X2 AND2X2_1182 ( .A(AES_CORE_DATAPATH__abc_16259_n4755), .B(AES_CORE_DATAPATH__abc_16259_n4475_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n4756) );
  AND2X2 AND2X2_1183 ( .A(AES_CORE_DATAPATH__abc_16259_n4474_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__30_), .Y(AES_CORE_DATAPATH__abc_16259_n4757_1) );
  AND2X2 AND2X2_1184 ( .A(AES_CORE_DATAPATH__abc_16259_n4468_1_bF_buf2), .B(AES_CORE_DATAPATH_key_host_0__31_), .Y(AES_CORE_DATAPATH__abc_16259_n4760) );
  AND2X2 AND2X2_1185 ( .A(key_en_0_bF_buf2), .B(\bus_in[31] ), .Y(AES_CORE_DATAPATH__abc_16259_n4761) );
  AND2X2 AND2X2_1186 ( .A(AES_CORE_DATAPATH__abc_16259_n4759), .B(AES_CORE_DATAPATH__abc_16259_n4763_1), .Y(AES_CORE_DATAPATH__abc_16259_n4764) );
  AND2X2 AND2X2_1187 ( .A(AES_CORE_DATAPATH__abc_16259_n4765), .B(AES_CORE_DATAPATH__abc_16259_n4766), .Y(AES_CORE_DATAPATH__0key_0__31_0__31_) );
  AND2X2 AND2X2_1188 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__0_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf10), .Y(AES_CORE_DATAPATH__abc_16259_n4768) );
  AND2X2 AND2X2_1189 ( .A(AES_CORE_DATAPATH__abc_16259_n4483_1), .B(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf10), .Y(AES_CORE_DATAPATH__abc_16259_n4770) );
  AND2X2 AND2X2_119 ( .A(AES_CORE_DATAPATH__abc_16259_n2504_1), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n2505) );
  AND2X2 AND2X2_1190 ( .A(AES_CORE_DATAPATH__abc_16259_n4772_1), .B(AES_CORE_DATAPATH__abc_16259_n4773), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__1_) );
  AND2X2 AND2X2_1191 ( .A(AES_CORE_DATAPATH__abc_16259_n4775), .B(AES_CORE_DATAPATH__abc_16259_n4776), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__2_) );
  AND2X2 AND2X2_1192 ( .A(AES_CORE_DATAPATH__abc_16259_n4778_1), .B(AES_CORE_DATAPATH__abc_16259_n4779), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__3_) );
  AND2X2 AND2X2_1193 ( .A(AES_CORE_DATAPATH__abc_16259_n4781), .B(AES_CORE_DATAPATH__abc_16259_n4782), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__4_) );
  AND2X2 AND2X2_1194 ( .A(AES_CORE_DATAPATH__abc_16259_n4784), .B(AES_CORE_DATAPATH__abc_16259_n4785_1), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__5_) );
  AND2X2 AND2X2_1195 ( .A(AES_CORE_DATAPATH__abc_16259_n4787), .B(AES_CORE_DATAPATH__abc_16259_n4788), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__6_) );
  AND2X2 AND2X2_1196 ( .A(AES_CORE_DATAPATH__abc_16259_n4790), .B(AES_CORE_DATAPATH__abc_16259_n4791_1), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__7_) );
  AND2X2 AND2X2_1197 ( .A(AES_CORE_DATAPATH__abc_16259_n4793), .B(AES_CORE_DATAPATH__abc_16259_n4794), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__8_) );
  AND2X2 AND2X2_1198 ( .A(AES_CORE_DATAPATH__abc_16259_n4796), .B(AES_CORE_DATAPATH__abc_16259_n4797), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__9_) );
  AND2X2 AND2X2_1199 ( .A(AES_CORE_DATAPATH__abc_16259_n4799_1), .B(AES_CORE_DATAPATH__abc_16259_n4800), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__10_) );
  AND2X2 AND2X2_12 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf14), .B(AES_CORE_CONTROL_UNIT__abc_15841_n84_1), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n85) );
  AND2X2 AND2X2_120 ( .A(AES_CORE_DATAPATH__abc_16259_n2503_1), .B(AES_CORE_DATAPATH__abc_16259_n2505), .Y(AES_CORE_DATAPATH__abc_16259_n2506_1) );
  AND2X2 AND2X2_1200 ( .A(AES_CORE_DATAPATH__abc_16259_n4802), .B(AES_CORE_DATAPATH__abc_16259_n4803), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__11_) );
  AND2X2 AND2X2_1201 ( .A(AES_CORE_DATAPATH__abc_16259_n4805_1), .B(AES_CORE_DATAPATH__abc_16259_n4806), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__12_) );
  AND2X2 AND2X2_1202 ( .A(AES_CORE_DATAPATH__abc_16259_n4808), .B(AES_CORE_DATAPATH__abc_16259_n4809), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__13_) );
  AND2X2 AND2X2_1203 ( .A(AES_CORE_DATAPATH__abc_16259_n4811), .B(AES_CORE_DATAPATH__abc_16259_n4812_1), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__14_) );
  AND2X2 AND2X2_1204 ( .A(AES_CORE_DATAPATH__abc_16259_n4814), .B(AES_CORE_DATAPATH__abc_16259_n4815), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__15_) );
  AND2X2 AND2X2_1205 ( .A(AES_CORE_DATAPATH__abc_16259_n4817), .B(AES_CORE_DATAPATH__abc_16259_n4818_1), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__16_) );
  AND2X2 AND2X2_1206 ( .A(AES_CORE_DATAPATH__abc_16259_n4820_1), .B(AES_CORE_DATAPATH__abc_16259_n4821_1), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__17_) );
  AND2X2 AND2X2_1207 ( .A(AES_CORE_DATAPATH__abc_16259_n4823_1), .B(AES_CORE_DATAPATH__abc_16259_n4824_1), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__18_) );
  AND2X2 AND2X2_1208 ( .A(AES_CORE_DATAPATH__abc_16259_n4826_1), .B(AES_CORE_DATAPATH__abc_16259_n4827_1), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__19_) );
  AND2X2 AND2X2_1209 ( .A(AES_CORE_DATAPATH__abc_16259_n4829_1), .B(AES_CORE_DATAPATH__abc_16259_n4830_1), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__20_) );
  AND2X2 AND2X2_121 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf4), .B(AES_CORE_DATAPATH_iv_3__2_), .Y(AES_CORE_DATAPATH__abc_16259_n2507) );
  AND2X2 AND2X2_1210 ( .A(AES_CORE_DATAPATH__abc_16259_n4832_1), .B(AES_CORE_DATAPATH__abc_16259_n4833_1), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__21_) );
  AND2X2 AND2X2_1211 ( .A(AES_CORE_DATAPATH__abc_16259_n4835_1), .B(AES_CORE_DATAPATH__abc_16259_n4836_1), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__22_) );
  AND2X2 AND2X2_1212 ( .A(AES_CORE_DATAPATH__abc_16259_n4838_1), .B(AES_CORE_DATAPATH__abc_16259_n4839_1), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__23_) );
  AND2X2 AND2X2_1213 ( .A(AES_CORE_DATAPATH__abc_16259_n4841_1), .B(AES_CORE_DATAPATH__abc_16259_n4842_1), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__24_) );
  AND2X2 AND2X2_1214 ( .A(AES_CORE_DATAPATH__abc_16259_n4844_1), .B(AES_CORE_DATAPATH__abc_16259_n4845_1), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__25_) );
  AND2X2 AND2X2_1215 ( .A(AES_CORE_DATAPATH__abc_16259_n4847_1), .B(AES_CORE_DATAPATH__abc_16259_n4848_1), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__26_) );
  AND2X2 AND2X2_1216 ( .A(AES_CORE_DATAPATH__abc_16259_n4850_1), .B(AES_CORE_DATAPATH__abc_16259_n4851_1), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__27_) );
  AND2X2 AND2X2_1217 ( .A(AES_CORE_DATAPATH__abc_16259_n4853_1), .B(AES_CORE_DATAPATH__abc_16259_n4854_1), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__28_) );
  AND2X2 AND2X2_1218 ( .A(AES_CORE_DATAPATH__abc_16259_n4856_1), .B(AES_CORE_DATAPATH__abc_16259_n4857_1), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__29_) );
  AND2X2 AND2X2_1219 ( .A(AES_CORE_DATAPATH__abc_16259_n4859_1), .B(AES_CORE_DATAPATH__abc_16259_n4860_1), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__30_) );
  AND2X2 AND2X2_122 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf4), .B(AES_CORE_DATAPATH_iv_0__3_), .Y(AES_CORE_DATAPATH__abc_16259_n2509_1) );
  AND2X2 AND2X2_1220 ( .A(AES_CORE_DATAPATH__abc_16259_n4863_1), .B(AES_CORE_DATAPATH__abc_16259_n4862_1), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__31_) );
  AND2X2 AND2X2_1221 ( .A(AES_CORE_CONTROL_UNIT_bypass_key_en), .B(AES_CORE_CONTROL_UNIT_key_en_1_), .Y(AES_CORE_DATAPATH__abc_16259_n4865_1) );
  AND2X2 AND2X2_1222 ( .A(AES_CORE_DATAPATH__abc_16259_n4469_1), .B(AES_CORE_DATAPATH__abc_16259_n4867_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n4868_1) );
  AND2X2 AND2X2_1223 ( .A(AES_CORE_DATAPATH__abc_16259_n2806_1), .B(AES_CORE_DATAPATH_key_en_pp1_1_), .Y(AES_CORE_DATAPATH__abc_16259_n4869_1) );
  AND2X2 AND2X2_1224 ( .A(AES_CORE_DATAPATH__abc_16259_n4870_1), .B(AES_CORE_DATAPATH__abc_16259_n4868_1), .Y(AES_CORE_DATAPATH__abc_16259_n4871_1) );
  AND2X2 AND2X2_1225 ( .A(AES_CORE_DATAPATH__abc_16259_n4871_1), .B(AES_CORE_DATAPATH__abc_16259_n4866_1), .Y(AES_CORE_DATAPATH__abc_16259_n4872_1) );
  AND2X2 AND2X2_1226 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf10), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_64_), .Y(AES_CORE_DATAPATH__abc_16259_n4874_1) );
  AND2X2 AND2X2_1227 ( .A(\bus_in[0] ), .B(key_en_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n4875_1) );
  AND2X2 AND2X2_1228 ( .A(AES_CORE_DATAPATH__abc_16259_n4867_1_bF_buf3), .B(AES_CORE_DATAPATH_key_host_1__0_), .Y(AES_CORE_DATAPATH__abc_16259_n4876_1) );
  AND2X2 AND2X2_1229 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n4877_1), .Y(AES_CORE_DATAPATH__abc_16259_n4878_1) );
  AND2X2 AND2X2_123 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf3), .B(AES_CORE_DATAPATH_iv_1__3_), .Y(AES_CORE_DATAPATH__abc_16259_n2510) );
  AND2X2 AND2X2_1230 ( .A(AES_CORE_DATAPATH__abc_16259_n4879_1), .B(AES_CORE_DATAPATH__abc_16259_n4873_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n4880_1) );
  AND2X2 AND2X2_1231 ( .A(AES_CORE_DATAPATH__abc_16259_n4872_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__0_), .Y(AES_CORE_DATAPATH__abc_16259_n4881_1) );
  AND2X2 AND2X2_1232 ( .A(AES_CORE_DATAPATH__abc_16259_n4867_1_bF_buf2), .B(AES_CORE_DATAPATH_key_host_1__1_), .Y(AES_CORE_DATAPATH__abc_16259_n4884) );
  AND2X2 AND2X2_1233 ( .A(\bus_in[1] ), .B(key_en_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n4885) );
  AND2X2 AND2X2_1234 ( .A(AES_CORE_DATAPATH__abc_16259_n4883_1), .B(AES_CORE_DATAPATH__abc_16259_n4887), .Y(AES_CORE_DATAPATH__abc_16259_n4888) );
  AND2X2 AND2X2_1235 ( .A(AES_CORE_DATAPATH__abc_16259_n4888), .B(AES_CORE_DATAPATH__abc_16259_n4873_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n4889_1) );
  AND2X2 AND2X2_1236 ( .A(AES_CORE_DATAPATH__abc_16259_n4872_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__1_), .Y(AES_CORE_DATAPATH__abc_16259_n4890) );
  AND2X2 AND2X2_1237 ( .A(AES_CORE_DATAPATH__abc_16259_n4867_1_bF_buf1), .B(AES_CORE_DATAPATH_key_host_1__2_), .Y(AES_CORE_DATAPATH__abc_16259_n4893) );
  AND2X2 AND2X2_1238 ( .A(\bus_in[2] ), .B(key_en_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n4894) );
  AND2X2 AND2X2_1239 ( .A(AES_CORE_DATAPATH__abc_16259_n4892_1), .B(AES_CORE_DATAPATH__abc_16259_n4896), .Y(AES_CORE_DATAPATH__abc_16259_n4897) );
  AND2X2 AND2X2_124 ( .A(AES_CORE_DATAPATH__abc_16259_n2513_1), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n2514_1) );
  AND2X2 AND2X2_1240 ( .A(AES_CORE_DATAPATH__abc_16259_n4898_1), .B(AES_CORE_DATAPATH__abc_16259_n4899), .Y(AES_CORE_DATAPATH__0key_1__31_0__2_) );
  AND2X2 AND2X2_1241 ( .A(AES_CORE_DATAPATH__abc_16259_n4867_1_bF_buf0), .B(AES_CORE_DATAPATH_key_host_1__3_), .Y(AES_CORE_DATAPATH__abc_16259_n4902) );
  AND2X2 AND2X2_1242 ( .A(\bus_in[3] ), .B(key_en_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n4903) );
  AND2X2 AND2X2_1243 ( .A(AES_CORE_DATAPATH__abc_16259_n4901_1), .B(AES_CORE_DATAPATH__abc_16259_n4905), .Y(AES_CORE_DATAPATH__abc_16259_n4906) );
  AND2X2 AND2X2_1244 ( .A(AES_CORE_DATAPATH__abc_16259_n4906), .B(AES_CORE_DATAPATH__abc_16259_n4873_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n4907_1) );
  AND2X2 AND2X2_1245 ( .A(AES_CORE_DATAPATH__abc_16259_n4872_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__3_), .Y(AES_CORE_DATAPATH__abc_16259_n4908) );
  AND2X2 AND2X2_1246 ( .A(AES_CORE_DATAPATH__abc_16259_n4867_1_bF_buf4), .B(AES_CORE_DATAPATH_key_host_1__4_), .Y(AES_CORE_DATAPATH__abc_16259_n4911) );
  AND2X2 AND2X2_1247 ( .A(\bus_in[4] ), .B(key_en_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n4912) );
  AND2X2 AND2X2_1248 ( .A(AES_CORE_DATAPATH__abc_16259_n4910_1), .B(AES_CORE_DATAPATH__abc_16259_n4914), .Y(AES_CORE_DATAPATH__abc_16259_n4915) );
  AND2X2 AND2X2_1249 ( .A(AES_CORE_DATAPATH__abc_16259_n4915), .B(AES_CORE_DATAPATH__abc_16259_n4873_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n4916_1) );
  AND2X2 AND2X2_125 ( .A(AES_CORE_DATAPATH__abc_16259_n2512), .B(AES_CORE_DATAPATH__abc_16259_n2514_1), .Y(AES_CORE_DATAPATH__abc_16259_n2515) );
  AND2X2 AND2X2_1250 ( .A(AES_CORE_DATAPATH__abc_16259_n4872_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__4_), .Y(AES_CORE_DATAPATH__abc_16259_n4917) );
  AND2X2 AND2X2_1251 ( .A(AES_CORE_DATAPATH__abc_16259_n4867_1_bF_buf3), .B(AES_CORE_DATAPATH_key_host_1__5_), .Y(AES_CORE_DATAPATH__abc_16259_n4920) );
  AND2X2 AND2X2_1252 ( .A(\bus_in[5] ), .B(key_en_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n4921) );
  AND2X2 AND2X2_1253 ( .A(AES_CORE_DATAPATH__abc_16259_n4919_1), .B(AES_CORE_DATAPATH__abc_16259_n4923), .Y(AES_CORE_DATAPATH__abc_16259_n4924) );
  AND2X2 AND2X2_1254 ( .A(AES_CORE_DATAPATH__abc_16259_n4925_1), .B(AES_CORE_DATAPATH__abc_16259_n4926), .Y(AES_CORE_DATAPATH__0key_1__31_0__5_) );
  AND2X2 AND2X2_1255 ( .A(AES_CORE_DATAPATH__abc_16259_n4867_1_bF_buf2), .B(AES_CORE_DATAPATH_key_host_1__6_), .Y(AES_CORE_DATAPATH__abc_16259_n4929) );
  AND2X2 AND2X2_1256 ( .A(\bus_in[6] ), .B(key_en_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n4930) );
  AND2X2 AND2X2_1257 ( .A(AES_CORE_DATAPATH__abc_16259_n4928_1), .B(AES_CORE_DATAPATH__abc_16259_n4932), .Y(AES_CORE_DATAPATH__abc_16259_n4933) );
  AND2X2 AND2X2_1258 ( .A(AES_CORE_DATAPATH__abc_16259_n4934_1), .B(AES_CORE_DATAPATH__abc_16259_n4935), .Y(AES_CORE_DATAPATH__0key_1__31_0__6_) );
  AND2X2 AND2X2_1259 ( .A(AES_CORE_DATAPATH__abc_16259_n4867_1_bF_buf1), .B(AES_CORE_DATAPATH_key_host_1__7_), .Y(AES_CORE_DATAPATH__abc_16259_n4938) );
  AND2X2 AND2X2_126 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf3), .B(AES_CORE_DATAPATH_iv_3__3_), .Y(AES_CORE_DATAPATH__abc_16259_n2516_1) );
  AND2X2 AND2X2_1260 ( .A(\bus_in[7] ), .B(key_en_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n4939) );
  AND2X2 AND2X2_1261 ( .A(AES_CORE_DATAPATH__abc_16259_n4937_1), .B(AES_CORE_DATAPATH__abc_16259_n4941), .Y(AES_CORE_DATAPATH__abc_16259_n4942) );
  AND2X2 AND2X2_1262 ( .A(AES_CORE_DATAPATH__abc_16259_n4942), .B(AES_CORE_DATAPATH__abc_16259_n4873_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n4943_1) );
  AND2X2 AND2X2_1263 ( .A(AES_CORE_DATAPATH__abc_16259_n4872_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__7_), .Y(AES_CORE_DATAPATH__abc_16259_n4944) );
  AND2X2 AND2X2_1264 ( .A(AES_CORE_DATAPATH__abc_16259_n4867_1_bF_buf0), .B(AES_CORE_DATAPATH_key_host_1__8_), .Y(AES_CORE_DATAPATH__abc_16259_n4947) );
  AND2X2 AND2X2_1265 ( .A(\bus_in[8] ), .B(key_en_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n4948) );
  AND2X2 AND2X2_1266 ( .A(AES_CORE_DATAPATH__abc_16259_n4946_1), .B(AES_CORE_DATAPATH__abc_16259_n4950), .Y(AES_CORE_DATAPATH__abc_16259_n4951) );
  AND2X2 AND2X2_1267 ( .A(AES_CORE_DATAPATH__abc_16259_n4951), .B(AES_CORE_DATAPATH__abc_16259_n4873_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n4952_1) );
  AND2X2 AND2X2_1268 ( .A(AES_CORE_DATAPATH__abc_16259_n4872_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__8_), .Y(AES_CORE_DATAPATH__abc_16259_n4953) );
  AND2X2 AND2X2_1269 ( .A(AES_CORE_DATAPATH__abc_16259_n4867_1_bF_buf4), .B(AES_CORE_DATAPATH_key_host_1__9_), .Y(AES_CORE_DATAPATH__abc_16259_n4956) );
  AND2X2 AND2X2_127 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf3), .B(AES_CORE_DATAPATH_iv_0__4_), .Y(AES_CORE_DATAPATH__abc_16259_n2518_1) );
  AND2X2 AND2X2_1270 ( .A(\bus_in[9] ), .B(key_en_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n4957) );
  AND2X2 AND2X2_1271 ( .A(AES_CORE_DATAPATH__abc_16259_n4955_1), .B(AES_CORE_DATAPATH__abc_16259_n4959), .Y(AES_CORE_DATAPATH__abc_16259_n4960) );
  AND2X2 AND2X2_1272 ( .A(AES_CORE_DATAPATH__abc_16259_n4960), .B(AES_CORE_DATAPATH__abc_16259_n4873_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n4961_1) );
  AND2X2 AND2X2_1273 ( .A(AES_CORE_DATAPATH__abc_16259_n4872_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__9_), .Y(AES_CORE_DATAPATH__abc_16259_n4962) );
  AND2X2 AND2X2_1274 ( .A(AES_CORE_DATAPATH__abc_16259_n4867_1_bF_buf3), .B(AES_CORE_DATAPATH_key_host_1__10_), .Y(AES_CORE_DATAPATH__abc_16259_n4965) );
  AND2X2 AND2X2_1275 ( .A(\bus_in[10] ), .B(key_en_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n4966) );
  AND2X2 AND2X2_1276 ( .A(AES_CORE_DATAPATH__abc_16259_n4964_1), .B(AES_CORE_DATAPATH__abc_16259_n4968), .Y(AES_CORE_DATAPATH__abc_16259_n4969) );
  AND2X2 AND2X2_1277 ( .A(AES_CORE_DATAPATH__abc_16259_n4970_1), .B(AES_CORE_DATAPATH__abc_16259_n4971), .Y(AES_CORE_DATAPATH__0key_1__31_0__10_) );
  AND2X2 AND2X2_1278 ( .A(AES_CORE_DATAPATH__abc_16259_n4867_1_bF_buf2), .B(AES_CORE_DATAPATH_key_host_1__11_), .Y(AES_CORE_DATAPATH__abc_16259_n4974) );
  AND2X2 AND2X2_1279 ( .A(\bus_in[11] ), .B(key_en_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n4975) );
  AND2X2 AND2X2_128 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf2), .B(AES_CORE_DATAPATH_iv_1__4_), .Y(AES_CORE_DATAPATH__abc_16259_n2519_1) );
  AND2X2 AND2X2_1280 ( .A(AES_CORE_DATAPATH__abc_16259_n4973_1), .B(AES_CORE_DATAPATH__abc_16259_n4977), .Y(AES_CORE_DATAPATH__abc_16259_n4978) );
  AND2X2 AND2X2_1281 ( .A(AES_CORE_DATAPATH__abc_16259_n4978), .B(AES_CORE_DATAPATH__abc_16259_n4873_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n4979_1) );
  AND2X2 AND2X2_1282 ( .A(AES_CORE_DATAPATH__abc_16259_n4872_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__11_), .Y(AES_CORE_DATAPATH__abc_16259_n4980_1) );
  AND2X2 AND2X2_1283 ( .A(AES_CORE_DATAPATH__abc_16259_n4867_1_bF_buf1), .B(AES_CORE_DATAPATH_key_host_1__12_), .Y(AES_CORE_DATAPATH__abc_16259_n4983_1) );
  AND2X2 AND2X2_1284 ( .A(\bus_in[12] ), .B(key_en_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n4984_1) );
  AND2X2 AND2X2_1285 ( .A(AES_CORE_DATAPATH__abc_16259_n4982_1), .B(AES_CORE_DATAPATH__abc_16259_n4986_1), .Y(AES_CORE_DATAPATH__abc_16259_n4987_1) );
  AND2X2 AND2X2_1286 ( .A(AES_CORE_DATAPATH__abc_16259_n4987_1), .B(AES_CORE_DATAPATH__abc_16259_n4873_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n4988_1) );
  AND2X2 AND2X2_1287 ( .A(AES_CORE_DATAPATH__abc_16259_n4872_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__12_), .Y(AES_CORE_DATAPATH__abc_16259_n4989_1) );
  AND2X2 AND2X2_1288 ( .A(AES_CORE_DATAPATH__abc_16259_n4867_1_bF_buf0), .B(AES_CORE_DATAPATH_key_host_1__13_), .Y(AES_CORE_DATAPATH__abc_16259_n4992_1) );
  AND2X2 AND2X2_1289 ( .A(\bus_in[13] ), .B(key_en_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n4993_1) );
  AND2X2 AND2X2_129 ( .A(AES_CORE_DATAPATH__abc_16259_n2522), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n2523_1) );
  AND2X2 AND2X2_1290 ( .A(AES_CORE_DATAPATH__abc_16259_n4991_1), .B(AES_CORE_DATAPATH__abc_16259_n4995_1), .Y(AES_CORE_DATAPATH__abc_16259_n4996_1) );
  AND2X2 AND2X2_1291 ( .A(AES_CORE_DATAPATH__abc_16259_n4997_1), .B(AES_CORE_DATAPATH__abc_16259_n4998_1), .Y(AES_CORE_DATAPATH__0key_1__31_0__13_) );
  AND2X2 AND2X2_1292 ( .A(AES_CORE_DATAPATH__abc_16259_n4867_1_bF_buf4), .B(AES_CORE_DATAPATH_key_host_1__14_), .Y(AES_CORE_DATAPATH__abc_16259_n5001_1) );
  AND2X2 AND2X2_1293 ( .A(\bus_in[14] ), .B(key_en_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5002_1) );
  AND2X2 AND2X2_1294 ( .A(AES_CORE_DATAPATH__abc_16259_n5000_1), .B(AES_CORE_DATAPATH__abc_16259_n5004_1), .Y(AES_CORE_DATAPATH__abc_16259_n5005_1) );
  AND2X2 AND2X2_1295 ( .A(AES_CORE_DATAPATH__abc_16259_n5005_1), .B(AES_CORE_DATAPATH__abc_16259_n4873_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n5006_1) );
  AND2X2 AND2X2_1296 ( .A(AES_CORE_DATAPATH__abc_16259_n4872_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__14_), .Y(AES_CORE_DATAPATH__abc_16259_n5007_1) );
  AND2X2 AND2X2_1297 ( .A(AES_CORE_DATAPATH__abc_16259_n4867_1_bF_buf3), .B(AES_CORE_DATAPATH_key_host_1__15_), .Y(AES_CORE_DATAPATH__abc_16259_n5010_1) );
  AND2X2 AND2X2_1298 ( .A(\bus_in[15] ), .B(key_en_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n5011_1) );
  AND2X2 AND2X2_1299 ( .A(AES_CORE_DATAPATH__abc_16259_n5009_1), .B(AES_CORE_DATAPATH__abc_16259_n5013), .Y(AES_CORE_DATAPATH__abc_16259_n5014_1) );
  AND2X2 AND2X2_13 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n85), .B(AES_CORE_CONTROL_UNIT_state_12_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n86_1) );
  AND2X2 AND2X2_130 ( .A(AES_CORE_DATAPATH__abc_16259_n2521_1), .B(AES_CORE_DATAPATH__abc_16259_n2523_1), .Y(AES_CORE_DATAPATH__abc_16259_n2524_1) );
  AND2X2 AND2X2_1300 ( .A(AES_CORE_DATAPATH__abc_16259_n5014_1), .B(AES_CORE_DATAPATH__abc_16259_n4873_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5015_1) );
  AND2X2 AND2X2_1301 ( .A(AES_CORE_DATAPATH__abc_16259_n4872_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__15_), .Y(AES_CORE_DATAPATH__abc_16259_n5016_1) );
  AND2X2 AND2X2_1302 ( .A(AES_CORE_DATAPATH__abc_16259_n4867_1_bF_buf2), .B(AES_CORE_DATAPATH_key_host_1__16_), .Y(AES_CORE_DATAPATH__abc_16259_n5019_1) );
  AND2X2 AND2X2_1303 ( .A(\bus_in[16] ), .B(key_en_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n5020_1) );
  AND2X2 AND2X2_1304 ( .A(AES_CORE_DATAPATH__abc_16259_n5018_1), .B(AES_CORE_DATAPATH__abc_16259_n5022_1), .Y(AES_CORE_DATAPATH__abc_16259_n5023_1) );
  AND2X2 AND2X2_1305 ( .A(AES_CORE_DATAPATH__abc_16259_n5023_1), .B(AES_CORE_DATAPATH__abc_16259_n4873_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n5024_1) );
  AND2X2 AND2X2_1306 ( .A(AES_CORE_DATAPATH__abc_16259_n4872_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__16_), .Y(AES_CORE_DATAPATH__abc_16259_n5025_1) );
  AND2X2 AND2X2_1307 ( .A(AES_CORE_DATAPATH__abc_16259_n4867_1_bF_buf1), .B(AES_CORE_DATAPATH_key_host_1__17_), .Y(AES_CORE_DATAPATH__abc_16259_n5028_1) );
  AND2X2 AND2X2_1308 ( .A(\bus_in[17] ), .B(key_en_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n5029_1) );
  AND2X2 AND2X2_1309 ( .A(AES_CORE_DATAPATH__abc_16259_n5027_1), .B(AES_CORE_DATAPATH__abc_16259_n5031_1), .Y(AES_CORE_DATAPATH__abc_16259_n5032_1) );
  AND2X2 AND2X2_131 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf2), .B(AES_CORE_DATAPATH_iv_3__4_), .Y(AES_CORE_DATAPATH__abc_16259_n2525) );
  AND2X2 AND2X2_1310 ( .A(AES_CORE_DATAPATH__abc_16259_n5033_1), .B(AES_CORE_DATAPATH__abc_16259_n5034_1), .Y(AES_CORE_DATAPATH__0key_1__31_0__17_) );
  AND2X2 AND2X2_1311 ( .A(AES_CORE_DATAPATH__abc_16259_n4867_1_bF_buf0), .B(AES_CORE_DATAPATH_key_host_1__18_), .Y(AES_CORE_DATAPATH__abc_16259_n5037_1) );
  AND2X2 AND2X2_1312 ( .A(\bus_in[18] ), .B(key_en_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n5038_1) );
  AND2X2 AND2X2_1313 ( .A(AES_CORE_DATAPATH__abc_16259_n5036_1), .B(AES_CORE_DATAPATH__abc_16259_n5040_1), .Y(AES_CORE_DATAPATH__abc_16259_n5041_1) );
  AND2X2 AND2X2_1314 ( .A(AES_CORE_DATAPATH__abc_16259_n5041_1), .B(AES_CORE_DATAPATH__abc_16259_n4873_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n5042_1) );
  AND2X2 AND2X2_1315 ( .A(AES_CORE_DATAPATH__abc_16259_n4872_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__18_), .Y(AES_CORE_DATAPATH__abc_16259_n5043_1) );
  AND2X2 AND2X2_1316 ( .A(AES_CORE_DATAPATH__abc_16259_n4867_1_bF_buf4), .B(AES_CORE_DATAPATH_key_host_1__19_), .Y(AES_CORE_DATAPATH__abc_16259_n5046_1) );
  AND2X2 AND2X2_1317 ( .A(\bus_in[19] ), .B(key_en_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5047_1) );
  AND2X2 AND2X2_1318 ( .A(AES_CORE_DATAPATH__abc_16259_n5045_1), .B(AES_CORE_DATAPATH__abc_16259_n5049_1), .Y(AES_CORE_DATAPATH__abc_16259_n5050_1) );
  AND2X2 AND2X2_1319 ( .A(AES_CORE_DATAPATH__abc_16259_n5051_1), .B(AES_CORE_DATAPATH__abc_16259_n5052_1), .Y(AES_CORE_DATAPATH__0key_1__31_0__19_) );
  AND2X2 AND2X2_132 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf2), .B(AES_CORE_DATAPATH_iv_0__5_), .Y(AES_CORE_DATAPATH__abc_16259_n2527) );
  AND2X2 AND2X2_1320 ( .A(AES_CORE_DATAPATH__abc_16259_n4867_1_bF_buf3), .B(AES_CORE_DATAPATH_key_host_1__20_), .Y(AES_CORE_DATAPATH__abc_16259_n5055_1) );
  AND2X2 AND2X2_1321 ( .A(\bus_in[20] ), .B(key_en_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n5056_1) );
  AND2X2 AND2X2_1322 ( .A(AES_CORE_DATAPATH__abc_16259_n5054_1), .B(AES_CORE_DATAPATH__abc_16259_n5058_1), .Y(AES_CORE_DATAPATH__abc_16259_n5059_1) );
  AND2X2 AND2X2_1323 ( .A(AES_CORE_DATAPATH__abc_16259_n5059_1), .B(AES_CORE_DATAPATH__abc_16259_n4873_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5060_1) );
  AND2X2 AND2X2_1324 ( .A(AES_CORE_DATAPATH__abc_16259_n4872_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__20_), .Y(AES_CORE_DATAPATH__abc_16259_n5061_1) );
  AND2X2 AND2X2_1325 ( .A(AES_CORE_DATAPATH__abc_16259_n4867_1_bF_buf2), .B(AES_CORE_DATAPATH_key_host_1__21_), .Y(AES_CORE_DATAPATH__abc_16259_n5064_1) );
  AND2X2 AND2X2_1326 ( .A(\bus_in[21] ), .B(key_en_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n5065_1) );
  AND2X2 AND2X2_1327 ( .A(AES_CORE_DATAPATH__abc_16259_n5063_1), .B(AES_CORE_DATAPATH__abc_16259_n5067_1), .Y(AES_CORE_DATAPATH__abc_16259_n5068_1) );
  AND2X2 AND2X2_1328 ( .A(AES_CORE_DATAPATH__abc_16259_n5069_1), .B(AES_CORE_DATAPATH__abc_16259_n5070_1), .Y(AES_CORE_DATAPATH__0key_1__31_0__21_) );
  AND2X2 AND2X2_1329 ( .A(AES_CORE_DATAPATH__abc_16259_n4867_1_bF_buf1), .B(AES_CORE_DATAPATH_key_host_1__22_), .Y(AES_CORE_DATAPATH__abc_16259_n5073_1) );
  AND2X2 AND2X2_133 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf1), .B(AES_CORE_DATAPATH_iv_1__5_), .Y(AES_CORE_DATAPATH__abc_16259_n2528_1) );
  AND2X2 AND2X2_1330 ( .A(\bus_in[22] ), .B(key_en_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n5074_1) );
  AND2X2 AND2X2_1331 ( .A(AES_CORE_DATAPATH__abc_16259_n5072_1), .B(AES_CORE_DATAPATH__abc_16259_n5076_1), .Y(AES_CORE_DATAPATH__abc_16259_n5077_1) );
  AND2X2 AND2X2_1332 ( .A(AES_CORE_DATAPATH__abc_16259_n5078), .B(AES_CORE_DATAPATH__abc_16259_n5079), .Y(AES_CORE_DATAPATH__0key_1__31_0__22_) );
  AND2X2 AND2X2_1333 ( .A(AES_CORE_DATAPATH__abc_16259_n4867_1_bF_buf0), .B(AES_CORE_DATAPATH_key_host_1__23_), .Y(AES_CORE_DATAPATH__abc_16259_n5082) );
  AND2X2 AND2X2_1334 ( .A(\bus_in[23] ), .B(key_en_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n5083_1) );
  AND2X2 AND2X2_1335 ( .A(AES_CORE_DATAPATH__abc_16259_n5081), .B(AES_CORE_DATAPATH__abc_16259_n5085), .Y(AES_CORE_DATAPATH__abc_16259_n5086_1) );
  AND2X2 AND2X2_1336 ( .A(AES_CORE_DATAPATH__abc_16259_n5086_1), .B(AES_CORE_DATAPATH__abc_16259_n4873_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n5087) );
  AND2X2 AND2X2_1337 ( .A(AES_CORE_DATAPATH__abc_16259_n4872_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__23_), .Y(AES_CORE_DATAPATH__abc_16259_n5088) );
  AND2X2 AND2X2_1338 ( .A(AES_CORE_DATAPATH__abc_16259_n4867_1_bF_buf4), .B(AES_CORE_DATAPATH_key_host_1__24_), .Y(AES_CORE_DATAPATH__abc_16259_n5091) );
  AND2X2 AND2X2_1339 ( .A(\bus_in[24] ), .B(key_en_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5092_1) );
  AND2X2 AND2X2_134 ( .A(AES_CORE_DATAPATH__abc_16259_n2531_1), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n2532) );
  AND2X2 AND2X2_1340 ( .A(AES_CORE_DATAPATH__abc_16259_n5090), .B(AES_CORE_DATAPATH__abc_16259_n5094), .Y(AES_CORE_DATAPATH__abc_16259_n5095_1) );
  AND2X2 AND2X2_1341 ( .A(AES_CORE_DATAPATH__abc_16259_n5096), .B(AES_CORE_DATAPATH__abc_16259_n5097), .Y(AES_CORE_DATAPATH__0key_1__31_0__24_) );
  AND2X2 AND2X2_1342 ( .A(AES_CORE_DATAPATH__abc_16259_n4867_1_bF_buf3), .B(AES_CORE_DATAPATH_key_host_1__25_), .Y(AES_CORE_DATAPATH__abc_16259_n5100) );
  AND2X2 AND2X2_1343 ( .A(\bus_in[25] ), .B(key_en_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n5101_1) );
  AND2X2 AND2X2_1344 ( .A(AES_CORE_DATAPATH__abc_16259_n5099), .B(AES_CORE_DATAPATH__abc_16259_n5103), .Y(AES_CORE_DATAPATH__abc_16259_n5104_1) );
  AND2X2 AND2X2_1345 ( .A(AES_CORE_DATAPATH__abc_16259_n5104_1), .B(AES_CORE_DATAPATH__abc_16259_n4873_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5105) );
  AND2X2 AND2X2_1346 ( .A(AES_CORE_DATAPATH__abc_16259_n4872_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__25_), .Y(AES_CORE_DATAPATH__abc_16259_n5106) );
  AND2X2 AND2X2_1347 ( .A(AES_CORE_DATAPATH__abc_16259_n4867_1_bF_buf2), .B(AES_CORE_DATAPATH_key_host_1__26_), .Y(AES_CORE_DATAPATH__abc_16259_n5109) );
  AND2X2 AND2X2_1348 ( .A(\bus_in[26] ), .B(key_en_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n5110_1) );
  AND2X2 AND2X2_1349 ( .A(AES_CORE_DATAPATH__abc_16259_n5108), .B(AES_CORE_DATAPATH__abc_16259_n5112), .Y(AES_CORE_DATAPATH__abc_16259_n5113_1) );
  AND2X2 AND2X2_135 ( .A(AES_CORE_DATAPATH__abc_16259_n2530), .B(AES_CORE_DATAPATH__abc_16259_n2532), .Y(AES_CORE_DATAPATH__abc_16259_n2533_1) );
  AND2X2 AND2X2_1350 ( .A(AES_CORE_DATAPATH__abc_16259_n5114), .B(AES_CORE_DATAPATH__abc_16259_n5115), .Y(AES_CORE_DATAPATH__0key_1__31_0__26_) );
  AND2X2 AND2X2_1351 ( .A(AES_CORE_DATAPATH__abc_16259_n4867_1_bF_buf1), .B(AES_CORE_DATAPATH_key_host_1__27_), .Y(AES_CORE_DATAPATH__abc_16259_n5118) );
  AND2X2 AND2X2_1352 ( .A(\bus_in[27] ), .B(key_en_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n5119_1) );
  AND2X2 AND2X2_1353 ( .A(AES_CORE_DATAPATH__abc_16259_n5117), .B(AES_CORE_DATAPATH__abc_16259_n5121), .Y(AES_CORE_DATAPATH__abc_16259_n5122_1) );
  AND2X2 AND2X2_1354 ( .A(AES_CORE_DATAPATH__abc_16259_n5122_1), .B(AES_CORE_DATAPATH__abc_16259_n4873_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n5123) );
  AND2X2 AND2X2_1355 ( .A(AES_CORE_DATAPATH__abc_16259_n4872_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__27_), .Y(AES_CORE_DATAPATH__abc_16259_n5124) );
  AND2X2 AND2X2_1356 ( .A(AES_CORE_DATAPATH__abc_16259_n4867_1_bF_buf0), .B(AES_CORE_DATAPATH_key_host_1__28_), .Y(AES_CORE_DATAPATH__abc_16259_n5127) );
  AND2X2 AND2X2_1357 ( .A(\bus_in[28] ), .B(key_en_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n5128_1) );
  AND2X2 AND2X2_1358 ( .A(AES_CORE_DATAPATH__abc_16259_n5126), .B(AES_CORE_DATAPATH__abc_16259_n5130), .Y(AES_CORE_DATAPATH__abc_16259_n5131_1) );
  AND2X2 AND2X2_1359 ( .A(AES_CORE_DATAPATH__abc_16259_n5132), .B(AES_CORE_DATAPATH__abc_16259_n5133), .Y(AES_CORE_DATAPATH__0key_1__31_0__28_) );
  AND2X2 AND2X2_136 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf1), .B(AES_CORE_DATAPATH_iv_3__5_), .Y(AES_CORE_DATAPATH__abc_16259_n2534_1) );
  AND2X2 AND2X2_1360 ( .A(AES_CORE_DATAPATH__abc_16259_n4867_1_bF_buf4), .B(AES_CORE_DATAPATH_key_host_1__29_), .Y(AES_CORE_DATAPATH__abc_16259_n5136) );
  AND2X2 AND2X2_1361 ( .A(\bus_in[29] ), .B(key_en_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5137_1) );
  AND2X2 AND2X2_1362 ( .A(AES_CORE_DATAPATH__abc_16259_n5135), .B(AES_CORE_DATAPATH__abc_16259_n5139), .Y(AES_CORE_DATAPATH__abc_16259_n5140_1) );
  AND2X2 AND2X2_1363 ( .A(AES_CORE_DATAPATH__abc_16259_n5141), .B(AES_CORE_DATAPATH__abc_16259_n5142), .Y(AES_CORE_DATAPATH__0key_1__31_0__29_) );
  AND2X2 AND2X2_1364 ( .A(AES_CORE_DATAPATH__abc_16259_n4867_1_bF_buf3), .B(AES_CORE_DATAPATH_key_host_1__30_), .Y(AES_CORE_DATAPATH__abc_16259_n5145) );
  AND2X2 AND2X2_1365 ( .A(\bus_in[30] ), .B(key_en_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n5146_1) );
  AND2X2 AND2X2_1366 ( .A(AES_CORE_DATAPATH__abc_16259_n5144), .B(AES_CORE_DATAPATH__abc_16259_n5148), .Y(AES_CORE_DATAPATH__abc_16259_n5149_1) );
  AND2X2 AND2X2_1367 ( .A(AES_CORE_DATAPATH__abc_16259_n5150), .B(AES_CORE_DATAPATH__abc_16259_n5151), .Y(AES_CORE_DATAPATH__0key_1__31_0__30_) );
  AND2X2 AND2X2_1368 ( .A(AES_CORE_DATAPATH__abc_16259_n4867_1_bF_buf2), .B(AES_CORE_DATAPATH_key_host_1__31_), .Y(AES_CORE_DATAPATH__abc_16259_n5153) );
  AND2X2 AND2X2_1369 ( .A(\bus_in[31] ), .B(key_en_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n5154) );
  AND2X2 AND2X2_137 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf1), .B(AES_CORE_DATAPATH_iv_0__6_), .Y(AES_CORE_DATAPATH__abc_16259_n2536_1) );
  AND2X2 AND2X2_1370 ( .A(AES_CORE_DATAPATH__abc_16259_n5157), .B(AES_CORE_DATAPATH__abc_16259_n5156), .Y(AES_CORE_DATAPATH__abc_16259_n5158_1) );
  AND2X2 AND2X2_1371 ( .A(AES_CORE_DATAPATH__abc_16259_n5158_1), .B(AES_CORE_DATAPATH__abc_16259_n4873_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n5159) );
  AND2X2 AND2X2_1372 ( .A(AES_CORE_DATAPATH__abc_16259_n4872_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__31_), .Y(AES_CORE_DATAPATH__abc_16259_n5160) );
  AND2X2 AND2X2_1373 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__0_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf10), .Y(AES_CORE_DATAPATH__abc_16259_n5162) );
  AND2X2 AND2X2_1374 ( .A(AES_CORE_DATAPATH__abc_16259_n4877_1), .B(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n5163) );
  AND2X2 AND2X2_1375 ( .A(AES_CORE_DATAPATH__abc_16259_n5166), .B(AES_CORE_DATAPATH__abc_16259_n5165), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__1_) );
  AND2X2 AND2X2_1376 ( .A(AES_CORE_DATAPATH__abc_16259_n5169), .B(AES_CORE_DATAPATH__abc_16259_n5168), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__2_) );
  AND2X2 AND2X2_1377 ( .A(AES_CORE_DATAPATH__abc_16259_n5172), .B(AES_CORE_DATAPATH__abc_16259_n5171), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__3_) );
  AND2X2 AND2X2_1378 ( .A(AES_CORE_DATAPATH__abc_16259_n5175_1), .B(AES_CORE_DATAPATH__abc_16259_n5174_1), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__4_) );
  AND2X2 AND2X2_1379 ( .A(AES_CORE_DATAPATH__abc_16259_n5178_1), .B(AES_CORE_DATAPATH__abc_16259_n5177_1), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__5_) );
  AND2X2 AND2X2_138 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf0), .B(AES_CORE_DATAPATH_iv_1__6_), .Y(AES_CORE_DATAPATH__abc_16259_n2537) );
  AND2X2 AND2X2_1380 ( .A(AES_CORE_DATAPATH__abc_16259_n5181_1), .B(AES_CORE_DATAPATH__abc_16259_n5180_1), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__6_) );
  AND2X2 AND2X2_1381 ( .A(AES_CORE_DATAPATH__abc_16259_n5184_1), .B(AES_CORE_DATAPATH__abc_16259_n5183_1), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__7_) );
  AND2X2 AND2X2_1382 ( .A(AES_CORE_DATAPATH__abc_16259_n5187_1), .B(AES_CORE_DATAPATH__abc_16259_n5186_1), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__8_) );
  AND2X2 AND2X2_1383 ( .A(AES_CORE_DATAPATH__abc_16259_n5190_1), .B(AES_CORE_DATAPATH__abc_16259_n5189_1), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__9_) );
  AND2X2 AND2X2_1384 ( .A(AES_CORE_DATAPATH__abc_16259_n5193_1), .B(AES_CORE_DATAPATH__abc_16259_n5192_1), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__10_) );
  AND2X2 AND2X2_1385 ( .A(AES_CORE_DATAPATH__abc_16259_n5196_1), .B(AES_CORE_DATAPATH__abc_16259_n5195_1), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__11_) );
  AND2X2 AND2X2_1386 ( .A(AES_CORE_DATAPATH__abc_16259_n5199_1), .B(AES_CORE_DATAPATH__abc_16259_n5198_1), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__12_) );
  AND2X2 AND2X2_1387 ( .A(AES_CORE_DATAPATH__abc_16259_n5202_1), .B(AES_CORE_DATAPATH__abc_16259_n5201_1), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__13_) );
  AND2X2 AND2X2_1388 ( .A(AES_CORE_DATAPATH__abc_16259_n5205_1), .B(AES_CORE_DATAPATH__abc_16259_n5204_1), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__14_) );
  AND2X2 AND2X2_1389 ( .A(AES_CORE_DATAPATH__abc_16259_n5208_1), .B(AES_CORE_DATAPATH__abc_16259_n5207), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__15_) );
  AND2X2 AND2X2_139 ( .A(AES_CORE_DATAPATH__abc_16259_n2540), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n2541_1) );
  AND2X2 AND2X2_1390 ( .A(AES_CORE_DATAPATH__abc_16259_n5211_1), .B(AES_CORE_DATAPATH__abc_16259_n5210_1), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__16_) );
  AND2X2 AND2X2_1391 ( .A(AES_CORE_DATAPATH__abc_16259_n5214_1), .B(AES_CORE_DATAPATH__abc_16259_n5213_1), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__17_) );
  AND2X2 AND2X2_1392 ( .A(AES_CORE_DATAPATH__abc_16259_n5217_1), .B(AES_CORE_DATAPATH__abc_16259_n5216_1), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__18_) );
  AND2X2 AND2X2_1393 ( .A(AES_CORE_DATAPATH__abc_16259_n5220_1), .B(AES_CORE_DATAPATH__abc_16259_n5219_1), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__19_) );
  AND2X2 AND2X2_1394 ( .A(AES_CORE_DATAPATH__abc_16259_n5223_1), .B(AES_CORE_DATAPATH__abc_16259_n5222_1), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__20_) );
  AND2X2 AND2X2_1395 ( .A(AES_CORE_DATAPATH__abc_16259_n5226_1), .B(AES_CORE_DATAPATH__abc_16259_n5225_1), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__21_) );
  AND2X2 AND2X2_1396 ( .A(AES_CORE_DATAPATH__abc_16259_n5229_1), .B(AES_CORE_DATAPATH__abc_16259_n5228_1), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__22_) );
  AND2X2 AND2X2_1397 ( .A(AES_CORE_DATAPATH__abc_16259_n5232_1), .B(AES_CORE_DATAPATH__abc_16259_n5231_1), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__23_) );
  AND2X2 AND2X2_1398 ( .A(AES_CORE_DATAPATH__abc_16259_n5235_1), .B(AES_CORE_DATAPATH__abc_16259_n5234_1), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__24_) );
  AND2X2 AND2X2_1399 ( .A(AES_CORE_DATAPATH__abc_16259_n5238_1), .B(AES_CORE_DATAPATH__abc_16259_n5237_1), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__25_) );
  AND2X2 AND2X2_14 ( .A(AES_CORE_CONTROL_UNIT_last_round_bF_buf5), .B(AES_CORE_CONTROL_UNIT__abc_15841_n84_1), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n87_1) );
  AND2X2 AND2X2_140 ( .A(AES_CORE_DATAPATH__abc_16259_n2539_1), .B(AES_CORE_DATAPATH__abc_16259_n2541_1), .Y(AES_CORE_DATAPATH__abc_16259_n2542) );
  AND2X2 AND2X2_1400 ( .A(AES_CORE_DATAPATH__abc_16259_n5241_1), .B(AES_CORE_DATAPATH__abc_16259_n5240_1), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__26_) );
  AND2X2 AND2X2_1401 ( .A(AES_CORE_DATAPATH__abc_16259_n5244_1), .B(AES_CORE_DATAPATH__abc_16259_n5243_1), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__27_) );
  AND2X2 AND2X2_1402 ( .A(AES_CORE_DATAPATH__abc_16259_n5247_1), .B(AES_CORE_DATAPATH__abc_16259_n5246_1), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__28_) );
  AND2X2 AND2X2_1403 ( .A(AES_CORE_DATAPATH__abc_16259_n5250_1), .B(AES_CORE_DATAPATH__abc_16259_n5249_1), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__29_) );
  AND2X2 AND2X2_1404 ( .A(AES_CORE_DATAPATH__abc_16259_n5253_1), .B(AES_CORE_DATAPATH__abc_16259_n5252_1), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__30_) );
  AND2X2 AND2X2_1405 ( .A(AES_CORE_DATAPATH__abc_16259_n5255_1), .B(AES_CORE_DATAPATH__abc_16259_n5256_1), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__31_) );
  AND2X2 AND2X2_1406 ( .A(AES_CORE_CONTROL_UNIT_bypass_key_en), .B(AES_CORE_CONTROL_UNIT_key_en_2_), .Y(AES_CORE_DATAPATH__abc_16259_n5258_1) );
  AND2X2 AND2X2_1407 ( .A(AES_CORE_DATAPATH__abc_16259_n4469_1), .B(AES_CORE_DATAPATH__abc_16259_n5260_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5261_1) );
  AND2X2 AND2X2_1408 ( .A(AES_CORE_DATAPATH__abc_16259_n2806_1), .B(AES_CORE_DATAPATH_key_en_pp1_2_), .Y(AES_CORE_DATAPATH__abc_16259_n5262_1) );
  AND2X2 AND2X2_1409 ( .A(AES_CORE_DATAPATH__abc_16259_n5263_1), .B(AES_CORE_DATAPATH__abc_16259_n5261_1), .Y(AES_CORE_DATAPATH__abc_16259_n5264_1) );
  AND2X2 AND2X2_141 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf0), .B(AES_CORE_DATAPATH_iv_3__6_), .Y(AES_CORE_DATAPATH__abc_16259_n2543_1) );
  AND2X2 AND2X2_1410 ( .A(AES_CORE_DATAPATH__abc_16259_n5264_1), .B(AES_CORE_DATAPATH__abc_16259_n5259_1), .Y(AES_CORE_DATAPATH__abc_16259_n5265_1) );
  AND2X2 AND2X2_1411 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_32_), .Y(AES_CORE_DATAPATH__abc_16259_n5267_1) );
  AND2X2 AND2X2_1412 ( .A(\bus_in[0] ), .B(key_en_2_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n5268_1) );
  AND2X2 AND2X2_1413 ( .A(AES_CORE_DATAPATH__abc_16259_n5260_1_bF_buf3), .B(AES_CORE_DATAPATH_key_host_2__0_), .Y(AES_CORE_DATAPATH__abc_16259_n5269_1) );
  AND2X2 AND2X2_1414 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n5270_1), .Y(AES_CORE_DATAPATH__abc_16259_n5271_1) );
  AND2X2 AND2X2_1415 ( .A(AES_CORE_DATAPATH__abc_16259_n5272), .B(AES_CORE_DATAPATH__abc_16259_n5266_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5273) );
  AND2X2 AND2X2_1416 ( .A(AES_CORE_DATAPATH__abc_16259_n5265_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__0_), .Y(AES_CORE_DATAPATH__abc_16259_n5274_1) );
  AND2X2 AND2X2_1417 ( .A(AES_CORE_DATAPATH__abc_16259_n5260_1_bF_buf2), .B(AES_CORE_DATAPATH_key_host_2__1_), .Y(AES_CORE_DATAPATH__abc_16259_n5277_1) );
  AND2X2 AND2X2_1418 ( .A(\bus_in[1] ), .B(key_en_2_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n5278) );
  AND2X2 AND2X2_1419 ( .A(AES_CORE_DATAPATH__abc_16259_n5276), .B(AES_CORE_DATAPATH__abc_16259_n5280_1), .Y(AES_CORE_DATAPATH__abc_16259_n5281) );
  AND2X2 AND2X2_142 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf0), .B(AES_CORE_DATAPATH_iv_0__7_), .Y(AES_CORE_DATAPATH__abc_16259_n2545) );
  AND2X2 AND2X2_1420 ( .A(AES_CORE_DATAPATH__abc_16259_n5281), .B(AES_CORE_DATAPATH__abc_16259_n5266_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n5282) );
  AND2X2 AND2X2_1421 ( .A(AES_CORE_DATAPATH__abc_16259_n5265_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__1_), .Y(AES_CORE_DATAPATH__abc_16259_n5283_1) );
  AND2X2 AND2X2_1422 ( .A(AES_CORE_DATAPATH__abc_16259_n5260_1_bF_buf1), .B(AES_CORE_DATAPATH_key_host_2__2_), .Y(AES_CORE_DATAPATH__abc_16259_n5286_1) );
  AND2X2 AND2X2_1423 ( .A(\bus_in[2] ), .B(key_en_2_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n5287) );
  AND2X2 AND2X2_1424 ( .A(AES_CORE_DATAPATH__abc_16259_n5285), .B(AES_CORE_DATAPATH__abc_16259_n5289_1), .Y(AES_CORE_DATAPATH__abc_16259_n5290) );
  AND2X2 AND2X2_1425 ( .A(AES_CORE_DATAPATH__abc_16259_n5290), .B(AES_CORE_DATAPATH__abc_16259_n5266_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n5291) );
  AND2X2 AND2X2_1426 ( .A(AES_CORE_DATAPATH__abc_16259_n5265_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__2_), .Y(AES_CORE_DATAPATH__abc_16259_n5292_1) );
  AND2X2 AND2X2_1427 ( .A(AES_CORE_DATAPATH__abc_16259_n5260_1_bF_buf0), .B(AES_CORE_DATAPATH_key_host_2__3_), .Y(AES_CORE_DATAPATH__abc_16259_n5295_1) );
  AND2X2 AND2X2_1428 ( .A(\bus_in[3] ), .B(key_en_2_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n5296) );
  AND2X2 AND2X2_1429 ( .A(AES_CORE_DATAPATH__abc_16259_n5294), .B(AES_CORE_DATAPATH__abc_16259_n5298_1), .Y(AES_CORE_DATAPATH__abc_16259_n5299) );
  AND2X2 AND2X2_143 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf7), .B(AES_CORE_DATAPATH_iv_1__7_), .Y(AES_CORE_DATAPATH__abc_16259_n2546_1) );
  AND2X2 AND2X2_1430 ( .A(AES_CORE_DATAPATH__abc_16259_n5299), .B(AES_CORE_DATAPATH__abc_16259_n5266_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n5300) );
  AND2X2 AND2X2_1431 ( .A(AES_CORE_DATAPATH__abc_16259_n5265_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__3_), .Y(AES_CORE_DATAPATH__abc_16259_n5301_1) );
  AND2X2 AND2X2_1432 ( .A(AES_CORE_DATAPATH__abc_16259_n5260_1_bF_buf4), .B(AES_CORE_DATAPATH_key_host_2__4_), .Y(AES_CORE_DATAPATH__abc_16259_n5304_1) );
  AND2X2 AND2X2_1433 ( .A(\bus_in[4] ), .B(key_en_2_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5305) );
  AND2X2 AND2X2_1434 ( .A(AES_CORE_DATAPATH__abc_16259_n5303), .B(AES_CORE_DATAPATH__abc_16259_n5307_1), .Y(AES_CORE_DATAPATH__abc_16259_n5308) );
  AND2X2 AND2X2_1435 ( .A(AES_CORE_DATAPATH__abc_16259_n5308), .B(AES_CORE_DATAPATH__abc_16259_n5266_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n5309) );
  AND2X2 AND2X2_1436 ( .A(AES_CORE_DATAPATH__abc_16259_n5265_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__4_), .Y(AES_CORE_DATAPATH__abc_16259_n5310_1) );
  AND2X2 AND2X2_1437 ( .A(AES_CORE_DATAPATH__abc_16259_n5260_1_bF_buf3), .B(AES_CORE_DATAPATH_key_host_2__5_), .Y(AES_CORE_DATAPATH__abc_16259_n5313_1) );
  AND2X2 AND2X2_1438 ( .A(\bus_in[5] ), .B(key_en_2_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n5314) );
  AND2X2 AND2X2_1439 ( .A(AES_CORE_DATAPATH__abc_16259_n5312), .B(AES_CORE_DATAPATH__abc_16259_n5316_1), .Y(AES_CORE_DATAPATH__abc_16259_n5317) );
  AND2X2 AND2X2_144 ( .A(AES_CORE_DATAPATH__abc_16259_n2549_1), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n2550) );
  AND2X2 AND2X2_1440 ( .A(AES_CORE_DATAPATH__abc_16259_n5317), .B(AES_CORE_DATAPATH__abc_16259_n5266_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5318) );
  AND2X2 AND2X2_1441 ( .A(AES_CORE_DATAPATH__abc_16259_n5265_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__5_), .Y(AES_CORE_DATAPATH__abc_16259_n5319_1) );
  AND2X2 AND2X2_1442 ( .A(AES_CORE_DATAPATH__abc_16259_n5260_1_bF_buf2), .B(AES_CORE_DATAPATH_key_host_2__6_), .Y(AES_CORE_DATAPATH__abc_16259_n5322_1) );
  AND2X2 AND2X2_1443 ( .A(\bus_in[6] ), .B(key_en_2_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n5323) );
  AND2X2 AND2X2_1444 ( .A(AES_CORE_DATAPATH__abc_16259_n5321), .B(AES_CORE_DATAPATH__abc_16259_n5325_1), .Y(AES_CORE_DATAPATH__abc_16259_n5326) );
  AND2X2 AND2X2_1445 ( .A(AES_CORE_DATAPATH__abc_16259_n5326), .B(AES_CORE_DATAPATH__abc_16259_n5266_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n5327) );
  AND2X2 AND2X2_1446 ( .A(AES_CORE_DATAPATH__abc_16259_n5265_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__6_), .Y(AES_CORE_DATAPATH__abc_16259_n5328_1) );
  AND2X2 AND2X2_1447 ( .A(AES_CORE_DATAPATH__abc_16259_n5260_1_bF_buf1), .B(AES_CORE_DATAPATH_key_host_2__7_), .Y(AES_CORE_DATAPATH__abc_16259_n5331_1) );
  AND2X2 AND2X2_1448 ( .A(\bus_in[7] ), .B(key_en_2_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n5332) );
  AND2X2 AND2X2_1449 ( .A(AES_CORE_DATAPATH__abc_16259_n5330), .B(AES_CORE_DATAPATH__abc_16259_n5334_1), .Y(AES_CORE_DATAPATH__abc_16259_n5335) );
  AND2X2 AND2X2_145 ( .A(AES_CORE_DATAPATH__abc_16259_n2548_1), .B(AES_CORE_DATAPATH__abc_16259_n2550), .Y(AES_CORE_DATAPATH__abc_16259_n2551_1) );
  AND2X2 AND2X2_1450 ( .A(AES_CORE_DATAPATH__abc_16259_n5335), .B(AES_CORE_DATAPATH__abc_16259_n5266_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n5336) );
  AND2X2 AND2X2_1451 ( .A(AES_CORE_DATAPATH__abc_16259_n5265_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__7_), .Y(AES_CORE_DATAPATH__abc_16259_n5337_1) );
  AND2X2 AND2X2_1452 ( .A(AES_CORE_DATAPATH__abc_16259_n5260_1_bF_buf0), .B(AES_CORE_DATAPATH_key_host_2__8_), .Y(AES_CORE_DATAPATH__abc_16259_n5340_1) );
  AND2X2 AND2X2_1453 ( .A(\bus_in[8] ), .B(key_en_2_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n5341) );
  AND2X2 AND2X2_1454 ( .A(AES_CORE_DATAPATH__abc_16259_n5339), .B(AES_CORE_DATAPATH__abc_16259_n5343_1), .Y(AES_CORE_DATAPATH__abc_16259_n5344) );
  AND2X2 AND2X2_1455 ( .A(AES_CORE_DATAPATH__abc_16259_n5344), .B(AES_CORE_DATAPATH__abc_16259_n5266_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n5345) );
  AND2X2 AND2X2_1456 ( .A(AES_CORE_DATAPATH__abc_16259_n5265_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__8_), .Y(AES_CORE_DATAPATH__abc_16259_n5346_1) );
  AND2X2 AND2X2_1457 ( .A(AES_CORE_DATAPATH__abc_16259_n5260_1_bF_buf4), .B(AES_CORE_DATAPATH_key_host_2__9_), .Y(AES_CORE_DATAPATH__abc_16259_n5349_1) );
  AND2X2 AND2X2_1458 ( .A(\bus_in[9] ), .B(key_en_2_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5350) );
  AND2X2 AND2X2_1459 ( .A(AES_CORE_DATAPATH__abc_16259_n5348), .B(AES_CORE_DATAPATH__abc_16259_n5352_1), .Y(AES_CORE_DATAPATH__abc_16259_n5353) );
  AND2X2 AND2X2_146 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf7), .B(AES_CORE_DATAPATH_iv_3__7_), .Y(AES_CORE_DATAPATH__abc_16259_n2552) );
  AND2X2 AND2X2_1460 ( .A(AES_CORE_DATAPATH__abc_16259_n5353), .B(AES_CORE_DATAPATH__abc_16259_n5266_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n5354) );
  AND2X2 AND2X2_1461 ( .A(AES_CORE_DATAPATH__abc_16259_n5265_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__9_), .Y(AES_CORE_DATAPATH__abc_16259_n5355_1) );
  AND2X2 AND2X2_1462 ( .A(AES_CORE_DATAPATH__abc_16259_n5260_1_bF_buf3), .B(AES_CORE_DATAPATH_key_host_2__10_), .Y(AES_CORE_DATAPATH__abc_16259_n5358_1) );
  AND2X2 AND2X2_1463 ( .A(\bus_in[10] ), .B(key_en_2_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n5359) );
  AND2X2 AND2X2_1464 ( .A(AES_CORE_DATAPATH__abc_16259_n5357), .B(AES_CORE_DATAPATH__abc_16259_n5361_1), .Y(AES_CORE_DATAPATH__abc_16259_n5362) );
  AND2X2 AND2X2_1465 ( .A(AES_CORE_DATAPATH__abc_16259_n5362), .B(AES_CORE_DATAPATH__abc_16259_n5266_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5363) );
  AND2X2 AND2X2_1466 ( .A(AES_CORE_DATAPATH__abc_16259_n5265_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__10_), .Y(AES_CORE_DATAPATH__abc_16259_n5364_1) );
  AND2X2 AND2X2_1467 ( .A(AES_CORE_DATAPATH__abc_16259_n5260_1_bF_buf2), .B(AES_CORE_DATAPATH_key_host_2__11_), .Y(AES_CORE_DATAPATH__abc_16259_n5367_1) );
  AND2X2 AND2X2_1468 ( .A(\bus_in[11] ), .B(key_en_2_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n5368_1) );
  AND2X2 AND2X2_1469 ( .A(AES_CORE_DATAPATH__abc_16259_n5366), .B(AES_CORE_DATAPATH__abc_16259_n5370_1), .Y(AES_CORE_DATAPATH__abc_16259_n5371_1) );
  AND2X2 AND2X2_147 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf7), .B(AES_CORE_DATAPATH_iv_0__8_), .Y(AES_CORE_DATAPATH__abc_16259_n2554_1) );
  AND2X2 AND2X2_1470 ( .A(AES_CORE_DATAPATH__abc_16259_n5371_1), .B(AES_CORE_DATAPATH__abc_16259_n5266_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n5372_1) );
  AND2X2 AND2X2_1471 ( .A(AES_CORE_DATAPATH__abc_16259_n5265_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__11_), .Y(AES_CORE_DATAPATH__abc_16259_n5373_1) );
  AND2X2 AND2X2_1472 ( .A(AES_CORE_DATAPATH__abc_16259_n5260_1_bF_buf1), .B(AES_CORE_DATAPATH_key_host_2__12_), .Y(AES_CORE_DATAPATH__abc_16259_n5376_1) );
  AND2X2 AND2X2_1473 ( .A(\bus_in[12] ), .B(key_en_2_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n5377_1) );
  AND2X2 AND2X2_1474 ( .A(AES_CORE_DATAPATH__abc_16259_n5375_1), .B(AES_CORE_DATAPATH__abc_16259_n5379_1), .Y(AES_CORE_DATAPATH__abc_16259_n5380_1) );
  AND2X2 AND2X2_1475 ( .A(AES_CORE_DATAPATH__abc_16259_n5380_1), .B(AES_CORE_DATAPATH__abc_16259_n5266_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n5381_1) );
  AND2X2 AND2X2_1476 ( .A(AES_CORE_DATAPATH__abc_16259_n5265_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__12_), .Y(AES_CORE_DATAPATH__abc_16259_n5382_1) );
  AND2X2 AND2X2_1477 ( .A(AES_CORE_DATAPATH__abc_16259_n5260_1_bF_buf0), .B(AES_CORE_DATAPATH_key_host_2__13_), .Y(AES_CORE_DATAPATH__abc_16259_n5385_1) );
  AND2X2 AND2X2_1478 ( .A(\bus_in[13] ), .B(key_en_2_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n5386_1) );
  AND2X2 AND2X2_1479 ( .A(AES_CORE_DATAPATH__abc_16259_n5384_1), .B(AES_CORE_DATAPATH__abc_16259_n5388_1), .Y(AES_CORE_DATAPATH__abc_16259_n5389_1) );
  AND2X2 AND2X2_148 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf6), .B(AES_CORE_DATAPATH_iv_1__8_), .Y(AES_CORE_DATAPATH__abc_16259_n2555) );
  AND2X2 AND2X2_1480 ( .A(AES_CORE_DATAPATH__abc_16259_n5389_1), .B(AES_CORE_DATAPATH__abc_16259_n5266_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n5390_1) );
  AND2X2 AND2X2_1481 ( .A(AES_CORE_DATAPATH__abc_16259_n5265_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__13_), .Y(AES_CORE_DATAPATH__abc_16259_n5391_1) );
  AND2X2 AND2X2_1482 ( .A(AES_CORE_DATAPATH__abc_16259_n5260_1_bF_buf4), .B(AES_CORE_DATAPATH_key_host_2__14_), .Y(AES_CORE_DATAPATH__abc_16259_n5394_1) );
  AND2X2 AND2X2_1483 ( .A(\bus_in[14] ), .B(key_en_2_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5395_1) );
  AND2X2 AND2X2_1484 ( .A(AES_CORE_DATAPATH__abc_16259_n5393_1), .B(AES_CORE_DATAPATH__abc_16259_n5397_1), .Y(AES_CORE_DATAPATH__abc_16259_n5398_1) );
  AND2X2 AND2X2_1485 ( .A(AES_CORE_DATAPATH__abc_16259_n5398_1), .B(AES_CORE_DATAPATH__abc_16259_n5266_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n5399_1) );
  AND2X2 AND2X2_1486 ( .A(AES_CORE_DATAPATH__abc_16259_n5265_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__14_), .Y(AES_CORE_DATAPATH__abc_16259_n5400_1) );
  AND2X2 AND2X2_1487 ( .A(AES_CORE_DATAPATH__abc_16259_n5260_1_bF_buf3), .B(AES_CORE_DATAPATH_key_host_2__15_), .Y(AES_CORE_DATAPATH__abc_16259_n5403_1) );
  AND2X2 AND2X2_1488 ( .A(\bus_in[15] ), .B(key_en_2_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n5404_1) );
  AND2X2 AND2X2_1489 ( .A(AES_CORE_DATAPATH__abc_16259_n5402_1), .B(AES_CORE_DATAPATH__abc_16259_n5406_1), .Y(AES_CORE_DATAPATH__abc_16259_n5407_1) );
  AND2X2 AND2X2_149 ( .A(AES_CORE_DATAPATH__abc_16259_n2558_1), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n2559_1) );
  AND2X2 AND2X2_1490 ( .A(AES_CORE_DATAPATH__abc_16259_n5407_1), .B(AES_CORE_DATAPATH__abc_16259_n5266_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5408_1) );
  AND2X2 AND2X2_1491 ( .A(AES_CORE_DATAPATH__abc_16259_n5265_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__15_), .Y(AES_CORE_DATAPATH__abc_16259_n5409_1) );
  AND2X2 AND2X2_1492 ( .A(AES_CORE_DATAPATH__abc_16259_n5260_1_bF_buf2), .B(AES_CORE_DATAPATH_key_host_2__16_), .Y(AES_CORE_DATAPATH__abc_16259_n5412_1) );
  AND2X2 AND2X2_1493 ( .A(\bus_in[16] ), .B(key_en_2_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n5413_1) );
  AND2X2 AND2X2_1494 ( .A(AES_CORE_DATAPATH__abc_16259_n5411_1), .B(AES_CORE_DATAPATH__abc_16259_n5415_1), .Y(AES_CORE_DATAPATH__abc_16259_n5416_1) );
  AND2X2 AND2X2_1495 ( .A(AES_CORE_DATAPATH__abc_16259_n5416_1), .B(AES_CORE_DATAPATH__abc_16259_n5266_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n5417_1) );
  AND2X2 AND2X2_1496 ( .A(AES_CORE_DATAPATH__abc_16259_n5265_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__16_), .Y(AES_CORE_DATAPATH__abc_16259_n5418_1) );
  AND2X2 AND2X2_1497 ( .A(AES_CORE_DATAPATH__abc_16259_n5260_1_bF_buf1), .B(AES_CORE_DATAPATH_key_host_2__17_), .Y(AES_CORE_DATAPATH__abc_16259_n5421_1) );
  AND2X2 AND2X2_1498 ( .A(\bus_in[17] ), .B(key_en_2_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n5422_1) );
  AND2X2 AND2X2_1499 ( .A(AES_CORE_DATAPATH__abc_16259_n5420_1), .B(AES_CORE_DATAPATH__abc_16259_n5424_1), .Y(AES_CORE_DATAPATH__abc_16259_n5425_1) );
  AND2X2 AND2X2_15 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n89_1), .B(\op_mode[0] ), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n90) );
  AND2X2 AND2X2_150 ( .A(AES_CORE_DATAPATH__abc_16259_n2557), .B(AES_CORE_DATAPATH__abc_16259_n2559_1), .Y(AES_CORE_DATAPATH__abc_16259_n2560) );
  AND2X2 AND2X2_1500 ( .A(AES_CORE_DATAPATH__abc_16259_n5425_1), .B(AES_CORE_DATAPATH__abc_16259_n5266_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n5426_1) );
  AND2X2 AND2X2_1501 ( .A(AES_CORE_DATAPATH__abc_16259_n5265_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__17_), .Y(AES_CORE_DATAPATH__abc_16259_n5427_1) );
  AND2X2 AND2X2_1502 ( .A(AES_CORE_DATAPATH__abc_16259_n5260_1_bF_buf0), .B(AES_CORE_DATAPATH_key_host_2__18_), .Y(AES_CORE_DATAPATH__abc_16259_n5430_1) );
  AND2X2 AND2X2_1503 ( .A(\bus_in[18] ), .B(key_en_2_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n5431_1) );
  AND2X2 AND2X2_1504 ( .A(AES_CORE_DATAPATH__abc_16259_n5429_1), .B(AES_CORE_DATAPATH__abc_16259_n5433_1), .Y(AES_CORE_DATAPATH__abc_16259_n5434_1) );
  AND2X2 AND2X2_1505 ( .A(AES_CORE_DATAPATH__abc_16259_n5434_1), .B(AES_CORE_DATAPATH__abc_16259_n5266_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n5435_1) );
  AND2X2 AND2X2_1506 ( .A(AES_CORE_DATAPATH__abc_16259_n5265_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__18_), .Y(AES_CORE_DATAPATH__abc_16259_n5436_1) );
  AND2X2 AND2X2_1507 ( .A(AES_CORE_DATAPATH__abc_16259_n5260_1_bF_buf4), .B(AES_CORE_DATAPATH_key_host_2__19_), .Y(AES_CORE_DATAPATH__abc_16259_n5439_1) );
  AND2X2 AND2X2_1508 ( .A(\bus_in[19] ), .B(key_en_2_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5440_1) );
  AND2X2 AND2X2_1509 ( .A(AES_CORE_DATAPATH__abc_16259_n5438_1), .B(AES_CORE_DATAPATH__abc_16259_n5442_1), .Y(AES_CORE_DATAPATH__abc_16259_n5443_1) );
  AND2X2 AND2X2_151 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf6), .B(AES_CORE_DATAPATH_iv_3__8_), .Y(AES_CORE_DATAPATH__abc_16259_n2561_1) );
  AND2X2 AND2X2_1510 ( .A(AES_CORE_DATAPATH__abc_16259_n5443_1), .B(AES_CORE_DATAPATH__abc_16259_n5266_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n5444_1) );
  AND2X2 AND2X2_1511 ( .A(AES_CORE_DATAPATH__abc_16259_n5265_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__19_), .Y(AES_CORE_DATAPATH__abc_16259_n5445_1) );
  AND2X2 AND2X2_1512 ( .A(AES_CORE_DATAPATH__abc_16259_n5260_1_bF_buf3), .B(AES_CORE_DATAPATH_key_host_2__20_), .Y(AES_CORE_DATAPATH__abc_16259_n5448_1) );
  AND2X2 AND2X2_1513 ( .A(\bus_in[20] ), .B(key_en_2_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n5449_1) );
  AND2X2 AND2X2_1514 ( .A(AES_CORE_DATAPATH__abc_16259_n5447_1), .B(AES_CORE_DATAPATH__abc_16259_n5451_1), .Y(AES_CORE_DATAPATH__abc_16259_n5452) );
  AND2X2 AND2X2_1515 ( .A(AES_CORE_DATAPATH__abc_16259_n5452), .B(AES_CORE_DATAPATH__abc_16259_n5266_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5453) );
  AND2X2 AND2X2_1516 ( .A(AES_CORE_DATAPATH__abc_16259_n5265_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__20_), .Y(AES_CORE_DATAPATH__abc_16259_n5454) );
  AND2X2 AND2X2_1517 ( .A(AES_CORE_DATAPATH__abc_16259_n5260_1_bF_buf2), .B(AES_CORE_DATAPATH_key_host_2__21_), .Y(AES_CORE_DATAPATH__abc_16259_n5457) );
  AND2X2 AND2X2_1518 ( .A(\bus_in[21] ), .B(key_en_2_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n5458) );
  AND2X2 AND2X2_1519 ( .A(AES_CORE_DATAPATH__abc_16259_n5456), .B(AES_CORE_DATAPATH__abc_16259_n5460), .Y(AES_CORE_DATAPATH__abc_16259_n5461) );
  AND2X2 AND2X2_152 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf6), .B(AES_CORE_DATAPATH_iv_0__9_), .Y(AES_CORE_DATAPATH__abc_16259_n2563_1) );
  AND2X2 AND2X2_1520 ( .A(AES_CORE_DATAPATH__abc_16259_n5461), .B(AES_CORE_DATAPATH__abc_16259_n5266_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n5462) );
  AND2X2 AND2X2_1521 ( .A(AES_CORE_DATAPATH__abc_16259_n5265_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__21_), .Y(AES_CORE_DATAPATH__abc_16259_n5463) );
  AND2X2 AND2X2_1522 ( .A(AES_CORE_DATAPATH__abc_16259_n5260_1_bF_buf1), .B(AES_CORE_DATAPATH_key_host_2__22_), .Y(AES_CORE_DATAPATH__abc_16259_n5466) );
  AND2X2 AND2X2_1523 ( .A(\bus_in[22] ), .B(key_en_2_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n5467) );
  AND2X2 AND2X2_1524 ( .A(AES_CORE_DATAPATH__abc_16259_n5465), .B(AES_CORE_DATAPATH__abc_16259_n5469), .Y(AES_CORE_DATAPATH__abc_16259_n5470) );
  AND2X2 AND2X2_1525 ( .A(AES_CORE_DATAPATH__abc_16259_n5470), .B(AES_CORE_DATAPATH__abc_16259_n5266_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n5471) );
  AND2X2 AND2X2_1526 ( .A(AES_CORE_DATAPATH__abc_16259_n5265_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__22_), .Y(AES_CORE_DATAPATH__abc_16259_n5472) );
  AND2X2 AND2X2_1527 ( .A(AES_CORE_DATAPATH__abc_16259_n5260_1_bF_buf0), .B(AES_CORE_DATAPATH_key_host_2__23_), .Y(AES_CORE_DATAPATH__abc_16259_n5475) );
  AND2X2 AND2X2_1528 ( .A(\bus_in[23] ), .B(key_en_2_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n5476) );
  AND2X2 AND2X2_1529 ( .A(AES_CORE_DATAPATH__abc_16259_n5474), .B(AES_CORE_DATAPATH__abc_16259_n5478), .Y(AES_CORE_DATAPATH__abc_16259_n5479) );
  AND2X2 AND2X2_153 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf5), .B(AES_CORE_DATAPATH_iv_1__9_), .Y(AES_CORE_DATAPATH__abc_16259_n2564_1) );
  AND2X2 AND2X2_1530 ( .A(AES_CORE_DATAPATH__abc_16259_n5479), .B(AES_CORE_DATAPATH__abc_16259_n5266_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n5480) );
  AND2X2 AND2X2_1531 ( .A(AES_CORE_DATAPATH__abc_16259_n5265_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__23_), .Y(AES_CORE_DATAPATH__abc_16259_n5481) );
  AND2X2 AND2X2_1532 ( .A(AES_CORE_DATAPATH__abc_16259_n5260_1_bF_buf4), .B(AES_CORE_DATAPATH_key_host_2__24_), .Y(AES_CORE_DATAPATH__abc_16259_n5484) );
  AND2X2 AND2X2_1533 ( .A(\bus_in[24] ), .B(key_en_2_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5485) );
  AND2X2 AND2X2_1534 ( .A(AES_CORE_DATAPATH__abc_16259_n5483), .B(AES_CORE_DATAPATH__abc_16259_n5487), .Y(AES_CORE_DATAPATH__abc_16259_n5488) );
  AND2X2 AND2X2_1535 ( .A(AES_CORE_DATAPATH__abc_16259_n5488), .B(AES_CORE_DATAPATH__abc_16259_n5266_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n5489) );
  AND2X2 AND2X2_1536 ( .A(AES_CORE_DATAPATH__abc_16259_n5265_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__24_), .Y(AES_CORE_DATAPATH__abc_16259_n5490) );
  AND2X2 AND2X2_1537 ( .A(AES_CORE_DATAPATH__abc_16259_n5260_1_bF_buf3), .B(AES_CORE_DATAPATH_key_host_2__25_), .Y(AES_CORE_DATAPATH__abc_16259_n5493) );
  AND2X2 AND2X2_1538 ( .A(\bus_in[25] ), .B(key_en_2_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n5494) );
  AND2X2 AND2X2_1539 ( .A(AES_CORE_DATAPATH__abc_16259_n5492), .B(AES_CORE_DATAPATH__abc_16259_n5496), .Y(AES_CORE_DATAPATH__abc_16259_n5497) );
  AND2X2 AND2X2_154 ( .A(AES_CORE_DATAPATH__abc_16259_n2567), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n2568_1) );
  AND2X2 AND2X2_1540 ( .A(AES_CORE_DATAPATH__abc_16259_n5497), .B(AES_CORE_DATAPATH__abc_16259_n5266_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5498) );
  AND2X2 AND2X2_1541 ( .A(AES_CORE_DATAPATH__abc_16259_n5265_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__25_), .Y(AES_CORE_DATAPATH__abc_16259_n5499) );
  AND2X2 AND2X2_1542 ( .A(AES_CORE_DATAPATH__abc_16259_n5260_1_bF_buf2), .B(AES_CORE_DATAPATH_key_host_2__26_), .Y(AES_CORE_DATAPATH__abc_16259_n5502) );
  AND2X2 AND2X2_1543 ( .A(\bus_in[26] ), .B(key_en_2_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n5503) );
  AND2X2 AND2X2_1544 ( .A(AES_CORE_DATAPATH__abc_16259_n5501), .B(AES_CORE_DATAPATH__abc_16259_n5505), .Y(AES_CORE_DATAPATH__abc_16259_n5506) );
  AND2X2 AND2X2_1545 ( .A(AES_CORE_DATAPATH__abc_16259_n5506), .B(AES_CORE_DATAPATH__abc_16259_n5266_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n5507) );
  AND2X2 AND2X2_1546 ( .A(AES_CORE_DATAPATH__abc_16259_n5265_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__26_), .Y(AES_CORE_DATAPATH__abc_16259_n5508) );
  AND2X2 AND2X2_1547 ( .A(AES_CORE_DATAPATH__abc_16259_n5260_1_bF_buf1), .B(AES_CORE_DATAPATH_key_host_2__27_), .Y(AES_CORE_DATAPATH__abc_16259_n5511) );
  AND2X2 AND2X2_1548 ( .A(\bus_in[27] ), .B(key_en_2_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n5512) );
  AND2X2 AND2X2_1549 ( .A(AES_CORE_DATAPATH__abc_16259_n5510), .B(AES_CORE_DATAPATH__abc_16259_n5514), .Y(AES_CORE_DATAPATH__abc_16259_n5515) );
  AND2X2 AND2X2_155 ( .A(AES_CORE_DATAPATH__abc_16259_n2566_1), .B(AES_CORE_DATAPATH__abc_16259_n2568_1), .Y(AES_CORE_DATAPATH__abc_16259_n2569_1) );
  AND2X2 AND2X2_1550 ( .A(AES_CORE_DATAPATH__abc_16259_n5515), .B(AES_CORE_DATAPATH__abc_16259_n5266_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n5516) );
  AND2X2 AND2X2_1551 ( .A(AES_CORE_DATAPATH__abc_16259_n5265_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__27_), .Y(AES_CORE_DATAPATH__abc_16259_n5517) );
  AND2X2 AND2X2_1552 ( .A(AES_CORE_DATAPATH__abc_16259_n5260_1_bF_buf0), .B(AES_CORE_DATAPATH_key_host_2__28_), .Y(AES_CORE_DATAPATH__abc_16259_n5520) );
  AND2X2 AND2X2_1553 ( .A(\bus_in[28] ), .B(key_en_2_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n5521) );
  AND2X2 AND2X2_1554 ( .A(AES_CORE_DATAPATH__abc_16259_n5519), .B(AES_CORE_DATAPATH__abc_16259_n5523), .Y(AES_CORE_DATAPATH__abc_16259_n5524) );
  AND2X2 AND2X2_1555 ( .A(AES_CORE_DATAPATH__abc_16259_n5524), .B(AES_CORE_DATAPATH__abc_16259_n5266_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n5525) );
  AND2X2 AND2X2_1556 ( .A(AES_CORE_DATAPATH__abc_16259_n5265_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__28_), .Y(AES_CORE_DATAPATH__abc_16259_n5526) );
  AND2X2 AND2X2_1557 ( .A(AES_CORE_DATAPATH__abc_16259_n5260_1_bF_buf4), .B(AES_CORE_DATAPATH_key_host_2__29_), .Y(AES_CORE_DATAPATH__abc_16259_n5529) );
  AND2X2 AND2X2_1558 ( .A(\bus_in[29] ), .B(key_en_2_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5530) );
  AND2X2 AND2X2_1559 ( .A(AES_CORE_DATAPATH__abc_16259_n5528), .B(AES_CORE_DATAPATH__abc_16259_n5532), .Y(AES_CORE_DATAPATH__abc_16259_n5533) );
  AND2X2 AND2X2_156 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf5), .B(AES_CORE_DATAPATH_iv_3__9_), .Y(AES_CORE_DATAPATH__abc_16259_n2570) );
  AND2X2 AND2X2_1560 ( .A(AES_CORE_DATAPATH__abc_16259_n5533), .B(AES_CORE_DATAPATH__abc_16259_n5266_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n5534) );
  AND2X2 AND2X2_1561 ( .A(AES_CORE_DATAPATH__abc_16259_n5265_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__29_), .Y(AES_CORE_DATAPATH__abc_16259_n5535) );
  AND2X2 AND2X2_1562 ( .A(AES_CORE_DATAPATH__abc_16259_n5260_1_bF_buf3), .B(AES_CORE_DATAPATH_key_host_2__30_), .Y(AES_CORE_DATAPATH__abc_16259_n5538) );
  AND2X2 AND2X2_1563 ( .A(\bus_in[30] ), .B(key_en_2_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n5539) );
  AND2X2 AND2X2_1564 ( .A(AES_CORE_DATAPATH__abc_16259_n5537), .B(AES_CORE_DATAPATH__abc_16259_n5541), .Y(AES_CORE_DATAPATH__abc_16259_n5542) );
  AND2X2 AND2X2_1565 ( .A(AES_CORE_DATAPATH__abc_16259_n5542), .B(AES_CORE_DATAPATH__abc_16259_n5266_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5543) );
  AND2X2 AND2X2_1566 ( .A(AES_CORE_DATAPATH__abc_16259_n5265_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__30_), .Y(AES_CORE_DATAPATH__abc_16259_n5544) );
  AND2X2 AND2X2_1567 ( .A(AES_CORE_DATAPATH__abc_16259_n5260_1_bF_buf2), .B(AES_CORE_DATAPATH_key_host_2__31_), .Y(AES_CORE_DATAPATH__abc_16259_n5546) );
  AND2X2 AND2X2_1568 ( .A(\bus_in[31] ), .B(key_en_2_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n5547) );
  AND2X2 AND2X2_1569 ( .A(AES_CORE_DATAPATH__abc_16259_n5550), .B(AES_CORE_DATAPATH__abc_16259_n5549), .Y(AES_CORE_DATAPATH__abc_16259_n5551) );
  AND2X2 AND2X2_157 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf5), .B(AES_CORE_DATAPATH_iv_0__10_), .Y(AES_CORE_DATAPATH__abc_16259_n2572) );
  AND2X2 AND2X2_1570 ( .A(AES_CORE_DATAPATH__abc_16259_n5551), .B(AES_CORE_DATAPATH__abc_16259_n5266_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n5552) );
  AND2X2 AND2X2_1571 ( .A(AES_CORE_DATAPATH__abc_16259_n5265_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__31_), .Y(AES_CORE_DATAPATH__abc_16259_n5553) );
  AND2X2 AND2X2_1572 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__0_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n5555) );
  AND2X2 AND2X2_1573 ( .A(AES_CORE_DATAPATH__abc_16259_n5270_1), .B(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n5556) );
  AND2X2 AND2X2_1574 ( .A(AES_CORE_DATAPATH__abc_16259_n5559), .B(AES_CORE_DATAPATH__abc_16259_n5558), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__1_) );
  AND2X2 AND2X2_1575 ( .A(AES_CORE_DATAPATH__abc_16259_n5562), .B(AES_CORE_DATAPATH__abc_16259_n5561), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__2_) );
  AND2X2 AND2X2_1576 ( .A(AES_CORE_DATAPATH__abc_16259_n5565), .B(AES_CORE_DATAPATH__abc_16259_n5564), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__3_) );
  AND2X2 AND2X2_1577 ( .A(AES_CORE_DATAPATH__abc_16259_n5568), .B(AES_CORE_DATAPATH__abc_16259_n5567), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__4_) );
  AND2X2 AND2X2_1578 ( .A(AES_CORE_DATAPATH__abc_16259_n5571), .B(AES_CORE_DATAPATH__abc_16259_n5570), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__5_) );
  AND2X2 AND2X2_1579 ( .A(AES_CORE_DATAPATH__abc_16259_n5574), .B(AES_CORE_DATAPATH__abc_16259_n5573), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__6_) );
  AND2X2 AND2X2_158 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf4), .B(AES_CORE_DATAPATH_iv_1__10_), .Y(AES_CORE_DATAPATH__abc_16259_n2573_1) );
  AND2X2 AND2X2_1580 ( .A(AES_CORE_DATAPATH__abc_16259_n5577), .B(AES_CORE_DATAPATH__abc_16259_n5576), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__7_) );
  AND2X2 AND2X2_1581 ( .A(AES_CORE_DATAPATH__abc_16259_n5580), .B(AES_CORE_DATAPATH__abc_16259_n5579), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__8_) );
  AND2X2 AND2X2_1582 ( .A(AES_CORE_DATAPATH__abc_16259_n5583), .B(AES_CORE_DATAPATH__abc_16259_n5582), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__9_) );
  AND2X2 AND2X2_1583 ( .A(AES_CORE_DATAPATH__abc_16259_n5586), .B(AES_CORE_DATAPATH__abc_16259_n5585), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__10_) );
  AND2X2 AND2X2_1584 ( .A(AES_CORE_DATAPATH__abc_16259_n5589), .B(AES_CORE_DATAPATH__abc_16259_n5588), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__11_) );
  AND2X2 AND2X2_1585 ( .A(AES_CORE_DATAPATH__abc_16259_n5592), .B(AES_CORE_DATAPATH__abc_16259_n5591), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__12_) );
  AND2X2 AND2X2_1586 ( .A(AES_CORE_DATAPATH__abc_16259_n5595), .B(AES_CORE_DATAPATH__abc_16259_n5594), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__13_) );
  AND2X2 AND2X2_1587 ( .A(AES_CORE_DATAPATH__abc_16259_n5598), .B(AES_CORE_DATAPATH__abc_16259_n5597), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__14_) );
  AND2X2 AND2X2_1588 ( .A(AES_CORE_DATAPATH__abc_16259_n5601), .B(AES_CORE_DATAPATH__abc_16259_n5600), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__15_) );
  AND2X2 AND2X2_1589 ( .A(AES_CORE_DATAPATH__abc_16259_n5604), .B(AES_CORE_DATAPATH__abc_16259_n5603), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__16_) );
  AND2X2 AND2X2_159 ( .A(AES_CORE_DATAPATH__abc_16259_n2576_1), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n2577) );
  AND2X2 AND2X2_1590 ( .A(AES_CORE_DATAPATH__abc_16259_n5607), .B(AES_CORE_DATAPATH__abc_16259_n5606), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__17_) );
  AND2X2 AND2X2_1591 ( .A(AES_CORE_DATAPATH__abc_16259_n5610), .B(AES_CORE_DATAPATH__abc_16259_n5609), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__18_) );
  AND2X2 AND2X2_1592 ( .A(AES_CORE_DATAPATH__abc_16259_n5613), .B(AES_CORE_DATAPATH__abc_16259_n5612), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__19_) );
  AND2X2 AND2X2_1593 ( .A(AES_CORE_DATAPATH__abc_16259_n5616), .B(AES_CORE_DATAPATH__abc_16259_n5615), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__20_) );
  AND2X2 AND2X2_1594 ( .A(AES_CORE_DATAPATH__abc_16259_n5619), .B(AES_CORE_DATAPATH__abc_16259_n5618), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__21_) );
  AND2X2 AND2X2_1595 ( .A(AES_CORE_DATAPATH__abc_16259_n5622), .B(AES_CORE_DATAPATH__abc_16259_n5621), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__22_) );
  AND2X2 AND2X2_1596 ( .A(AES_CORE_DATAPATH__abc_16259_n5625), .B(AES_CORE_DATAPATH__abc_16259_n5624), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__23_) );
  AND2X2 AND2X2_1597 ( .A(AES_CORE_DATAPATH__abc_16259_n5628), .B(AES_CORE_DATAPATH__abc_16259_n5627), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__24_) );
  AND2X2 AND2X2_1598 ( .A(AES_CORE_DATAPATH__abc_16259_n5631), .B(AES_CORE_DATAPATH__abc_16259_n5630), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__25_) );
  AND2X2 AND2X2_1599 ( .A(AES_CORE_DATAPATH__abc_16259_n5634), .B(AES_CORE_DATAPATH__abc_16259_n5633), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__26_) );
  AND2X2 AND2X2_16 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n90), .B(AES_CORE_CONTROL_UNIT__abc_15841_n77), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n91) );
  AND2X2 AND2X2_160 ( .A(AES_CORE_DATAPATH__abc_16259_n2575), .B(AES_CORE_DATAPATH__abc_16259_n2577), .Y(AES_CORE_DATAPATH__abc_16259_n2578_1) );
  AND2X2 AND2X2_1600 ( .A(AES_CORE_DATAPATH__abc_16259_n5637), .B(AES_CORE_DATAPATH__abc_16259_n5636), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__27_) );
  AND2X2 AND2X2_1601 ( .A(AES_CORE_DATAPATH__abc_16259_n5640), .B(AES_CORE_DATAPATH__abc_16259_n5639), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__28_) );
  AND2X2 AND2X2_1602 ( .A(AES_CORE_DATAPATH__abc_16259_n5643), .B(AES_CORE_DATAPATH__abc_16259_n5642), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__29_) );
  AND2X2 AND2X2_1603 ( .A(AES_CORE_DATAPATH__abc_16259_n5646), .B(AES_CORE_DATAPATH__abc_16259_n5645), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__30_) );
  AND2X2 AND2X2_1604 ( .A(AES_CORE_DATAPATH__abc_16259_n5648), .B(AES_CORE_DATAPATH__abc_16259_n5649), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__31_) );
  AND2X2 AND2X2_1605 ( .A(AES_CORE_CONTROL_UNIT_bypass_key_en), .B(AES_CORE_CONTROL_UNIT_key_en_3_), .Y(AES_CORE_DATAPATH__abc_16259_n5651) );
  AND2X2 AND2X2_1606 ( .A(AES_CORE_DATAPATH__abc_16259_n4469_1), .B(AES_CORE_DATAPATH__abc_16259_n5653_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5654) );
  AND2X2 AND2X2_1607 ( .A(AES_CORE_DATAPATH__abc_16259_n2806_1), .B(AES_CORE_DATAPATH_key_en_pp1_3_), .Y(AES_CORE_DATAPATH__abc_16259_n5655) );
  AND2X2 AND2X2_1608 ( .A(AES_CORE_DATAPATH__abc_16259_n5656), .B(AES_CORE_DATAPATH__abc_16259_n5654), .Y(AES_CORE_DATAPATH__abc_16259_n5657) );
  AND2X2 AND2X2_1609 ( .A(AES_CORE_DATAPATH__abc_16259_n5657), .B(AES_CORE_DATAPATH__abc_16259_n5652), .Y(AES_CORE_DATAPATH__abc_16259_n5658) );
  AND2X2 AND2X2_161 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf4), .B(AES_CORE_DATAPATH_iv_3__10_), .Y(AES_CORE_DATAPATH__abc_16259_n2579_1) );
  AND2X2 AND2X2_1610 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_0_), .Y(AES_CORE_DATAPATH__abc_16259_n5660) );
  AND2X2 AND2X2_1611 ( .A(\bus_in[0] ), .B(key_en_3_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n5661) );
  AND2X2 AND2X2_1612 ( .A(AES_CORE_DATAPATH__abc_16259_n5653_bF_buf3), .B(AES_CORE_DATAPATH_key_host_3__0_), .Y(AES_CORE_DATAPATH__abc_16259_n5662) );
  AND2X2 AND2X2_1613 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n5663), .Y(AES_CORE_DATAPATH__abc_16259_n5664) );
  AND2X2 AND2X2_1614 ( .A(AES_CORE_DATAPATH__abc_16259_n5665), .B(AES_CORE_DATAPATH__abc_16259_n5659_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5666) );
  AND2X2 AND2X2_1615 ( .A(AES_CORE_DATAPATH__abc_16259_n5658_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__0_), .Y(AES_CORE_DATAPATH__abc_16259_n5667) );
  AND2X2 AND2X2_1616 ( .A(AES_CORE_DATAPATH__abc_16259_n5653_bF_buf2), .B(AES_CORE_DATAPATH_key_host_3__1_), .Y(AES_CORE_DATAPATH__abc_16259_n5670) );
  AND2X2 AND2X2_1617 ( .A(\bus_in[1] ), .B(key_en_3_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n5671) );
  AND2X2 AND2X2_1618 ( .A(AES_CORE_DATAPATH__abc_16259_n5669), .B(AES_CORE_DATAPATH__abc_16259_n5673), .Y(AES_CORE_DATAPATH__abc_16259_n5674) );
  AND2X2 AND2X2_1619 ( .A(AES_CORE_DATAPATH__abc_16259_n5674), .B(AES_CORE_DATAPATH__abc_16259_n5659_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n5675) );
  AND2X2 AND2X2_162 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf4), .B(AES_CORE_DATAPATH_iv_0__11_), .Y(AES_CORE_DATAPATH__abc_16259_n2581_1) );
  AND2X2 AND2X2_1620 ( .A(AES_CORE_DATAPATH__abc_16259_n5658_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__1_), .Y(AES_CORE_DATAPATH__abc_16259_n5676) );
  AND2X2 AND2X2_1621 ( .A(AES_CORE_DATAPATH__abc_16259_n5653_bF_buf1), .B(AES_CORE_DATAPATH_key_host_3__2_), .Y(AES_CORE_DATAPATH__abc_16259_n5679) );
  AND2X2 AND2X2_1622 ( .A(\bus_in[2] ), .B(key_en_3_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n5680) );
  AND2X2 AND2X2_1623 ( .A(AES_CORE_DATAPATH__abc_16259_n5678), .B(AES_CORE_DATAPATH__abc_16259_n5682), .Y(AES_CORE_DATAPATH__abc_16259_n5683) );
  AND2X2 AND2X2_1624 ( .A(AES_CORE_DATAPATH__abc_16259_n5683), .B(AES_CORE_DATAPATH__abc_16259_n5659_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n5684) );
  AND2X2 AND2X2_1625 ( .A(AES_CORE_DATAPATH__abc_16259_n5658_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__2_), .Y(AES_CORE_DATAPATH__abc_16259_n5685) );
  AND2X2 AND2X2_1626 ( .A(AES_CORE_DATAPATH__abc_16259_n5653_bF_buf0), .B(AES_CORE_DATAPATH_key_host_3__3_), .Y(AES_CORE_DATAPATH__abc_16259_n5688) );
  AND2X2 AND2X2_1627 ( .A(\bus_in[3] ), .B(key_en_3_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n5689) );
  AND2X2 AND2X2_1628 ( .A(AES_CORE_DATAPATH__abc_16259_n5687), .B(AES_CORE_DATAPATH__abc_16259_n5691), .Y(AES_CORE_DATAPATH__abc_16259_n5692) );
  AND2X2 AND2X2_1629 ( .A(AES_CORE_DATAPATH__abc_16259_n5692), .B(AES_CORE_DATAPATH__abc_16259_n5659_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n5693) );
  AND2X2 AND2X2_163 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf3), .B(AES_CORE_DATAPATH_iv_1__11_), .Y(AES_CORE_DATAPATH__abc_16259_n2582) );
  AND2X2 AND2X2_1630 ( .A(AES_CORE_DATAPATH__abc_16259_n5658_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__3_), .Y(AES_CORE_DATAPATH__abc_16259_n5694) );
  AND2X2 AND2X2_1631 ( .A(AES_CORE_DATAPATH__abc_16259_n5653_bF_buf4), .B(AES_CORE_DATAPATH_key_host_3__4_), .Y(AES_CORE_DATAPATH__abc_16259_n5697) );
  AND2X2 AND2X2_1632 ( .A(\bus_in[4] ), .B(key_en_3_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5698) );
  AND2X2 AND2X2_1633 ( .A(AES_CORE_DATAPATH__abc_16259_n5696), .B(AES_CORE_DATAPATH__abc_16259_n5700), .Y(AES_CORE_DATAPATH__abc_16259_n5701) );
  AND2X2 AND2X2_1634 ( .A(AES_CORE_DATAPATH__abc_16259_n5701), .B(AES_CORE_DATAPATH__abc_16259_n5659_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n5702) );
  AND2X2 AND2X2_1635 ( .A(AES_CORE_DATAPATH__abc_16259_n5658_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__4_), .Y(AES_CORE_DATAPATH__abc_16259_n5703) );
  AND2X2 AND2X2_1636 ( .A(AES_CORE_DATAPATH__abc_16259_n5653_bF_buf3), .B(AES_CORE_DATAPATH_key_host_3__5_), .Y(AES_CORE_DATAPATH__abc_16259_n5706) );
  AND2X2 AND2X2_1637 ( .A(\bus_in[5] ), .B(key_en_3_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n5707) );
  AND2X2 AND2X2_1638 ( .A(AES_CORE_DATAPATH__abc_16259_n5705), .B(AES_CORE_DATAPATH__abc_16259_n5709), .Y(AES_CORE_DATAPATH__abc_16259_n5710) );
  AND2X2 AND2X2_1639 ( .A(AES_CORE_DATAPATH__abc_16259_n5710), .B(AES_CORE_DATAPATH__abc_16259_n5659_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5711) );
  AND2X2 AND2X2_164 ( .A(AES_CORE_DATAPATH__abc_16259_n2585), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n2586_1) );
  AND2X2 AND2X2_1640 ( .A(AES_CORE_DATAPATH__abc_16259_n5658_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__5_), .Y(AES_CORE_DATAPATH__abc_16259_n5712) );
  AND2X2 AND2X2_1641 ( .A(AES_CORE_DATAPATH__abc_16259_n5653_bF_buf2), .B(AES_CORE_DATAPATH_key_host_3__6_), .Y(AES_CORE_DATAPATH__abc_16259_n5715) );
  AND2X2 AND2X2_1642 ( .A(\bus_in[6] ), .B(key_en_3_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n5716) );
  AND2X2 AND2X2_1643 ( .A(AES_CORE_DATAPATH__abc_16259_n5714), .B(AES_CORE_DATAPATH__abc_16259_n5718), .Y(AES_CORE_DATAPATH__abc_16259_n5719) );
  AND2X2 AND2X2_1644 ( .A(AES_CORE_DATAPATH__abc_16259_n5720), .B(AES_CORE_DATAPATH__abc_16259_n5721), .Y(AES_CORE_DATAPATH__0key_3__31_0__6_) );
  AND2X2 AND2X2_1645 ( .A(AES_CORE_DATAPATH__abc_16259_n5653_bF_buf1), .B(AES_CORE_DATAPATH_key_host_3__7_), .Y(AES_CORE_DATAPATH__abc_16259_n5724) );
  AND2X2 AND2X2_1646 ( .A(\bus_in[7] ), .B(key_en_3_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n5725) );
  AND2X2 AND2X2_1647 ( .A(AES_CORE_DATAPATH__abc_16259_n5723), .B(AES_CORE_DATAPATH__abc_16259_n5727), .Y(AES_CORE_DATAPATH__abc_16259_n5728) );
  AND2X2 AND2X2_1648 ( .A(AES_CORE_DATAPATH__abc_16259_n5728), .B(AES_CORE_DATAPATH__abc_16259_n5659_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n5729) );
  AND2X2 AND2X2_1649 ( .A(AES_CORE_DATAPATH__abc_16259_n5658_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__7_), .Y(AES_CORE_DATAPATH__abc_16259_n5730) );
  AND2X2 AND2X2_165 ( .A(AES_CORE_DATAPATH__abc_16259_n2584_1), .B(AES_CORE_DATAPATH__abc_16259_n2586_1), .Y(AES_CORE_DATAPATH__abc_16259_n2587) );
  AND2X2 AND2X2_1650 ( .A(AES_CORE_DATAPATH__abc_16259_n5653_bF_buf0), .B(AES_CORE_DATAPATH_key_host_3__8_), .Y(AES_CORE_DATAPATH__abc_16259_n5733) );
  AND2X2 AND2X2_1651 ( .A(\bus_in[8] ), .B(key_en_3_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n5734) );
  AND2X2 AND2X2_1652 ( .A(AES_CORE_DATAPATH__abc_16259_n5732), .B(AES_CORE_DATAPATH__abc_16259_n5736), .Y(AES_CORE_DATAPATH__abc_16259_n5737) );
  AND2X2 AND2X2_1653 ( .A(AES_CORE_DATAPATH__abc_16259_n5738), .B(AES_CORE_DATAPATH__abc_16259_n5739), .Y(AES_CORE_DATAPATH__0key_3__31_0__8_) );
  AND2X2 AND2X2_1654 ( .A(AES_CORE_DATAPATH__abc_16259_n5653_bF_buf4), .B(AES_CORE_DATAPATH_key_host_3__9_), .Y(AES_CORE_DATAPATH__abc_16259_n5742) );
  AND2X2 AND2X2_1655 ( .A(\bus_in[9] ), .B(key_en_3_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5743) );
  AND2X2 AND2X2_1656 ( .A(AES_CORE_DATAPATH__abc_16259_n5741), .B(AES_CORE_DATAPATH__abc_16259_n5745), .Y(AES_CORE_DATAPATH__abc_16259_n5746) );
  AND2X2 AND2X2_1657 ( .A(AES_CORE_DATAPATH__abc_16259_n5746), .B(AES_CORE_DATAPATH__abc_16259_n5659_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n5747) );
  AND2X2 AND2X2_1658 ( .A(AES_CORE_DATAPATH__abc_16259_n5658_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__9_), .Y(AES_CORE_DATAPATH__abc_16259_n5748) );
  AND2X2 AND2X2_1659 ( .A(AES_CORE_DATAPATH__abc_16259_n5653_bF_buf3), .B(AES_CORE_DATAPATH_key_host_3__10_), .Y(AES_CORE_DATAPATH__abc_16259_n5751) );
  AND2X2 AND2X2_166 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf3), .B(AES_CORE_DATAPATH_iv_3__11_), .Y(AES_CORE_DATAPATH__abc_16259_n2588_1) );
  AND2X2 AND2X2_1660 ( .A(\bus_in[10] ), .B(key_en_3_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n5752) );
  AND2X2 AND2X2_1661 ( .A(AES_CORE_DATAPATH__abc_16259_n5750), .B(AES_CORE_DATAPATH__abc_16259_n5754), .Y(AES_CORE_DATAPATH__abc_16259_n5755) );
  AND2X2 AND2X2_1662 ( .A(AES_CORE_DATAPATH__abc_16259_n5755), .B(AES_CORE_DATAPATH__abc_16259_n5659_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5756) );
  AND2X2 AND2X2_1663 ( .A(AES_CORE_DATAPATH__abc_16259_n5658_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__10_), .Y(AES_CORE_DATAPATH__abc_16259_n5757) );
  AND2X2 AND2X2_1664 ( .A(AES_CORE_DATAPATH__abc_16259_n5653_bF_buf2), .B(AES_CORE_DATAPATH_key_host_3__11_), .Y(AES_CORE_DATAPATH__abc_16259_n5760) );
  AND2X2 AND2X2_1665 ( .A(\bus_in[11] ), .B(key_en_3_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n5761) );
  AND2X2 AND2X2_1666 ( .A(AES_CORE_DATAPATH__abc_16259_n5759), .B(AES_CORE_DATAPATH__abc_16259_n5763), .Y(AES_CORE_DATAPATH__abc_16259_n5764) );
  AND2X2 AND2X2_1667 ( .A(AES_CORE_DATAPATH__abc_16259_n5764), .B(AES_CORE_DATAPATH__abc_16259_n5659_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n5765) );
  AND2X2 AND2X2_1668 ( .A(AES_CORE_DATAPATH__abc_16259_n5658_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__11_), .Y(AES_CORE_DATAPATH__abc_16259_n5766) );
  AND2X2 AND2X2_1669 ( .A(AES_CORE_DATAPATH__abc_16259_n5653_bF_buf1), .B(AES_CORE_DATAPATH_key_host_3__12_), .Y(AES_CORE_DATAPATH__abc_16259_n5769) );
  AND2X2 AND2X2_167 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf3), .B(AES_CORE_DATAPATH_iv_0__12_), .Y(AES_CORE_DATAPATH__abc_16259_n2590) );
  AND2X2 AND2X2_1670 ( .A(\bus_in[12] ), .B(key_en_3_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n5770) );
  AND2X2 AND2X2_1671 ( .A(AES_CORE_DATAPATH__abc_16259_n5768), .B(AES_CORE_DATAPATH__abc_16259_n5772), .Y(AES_CORE_DATAPATH__abc_16259_n5773) );
  AND2X2 AND2X2_1672 ( .A(AES_CORE_DATAPATH__abc_16259_n5774), .B(AES_CORE_DATAPATH__abc_16259_n5775), .Y(AES_CORE_DATAPATH__0key_3__31_0__12_) );
  AND2X2 AND2X2_1673 ( .A(AES_CORE_DATAPATH__abc_16259_n5653_bF_buf0), .B(AES_CORE_DATAPATH_key_host_3__13_), .Y(AES_CORE_DATAPATH__abc_16259_n5778) );
  AND2X2 AND2X2_1674 ( .A(\bus_in[13] ), .B(key_en_3_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n5779) );
  AND2X2 AND2X2_1675 ( .A(AES_CORE_DATAPATH__abc_16259_n5777), .B(AES_CORE_DATAPATH__abc_16259_n5781), .Y(AES_CORE_DATAPATH__abc_16259_n5782) );
  AND2X2 AND2X2_1676 ( .A(AES_CORE_DATAPATH__abc_16259_n5782), .B(AES_CORE_DATAPATH__abc_16259_n5659_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n5783) );
  AND2X2 AND2X2_1677 ( .A(AES_CORE_DATAPATH__abc_16259_n5658_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__13_), .Y(AES_CORE_DATAPATH__abc_16259_n5784) );
  AND2X2 AND2X2_1678 ( .A(AES_CORE_DATAPATH__abc_16259_n5653_bF_buf4), .B(AES_CORE_DATAPATH_key_host_3__14_), .Y(AES_CORE_DATAPATH__abc_16259_n5787) );
  AND2X2 AND2X2_1679 ( .A(\bus_in[14] ), .B(key_en_3_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5788) );
  AND2X2 AND2X2_168 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf2), .B(AES_CORE_DATAPATH_iv_1__12_), .Y(AES_CORE_DATAPATH__abc_16259_n2591_1) );
  AND2X2 AND2X2_1680 ( .A(AES_CORE_DATAPATH__abc_16259_n5786), .B(AES_CORE_DATAPATH__abc_16259_n5790), .Y(AES_CORE_DATAPATH__abc_16259_n5791) );
  AND2X2 AND2X2_1681 ( .A(AES_CORE_DATAPATH__abc_16259_n5792), .B(AES_CORE_DATAPATH__abc_16259_n5793), .Y(AES_CORE_DATAPATH__0key_3__31_0__14_) );
  AND2X2 AND2X2_1682 ( .A(AES_CORE_DATAPATH__abc_16259_n5653_bF_buf3), .B(AES_CORE_DATAPATH_key_host_3__15_), .Y(AES_CORE_DATAPATH__abc_16259_n5796) );
  AND2X2 AND2X2_1683 ( .A(\bus_in[15] ), .B(key_en_3_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n5797) );
  AND2X2 AND2X2_1684 ( .A(AES_CORE_DATAPATH__abc_16259_n5795), .B(AES_CORE_DATAPATH__abc_16259_n5799), .Y(AES_CORE_DATAPATH__abc_16259_n5800) );
  AND2X2 AND2X2_1685 ( .A(AES_CORE_DATAPATH__abc_16259_n5800), .B(AES_CORE_DATAPATH__abc_16259_n5659_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5801) );
  AND2X2 AND2X2_1686 ( .A(AES_CORE_DATAPATH__abc_16259_n5658_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__15_), .Y(AES_CORE_DATAPATH__abc_16259_n5802) );
  AND2X2 AND2X2_1687 ( .A(AES_CORE_DATAPATH__abc_16259_n5653_bF_buf2), .B(AES_CORE_DATAPATH_key_host_3__16_), .Y(AES_CORE_DATAPATH__abc_16259_n5805) );
  AND2X2 AND2X2_1688 ( .A(\bus_in[16] ), .B(key_en_3_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n5806) );
  AND2X2 AND2X2_1689 ( .A(AES_CORE_DATAPATH__abc_16259_n5804), .B(AES_CORE_DATAPATH__abc_16259_n5808), .Y(AES_CORE_DATAPATH__abc_16259_n5809) );
  AND2X2 AND2X2_169 ( .A(AES_CORE_DATAPATH__abc_16259_n2594_1), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n2595) );
  AND2X2 AND2X2_1690 ( .A(AES_CORE_DATAPATH__abc_16259_n5810), .B(AES_CORE_DATAPATH__abc_16259_n5811), .Y(AES_CORE_DATAPATH__0key_3__31_0__16_) );
  AND2X2 AND2X2_1691 ( .A(AES_CORE_DATAPATH__abc_16259_n5653_bF_buf1), .B(AES_CORE_DATAPATH_key_host_3__17_), .Y(AES_CORE_DATAPATH__abc_16259_n5814) );
  AND2X2 AND2X2_1692 ( .A(\bus_in[17] ), .B(key_en_3_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n5815) );
  AND2X2 AND2X2_1693 ( .A(AES_CORE_DATAPATH__abc_16259_n5813), .B(AES_CORE_DATAPATH__abc_16259_n5817), .Y(AES_CORE_DATAPATH__abc_16259_n5818) );
  AND2X2 AND2X2_1694 ( .A(AES_CORE_DATAPATH__abc_16259_n5818), .B(AES_CORE_DATAPATH__abc_16259_n5659_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n5819) );
  AND2X2 AND2X2_1695 ( .A(AES_CORE_DATAPATH__abc_16259_n5658_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__17_), .Y(AES_CORE_DATAPATH__abc_16259_n5820) );
  AND2X2 AND2X2_1696 ( .A(AES_CORE_DATAPATH__abc_16259_n5653_bF_buf0), .B(AES_CORE_DATAPATH_key_host_3__18_), .Y(AES_CORE_DATAPATH__abc_16259_n5823) );
  AND2X2 AND2X2_1697 ( .A(\bus_in[18] ), .B(key_en_3_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n5824) );
  AND2X2 AND2X2_1698 ( .A(AES_CORE_DATAPATH__abc_16259_n5822), .B(AES_CORE_DATAPATH__abc_16259_n5826), .Y(AES_CORE_DATAPATH__abc_16259_n5827) );
  AND2X2 AND2X2_1699 ( .A(AES_CORE_DATAPATH__abc_16259_n5827), .B(AES_CORE_DATAPATH__abc_16259_n5659_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n5828) );
  AND2X2 AND2X2_17 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n92), .B(AES_CORE_CONTROL_UNIT_state_7_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n93_1) );
  AND2X2 AND2X2_170 ( .A(AES_CORE_DATAPATH__abc_16259_n2593_1), .B(AES_CORE_DATAPATH__abc_16259_n2595), .Y(AES_CORE_DATAPATH__abc_16259_n2596_1) );
  AND2X2 AND2X2_1700 ( .A(AES_CORE_DATAPATH__abc_16259_n5658_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__18_), .Y(AES_CORE_DATAPATH__abc_16259_n5829) );
  AND2X2 AND2X2_1701 ( .A(AES_CORE_DATAPATH__abc_16259_n5653_bF_buf4), .B(AES_CORE_DATAPATH_key_host_3__19_), .Y(AES_CORE_DATAPATH__abc_16259_n5832) );
  AND2X2 AND2X2_1702 ( .A(\bus_in[19] ), .B(key_en_3_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5833) );
  AND2X2 AND2X2_1703 ( .A(AES_CORE_DATAPATH__abc_16259_n5831), .B(AES_CORE_DATAPATH__abc_16259_n5835), .Y(AES_CORE_DATAPATH__abc_16259_n5836) );
  AND2X2 AND2X2_1704 ( .A(AES_CORE_DATAPATH__abc_16259_n5836), .B(AES_CORE_DATAPATH__abc_16259_n5659_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n5837) );
  AND2X2 AND2X2_1705 ( .A(AES_CORE_DATAPATH__abc_16259_n5658_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__19_), .Y(AES_CORE_DATAPATH__abc_16259_n5838) );
  AND2X2 AND2X2_1706 ( .A(AES_CORE_DATAPATH__abc_16259_n5653_bF_buf3), .B(AES_CORE_DATAPATH_key_host_3__20_), .Y(AES_CORE_DATAPATH__abc_16259_n5841) );
  AND2X2 AND2X2_1707 ( .A(\bus_in[20] ), .B(key_en_3_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n5842) );
  AND2X2 AND2X2_1708 ( .A(AES_CORE_DATAPATH__abc_16259_n5840), .B(AES_CORE_DATAPATH__abc_16259_n5844), .Y(AES_CORE_DATAPATH__abc_16259_n5845) );
  AND2X2 AND2X2_1709 ( .A(AES_CORE_DATAPATH__abc_16259_n5845), .B(AES_CORE_DATAPATH__abc_16259_n5659_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5846) );
  AND2X2 AND2X2_171 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf2), .B(AES_CORE_DATAPATH_iv_3__12_), .Y(AES_CORE_DATAPATH__abc_16259_n2597) );
  AND2X2 AND2X2_1710 ( .A(AES_CORE_DATAPATH__abc_16259_n5658_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__20_), .Y(AES_CORE_DATAPATH__abc_16259_n5847) );
  AND2X2 AND2X2_1711 ( .A(AES_CORE_DATAPATH__abc_16259_n5653_bF_buf2), .B(AES_CORE_DATAPATH_key_host_3__21_), .Y(AES_CORE_DATAPATH__abc_16259_n5850) );
  AND2X2 AND2X2_1712 ( .A(\bus_in[21] ), .B(key_en_3_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n5851) );
  AND2X2 AND2X2_1713 ( .A(AES_CORE_DATAPATH__abc_16259_n5849), .B(AES_CORE_DATAPATH__abc_16259_n5853), .Y(AES_CORE_DATAPATH__abc_16259_n5854) );
  AND2X2 AND2X2_1714 ( .A(AES_CORE_DATAPATH__abc_16259_n5855), .B(AES_CORE_DATAPATH__abc_16259_n5856), .Y(AES_CORE_DATAPATH__0key_3__31_0__21_) );
  AND2X2 AND2X2_1715 ( .A(AES_CORE_DATAPATH__abc_16259_n5653_bF_buf1), .B(AES_CORE_DATAPATH_key_host_3__22_), .Y(AES_CORE_DATAPATH__abc_16259_n5859) );
  AND2X2 AND2X2_1716 ( .A(\bus_in[22] ), .B(key_en_3_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n5860) );
  AND2X2 AND2X2_1717 ( .A(AES_CORE_DATAPATH__abc_16259_n5858), .B(AES_CORE_DATAPATH__abc_16259_n5862), .Y(AES_CORE_DATAPATH__abc_16259_n5863) );
  AND2X2 AND2X2_1718 ( .A(AES_CORE_DATAPATH__abc_16259_n5863), .B(AES_CORE_DATAPATH__abc_16259_n5659_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n5864) );
  AND2X2 AND2X2_1719 ( .A(AES_CORE_DATAPATH__abc_16259_n5658_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__22_), .Y(AES_CORE_DATAPATH__abc_16259_n5865) );
  AND2X2 AND2X2_172 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf2), .B(AES_CORE_DATAPATH_iv_0__13_), .Y(AES_CORE_DATAPATH__abc_16259_n2599_1) );
  AND2X2 AND2X2_1720 ( .A(AES_CORE_DATAPATH__abc_16259_n5653_bF_buf0), .B(AES_CORE_DATAPATH_key_host_3__23_), .Y(AES_CORE_DATAPATH__abc_16259_n5868) );
  AND2X2 AND2X2_1721 ( .A(\bus_in[23] ), .B(key_en_3_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n5869) );
  AND2X2 AND2X2_1722 ( .A(AES_CORE_DATAPATH__abc_16259_n5867), .B(AES_CORE_DATAPATH__abc_16259_n5871), .Y(AES_CORE_DATAPATH__abc_16259_n5872) );
  AND2X2 AND2X2_1723 ( .A(AES_CORE_DATAPATH__abc_16259_n5873), .B(AES_CORE_DATAPATH__abc_16259_n5874), .Y(AES_CORE_DATAPATH__0key_3__31_0__23_) );
  AND2X2 AND2X2_1724 ( .A(AES_CORE_DATAPATH__abc_16259_n5653_bF_buf4), .B(AES_CORE_DATAPATH_key_host_3__24_), .Y(AES_CORE_DATAPATH__abc_16259_n5877) );
  AND2X2 AND2X2_1725 ( .A(\bus_in[24] ), .B(key_en_3_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5878) );
  AND2X2 AND2X2_1726 ( .A(AES_CORE_DATAPATH__abc_16259_n5876), .B(AES_CORE_DATAPATH__abc_16259_n5880), .Y(AES_CORE_DATAPATH__abc_16259_n5881) );
  AND2X2 AND2X2_1727 ( .A(AES_CORE_DATAPATH__abc_16259_n5881), .B(AES_CORE_DATAPATH__abc_16259_n5659_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n5882) );
  AND2X2 AND2X2_1728 ( .A(AES_CORE_DATAPATH__abc_16259_n5658_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__24_), .Y(AES_CORE_DATAPATH__abc_16259_n5883) );
  AND2X2 AND2X2_1729 ( .A(AES_CORE_DATAPATH__abc_16259_n5653_bF_buf3), .B(AES_CORE_DATAPATH_key_host_3__25_), .Y(AES_CORE_DATAPATH__abc_16259_n5886) );
  AND2X2 AND2X2_173 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf1), .B(AES_CORE_DATAPATH_iv_1__13_), .Y(AES_CORE_DATAPATH__abc_16259_n2600) );
  AND2X2 AND2X2_1730 ( .A(\bus_in[25] ), .B(key_en_3_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n5887) );
  AND2X2 AND2X2_1731 ( .A(AES_CORE_DATAPATH__abc_16259_n5885), .B(AES_CORE_DATAPATH__abc_16259_n5889), .Y(AES_CORE_DATAPATH__abc_16259_n5890) );
  AND2X2 AND2X2_1732 ( .A(AES_CORE_DATAPATH__abc_16259_n5891), .B(AES_CORE_DATAPATH__abc_16259_n5892), .Y(AES_CORE_DATAPATH__0key_3__31_0__25_) );
  AND2X2 AND2X2_1733 ( .A(AES_CORE_DATAPATH__abc_16259_n5653_bF_buf2), .B(AES_CORE_DATAPATH_key_host_3__26_), .Y(AES_CORE_DATAPATH__abc_16259_n5895) );
  AND2X2 AND2X2_1734 ( .A(\bus_in[26] ), .B(key_en_3_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n5896) );
  AND2X2 AND2X2_1735 ( .A(AES_CORE_DATAPATH__abc_16259_n5894), .B(AES_CORE_DATAPATH__abc_16259_n5898), .Y(AES_CORE_DATAPATH__abc_16259_n5899) );
  AND2X2 AND2X2_1736 ( .A(AES_CORE_DATAPATH__abc_16259_n5899), .B(AES_CORE_DATAPATH__abc_16259_n5659_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n5900) );
  AND2X2 AND2X2_1737 ( .A(AES_CORE_DATAPATH__abc_16259_n5658_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__26_), .Y(AES_CORE_DATAPATH__abc_16259_n5901) );
  AND2X2 AND2X2_1738 ( .A(AES_CORE_DATAPATH__abc_16259_n5653_bF_buf1), .B(AES_CORE_DATAPATH_key_host_3__27_), .Y(AES_CORE_DATAPATH__abc_16259_n5904) );
  AND2X2 AND2X2_1739 ( .A(\bus_in[27] ), .B(key_en_3_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n5905) );
  AND2X2 AND2X2_174 ( .A(AES_CORE_DATAPATH__abc_16259_n2603_1), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n2604_1) );
  AND2X2 AND2X2_1740 ( .A(AES_CORE_DATAPATH__abc_16259_n5903), .B(AES_CORE_DATAPATH__abc_16259_n5907), .Y(AES_CORE_DATAPATH__abc_16259_n5908) );
  AND2X2 AND2X2_1741 ( .A(AES_CORE_DATAPATH__abc_16259_n5908), .B(AES_CORE_DATAPATH__abc_16259_n5659_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n5909) );
  AND2X2 AND2X2_1742 ( .A(AES_CORE_DATAPATH__abc_16259_n5658_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__27_), .Y(AES_CORE_DATAPATH__abc_16259_n5910) );
  AND2X2 AND2X2_1743 ( .A(AES_CORE_DATAPATH__abc_16259_n5653_bF_buf0), .B(AES_CORE_DATAPATH_key_host_3__28_), .Y(AES_CORE_DATAPATH__abc_16259_n5913) );
  AND2X2 AND2X2_1744 ( .A(\bus_in[28] ), .B(key_en_3_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n5914) );
  AND2X2 AND2X2_1745 ( .A(AES_CORE_DATAPATH__abc_16259_n5912), .B(AES_CORE_DATAPATH__abc_16259_n5916), .Y(AES_CORE_DATAPATH__abc_16259_n5917) );
  AND2X2 AND2X2_1746 ( .A(AES_CORE_DATAPATH__abc_16259_n5917), .B(AES_CORE_DATAPATH__abc_16259_n5659_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n5918) );
  AND2X2 AND2X2_1747 ( .A(AES_CORE_DATAPATH__abc_16259_n5658_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__28_), .Y(AES_CORE_DATAPATH__abc_16259_n5919) );
  AND2X2 AND2X2_1748 ( .A(AES_CORE_DATAPATH__abc_16259_n5653_bF_buf4), .B(AES_CORE_DATAPATH_key_host_3__29_), .Y(AES_CORE_DATAPATH__abc_16259_n5922) );
  AND2X2 AND2X2_1749 ( .A(\bus_in[29] ), .B(key_en_3_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5923) );
  AND2X2 AND2X2_175 ( .A(AES_CORE_DATAPATH__abc_16259_n2602), .B(AES_CORE_DATAPATH__abc_16259_n2604_1), .Y(AES_CORE_DATAPATH__abc_16259_n2605) );
  AND2X2 AND2X2_1750 ( .A(AES_CORE_DATAPATH__abc_16259_n5921), .B(AES_CORE_DATAPATH__abc_16259_n5925), .Y(AES_CORE_DATAPATH__abc_16259_n5926) );
  AND2X2 AND2X2_1751 ( .A(AES_CORE_DATAPATH__abc_16259_n5926), .B(AES_CORE_DATAPATH__abc_16259_n5659_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n5927) );
  AND2X2 AND2X2_1752 ( .A(AES_CORE_DATAPATH__abc_16259_n5658_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__29_), .Y(AES_CORE_DATAPATH__abc_16259_n5928) );
  AND2X2 AND2X2_1753 ( .A(AES_CORE_DATAPATH__abc_16259_n5653_bF_buf3), .B(AES_CORE_DATAPATH_key_host_3__30_), .Y(AES_CORE_DATAPATH__abc_16259_n5931) );
  AND2X2 AND2X2_1754 ( .A(\bus_in[30] ), .B(key_en_3_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n5932) );
  AND2X2 AND2X2_1755 ( .A(AES_CORE_DATAPATH__abc_16259_n5930), .B(AES_CORE_DATAPATH__abc_16259_n5934), .Y(AES_CORE_DATAPATH__abc_16259_n5935) );
  AND2X2 AND2X2_1756 ( .A(AES_CORE_DATAPATH__abc_16259_n5935), .B(AES_CORE_DATAPATH__abc_16259_n5659_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5936) );
  AND2X2 AND2X2_1757 ( .A(AES_CORE_DATAPATH__abc_16259_n5658_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__30_), .Y(AES_CORE_DATAPATH__abc_16259_n5937) );
  AND2X2 AND2X2_1758 ( .A(AES_CORE_DATAPATH__abc_16259_n5653_bF_buf2), .B(AES_CORE_DATAPATH_key_host_3__31_), .Y(AES_CORE_DATAPATH__abc_16259_n5939) );
  AND2X2 AND2X2_1759 ( .A(\bus_in[31] ), .B(key_en_3_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n5940) );
  AND2X2 AND2X2_176 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf1), .B(AES_CORE_DATAPATH_iv_3__13_), .Y(AES_CORE_DATAPATH__abc_16259_n2606_1) );
  AND2X2 AND2X2_1760 ( .A(AES_CORE_DATAPATH__abc_16259_n5943), .B(AES_CORE_DATAPATH__abc_16259_n5942), .Y(AES_CORE_DATAPATH__abc_16259_n5944) );
  AND2X2 AND2X2_1761 ( .A(AES_CORE_DATAPATH__abc_16259_n5944), .B(AES_CORE_DATAPATH__abc_16259_n5659_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n5945) );
  AND2X2 AND2X2_1762 ( .A(AES_CORE_DATAPATH__abc_16259_n5658_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__31_), .Y(AES_CORE_DATAPATH__abc_16259_n5946) );
  AND2X2 AND2X2_1763 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__0_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n5948) );
  AND2X2 AND2X2_1764 ( .A(AES_CORE_DATAPATH__abc_16259_n5663), .B(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n5949) );
  AND2X2 AND2X2_1765 ( .A(AES_CORE_DATAPATH__abc_16259_n5951), .B(AES_CORE_DATAPATH__abc_16259_n5952), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__1_) );
  AND2X2 AND2X2_1766 ( .A(AES_CORE_DATAPATH__abc_16259_n5954), .B(AES_CORE_DATAPATH__abc_16259_n5955), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__2_) );
  AND2X2 AND2X2_1767 ( .A(AES_CORE_DATAPATH__abc_16259_n5957), .B(AES_CORE_DATAPATH__abc_16259_n5958), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__3_) );
  AND2X2 AND2X2_1768 ( .A(AES_CORE_DATAPATH__abc_16259_n5960), .B(AES_CORE_DATAPATH__abc_16259_n5961), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__4_) );
  AND2X2 AND2X2_1769 ( .A(AES_CORE_DATAPATH__abc_16259_n5963), .B(AES_CORE_DATAPATH__abc_16259_n5964), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__5_) );
  AND2X2 AND2X2_177 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf1), .B(AES_CORE_DATAPATH_iv_0__14_), .Y(AES_CORE_DATAPATH__abc_16259_n2608_1) );
  AND2X2 AND2X2_1770 ( .A(AES_CORE_DATAPATH__abc_16259_n5966), .B(AES_CORE_DATAPATH__abc_16259_n5967), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__6_) );
  AND2X2 AND2X2_1771 ( .A(AES_CORE_DATAPATH__abc_16259_n5969), .B(AES_CORE_DATAPATH__abc_16259_n5970), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__7_) );
  AND2X2 AND2X2_1772 ( .A(AES_CORE_DATAPATH__abc_16259_n5972), .B(AES_CORE_DATAPATH__abc_16259_n5973), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__8_) );
  AND2X2 AND2X2_1773 ( .A(AES_CORE_DATAPATH__abc_16259_n5975), .B(AES_CORE_DATAPATH__abc_16259_n5976), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__9_) );
  AND2X2 AND2X2_1774 ( .A(AES_CORE_DATAPATH__abc_16259_n5978), .B(AES_CORE_DATAPATH__abc_16259_n5979), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__10_) );
  AND2X2 AND2X2_1775 ( .A(AES_CORE_DATAPATH__abc_16259_n5981), .B(AES_CORE_DATAPATH__abc_16259_n5982), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__11_) );
  AND2X2 AND2X2_1776 ( .A(AES_CORE_DATAPATH__abc_16259_n5984), .B(AES_CORE_DATAPATH__abc_16259_n5985), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__12_) );
  AND2X2 AND2X2_1777 ( .A(AES_CORE_DATAPATH__abc_16259_n5987), .B(AES_CORE_DATAPATH__abc_16259_n5988), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__13_) );
  AND2X2 AND2X2_1778 ( .A(AES_CORE_DATAPATH__abc_16259_n5990), .B(AES_CORE_DATAPATH__abc_16259_n5991), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__14_) );
  AND2X2 AND2X2_1779 ( .A(AES_CORE_DATAPATH__abc_16259_n5993), .B(AES_CORE_DATAPATH__abc_16259_n5994), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__15_) );
  AND2X2 AND2X2_178 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf0), .B(AES_CORE_DATAPATH_iv_1__14_), .Y(AES_CORE_DATAPATH__abc_16259_n2609_1) );
  AND2X2 AND2X2_1780 ( .A(AES_CORE_DATAPATH__abc_16259_n5996), .B(AES_CORE_DATAPATH__abc_16259_n5997), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__16_) );
  AND2X2 AND2X2_1781 ( .A(AES_CORE_DATAPATH__abc_16259_n5999), .B(AES_CORE_DATAPATH__abc_16259_n6000), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__17_) );
  AND2X2 AND2X2_1782 ( .A(AES_CORE_DATAPATH__abc_16259_n6002), .B(AES_CORE_DATAPATH__abc_16259_n6003), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__18_) );
  AND2X2 AND2X2_1783 ( .A(AES_CORE_DATAPATH__abc_16259_n6005), .B(AES_CORE_DATAPATH__abc_16259_n6006), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__19_) );
  AND2X2 AND2X2_1784 ( .A(AES_CORE_DATAPATH__abc_16259_n6008), .B(AES_CORE_DATAPATH__abc_16259_n6009), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__20_) );
  AND2X2 AND2X2_1785 ( .A(AES_CORE_DATAPATH__abc_16259_n6011), .B(AES_CORE_DATAPATH__abc_16259_n6012), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__21_) );
  AND2X2 AND2X2_1786 ( .A(AES_CORE_DATAPATH__abc_16259_n6014), .B(AES_CORE_DATAPATH__abc_16259_n6015), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__22_) );
  AND2X2 AND2X2_1787 ( .A(AES_CORE_DATAPATH__abc_16259_n6017), .B(AES_CORE_DATAPATH__abc_16259_n6018), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__23_) );
  AND2X2 AND2X2_1788 ( .A(AES_CORE_DATAPATH__abc_16259_n6020), .B(AES_CORE_DATAPATH__abc_16259_n6021), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__24_) );
  AND2X2 AND2X2_1789 ( .A(AES_CORE_DATAPATH__abc_16259_n6023), .B(AES_CORE_DATAPATH__abc_16259_n6024), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__25_) );
  AND2X2 AND2X2_179 ( .A(AES_CORE_DATAPATH__abc_16259_n2612), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n2613_1) );
  AND2X2 AND2X2_1790 ( .A(AES_CORE_DATAPATH__abc_16259_n6026), .B(AES_CORE_DATAPATH__abc_16259_n6027), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__26_) );
  AND2X2 AND2X2_1791 ( .A(AES_CORE_DATAPATH__abc_16259_n6029), .B(AES_CORE_DATAPATH__abc_16259_n6030), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__27_) );
  AND2X2 AND2X2_1792 ( .A(AES_CORE_DATAPATH__abc_16259_n6032), .B(AES_CORE_DATAPATH__abc_16259_n6033), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__28_) );
  AND2X2 AND2X2_1793 ( .A(AES_CORE_DATAPATH__abc_16259_n6035), .B(AES_CORE_DATAPATH__abc_16259_n6036), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__29_) );
  AND2X2 AND2X2_1794 ( .A(AES_CORE_DATAPATH__abc_16259_n6038), .B(AES_CORE_DATAPATH__abc_16259_n6039), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__30_) );
  AND2X2 AND2X2_1795 ( .A(AES_CORE_DATAPATH__abc_16259_n6042), .B(AES_CORE_DATAPATH__abc_16259_n6041), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__31_) );
  AND2X2 AND2X2_1796 ( .A(AES_CORE_DATAPATH__abc_16259_n6044_bF_buf4), .B(AES_CORE_DATAPATH_col_0__0_), .Y(AES_CORE_DATAPATH__abc_16259_n6045) );
  AND2X2 AND2X2_1797 ( .A(AES_CORE_DATAPATH__abc_16259_n2457_1), .B(AES_CORE_DATAPATH_col_sel_pp2_1_), .Y(AES_CORE_DATAPATH__abc_16259_n6046) );
  AND2X2 AND2X2_1798 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk_bF_buf1), .B(AES_CORE_CONTROL_UNIT_col_sel_1_), .Y(AES_CORE_DATAPATH__abc_16259_n6047) );
  AND2X2 AND2X2_1799 ( .A(AES_CORE_DATAPATH__abc_16259_n2457_1), .B(AES_CORE_DATAPATH_col_sel_pp2_0_), .Y(AES_CORE_DATAPATH__abc_16259_n6050) );
  AND2X2 AND2X2_18 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n93_1), .B(AES_CORE_CONTROL_UNIT__abc_15841_n87_1), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n94) );
  AND2X2 AND2X2_180 ( .A(AES_CORE_DATAPATH__abc_16259_n2611_1), .B(AES_CORE_DATAPATH__abc_16259_n2613_1), .Y(AES_CORE_DATAPATH__abc_16259_n2614_1) );
  AND2X2 AND2X2_1800 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk_bF_buf0), .B(AES_CORE_CONTROL_UNIT_col_sel_0_), .Y(AES_CORE_DATAPATH__abc_16259_n6051) );
  AND2X2 AND2X2_1801 ( .A(AES_CORE_DATAPATH__abc_16259_n6049), .B(AES_CORE_DATAPATH__abc_16259_n6052), .Y(AES_CORE_DATAPATH__abc_16259_n6053) );
  AND2X2 AND2X2_1802 ( .A(AES_CORE_DATAPATH__abc_16259_n2868_1), .B(AES_CORE_DATAPATH__abc_16259_n6053_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6054) );
  AND2X2 AND2X2_1803 ( .A(AES_CORE_DATAPATH__abc_16259_n6055), .B(AES_CORE_DATAPATH__abc_16259_n6048), .Y(AES_CORE_DATAPATH__abc_16259_n6056) );
  AND2X2 AND2X2_1804 ( .A(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf9), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n6058) );
  AND2X2 AND2X2_1805 ( .A(AES_CORE_DATAPATH__abc_16259_n2868_1), .B(AES_CORE_DATAPATH__abc_16259_n6059_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n6060) );
  AND2X2 AND2X2_1806 ( .A(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf5), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_0_), .Y(AES_CORE_DATAPATH__abc_16259_n6061) );
  AND2X2 AND2X2_1807 ( .A(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf8), .B(first_block), .Y(AES_CORE_DATAPATH__abc_16259_n6063) );
  AND2X2 AND2X2_1808 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf6), .B(AES_CORE_DATAPATH_bkp_3__0_), .Y(AES_CORE_DATAPATH__abc_16259_n6064) );
  AND2X2 AND2X2_1809 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf7), .B(AES_CORE_DATAPATH_bkp_0__0_), .Y(AES_CORE_DATAPATH__abc_16259_n6065) );
  AND2X2 AND2X2_181 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf0), .B(AES_CORE_DATAPATH_iv_3__14_), .Y(AES_CORE_DATAPATH__abc_16259_n2615) );
  AND2X2 AND2X2_1810 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf6), .B(AES_CORE_DATAPATH_bkp_1__0_), .Y(AES_CORE_DATAPATH__abc_16259_n6066) );
  AND2X2 AND2X2_1811 ( .A(AES_CORE_DATAPATH__abc_16259_n6069), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n6070) );
  AND2X2 AND2X2_1812 ( .A(AES_CORE_DATAPATH__abc_16259_n6068), .B(AES_CORE_DATAPATH__abc_16259_n6070), .Y(AES_CORE_DATAPATH__abc_16259_n6071) );
  AND2X2 AND2X2_1813 ( .A(AES_CORE_DATAPATH__abc_16259_n6073), .B(AES_CORE_DATAPATH__abc_16259_n6075), .Y(AES_CORE_DATAPATH__abc_16259_n6076) );
  AND2X2 AND2X2_1814 ( .A(AES_CORE_DATAPATH__abc_16259_n2862_1), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n6080) );
  AND2X2 AND2X2_1815 ( .A(AES_CORE_DATAPATH__abc_16259_n6080), .B(AES_CORE_DATAPATH__abc_16259_n6079), .Y(AES_CORE_DATAPATH__abc_16259_n6081) );
  AND2X2 AND2X2_1816 ( .A(AES_CORE_DATAPATH__abc_16259_n6083), .B(AES_CORE_DATAPATH__abc_16259_n6084), .Y(AES_CORE_DATAPATH__abc_16259_n6085) );
  AND2X2 AND2X2_1817 ( .A(AES_CORE_DATAPATH__abc_16259_n6077), .B(AES_CORE_DATAPATH__abc_16259_n6087), .Y(AES_CORE_DATAPATH__abc_16259_n6088) );
  AND2X2 AND2X2_1818 ( .A(AES_CORE_DATAPATH__abc_16259_n6091), .B(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6092) );
  AND2X2 AND2X2_1819 ( .A(AES_CORE_DATAPATH__abc_16259_n6090), .B(AES_CORE_DATAPATH__abc_16259_n6092_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6093) );
  AND2X2 AND2X2_182 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf0), .B(AES_CORE_DATAPATH_iv_0__15_), .Y(AES_CORE_DATAPATH__abc_16259_n2617) );
  AND2X2 AND2X2_1820 ( .A(AES_CORE_DATAPATH__abc_16259_n6089), .B(AES_CORE_DATAPATH__abc_16259_n6093), .Y(AES_CORE_DATAPATH__abc_16259_n6094) );
  AND2X2 AND2X2_1821 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf12), .B(AES_CORE_DATAPATH__abc_16259_n6057_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6095) );
  AND2X2 AND2X2_1822 ( .A(AES_CORE_DATAPATH__abc_16259_n6098), .B(AES_CORE_CONTROL_UNIT_mode_cbc_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6099) );
  AND2X2 AND2X2_1823 ( .A(AES_CORE_DATAPATH__abc_16259_n6096), .B(AES_CORE_DATAPATH__abc_16259_n6099), .Y(AES_CORE_DATAPATH__abc_16259_n6100) );
  AND2X2 AND2X2_1824 ( .A(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf7), .B(AES_CORE_DATAPATH__abc_16259_n6091), .Y(AES_CORE_DATAPATH__abc_16259_n6101) );
  AND2X2 AND2X2_1825 ( .A(AES_CORE_DATAPATH__abc_16259_n6101_bF_buf4), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_0_), .Y(AES_CORE_DATAPATH__abc_16259_n6102) );
  AND2X2 AND2X2_1826 ( .A(AES_CORE_DATAPATH__abc_16259_n6104), .B(AES_CORE_DATAPATH__abc_16259_n6056_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6105) );
  AND2X2 AND2X2_1827 ( .A(AES_CORE_DATAPATH__abc_16259_n6049), .B(AES_CORE_DATAPATH__abc_16259_n6055), .Y(AES_CORE_DATAPATH__abc_16259_n6107) );
  AND2X2 AND2X2_1828 ( .A(AES_CORE_DATAPATH__abc_16259_n6108), .B(AES_CORE_DATAPATH__abc_16259_n6109), .Y(AES_CORE_DATAPATH__abc_16259_n6110) );
  AND2X2 AND2X2_1829 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf9), .B(AES_CORE_DATAPATH__abc_16259_n6110), .Y(AES_CORE_DATAPATH__abc_16259_n6111) );
  AND2X2 AND2X2_183 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf7), .B(AES_CORE_DATAPATH_iv_1__15_), .Y(AES_CORE_DATAPATH__abc_16259_n2618_1) );
  AND2X2 AND2X2_1830 ( .A(AES_CORE_DATAPATH__abc_16259_n6112), .B(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6113) );
  AND2X2 AND2X2_1831 ( .A(AES_CORE_DATAPATH__abc_16259_n6044_bF_buf3), .B(AES_CORE_DATAPATH_col_0__1_), .Y(AES_CORE_DATAPATH__abc_16259_n6115) );
  AND2X2 AND2X2_1832 ( .A(AES_CORE_DATAPATH__abc_16259_n6116), .B(AES_CORE_DATAPATH__abc_16259_n6117), .Y(AES_CORE_DATAPATH__abc_16259_n6118) );
  AND2X2 AND2X2_1833 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf6), .B(AES_CORE_DATAPATH_bkp_0__1_), .Y(AES_CORE_DATAPATH__abc_16259_n6119) );
  AND2X2 AND2X2_1834 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf5), .B(AES_CORE_DATAPATH_bkp_1__1_), .Y(AES_CORE_DATAPATH__abc_16259_n6120) );
  AND2X2 AND2X2_1835 ( .A(AES_CORE_DATAPATH__abc_16259_n6123), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n6124) );
  AND2X2 AND2X2_1836 ( .A(AES_CORE_DATAPATH__abc_16259_n6122), .B(AES_CORE_DATAPATH__abc_16259_n6124), .Y(AES_CORE_DATAPATH__abc_16259_n6125) );
  AND2X2 AND2X2_1837 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf5), .B(AES_CORE_DATAPATH_bkp_3__1_), .Y(AES_CORE_DATAPATH__abc_16259_n6126) );
  AND2X2 AND2X2_1838 ( .A(AES_CORE_DATAPATH__abc_16259_n6128), .B(AES_CORE_DATAPATH__abc_16259_n6129), .Y(AES_CORE_DATAPATH__abc_16259_n6130) );
  AND2X2 AND2X2_1839 ( .A(AES_CORE_DATAPATH__abc_16259_n2900), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n6133) );
  AND2X2 AND2X2_184 ( .A(AES_CORE_DATAPATH__abc_16259_n2621_1), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n2622) );
  AND2X2 AND2X2_1840 ( .A(AES_CORE_DATAPATH__abc_16259_n6133), .B(AES_CORE_DATAPATH__abc_16259_n6132), .Y(AES_CORE_DATAPATH__abc_16259_n6134) );
  AND2X2 AND2X2_1841 ( .A(AES_CORE_DATAPATH__abc_16259_n6136), .B(AES_CORE_DATAPATH__abc_16259_n6059_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6137) );
  AND2X2 AND2X2_1842 ( .A(AES_CORE_DATAPATH__abc_16259_n6131), .B(AES_CORE_DATAPATH__abc_16259_n6141), .Y(AES_CORE_DATAPATH__abc_16259_n6142) );
  AND2X2 AND2X2_1843 ( .A(AES_CORE_DATAPATH__abc_16259_n6144), .B(AES_CORE_DATAPATH__abc_16259_n6092_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6145) );
  AND2X2 AND2X2_1844 ( .A(AES_CORE_DATAPATH__abc_16259_n6143), .B(AES_CORE_DATAPATH__abc_16259_n6145), .Y(AES_CORE_DATAPATH__abc_16259_n6146) );
  AND2X2 AND2X2_1845 ( .A(AES_CORE_DATAPATH__abc_16259_n6148), .B(AES_CORE_CONTROL_UNIT_mode_cbc_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6149) );
  AND2X2 AND2X2_1846 ( .A(AES_CORE_DATAPATH__abc_16259_n6147), .B(AES_CORE_DATAPATH__abc_16259_n6149), .Y(AES_CORE_DATAPATH__abc_16259_n6150) );
  AND2X2 AND2X2_1847 ( .A(AES_CORE_DATAPATH__abc_16259_n6101_bF_buf3), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_1_), .Y(AES_CORE_DATAPATH__abc_16259_n6151) );
  AND2X2 AND2X2_1848 ( .A(AES_CORE_DATAPATH__abc_16259_n6153), .B(AES_CORE_DATAPATH__abc_16259_n6056_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6154) );
  AND2X2 AND2X2_1849 ( .A(AES_CORE_DATAPATH__abc_16259_n2909_1), .B(AES_CORE_DATAPATH__abc_16259_n6053_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6155) );
  AND2X2 AND2X2_185 ( .A(AES_CORE_DATAPATH__abc_16259_n2620), .B(AES_CORE_DATAPATH__abc_16259_n2622), .Y(AES_CORE_DATAPATH__abc_16259_n2623_1) );
  AND2X2 AND2X2_1850 ( .A(AES_CORE_DATAPATH__abc_16259_n6157), .B(AES_CORE_DATAPATH__abc_16259_n6158), .Y(AES_CORE_DATAPATH__abc_16259_n6159) );
  AND2X2 AND2X2_1851 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf8), .B(AES_CORE_DATAPATH__abc_16259_n6159), .Y(AES_CORE_DATAPATH__abc_16259_n6160) );
  AND2X2 AND2X2_1852 ( .A(AES_CORE_DATAPATH__abc_16259_n6161), .B(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6162) );
  AND2X2 AND2X2_1853 ( .A(AES_CORE_DATAPATH__abc_16259_n6044_bF_buf2), .B(AES_CORE_DATAPATH_col_0__2_), .Y(AES_CORE_DATAPATH__abc_16259_n6164) );
  AND2X2 AND2X2_1854 ( .A(AES_CORE_DATAPATH__abc_16259_n2949_1), .B(AES_CORE_DATAPATH__abc_16259_n6059_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6165) );
  AND2X2 AND2X2_1855 ( .A(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf2), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_2_), .Y(AES_CORE_DATAPATH__abc_16259_n6166) );
  AND2X2 AND2X2_1856 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf5), .B(AES_CORE_DATAPATH_bkp_0__2_), .Y(AES_CORE_DATAPATH__abc_16259_n6168) );
  AND2X2 AND2X2_1857 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf4), .B(AES_CORE_DATAPATH_bkp_1__2_), .Y(AES_CORE_DATAPATH__abc_16259_n6169) );
  AND2X2 AND2X2_1858 ( .A(AES_CORE_DATAPATH__abc_16259_n6172), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n6173) );
  AND2X2 AND2X2_1859 ( .A(AES_CORE_DATAPATH__abc_16259_n6171), .B(AES_CORE_DATAPATH__abc_16259_n6173), .Y(AES_CORE_DATAPATH__abc_16259_n6174) );
  AND2X2 AND2X2_186 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf7), .B(AES_CORE_DATAPATH_iv_3__15_), .Y(AES_CORE_DATAPATH__abc_16259_n2624_1) );
  AND2X2 AND2X2_1860 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf4), .B(AES_CORE_DATAPATH_bkp_3__2_), .Y(AES_CORE_DATAPATH__abc_16259_n6175) );
  AND2X2 AND2X2_1861 ( .A(AES_CORE_DATAPATH__abc_16259_n6177), .B(AES_CORE_DATAPATH__abc_16259_n6178), .Y(AES_CORE_DATAPATH__abc_16259_n6179) );
  AND2X2 AND2X2_1862 ( .A(AES_CORE_DATAPATH__abc_16259_n2940_1), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6182) );
  AND2X2 AND2X2_1863 ( .A(AES_CORE_DATAPATH__abc_16259_n6182), .B(AES_CORE_DATAPATH__abc_16259_n6181), .Y(AES_CORE_DATAPATH__abc_16259_n6183) );
  AND2X2 AND2X2_1864 ( .A(AES_CORE_DATAPATH__abc_16259_n6186), .B(AES_CORE_DATAPATH__abc_16259_n6187), .Y(AES_CORE_DATAPATH__abc_16259_n6188) );
  AND2X2 AND2X2_1865 ( .A(AES_CORE_DATAPATH__abc_16259_n6180), .B(AES_CORE_DATAPATH__abc_16259_n6190), .Y(AES_CORE_DATAPATH__abc_16259_n6191) );
  AND2X2 AND2X2_1866 ( .A(AES_CORE_DATAPATH__abc_16259_n6193), .B(AES_CORE_DATAPATH__abc_16259_n6092_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6194) );
  AND2X2 AND2X2_1867 ( .A(AES_CORE_DATAPATH__abc_16259_n6192), .B(AES_CORE_DATAPATH__abc_16259_n6194), .Y(AES_CORE_DATAPATH__abc_16259_n6195) );
  AND2X2 AND2X2_1868 ( .A(AES_CORE_DATAPATH__abc_16259_n6197), .B(AES_CORE_CONTROL_UNIT_mode_cbc_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n6198) );
  AND2X2 AND2X2_1869 ( .A(AES_CORE_DATAPATH__abc_16259_n6196), .B(AES_CORE_DATAPATH__abc_16259_n6198), .Y(AES_CORE_DATAPATH__abc_16259_n6199) );
  AND2X2 AND2X2_187 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf7), .B(AES_CORE_DATAPATH_iv_0__16_), .Y(AES_CORE_DATAPATH__abc_16259_n2626_1) );
  AND2X2 AND2X2_1870 ( .A(AES_CORE_DATAPATH__abc_16259_n6101_bF_buf2), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_2_), .Y(AES_CORE_DATAPATH__abc_16259_n6200) );
  AND2X2 AND2X2_1871 ( .A(AES_CORE_DATAPATH__abc_16259_n6202), .B(AES_CORE_DATAPATH__abc_16259_n6056_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6203) );
  AND2X2 AND2X2_1872 ( .A(AES_CORE_DATAPATH__abc_16259_n2949_1), .B(AES_CORE_DATAPATH__abc_16259_n6053_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6204) );
  AND2X2 AND2X2_1873 ( .A(AES_CORE_DATAPATH__abc_16259_n6206), .B(AES_CORE_DATAPATH__abc_16259_n6207), .Y(AES_CORE_DATAPATH__abc_16259_n6208) );
  AND2X2 AND2X2_1874 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf7), .B(AES_CORE_DATAPATH__abc_16259_n6208), .Y(AES_CORE_DATAPATH__abc_16259_n6209) );
  AND2X2 AND2X2_1875 ( .A(AES_CORE_DATAPATH__abc_16259_n6210), .B(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6211) );
  AND2X2 AND2X2_1876 ( .A(AES_CORE_DATAPATH__abc_16259_n6044_bF_buf1), .B(AES_CORE_DATAPATH_col_0__3_), .Y(AES_CORE_DATAPATH__abc_16259_n6213) );
  AND2X2 AND2X2_1877 ( .A(AES_CORE_DATAPATH__abc_16259_n2989), .B(AES_CORE_DATAPATH__abc_16259_n6059_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6214) );
  AND2X2 AND2X2_1878 ( .A(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf0), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_3_), .Y(AES_CORE_DATAPATH__abc_16259_n6215) );
  AND2X2 AND2X2_1879 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf4), .B(AES_CORE_DATAPATH_bkp_0__3_), .Y(AES_CORE_DATAPATH__abc_16259_n6217) );
  AND2X2 AND2X2_188 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf6), .B(AES_CORE_DATAPATH_iv_1__16_), .Y(AES_CORE_DATAPATH__abc_16259_n2627) );
  AND2X2 AND2X2_1880 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1__3_), .Y(AES_CORE_DATAPATH__abc_16259_n6218) );
  AND2X2 AND2X2_1881 ( .A(AES_CORE_DATAPATH__abc_16259_n6221), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6222) );
  AND2X2 AND2X2_1882 ( .A(AES_CORE_DATAPATH__abc_16259_n6220), .B(AES_CORE_DATAPATH__abc_16259_n6222), .Y(AES_CORE_DATAPATH__abc_16259_n6223) );
  AND2X2 AND2X2_1883 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf3), .B(AES_CORE_DATAPATH_bkp_3__3_), .Y(AES_CORE_DATAPATH__abc_16259_n6224) );
  AND2X2 AND2X2_1884 ( .A(AES_CORE_DATAPATH__abc_16259_n6227), .B(AES_CORE_DATAPATH__abc_16259_n6226), .Y(AES_CORE_DATAPATH__abc_16259_n6228) );
  AND2X2 AND2X2_1885 ( .A(AES_CORE_DATAPATH__abc_16259_n2980_1), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6231) );
  AND2X2 AND2X2_1886 ( .A(AES_CORE_DATAPATH__abc_16259_n6231), .B(AES_CORE_DATAPATH__abc_16259_n6230), .Y(AES_CORE_DATAPATH__abc_16259_n6232) );
  AND2X2 AND2X2_1887 ( .A(AES_CORE_DATAPATH__abc_16259_n6235), .B(AES_CORE_DATAPATH__abc_16259_n6236), .Y(AES_CORE_DATAPATH__abc_16259_n6237) );
  AND2X2 AND2X2_1888 ( .A(AES_CORE_DATAPATH__abc_16259_n6229), .B(AES_CORE_DATAPATH__abc_16259_n6239), .Y(AES_CORE_DATAPATH__abc_16259_n6240) );
  AND2X2 AND2X2_1889 ( .A(AES_CORE_DATAPATH__abc_16259_n6242), .B(AES_CORE_DATAPATH__abc_16259_n6092_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6243) );
  AND2X2 AND2X2_189 ( .A(AES_CORE_DATAPATH__abc_16259_n2630), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n2631_1) );
  AND2X2 AND2X2_1890 ( .A(AES_CORE_DATAPATH__abc_16259_n6241), .B(AES_CORE_DATAPATH__abc_16259_n6243), .Y(AES_CORE_DATAPATH__abc_16259_n6244) );
  AND2X2 AND2X2_1891 ( .A(AES_CORE_DATAPATH__abc_16259_n6246), .B(AES_CORE_CONTROL_UNIT_mode_cbc_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6247) );
  AND2X2 AND2X2_1892 ( .A(AES_CORE_DATAPATH__abc_16259_n6245), .B(AES_CORE_DATAPATH__abc_16259_n6247), .Y(AES_CORE_DATAPATH__abc_16259_n6248) );
  AND2X2 AND2X2_1893 ( .A(AES_CORE_DATAPATH__abc_16259_n6101_bF_buf1), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_3_), .Y(AES_CORE_DATAPATH__abc_16259_n6249) );
  AND2X2 AND2X2_1894 ( .A(AES_CORE_DATAPATH__abc_16259_n6251), .B(AES_CORE_DATAPATH__abc_16259_n6056_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6252) );
  AND2X2 AND2X2_1895 ( .A(AES_CORE_DATAPATH__abc_16259_n2989), .B(AES_CORE_DATAPATH__abc_16259_n6053_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6253) );
  AND2X2 AND2X2_1896 ( .A(AES_CORE_DATAPATH__abc_16259_n6255), .B(AES_CORE_DATAPATH__abc_16259_n6256), .Y(AES_CORE_DATAPATH__abc_16259_n6257) );
  AND2X2 AND2X2_1897 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf6), .B(AES_CORE_DATAPATH__abc_16259_n6257), .Y(AES_CORE_DATAPATH__abc_16259_n6258) );
  AND2X2 AND2X2_1898 ( .A(AES_CORE_DATAPATH__abc_16259_n6259), .B(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n6260) );
  AND2X2 AND2X2_1899 ( .A(AES_CORE_DATAPATH__abc_16259_n6044_bF_buf0), .B(AES_CORE_DATAPATH_col_0__4_), .Y(AES_CORE_DATAPATH__abc_16259_n6262) );
  AND2X2 AND2X2_19 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n89_1), .B(\op_mode[1] ), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n95) );
  AND2X2 AND2X2_190 ( .A(AES_CORE_DATAPATH__abc_16259_n2629_1), .B(AES_CORE_DATAPATH__abc_16259_n2631_1), .Y(AES_CORE_DATAPATH__abc_16259_n2632) );
  AND2X2 AND2X2_1900 ( .A(AES_CORE_DATAPATH__abc_16259_n3029), .B(AES_CORE_DATAPATH__abc_16259_n6059_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n6263) );
  AND2X2 AND2X2_1901 ( .A(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf5), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_4_), .Y(AES_CORE_DATAPATH__abc_16259_n6264) );
  AND2X2 AND2X2_1902 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf3), .B(AES_CORE_DATAPATH_bkp_0__4_), .Y(AES_CORE_DATAPATH__abc_16259_n6266) );
  AND2X2 AND2X2_1903 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf2), .B(AES_CORE_DATAPATH_bkp_1__4_), .Y(AES_CORE_DATAPATH__abc_16259_n6267) );
  AND2X2 AND2X2_1904 ( .A(AES_CORE_DATAPATH__abc_16259_n6270), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6271) );
  AND2X2 AND2X2_1905 ( .A(AES_CORE_DATAPATH__abc_16259_n6269), .B(AES_CORE_DATAPATH__abc_16259_n6271), .Y(AES_CORE_DATAPATH__abc_16259_n6272) );
  AND2X2 AND2X2_1906 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf2), .B(AES_CORE_DATAPATH_bkp_3__4_), .Y(AES_CORE_DATAPATH__abc_16259_n6273) );
  AND2X2 AND2X2_1907 ( .A(AES_CORE_DATAPATH__abc_16259_n6275), .B(AES_CORE_DATAPATH__abc_16259_n6276), .Y(AES_CORE_DATAPATH__abc_16259_n6277) );
  AND2X2 AND2X2_1908 ( .A(AES_CORE_DATAPATH__abc_16259_n3020), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6280) );
  AND2X2 AND2X2_1909 ( .A(AES_CORE_DATAPATH__abc_16259_n6280), .B(AES_CORE_DATAPATH__abc_16259_n6279), .Y(AES_CORE_DATAPATH__abc_16259_n6281) );
  AND2X2 AND2X2_191 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf6), .B(AES_CORE_DATAPATH_iv_3__16_), .Y(AES_CORE_DATAPATH__abc_16259_n2633_1) );
  AND2X2 AND2X2_1910 ( .A(AES_CORE_DATAPATH__abc_16259_n6284), .B(AES_CORE_DATAPATH__abc_16259_n6285), .Y(AES_CORE_DATAPATH__abc_16259_n6286) );
  AND2X2 AND2X2_1911 ( .A(AES_CORE_DATAPATH__abc_16259_n6278), .B(AES_CORE_DATAPATH__abc_16259_n6288), .Y(AES_CORE_DATAPATH__abc_16259_n6289) );
  AND2X2 AND2X2_1912 ( .A(AES_CORE_DATAPATH__abc_16259_n6291), .B(AES_CORE_DATAPATH__abc_16259_n6092_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n6292) );
  AND2X2 AND2X2_1913 ( .A(AES_CORE_DATAPATH__abc_16259_n6290), .B(AES_CORE_DATAPATH__abc_16259_n6292), .Y(AES_CORE_DATAPATH__abc_16259_n6293) );
  AND2X2 AND2X2_1914 ( .A(AES_CORE_DATAPATH__abc_16259_n6295), .B(AES_CORE_CONTROL_UNIT_mode_cbc_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6296) );
  AND2X2 AND2X2_1915 ( .A(AES_CORE_DATAPATH__abc_16259_n6294), .B(AES_CORE_DATAPATH__abc_16259_n6296), .Y(AES_CORE_DATAPATH__abc_16259_n6297) );
  AND2X2 AND2X2_1916 ( .A(AES_CORE_DATAPATH__abc_16259_n6101_bF_buf0), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_4_), .Y(AES_CORE_DATAPATH__abc_16259_n6298) );
  AND2X2 AND2X2_1917 ( .A(AES_CORE_DATAPATH__abc_16259_n6300), .B(AES_CORE_DATAPATH__abc_16259_n6056_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n6301) );
  AND2X2 AND2X2_1918 ( .A(AES_CORE_DATAPATH__abc_16259_n3029), .B(AES_CORE_DATAPATH__abc_16259_n6053_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n6302) );
  AND2X2 AND2X2_1919 ( .A(AES_CORE_DATAPATH__abc_16259_n6304), .B(AES_CORE_DATAPATH__abc_16259_n6305), .Y(AES_CORE_DATAPATH__abc_16259_n6306) );
  AND2X2 AND2X2_192 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf6), .B(AES_CORE_DATAPATH_iv_0__17_), .Y(AES_CORE_DATAPATH__abc_16259_n2635) );
  AND2X2 AND2X2_1920 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf5), .B(AES_CORE_DATAPATH__abc_16259_n6306), .Y(AES_CORE_DATAPATH__abc_16259_n6307) );
  AND2X2 AND2X2_1921 ( .A(AES_CORE_DATAPATH__abc_16259_n6308), .B(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n6309) );
  AND2X2 AND2X2_1922 ( .A(AES_CORE_DATAPATH__abc_16259_n6044_bF_buf4), .B(AES_CORE_DATAPATH_col_0__5_), .Y(AES_CORE_DATAPATH__abc_16259_n6311) );
  AND2X2 AND2X2_1923 ( .A(AES_CORE_DATAPATH__abc_16259_n3069_1), .B(AES_CORE_DATAPATH__abc_16259_n6059_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n6312) );
  AND2X2 AND2X2_1924 ( .A(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf3), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_5_), .Y(AES_CORE_DATAPATH__abc_16259_n6313) );
  AND2X2 AND2X2_1925 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf2), .B(AES_CORE_DATAPATH_bkp_0__5_), .Y(AES_CORE_DATAPATH__abc_16259_n6315) );
  AND2X2 AND2X2_1926 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf1), .B(AES_CORE_DATAPATH_bkp_1__5_), .Y(AES_CORE_DATAPATH__abc_16259_n6316) );
  AND2X2 AND2X2_1927 ( .A(AES_CORE_DATAPATH__abc_16259_n6319), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6320) );
  AND2X2 AND2X2_1928 ( .A(AES_CORE_DATAPATH__abc_16259_n6318), .B(AES_CORE_DATAPATH__abc_16259_n6320), .Y(AES_CORE_DATAPATH__abc_16259_n6321) );
  AND2X2 AND2X2_1929 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf1), .B(AES_CORE_DATAPATH_bkp_3__5_), .Y(AES_CORE_DATAPATH__abc_16259_n6322) );
  AND2X2 AND2X2_193 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf5), .B(AES_CORE_DATAPATH_iv_1__17_), .Y(AES_CORE_DATAPATH__abc_16259_n2636_1) );
  AND2X2 AND2X2_1930 ( .A(AES_CORE_DATAPATH__abc_16259_n6325), .B(AES_CORE_DATAPATH__abc_16259_n6324), .Y(AES_CORE_DATAPATH__abc_16259_n6326) );
  AND2X2 AND2X2_1931 ( .A(AES_CORE_DATAPATH__abc_16259_n3060), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6329) );
  AND2X2 AND2X2_1932 ( .A(AES_CORE_DATAPATH__abc_16259_n6329), .B(AES_CORE_DATAPATH__abc_16259_n6328), .Y(AES_CORE_DATAPATH__abc_16259_n6330) );
  AND2X2 AND2X2_1933 ( .A(AES_CORE_DATAPATH__abc_16259_n6333), .B(AES_CORE_DATAPATH__abc_16259_n6334), .Y(AES_CORE_DATAPATH__abc_16259_n6335) );
  AND2X2 AND2X2_1934 ( .A(AES_CORE_DATAPATH__abc_16259_n6327), .B(AES_CORE_DATAPATH__abc_16259_n6337), .Y(AES_CORE_DATAPATH__abc_16259_n6338) );
  AND2X2 AND2X2_1935 ( .A(AES_CORE_DATAPATH__abc_16259_n6340), .B(AES_CORE_DATAPATH__abc_16259_n6092_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6341) );
  AND2X2 AND2X2_1936 ( .A(AES_CORE_DATAPATH__abc_16259_n6339), .B(AES_CORE_DATAPATH__abc_16259_n6341), .Y(AES_CORE_DATAPATH__abc_16259_n6342) );
  AND2X2 AND2X2_1937 ( .A(AES_CORE_DATAPATH__abc_16259_n6344), .B(AES_CORE_CONTROL_UNIT_mode_cbc_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6345) );
  AND2X2 AND2X2_1938 ( .A(AES_CORE_DATAPATH__abc_16259_n6343), .B(AES_CORE_DATAPATH__abc_16259_n6345), .Y(AES_CORE_DATAPATH__abc_16259_n6346) );
  AND2X2 AND2X2_1939 ( .A(AES_CORE_DATAPATH__abc_16259_n6101_bF_buf4), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_5_), .Y(AES_CORE_DATAPATH__abc_16259_n6347) );
  AND2X2 AND2X2_194 ( .A(AES_CORE_DATAPATH__abc_16259_n2639_1), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n2640) );
  AND2X2 AND2X2_1940 ( .A(AES_CORE_DATAPATH__abc_16259_n6349), .B(AES_CORE_DATAPATH__abc_16259_n6056_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6350) );
  AND2X2 AND2X2_1941 ( .A(AES_CORE_DATAPATH__abc_16259_n3069_1), .B(AES_CORE_DATAPATH__abc_16259_n6053_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6351) );
  AND2X2 AND2X2_1942 ( .A(AES_CORE_DATAPATH__abc_16259_n6353), .B(AES_CORE_DATAPATH__abc_16259_n6354), .Y(AES_CORE_DATAPATH__abc_16259_n6355) );
  AND2X2 AND2X2_1943 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n6355), .Y(AES_CORE_DATAPATH__abc_16259_n6356) );
  AND2X2 AND2X2_1944 ( .A(AES_CORE_DATAPATH__abc_16259_n6357), .B(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6358) );
  AND2X2 AND2X2_1945 ( .A(AES_CORE_DATAPATH__abc_16259_n6044_bF_buf3), .B(AES_CORE_DATAPATH_col_0__6_), .Y(AES_CORE_DATAPATH__abc_16259_n6360) );
  AND2X2 AND2X2_1946 ( .A(AES_CORE_DATAPATH__abc_16259_n3109), .B(AES_CORE_DATAPATH__abc_16259_n6059_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6361) );
  AND2X2 AND2X2_1947 ( .A(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf1), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_6_), .Y(AES_CORE_DATAPATH__abc_16259_n6362) );
  AND2X2 AND2X2_1948 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf1), .B(AES_CORE_DATAPATH_bkp_0__6_), .Y(AES_CORE_DATAPATH__abc_16259_n6364) );
  AND2X2 AND2X2_1949 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf0), .B(AES_CORE_DATAPATH_bkp_1__6_), .Y(AES_CORE_DATAPATH__abc_16259_n6365) );
  AND2X2 AND2X2_195 ( .A(AES_CORE_DATAPATH__abc_16259_n2638_1), .B(AES_CORE_DATAPATH__abc_16259_n2640), .Y(AES_CORE_DATAPATH__abc_16259_n2641_1) );
  AND2X2 AND2X2_1950 ( .A(AES_CORE_DATAPATH__abc_16259_n6368), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6369) );
  AND2X2 AND2X2_1951 ( .A(AES_CORE_DATAPATH__abc_16259_n6367), .B(AES_CORE_DATAPATH__abc_16259_n6369), .Y(AES_CORE_DATAPATH__abc_16259_n6370) );
  AND2X2 AND2X2_1952 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf0), .B(AES_CORE_DATAPATH_bkp_3__6_), .Y(AES_CORE_DATAPATH__abc_16259_n6371) );
  AND2X2 AND2X2_1953 ( .A(AES_CORE_DATAPATH__abc_16259_n6373), .B(AES_CORE_DATAPATH__abc_16259_n6374), .Y(AES_CORE_DATAPATH__abc_16259_n6375) );
  AND2X2 AND2X2_1954 ( .A(AES_CORE_DATAPATH__abc_16259_n3100_1), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n6378) );
  AND2X2 AND2X2_1955 ( .A(AES_CORE_DATAPATH__abc_16259_n6378), .B(AES_CORE_DATAPATH__abc_16259_n6377), .Y(AES_CORE_DATAPATH__abc_16259_n6379) );
  AND2X2 AND2X2_1956 ( .A(AES_CORE_DATAPATH__abc_16259_n6382), .B(AES_CORE_DATAPATH__abc_16259_n6383), .Y(AES_CORE_DATAPATH__abc_16259_n6384) );
  AND2X2 AND2X2_1957 ( .A(AES_CORE_DATAPATH__abc_16259_n6376), .B(AES_CORE_DATAPATH__abc_16259_n6386), .Y(AES_CORE_DATAPATH__abc_16259_n6387) );
  AND2X2 AND2X2_1958 ( .A(AES_CORE_DATAPATH__abc_16259_n6389), .B(AES_CORE_DATAPATH__abc_16259_n6092_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6390) );
  AND2X2 AND2X2_1959 ( .A(AES_CORE_DATAPATH__abc_16259_n6388), .B(AES_CORE_DATAPATH__abc_16259_n6390), .Y(AES_CORE_DATAPATH__abc_16259_n6391) );
  AND2X2 AND2X2_196 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf5), .B(AES_CORE_DATAPATH_iv_3__17_), .Y(AES_CORE_DATAPATH__abc_16259_n2642) );
  AND2X2 AND2X2_1960 ( .A(AES_CORE_DATAPATH__abc_16259_n6393), .B(AES_CORE_CONTROL_UNIT_mode_cbc_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6394) );
  AND2X2 AND2X2_1961 ( .A(AES_CORE_DATAPATH__abc_16259_n6392), .B(AES_CORE_DATAPATH__abc_16259_n6394), .Y(AES_CORE_DATAPATH__abc_16259_n6395) );
  AND2X2 AND2X2_1962 ( .A(AES_CORE_DATAPATH__abc_16259_n6101_bF_buf3), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_6_), .Y(AES_CORE_DATAPATH__abc_16259_n6396) );
  AND2X2 AND2X2_1963 ( .A(AES_CORE_DATAPATH__abc_16259_n6398), .B(AES_CORE_DATAPATH__abc_16259_n6056_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6399) );
  AND2X2 AND2X2_1964 ( .A(AES_CORE_DATAPATH__abc_16259_n3109), .B(AES_CORE_DATAPATH__abc_16259_n6053_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6400) );
  AND2X2 AND2X2_1965 ( .A(AES_CORE_DATAPATH__abc_16259_n6402), .B(AES_CORE_DATAPATH__abc_16259_n6403), .Y(AES_CORE_DATAPATH__abc_16259_n6404) );
  AND2X2 AND2X2_1966 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n6404), .Y(AES_CORE_DATAPATH__abc_16259_n6405) );
  AND2X2 AND2X2_1967 ( .A(AES_CORE_DATAPATH__abc_16259_n6406), .B(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6407) );
  AND2X2 AND2X2_1968 ( .A(AES_CORE_DATAPATH__abc_16259_n6044_bF_buf2), .B(AES_CORE_DATAPATH_col_0__7_), .Y(AES_CORE_DATAPATH__abc_16259_n6409) );
  AND2X2 AND2X2_1969 ( .A(AES_CORE_DATAPATH__abc_16259_n3149_1), .B(AES_CORE_DATAPATH__abc_16259_n6059_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6410) );
  AND2X2 AND2X2_197 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf5), .B(AES_CORE_DATAPATH_iv_0__18_), .Y(AES_CORE_DATAPATH__abc_16259_n2644_1) );
  AND2X2 AND2X2_1970 ( .A(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf6), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_7_), .Y(AES_CORE_DATAPATH__abc_16259_n6411) );
  AND2X2 AND2X2_1971 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf0), .B(AES_CORE_DATAPATH_bkp_0__7_), .Y(AES_CORE_DATAPATH__abc_16259_n6413) );
  AND2X2 AND2X2_1972 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf7), .B(AES_CORE_DATAPATH_bkp_1__7_), .Y(AES_CORE_DATAPATH__abc_16259_n6414) );
  AND2X2 AND2X2_1973 ( .A(AES_CORE_DATAPATH__abc_16259_n6417), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n6418) );
  AND2X2 AND2X2_1974 ( .A(AES_CORE_DATAPATH__abc_16259_n6416), .B(AES_CORE_DATAPATH__abc_16259_n6418), .Y(AES_CORE_DATAPATH__abc_16259_n6419) );
  AND2X2 AND2X2_1975 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf7), .B(AES_CORE_DATAPATH_bkp_3__7_), .Y(AES_CORE_DATAPATH__abc_16259_n6420) );
  AND2X2 AND2X2_1976 ( .A(AES_CORE_DATAPATH__abc_16259_n6422), .B(AES_CORE_DATAPATH__abc_16259_n6423), .Y(AES_CORE_DATAPATH__abc_16259_n6424) );
  AND2X2 AND2X2_1977 ( .A(AES_CORE_DATAPATH__abc_16259_n3140), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n6427) );
  AND2X2 AND2X2_1978 ( .A(AES_CORE_DATAPATH__abc_16259_n6427), .B(AES_CORE_DATAPATH__abc_16259_n6426), .Y(AES_CORE_DATAPATH__abc_16259_n6428) );
  AND2X2 AND2X2_1979 ( .A(AES_CORE_DATAPATH__abc_16259_n6431), .B(AES_CORE_DATAPATH__abc_16259_n6432), .Y(AES_CORE_DATAPATH__abc_16259_n6433) );
  AND2X2 AND2X2_198 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf4), .B(AES_CORE_DATAPATH_iv_1__18_), .Y(AES_CORE_DATAPATH__abc_16259_n2645) );
  AND2X2 AND2X2_1980 ( .A(AES_CORE_DATAPATH__abc_16259_n6425), .B(AES_CORE_DATAPATH__abc_16259_n6435), .Y(AES_CORE_DATAPATH__abc_16259_n6436) );
  AND2X2 AND2X2_1981 ( .A(AES_CORE_DATAPATH__abc_16259_n6438), .B(AES_CORE_DATAPATH__abc_16259_n6092_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6439) );
  AND2X2 AND2X2_1982 ( .A(AES_CORE_DATAPATH__abc_16259_n6437), .B(AES_CORE_DATAPATH__abc_16259_n6439), .Y(AES_CORE_DATAPATH__abc_16259_n6440) );
  AND2X2 AND2X2_1983 ( .A(AES_CORE_DATAPATH__abc_16259_n6442), .B(AES_CORE_CONTROL_UNIT_mode_cbc_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n6443) );
  AND2X2 AND2X2_1984 ( .A(AES_CORE_DATAPATH__abc_16259_n6441), .B(AES_CORE_DATAPATH__abc_16259_n6443), .Y(AES_CORE_DATAPATH__abc_16259_n6444) );
  AND2X2 AND2X2_1985 ( .A(AES_CORE_DATAPATH__abc_16259_n6101_bF_buf2), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_7_), .Y(AES_CORE_DATAPATH__abc_16259_n6445) );
  AND2X2 AND2X2_1986 ( .A(AES_CORE_DATAPATH__abc_16259_n6447), .B(AES_CORE_DATAPATH__abc_16259_n6056_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6448) );
  AND2X2 AND2X2_1987 ( .A(AES_CORE_DATAPATH__abc_16259_n3149_1), .B(AES_CORE_DATAPATH__abc_16259_n6053_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6449) );
  AND2X2 AND2X2_1988 ( .A(AES_CORE_DATAPATH__abc_16259_n6451), .B(AES_CORE_DATAPATH__abc_16259_n6452), .Y(AES_CORE_DATAPATH__abc_16259_n6453) );
  AND2X2 AND2X2_1989 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n6453), .Y(AES_CORE_DATAPATH__abc_16259_n6454) );
  AND2X2 AND2X2_199 ( .A(AES_CORE_DATAPATH__abc_16259_n2648_1), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n2649_1) );
  AND2X2 AND2X2_1990 ( .A(AES_CORE_DATAPATH__abc_16259_n6455), .B(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6456) );
  AND2X2 AND2X2_1991 ( .A(AES_CORE_DATAPATH__abc_16259_n6044_bF_buf1), .B(AES_CORE_DATAPATH_col_0__8_), .Y(AES_CORE_DATAPATH__abc_16259_n6458) );
  AND2X2 AND2X2_1992 ( .A(AES_CORE_DATAPATH__abc_16259_n3189), .B(AES_CORE_DATAPATH__abc_16259_n6059_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6459) );
  AND2X2 AND2X2_1993 ( .A(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf4), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_8_), .Y(AES_CORE_DATAPATH__abc_16259_n6460) );
  AND2X2 AND2X2_1994 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf7), .B(AES_CORE_DATAPATH_bkp_0__8_), .Y(AES_CORE_DATAPATH__abc_16259_n6462) );
  AND2X2 AND2X2_1995 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf6), .B(AES_CORE_DATAPATH_bkp_1__8_), .Y(AES_CORE_DATAPATH__abc_16259_n6463) );
  AND2X2 AND2X2_1996 ( .A(AES_CORE_DATAPATH__abc_16259_n6466), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n6467) );
  AND2X2 AND2X2_1997 ( .A(AES_CORE_DATAPATH__abc_16259_n6465), .B(AES_CORE_DATAPATH__abc_16259_n6467), .Y(AES_CORE_DATAPATH__abc_16259_n6468) );
  AND2X2 AND2X2_1998 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf6), .B(AES_CORE_DATAPATH_bkp_3__8_), .Y(AES_CORE_DATAPATH__abc_16259_n6469) );
  AND2X2 AND2X2_1999 ( .A(AES_CORE_DATAPATH__abc_16259_n6471), .B(AES_CORE_DATAPATH__abc_16259_n6472), .Y(AES_CORE_DATAPATH__abc_16259_n6473) );
  AND2X2 AND2X2_2 ( .A(_abc_15830_n13_1), .B(_abc_15830_n11_1), .Y(AES_CORE_DATAPATH_col_en_host_0_) );
  AND2X2 AND2X2_20 ( .A(start), .B(AES_CORE_CONTROL_UNIT_state_0_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n97) );
  AND2X2 AND2X2_200 ( .A(AES_CORE_DATAPATH__abc_16259_n2647), .B(AES_CORE_DATAPATH__abc_16259_n2649_1), .Y(AES_CORE_DATAPATH__abc_16259_n2650) );
  AND2X2 AND2X2_2000 ( .A(AES_CORE_DATAPATH__abc_16259_n3180), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n6476) );
  AND2X2 AND2X2_2001 ( .A(AES_CORE_DATAPATH__abc_16259_n6476), .B(AES_CORE_DATAPATH__abc_16259_n6475), .Y(AES_CORE_DATAPATH__abc_16259_n6477) );
  AND2X2 AND2X2_2002 ( .A(AES_CORE_DATAPATH__abc_16259_n6480), .B(AES_CORE_DATAPATH__abc_16259_n6481), .Y(AES_CORE_DATAPATH__abc_16259_n6482) );
  AND2X2 AND2X2_2003 ( .A(AES_CORE_DATAPATH__abc_16259_n6474), .B(AES_CORE_DATAPATH__abc_16259_n6484), .Y(AES_CORE_DATAPATH__abc_16259_n6485) );
  AND2X2 AND2X2_2004 ( .A(AES_CORE_DATAPATH__abc_16259_n6487), .B(AES_CORE_DATAPATH__abc_16259_n6092_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6488) );
  AND2X2 AND2X2_2005 ( .A(AES_CORE_DATAPATH__abc_16259_n6486), .B(AES_CORE_DATAPATH__abc_16259_n6488), .Y(AES_CORE_DATAPATH__abc_16259_n6489) );
  AND2X2 AND2X2_2006 ( .A(AES_CORE_DATAPATH__abc_16259_n6491), .B(AES_CORE_CONTROL_UNIT_mode_cbc_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6492) );
  AND2X2 AND2X2_2007 ( .A(AES_CORE_DATAPATH__abc_16259_n6490), .B(AES_CORE_DATAPATH__abc_16259_n6492), .Y(AES_CORE_DATAPATH__abc_16259_n6493) );
  AND2X2 AND2X2_2008 ( .A(AES_CORE_DATAPATH__abc_16259_n6101_bF_buf1), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_8_), .Y(AES_CORE_DATAPATH__abc_16259_n6494) );
  AND2X2 AND2X2_2009 ( .A(AES_CORE_DATAPATH__abc_16259_n6496), .B(AES_CORE_DATAPATH__abc_16259_n6056_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6497) );
  AND2X2 AND2X2_201 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf4), .B(AES_CORE_DATAPATH_iv_3__18_), .Y(AES_CORE_DATAPATH__abc_16259_n2651_1) );
  AND2X2 AND2X2_2010 ( .A(AES_CORE_DATAPATH__abc_16259_n3189), .B(AES_CORE_DATAPATH__abc_16259_n6053_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6498) );
  AND2X2 AND2X2_2011 ( .A(AES_CORE_DATAPATH__abc_16259_n6500), .B(AES_CORE_DATAPATH__abc_16259_n6501), .Y(AES_CORE_DATAPATH__abc_16259_n6502) );
  AND2X2 AND2X2_2012 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n6502), .Y(AES_CORE_DATAPATH__abc_16259_n6503) );
  AND2X2 AND2X2_2013 ( .A(AES_CORE_DATAPATH__abc_16259_n6504), .B(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6505) );
  AND2X2 AND2X2_2014 ( .A(AES_CORE_DATAPATH__abc_16259_n6044_bF_buf0), .B(AES_CORE_DATAPATH_col_0__9_), .Y(AES_CORE_DATAPATH__abc_16259_n6507) );
  AND2X2 AND2X2_2015 ( .A(AES_CORE_DATAPATH__abc_16259_n3229), .B(AES_CORE_DATAPATH__abc_16259_n6059_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6508) );
  AND2X2 AND2X2_2016 ( .A(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf2), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_9_), .Y(AES_CORE_DATAPATH__abc_16259_n6509) );
  AND2X2 AND2X2_2017 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf6), .B(AES_CORE_DATAPATH_bkp_0__9_), .Y(AES_CORE_DATAPATH__abc_16259_n6511) );
  AND2X2 AND2X2_2018 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf5), .B(AES_CORE_DATAPATH_bkp_1__9_), .Y(AES_CORE_DATAPATH__abc_16259_n6512) );
  AND2X2 AND2X2_2019 ( .A(AES_CORE_DATAPATH__abc_16259_n6515), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n6516) );
  AND2X2 AND2X2_202 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf4), .B(AES_CORE_DATAPATH_iv_0__19_), .Y(AES_CORE_DATAPATH__abc_16259_n2653_1) );
  AND2X2 AND2X2_2020 ( .A(AES_CORE_DATAPATH__abc_16259_n6514), .B(AES_CORE_DATAPATH__abc_16259_n6516), .Y(AES_CORE_DATAPATH__abc_16259_n6517) );
  AND2X2 AND2X2_2021 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf5), .B(AES_CORE_DATAPATH_bkp_3__9_), .Y(AES_CORE_DATAPATH__abc_16259_n6518) );
  AND2X2 AND2X2_2022 ( .A(AES_CORE_DATAPATH__abc_16259_n6520), .B(AES_CORE_DATAPATH__abc_16259_n6521), .Y(AES_CORE_DATAPATH__abc_16259_n6522) );
  AND2X2 AND2X2_2023 ( .A(AES_CORE_DATAPATH__abc_16259_n3220), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n6525) );
  AND2X2 AND2X2_2024 ( .A(AES_CORE_DATAPATH__abc_16259_n6525), .B(AES_CORE_DATAPATH__abc_16259_n6524), .Y(AES_CORE_DATAPATH__abc_16259_n6526) );
  AND2X2 AND2X2_2025 ( .A(AES_CORE_DATAPATH__abc_16259_n6529), .B(AES_CORE_DATAPATH__abc_16259_n6530), .Y(AES_CORE_DATAPATH__abc_16259_n6531) );
  AND2X2 AND2X2_2026 ( .A(AES_CORE_DATAPATH__abc_16259_n6523), .B(AES_CORE_DATAPATH__abc_16259_n6533), .Y(AES_CORE_DATAPATH__abc_16259_n6534) );
  AND2X2 AND2X2_2027 ( .A(AES_CORE_DATAPATH__abc_16259_n6536), .B(AES_CORE_DATAPATH__abc_16259_n6092_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n6537) );
  AND2X2 AND2X2_2028 ( .A(AES_CORE_DATAPATH__abc_16259_n6535), .B(AES_CORE_DATAPATH__abc_16259_n6537), .Y(AES_CORE_DATAPATH__abc_16259_n6538) );
  AND2X2 AND2X2_2029 ( .A(AES_CORE_DATAPATH__abc_16259_n6540), .B(AES_CORE_CONTROL_UNIT_mode_cbc_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6541) );
  AND2X2 AND2X2_203 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf3), .B(AES_CORE_DATAPATH_iv_1__19_), .Y(AES_CORE_DATAPATH__abc_16259_n2654_1) );
  AND2X2 AND2X2_2030 ( .A(AES_CORE_DATAPATH__abc_16259_n6539), .B(AES_CORE_DATAPATH__abc_16259_n6541), .Y(AES_CORE_DATAPATH__abc_16259_n6542) );
  AND2X2 AND2X2_2031 ( .A(AES_CORE_DATAPATH__abc_16259_n6101_bF_buf0), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_9_), .Y(AES_CORE_DATAPATH__abc_16259_n6543) );
  AND2X2 AND2X2_2032 ( .A(AES_CORE_DATAPATH__abc_16259_n6545), .B(AES_CORE_DATAPATH__abc_16259_n6056_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n6546) );
  AND2X2 AND2X2_2033 ( .A(AES_CORE_DATAPATH__abc_16259_n3229), .B(AES_CORE_DATAPATH__abc_16259_n6053_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n6547) );
  AND2X2 AND2X2_2034 ( .A(AES_CORE_DATAPATH__abc_16259_n6549), .B(AES_CORE_DATAPATH__abc_16259_n6550), .Y(AES_CORE_DATAPATH__abc_16259_n6551) );
  AND2X2 AND2X2_2035 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n6551), .Y(AES_CORE_DATAPATH__abc_16259_n6552) );
  AND2X2 AND2X2_2036 ( .A(AES_CORE_DATAPATH__abc_16259_n6553), .B(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n6554) );
  AND2X2 AND2X2_2037 ( .A(AES_CORE_DATAPATH__abc_16259_n3260), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6558) );
  AND2X2 AND2X2_2038 ( .A(AES_CORE_DATAPATH__abc_16259_n6558), .B(AES_CORE_DATAPATH__abc_16259_n6557), .Y(AES_CORE_DATAPATH__abc_16259_n6559) );
  AND2X2 AND2X2_2039 ( .A(AES_CORE_DATAPATH__abc_16259_n6561), .B(AES_CORE_DATAPATH__abc_16259_n6059_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n6562) );
  AND2X2 AND2X2_204 ( .A(AES_CORE_DATAPATH__abc_16259_n2657), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n2658_1) );
  AND2X2 AND2X2_2040 ( .A(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n6563), .Y(AES_CORE_DATAPATH__abc_16259_n6564) );
  AND2X2 AND2X2_2041 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf5), .B(AES_CORE_DATAPATH_bkp_0__10_), .Y(AES_CORE_DATAPATH__abc_16259_n6566) );
  AND2X2 AND2X2_2042 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf4), .B(AES_CORE_DATAPATH_bkp_1__10_), .Y(AES_CORE_DATAPATH__abc_16259_n6567) );
  AND2X2 AND2X2_2043 ( .A(AES_CORE_DATAPATH__abc_16259_n6570), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n6571) );
  AND2X2 AND2X2_2044 ( .A(AES_CORE_DATAPATH__abc_16259_n6569), .B(AES_CORE_DATAPATH__abc_16259_n6571), .Y(AES_CORE_DATAPATH__abc_16259_n6572) );
  AND2X2 AND2X2_2045 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf4), .B(AES_CORE_DATAPATH_bkp_3__10_), .Y(AES_CORE_DATAPATH__abc_16259_n6573) );
  AND2X2 AND2X2_2046 ( .A(AES_CORE_DATAPATH__abc_16259_n6576), .B(AES_CORE_DATAPATH__abc_16259_n6575), .Y(AES_CORE_DATAPATH__abc_16259_n6577) );
  AND2X2 AND2X2_2047 ( .A(AES_CORE_DATAPATH__abc_16259_n6579), .B(AES_CORE_DATAPATH__abc_16259_n6580), .Y(AES_CORE_DATAPATH__abc_16259_n6581) );
  AND2X2 AND2X2_2048 ( .A(AES_CORE_DATAPATH__abc_16259_n6578), .B(AES_CORE_DATAPATH__abc_16259_n6583), .Y(AES_CORE_DATAPATH__abc_16259_n6584) );
  AND2X2 AND2X2_2049 ( .A(AES_CORE_DATAPATH__abc_16259_n6584), .B(AES_CORE_CONTROL_UNIT_last_round_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6585) );
  AND2X2 AND2X2_205 ( .A(AES_CORE_DATAPATH__abc_16259_n2656_1), .B(AES_CORE_DATAPATH__abc_16259_n2658_1), .Y(AES_CORE_DATAPATH__abc_16259_n2659) );
  AND2X2 AND2X2_2050 ( .A(AES_CORE_DATAPATH__abc_16259_n6587), .B(AES_CORE_DATAPATH__abc_16259_n6057_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6588) );
  AND2X2 AND2X2_2051 ( .A(AES_CORE_DATAPATH__abc_16259_n6584), .B(AES_CORE_DATAPATH__abc_16259_n6097_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6591) );
  AND2X2 AND2X2_2052 ( .A(AES_CORE_DATAPATH__abc_16259_n6095_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n6563), .Y(AES_CORE_DATAPATH__abc_16259_n6592) );
  AND2X2 AND2X2_2053 ( .A(AES_CORE_DATAPATH__abc_16259_n6594), .B(AES_CORE_DATAPATH__abc_16259_n6596), .Y(AES_CORE_DATAPATH__abc_16259_n6597) );
  AND2X2 AND2X2_2054 ( .A(AES_CORE_DATAPATH__abc_16259_n6597), .B(AES_CORE_DATAPATH__abc_16259_n6590), .Y(AES_CORE_DATAPATH__abc_16259_n6598) );
  AND2X2 AND2X2_2055 ( .A(AES_CORE_DATAPATH__abc_16259_n6599), .B(AES_CORE_DATAPATH__abc_16259_n6601), .Y(AES_CORE_DATAPATH__abc_16259_n6602) );
  AND2X2 AND2X2_2056 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf3), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_42_), .Y(AES_CORE_DATAPATH__abc_16259_n6606) );
  AND2X2 AND2X2_2057 ( .A(AES_CORE_DATAPATH__abc_16259_n6605), .B(AES_CORE_DATAPATH__abc_16259_n6607), .Y(AES_CORE_DATAPATH__abc_16259_n6608) );
  AND2X2 AND2X2_2058 ( .A(AES_CORE_DATAPATH__abc_16259_n6602), .B(AES_CORE_DATAPATH__abc_16259_n6609), .Y(AES_CORE_DATAPATH__abc_16259_n6610) );
  AND2X2 AND2X2_2059 ( .A(AES_CORE_DATAPATH__abc_16259_n6610), .B(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n6611) );
  AND2X2 AND2X2_206 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf3), .B(AES_CORE_DATAPATH_iv_3__19_), .Y(AES_CORE_DATAPATH__abc_16259_n2660) );
  AND2X2 AND2X2_2060 ( .A(AES_CORE_DATAPATH__abc_16259_n6612), .B(AES_CORE_DATAPATH__abc_16259_n6613), .Y(AES_CORE_DATAPATH__0col_0__31_0__10_) );
  AND2X2 AND2X2_2061 ( .A(AES_CORE_DATAPATH__abc_16259_n3300), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6616) );
  AND2X2 AND2X2_2062 ( .A(AES_CORE_DATAPATH__abc_16259_n6616), .B(AES_CORE_DATAPATH__abc_16259_n6615), .Y(AES_CORE_DATAPATH__abc_16259_n6617) );
  AND2X2 AND2X2_2063 ( .A(AES_CORE_DATAPATH__abc_16259_n6619), .B(AES_CORE_DATAPATH__abc_16259_n6059_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n6620) );
  AND2X2 AND2X2_2064 ( .A(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf5), .B(AES_CORE_DATAPATH__abc_16259_n6621), .Y(AES_CORE_DATAPATH__abc_16259_n6622) );
  AND2X2 AND2X2_2065 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf4), .B(AES_CORE_DATAPATH_bkp_0__11_), .Y(AES_CORE_DATAPATH__abc_16259_n6624) );
  AND2X2 AND2X2_2066 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1__11_), .Y(AES_CORE_DATAPATH__abc_16259_n6625) );
  AND2X2 AND2X2_2067 ( .A(AES_CORE_DATAPATH__abc_16259_n6628), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6629) );
  AND2X2 AND2X2_2068 ( .A(AES_CORE_DATAPATH__abc_16259_n6627), .B(AES_CORE_DATAPATH__abc_16259_n6629), .Y(AES_CORE_DATAPATH__abc_16259_n6630) );
  AND2X2 AND2X2_2069 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf3), .B(AES_CORE_DATAPATH_bkp_3__11_), .Y(AES_CORE_DATAPATH__abc_16259_n6631) );
  AND2X2 AND2X2_207 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf3), .B(AES_CORE_DATAPATH_iv_0__20_), .Y(AES_CORE_DATAPATH__abc_16259_n2662) );
  AND2X2 AND2X2_2070 ( .A(AES_CORE_DATAPATH__abc_16259_n6633), .B(AES_CORE_DATAPATH__abc_16259_n6634), .Y(AES_CORE_DATAPATH__abc_16259_n6635) );
  AND2X2 AND2X2_2071 ( .A(AES_CORE_DATAPATH__abc_16259_n6637), .B(AES_CORE_DATAPATH__abc_16259_n6638), .Y(AES_CORE_DATAPATH__abc_16259_n6639) );
  AND2X2 AND2X2_2072 ( .A(AES_CORE_DATAPATH__abc_16259_n6636), .B(AES_CORE_DATAPATH__abc_16259_n6641), .Y(AES_CORE_DATAPATH__abc_16259_n6642) );
  AND2X2 AND2X2_2073 ( .A(AES_CORE_DATAPATH__abc_16259_n6642), .B(AES_CORE_CONTROL_UNIT_last_round_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6643) );
  AND2X2 AND2X2_2074 ( .A(AES_CORE_DATAPATH__abc_16259_n6644), .B(AES_CORE_DATAPATH__abc_16259_n6057_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6645) );
  AND2X2 AND2X2_2075 ( .A(AES_CORE_DATAPATH__abc_16259_n6642), .B(AES_CORE_DATAPATH__abc_16259_n6097_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6648) );
  AND2X2 AND2X2_2076 ( .A(AES_CORE_DATAPATH__abc_16259_n6095_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n6621), .Y(AES_CORE_DATAPATH__abc_16259_n6649) );
  AND2X2 AND2X2_2077 ( .A(AES_CORE_DATAPATH__abc_16259_n6651), .B(AES_CORE_DATAPATH__abc_16259_n6652), .Y(AES_CORE_DATAPATH__abc_16259_n6653) );
  AND2X2 AND2X2_2078 ( .A(AES_CORE_DATAPATH__abc_16259_n6653), .B(AES_CORE_DATAPATH__abc_16259_n6647), .Y(AES_CORE_DATAPATH__abc_16259_n6654) );
  AND2X2 AND2X2_2079 ( .A(AES_CORE_DATAPATH__abc_16259_n6655), .B(AES_CORE_DATAPATH__abc_16259_n6656), .Y(AES_CORE_DATAPATH__abc_16259_n6657) );
  AND2X2 AND2X2_208 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf2), .B(AES_CORE_DATAPATH_iv_1__20_), .Y(AES_CORE_DATAPATH__abc_16259_n2663_1) );
  AND2X2 AND2X2_2080 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf1), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_43_), .Y(AES_CORE_DATAPATH__abc_16259_n6660) );
  AND2X2 AND2X2_2081 ( .A(AES_CORE_DATAPATH__abc_16259_n6659), .B(AES_CORE_DATAPATH__abc_16259_n6661), .Y(AES_CORE_DATAPATH__abc_16259_n6662) );
  AND2X2 AND2X2_2082 ( .A(AES_CORE_DATAPATH__abc_16259_n6657), .B(AES_CORE_DATAPATH__abc_16259_n6663), .Y(AES_CORE_DATAPATH__abc_16259_n6664) );
  AND2X2 AND2X2_2083 ( .A(AES_CORE_DATAPATH__abc_16259_n6664), .B(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6665) );
  AND2X2 AND2X2_2084 ( .A(AES_CORE_DATAPATH__abc_16259_n6666), .B(AES_CORE_DATAPATH__abc_16259_n6667), .Y(AES_CORE_DATAPATH__0col_0__31_0__11_) );
  AND2X2 AND2X2_2085 ( .A(AES_CORE_DATAPATH__abc_16259_n6044_bF_buf4), .B(AES_CORE_DATAPATH_col_0__12_), .Y(AES_CORE_DATAPATH__abc_16259_n6669) );
  AND2X2 AND2X2_2086 ( .A(AES_CORE_DATAPATH__abc_16259_n3349), .B(AES_CORE_DATAPATH__abc_16259_n6059_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6670) );
  AND2X2 AND2X2_2087 ( .A(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf3), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_12_), .Y(AES_CORE_DATAPATH__abc_16259_n6671) );
  AND2X2 AND2X2_2088 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf3), .B(AES_CORE_DATAPATH_bkp_0__12_), .Y(AES_CORE_DATAPATH__abc_16259_n6673) );
  AND2X2 AND2X2_2089 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf2), .B(AES_CORE_DATAPATH_bkp_1__12_), .Y(AES_CORE_DATAPATH__abc_16259_n6674) );
  AND2X2 AND2X2_209 ( .A(AES_CORE_DATAPATH__abc_16259_n2666), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n2667_1) );
  AND2X2 AND2X2_2090 ( .A(AES_CORE_DATAPATH__abc_16259_n6677), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6678) );
  AND2X2 AND2X2_2091 ( .A(AES_CORE_DATAPATH__abc_16259_n6676), .B(AES_CORE_DATAPATH__abc_16259_n6678), .Y(AES_CORE_DATAPATH__abc_16259_n6679) );
  AND2X2 AND2X2_2092 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf2), .B(AES_CORE_DATAPATH_bkp_3__12_), .Y(AES_CORE_DATAPATH__abc_16259_n6680) );
  AND2X2 AND2X2_2093 ( .A(AES_CORE_DATAPATH__abc_16259_n6682), .B(AES_CORE_DATAPATH__abc_16259_n6683), .Y(AES_CORE_DATAPATH__abc_16259_n6684) );
  AND2X2 AND2X2_2094 ( .A(AES_CORE_DATAPATH__abc_16259_n3340), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6687) );
  AND2X2 AND2X2_2095 ( .A(AES_CORE_DATAPATH__abc_16259_n6687), .B(AES_CORE_DATAPATH__abc_16259_n6686), .Y(AES_CORE_DATAPATH__abc_16259_n6688) );
  AND2X2 AND2X2_2096 ( .A(AES_CORE_DATAPATH__abc_16259_n6691), .B(AES_CORE_DATAPATH__abc_16259_n6692), .Y(AES_CORE_DATAPATH__abc_16259_n6693) );
  AND2X2 AND2X2_2097 ( .A(AES_CORE_DATAPATH__abc_16259_n6685), .B(AES_CORE_DATAPATH__abc_16259_n6695), .Y(AES_CORE_DATAPATH__abc_16259_n6696) );
  AND2X2 AND2X2_2098 ( .A(AES_CORE_DATAPATH__abc_16259_n6698), .B(AES_CORE_DATAPATH__abc_16259_n6092_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6699) );
  AND2X2 AND2X2_2099 ( .A(AES_CORE_DATAPATH__abc_16259_n6697), .B(AES_CORE_DATAPATH__abc_16259_n6699), .Y(AES_CORE_DATAPATH__abc_16259_n6700) );
  AND2X2 AND2X2_21 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n97), .B(AES_CORE_CONTROL_UNIT__abc_15841_n84_1), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n98) );
  AND2X2 AND2X2_210 ( .A(AES_CORE_DATAPATH__abc_16259_n2665_1), .B(AES_CORE_DATAPATH__abc_16259_n2667_1), .Y(AES_CORE_DATAPATH__abc_16259_n2668) );
  AND2X2 AND2X2_2100 ( .A(AES_CORE_DATAPATH__abc_16259_n6702), .B(AES_CORE_CONTROL_UNIT_mode_cbc_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6703) );
  AND2X2 AND2X2_2101 ( .A(AES_CORE_DATAPATH__abc_16259_n6701), .B(AES_CORE_DATAPATH__abc_16259_n6703), .Y(AES_CORE_DATAPATH__abc_16259_n6704) );
  AND2X2 AND2X2_2102 ( .A(AES_CORE_DATAPATH__abc_16259_n6101_bF_buf3), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_12_), .Y(AES_CORE_DATAPATH__abc_16259_n6705) );
  AND2X2 AND2X2_2103 ( .A(AES_CORE_DATAPATH__abc_16259_n6707), .B(AES_CORE_DATAPATH__abc_16259_n6056_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6708) );
  AND2X2 AND2X2_2104 ( .A(AES_CORE_DATAPATH__abc_16259_n3349), .B(AES_CORE_DATAPATH__abc_16259_n6053_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6709) );
  AND2X2 AND2X2_2105 ( .A(AES_CORE_DATAPATH__abc_16259_n6711), .B(AES_CORE_DATAPATH__abc_16259_n6712), .Y(AES_CORE_DATAPATH__abc_16259_n6713) );
  AND2X2 AND2X2_2106 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf8), .B(AES_CORE_DATAPATH__abc_16259_n6713), .Y(AES_CORE_DATAPATH__abc_16259_n6714) );
  AND2X2 AND2X2_2107 ( .A(AES_CORE_DATAPATH__abc_16259_n6715), .B(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6716) );
  AND2X2 AND2X2_2108 ( .A(AES_CORE_DATAPATH__abc_16259_n3380_1), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6719) );
  AND2X2 AND2X2_2109 ( .A(AES_CORE_DATAPATH__abc_16259_n6719), .B(AES_CORE_DATAPATH__abc_16259_n6718), .Y(AES_CORE_DATAPATH__abc_16259_n6720) );
  AND2X2 AND2X2_211 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf2), .B(AES_CORE_DATAPATH_iv_3__20_), .Y(AES_CORE_DATAPATH__abc_16259_n2669_1) );
  AND2X2 AND2X2_2110 ( .A(AES_CORE_DATAPATH__abc_16259_n6722), .B(AES_CORE_DATAPATH__abc_16259_n6059_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6723) );
  AND2X2 AND2X2_2111 ( .A(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n6724), .Y(AES_CORE_DATAPATH__abc_16259_n6725) );
  AND2X2 AND2X2_2112 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf2), .B(AES_CORE_DATAPATH_bkp_0__13_), .Y(AES_CORE_DATAPATH__abc_16259_n6727) );
  AND2X2 AND2X2_2113 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf1), .B(AES_CORE_DATAPATH_bkp_1__13_), .Y(AES_CORE_DATAPATH__abc_16259_n6728) );
  AND2X2 AND2X2_2114 ( .A(AES_CORE_DATAPATH__abc_16259_n6731), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6732) );
  AND2X2 AND2X2_2115 ( .A(AES_CORE_DATAPATH__abc_16259_n6730), .B(AES_CORE_DATAPATH__abc_16259_n6732), .Y(AES_CORE_DATAPATH__abc_16259_n6733) );
  AND2X2 AND2X2_2116 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf1), .B(AES_CORE_DATAPATH_bkp_3__13_), .Y(AES_CORE_DATAPATH__abc_16259_n6734) );
  AND2X2 AND2X2_2117 ( .A(AES_CORE_DATAPATH__abc_16259_n6736), .B(AES_CORE_DATAPATH__abc_16259_n6737), .Y(AES_CORE_DATAPATH__abc_16259_n6738) );
  AND2X2 AND2X2_2118 ( .A(AES_CORE_DATAPATH__abc_16259_n6740), .B(AES_CORE_DATAPATH__abc_16259_n6741), .Y(AES_CORE_DATAPATH__abc_16259_n6742) );
  AND2X2 AND2X2_2119 ( .A(AES_CORE_DATAPATH__abc_16259_n6739), .B(AES_CORE_DATAPATH__abc_16259_n6744), .Y(AES_CORE_DATAPATH__abc_16259_n6745) );
  AND2X2 AND2X2_212 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf2), .B(AES_CORE_DATAPATH_iv_0__21_), .Y(AES_CORE_DATAPATH__abc_16259_n2671_1) );
  AND2X2 AND2X2_2120 ( .A(AES_CORE_DATAPATH__abc_16259_n6745), .B(AES_CORE_CONTROL_UNIT_last_round_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6746) );
  AND2X2 AND2X2_2121 ( .A(AES_CORE_DATAPATH__abc_16259_n6747), .B(AES_CORE_DATAPATH__abc_16259_n6057_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n6748) );
  AND2X2 AND2X2_2122 ( .A(AES_CORE_DATAPATH__abc_16259_n6745), .B(AES_CORE_DATAPATH__abc_16259_n6097_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6751) );
  AND2X2 AND2X2_2123 ( .A(AES_CORE_DATAPATH__abc_16259_n6095_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n6724), .Y(AES_CORE_DATAPATH__abc_16259_n6752) );
  AND2X2 AND2X2_2124 ( .A(AES_CORE_DATAPATH__abc_16259_n6754), .B(AES_CORE_DATAPATH__abc_16259_n6755), .Y(AES_CORE_DATAPATH__abc_16259_n6756) );
  AND2X2 AND2X2_2125 ( .A(AES_CORE_DATAPATH__abc_16259_n6756), .B(AES_CORE_DATAPATH__abc_16259_n6750), .Y(AES_CORE_DATAPATH__abc_16259_n6757) );
  AND2X2 AND2X2_2126 ( .A(AES_CORE_DATAPATH__abc_16259_n6758), .B(AES_CORE_DATAPATH__abc_16259_n6759), .Y(AES_CORE_DATAPATH__abc_16259_n6760) );
  AND2X2 AND2X2_2127 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf13), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_45_), .Y(AES_CORE_DATAPATH__abc_16259_n6763) );
  AND2X2 AND2X2_2128 ( .A(AES_CORE_DATAPATH__abc_16259_n6762), .B(AES_CORE_DATAPATH__abc_16259_n6764), .Y(AES_CORE_DATAPATH__abc_16259_n6765) );
  AND2X2 AND2X2_2129 ( .A(AES_CORE_DATAPATH__abc_16259_n6760), .B(AES_CORE_DATAPATH__abc_16259_n6766), .Y(AES_CORE_DATAPATH__abc_16259_n6767) );
  AND2X2 AND2X2_213 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf1), .B(AES_CORE_DATAPATH_iv_1__21_), .Y(AES_CORE_DATAPATH__abc_16259_n2672) );
  AND2X2 AND2X2_2130 ( .A(AES_CORE_DATAPATH__abc_16259_n6767), .B(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n6768) );
  AND2X2 AND2X2_2131 ( .A(AES_CORE_DATAPATH__abc_16259_n6769), .B(AES_CORE_DATAPATH__abc_16259_n6770), .Y(AES_CORE_DATAPATH__0col_0__31_0__13_) );
  AND2X2 AND2X2_2132 ( .A(AES_CORE_DATAPATH__abc_16259_n6044_bF_buf3), .B(AES_CORE_DATAPATH_col_0__14_), .Y(AES_CORE_DATAPATH__abc_16259_n6772) );
  AND2X2 AND2X2_2133 ( .A(AES_CORE_DATAPATH__abc_16259_n3429), .B(AES_CORE_DATAPATH__abc_16259_n6059_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6773) );
  AND2X2 AND2X2_2134 ( .A(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf6), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_14_), .Y(AES_CORE_DATAPATH__abc_16259_n6774) );
  AND2X2 AND2X2_2135 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf1), .B(AES_CORE_DATAPATH_bkp_0__14_), .Y(AES_CORE_DATAPATH__abc_16259_n6776) );
  AND2X2 AND2X2_2136 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf0), .B(AES_CORE_DATAPATH_bkp_1__14_), .Y(AES_CORE_DATAPATH__abc_16259_n6777) );
  AND2X2 AND2X2_2137 ( .A(AES_CORE_DATAPATH__abc_16259_n6780), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6781) );
  AND2X2 AND2X2_2138 ( .A(AES_CORE_DATAPATH__abc_16259_n6779), .B(AES_CORE_DATAPATH__abc_16259_n6781), .Y(AES_CORE_DATAPATH__abc_16259_n6782) );
  AND2X2 AND2X2_2139 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf0), .B(AES_CORE_DATAPATH_bkp_3__14_), .Y(AES_CORE_DATAPATH__abc_16259_n6783) );
  AND2X2 AND2X2_214 ( .A(AES_CORE_DATAPATH__abc_16259_n2675_1), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n2676) );
  AND2X2 AND2X2_2140 ( .A(AES_CORE_DATAPATH__abc_16259_n6785), .B(AES_CORE_DATAPATH__abc_16259_n6786), .Y(AES_CORE_DATAPATH__abc_16259_n6787) );
  AND2X2 AND2X2_2141 ( .A(AES_CORE_DATAPATH__abc_16259_n3420), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n6790) );
  AND2X2 AND2X2_2142 ( .A(AES_CORE_DATAPATH__abc_16259_n6790), .B(AES_CORE_DATAPATH__abc_16259_n6789), .Y(AES_CORE_DATAPATH__abc_16259_n6791) );
  AND2X2 AND2X2_2143 ( .A(AES_CORE_DATAPATH__abc_16259_n6794), .B(AES_CORE_DATAPATH__abc_16259_n6795), .Y(AES_CORE_DATAPATH__abc_16259_n6796) );
  AND2X2 AND2X2_2144 ( .A(AES_CORE_DATAPATH__abc_16259_n6788), .B(AES_CORE_DATAPATH__abc_16259_n6798), .Y(AES_CORE_DATAPATH__abc_16259_n6799) );
  AND2X2 AND2X2_2145 ( .A(AES_CORE_DATAPATH__abc_16259_n6801), .B(AES_CORE_DATAPATH__abc_16259_n6092_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6802) );
  AND2X2 AND2X2_2146 ( .A(AES_CORE_DATAPATH__abc_16259_n6800), .B(AES_CORE_DATAPATH__abc_16259_n6802), .Y(AES_CORE_DATAPATH__abc_16259_n6803) );
  AND2X2 AND2X2_2147 ( .A(AES_CORE_DATAPATH__abc_16259_n6805), .B(AES_CORE_CONTROL_UNIT_mode_cbc_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6806) );
  AND2X2 AND2X2_2148 ( .A(AES_CORE_DATAPATH__abc_16259_n6804), .B(AES_CORE_DATAPATH__abc_16259_n6806), .Y(AES_CORE_DATAPATH__abc_16259_n6807) );
  AND2X2 AND2X2_2149 ( .A(AES_CORE_DATAPATH__abc_16259_n6101_bF_buf2), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_14_), .Y(AES_CORE_DATAPATH__abc_16259_n6808) );
  AND2X2 AND2X2_215 ( .A(AES_CORE_DATAPATH__abc_16259_n2674), .B(AES_CORE_DATAPATH__abc_16259_n2676), .Y(AES_CORE_DATAPATH__abc_16259_n2677_1) );
  AND2X2 AND2X2_2150 ( .A(AES_CORE_DATAPATH__abc_16259_n6810), .B(AES_CORE_DATAPATH__abc_16259_n6056_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6811) );
  AND2X2 AND2X2_2151 ( .A(AES_CORE_DATAPATH__abc_16259_n3429), .B(AES_CORE_DATAPATH__abc_16259_n6053_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6812) );
  AND2X2 AND2X2_2152 ( .A(AES_CORE_DATAPATH__abc_16259_n6814), .B(AES_CORE_DATAPATH__abc_16259_n6815), .Y(AES_CORE_DATAPATH__abc_16259_n6816) );
  AND2X2 AND2X2_2153 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf7), .B(AES_CORE_DATAPATH__abc_16259_n6816), .Y(AES_CORE_DATAPATH__abc_16259_n6817) );
  AND2X2 AND2X2_2154 ( .A(AES_CORE_DATAPATH__abc_16259_n6818), .B(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6819) );
  AND2X2 AND2X2_2155 ( .A(AES_CORE_DATAPATH__abc_16259_n3460_1), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n6822) );
  AND2X2 AND2X2_2156 ( .A(AES_CORE_DATAPATH__abc_16259_n6822), .B(AES_CORE_DATAPATH__abc_16259_n6821), .Y(AES_CORE_DATAPATH__abc_16259_n6823) );
  AND2X2 AND2X2_2157 ( .A(AES_CORE_DATAPATH__abc_16259_n6825), .B(AES_CORE_DATAPATH__abc_16259_n6059_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6826) );
  AND2X2 AND2X2_2158 ( .A(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n6827), .Y(AES_CORE_DATAPATH__abc_16259_n6828) );
  AND2X2 AND2X2_2159 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf0), .B(AES_CORE_DATAPATH_bkp_0__15_), .Y(AES_CORE_DATAPATH__abc_16259_n6830) );
  AND2X2 AND2X2_216 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf1), .B(AES_CORE_DATAPATH_iv_3__21_), .Y(AES_CORE_DATAPATH__abc_16259_n2678) );
  AND2X2 AND2X2_2160 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf7), .B(AES_CORE_DATAPATH_bkp_1__15_), .Y(AES_CORE_DATAPATH__abc_16259_n6831) );
  AND2X2 AND2X2_2161 ( .A(AES_CORE_DATAPATH__abc_16259_n6834), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n6835) );
  AND2X2 AND2X2_2162 ( .A(AES_CORE_DATAPATH__abc_16259_n6833), .B(AES_CORE_DATAPATH__abc_16259_n6835), .Y(AES_CORE_DATAPATH__abc_16259_n6836) );
  AND2X2 AND2X2_2163 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf7), .B(AES_CORE_DATAPATH_bkp_3__15_), .Y(AES_CORE_DATAPATH__abc_16259_n6837) );
  AND2X2 AND2X2_2164 ( .A(AES_CORE_DATAPATH__abc_16259_n6840), .B(AES_CORE_DATAPATH__abc_16259_n6839), .Y(AES_CORE_DATAPATH__abc_16259_n6841) );
  AND2X2 AND2X2_2165 ( .A(AES_CORE_DATAPATH__abc_16259_n6843), .B(AES_CORE_DATAPATH__abc_16259_n6844), .Y(AES_CORE_DATAPATH__abc_16259_n6845) );
  AND2X2 AND2X2_2166 ( .A(AES_CORE_DATAPATH__abc_16259_n6842), .B(AES_CORE_DATAPATH__abc_16259_n6847), .Y(AES_CORE_DATAPATH__abc_16259_n6848) );
  AND2X2 AND2X2_2167 ( .A(AES_CORE_DATAPATH__abc_16259_n6848), .B(AES_CORE_CONTROL_UNIT_last_round_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n6849) );
  AND2X2 AND2X2_2168 ( .A(AES_CORE_DATAPATH__abc_16259_n6850), .B(AES_CORE_DATAPATH__abc_16259_n6057_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6851) );
  AND2X2 AND2X2_2169 ( .A(AES_CORE_DATAPATH__abc_16259_n6848), .B(AES_CORE_DATAPATH__abc_16259_n6097_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6854) );
  AND2X2 AND2X2_217 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf1), .B(AES_CORE_DATAPATH_iv_0__22_), .Y(AES_CORE_DATAPATH__abc_16259_n2680) );
  AND2X2 AND2X2_2170 ( .A(AES_CORE_DATAPATH__abc_16259_n6095_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n6827), .Y(AES_CORE_DATAPATH__abc_16259_n6855) );
  AND2X2 AND2X2_2171 ( .A(AES_CORE_DATAPATH__abc_16259_n6857), .B(AES_CORE_DATAPATH__abc_16259_n6858), .Y(AES_CORE_DATAPATH__abc_16259_n6859) );
  AND2X2 AND2X2_2172 ( .A(AES_CORE_DATAPATH__abc_16259_n6859), .B(AES_CORE_DATAPATH__abc_16259_n6853), .Y(AES_CORE_DATAPATH__abc_16259_n6860) );
  AND2X2 AND2X2_2173 ( .A(AES_CORE_DATAPATH__abc_16259_n6861), .B(AES_CORE_DATAPATH__abc_16259_n6862), .Y(AES_CORE_DATAPATH__abc_16259_n6863) );
  AND2X2 AND2X2_2174 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf10), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_47_), .Y(AES_CORE_DATAPATH__abc_16259_n6866) );
  AND2X2 AND2X2_2175 ( .A(AES_CORE_DATAPATH__abc_16259_n6865), .B(AES_CORE_DATAPATH__abc_16259_n6867), .Y(AES_CORE_DATAPATH__abc_16259_n6868) );
  AND2X2 AND2X2_2176 ( .A(AES_CORE_DATAPATH__abc_16259_n6863), .B(AES_CORE_DATAPATH__abc_16259_n6869), .Y(AES_CORE_DATAPATH__abc_16259_n6870) );
  AND2X2 AND2X2_2177 ( .A(AES_CORE_DATAPATH__abc_16259_n6870), .B(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6871) );
  AND2X2 AND2X2_2178 ( .A(AES_CORE_DATAPATH__abc_16259_n6872), .B(AES_CORE_DATAPATH__abc_16259_n6873), .Y(AES_CORE_DATAPATH__0col_0__31_0__15_) );
  AND2X2 AND2X2_2179 ( .A(AES_CORE_DATAPATH__abc_16259_n6044_bF_buf2), .B(AES_CORE_DATAPATH_col_0__16_), .Y(AES_CORE_DATAPATH__abc_16259_n6875) );
  AND2X2 AND2X2_218 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf0), .B(AES_CORE_DATAPATH_iv_1__22_), .Y(AES_CORE_DATAPATH__abc_16259_n2681_1) );
  AND2X2 AND2X2_2180 ( .A(AES_CORE_DATAPATH__abc_16259_n3500_1), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n6877) );
  AND2X2 AND2X2_2181 ( .A(AES_CORE_DATAPATH__abc_16259_n6877), .B(AES_CORE_DATAPATH__abc_16259_n6876), .Y(AES_CORE_DATAPATH__abc_16259_n6878) );
  AND2X2 AND2X2_2182 ( .A(AES_CORE_DATAPATH__abc_16259_n6880), .B(AES_CORE_DATAPATH__abc_16259_n6059_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n6881) );
  AND2X2 AND2X2_2183 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf7), .B(AES_CORE_DATAPATH_bkp_0__16_), .Y(AES_CORE_DATAPATH__abc_16259_n6885) );
  AND2X2 AND2X2_2184 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf6), .B(AES_CORE_DATAPATH_bkp_1__16_), .Y(AES_CORE_DATAPATH__abc_16259_n6886) );
  AND2X2 AND2X2_2185 ( .A(AES_CORE_DATAPATH__abc_16259_n6889), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n6890) );
  AND2X2 AND2X2_2186 ( .A(AES_CORE_DATAPATH__abc_16259_n6888), .B(AES_CORE_DATAPATH__abc_16259_n6890), .Y(AES_CORE_DATAPATH__abc_16259_n6891) );
  AND2X2 AND2X2_2187 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf6), .B(AES_CORE_DATAPATH_bkp_3__16_), .Y(AES_CORE_DATAPATH__abc_16259_n6892) );
  AND2X2 AND2X2_2188 ( .A(AES_CORE_DATAPATH__abc_16259_n6894), .B(AES_CORE_DATAPATH__abc_16259_n6895), .Y(AES_CORE_DATAPATH__abc_16259_n6896) );
  AND2X2 AND2X2_2189 ( .A(AES_CORE_DATAPATH__abc_16259_n6899), .B(AES_CORE_DATAPATH__abc_16259_n6882), .Y(AES_CORE_DATAPATH__abc_16259_n6900) );
  AND2X2 AND2X2_219 ( .A(AES_CORE_DATAPATH__abc_16259_n2684), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n2685_1) );
  AND2X2 AND2X2_2190 ( .A(AES_CORE_DATAPATH__abc_16259_n6898), .B(AES_CORE_DATAPATH__abc_16259_n6901), .Y(AES_CORE_DATAPATH__abc_16259_n6902) );
  AND2X2 AND2X2_2191 ( .A(AES_CORE_DATAPATH__abc_16259_n6904), .B(AES_CORE_DATAPATH__abc_16259_n6092_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6905) );
  AND2X2 AND2X2_2192 ( .A(AES_CORE_DATAPATH__abc_16259_n6903), .B(AES_CORE_DATAPATH__abc_16259_n6905), .Y(AES_CORE_DATAPATH__abc_16259_n6906) );
  AND2X2 AND2X2_2193 ( .A(AES_CORE_DATAPATH__abc_16259_n6908), .B(AES_CORE_CONTROL_UNIT_mode_cbc_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n6909) );
  AND2X2 AND2X2_2194 ( .A(AES_CORE_DATAPATH__abc_16259_n6907), .B(AES_CORE_DATAPATH__abc_16259_n6909), .Y(AES_CORE_DATAPATH__abc_16259_n6910) );
  AND2X2 AND2X2_2195 ( .A(AES_CORE_DATAPATH__abc_16259_n6101_bF_buf1), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_16_), .Y(AES_CORE_DATAPATH__abc_16259_n6911) );
  AND2X2 AND2X2_2196 ( .A(AES_CORE_DATAPATH__abc_16259_n6913), .B(AES_CORE_DATAPATH__abc_16259_n6056_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6914) );
  AND2X2 AND2X2_2197 ( .A(AES_CORE_DATAPATH__abc_16259_n3509), .B(AES_CORE_DATAPATH__abc_16259_n6053_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6915) );
  AND2X2 AND2X2_2198 ( .A(AES_CORE_DATAPATH__abc_16259_n6917), .B(AES_CORE_DATAPATH__abc_16259_n6918), .Y(AES_CORE_DATAPATH__abc_16259_n6919) );
  AND2X2 AND2X2_2199 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf6), .B(AES_CORE_DATAPATH__abc_16259_n6919), .Y(AES_CORE_DATAPATH__abc_16259_n6920) );
  AND2X2 AND2X2_22 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n96_1), .B(AES_CORE_CONTROL_UNIT__abc_15841_n98), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n99_1) );
  AND2X2 AND2X2_220 ( .A(AES_CORE_DATAPATH__abc_16259_n2683_1), .B(AES_CORE_DATAPATH__abc_16259_n2685_1), .Y(AES_CORE_DATAPATH__abc_16259_n2686) );
  AND2X2 AND2X2_2200 ( .A(AES_CORE_DATAPATH__abc_16259_n6921), .B(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6922) );
  AND2X2 AND2X2_2201 ( .A(AES_CORE_DATAPATH__abc_16259_n3540), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n6925) );
  AND2X2 AND2X2_2202 ( .A(AES_CORE_DATAPATH__abc_16259_n6925), .B(AES_CORE_DATAPATH__abc_16259_n6924), .Y(AES_CORE_DATAPATH__abc_16259_n6926) );
  AND2X2 AND2X2_2203 ( .A(AES_CORE_DATAPATH__abc_16259_n6928), .B(AES_CORE_DATAPATH__abc_16259_n6059_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6929) );
  AND2X2 AND2X2_2204 ( .A(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n6930), .Y(AES_CORE_DATAPATH__abc_16259_n6931) );
  AND2X2 AND2X2_2205 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf6), .B(AES_CORE_DATAPATH_bkp_0__17_), .Y(AES_CORE_DATAPATH__abc_16259_n6933) );
  AND2X2 AND2X2_2206 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf5), .B(AES_CORE_DATAPATH_bkp_1__17_), .Y(AES_CORE_DATAPATH__abc_16259_n6934) );
  AND2X2 AND2X2_2207 ( .A(AES_CORE_DATAPATH__abc_16259_n6937), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n6938) );
  AND2X2 AND2X2_2208 ( .A(AES_CORE_DATAPATH__abc_16259_n6936), .B(AES_CORE_DATAPATH__abc_16259_n6938), .Y(AES_CORE_DATAPATH__abc_16259_n6939) );
  AND2X2 AND2X2_2209 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf5), .B(AES_CORE_DATAPATH_bkp_3__17_), .Y(AES_CORE_DATAPATH__abc_16259_n6940) );
  AND2X2 AND2X2_221 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf0), .B(AES_CORE_DATAPATH_iv_3__22_), .Y(AES_CORE_DATAPATH__abc_16259_n2687_1) );
  AND2X2 AND2X2_2210 ( .A(AES_CORE_DATAPATH__abc_16259_n6943), .B(AES_CORE_DATAPATH__abc_16259_n6942), .Y(AES_CORE_DATAPATH__abc_16259_n6944) );
  AND2X2 AND2X2_2211 ( .A(AES_CORE_DATAPATH__abc_16259_n6946), .B(AES_CORE_DATAPATH__abc_16259_n6947), .Y(AES_CORE_DATAPATH__abc_16259_n6948) );
  AND2X2 AND2X2_2212 ( .A(AES_CORE_DATAPATH__abc_16259_n6945), .B(AES_CORE_DATAPATH__abc_16259_n6950), .Y(AES_CORE_DATAPATH__abc_16259_n6951) );
  AND2X2 AND2X2_2213 ( .A(AES_CORE_DATAPATH__abc_16259_n6951), .B(AES_CORE_CONTROL_UNIT_last_round_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6952) );
  AND2X2 AND2X2_2214 ( .A(AES_CORE_DATAPATH__abc_16259_n6953), .B(AES_CORE_DATAPATH__abc_16259_n6057_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6954) );
  AND2X2 AND2X2_2215 ( .A(AES_CORE_DATAPATH__abc_16259_n6951), .B(AES_CORE_DATAPATH__abc_16259_n6097_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6957) );
  AND2X2 AND2X2_2216 ( .A(AES_CORE_DATAPATH__abc_16259_n6095_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n6930), .Y(AES_CORE_DATAPATH__abc_16259_n6958) );
  AND2X2 AND2X2_2217 ( .A(AES_CORE_DATAPATH__abc_16259_n6960), .B(AES_CORE_DATAPATH__abc_16259_n6961), .Y(AES_CORE_DATAPATH__abc_16259_n6962) );
  AND2X2 AND2X2_2218 ( .A(AES_CORE_DATAPATH__abc_16259_n6962), .B(AES_CORE_DATAPATH__abc_16259_n6956), .Y(AES_CORE_DATAPATH__abc_16259_n6963) );
  AND2X2 AND2X2_2219 ( .A(AES_CORE_DATAPATH__abc_16259_n6964), .B(AES_CORE_DATAPATH__abc_16259_n6965), .Y(AES_CORE_DATAPATH__abc_16259_n6966) );
  AND2X2 AND2X2_222 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf0), .B(AES_CORE_DATAPATH_iv_0__23_), .Y(AES_CORE_DATAPATH__abc_16259_n2689_1) );
  AND2X2 AND2X2_2220 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf7), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_81_), .Y(AES_CORE_DATAPATH__abc_16259_n6969) );
  AND2X2 AND2X2_2221 ( .A(AES_CORE_DATAPATH__abc_16259_n6968), .B(AES_CORE_DATAPATH__abc_16259_n6970), .Y(AES_CORE_DATAPATH__abc_16259_n6971) );
  AND2X2 AND2X2_2222 ( .A(AES_CORE_DATAPATH__abc_16259_n6966), .B(AES_CORE_DATAPATH__abc_16259_n6972), .Y(AES_CORE_DATAPATH__abc_16259_n6973) );
  AND2X2 AND2X2_2223 ( .A(AES_CORE_DATAPATH__abc_16259_n6973), .B(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n6974) );
  AND2X2 AND2X2_2224 ( .A(AES_CORE_DATAPATH__abc_16259_n6975), .B(AES_CORE_DATAPATH__abc_16259_n6976), .Y(AES_CORE_DATAPATH__0col_0__31_0__17_) );
  AND2X2 AND2X2_2225 ( .A(AES_CORE_DATAPATH__abc_16259_n6044_bF_buf1), .B(AES_CORE_DATAPATH_col_0__18_), .Y(AES_CORE_DATAPATH__abc_16259_n6978) );
  AND2X2 AND2X2_2226 ( .A(AES_CORE_DATAPATH__abc_16259_n3589_1), .B(AES_CORE_DATAPATH__abc_16259_n6059_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6979) );
  AND2X2 AND2X2_2227 ( .A(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf6), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_18_), .Y(AES_CORE_DATAPATH__abc_16259_n6980) );
  AND2X2 AND2X2_2228 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf5), .B(AES_CORE_DATAPATH_bkp_0__18_), .Y(AES_CORE_DATAPATH__abc_16259_n6982) );
  AND2X2 AND2X2_2229 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf4), .B(AES_CORE_DATAPATH_bkp_1__18_), .Y(AES_CORE_DATAPATH__abc_16259_n6983) );
  AND2X2 AND2X2_223 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf7), .B(AES_CORE_DATAPATH_iv_1__23_), .Y(AES_CORE_DATAPATH__abc_16259_n2690) );
  AND2X2 AND2X2_2230 ( .A(AES_CORE_DATAPATH__abc_16259_n6986), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n6987) );
  AND2X2 AND2X2_2231 ( .A(AES_CORE_DATAPATH__abc_16259_n6985), .B(AES_CORE_DATAPATH__abc_16259_n6987), .Y(AES_CORE_DATAPATH__abc_16259_n6988) );
  AND2X2 AND2X2_2232 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf4), .B(AES_CORE_DATAPATH_bkp_3__18_), .Y(AES_CORE_DATAPATH__abc_16259_n6989) );
  AND2X2 AND2X2_2233 ( .A(AES_CORE_DATAPATH__abc_16259_n6991), .B(AES_CORE_DATAPATH__abc_16259_n6992), .Y(AES_CORE_DATAPATH__abc_16259_n6993) );
  AND2X2 AND2X2_2234 ( .A(AES_CORE_DATAPATH__abc_16259_n3580), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6996) );
  AND2X2 AND2X2_2235 ( .A(AES_CORE_DATAPATH__abc_16259_n6996), .B(AES_CORE_DATAPATH__abc_16259_n6995), .Y(AES_CORE_DATAPATH__abc_16259_n6997) );
  AND2X2 AND2X2_2236 ( .A(AES_CORE_DATAPATH__abc_16259_n7000), .B(AES_CORE_DATAPATH__abc_16259_n7001), .Y(AES_CORE_DATAPATH__abc_16259_n7002) );
  AND2X2 AND2X2_2237 ( .A(AES_CORE_DATAPATH__abc_16259_n6994), .B(AES_CORE_DATAPATH__abc_16259_n7004), .Y(AES_CORE_DATAPATH__abc_16259_n7005) );
  AND2X2 AND2X2_2238 ( .A(AES_CORE_DATAPATH__abc_16259_n7007), .B(AES_CORE_DATAPATH__abc_16259_n6092_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n7008) );
  AND2X2 AND2X2_2239 ( .A(AES_CORE_DATAPATH__abc_16259_n7006), .B(AES_CORE_DATAPATH__abc_16259_n7008), .Y(AES_CORE_DATAPATH__abc_16259_n7009) );
  AND2X2 AND2X2_224 ( .A(AES_CORE_DATAPATH__abc_16259_n2693_1), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n2694) );
  AND2X2 AND2X2_2240 ( .A(AES_CORE_DATAPATH__abc_16259_n7011), .B(AES_CORE_CONTROL_UNIT_mode_cbc_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7012) );
  AND2X2 AND2X2_2241 ( .A(AES_CORE_DATAPATH__abc_16259_n7010), .B(AES_CORE_DATAPATH__abc_16259_n7012), .Y(AES_CORE_DATAPATH__abc_16259_n7013) );
  AND2X2 AND2X2_2242 ( .A(AES_CORE_DATAPATH__abc_16259_n6101_bF_buf0), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_18_), .Y(AES_CORE_DATAPATH__abc_16259_n7014) );
  AND2X2 AND2X2_2243 ( .A(AES_CORE_DATAPATH__abc_16259_n7016), .B(AES_CORE_DATAPATH__abc_16259_n6056_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n7017) );
  AND2X2 AND2X2_2244 ( .A(AES_CORE_DATAPATH__abc_16259_n3589_1), .B(AES_CORE_DATAPATH__abc_16259_n6053_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n7018) );
  AND2X2 AND2X2_2245 ( .A(AES_CORE_DATAPATH__abc_16259_n7020), .B(AES_CORE_DATAPATH__abc_16259_n7021), .Y(AES_CORE_DATAPATH__abc_16259_n7022) );
  AND2X2 AND2X2_2246 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf5), .B(AES_CORE_DATAPATH__abc_16259_n7022), .Y(AES_CORE_DATAPATH__abc_16259_n7023) );
  AND2X2 AND2X2_2247 ( .A(AES_CORE_DATAPATH__abc_16259_n7024), .B(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7025) );
  AND2X2 AND2X2_2248 ( .A(AES_CORE_DATAPATH__abc_16259_n6044_bF_buf0), .B(AES_CORE_DATAPATH_col_0__19_), .Y(AES_CORE_DATAPATH__abc_16259_n7027) );
  AND2X2 AND2X2_2249 ( .A(AES_CORE_DATAPATH__abc_16259_n3629), .B(AES_CORE_DATAPATH__abc_16259_n6059_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n7028) );
  AND2X2 AND2X2_225 ( .A(AES_CORE_DATAPATH__abc_16259_n2692), .B(AES_CORE_DATAPATH__abc_16259_n2694), .Y(AES_CORE_DATAPATH__abc_16259_n2695_1) );
  AND2X2 AND2X2_2250 ( .A(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf4), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_19_), .Y(AES_CORE_DATAPATH__abc_16259_n7029) );
  AND2X2 AND2X2_2251 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf4), .B(AES_CORE_DATAPATH_bkp_0__19_), .Y(AES_CORE_DATAPATH__abc_16259_n7031) );
  AND2X2 AND2X2_2252 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1__19_), .Y(AES_CORE_DATAPATH__abc_16259_n7032) );
  AND2X2 AND2X2_2253 ( .A(AES_CORE_DATAPATH__abc_16259_n7035), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7036) );
  AND2X2 AND2X2_2254 ( .A(AES_CORE_DATAPATH__abc_16259_n7034), .B(AES_CORE_DATAPATH__abc_16259_n7036), .Y(AES_CORE_DATAPATH__abc_16259_n7037) );
  AND2X2 AND2X2_2255 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf3), .B(AES_CORE_DATAPATH_bkp_3__19_), .Y(AES_CORE_DATAPATH__abc_16259_n7038) );
  AND2X2 AND2X2_2256 ( .A(AES_CORE_DATAPATH__abc_16259_n7040), .B(AES_CORE_DATAPATH__abc_16259_n7041), .Y(AES_CORE_DATAPATH__abc_16259_n7042) );
  AND2X2 AND2X2_2257 ( .A(AES_CORE_DATAPATH__abc_16259_n3620_1), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7045) );
  AND2X2 AND2X2_2258 ( .A(AES_CORE_DATAPATH__abc_16259_n7045), .B(AES_CORE_DATAPATH__abc_16259_n7044), .Y(AES_CORE_DATAPATH__abc_16259_n7046) );
  AND2X2 AND2X2_2259 ( .A(AES_CORE_DATAPATH__abc_16259_n7049), .B(AES_CORE_DATAPATH__abc_16259_n7050), .Y(AES_CORE_DATAPATH__abc_16259_n7051) );
  AND2X2 AND2X2_226 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf7), .B(AES_CORE_DATAPATH_iv_3__23_), .Y(AES_CORE_DATAPATH__abc_16259_n2696) );
  AND2X2 AND2X2_2260 ( .A(AES_CORE_DATAPATH__abc_16259_n7043), .B(AES_CORE_DATAPATH__abc_16259_n7053), .Y(AES_CORE_DATAPATH__abc_16259_n7054) );
  AND2X2 AND2X2_2261 ( .A(AES_CORE_DATAPATH__abc_16259_n7056), .B(AES_CORE_DATAPATH__abc_16259_n6092_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7057) );
  AND2X2 AND2X2_2262 ( .A(AES_CORE_DATAPATH__abc_16259_n7055), .B(AES_CORE_DATAPATH__abc_16259_n7057), .Y(AES_CORE_DATAPATH__abc_16259_n7058) );
  AND2X2 AND2X2_2263 ( .A(AES_CORE_DATAPATH__abc_16259_n7060), .B(AES_CORE_CONTROL_UNIT_mode_cbc_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7061) );
  AND2X2 AND2X2_2264 ( .A(AES_CORE_DATAPATH__abc_16259_n7059), .B(AES_CORE_DATAPATH__abc_16259_n7061), .Y(AES_CORE_DATAPATH__abc_16259_n7062) );
  AND2X2 AND2X2_2265 ( .A(AES_CORE_DATAPATH__abc_16259_n6101_bF_buf4), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_19_), .Y(AES_CORE_DATAPATH__abc_16259_n7063) );
  AND2X2 AND2X2_2266 ( .A(AES_CORE_DATAPATH__abc_16259_n7065), .B(AES_CORE_DATAPATH__abc_16259_n6056_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7066) );
  AND2X2 AND2X2_2267 ( .A(AES_CORE_DATAPATH__abc_16259_n3629), .B(AES_CORE_DATAPATH__abc_16259_n6053_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7067) );
  AND2X2 AND2X2_2268 ( .A(AES_CORE_DATAPATH__abc_16259_n7069), .B(AES_CORE_DATAPATH__abc_16259_n7070), .Y(AES_CORE_DATAPATH__abc_16259_n7071) );
  AND2X2 AND2X2_2269 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n7071), .Y(AES_CORE_DATAPATH__abc_16259_n7072) );
  AND2X2 AND2X2_227 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf7), .B(AES_CORE_DATAPATH_iv_0__24_), .Y(AES_CORE_DATAPATH__abc_16259_n2698) );
  AND2X2 AND2X2_2270 ( .A(AES_CORE_DATAPATH__abc_16259_n7073), .B(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7074) );
  AND2X2 AND2X2_2271 ( .A(AES_CORE_DATAPATH__abc_16259_n6044_bF_buf4), .B(AES_CORE_DATAPATH_col_0__20_), .Y(AES_CORE_DATAPATH__abc_16259_n7076) );
  AND2X2 AND2X2_2272 ( .A(AES_CORE_DATAPATH__abc_16259_n7077), .B(AES_CORE_DATAPATH__abc_16259_n7078), .Y(AES_CORE_DATAPATH__abc_16259_n7079) );
  AND2X2 AND2X2_2273 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf3), .B(AES_CORE_DATAPATH_bkp_0__20_), .Y(AES_CORE_DATAPATH__abc_16259_n7080) );
  AND2X2 AND2X2_2274 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf2), .B(AES_CORE_DATAPATH_bkp_1__20_), .Y(AES_CORE_DATAPATH__abc_16259_n7081) );
  AND2X2 AND2X2_2275 ( .A(AES_CORE_DATAPATH__abc_16259_n7084), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7085) );
  AND2X2 AND2X2_2276 ( .A(AES_CORE_DATAPATH__abc_16259_n7083), .B(AES_CORE_DATAPATH__abc_16259_n7085), .Y(AES_CORE_DATAPATH__abc_16259_n7086) );
  AND2X2 AND2X2_2277 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf2), .B(AES_CORE_DATAPATH_bkp_3__20_), .Y(AES_CORE_DATAPATH__abc_16259_n7087) );
  AND2X2 AND2X2_2278 ( .A(AES_CORE_DATAPATH__abc_16259_n7089), .B(AES_CORE_DATAPATH__abc_16259_n7090), .Y(AES_CORE_DATAPATH__abc_16259_n7091) );
  AND2X2 AND2X2_2279 ( .A(AES_CORE_DATAPATH__abc_16259_n3660), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n7094) );
  AND2X2 AND2X2_228 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf6), .B(AES_CORE_DATAPATH_iv_1__24_), .Y(AES_CORE_DATAPATH__abc_16259_n2699_1) );
  AND2X2 AND2X2_2280 ( .A(AES_CORE_DATAPATH__abc_16259_n7094), .B(AES_CORE_DATAPATH__abc_16259_n7093), .Y(AES_CORE_DATAPATH__abc_16259_n7095) );
  AND2X2 AND2X2_2281 ( .A(AES_CORE_DATAPATH__abc_16259_n7097), .B(AES_CORE_DATAPATH__abc_16259_n6059_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n7098) );
  AND2X2 AND2X2_2282 ( .A(AES_CORE_DATAPATH__abc_16259_n7092), .B(AES_CORE_DATAPATH__abc_16259_n7102), .Y(AES_CORE_DATAPATH__abc_16259_n7103) );
  AND2X2 AND2X2_2283 ( .A(AES_CORE_DATAPATH__abc_16259_n7105), .B(AES_CORE_DATAPATH__abc_16259_n6092_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7106) );
  AND2X2 AND2X2_2284 ( .A(AES_CORE_DATAPATH__abc_16259_n7104), .B(AES_CORE_DATAPATH__abc_16259_n7106), .Y(AES_CORE_DATAPATH__abc_16259_n7107) );
  AND2X2 AND2X2_2285 ( .A(AES_CORE_DATAPATH__abc_16259_n7109), .B(AES_CORE_CONTROL_UNIT_mode_cbc_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n7110) );
  AND2X2 AND2X2_2286 ( .A(AES_CORE_DATAPATH__abc_16259_n7108), .B(AES_CORE_DATAPATH__abc_16259_n7110), .Y(AES_CORE_DATAPATH__abc_16259_n7111) );
  AND2X2 AND2X2_2287 ( .A(AES_CORE_DATAPATH__abc_16259_n6101_bF_buf3), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_20_), .Y(AES_CORE_DATAPATH__abc_16259_n7112) );
  AND2X2 AND2X2_2288 ( .A(AES_CORE_DATAPATH__abc_16259_n7114), .B(AES_CORE_DATAPATH__abc_16259_n6056_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7115) );
  AND2X2 AND2X2_2289 ( .A(AES_CORE_DATAPATH__abc_16259_n3669), .B(AES_CORE_DATAPATH__abc_16259_n6053_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7116) );
  AND2X2 AND2X2_229 ( .A(AES_CORE_DATAPATH__abc_16259_n2702), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n2703_1) );
  AND2X2 AND2X2_2290 ( .A(AES_CORE_DATAPATH__abc_16259_n7118), .B(AES_CORE_DATAPATH__abc_16259_n7119), .Y(AES_CORE_DATAPATH__abc_16259_n7120) );
  AND2X2 AND2X2_2291 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n7120), .Y(AES_CORE_DATAPATH__abc_16259_n7121) );
  AND2X2 AND2X2_2292 ( .A(AES_CORE_DATAPATH__abc_16259_n7122), .B(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n7123) );
  AND2X2 AND2X2_2293 ( .A(AES_CORE_DATAPATH__abc_16259_n3700), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n7126) );
  AND2X2 AND2X2_2294 ( .A(AES_CORE_DATAPATH__abc_16259_n7126), .B(AES_CORE_DATAPATH__abc_16259_n7125), .Y(AES_CORE_DATAPATH__abc_16259_n7127) );
  AND2X2 AND2X2_2295 ( .A(AES_CORE_DATAPATH__abc_16259_n7129), .B(AES_CORE_DATAPATH__abc_16259_n6059_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n7130) );
  AND2X2 AND2X2_2296 ( .A(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n7131), .Y(AES_CORE_DATAPATH__abc_16259_n7132) );
  AND2X2 AND2X2_2297 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf2), .B(AES_CORE_DATAPATH_bkp_0__21_), .Y(AES_CORE_DATAPATH__abc_16259_n7134) );
  AND2X2 AND2X2_2298 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf1), .B(AES_CORE_DATAPATH_bkp_1__21_), .Y(AES_CORE_DATAPATH__abc_16259_n7135) );
  AND2X2 AND2X2_2299 ( .A(AES_CORE_DATAPATH__abc_16259_n7138), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n7139) );
  AND2X2 AND2X2_23 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n99_1), .B(AES_CORE_CONTROL_UNIT__abc_15841_n95), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n100) );
  AND2X2 AND2X2_230 ( .A(AES_CORE_DATAPATH__abc_16259_n2701_1), .B(AES_CORE_DATAPATH__abc_16259_n2703_1), .Y(AES_CORE_DATAPATH__abc_16259_n2704) );
  AND2X2 AND2X2_2300 ( .A(AES_CORE_DATAPATH__abc_16259_n7137), .B(AES_CORE_DATAPATH__abc_16259_n7139), .Y(AES_CORE_DATAPATH__abc_16259_n7140) );
  AND2X2 AND2X2_2301 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf1), .B(AES_CORE_DATAPATH_bkp_3__21_), .Y(AES_CORE_DATAPATH__abc_16259_n7141) );
  AND2X2 AND2X2_2302 ( .A(AES_CORE_DATAPATH__abc_16259_n7144), .B(AES_CORE_DATAPATH__abc_16259_n7143), .Y(AES_CORE_DATAPATH__abc_16259_n7145) );
  AND2X2 AND2X2_2303 ( .A(AES_CORE_DATAPATH__abc_16259_n7147), .B(AES_CORE_DATAPATH__abc_16259_n7148), .Y(AES_CORE_DATAPATH__abc_16259_n7149) );
  AND2X2 AND2X2_2304 ( .A(AES_CORE_DATAPATH__abc_16259_n7146), .B(AES_CORE_DATAPATH__abc_16259_n7151), .Y(AES_CORE_DATAPATH__abc_16259_n7152) );
  AND2X2 AND2X2_2305 ( .A(AES_CORE_DATAPATH__abc_16259_n7152), .B(AES_CORE_CONTROL_UNIT_last_round_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n7153) );
  AND2X2 AND2X2_2306 ( .A(AES_CORE_DATAPATH__abc_16259_n7154), .B(AES_CORE_DATAPATH__abc_16259_n6057_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n7155) );
  AND2X2 AND2X2_2307 ( .A(AES_CORE_DATAPATH__abc_16259_n7152), .B(AES_CORE_DATAPATH__abc_16259_n6097_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7158) );
  AND2X2 AND2X2_2308 ( .A(AES_CORE_DATAPATH__abc_16259_n6095_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n7131), .Y(AES_CORE_DATAPATH__abc_16259_n7159) );
  AND2X2 AND2X2_2309 ( .A(AES_CORE_DATAPATH__abc_16259_n7161), .B(AES_CORE_DATAPATH__abc_16259_n7162), .Y(AES_CORE_DATAPATH__abc_16259_n7163) );
  AND2X2 AND2X2_231 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf6), .B(AES_CORE_DATAPATH_iv_3__24_), .Y(AES_CORE_DATAPATH__abc_16259_n2705_1) );
  AND2X2 AND2X2_2310 ( .A(AES_CORE_DATAPATH__abc_16259_n7163), .B(AES_CORE_DATAPATH__abc_16259_n7157), .Y(AES_CORE_DATAPATH__abc_16259_n7164) );
  AND2X2 AND2X2_2311 ( .A(AES_CORE_DATAPATH__abc_16259_n7165), .B(AES_CORE_DATAPATH__abc_16259_n7166), .Y(AES_CORE_DATAPATH__abc_16259_n7167) );
  AND2X2 AND2X2_2312 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf2), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_85_), .Y(AES_CORE_DATAPATH__abc_16259_n7170) );
  AND2X2 AND2X2_2313 ( .A(AES_CORE_DATAPATH__abc_16259_n7169), .B(AES_CORE_DATAPATH__abc_16259_n7171), .Y(AES_CORE_DATAPATH__abc_16259_n7172) );
  AND2X2 AND2X2_2314 ( .A(AES_CORE_DATAPATH__abc_16259_n7167), .B(AES_CORE_DATAPATH__abc_16259_n7173), .Y(AES_CORE_DATAPATH__abc_16259_n7174) );
  AND2X2 AND2X2_2315 ( .A(AES_CORE_DATAPATH__abc_16259_n7174), .B(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n7175) );
  AND2X2 AND2X2_2316 ( .A(AES_CORE_DATAPATH__abc_16259_n7176), .B(AES_CORE_DATAPATH__abc_16259_n7177), .Y(AES_CORE_DATAPATH__0col_0__31_0__21_) );
  AND2X2 AND2X2_2317 ( .A(AES_CORE_DATAPATH__abc_16259_n6044_bF_buf3), .B(AES_CORE_DATAPATH_col_0__22_), .Y(AES_CORE_DATAPATH__abc_16259_n7179) );
  AND2X2 AND2X2_2318 ( .A(AES_CORE_DATAPATH__abc_16259_n3749), .B(AES_CORE_DATAPATH__abc_16259_n6059_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7180) );
  AND2X2 AND2X2_2319 ( .A(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf6), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_22_), .Y(AES_CORE_DATAPATH__abc_16259_n7181) );
  AND2X2 AND2X2_232 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf6), .B(AES_CORE_DATAPATH_iv_0__25_), .Y(AES_CORE_DATAPATH__abc_16259_n2707_1) );
  AND2X2 AND2X2_2320 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf1), .B(AES_CORE_DATAPATH_bkp_0__22_), .Y(AES_CORE_DATAPATH__abc_16259_n7183) );
  AND2X2 AND2X2_2321 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf0), .B(AES_CORE_DATAPATH_bkp_1__22_), .Y(AES_CORE_DATAPATH__abc_16259_n7184) );
  AND2X2 AND2X2_2322 ( .A(AES_CORE_DATAPATH__abc_16259_n7187), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n7188) );
  AND2X2 AND2X2_2323 ( .A(AES_CORE_DATAPATH__abc_16259_n7186), .B(AES_CORE_DATAPATH__abc_16259_n7188), .Y(AES_CORE_DATAPATH__abc_16259_n7189) );
  AND2X2 AND2X2_2324 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf0), .B(AES_CORE_DATAPATH_bkp_3__22_), .Y(AES_CORE_DATAPATH__abc_16259_n7190) );
  AND2X2 AND2X2_2325 ( .A(AES_CORE_DATAPATH__abc_16259_n7192), .B(AES_CORE_DATAPATH__abc_16259_n7193), .Y(AES_CORE_DATAPATH__abc_16259_n7194) );
  AND2X2 AND2X2_2326 ( .A(AES_CORE_DATAPATH__abc_16259_n3740), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n7197) );
  AND2X2 AND2X2_2327 ( .A(AES_CORE_DATAPATH__abc_16259_n7197), .B(AES_CORE_DATAPATH__abc_16259_n7196), .Y(AES_CORE_DATAPATH__abc_16259_n7198) );
  AND2X2 AND2X2_2328 ( .A(AES_CORE_DATAPATH__abc_16259_n7201), .B(AES_CORE_DATAPATH__abc_16259_n7202), .Y(AES_CORE_DATAPATH__abc_16259_n7203) );
  AND2X2 AND2X2_2329 ( .A(AES_CORE_DATAPATH__abc_16259_n7195), .B(AES_CORE_DATAPATH__abc_16259_n7205), .Y(AES_CORE_DATAPATH__abc_16259_n7206) );
  AND2X2 AND2X2_233 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf5), .B(AES_CORE_DATAPATH_iv_1__25_), .Y(AES_CORE_DATAPATH__abc_16259_n2708) );
  AND2X2 AND2X2_2330 ( .A(AES_CORE_DATAPATH__abc_16259_n7208), .B(AES_CORE_DATAPATH__abc_16259_n6092_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n7209) );
  AND2X2 AND2X2_2331 ( .A(AES_CORE_DATAPATH__abc_16259_n7207), .B(AES_CORE_DATAPATH__abc_16259_n7209), .Y(AES_CORE_DATAPATH__abc_16259_n7210) );
  AND2X2 AND2X2_2332 ( .A(AES_CORE_DATAPATH__abc_16259_n7212), .B(AES_CORE_CONTROL_UNIT_mode_cbc_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n7213) );
  AND2X2 AND2X2_2333 ( .A(AES_CORE_DATAPATH__abc_16259_n7211), .B(AES_CORE_DATAPATH__abc_16259_n7213), .Y(AES_CORE_DATAPATH__abc_16259_n7214) );
  AND2X2 AND2X2_2334 ( .A(AES_CORE_DATAPATH__abc_16259_n6101_bF_buf2), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_22_), .Y(AES_CORE_DATAPATH__abc_16259_n7215) );
  AND2X2 AND2X2_2335 ( .A(AES_CORE_DATAPATH__abc_16259_n7217), .B(AES_CORE_DATAPATH__abc_16259_n6056_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n7218) );
  AND2X2 AND2X2_2336 ( .A(AES_CORE_DATAPATH__abc_16259_n3749), .B(AES_CORE_DATAPATH__abc_16259_n6053_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n7219) );
  AND2X2 AND2X2_2337 ( .A(AES_CORE_DATAPATH__abc_16259_n7221), .B(AES_CORE_DATAPATH__abc_16259_n7222), .Y(AES_CORE_DATAPATH__abc_16259_n7223) );
  AND2X2 AND2X2_2338 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n7223), .Y(AES_CORE_DATAPATH__abc_16259_n7224) );
  AND2X2 AND2X2_2339 ( .A(AES_CORE_DATAPATH__abc_16259_n7225), .B(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n7226) );
  AND2X2 AND2X2_234 ( .A(AES_CORE_DATAPATH__abc_16259_n2711_1), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n2712) );
  AND2X2 AND2X2_2340 ( .A(AES_CORE_DATAPATH__abc_16259_n6044_bF_buf2), .B(AES_CORE_DATAPATH_col_0__23_), .Y(AES_CORE_DATAPATH__abc_16259_n7228) );
  AND2X2 AND2X2_2341 ( .A(AES_CORE_DATAPATH__abc_16259_n3780), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n7230) );
  AND2X2 AND2X2_2342 ( .A(AES_CORE_DATAPATH__abc_16259_n7230), .B(AES_CORE_DATAPATH__abc_16259_n7229), .Y(AES_CORE_DATAPATH__abc_16259_n7231) );
  AND2X2 AND2X2_2343 ( .A(AES_CORE_DATAPATH__abc_16259_n7233), .B(AES_CORE_DATAPATH__abc_16259_n6059_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7234) );
  AND2X2 AND2X2_2344 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf0), .B(AES_CORE_DATAPATH_bkp_0__23_), .Y(AES_CORE_DATAPATH__abc_16259_n7238) );
  AND2X2 AND2X2_2345 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf7), .B(AES_CORE_DATAPATH_bkp_1__23_), .Y(AES_CORE_DATAPATH__abc_16259_n7239) );
  AND2X2 AND2X2_2346 ( .A(AES_CORE_DATAPATH__abc_16259_n7242), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n7243) );
  AND2X2 AND2X2_2347 ( .A(AES_CORE_DATAPATH__abc_16259_n7241), .B(AES_CORE_DATAPATH__abc_16259_n7243), .Y(AES_CORE_DATAPATH__abc_16259_n7244) );
  AND2X2 AND2X2_2348 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf7), .B(AES_CORE_DATAPATH_bkp_3__23_), .Y(AES_CORE_DATAPATH__abc_16259_n7245) );
  AND2X2 AND2X2_2349 ( .A(AES_CORE_DATAPATH__abc_16259_n7247), .B(AES_CORE_DATAPATH__abc_16259_n7248), .Y(AES_CORE_DATAPATH__abc_16259_n7249) );
  AND2X2 AND2X2_235 ( .A(AES_CORE_DATAPATH__abc_16259_n2710), .B(AES_CORE_DATAPATH__abc_16259_n2712), .Y(AES_CORE_DATAPATH__abc_16259_n2713_1) );
  AND2X2 AND2X2_2350 ( .A(AES_CORE_DATAPATH__abc_16259_n7252), .B(AES_CORE_DATAPATH__abc_16259_n7235), .Y(AES_CORE_DATAPATH__abc_16259_n7253) );
  AND2X2 AND2X2_2351 ( .A(AES_CORE_DATAPATH__abc_16259_n7251), .B(AES_CORE_DATAPATH__abc_16259_n7254), .Y(AES_CORE_DATAPATH__abc_16259_n7255) );
  AND2X2 AND2X2_2352 ( .A(AES_CORE_DATAPATH__abc_16259_n7257), .B(AES_CORE_DATAPATH__abc_16259_n6092_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n7258) );
  AND2X2 AND2X2_2353 ( .A(AES_CORE_DATAPATH__abc_16259_n7256), .B(AES_CORE_DATAPATH__abc_16259_n7258), .Y(AES_CORE_DATAPATH__abc_16259_n7259) );
  AND2X2 AND2X2_2354 ( .A(AES_CORE_DATAPATH__abc_16259_n7261), .B(AES_CORE_CONTROL_UNIT_mode_cbc_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n7262) );
  AND2X2 AND2X2_2355 ( .A(AES_CORE_DATAPATH__abc_16259_n7260), .B(AES_CORE_DATAPATH__abc_16259_n7262), .Y(AES_CORE_DATAPATH__abc_16259_n7263) );
  AND2X2 AND2X2_2356 ( .A(AES_CORE_DATAPATH__abc_16259_n6101_bF_buf1), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_23_), .Y(AES_CORE_DATAPATH__abc_16259_n7264) );
  AND2X2 AND2X2_2357 ( .A(AES_CORE_DATAPATH__abc_16259_n7266), .B(AES_CORE_DATAPATH__abc_16259_n6056_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n7267) );
  AND2X2 AND2X2_2358 ( .A(AES_CORE_DATAPATH__abc_16259_n3789), .B(AES_CORE_DATAPATH__abc_16259_n6053_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n7268) );
  AND2X2 AND2X2_2359 ( .A(AES_CORE_DATAPATH__abc_16259_n7270), .B(AES_CORE_DATAPATH__abc_16259_n7271), .Y(AES_CORE_DATAPATH__abc_16259_n7272) );
  AND2X2 AND2X2_236 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf5), .B(AES_CORE_DATAPATH_iv_3__25_), .Y(AES_CORE_DATAPATH__abc_16259_n2714) );
  AND2X2 AND2X2_2360 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n7272), .Y(AES_CORE_DATAPATH__abc_16259_n7273) );
  AND2X2 AND2X2_2361 ( .A(AES_CORE_DATAPATH__abc_16259_n7274), .B(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7275) );
  AND2X2 AND2X2_2362 ( .A(AES_CORE_DATAPATH__abc_16259_n6044_bF_buf1), .B(AES_CORE_DATAPATH_col_0__24_), .Y(AES_CORE_DATAPATH__abc_16259_n7277) );
  AND2X2 AND2X2_2363 ( .A(AES_CORE_DATAPATH__abc_16259_n3829), .B(AES_CORE_DATAPATH__abc_16259_n6059_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n7278) );
  AND2X2 AND2X2_2364 ( .A(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf3), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_24_), .Y(AES_CORE_DATAPATH__abc_16259_n7279) );
  AND2X2 AND2X2_2365 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf7), .B(AES_CORE_DATAPATH_bkp_0__24_), .Y(AES_CORE_DATAPATH__abc_16259_n7281) );
  AND2X2 AND2X2_2366 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf6), .B(AES_CORE_DATAPATH_bkp_1__24_), .Y(AES_CORE_DATAPATH__abc_16259_n7282) );
  AND2X2 AND2X2_2367 ( .A(AES_CORE_DATAPATH__abc_16259_n7285), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n7286) );
  AND2X2 AND2X2_2368 ( .A(AES_CORE_DATAPATH__abc_16259_n7284), .B(AES_CORE_DATAPATH__abc_16259_n7286), .Y(AES_CORE_DATAPATH__abc_16259_n7287) );
  AND2X2 AND2X2_2369 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf6), .B(AES_CORE_DATAPATH_bkp_3__24_), .Y(AES_CORE_DATAPATH__abc_16259_n7288) );
  AND2X2 AND2X2_237 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf5), .B(AES_CORE_DATAPATH_iv_0__26_), .Y(AES_CORE_DATAPATH__abc_16259_n2716) );
  AND2X2 AND2X2_2370 ( .A(AES_CORE_DATAPATH__abc_16259_n7290), .B(AES_CORE_DATAPATH__abc_16259_n7291), .Y(AES_CORE_DATAPATH__abc_16259_n7292) );
  AND2X2 AND2X2_2371 ( .A(AES_CORE_DATAPATH__abc_16259_n3820), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n7295) );
  AND2X2 AND2X2_2372 ( .A(AES_CORE_DATAPATH__abc_16259_n7295), .B(AES_CORE_DATAPATH__abc_16259_n7294), .Y(AES_CORE_DATAPATH__abc_16259_n7296) );
  AND2X2 AND2X2_2373 ( .A(AES_CORE_DATAPATH__abc_16259_n7299), .B(AES_CORE_DATAPATH__abc_16259_n7300), .Y(AES_CORE_DATAPATH__abc_16259_n7301) );
  AND2X2 AND2X2_2374 ( .A(AES_CORE_DATAPATH__abc_16259_n7293), .B(AES_CORE_DATAPATH__abc_16259_n7303), .Y(AES_CORE_DATAPATH__abc_16259_n7304) );
  AND2X2 AND2X2_2375 ( .A(AES_CORE_DATAPATH__abc_16259_n7306), .B(AES_CORE_DATAPATH__abc_16259_n6092_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n7307) );
  AND2X2 AND2X2_2376 ( .A(AES_CORE_DATAPATH__abc_16259_n7305), .B(AES_CORE_DATAPATH__abc_16259_n7307), .Y(AES_CORE_DATAPATH__abc_16259_n7308) );
  AND2X2 AND2X2_2377 ( .A(AES_CORE_DATAPATH__abc_16259_n7310), .B(AES_CORE_CONTROL_UNIT_mode_cbc_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7311) );
  AND2X2 AND2X2_2378 ( .A(AES_CORE_DATAPATH__abc_16259_n7309), .B(AES_CORE_DATAPATH__abc_16259_n7311), .Y(AES_CORE_DATAPATH__abc_16259_n7312) );
  AND2X2 AND2X2_2379 ( .A(AES_CORE_DATAPATH__abc_16259_n6101_bF_buf0), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_24_), .Y(AES_CORE_DATAPATH__abc_16259_n7313) );
  AND2X2 AND2X2_238 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf4), .B(AES_CORE_DATAPATH_iv_1__26_), .Y(AES_CORE_DATAPATH__abc_16259_n2717_1) );
  AND2X2 AND2X2_2380 ( .A(AES_CORE_DATAPATH__abc_16259_n7315), .B(AES_CORE_DATAPATH__abc_16259_n6056_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n7316) );
  AND2X2 AND2X2_2381 ( .A(AES_CORE_DATAPATH__abc_16259_n3829), .B(AES_CORE_DATAPATH__abc_16259_n6053_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n7317) );
  AND2X2 AND2X2_2382 ( .A(AES_CORE_DATAPATH__abc_16259_n7319), .B(AES_CORE_DATAPATH__abc_16259_n7320), .Y(AES_CORE_DATAPATH__abc_16259_n7321) );
  AND2X2 AND2X2_2383 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n7321), .Y(AES_CORE_DATAPATH__abc_16259_n7322) );
  AND2X2 AND2X2_2384 ( .A(AES_CORE_DATAPATH__abc_16259_n7323), .B(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7324) );
  AND2X2 AND2X2_2385 ( .A(AES_CORE_DATAPATH__abc_16259_n6044_bF_buf0), .B(AES_CORE_DATAPATH_col_0__25_), .Y(AES_CORE_DATAPATH__abc_16259_n7326) );
  AND2X2 AND2X2_2386 ( .A(AES_CORE_DATAPATH__abc_16259_n3869), .B(AES_CORE_DATAPATH__abc_16259_n6059_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n7327) );
  AND2X2 AND2X2_2387 ( .A(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf1), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_25_), .Y(AES_CORE_DATAPATH__abc_16259_n7328) );
  AND2X2 AND2X2_2388 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf6), .B(AES_CORE_DATAPATH_bkp_0__25_), .Y(AES_CORE_DATAPATH__abc_16259_n7330) );
  AND2X2 AND2X2_2389 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf5), .B(AES_CORE_DATAPATH_bkp_1__25_), .Y(AES_CORE_DATAPATH__abc_16259_n7331) );
  AND2X2 AND2X2_239 ( .A(AES_CORE_DATAPATH__abc_16259_n2720), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n2721_1) );
  AND2X2 AND2X2_2390 ( .A(AES_CORE_DATAPATH__abc_16259_n7334), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n7335) );
  AND2X2 AND2X2_2391 ( .A(AES_CORE_DATAPATH__abc_16259_n7333), .B(AES_CORE_DATAPATH__abc_16259_n7335), .Y(AES_CORE_DATAPATH__abc_16259_n7336) );
  AND2X2 AND2X2_2392 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf5), .B(AES_CORE_DATAPATH_bkp_3__25_), .Y(AES_CORE_DATAPATH__abc_16259_n7337) );
  AND2X2 AND2X2_2393 ( .A(AES_CORE_DATAPATH__abc_16259_n7339), .B(AES_CORE_DATAPATH__abc_16259_n7340), .Y(AES_CORE_DATAPATH__abc_16259_n7341) );
  AND2X2 AND2X2_2394 ( .A(AES_CORE_DATAPATH__abc_16259_n3860), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n7344) );
  AND2X2 AND2X2_2395 ( .A(AES_CORE_DATAPATH__abc_16259_n7344), .B(AES_CORE_DATAPATH__abc_16259_n7343), .Y(AES_CORE_DATAPATH__abc_16259_n7345) );
  AND2X2 AND2X2_2396 ( .A(AES_CORE_DATAPATH__abc_16259_n7348), .B(AES_CORE_DATAPATH__abc_16259_n7349), .Y(AES_CORE_DATAPATH__abc_16259_n7350) );
  AND2X2 AND2X2_2397 ( .A(AES_CORE_DATAPATH__abc_16259_n7342), .B(AES_CORE_DATAPATH__abc_16259_n7352), .Y(AES_CORE_DATAPATH__abc_16259_n7353) );
  AND2X2 AND2X2_2398 ( .A(AES_CORE_DATAPATH__abc_16259_n7355), .B(AES_CORE_DATAPATH__abc_16259_n6092_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7356) );
  AND2X2 AND2X2_2399 ( .A(AES_CORE_DATAPATH__abc_16259_n7354), .B(AES_CORE_DATAPATH__abc_16259_n7356), .Y(AES_CORE_DATAPATH__abc_16259_n7357) );
  AND2X2 AND2X2_24 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n95), .B(AES_CORE_CONTROL_UNIT__abc_15841_n104), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n105) );
  AND2X2 AND2X2_240 ( .A(AES_CORE_DATAPATH__abc_16259_n2719_1), .B(AES_CORE_DATAPATH__abc_16259_n2721_1), .Y(AES_CORE_DATAPATH__abc_16259_n2722) );
  AND2X2 AND2X2_2400 ( .A(AES_CORE_DATAPATH__abc_16259_n7359), .B(AES_CORE_CONTROL_UNIT_mode_cbc_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7360) );
  AND2X2 AND2X2_2401 ( .A(AES_CORE_DATAPATH__abc_16259_n7358), .B(AES_CORE_DATAPATH__abc_16259_n7360), .Y(AES_CORE_DATAPATH__abc_16259_n7361) );
  AND2X2 AND2X2_2402 ( .A(AES_CORE_DATAPATH__abc_16259_n6101_bF_buf4), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_25_), .Y(AES_CORE_DATAPATH__abc_16259_n7362) );
  AND2X2 AND2X2_2403 ( .A(AES_CORE_DATAPATH__abc_16259_n7364), .B(AES_CORE_DATAPATH__abc_16259_n6056_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7365) );
  AND2X2 AND2X2_2404 ( .A(AES_CORE_DATAPATH__abc_16259_n3869), .B(AES_CORE_DATAPATH__abc_16259_n6053_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7366) );
  AND2X2 AND2X2_2405 ( .A(AES_CORE_DATAPATH__abc_16259_n7368), .B(AES_CORE_DATAPATH__abc_16259_n7369), .Y(AES_CORE_DATAPATH__abc_16259_n7370) );
  AND2X2 AND2X2_2406 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf9), .B(AES_CORE_DATAPATH__abc_16259_n7370), .Y(AES_CORE_DATAPATH__abc_16259_n7371) );
  AND2X2 AND2X2_2407 ( .A(AES_CORE_DATAPATH__abc_16259_n7372), .B(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n7373) );
  AND2X2 AND2X2_2408 ( .A(AES_CORE_DATAPATH__abc_16259_n6044_bF_buf4), .B(AES_CORE_DATAPATH_col_0__26_), .Y(AES_CORE_DATAPATH__abc_16259_n7375) );
  AND2X2 AND2X2_2409 ( .A(AES_CORE_DATAPATH__abc_16259_n3900), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7377) );
  AND2X2 AND2X2_241 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf4), .B(AES_CORE_DATAPATH_iv_3__26_), .Y(AES_CORE_DATAPATH__abc_16259_n2723_1) );
  AND2X2 AND2X2_2410 ( .A(AES_CORE_DATAPATH__abc_16259_n7377), .B(AES_CORE_DATAPATH__abc_16259_n7376), .Y(AES_CORE_DATAPATH__abc_16259_n7378) );
  AND2X2 AND2X2_2411 ( .A(AES_CORE_DATAPATH__abc_16259_n7380), .B(AES_CORE_DATAPATH__abc_16259_n6059_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n7381) );
  AND2X2 AND2X2_2412 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf5), .B(AES_CORE_DATAPATH_bkp_0__26_), .Y(AES_CORE_DATAPATH__abc_16259_n7385) );
  AND2X2 AND2X2_2413 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf4), .B(AES_CORE_DATAPATH_bkp_1__26_), .Y(AES_CORE_DATAPATH__abc_16259_n7386) );
  AND2X2 AND2X2_2414 ( .A(AES_CORE_DATAPATH__abc_16259_n7389), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n7390) );
  AND2X2 AND2X2_2415 ( .A(AES_CORE_DATAPATH__abc_16259_n7388), .B(AES_CORE_DATAPATH__abc_16259_n7390), .Y(AES_CORE_DATAPATH__abc_16259_n7391) );
  AND2X2 AND2X2_2416 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf4), .B(AES_CORE_DATAPATH_bkp_3__26_), .Y(AES_CORE_DATAPATH__abc_16259_n7392) );
  AND2X2 AND2X2_2417 ( .A(AES_CORE_DATAPATH__abc_16259_n7394), .B(AES_CORE_DATAPATH__abc_16259_n7395), .Y(AES_CORE_DATAPATH__abc_16259_n7396) );
  AND2X2 AND2X2_2418 ( .A(AES_CORE_DATAPATH__abc_16259_n7399), .B(AES_CORE_DATAPATH__abc_16259_n7382), .Y(AES_CORE_DATAPATH__abc_16259_n7400) );
  AND2X2 AND2X2_2419 ( .A(AES_CORE_DATAPATH__abc_16259_n7398), .B(AES_CORE_DATAPATH__abc_16259_n7401), .Y(AES_CORE_DATAPATH__abc_16259_n7402) );
  AND2X2 AND2X2_242 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf4), .B(AES_CORE_DATAPATH_iv_0__27_), .Y(AES_CORE_DATAPATH__abc_16259_n2725) );
  AND2X2 AND2X2_2420 ( .A(AES_CORE_DATAPATH__abc_16259_n7404), .B(AES_CORE_DATAPATH__abc_16259_n6092_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7405) );
  AND2X2 AND2X2_2421 ( .A(AES_CORE_DATAPATH__abc_16259_n7403), .B(AES_CORE_DATAPATH__abc_16259_n7405), .Y(AES_CORE_DATAPATH__abc_16259_n7406) );
  AND2X2 AND2X2_2422 ( .A(AES_CORE_DATAPATH__abc_16259_n7408), .B(AES_CORE_CONTROL_UNIT_mode_cbc_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n7409) );
  AND2X2 AND2X2_2423 ( .A(AES_CORE_DATAPATH__abc_16259_n7407), .B(AES_CORE_DATAPATH__abc_16259_n7409), .Y(AES_CORE_DATAPATH__abc_16259_n7410) );
  AND2X2 AND2X2_2424 ( .A(AES_CORE_DATAPATH__abc_16259_n6101_bF_buf3), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_26_), .Y(AES_CORE_DATAPATH__abc_16259_n7411) );
  AND2X2 AND2X2_2425 ( .A(AES_CORE_DATAPATH__abc_16259_n7413), .B(AES_CORE_DATAPATH__abc_16259_n6056_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7414) );
  AND2X2 AND2X2_2426 ( .A(AES_CORE_DATAPATH__abc_16259_n3909), .B(AES_CORE_DATAPATH__abc_16259_n6053_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7415) );
  AND2X2 AND2X2_2427 ( .A(AES_CORE_DATAPATH__abc_16259_n7417), .B(AES_CORE_DATAPATH__abc_16259_n7418), .Y(AES_CORE_DATAPATH__abc_16259_n7419) );
  AND2X2 AND2X2_2428 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf8), .B(AES_CORE_DATAPATH__abc_16259_n7419), .Y(AES_CORE_DATAPATH__abc_16259_n7420) );
  AND2X2 AND2X2_2429 ( .A(AES_CORE_DATAPATH__abc_16259_n7421), .B(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n7422) );
  AND2X2 AND2X2_243 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf3), .B(AES_CORE_DATAPATH_iv_1__27_), .Y(AES_CORE_DATAPATH__abc_16259_n2726) );
  AND2X2 AND2X2_2430 ( .A(AES_CORE_DATAPATH__abc_16259_n6044_bF_buf3), .B(AES_CORE_DATAPATH_col_0__27_), .Y(AES_CORE_DATAPATH__abc_16259_n7424) );
  AND2X2 AND2X2_2431 ( .A(AES_CORE_DATAPATH__abc_16259_n3949), .B(AES_CORE_DATAPATH__abc_16259_n6059_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7425) );
  AND2X2 AND2X2_2432 ( .A(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf5), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_27_), .Y(AES_CORE_DATAPATH__abc_16259_n7426) );
  AND2X2 AND2X2_2433 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf4), .B(AES_CORE_DATAPATH_bkp_0__27_), .Y(AES_CORE_DATAPATH__abc_16259_n7428) );
  AND2X2 AND2X2_2434 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1__27_), .Y(AES_CORE_DATAPATH__abc_16259_n7429) );
  AND2X2 AND2X2_2435 ( .A(AES_CORE_DATAPATH__abc_16259_n7432), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7433) );
  AND2X2 AND2X2_2436 ( .A(AES_CORE_DATAPATH__abc_16259_n7431), .B(AES_CORE_DATAPATH__abc_16259_n7433), .Y(AES_CORE_DATAPATH__abc_16259_n7434) );
  AND2X2 AND2X2_2437 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf3), .B(AES_CORE_DATAPATH_bkp_3__27_), .Y(AES_CORE_DATAPATH__abc_16259_n7435) );
  AND2X2 AND2X2_2438 ( .A(AES_CORE_DATAPATH__abc_16259_n7437), .B(AES_CORE_DATAPATH__abc_16259_n7438), .Y(AES_CORE_DATAPATH__abc_16259_n7439) );
  AND2X2 AND2X2_2439 ( .A(AES_CORE_DATAPATH__abc_16259_n3940), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7442) );
  AND2X2 AND2X2_244 ( .A(AES_CORE_DATAPATH__abc_16259_n2729), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n2730) );
  AND2X2 AND2X2_2440 ( .A(AES_CORE_DATAPATH__abc_16259_n7442), .B(AES_CORE_DATAPATH__abc_16259_n7441), .Y(AES_CORE_DATAPATH__abc_16259_n7443) );
  AND2X2 AND2X2_2441 ( .A(AES_CORE_DATAPATH__abc_16259_n7446), .B(AES_CORE_DATAPATH__abc_16259_n7447), .Y(AES_CORE_DATAPATH__abc_16259_n7448) );
  AND2X2 AND2X2_2442 ( .A(AES_CORE_DATAPATH__abc_16259_n7440), .B(AES_CORE_DATAPATH__abc_16259_n7450), .Y(AES_CORE_DATAPATH__abc_16259_n7451) );
  AND2X2 AND2X2_2443 ( .A(AES_CORE_DATAPATH__abc_16259_n7453), .B(AES_CORE_DATAPATH__abc_16259_n6092_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n7454) );
  AND2X2 AND2X2_2444 ( .A(AES_CORE_DATAPATH__abc_16259_n7452), .B(AES_CORE_DATAPATH__abc_16259_n7454), .Y(AES_CORE_DATAPATH__abc_16259_n7455) );
  AND2X2 AND2X2_2445 ( .A(AES_CORE_DATAPATH__abc_16259_n7457), .B(AES_CORE_CONTROL_UNIT_mode_cbc_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n7458) );
  AND2X2 AND2X2_2446 ( .A(AES_CORE_DATAPATH__abc_16259_n7456), .B(AES_CORE_DATAPATH__abc_16259_n7458), .Y(AES_CORE_DATAPATH__abc_16259_n7459) );
  AND2X2 AND2X2_2447 ( .A(AES_CORE_DATAPATH__abc_16259_n6101_bF_buf2), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_27_), .Y(AES_CORE_DATAPATH__abc_16259_n7460) );
  AND2X2 AND2X2_2448 ( .A(AES_CORE_DATAPATH__abc_16259_n7462), .B(AES_CORE_DATAPATH__abc_16259_n6056_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n7463) );
  AND2X2 AND2X2_2449 ( .A(AES_CORE_DATAPATH__abc_16259_n3949), .B(AES_CORE_DATAPATH__abc_16259_n6053_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n7464) );
  AND2X2 AND2X2_245 ( .A(AES_CORE_DATAPATH__abc_16259_n2728), .B(AES_CORE_DATAPATH__abc_16259_n2730), .Y(AES_CORE_DATAPATH__abc_16259_n2731_1) );
  AND2X2 AND2X2_2450 ( .A(AES_CORE_DATAPATH__abc_16259_n7466), .B(AES_CORE_DATAPATH__abc_16259_n7467), .Y(AES_CORE_DATAPATH__abc_16259_n7468) );
  AND2X2 AND2X2_2451 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf7), .B(AES_CORE_DATAPATH__abc_16259_n7468), .Y(AES_CORE_DATAPATH__abc_16259_n7469) );
  AND2X2 AND2X2_2452 ( .A(AES_CORE_DATAPATH__abc_16259_n7470), .B(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n7471) );
  AND2X2 AND2X2_2453 ( .A(AES_CORE_DATAPATH__abc_16259_n6044_bF_buf2), .B(AES_CORE_DATAPATH_col_0__28_), .Y(AES_CORE_DATAPATH__abc_16259_n7473) );
  AND2X2 AND2X2_2454 ( .A(AES_CORE_DATAPATH__abc_16259_n3980), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n7475) );
  AND2X2 AND2X2_2455 ( .A(AES_CORE_DATAPATH__abc_16259_n7475), .B(AES_CORE_DATAPATH__abc_16259_n7474), .Y(AES_CORE_DATAPATH__abc_16259_n7476) );
  AND2X2 AND2X2_2456 ( .A(AES_CORE_DATAPATH__abc_16259_n7478), .B(AES_CORE_DATAPATH__abc_16259_n6059_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n7479) );
  AND2X2 AND2X2_2457 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf3), .B(AES_CORE_DATAPATH_bkp_0__28_), .Y(AES_CORE_DATAPATH__abc_16259_n7483) );
  AND2X2 AND2X2_2458 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf2), .B(AES_CORE_DATAPATH_bkp_1__28_), .Y(AES_CORE_DATAPATH__abc_16259_n7484) );
  AND2X2 AND2X2_2459 ( .A(AES_CORE_DATAPATH__abc_16259_n7487), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7488) );
  AND2X2 AND2X2_246 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf3), .B(AES_CORE_DATAPATH_iv_3__27_), .Y(AES_CORE_DATAPATH__abc_16259_n2732) );
  AND2X2 AND2X2_2460 ( .A(AES_CORE_DATAPATH__abc_16259_n7486), .B(AES_CORE_DATAPATH__abc_16259_n7488), .Y(AES_CORE_DATAPATH__abc_16259_n7489) );
  AND2X2 AND2X2_2461 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf2), .B(AES_CORE_DATAPATH_bkp_3__28_), .Y(AES_CORE_DATAPATH__abc_16259_n7490) );
  AND2X2 AND2X2_2462 ( .A(AES_CORE_DATAPATH__abc_16259_n7492), .B(AES_CORE_DATAPATH__abc_16259_n7493), .Y(AES_CORE_DATAPATH__abc_16259_n7494) );
  AND2X2 AND2X2_2463 ( .A(AES_CORE_DATAPATH__abc_16259_n7497), .B(AES_CORE_DATAPATH__abc_16259_n7480), .Y(AES_CORE_DATAPATH__abc_16259_n7498) );
  AND2X2 AND2X2_2464 ( .A(AES_CORE_DATAPATH__abc_16259_n7496), .B(AES_CORE_DATAPATH__abc_16259_n7499), .Y(AES_CORE_DATAPATH__abc_16259_n7500) );
  AND2X2 AND2X2_2465 ( .A(AES_CORE_DATAPATH__abc_16259_n7502), .B(AES_CORE_DATAPATH__abc_16259_n6092_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n7503) );
  AND2X2 AND2X2_2466 ( .A(AES_CORE_DATAPATH__abc_16259_n7501), .B(AES_CORE_DATAPATH__abc_16259_n7503), .Y(AES_CORE_DATAPATH__abc_16259_n7504) );
  AND2X2 AND2X2_2467 ( .A(AES_CORE_DATAPATH__abc_16259_n7506), .B(AES_CORE_CONTROL_UNIT_mode_cbc_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n7507) );
  AND2X2 AND2X2_2468 ( .A(AES_CORE_DATAPATH__abc_16259_n7505), .B(AES_CORE_DATAPATH__abc_16259_n7507), .Y(AES_CORE_DATAPATH__abc_16259_n7508) );
  AND2X2 AND2X2_2469 ( .A(AES_CORE_DATAPATH__abc_16259_n6101_bF_buf1), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_28_), .Y(AES_CORE_DATAPATH__abc_16259_n7509) );
  AND2X2 AND2X2_247 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf3), .B(AES_CORE_DATAPATH_iv_0__28_), .Y(AES_CORE_DATAPATH__abc_16259_n2734) );
  AND2X2 AND2X2_2470 ( .A(AES_CORE_DATAPATH__abc_16259_n7511), .B(AES_CORE_DATAPATH__abc_16259_n6056_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n7512) );
  AND2X2 AND2X2_2471 ( .A(AES_CORE_DATAPATH__abc_16259_n3989), .B(AES_CORE_DATAPATH__abc_16259_n6053_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n7513) );
  AND2X2 AND2X2_2472 ( .A(AES_CORE_DATAPATH__abc_16259_n7515), .B(AES_CORE_DATAPATH__abc_16259_n7516), .Y(AES_CORE_DATAPATH__abc_16259_n7517) );
  AND2X2 AND2X2_2473 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf6), .B(AES_CORE_DATAPATH__abc_16259_n7517), .Y(AES_CORE_DATAPATH__abc_16259_n7518) );
  AND2X2 AND2X2_2474 ( .A(AES_CORE_DATAPATH__abc_16259_n7519), .B(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n7520) );
  AND2X2 AND2X2_2475 ( .A(AES_CORE_DATAPATH__abc_16259_n6044_bF_buf1), .B(AES_CORE_DATAPATH_col_0__29_), .Y(AES_CORE_DATAPATH__abc_16259_n7522) );
  AND2X2 AND2X2_2476 ( .A(AES_CORE_DATAPATH__abc_16259_n4029), .B(AES_CORE_DATAPATH__abc_16259_n6059_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n7523) );
  AND2X2 AND2X2_2477 ( .A(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf2), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_29_), .Y(AES_CORE_DATAPATH__abc_16259_n7524) );
  AND2X2 AND2X2_2478 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf2), .B(AES_CORE_DATAPATH_bkp_0__29_), .Y(AES_CORE_DATAPATH__abc_16259_n7526) );
  AND2X2 AND2X2_2479 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf1), .B(AES_CORE_DATAPATH_bkp_1__29_), .Y(AES_CORE_DATAPATH__abc_16259_n7527) );
  AND2X2 AND2X2_248 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf2), .B(AES_CORE_DATAPATH_iv_1__28_), .Y(AES_CORE_DATAPATH__abc_16259_n2735_1) );
  AND2X2 AND2X2_2480 ( .A(AES_CORE_DATAPATH__abc_16259_n7530), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n7531) );
  AND2X2 AND2X2_2481 ( .A(AES_CORE_DATAPATH__abc_16259_n7529), .B(AES_CORE_DATAPATH__abc_16259_n7531), .Y(AES_CORE_DATAPATH__abc_16259_n7532) );
  AND2X2 AND2X2_2482 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf1), .B(AES_CORE_DATAPATH_bkp_3__29_), .Y(AES_CORE_DATAPATH__abc_16259_n7533) );
  AND2X2 AND2X2_2483 ( .A(AES_CORE_DATAPATH__abc_16259_n7535), .B(AES_CORE_DATAPATH__abc_16259_n7536), .Y(AES_CORE_DATAPATH__abc_16259_n7537) );
  AND2X2 AND2X2_2484 ( .A(AES_CORE_DATAPATH__abc_16259_n4020), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n7540) );
  AND2X2 AND2X2_2485 ( .A(AES_CORE_DATAPATH__abc_16259_n7540), .B(AES_CORE_DATAPATH__abc_16259_n7539), .Y(AES_CORE_DATAPATH__abc_16259_n7541) );
  AND2X2 AND2X2_2486 ( .A(AES_CORE_DATAPATH__abc_16259_n7544), .B(AES_CORE_DATAPATH__abc_16259_n7545), .Y(AES_CORE_DATAPATH__abc_16259_n7546) );
  AND2X2 AND2X2_2487 ( .A(AES_CORE_DATAPATH__abc_16259_n7538), .B(AES_CORE_DATAPATH__abc_16259_n7548), .Y(AES_CORE_DATAPATH__abc_16259_n7549) );
  AND2X2 AND2X2_2488 ( .A(AES_CORE_DATAPATH__abc_16259_n7551), .B(AES_CORE_DATAPATH__abc_16259_n6092_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n7552) );
  AND2X2 AND2X2_2489 ( .A(AES_CORE_DATAPATH__abc_16259_n7550), .B(AES_CORE_DATAPATH__abc_16259_n7552), .Y(AES_CORE_DATAPATH__abc_16259_n7553) );
  AND2X2 AND2X2_249 ( .A(AES_CORE_DATAPATH__abc_16259_n2738), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n2739) );
  AND2X2 AND2X2_2490 ( .A(AES_CORE_DATAPATH__abc_16259_n7555), .B(AES_CORE_CONTROL_UNIT_mode_cbc_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7556) );
  AND2X2 AND2X2_2491 ( .A(AES_CORE_DATAPATH__abc_16259_n7554), .B(AES_CORE_DATAPATH__abc_16259_n7556), .Y(AES_CORE_DATAPATH__abc_16259_n7557) );
  AND2X2 AND2X2_2492 ( .A(AES_CORE_DATAPATH__abc_16259_n6101_bF_buf0), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_29_), .Y(AES_CORE_DATAPATH__abc_16259_n7558) );
  AND2X2 AND2X2_2493 ( .A(AES_CORE_DATAPATH__abc_16259_n7560), .B(AES_CORE_DATAPATH__abc_16259_n6056_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n7561) );
  AND2X2 AND2X2_2494 ( .A(AES_CORE_DATAPATH__abc_16259_n4029), .B(AES_CORE_DATAPATH__abc_16259_n6053_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n7562) );
  AND2X2 AND2X2_2495 ( .A(AES_CORE_DATAPATH__abc_16259_n7564), .B(AES_CORE_DATAPATH__abc_16259_n7565), .Y(AES_CORE_DATAPATH__abc_16259_n7566) );
  AND2X2 AND2X2_2496 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf5), .B(AES_CORE_DATAPATH__abc_16259_n7566), .Y(AES_CORE_DATAPATH__abc_16259_n7567) );
  AND2X2 AND2X2_2497 ( .A(AES_CORE_DATAPATH__abc_16259_n7568), .B(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7569) );
  AND2X2 AND2X2_2498 ( .A(AES_CORE_DATAPATH__abc_16259_n6044_bF_buf0), .B(AES_CORE_DATAPATH_col_0__30_), .Y(AES_CORE_DATAPATH__abc_16259_n7571) );
  AND2X2 AND2X2_2499 ( .A(AES_CORE_DATAPATH__abc_16259_n4069), .B(AES_CORE_DATAPATH__abc_16259_n6059_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n7572) );
  AND2X2 AND2X2_25 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n105), .B(AES_CORE_CONTROL_UNIT__abc_15841_n103), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n106_1) );
  AND2X2 AND2X2_250 ( .A(AES_CORE_DATAPATH__abc_16259_n2737_1), .B(AES_CORE_DATAPATH__abc_16259_n2739), .Y(AES_CORE_DATAPATH__abc_16259_n2740) );
  AND2X2 AND2X2_2500 ( .A(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf0), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_30_), .Y(AES_CORE_DATAPATH__abc_16259_n7573) );
  AND2X2 AND2X2_2501 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf1), .B(AES_CORE_DATAPATH_bkp_0__30_), .Y(AES_CORE_DATAPATH__abc_16259_n7575) );
  AND2X2 AND2X2_2502 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf0), .B(AES_CORE_DATAPATH_bkp_1__30_), .Y(AES_CORE_DATAPATH__abc_16259_n7576) );
  AND2X2 AND2X2_2503 ( .A(AES_CORE_DATAPATH__abc_16259_n7579), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n7580) );
  AND2X2 AND2X2_2504 ( .A(AES_CORE_DATAPATH__abc_16259_n7578), .B(AES_CORE_DATAPATH__abc_16259_n7580), .Y(AES_CORE_DATAPATH__abc_16259_n7581) );
  AND2X2 AND2X2_2505 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf0), .B(AES_CORE_DATAPATH_bkp_3__30_), .Y(AES_CORE_DATAPATH__abc_16259_n7582) );
  AND2X2 AND2X2_2506 ( .A(AES_CORE_DATAPATH__abc_16259_n7585), .B(AES_CORE_DATAPATH__abc_16259_n7584), .Y(AES_CORE_DATAPATH__abc_16259_n7586) );
  AND2X2 AND2X2_2507 ( .A(AES_CORE_DATAPATH__abc_16259_n4060), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n7589) );
  AND2X2 AND2X2_2508 ( .A(AES_CORE_DATAPATH__abc_16259_n7589), .B(AES_CORE_DATAPATH__abc_16259_n7588), .Y(AES_CORE_DATAPATH__abc_16259_n7590) );
  AND2X2 AND2X2_2509 ( .A(AES_CORE_DATAPATH__abc_16259_n7593), .B(AES_CORE_DATAPATH__abc_16259_n7594), .Y(AES_CORE_DATAPATH__abc_16259_n7595) );
  AND2X2 AND2X2_251 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf2), .B(AES_CORE_DATAPATH_iv_3__28_), .Y(AES_CORE_DATAPATH__abc_16259_n2741) );
  AND2X2 AND2X2_2510 ( .A(AES_CORE_DATAPATH__abc_16259_n7587), .B(AES_CORE_DATAPATH__abc_16259_n7597), .Y(AES_CORE_DATAPATH__abc_16259_n7598) );
  AND2X2 AND2X2_2511 ( .A(AES_CORE_DATAPATH__abc_16259_n7600), .B(AES_CORE_DATAPATH__abc_16259_n6092_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7601) );
  AND2X2 AND2X2_2512 ( .A(AES_CORE_DATAPATH__abc_16259_n7599), .B(AES_CORE_DATAPATH__abc_16259_n7601), .Y(AES_CORE_DATAPATH__abc_16259_n7602) );
  AND2X2 AND2X2_2513 ( .A(AES_CORE_DATAPATH__abc_16259_n7604), .B(AES_CORE_CONTROL_UNIT_mode_cbc_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7605) );
  AND2X2 AND2X2_2514 ( .A(AES_CORE_DATAPATH__abc_16259_n7603), .B(AES_CORE_DATAPATH__abc_16259_n7605), .Y(AES_CORE_DATAPATH__abc_16259_n7606) );
  AND2X2 AND2X2_2515 ( .A(AES_CORE_DATAPATH__abc_16259_n6101_bF_buf4), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_30_), .Y(AES_CORE_DATAPATH__abc_16259_n7607) );
  AND2X2 AND2X2_2516 ( .A(AES_CORE_DATAPATH__abc_16259_n7609), .B(AES_CORE_DATAPATH__abc_16259_n6056_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7610) );
  AND2X2 AND2X2_2517 ( .A(AES_CORE_DATAPATH__abc_16259_n4069), .B(AES_CORE_DATAPATH__abc_16259_n6053_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7611) );
  AND2X2 AND2X2_2518 ( .A(AES_CORE_DATAPATH__abc_16259_n7613), .B(AES_CORE_DATAPATH__abc_16259_n7614), .Y(AES_CORE_DATAPATH__abc_16259_n7615) );
  AND2X2 AND2X2_2519 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n7615), .Y(AES_CORE_DATAPATH__abc_16259_n7616) );
  AND2X2 AND2X2_252 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf2), .B(AES_CORE_DATAPATH_iv_0__29_), .Y(AES_CORE_DATAPATH__abc_16259_n2743) );
  AND2X2 AND2X2_2520 ( .A(AES_CORE_DATAPATH__abc_16259_n7617), .B(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7618) );
  AND2X2 AND2X2_2521 ( .A(AES_CORE_DATAPATH__abc_16259_n6044_bF_buf4), .B(AES_CORE_DATAPATH_col_0__31_), .Y(AES_CORE_DATAPATH__abc_16259_n7620) );
  AND2X2 AND2X2_2522 ( .A(AES_CORE_DATAPATH__abc_16259_n4109), .B(AES_CORE_DATAPATH__abc_16259_n6059_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7621) );
  AND2X2 AND2X2_2523 ( .A(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf5), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_31_), .Y(AES_CORE_DATAPATH__abc_16259_n7622) );
  AND2X2 AND2X2_2524 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf0), .B(AES_CORE_DATAPATH_bkp_0__31_), .Y(AES_CORE_DATAPATH__abc_16259_n7624) );
  AND2X2 AND2X2_2525 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf7), .B(AES_CORE_DATAPATH_bkp_1__31_), .Y(AES_CORE_DATAPATH__abc_16259_n7625) );
  AND2X2 AND2X2_2526 ( .A(AES_CORE_DATAPATH__abc_16259_n7628), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n7629) );
  AND2X2 AND2X2_2527 ( .A(AES_CORE_DATAPATH__abc_16259_n7627), .B(AES_CORE_DATAPATH__abc_16259_n7629), .Y(AES_CORE_DATAPATH__abc_16259_n7630) );
  AND2X2 AND2X2_2528 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf7), .B(AES_CORE_DATAPATH_bkp_3__31_), .Y(AES_CORE_DATAPATH__abc_16259_n7631) );
  AND2X2 AND2X2_2529 ( .A(AES_CORE_DATAPATH__abc_16259_n7633), .B(AES_CORE_DATAPATH__abc_16259_n7634), .Y(AES_CORE_DATAPATH__abc_16259_n7635) );
  AND2X2 AND2X2_253 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf1), .B(AES_CORE_DATAPATH_iv_1__29_), .Y(AES_CORE_DATAPATH__abc_16259_n2744) );
  AND2X2 AND2X2_2530 ( .A(AES_CORE_DATAPATH__abc_16259_n4100), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n7638) );
  AND2X2 AND2X2_2531 ( .A(AES_CORE_DATAPATH__abc_16259_n7638), .B(AES_CORE_DATAPATH__abc_16259_n7637), .Y(AES_CORE_DATAPATH__abc_16259_n7639) );
  AND2X2 AND2X2_2532 ( .A(AES_CORE_DATAPATH__abc_16259_n7642), .B(AES_CORE_DATAPATH__abc_16259_n7643), .Y(AES_CORE_DATAPATH__abc_16259_n7644) );
  AND2X2 AND2X2_2533 ( .A(AES_CORE_DATAPATH__abc_16259_n7636), .B(AES_CORE_DATAPATH__abc_16259_n7646), .Y(AES_CORE_DATAPATH__abc_16259_n7647) );
  AND2X2 AND2X2_2534 ( .A(AES_CORE_DATAPATH__abc_16259_n7649), .B(AES_CORE_DATAPATH__abc_16259_n6092_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7650) );
  AND2X2 AND2X2_2535 ( .A(AES_CORE_DATAPATH__abc_16259_n7648), .B(AES_CORE_DATAPATH__abc_16259_n7650), .Y(AES_CORE_DATAPATH__abc_16259_n7651) );
  AND2X2 AND2X2_2536 ( .A(AES_CORE_DATAPATH__abc_16259_n7653), .B(AES_CORE_CONTROL_UNIT_mode_cbc_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n7654) );
  AND2X2 AND2X2_2537 ( .A(AES_CORE_DATAPATH__abc_16259_n7652), .B(AES_CORE_DATAPATH__abc_16259_n7654), .Y(AES_CORE_DATAPATH__abc_16259_n7655) );
  AND2X2 AND2X2_2538 ( .A(AES_CORE_DATAPATH__abc_16259_n6101_bF_buf3), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_31_), .Y(AES_CORE_DATAPATH__abc_16259_n7656) );
  AND2X2 AND2X2_2539 ( .A(AES_CORE_DATAPATH__abc_16259_n7658), .B(AES_CORE_DATAPATH__abc_16259_n6056_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7659) );
  AND2X2 AND2X2_254 ( .A(AES_CORE_DATAPATH__abc_16259_n2747), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n2748) );
  AND2X2 AND2X2_2540 ( .A(AES_CORE_DATAPATH__abc_16259_n4109), .B(AES_CORE_DATAPATH__abc_16259_n6053_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7660) );
  AND2X2 AND2X2_2541 ( .A(AES_CORE_DATAPATH__abc_16259_n7662), .B(AES_CORE_DATAPATH__abc_16259_n7663), .Y(AES_CORE_DATAPATH__abc_16259_n7664) );
  AND2X2 AND2X2_2542 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n7664), .Y(AES_CORE_DATAPATH__abc_16259_n7665) );
  AND2X2 AND2X2_2543 ( .A(AES_CORE_DATAPATH__abc_16259_n7666), .B(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n7667) );
  AND2X2 AND2X2_2544 ( .A(AES_CORE_DATAPATH__abc_16259_n7669_bF_buf4), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_64_), .Y(AES_CORE_DATAPATH__abc_16259_n7670) );
  AND2X2 AND2X2_2545 ( .A(AES_CORE_DATAPATH__abc_16259_n7671), .B(AES_CORE_DATAPATH__abc_16259_n7672), .Y(AES_CORE_DATAPATH__abc_16259_n7673) );
  AND2X2 AND2X2_2546 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n7673), .Y(AES_CORE_DATAPATH__abc_16259_n7674) );
  AND2X2 AND2X2_2547 ( .A(AES_CORE_DATAPATH__abc_16259_n7675), .B(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7676) );
  AND2X2 AND2X2_2548 ( .A(AES_CORE_DATAPATH__abc_16259_n7669_bF_buf3), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_65_), .Y(AES_CORE_DATAPATH__abc_16259_n7678) );
  AND2X2 AND2X2_2549 ( .A(AES_CORE_DATAPATH__abc_16259_n7679), .B(AES_CORE_DATAPATH__abc_16259_n7680), .Y(AES_CORE_DATAPATH__abc_16259_n7681) );
  AND2X2 AND2X2_255 ( .A(AES_CORE_DATAPATH__abc_16259_n2746_1), .B(AES_CORE_DATAPATH__abc_16259_n2748), .Y(AES_CORE_DATAPATH__abc_16259_n2749) );
  AND2X2 AND2X2_2550 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n7681), .Y(AES_CORE_DATAPATH__abc_16259_n7682) );
  AND2X2 AND2X2_2551 ( .A(AES_CORE_DATAPATH__abc_16259_n7683), .B(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n7684) );
  AND2X2 AND2X2_2552 ( .A(AES_CORE_DATAPATH__abc_16259_n7669_bF_buf2), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_66_), .Y(AES_CORE_DATAPATH__abc_16259_n7686) );
  AND2X2 AND2X2_2553 ( .A(AES_CORE_DATAPATH__abc_16259_n7687), .B(AES_CORE_DATAPATH__abc_16259_n7688), .Y(AES_CORE_DATAPATH__abc_16259_n7689) );
  AND2X2 AND2X2_2554 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n7689), .Y(AES_CORE_DATAPATH__abc_16259_n7690) );
  AND2X2 AND2X2_2555 ( .A(AES_CORE_DATAPATH__abc_16259_n7691), .B(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n7692) );
  AND2X2 AND2X2_2556 ( .A(AES_CORE_DATAPATH__abc_16259_n7669_bF_buf1), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_67_), .Y(AES_CORE_DATAPATH__abc_16259_n7694) );
  AND2X2 AND2X2_2557 ( .A(AES_CORE_DATAPATH__abc_16259_n7695), .B(AES_CORE_DATAPATH__abc_16259_n7696), .Y(AES_CORE_DATAPATH__abc_16259_n7697) );
  AND2X2 AND2X2_2558 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf9), .B(AES_CORE_DATAPATH__abc_16259_n7697), .Y(AES_CORE_DATAPATH__abc_16259_n7698) );
  AND2X2 AND2X2_2559 ( .A(AES_CORE_DATAPATH__abc_16259_n7699), .B(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n7700) );
  AND2X2 AND2X2_256 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf1), .B(AES_CORE_DATAPATH_iv_3__29_), .Y(AES_CORE_DATAPATH__abc_16259_n2750) );
  AND2X2 AND2X2_2560 ( .A(AES_CORE_DATAPATH__abc_16259_n7669_bF_buf0), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_68_), .Y(AES_CORE_DATAPATH__abc_16259_n7702) );
  AND2X2 AND2X2_2561 ( .A(AES_CORE_DATAPATH__abc_16259_n7703), .B(AES_CORE_DATAPATH__abc_16259_n7704), .Y(AES_CORE_DATAPATH__abc_16259_n7705) );
  AND2X2 AND2X2_2562 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf8), .B(AES_CORE_DATAPATH__abc_16259_n7705), .Y(AES_CORE_DATAPATH__abc_16259_n7706) );
  AND2X2 AND2X2_2563 ( .A(AES_CORE_DATAPATH__abc_16259_n7707), .B(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n7708) );
  AND2X2 AND2X2_2564 ( .A(AES_CORE_DATAPATH__abc_16259_n7669_bF_buf4), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_69_), .Y(AES_CORE_DATAPATH__abc_16259_n7710) );
  AND2X2 AND2X2_2565 ( .A(AES_CORE_DATAPATH__abc_16259_n7711), .B(AES_CORE_DATAPATH__abc_16259_n7712), .Y(AES_CORE_DATAPATH__abc_16259_n7713) );
  AND2X2 AND2X2_2566 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf7), .B(AES_CORE_DATAPATH__abc_16259_n7713), .Y(AES_CORE_DATAPATH__abc_16259_n7714) );
  AND2X2 AND2X2_2567 ( .A(AES_CORE_DATAPATH__abc_16259_n7715), .B(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7716) );
  AND2X2 AND2X2_2568 ( .A(AES_CORE_DATAPATH__abc_16259_n7669_bF_buf3), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_70_), .Y(AES_CORE_DATAPATH__abc_16259_n7718) );
  AND2X2 AND2X2_2569 ( .A(AES_CORE_DATAPATH__abc_16259_n7719), .B(AES_CORE_DATAPATH__abc_16259_n7720), .Y(AES_CORE_DATAPATH__abc_16259_n7721) );
  AND2X2 AND2X2_257 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf1), .B(AES_CORE_DATAPATH_iv_0__30_), .Y(AES_CORE_DATAPATH__abc_16259_n2752_1) );
  AND2X2 AND2X2_2570 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf6), .B(AES_CORE_DATAPATH__abc_16259_n7721), .Y(AES_CORE_DATAPATH__abc_16259_n7722) );
  AND2X2 AND2X2_2571 ( .A(AES_CORE_DATAPATH__abc_16259_n7723), .B(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7724) );
  AND2X2 AND2X2_2572 ( .A(AES_CORE_DATAPATH__abc_16259_n7669_bF_buf2), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_71_), .Y(AES_CORE_DATAPATH__abc_16259_n7726) );
  AND2X2 AND2X2_2573 ( .A(AES_CORE_DATAPATH__abc_16259_n7727), .B(AES_CORE_DATAPATH__abc_16259_n7728), .Y(AES_CORE_DATAPATH__abc_16259_n7729) );
  AND2X2 AND2X2_2574 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf5), .B(AES_CORE_DATAPATH__abc_16259_n7729), .Y(AES_CORE_DATAPATH__abc_16259_n7730) );
  AND2X2 AND2X2_2575 ( .A(AES_CORE_DATAPATH__abc_16259_n7731), .B(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n7732) );
  AND2X2 AND2X2_2576 ( .A(AES_CORE_DATAPATH__abc_16259_n7669_bF_buf1), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_72_), .Y(AES_CORE_DATAPATH__abc_16259_n7734) );
  AND2X2 AND2X2_2577 ( .A(AES_CORE_DATAPATH__abc_16259_n7735), .B(AES_CORE_DATAPATH__abc_16259_n7736), .Y(AES_CORE_DATAPATH__abc_16259_n7737) );
  AND2X2 AND2X2_2578 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n7737), .Y(AES_CORE_DATAPATH__abc_16259_n7738) );
  AND2X2 AND2X2_2579 ( .A(AES_CORE_DATAPATH__abc_16259_n7739), .B(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n7740) );
  AND2X2 AND2X2_258 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf0), .B(AES_CORE_DATAPATH_iv_1__30_), .Y(AES_CORE_DATAPATH__abc_16259_n2753_1) );
  AND2X2 AND2X2_2580 ( .A(AES_CORE_DATAPATH__abc_16259_n7669_bF_buf0), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_73_), .Y(AES_CORE_DATAPATH__abc_16259_n7742) );
  AND2X2 AND2X2_2581 ( .A(AES_CORE_DATAPATH__abc_16259_n7743), .B(AES_CORE_DATAPATH__abc_16259_n7744), .Y(AES_CORE_DATAPATH__abc_16259_n7745) );
  AND2X2 AND2X2_2582 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n7745), .Y(AES_CORE_DATAPATH__abc_16259_n7746) );
  AND2X2 AND2X2_2583 ( .A(AES_CORE_DATAPATH__abc_16259_n7747), .B(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n7748) );
  AND2X2 AND2X2_2584 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf10), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_10_), .Y(AES_CORE_DATAPATH__abc_16259_n7753) );
  AND2X2 AND2X2_2585 ( .A(AES_CORE_DATAPATH__abc_16259_n7752), .B(AES_CORE_DATAPATH__abc_16259_n7754), .Y(AES_CORE_DATAPATH__abc_16259_n7755) );
  AND2X2 AND2X2_2586 ( .A(AES_CORE_DATAPATH__abc_16259_n6602), .B(AES_CORE_DATAPATH__abc_16259_n7756), .Y(AES_CORE_DATAPATH__abc_16259_n7757) );
  AND2X2 AND2X2_2587 ( .A(AES_CORE_DATAPATH__abc_16259_n7757), .B(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7758) );
  AND2X2 AND2X2_2588 ( .A(AES_CORE_DATAPATH__abc_16259_n7759), .B(AES_CORE_DATAPATH__abc_16259_n7750), .Y(AES_CORE_DATAPATH__0col_1__31_0__10_) );
  AND2X2 AND2X2_2589 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf8), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_11_), .Y(AES_CORE_DATAPATH__abc_16259_n7763) );
  AND2X2 AND2X2_259 ( .A(AES_CORE_DATAPATH__abc_16259_n2756_1), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n2757) );
  AND2X2 AND2X2_2590 ( .A(AES_CORE_DATAPATH__abc_16259_n7762), .B(AES_CORE_DATAPATH__abc_16259_n7764), .Y(AES_CORE_DATAPATH__abc_16259_n7765) );
  AND2X2 AND2X2_2591 ( .A(AES_CORE_DATAPATH__abc_16259_n6657), .B(AES_CORE_DATAPATH__abc_16259_n7766), .Y(AES_CORE_DATAPATH__abc_16259_n7767) );
  AND2X2 AND2X2_2592 ( .A(AES_CORE_DATAPATH__abc_16259_n7767), .B(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7768) );
  AND2X2 AND2X2_2593 ( .A(AES_CORE_DATAPATH__abc_16259_n7769), .B(AES_CORE_DATAPATH__abc_16259_n7770), .Y(AES_CORE_DATAPATH__0col_1__31_0__11_) );
  AND2X2 AND2X2_2594 ( .A(AES_CORE_DATAPATH__abc_16259_n7669_bF_buf4), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_76_), .Y(AES_CORE_DATAPATH__abc_16259_n7772) );
  AND2X2 AND2X2_2595 ( .A(AES_CORE_DATAPATH__abc_16259_n7773), .B(AES_CORE_DATAPATH__abc_16259_n7774), .Y(AES_CORE_DATAPATH__abc_16259_n7775) );
  AND2X2 AND2X2_2596 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n7775), .Y(AES_CORE_DATAPATH__abc_16259_n7776) );
  AND2X2 AND2X2_2597 ( .A(AES_CORE_DATAPATH__abc_16259_n7777), .B(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n7778) );
  AND2X2 AND2X2_2598 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf5), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_13_), .Y(AES_CORE_DATAPATH__abc_16259_n7782) );
  AND2X2 AND2X2_2599 ( .A(AES_CORE_DATAPATH__abc_16259_n7781), .B(AES_CORE_DATAPATH__abc_16259_n7783), .Y(AES_CORE_DATAPATH__abc_16259_n7784) );
  AND2X2 AND2X2_26 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n106_1), .B(AES_CORE_CONTROL_UNIT__abc_15841_n84_1), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n107) );
  AND2X2 AND2X2_260 ( .A(AES_CORE_DATAPATH__abc_16259_n2755_1), .B(AES_CORE_DATAPATH__abc_16259_n2757), .Y(AES_CORE_DATAPATH__abc_16259_n2758) );
  AND2X2 AND2X2_2600 ( .A(AES_CORE_DATAPATH__abc_16259_n6760), .B(AES_CORE_DATAPATH__abc_16259_n7785), .Y(AES_CORE_DATAPATH__abc_16259_n7786) );
  AND2X2 AND2X2_2601 ( .A(AES_CORE_DATAPATH__abc_16259_n7786), .B(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n7787) );
  AND2X2 AND2X2_2602 ( .A(AES_CORE_DATAPATH__abc_16259_n7788), .B(AES_CORE_DATAPATH__abc_16259_n7789), .Y(AES_CORE_DATAPATH__0col_1__31_0__13_) );
  AND2X2 AND2X2_2603 ( .A(AES_CORE_DATAPATH__abc_16259_n7669_bF_buf3), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_78_), .Y(AES_CORE_DATAPATH__abc_16259_n7791) );
  AND2X2 AND2X2_2604 ( .A(AES_CORE_DATAPATH__abc_16259_n7792), .B(AES_CORE_DATAPATH__abc_16259_n7793), .Y(AES_CORE_DATAPATH__abc_16259_n7794) );
  AND2X2 AND2X2_2605 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n7794), .Y(AES_CORE_DATAPATH__abc_16259_n7795) );
  AND2X2 AND2X2_2606 ( .A(AES_CORE_DATAPATH__abc_16259_n7796), .B(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7797) );
  AND2X2 AND2X2_2607 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf2), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_15_), .Y(AES_CORE_DATAPATH__abc_16259_n7801) );
  AND2X2 AND2X2_2608 ( .A(AES_CORE_DATAPATH__abc_16259_n7800), .B(AES_CORE_DATAPATH__abc_16259_n7802), .Y(AES_CORE_DATAPATH__abc_16259_n7803) );
  AND2X2 AND2X2_2609 ( .A(AES_CORE_DATAPATH__abc_16259_n6863), .B(AES_CORE_DATAPATH__abc_16259_n7804), .Y(AES_CORE_DATAPATH__abc_16259_n7805) );
  AND2X2 AND2X2_261 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf0), .B(AES_CORE_DATAPATH_iv_3__30_), .Y(AES_CORE_DATAPATH__abc_16259_n2759) );
  AND2X2 AND2X2_2610 ( .A(AES_CORE_DATAPATH__abc_16259_n7805), .B(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7806) );
  AND2X2 AND2X2_2611 ( .A(AES_CORE_DATAPATH__abc_16259_n7807), .B(AES_CORE_DATAPATH__abc_16259_n7808), .Y(AES_CORE_DATAPATH__0col_1__31_0__15_) );
  AND2X2 AND2X2_2612 ( .A(AES_CORE_DATAPATH__abc_16259_n7669_bF_buf2), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_80_), .Y(AES_CORE_DATAPATH__abc_16259_n7810) );
  AND2X2 AND2X2_2613 ( .A(AES_CORE_DATAPATH__abc_16259_n7811), .B(AES_CORE_DATAPATH__abc_16259_n7812), .Y(AES_CORE_DATAPATH__abc_16259_n7813) );
  AND2X2 AND2X2_2614 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n7813), .Y(AES_CORE_DATAPATH__abc_16259_n7814) );
  AND2X2 AND2X2_2615 ( .A(AES_CORE_DATAPATH__abc_16259_n7815), .B(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n7816) );
  AND2X2 AND2X2_2616 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf14), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_49_), .Y(AES_CORE_DATAPATH__abc_16259_n7820) );
  AND2X2 AND2X2_2617 ( .A(AES_CORE_DATAPATH__abc_16259_n7819), .B(AES_CORE_DATAPATH__abc_16259_n7821), .Y(AES_CORE_DATAPATH__abc_16259_n7822) );
  AND2X2 AND2X2_2618 ( .A(AES_CORE_DATAPATH__abc_16259_n6966), .B(AES_CORE_DATAPATH__abc_16259_n7823), .Y(AES_CORE_DATAPATH__abc_16259_n7824) );
  AND2X2 AND2X2_2619 ( .A(AES_CORE_DATAPATH__abc_16259_n7824), .B(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n7825) );
  AND2X2 AND2X2_262 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf0), .B(AES_CORE_DATAPATH_iv_0__31_), .Y(AES_CORE_DATAPATH__abc_16259_n2761) );
  AND2X2 AND2X2_2620 ( .A(AES_CORE_DATAPATH__abc_16259_n7826), .B(AES_CORE_DATAPATH__abc_16259_n7827), .Y(AES_CORE_DATAPATH__0col_1__31_0__17_) );
  AND2X2 AND2X2_2621 ( .A(AES_CORE_DATAPATH__abc_16259_n7669_bF_buf1), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_82_), .Y(AES_CORE_DATAPATH__abc_16259_n7829) );
  AND2X2 AND2X2_2622 ( .A(AES_CORE_DATAPATH__abc_16259_n7830), .B(AES_CORE_DATAPATH__abc_16259_n7831), .Y(AES_CORE_DATAPATH__abc_16259_n7832) );
  AND2X2 AND2X2_2623 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf9), .B(AES_CORE_DATAPATH__abc_16259_n7832), .Y(AES_CORE_DATAPATH__abc_16259_n7833) );
  AND2X2 AND2X2_2624 ( .A(AES_CORE_DATAPATH__abc_16259_n7834), .B(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7835) );
  AND2X2 AND2X2_2625 ( .A(AES_CORE_DATAPATH__abc_16259_n7669_bF_buf0), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_83_), .Y(AES_CORE_DATAPATH__abc_16259_n7837) );
  AND2X2 AND2X2_2626 ( .A(AES_CORE_DATAPATH__abc_16259_n7838), .B(AES_CORE_DATAPATH__abc_16259_n7839), .Y(AES_CORE_DATAPATH__abc_16259_n7840) );
  AND2X2 AND2X2_2627 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf8), .B(AES_CORE_DATAPATH__abc_16259_n7840), .Y(AES_CORE_DATAPATH__abc_16259_n7841) );
  AND2X2 AND2X2_2628 ( .A(AES_CORE_DATAPATH__abc_16259_n7842), .B(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7843) );
  AND2X2 AND2X2_2629 ( .A(AES_CORE_DATAPATH__abc_16259_n7669_bF_buf4), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_84_), .Y(AES_CORE_DATAPATH__abc_16259_n7845) );
  AND2X2 AND2X2_263 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf7), .B(AES_CORE_DATAPATH_iv_1__31_), .Y(AES_CORE_DATAPATH__abc_16259_n2762_1) );
  AND2X2 AND2X2_2630 ( .A(AES_CORE_DATAPATH__abc_16259_n7846), .B(AES_CORE_DATAPATH__abc_16259_n7847), .Y(AES_CORE_DATAPATH__abc_16259_n7848) );
  AND2X2 AND2X2_2631 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf7), .B(AES_CORE_DATAPATH__abc_16259_n7848), .Y(AES_CORE_DATAPATH__abc_16259_n7849) );
  AND2X2 AND2X2_2632 ( .A(AES_CORE_DATAPATH__abc_16259_n7850), .B(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n7851) );
  AND2X2 AND2X2_2633 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf9), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_53_), .Y(AES_CORE_DATAPATH__abc_16259_n7855) );
  AND2X2 AND2X2_2634 ( .A(AES_CORE_DATAPATH__abc_16259_n7854), .B(AES_CORE_DATAPATH__abc_16259_n7856), .Y(AES_CORE_DATAPATH__abc_16259_n7857) );
  AND2X2 AND2X2_2635 ( .A(AES_CORE_DATAPATH__abc_16259_n7167), .B(AES_CORE_DATAPATH__abc_16259_n7858), .Y(AES_CORE_DATAPATH__abc_16259_n7859) );
  AND2X2 AND2X2_2636 ( .A(AES_CORE_DATAPATH__abc_16259_n7859), .B(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n7860) );
  AND2X2 AND2X2_2637 ( .A(AES_CORE_DATAPATH__abc_16259_n7861), .B(AES_CORE_DATAPATH__abc_16259_n7862), .Y(AES_CORE_DATAPATH__0col_1__31_0__21_) );
  AND2X2 AND2X2_2638 ( .A(AES_CORE_DATAPATH__abc_16259_n7669_bF_buf3), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_86_), .Y(AES_CORE_DATAPATH__abc_16259_n7864) );
  AND2X2 AND2X2_2639 ( .A(AES_CORE_DATAPATH__abc_16259_n7865), .B(AES_CORE_DATAPATH__abc_16259_n7866), .Y(AES_CORE_DATAPATH__abc_16259_n7867) );
  AND2X2 AND2X2_264 ( .A(AES_CORE_DATAPATH__abc_16259_n2765), .B(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n2766) );
  AND2X2 AND2X2_2640 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf6), .B(AES_CORE_DATAPATH__abc_16259_n7867), .Y(AES_CORE_DATAPATH__abc_16259_n7868) );
  AND2X2 AND2X2_2641 ( .A(AES_CORE_DATAPATH__abc_16259_n7869), .B(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n7870) );
  AND2X2 AND2X2_2642 ( .A(AES_CORE_DATAPATH__abc_16259_n7669_bF_buf2), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_87_), .Y(AES_CORE_DATAPATH__abc_16259_n7872) );
  AND2X2 AND2X2_2643 ( .A(AES_CORE_DATAPATH__abc_16259_n7873), .B(AES_CORE_DATAPATH__abc_16259_n7874), .Y(AES_CORE_DATAPATH__abc_16259_n7875) );
  AND2X2 AND2X2_2644 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf5), .B(AES_CORE_DATAPATH__abc_16259_n7875), .Y(AES_CORE_DATAPATH__abc_16259_n7876) );
  AND2X2 AND2X2_2645 ( .A(AES_CORE_DATAPATH__abc_16259_n7877), .B(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7878) );
  AND2X2 AND2X2_2646 ( .A(AES_CORE_DATAPATH__abc_16259_n7669_bF_buf1), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_88_), .Y(AES_CORE_DATAPATH__abc_16259_n7880) );
  AND2X2 AND2X2_2647 ( .A(AES_CORE_DATAPATH__abc_16259_n7881), .B(AES_CORE_DATAPATH__abc_16259_n7882), .Y(AES_CORE_DATAPATH__abc_16259_n7883) );
  AND2X2 AND2X2_2648 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n7883), .Y(AES_CORE_DATAPATH__abc_16259_n7884) );
  AND2X2 AND2X2_2649 ( .A(AES_CORE_DATAPATH__abc_16259_n7885), .B(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7886) );
  AND2X2 AND2X2_265 ( .A(AES_CORE_DATAPATH__abc_16259_n2764_1), .B(AES_CORE_DATAPATH__abc_16259_n2766), .Y(AES_CORE_DATAPATH__abc_16259_n2767) );
  AND2X2 AND2X2_2650 ( .A(AES_CORE_DATAPATH__abc_16259_n7669_bF_buf0), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_89_), .Y(AES_CORE_DATAPATH__abc_16259_n7888) );
  AND2X2 AND2X2_2651 ( .A(AES_CORE_DATAPATH__abc_16259_n7889), .B(AES_CORE_DATAPATH__abc_16259_n7890), .Y(AES_CORE_DATAPATH__abc_16259_n7891) );
  AND2X2 AND2X2_2652 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n7891), .Y(AES_CORE_DATAPATH__abc_16259_n7892) );
  AND2X2 AND2X2_2653 ( .A(AES_CORE_DATAPATH__abc_16259_n7893), .B(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n7894) );
  AND2X2 AND2X2_2654 ( .A(AES_CORE_DATAPATH__abc_16259_n7669_bF_buf4), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_90_), .Y(AES_CORE_DATAPATH__abc_16259_n7896) );
  AND2X2 AND2X2_2655 ( .A(AES_CORE_DATAPATH__abc_16259_n7897), .B(AES_CORE_DATAPATH__abc_16259_n7898), .Y(AES_CORE_DATAPATH__abc_16259_n7899) );
  AND2X2 AND2X2_2656 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n7899), .Y(AES_CORE_DATAPATH__abc_16259_n7900) );
  AND2X2 AND2X2_2657 ( .A(AES_CORE_DATAPATH__abc_16259_n7901), .B(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n7902) );
  AND2X2 AND2X2_2658 ( .A(AES_CORE_DATAPATH__abc_16259_n7669_bF_buf3), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_91_), .Y(AES_CORE_DATAPATH__abc_16259_n7904) );
  AND2X2 AND2X2_2659 ( .A(AES_CORE_DATAPATH__abc_16259_n7905), .B(AES_CORE_DATAPATH__abc_16259_n7906), .Y(AES_CORE_DATAPATH__abc_16259_n7907) );
  AND2X2 AND2X2_266 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf7), .B(AES_CORE_DATAPATH_iv_3__31_), .Y(AES_CORE_DATAPATH__abc_16259_n2768) );
  AND2X2 AND2X2_2660 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n7907), .Y(AES_CORE_DATAPATH__abc_16259_n7908) );
  AND2X2 AND2X2_2661 ( .A(AES_CORE_DATAPATH__abc_16259_n7909), .B(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n7910) );
  AND2X2 AND2X2_2662 ( .A(AES_CORE_DATAPATH__abc_16259_n7669_bF_buf2), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_92_), .Y(AES_CORE_DATAPATH__abc_16259_n7912) );
  AND2X2 AND2X2_2663 ( .A(AES_CORE_DATAPATH__abc_16259_n7913), .B(AES_CORE_DATAPATH__abc_16259_n7914), .Y(AES_CORE_DATAPATH__abc_16259_n7915) );
  AND2X2 AND2X2_2664 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n7915), .Y(AES_CORE_DATAPATH__abc_16259_n7916) );
  AND2X2 AND2X2_2665 ( .A(AES_CORE_DATAPATH__abc_16259_n7917), .B(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n7918) );
  AND2X2 AND2X2_2666 ( .A(AES_CORE_DATAPATH__abc_16259_n7669_bF_buf1), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_93_), .Y(AES_CORE_DATAPATH__abc_16259_n7920) );
  AND2X2 AND2X2_2667 ( .A(AES_CORE_DATAPATH__abc_16259_n7921), .B(AES_CORE_DATAPATH__abc_16259_n7922), .Y(AES_CORE_DATAPATH__abc_16259_n7923) );
  AND2X2 AND2X2_2668 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf9), .B(AES_CORE_DATAPATH__abc_16259_n7923), .Y(AES_CORE_DATAPATH__abc_16259_n7924) );
  AND2X2 AND2X2_2669 ( .A(AES_CORE_DATAPATH__abc_16259_n7925), .B(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7926) );
  AND2X2 AND2X2_267 ( .A(AES_CORE_DATAPATH__abc_16259_n2775_1), .B(AES_CORE_DATAPATH__abc_16259_n2779_1), .Y(AES_CORE_DATAPATH__abc_16259_n2780) );
  AND2X2 AND2X2_2670 ( .A(AES_CORE_DATAPATH__abc_16259_n7669_bF_buf0), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_94_), .Y(AES_CORE_DATAPATH__abc_16259_n7928) );
  AND2X2 AND2X2_2671 ( .A(AES_CORE_DATAPATH__abc_16259_n7929), .B(AES_CORE_DATAPATH__abc_16259_n7930), .Y(AES_CORE_DATAPATH__abc_16259_n7931) );
  AND2X2 AND2X2_2672 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf8), .B(AES_CORE_DATAPATH__abc_16259_n7931), .Y(AES_CORE_DATAPATH__abc_16259_n7932) );
  AND2X2 AND2X2_2673 ( .A(AES_CORE_DATAPATH__abc_16259_n7933), .B(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7934) );
  AND2X2 AND2X2_2674 ( .A(AES_CORE_DATAPATH__abc_16259_n7669_bF_buf4), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_95_), .Y(AES_CORE_DATAPATH__abc_16259_n7936) );
  AND2X2 AND2X2_2675 ( .A(AES_CORE_DATAPATH__abc_16259_n7937), .B(AES_CORE_DATAPATH__abc_16259_n7938), .Y(AES_CORE_DATAPATH__abc_16259_n7939) );
  AND2X2 AND2X2_2676 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf7), .B(AES_CORE_DATAPATH__abc_16259_n7939), .Y(AES_CORE_DATAPATH__abc_16259_n7940) );
  AND2X2 AND2X2_2677 ( .A(AES_CORE_DATAPATH__abc_16259_n7941), .B(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n7942) );
  AND2X2 AND2X2_2678 ( .A(AES_CORE_DATAPATH__abc_16259_n7944_bF_buf4), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_32_), .Y(AES_CORE_DATAPATH__abc_16259_n7945) );
  AND2X2 AND2X2_2679 ( .A(AES_CORE_DATAPATH__abc_16259_n7946), .B(AES_CORE_DATAPATH__abc_16259_n7947), .Y(AES_CORE_DATAPATH__abc_16259_n7948) );
  AND2X2 AND2X2_268 ( .A(AES_CORE_DATAPATH__abc_16259_n2772_1), .B(AES_CORE_DATAPATH__abc_16259_n2777_1), .Y(AES_CORE_DATAPATH__abc_16259_n2781_1) );
  AND2X2 AND2X2_2680 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf6), .B(AES_CORE_DATAPATH__abc_16259_n7948), .Y(AES_CORE_DATAPATH__abc_16259_n7949) );
  AND2X2 AND2X2_2681 ( .A(AES_CORE_DATAPATH__abc_16259_n7950), .B(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7951) );
  AND2X2 AND2X2_2682 ( .A(AES_CORE_DATAPATH__abc_16259_n7944_bF_buf3), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_33_), .Y(AES_CORE_DATAPATH__abc_16259_n7953) );
  AND2X2 AND2X2_2683 ( .A(AES_CORE_DATAPATH__abc_16259_n7954), .B(AES_CORE_DATAPATH__abc_16259_n7955), .Y(AES_CORE_DATAPATH__abc_16259_n7956) );
  AND2X2 AND2X2_2684 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf5), .B(AES_CORE_DATAPATH__abc_16259_n7956), .Y(AES_CORE_DATAPATH__abc_16259_n7957) );
  AND2X2 AND2X2_2685 ( .A(AES_CORE_DATAPATH__abc_16259_n7958), .B(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n7959) );
  AND2X2 AND2X2_2686 ( .A(AES_CORE_DATAPATH__abc_16259_n7944_bF_buf2), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_34_), .Y(AES_CORE_DATAPATH__abc_16259_n7961) );
  AND2X2 AND2X2_2687 ( .A(AES_CORE_DATAPATH__abc_16259_n7962), .B(AES_CORE_DATAPATH__abc_16259_n7963), .Y(AES_CORE_DATAPATH__abc_16259_n7964) );
  AND2X2 AND2X2_2688 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n7964), .Y(AES_CORE_DATAPATH__abc_16259_n7965) );
  AND2X2 AND2X2_2689 ( .A(AES_CORE_DATAPATH__abc_16259_n7966), .B(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n7967) );
  AND2X2 AND2X2_269 ( .A(AES_CORE_DATAPATH__abc_16259_n2781_1), .B(AES_CORE_DATAPATH__abc_16259_n2771_1), .Y(AES_CORE_DATAPATH__abc_16259_n2782) );
  AND2X2 AND2X2_2690 ( .A(AES_CORE_DATAPATH__abc_16259_n7944_bF_buf1), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_35_), .Y(AES_CORE_DATAPATH__abc_16259_n7969) );
  AND2X2 AND2X2_2691 ( .A(AES_CORE_DATAPATH__abc_16259_n7970), .B(AES_CORE_DATAPATH__abc_16259_n7971), .Y(AES_CORE_DATAPATH__abc_16259_n7972) );
  AND2X2 AND2X2_2692 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n7972), .Y(AES_CORE_DATAPATH__abc_16259_n7973) );
  AND2X2 AND2X2_2693 ( .A(AES_CORE_DATAPATH__abc_16259_n7974), .B(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n7975) );
  AND2X2 AND2X2_2694 ( .A(AES_CORE_DATAPATH__abc_16259_n7944_bF_buf0), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_36_), .Y(AES_CORE_DATAPATH__abc_16259_n7977) );
  AND2X2 AND2X2_2695 ( .A(AES_CORE_DATAPATH__abc_16259_n7978), .B(AES_CORE_DATAPATH__abc_16259_n7979), .Y(AES_CORE_DATAPATH__abc_16259_n7980) );
  AND2X2 AND2X2_2696 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n7980), .Y(AES_CORE_DATAPATH__abc_16259_n7981) );
  AND2X2 AND2X2_2697 ( .A(AES_CORE_DATAPATH__abc_16259_n7982), .B(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n7983) );
  AND2X2 AND2X2_2698 ( .A(AES_CORE_DATAPATH__abc_16259_n7944_bF_buf4), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_37_), .Y(AES_CORE_DATAPATH__abc_16259_n7985) );
  AND2X2 AND2X2_2699 ( .A(AES_CORE_DATAPATH__abc_16259_n7986), .B(AES_CORE_DATAPATH__abc_16259_n7987), .Y(AES_CORE_DATAPATH__abc_16259_n7988) );
  AND2X2 AND2X2_27 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n107), .B(AES_CORE_CONTROL_UNIT_state_14_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n108) );
  AND2X2 AND2X2_270 ( .A(AES_CORE_DATAPATH__abc_16259_n2782_bF_buf4), .B(AES_CORE_DATAPATH_col_3__0_), .Y(AES_CORE_DATAPATH__abc_16259_n2783) );
  AND2X2 AND2X2_2700 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n7988), .Y(AES_CORE_DATAPATH__abc_16259_n7989) );
  AND2X2 AND2X2_2701 ( .A(AES_CORE_DATAPATH__abc_16259_n7990), .B(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7991) );
  AND2X2 AND2X2_2702 ( .A(AES_CORE_DATAPATH__abc_16259_n7944_bF_buf3), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_38_), .Y(AES_CORE_DATAPATH__abc_16259_n7993) );
  AND2X2 AND2X2_2703 ( .A(AES_CORE_DATAPATH__abc_16259_n7994), .B(AES_CORE_DATAPATH__abc_16259_n7995), .Y(AES_CORE_DATAPATH__abc_16259_n7996) );
  AND2X2 AND2X2_2704 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n7996), .Y(AES_CORE_DATAPATH__abc_16259_n7997) );
  AND2X2 AND2X2_2705 ( .A(AES_CORE_DATAPATH__abc_16259_n7998), .B(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7999) );
  AND2X2 AND2X2_2706 ( .A(AES_CORE_DATAPATH__abc_16259_n7944_bF_buf2), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_39_), .Y(AES_CORE_DATAPATH__abc_16259_n8001) );
  AND2X2 AND2X2_2707 ( .A(AES_CORE_DATAPATH__abc_16259_n8002), .B(AES_CORE_DATAPATH__abc_16259_n8003), .Y(AES_CORE_DATAPATH__abc_16259_n8004) );
  AND2X2 AND2X2_2708 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf9), .B(AES_CORE_DATAPATH__abc_16259_n8004), .Y(AES_CORE_DATAPATH__abc_16259_n8005) );
  AND2X2 AND2X2_2709 ( .A(AES_CORE_DATAPATH__abc_16259_n8006), .B(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n8007) );
  AND2X2 AND2X2_271 ( .A(AES_CORE_DATAPATH__abc_16259_n2771_1), .B(AES_CORE_DATAPATH__abc_16259_n2777_1), .Y(AES_CORE_DATAPATH__abc_16259_n2785) );
  AND2X2 AND2X2_2710 ( .A(AES_CORE_DATAPATH__abc_16259_n7944_bF_buf1), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_40_), .Y(AES_CORE_DATAPATH__abc_16259_n8009) );
  AND2X2 AND2X2_2711 ( .A(AES_CORE_DATAPATH__abc_16259_n8010), .B(AES_CORE_DATAPATH__abc_16259_n8011), .Y(AES_CORE_DATAPATH__abc_16259_n8012) );
  AND2X2 AND2X2_2712 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf8), .B(AES_CORE_DATAPATH__abc_16259_n8012), .Y(AES_CORE_DATAPATH__abc_16259_n8013) );
  AND2X2 AND2X2_2713 ( .A(AES_CORE_DATAPATH__abc_16259_n8014), .B(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n8015) );
  AND2X2 AND2X2_2714 ( .A(AES_CORE_DATAPATH__abc_16259_n7944_bF_buf0), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_41_), .Y(AES_CORE_DATAPATH__abc_16259_n8017) );
  AND2X2 AND2X2_2715 ( .A(AES_CORE_DATAPATH__abc_16259_n8018), .B(AES_CORE_DATAPATH__abc_16259_n8019), .Y(AES_CORE_DATAPATH__abc_16259_n8020) );
  AND2X2 AND2X2_2716 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf7), .B(AES_CORE_DATAPATH__abc_16259_n8020), .Y(AES_CORE_DATAPATH__abc_16259_n8021) );
  AND2X2 AND2X2_2717 ( .A(AES_CORE_DATAPATH__abc_16259_n8022), .B(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n8023) );
  AND2X2 AND2X2_2718 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf2), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_106_), .Y(AES_CORE_DATAPATH__abc_16259_n8027) );
  AND2X2 AND2X2_2719 ( .A(AES_CORE_DATAPATH__abc_16259_n8026), .B(AES_CORE_DATAPATH__abc_16259_n8028), .Y(AES_CORE_DATAPATH__abc_16259_n8029) );
  AND2X2 AND2X2_272 ( .A(AES_CORE_DATAPATH__abc_16259_n2785), .B(AES_CORE_DATAPATH__abc_16259_n2784), .Y(AES_CORE_DATAPATH__abc_16259_n2786) );
  AND2X2 AND2X2_2720 ( .A(AES_CORE_DATAPATH__abc_16259_n6602), .B(AES_CORE_DATAPATH__abc_16259_n8030), .Y(AES_CORE_DATAPATH__abc_16259_n8031) );
  AND2X2 AND2X2_2721 ( .A(AES_CORE_DATAPATH__abc_16259_n8031), .B(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n8032) );
  AND2X2 AND2X2_2722 ( .A(AES_CORE_DATAPATH__abc_16259_n8033), .B(AES_CORE_DATAPATH__abc_16259_n8034), .Y(AES_CORE_DATAPATH__0col_2__31_0__10_) );
  AND2X2 AND2X2_2723 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf0), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_107_), .Y(AES_CORE_DATAPATH__abc_16259_n8039) );
  AND2X2 AND2X2_2724 ( .A(AES_CORE_DATAPATH__abc_16259_n8038), .B(AES_CORE_DATAPATH__abc_16259_n8040), .Y(AES_CORE_DATAPATH__abc_16259_n8041) );
  AND2X2 AND2X2_2725 ( .A(AES_CORE_DATAPATH__abc_16259_n6657), .B(AES_CORE_DATAPATH__abc_16259_n8042), .Y(AES_CORE_DATAPATH__abc_16259_n8043) );
  AND2X2 AND2X2_2726 ( .A(AES_CORE_DATAPATH__abc_16259_n8043), .B(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n8044) );
  AND2X2 AND2X2_2727 ( .A(AES_CORE_DATAPATH__abc_16259_n8045), .B(AES_CORE_DATAPATH__abc_16259_n8036), .Y(AES_CORE_DATAPATH__0col_2__31_0__11_) );
  AND2X2 AND2X2_2728 ( .A(AES_CORE_DATAPATH__abc_16259_n7944_bF_buf4), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_44_), .Y(AES_CORE_DATAPATH__abc_16259_n8047) );
  AND2X2 AND2X2_2729 ( .A(AES_CORE_DATAPATH__abc_16259_n8048), .B(AES_CORE_DATAPATH__abc_16259_n8049), .Y(AES_CORE_DATAPATH__abc_16259_n8050) );
  AND2X2 AND2X2_273 ( .A(AES_CORE_DATAPATH__abc_16259_n2786_bF_buf4), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_64_), .Y(AES_CORE_DATAPATH__abc_16259_n2787) );
  AND2X2 AND2X2_2730 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf6), .B(AES_CORE_DATAPATH__abc_16259_n8050), .Y(AES_CORE_DATAPATH__abc_16259_n8051) );
  AND2X2 AND2X2_2731 ( .A(AES_CORE_DATAPATH__abc_16259_n8052), .B(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n8053) );
  AND2X2 AND2X2_2732 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf12), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_109_), .Y(AES_CORE_DATAPATH__abc_16259_n8057) );
  AND2X2 AND2X2_2733 ( .A(AES_CORE_DATAPATH__abc_16259_n8056), .B(AES_CORE_DATAPATH__abc_16259_n8058), .Y(AES_CORE_DATAPATH__abc_16259_n8059) );
  AND2X2 AND2X2_2734 ( .A(AES_CORE_DATAPATH__abc_16259_n6760), .B(AES_CORE_DATAPATH__abc_16259_n8060), .Y(AES_CORE_DATAPATH__abc_16259_n8061) );
  AND2X2 AND2X2_2735 ( .A(AES_CORE_DATAPATH__abc_16259_n8061), .B(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n8062) );
  AND2X2 AND2X2_2736 ( .A(AES_CORE_DATAPATH__abc_16259_n8063), .B(AES_CORE_DATAPATH__abc_16259_n8064), .Y(AES_CORE_DATAPATH__0col_2__31_0__13_) );
  AND2X2 AND2X2_2737 ( .A(AES_CORE_DATAPATH__abc_16259_n7944_bF_buf3), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_46_), .Y(AES_CORE_DATAPATH__abc_16259_n8066) );
  AND2X2 AND2X2_2738 ( .A(AES_CORE_DATAPATH__abc_16259_n8067), .B(AES_CORE_DATAPATH__abc_16259_n8068), .Y(AES_CORE_DATAPATH__abc_16259_n8069) );
  AND2X2 AND2X2_2739 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf5), .B(AES_CORE_DATAPATH__abc_16259_n8069), .Y(AES_CORE_DATAPATH__abc_16259_n8070) );
  AND2X2 AND2X2_274 ( .A(AES_CORE_DATAPATH__abc_16259_n2781_1), .B(AES_CORE_DATAPATH__abc_16259_n2788), .Y(AES_CORE_DATAPATH__abc_16259_n2789) );
  AND2X2 AND2X2_2740 ( .A(AES_CORE_DATAPATH__abc_16259_n8071), .B(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n8072) );
  AND2X2 AND2X2_2741 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf9), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_111_), .Y(AES_CORE_DATAPATH__abc_16259_n8076) );
  AND2X2 AND2X2_2742 ( .A(AES_CORE_DATAPATH__abc_16259_n8075), .B(AES_CORE_DATAPATH__abc_16259_n8077), .Y(AES_CORE_DATAPATH__abc_16259_n8078) );
  AND2X2 AND2X2_2743 ( .A(AES_CORE_DATAPATH__abc_16259_n6863), .B(AES_CORE_DATAPATH__abc_16259_n8079), .Y(AES_CORE_DATAPATH__abc_16259_n8080) );
  AND2X2 AND2X2_2744 ( .A(AES_CORE_DATAPATH__abc_16259_n8080), .B(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n8081) );
  AND2X2 AND2X2_2745 ( .A(AES_CORE_DATAPATH__abc_16259_n8082), .B(AES_CORE_DATAPATH__abc_16259_n8083), .Y(AES_CORE_DATAPATH__0col_2__31_0__15_) );
  AND2X2 AND2X2_2746 ( .A(AES_CORE_DATAPATH__abc_16259_n7944_bF_buf2), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_48_), .Y(AES_CORE_DATAPATH__abc_16259_n8085) );
  AND2X2 AND2X2_2747 ( .A(AES_CORE_DATAPATH__abc_16259_n8086), .B(AES_CORE_DATAPATH__abc_16259_n8087), .Y(AES_CORE_DATAPATH__abc_16259_n8088) );
  AND2X2 AND2X2_2748 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n8088), .Y(AES_CORE_DATAPATH__abc_16259_n8089) );
  AND2X2 AND2X2_2749 ( .A(AES_CORE_DATAPATH__abc_16259_n8090), .B(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n8091) );
  AND2X2 AND2X2_275 ( .A(AES_CORE_DATAPATH__abc_16259_n2789_bF_buf4), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_32_), .Y(AES_CORE_DATAPATH__abc_16259_n2790) );
  AND2X2 AND2X2_2750 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf6), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_17_), .Y(AES_CORE_DATAPATH__abc_16259_n8095) );
  AND2X2 AND2X2_2751 ( .A(AES_CORE_DATAPATH__abc_16259_n8094), .B(AES_CORE_DATAPATH__abc_16259_n8096), .Y(AES_CORE_DATAPATH__abc_16259_n8097) );
  AND2X2 AND2X2_2752 ( .A(AES_CORE_DATAPATH__abc_16259_n6966), .B(AES_CORE_DATAPATH__abc_16259_n8098), .Y(AES_CORE_DATAPATH__abc_16259_n8099) );
  AND2X2 AND2X2_2753 ( .A(AES_CORE_DATAPATH__abc_16259_n8099), .B(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n8100) );
  AND2X2 AND2X2_2754 ( .A(AES_CORE_DATAPATH__abc_16259_n8101), .B(AES_CORE_DATAPATH__abc_16259_n8102), .Y(AES_CORE_DATAPATH__0col_2__31_0__17_) );
  AND2X2 AND2X2_2755 ( .A(AES_CORE_DATAPATH__abc_16259_n7944_bF_buf1), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_50_), .Y(AES_CORE_DATAPATH__abc_16259_n8104) );
  AND2X2 AND2X2_2756 ( .A(AES_CORE_DATAPATH__abc_16259_n8105), .B(AES_CORE_DATAPATH__abc_16259_n8106), .Y(AES_CORE_DATAPATH__abc_16259_n8107) );
  AND2X2 AND2X2_2757 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n8107), .Y(AES_CORE_DATAPATH__abc_16259_n8108) );
  AND2X2 AND2X2_2758 ( .A(AES_CORE_DATAPATH__abc_16259_n8109), .B(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n8110) );
  AND2X2 AND2X2_2759 ( .A(AES_CORE_DATAPATH__abc_16259_n7944_bF_buf0), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_51_), .Y(AES_CORE_DATAPATH__abc_16259_n8112) );
  AND2X2 AND2X2_276 ( .A(AES_CORE_DATAPATH__abc_16259_n2793_1), .B(AES_CORE_DATAPATH__abc_16259_n2780), .Y(AES_CORE_DATAPATH__abc_16259_n2794) );
  AND2X2 AND2X2_2760 ( .A(AES_CORE_DATAPATH__abc_16259_n8113), .B(AES_CORE_DATAPATH__abc_16259_n8114), .Y(AES_CORE_DATAPATH__abc_16259_n8115) );
  AND2X2 AND2X2_2761 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n8115), .Y(AES_CORE_DATAPATH__abc_16259_n8116) );
  AND2X2 AND2X2_2762 ( .A(AES_CORE_DATAPATH__abc_16259_n8117), .B(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n8118) );
  AND2X2 AND2X2_2763 ( .A(AES_CORE_DATAPATH__abc_16259_n7944_bF_buf4), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_52_), .Y(AES_CORE_DATAPATH__abc_16259_n8120) );
  AND2X2 AND2X2_2764 ( .A(AES_CORE_DATAPATH__abc_16259_n8121), .B(AES_CORE_DATAPATH__abc_16259_n8122), .Y(AES_CORE_DATAPATH__abc_16259_n8123) );
  AND2X2 AND2X2_2765 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n8123), .Y(AES_CORE_DATAPATH__abc_16259_n8124) );
  AND2X2 AND2X2_2766 ( .A(AES_CORE_DATAPATH__abc_16259_n8125), .B(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n8126) );
  AND2X2 AND2X2_2767 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf1), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_21_), .Y(AES_CORE_DATAPATH__abc_16259_n8130) );
  AND2X2 AND2X2_2768 ( .A(AES_CORE_DATAPATH__abc_16259_n8129), .B(AES_CORE_DATAPATH__abc_16259_n8131), .Y(AES_CORE_DATAPATH__abc_16259_n8132) );
  AND2X2 AND2X2_2769 ( .A(AES_CORE_DATAPATH__abc_16259_n7167), .B(AES_CORE_DATAPATH__abc_16259_n8133), .Y(AES_CORE_DATAPATH__abc_16259_n8134) );
  AND2X2 AND2X2_277 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__0_), .B(AES_CORE_DATAPATH_last_round_pp2_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n2797) );
  AND2X2 AND2X2_2770 ( .A(AES_CORE_DATAPATH__abc_16259_n8134), .B(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n8135) );
  AND2X2 AND2X2_2771 ( .A(AES_CORE_DATAPATH__abc_16259_n8136), .B(AES_CORE_DATAPATH__abc_16259_n8137), .Y(AES_CORE_DATAPATH__0col_2__31_0__21_) );
  AND2X2 AND2X2_2772 ( .A(AES_CORE_DATAPATH__abc_16259_n7944_bF_buf3), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_54_), .Y(AES_CORE_DATAPATH__abc_16259_n8139) );
  AND2X2 AND2X2_2773 ( .A(AES_CORE_DATAPATH__abc_16259_n8140), .B(AES_CORE_DATAPATH__abc_16259_n8141), .Y(AES_CORE_DATAPATH__abc_16259_n8142) );
  AND2X2 AND2X2_2774 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n8142), .Y(AES_CORE_DATAPATH__abc_16259_n8143) );
  AND2X2 AND2X2_2775 ( .A(AES_CORE_DATAPATH__abc_16259_n8144), .B(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n8145) );
  AND2X2 AND2X2_2776 ( .A(AES_CORE_DATAPATH__abc_16259_n7944_bF_buf2), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_55_), .Y(AES_CORE_DATAPATH__abc_16259_n8147) );
  AND2X2 AND2X2_2777 ( .A(AES_CORE_DATAPATH__abc_16259_n8148), .B(AES_CORE_DATAPATH__abc_16259_n8149), .Y(AES_CORE_DATAPATH__abc_16259_n8150) );
  AND2X2 AND2X2_2778 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf9), .B(AES_CORE_DATAPATH__abc_16259_n8150), .Y(AES_CORE_DATAPATH__abc_16259_n8151) );
  AND2X2 AND2X2_2779 ( .A(AES_CORE_DATAPATH__abc_16259_n8152), .B(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n8153) );
  AND2X2 AND2X2_278 ( .A(AES_CORE_DATAPATH__abc_16259_n2798_bF_buf4), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_0_), .Y(AES_CORE_DATAPATH__abc_16259_n2799) );
  AND2X2 AND2X2_2780 ( .A(AES_CORE_DATAPATH__abc_16259_n7944_bF_buf1), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_56_), .Y(AES_CORE_DATAPATH__abc_16259_n8155) );
  AND2X2 AND2X2_2781 ( .A(AES_CORE_DATAPATH__abc_16259_n8156), .B(AES_CORE_DATAPATH__abc_16259_n8157), .Y(AES_CORE_DATAPATH__abc_16259_n8158) );
  AND2X2 AND2X2_2782 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf8), .B(AES_CORE_DATAPATH__abc_16259_n8158), .Y(AES_CORE_DATAPATH__abc_16259_n8159) );
  AND2X2 AND2X2_2783 ( .A(AES_CORE_DATAPATH__abc_16259_n8160), .B(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n8161) );
  AND2X2 AND2X2_2784 ( .A(AES_CORE_DATAPATH__abc_16259_n7944_bF_buf0), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_57_), .Y(AES_CORE_DATAPATH__abc_16259_n8163) );
  AND2X2 AND2X2_2785 ( .A(AES_CORE_DATAPATH__abc_16259_n8164), .B(AES_CORE_DATAPATH__abc_16259_n8165), .Y(AES_CORE_DATAPATH__abc_16259_n8166) );
  AND2X2 AND2X2_2786 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf7), .B(AES_CORE_DATAPATH__abc_16259_n8166), .Y(AES_CORE_DATAPATH__abc_16259_n8167) );
  AND2X2 AND2X2_2787 ( .A(AES_CORE_DATAPATH__abc_16259_n8168), .B(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n8169) );
  AND2X2 AND2X2_2788 ( .A(AES_CORE_DATAPATH__abc_16259_n7944_bF_buf4), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_58_), .Y(AES_CORE_DATAPATH__abc_16259_n8171) );
  AND2X2 AND2X2_2789 ( .A(AES_CORE_DATAPATH__abc_16259_n8172), .B(AES_CORE_DATAPATH__abc_16259_n8173), .Y(AES_CORE_DATAPATH__abc_16259_n8174) );
  AND2X2 AND2X2_279 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf12), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf10), .Y(AES_CORE_DATAPATH__abc_16259_n2804_1) );
  AND2X2 AND2X2_2790 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf6), .B(AES_CORE_DATAPATH__abc_16259_n8174), .Y(AES_CORE_DATAPATH__abc_16259_n8175) );
  AND2X2 AND2X2_2791 ( .A(AES_CORE_DATAPATH__abc_16259_n8176), .B(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n8177) );
  AND2X2 AND2X2_2792 ( .A(AES_CORE_DATAPATH__abc_16259_n7944_bF_buf3), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_59_), .Y(AES_CORE_DATAPATH__abc_16259_n8179) );
  AND2X2 AND2X2_2793 ( .A(AES_CORE_DATAPATH__abc_16259_n8180), .B(AES_CORE_DATAPATH__abc_16259_n8181), .Y(AES_CORE_DATAPATH__abc_16259_n8182) );
  AND2X2 AND2X2_2794 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf5), .B(AES_CORE_DATAPATH__abc_16259_n8182), .Y(AES_CORE_DATAPATH__abc_16259_n8183) );
  AND2X2 AND2X2_2795 ( .A(AES_CORE_DATAPATH__abc_16259_n8184), .B(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n8185) );
  AND2X2 AND2X2_2796 ( .A(AES_CORE_DATAPATH__abc_16259_n7944_bF_buf2), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_60_), .Y(AES_CORE_DATAPATH__abc_16259_n8187) );
  AND2X2 AND2X2_2797 ( .A(AES_CORE_DATAPATH__abc_16259_n8188), .B(AES_CORE_DATAPATH__abc_16259_n8189), .Y(AES_CORE_DATAPATH__abc_16259_n8190) );
  AND2X2 AND2X2_2798 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n8190), .Y(AES_CORE_DATAPATH__abc_16259_n8191) );
  AND2X2 AND2X2_2799 ( .A(AES_CORE_DATAPATH__abc_16259_n8192), .B(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n8193) );
  AND2X2 AND2X2_28 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n112), .B(AES_CORE_CONTROL_UNIT_key_gen), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n113) );
  AND2X2 AND2X2_280 ( .A(AES_CORE_DATAPATH__abc_16259_n2808_1), .B(AES_CORE_DATAPATH__abc_16259_n2806_1), .Y(AES_CORE_DATAPATH__abc_16259_n2809) );
  AND2X2 AND2X2_2800 ( .A(AES_CORE_DATAPATH__abc_16259_n7944_bF_buf1), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_61_), .Y(AES_CORE_DATAPATH__abc_16259_n8195) );
  AND2X2 AND2X2_2801 ( .A(AES_CORE_DATAPATH__abc_16259_n8196), .B(AES_CORE_DATAPATH__abc_16259_n8197), .Y(AES_CORE_DATAPATH__abc_16259_n8198) );
  AND2X2 AND2X2_2802 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n8198), .Y(AES_CORE_DATAPATH__abc_16259_n8199) );
  AND2X2 AND2X2_2803 ( .A(AES_CORE_DATAPATH__abc_16259_n8200), .B(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n8201) );
  AND2X2 AND2X2_2804 ( .A(AES_CORE_DATAPATH__abc_16259_n7944_bF_buf0), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_62_), .Y(AES_CORE_DATAPATH__abc_16259_n8203) );
  AND2X2 AND2X2_2805 ( .A(AES_CORE_DATAPATH__abc_16259_n8204), .B(AES_CORE_DATAPATH__abc_16259_n8205), .Y(AES_CORE_DATAPATH__abc_16259_n8206) );
  AND2X2 AND2X2_2806 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n8206), .Y(AES_CORE_DATAPATH__abc_16259_n8207) );
  AND2X2 AND2X2_2807 ( .A(AES_CORE_DATAPATH__abc_16259_n8208), .B(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n8209) );
  AND2X2 AND2X2_2808 ( .A(AES_CORE_DATAPATH__abc_16259_n7944_bF_buf4), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_63_), .Y(AES_CORE_DATAPATH__abc_16259_n8211) );
  AND2X2 AND2X2_2809 ( .A(AES_CORE_DATAPATH__abc_16259_n8212), .B(AES_CORE_DATAPATH__abc_16259_n8213), .Y(AES_CORE_DATAPATH__abc_16259_n8214) );
  AND2X2 AND2X2_281 ( .A(AES_CORE_DATAPATH__abc_16259_n2809), .B(AES_CORE_DATAPATH__abc_16259_n2805), .Y(AES_CORE_DATAPATH__abc_16259_n2810_1) );
  AND2X2 AND2X2_2810 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n8214), .Y(AES_CORE_DATAPATH__abc_16259_n8215) );
  AND2X2 AND2X2_2811 ( .A(AES_CORE_DATAPATH__abc_16259_n8216), .B(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n8217) );
  AND2X2 AND2X2_2812 ( .A(AES_CORE_DATAPATH__abc_16259_n8219_bF_buf4), .B(AES_CORE_DATAPATH_col_3__0_), .Y(AES_CORE_DATAPATH__abc_16259_n8220) );
  AND2X2 AND2X2_2813 ( .A(AES_CORE_DATAPATH__abc_16259_n8221), .B(AES_CORE_DATAPATH__abc_16259_n8222), .Y(AES_CORE_DATAPATH__abc_16259_n8223) );
  AND2X2 AND2X2_2814 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n8223), .Y(AES_CORE_DATAPATH__abc_16259_n8224) );
  AND2X2 AND2X2_2815 ( .A(AES_CORE_DATAPATH__abc_16259_n8225), .B(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n8226) );
  AND2X2 AND2X2_2816 ( .A(AES_CORE_DATAPATH__abc_16259_n8219_bF_buf3), .B(AES_CORE_DATAPATH_col_3__1_), .Y(AES_CORE_DATAPATH__abc_16259_n8228) );
  AND2X2 AND2X2_2817 ( .A(AES_CORE_DATAPATH__abc_16259_n8229), .B(AES_CORE_DATAPATH__abc_16259_n8230), .Y(AES_CORE_DATAPATH__abc_16259_n8231) );
  AND2X2 AND2X2_2818 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf9), .B(AES_CORE_DATAPATH__abc_16259_n8231), .Y(AES_CORE_DATAPATH__abc_16259_n8232) );
  AND2X2 AND2X2_2819 ( .A(AES_CORE_DATAPATH__abc_16259_n8233), .B(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n8234) );
  AND2X2 AND2X2_282 ( .A(AES_CORE_CONTROL_UNIT_bypass_key_en), .B(AES_CORE_CONTROL_UNIT_key_out_sel_1_), .Y(AES_CORE_DATAPATH__abc_16259_n2812) );
  AND2X2 AND2X2_2820 ( .A(AES_CORE_DATAPATH__abc_16259_n8219_bF_buf2), .B(AES_CORE_DATAPATH_col_3__2_), .Y(AES_CORE_DATAPATH__abc_16259_n8236) );
  AND2X2 AND2X2_2821 ( .A(AES_CORE_DATAPATH__abc_16259_n8237), .B(AES_CORE_DATAPATH__abc_16259_n8238), .Y(AES_CORE_DATAPATH__abc_16259_n8239) );
  AND2X2 AND2X2_2822 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf8), .B(AES_CORE_DATAPATH__abc_16259_n8239), .Y(AES_CORE_DATAPATH__abc_16259_n8240) );
  AND2X2 AND2X2_2823 ( .A(AES_CORE_DATAPATH__abc_16259_n8241), .B(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n8242) );
  AND2X2 AND2X2_2824 ( .A(AES_CORE_DATAPATH__abc_16259_n8219_bF_buf1), .B(AES_CORE_DATAPATH_col_3__3_), .Y(AES_CORE_DATAPATH__abc_16259_n8244) );
  AND2X2 AND2X2_2825 ( .A(AES_CORE_DATAPATH__abc_16259_n8245), .B(AES_CORE_DATAPATH__abc_16259_n8246), .Y(AES_CORE_DATAPATH__abc_16259_n8247) );
  AND2X2 AND2X2_2826 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf7), .B(AES_CORE_DATAPATH__abc_16259_n8247), .Y(AES_CORE_DATAPATH__abc_16259_n8248) );
  AND2X2 AND2X2_2827 ( .A(AES_CORE_DATAPATH__abc_16259_n8249), .B(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n8250) );
  AND2X2 AND2X2_2828 ( .A(AES_CORE_DATAPATH__abc_16259_n8219_bF_buf0), .B(AES_CORE_DATAPATH_col_3__4_), .Y(AES_CORE_DATAPATH__abc_16259_n8252) );
  AND2X2 AND2X2_2829 ( .A(AES_CORE_DATAPATH__abc_16259_n8253), .B(AES_CORE_DATAPATH__abc_16259_n8254), .Y(AES_CORE_DATAPATH__abc_16259_n8255) );
  AND2X2 AND2X2_283 ( .A(AES_CORE_DATAPATH__abc_16259_n2811), .B(AES_CORE_DATAPATH__abc_16259_n2814), .Y(AES_CORE_DATAPATH__abc_16259_n2815) );
  AND2X2 AND2X2_2830 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf6), .B(AES_CORE_DATAPATH__abc_16259_n8255), .Y(AES_CORE_DATAPATH__abc_16259_n8256) );
  AND2X2 AND2X2_2831 ( .A(AES_CORE_DATAPATH__abc_16259_n8257), .B(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n8258) );
  AND2X2 AND2X2_2832 ( .A(AES_CORE_DATAPATH__abc_16259_n8219_bF_buf4), .B(AES_CORE_DATAPATH_col_3__5_), .Y(AES_CORE_DATAPATH__abc_16259_n8260) );
  AND2X2 AND2X2_2833 ( .A(AES_CORE_DATAPATH__abc_16259_n8261), .B(AES_CORE_DATAPATH__abc_16259_n8262), .Y(AES_CORE_DATAPATH__abc_16259_n8263) );
  AND2X2 AND2X2_2834 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf5), .B(AES_CORE_DATAPATH__abc_16259_n8263), .Y(AES_CORE_DATAPATH__abc_16259_n8264) );
  AND2X2 AND2X2_2835 ( .A(AES_CORE_DATAPATH__abc_16259_n8265), .B(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n8266) );
  AND2X2 AND2X2_2836 ( .A(AES_CORE_DATAPATH__abc_16259_n8219_bF_buf3), .B(AES_CORE_DATAPATH_col_3__6_), .Y(AES_CORE_DATAPATH__abc_16259_n8268) );
  AND2X2 AND2X2_2837 ( .A(AES_CORE_DATAPATH__abc_16259_n8269), .B(AES_CORE_DATAPATH__abc_16259_n8270), .Y(AES_CORE_DATAPATH__abc_16259_n8271) );
  AND2X2 AND2X2_2838 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n8271), .Y(AES_CORE_DATAPATH__abc_16259_n8272) );
  AND2X2 AND2X2_2839 ( .A(AES_CORE_DATAPATH__abc_16259_n8273), .B(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n8274) );
  AND2X2 AND2X2_284 ( .A(AES_CORE_DATAPATH__abc_16259_n2819), .B(AES_CORE_DATAPATH__abc_16259_n2817), .Y(AES_CORE_DATAPATH__abc_16259_n2820) );
  AND2X2 AND2X2_2840 ( .A(AES_CORE_DATAPATH__abc_16259_n8219_bF_buf2), .B(AES_CORE_DATAPATH_col_3__7_), .Y(AES_CORE_DATAPATH__abc_16259_n8276) );
  AND2X2 AND2X2_2841 ( .A(AES_CORE_DATAPATH__abc_16259_n8277), .B(AES_CORE_DATAPATH__abc_16259_n8278), .Y(AES_CORE_DATAPATH__abc_16259_n8279) );
  AND2X2 AND2X2_2842 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n8279), .Y(AES_CORE_DATAPATH__abc_16259_n8280) );
  AND2X2 AND2X2_2843 ( .A(AES_CORE_DATAPATH__abc_16259_n8281), .B(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n8282) );
  AND2X2 AND2X2_2844 ( .A(AES_CORE_DATAPATH__abc_16259_n8219_bF_buf1), .B(AES_CORE_DATAPATH_col_3__8_), .Y(AES_CORE_DATAPATH__abc_16259_n8284) );
  AND2X2 AND2X2_2845 ( .A(AES_CORE_DATAPATH__abc_16259_n8285), .B(AES_CORE_DATAPATH__abc_16259_n8286), .Y(AES_CORE_DATAPATH__abc_16259_n8287) );
  AND2X2 AND2X2_2846 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n8287), .Y(AES_CORE_DATAPATH__abc_16259_n8288) );
  AND2X2 AND2X2_2847 ( .A(AES_CORE_DATAPATH__abc_16259_n8289), .B(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n8290) );
  AND2X2 AND2X2_2848 ( .A(AES_CORE_DATAPATH__abc_16259_n8219_bF_buf0), .B(AES_CORE_DATAPATH_col_3__9_), .Y(AES_CORE_DATAPATH__abc_16259_n8292) );
  AND2X2 AND2X2_2849 ( .A(AES_CORE_DATAPATH__abc_16259_n8293), .B(AES_CORE_DATAPATH__abc_16259_n8294), .Y(AES_CORE_DATAPATH__abc_16259_n8295) );
  AND2X2 AND2X2_285 ( .A(AES_CORE_CONTROL_UNIT_bypass_key_en), .B(AES_CORE_CONTROL_UNIT_key_out_sel_0_), .Y(AES_CORE_DATAPATH__abc_16259_n2822_1) );
  AND2X2 AND2X2_2850 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n8295), .Y(AES_CORE_DATAPATH__abc_16259_n8296) );
  AND2X2 AND2X2_2851 ( .A(AES_CORE_DATAPATH__abc_16259_n8297), .B(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n8298) );
  AND2X2 AND2X2_2852 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf9), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_74_), .Y(AES_CORE_DATAPATH__abc_16259_n8302) );
  AND2X2 AND2X2_2853 ( .A(AES_CORE_DATAPATH__abc_16259_n8301), .B(AES_CORE_DATAPATH__abc_16259_n8303), .Y(AES_CORE_DATAPATH__abc_16259_n8304) );
  AND2X2 AND2X2_2854 ( .A(AES_CORE_DATAPATH__abc_16259_n6602), .B(AES_CORE_DATAPATH__abc_16259_n8305), .Y(AES_CORE_DATAPATH__abc_16259_n8306) );
  AND2X2 AND2X2_2855 ( .A(AES_CORE_DATAPATH__abc_16259_n8306), .B(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n8307) );
  AND2X2 AND2X2_2856 ( .A(AES_CORE_DATAPATH__abc_16259_n8308), .B(AES_CORE_DATAPATH__abc_16259_n8309), .Y(AES_CORE_DATAPATH__0col_3__31_0__10_) );
  AND2X2 AND2X2_2857 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf7), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_75_), .Y(AES_CORE_DATAPATH__abc_16259_n8313) );
  AND2X2 AND2X2_2858 ( .A(AES_CORE_DATAPATH__abc_16259_n8312), .B(AES_CORE_DATAPATH__abc_16259_n8314), .Y(AES_CORE_DATAPATH__abc_16259_n8315) );
  AND2X2 AND2X2_2859 ( .A(AES_CORE_DATAPATH__abc_16259_n6657), .B(AES_CORE_DATAPATH__abc_16259_n8316), .Y(AES_CORE_DATAPATH__abc_16259_n8317) );
  AND2X2 AND2X2_286 ( .A(AES_CORE_DATAPATH__abc_16259_n2821), .B(AES_CORE_DATAPATH__abc_16259_n2824_1), .Y(AES_CORE_DATAPATH__abc_16259_n2825) );
  AND2X2 AND2X2_2860 ( .A(AES_CORE_DATAPATH__abc_16259_n8317), .B(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n8318) );
  AND2X2 AND2X2_2861 ( .A(AES_CORE_DATAPATH__abc_16259_n8319), .B(AES_CORE_DATAPATH__abc_16259_n8320), .Y(AES_CORE_DATAPATH__0col_3__31_0__11_) );
  AND2X2 AND2X2_2862 ( .A(AES_CORE_DATAPATH__abc_16259_n8219_bF_buf4), .B(AES_CORE_DATAPATH_col_3__12_), .Y(AES_CORE_DATAPATH__abc_16259_n8322) );
  AND2X2 AND2X2_2863 ( .A(AES_CORE_DATAPATH__abc_16259_n8323), .B(AES_CORE_DATAPATH__abc_16259_n8324), .Y(AES_CORE_DATAPATH__abc_16259_n8325) );
  AND2X2 AND2X2_2864 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n8325), .Y(AES_CORE_DATAPATH__abc_16259_n8326) );
  AND2X2 AND2X2_2865 ( .A(AES_CORE_DATAPATH__abc_16259_n8327), .B(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n8328) );
  AND2X2 AND2X2_2866 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf4), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_77_), .Y(AES_CORE_DATAPATH__abc_16259_n8332) );
  AND2X2 AND2X2_2867 ( .A(AES_CORE_DATAPATH__abc_16259_n8331), .B(AES_CORE_DATAPATH__abc_16259_n8333), .Y(AES_CORE_DATAPATH__abc_16259_n8334) );
  AND2X2 AND2X2_2868 ( .A(AES_CORE_DATAPATH__abc_16259_n6760), .B(AES_CORE_DATAPATH__abc_16259_n8335), .Y(AES_CORE_DATAPATH__abc_16259_n8336) );
  AND2X2 AND2X2_2869 ( .A(AES_CORE_DATAPATH__abc_16259_n8336), .B(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n8337) );
  AND2X2 AND2X2_287 ( .A(AES_CORE_DATAPATH__abc_16259_n2815), .B(AES_CORE_DATAPATH__abc_16259_n2825), .Y(AES_CORE_DATAPATH__abc_16259_n2826) );
  AND2X2 AND2X2_2870 ( .A(AES_CORE_DATAPATH__abc_16259_n8338), .B(AES_CORE_DATAPATH__abc_16259_n8339), .Y(AES_CORE_DATAPATH__0col_3__31_0__13_) );
  AND2X2 AND2X2_2871 ( .A(AES_CORE_DATAPATH__abc_16259_n8219_bF_buf3), .B(AES_CORE_DATAPATH_col_3__14_), .Y(AES_CORE_DATAPATH__abc_16259_n8341) );
  AND2X2 AND2X2_2872 ( .A(AES_CORE_DATAPATH__abc_16259_n8342), .B(AES_CORE_DATAPATH__abc_16259_n8343), .Y(AES_CORE_DATAPATH__abc_16259_n8344) );
  AND2X2 AND2X2_2873 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf9), .B(AES_CORE_DATAPATH__abc_16259_n8344), .Y(AES_CORE_DATAPATH__abc_16259_n8345) );
  AND2X2 AND2X2_2874 ( .A(AES_CORE_DATAPATH__abc_16259_n8346), .B(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n8347) );
  AND2X2 AND2X2_2875 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf1), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_79_), .Y(AES_CORE_DATAPATH__abc_16259_n8351) );
  AND2X2 AND2X2_2876 ( .A(AES_CORE_DATAPATH__abc_16259_n8350), .B(AES_CORE_DATAPATH__abc_16259_n8352), .Y(AES_CORE_DATAPATH__abc_16259_n8353) );
  AND2X2 AND2X2_2877 ( .A(AES_CORE_DATAPATH__abc_16259_n6863), .B(AES_CORE_DATAPATH__abc_16259_n8354), .Y(AES_CORE_DATAPATH__abc_16259_n8355) );
  AND2X2 AND2X2_2878 ( .A(AES_CORE_DATAPATH__abc_16259_n8355), .B(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n8356) );
  AND2X2 AND2X2_2879 ( .A(AES_CORE_DATAPATH__abc_16259_n8357), .B(AES_CORE_DATAPATH__abc_16259_n8358), .Y(AES_CORE_DATAPATH__0col_3__31_0__15_) );
  AND2X2 AND2X2_288 ( .A(AES_CORE_DATAPATH__abc_16259_n2815), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__0_), .Y(AES_CORE_DATAPATH__abc_16259_n2827) );
  AND2X2 AND2X2_2880 ( .A(AES_CORE_DATAPATH__abc_16259_n8219_bF_buf2), .B(AES_CORE_DATAPATH_col_3__16_), .Y(AES_CORE_DATAPATH__abc_16259_n8360) );
  AND2X2 AND2X2_2881 ( .A(AES_CORE_DATAPATH__abc_16259_n8361), .B(AES_CORE_DATAPATH__abc_16259_n8362), .Y(AES_CORE_DATAPATH__abc_16259_n8363) );
  AND2X2 AND2X2_2882 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf8), .B(AES_CORE_DATAPATH__abc_16259_n8363), .Y(AES_CORE_DATAPATH__abc_16259_n8364) );
  AND2X2 AND2X2_2883 ( .A(AES_CORE_DATAPATH__abc_16259_n8365), .B(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n8366) );
  AND2X2 AND2X2_2884 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf13), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_113_), .Y(AES_CORE_DATAPATH__abc_16259_n8370) );
  AND2X2 AND2X2_2885 ( .A(AES_CORE_DATAPATH__abc_16259_n8369), .B(AES_CORE_DATAPATH__abc_16259_n8371), .Y(AES_CORE_DATAPATH__abc_16259_n8372) );
  AND2X2 AND2X2_2886 ( .A(AES_CORE_DATAPATH__abc_16259_n6966), .B(AES_CORE_DATAPATH__abc_16259_n8373), .Y(AES_CORE_DATAPATH__abc_16259_n8374) );
  AND2X2 AND2X2_2887 ( .A(AES_CORE_DATAPATH__abc_16259_n8374), .B(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n8375) );
  AND2X2 AND2X2_2888 ( .A(AES_CORE_DATAPATH__abc_16259_n8376), .B(AES_CORE_DATAPATH__abc_16259_n8377), .Y(AES_CORE_DATAPATH__0col_3__31_0__17_) );
  AND2X2 AND2X2_2889 ( .A(AES_CORE_DATAPATH__abc_16259_n8219_bF_buf1), .B(AES_CORE_DATAPATH_col_3__18_), .Y(AES_CORE_DATAPATH__abc_16259_n8379) );
  AND2X2 AND2X2_289 ( .A(AES_CORE_DATAPATH__abc_16259_n2825), .B(AES_CORE_DATAPATH__abc_16259_n2829_1), .Y(AES_CORE_DATAPATH__abc_16259_n2830_1) );
  AND2X2 AND2X2_2890 ( .A(AES_CORE_DATAPATH__abc_16259_n8380), .B(AES_CORE_DATAPATH__abc_16259_n8381), .Y(AES_CORE_DATAPATH__abc_16259_n8382) );
  AND2X2 AND2X2_2891 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf7), .B(AES_CORE_DATAPATH__abc_16259_n8382), .Y(AES_CORE_DATAPATH__abc_16259_n8383) );
  AND2X2 AND2X2_2892 ( .A(AES_CORE_DATAPATH__abc_16259_n8384), .B(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n8385) );
  AND2X2 AND2X2_2893 ( .A(AES_CORE_DATAPATH__abc_16259_n8219_bF_buf0), .B(AES_CORE_DATAPATH_col_3__19_), .Y(AES_CORE_DATAPATH__abc_16259_n8387) );
  AND2X2 AND2X2_2894 ( .A(AES_CORE_DATAPATH__abc_16259_n8388), .B(AES_CORE_DATAPATH__abc_16259_n8389), .Y(AES_CORE_DATAPATH__abc_16259_n8390) );
  AND2X2 AND2X2_2895 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf6), .B(AES_CORE_DATAPATH__abc_16259_n8390), .Y(AES_CORE_DATAPATH__abc_16259_n8391) );
  AND2X2 AND2X2_2896 ( .A(AES_CORE_DATAPATH__abc_16259_n8392), .B(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n8393) );
  AND2X2 AND2X2_2897 ( .A(AES_CORE_DATAPATH__abc_16259_n8219_bF_buf4), .B(AES_CORE_DATAPATH_col_3__20_), .Y(AES_CORE_DATAPATH__abc_16259_n8395) );
  AND2X2 AND2X2_2898 ( .A(AES_CORE_DATAPATH__abc_16259_n8396), .B(AES_CORE_DATAPATH__abc_16259_n8397), .Y(AES_CORE_DATAPATH__abc_16259_n8398) );
  AND2X2 AND2X2_2899 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf5), .B(AES_CORE_DATAPATH__abc_16259_n8398), .Y(AES_CORE_DATAPATH__abc_16259_n8399) );
  AND2X2 AND2X2_29 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n85), .B(AES_CORE_CONTROL_UNIT__abc_15841_n114_1), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n115) );
  AND2X2 AND2X2_290 ( .A(AES_CORE_DATAPATH__abc_16259_n2830_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__0_), .Y(AES_CORE_DATAPATH__abc_16259_n2831) );
  AND2X2 AND2X2_2900 ( .A(AES_CORE_DATAPATH__abc_16259_n8400), .B(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n8401) );
  AND2X2 AND2X2_2901 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf8), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_117_), .Y(AES_CORE_DATAPATH__abc_16259_n8405) );
  AND2X2 AND2X2_2902 ( .A(AES_CORE_DATAPATH__abc_16259_n8404), .B(AES_CORE_DATAPATH__abc_16259_n8406), .Y(AES_CORE_DATAPATH__abc_16259_n8407) );
  AND2X2 AND2X2_2903 ( .A(AES_CORE_DATAPATH__abc_16259_n7167), .B(AES_CORE_DATAPATH__abc_16259_n8408), .Y(AES_CORE_DATAPATH__abc_16259_n8409) );
  AND2X2 AND2X2_2904 ( .A(AES_CORE_DATAPATH__abc_16259_n8409), .B(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n8410) );
  AND2X2 AND2X2_2905 ( .A(AES_CORE_DATAPATH__abc_16259_n8411), .B(AES_CORE_DATAPATH__abc_16259_n8412), .Y(AES_CORE_DATAPATH__0col_3__31_0__21_) );
  AND2X2 AND2X2_2906 ( .A(AES_CORE_DATAPATH__abc_16259_n8219_bF_buf3), .B(AES_CORE_DATAPATH_col_3__22_), .Y(AES_CORE_DATAPATH__abc_16259_n8414) );
  AND2X2 AND2X2_2907 ( .A(AES_CORE_DATAPATH__abc_16259_n8415), .B(AES_CORE_DATAPATH__abc_16259_n8416), .Y(AES_CORE_DATAPATH__abc_16259_n8417) );
  AND2X2 AND2X2_2908 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n8417), .Y(AES_CORE_DATAPATH__abc_16259_n8418) );
  AND2X2 AND2X2_2909 ( .A(AES_CORE_DATAPATH__abc_16259_n8419), .B(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n8420) );
  AND2X2 AND2X2_291 ( .A(AES_CORE_DATAPATH__abc_16259_n2804_1_bF_buf2), .B(AES_CORE_DATAPATH_key_out_sel_pp1_0_), .Y(AES_CORE_DATAPATH__abc_16259_n2832) );
  AND2X2 AND2X2_2910 ( .A(AES_CORE_DATAPATH__abc_16259_n8219_bF_buf2), .B(AES_CORE_DATAPATH_col_3__23_), .Y(AES_CORE_DATAPATH__abc_16259_n8422) );
  AND2X2 AND2X2_2911 ( .A(AES_CORE_DATAPATH__abc_16259_n8423), .B(AES_CORE_DATAPATH__abc_16259_n8424), .Y(AES_CORE_DATAPATH__abc_16259_n8425) );
  AND2X2 AND2X2_2912 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n8425), .Y(AES_CORE_DATAPATH__abc_16259_n8426) );
  AND2X2 AND2X2_2913 ( .A(AES_CORE_DATAPATH__abc_16259_n8427), .B(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n8428) );
  AND2X2 AND2X2_2914 ( .A(AES_CORE_DATAPATH__abc_16259_n8219_bF_buf1), .B(AES_CORE_DATAPATH_col_3__24_), .Y(AES_CORE_DATAPATH__abc_16259_n8430) );
  AND2X2 AND2X2_2915 ( .A(AES_CORE_DATAPATH__abc_16259_n8431), .B(AES_CORE_DATAPATH__abc_16259_n8432), .Y(AES_CORE_DATAPATH__abc_16259_n8433) );
  AND2X2 AND2X2_2916 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n8433), .Y(AES_CORE_DATAPATH__abc_16259_n8434) );
  AND2X2 AND2X2_2917 ( .A(AES_CORE_DATAPATH__abc_16259_n8435), .B(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n8436) );
  AND2X2 AND2X2_2918 ( .A(AES_CORE_DATAPATH__abc_16259_n8219_bF_buf0), .B(AES_CORE_DATAPATH_col_3__25_), .Y(AES_CORE_DATAPATH__abc_16259_n8438) );
  AND2X2 AND2X2_2919 ( .A(AES_CORE_DATAPATH__abc_16259_n8439), .B(AES_CORE_DATAPATH__abc_16259_n8440), .Y(AES_CORE_DATAPATH__abc_16259_n8441) );
  AND2X2 AND2X2_292 ( .A(AES_CORE_DATAPATH__abc_16259_n2807_bF_buf3), .B(AES_CORE_DATAPATH_key_out_sel_pp2_0_), .Y(AES_CORE_DATAPATH__abc_16259_n2833_1) );
  AND2X2 AND2X2_2920 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n8441), .Y(AES_CORE_DATAPATH__abc_16259_n8442) );
  AND2X2 AND2X2_2921 ( .A(AES_CORE_DATAPATH__abc_16259_n8443), .B(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n8444) );
  AND2X2 AND2X2_2922 ( .A(AES_CORE_DATAPATH__abc_16259_n8219_bF_buf4), .B(AES_CORE_DATAPATH_col_3__26_), .Y(AES_CORE_DATAPATH__abc_16259_n8446) );
  AND2X2 AND2X2_2923 ( .A(AES_CORE_DATAPATH__abc_16259_n8447), .B(AES_CORE_DATAPATH__abc_16259_n8448), .Y(AES_CORE_DATAPATH__abc_16259_n8449) );
  AND2X2 AND2X2_2924 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n8449), .Y(AES_CORE_DATAPATH__abc_16259_n8450) );
  AND2X2 AND2X2_2925 ( .A(AES_CORE_DATAPATH__abc_16259_n8451), .B(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n8452) );
  AND2X2 AND2X2_2926 ( .A(AES_CORE_DATAPATH__abc_16259_n8219_bF_buf3), .B(AES_CORE_DATAPATH_col_3__27_), .Y(AES_CORE_DATAPATH__abc_16259_n8454) );
  AND2X2 AND2X2_2927 ( .A(AES_CORE_DATAPATH__abc_16259_n8455), .B(AES_CORE_DATAPATH__abc_16259_n8456), .Y(AES_CORE_DATAPATH__abc_16259_n8457) );
  AND2X2 AND2X2_2928 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf9), .B(AES_CORE_DATAPATH__abc_16259_n8457), .Y(AES_CORE_DATAPATH__abc_16259_n8458) );
  AND2X2 AND2X2_2929 ( .A(AES_CORE_DATAPATH__abc_16259_n8459), .B(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n8460) );
  AND2X2 AND2X2_293 ( .A(AES_CORE_DATAPATH__abc_16259_n2834), .B(AES_CORE_DATAPATH__abc_16259_n2806_1), .Y(AES_CORE_DATAPATH__abc_16259_n2835_1) );
  AND2X2 AND2X2_2930 ( .A(AES_CORE_DATAPATH__abc_16259_n8219_bF_buf2), .B(AES_CORE_DATAPATH_col_3__28_), .Y(AES_CORE_DATAPATH__abc_16259_n8462) );
  AND2X2 AND2X2_2931 ( .A(AES_CORE_DATAPATH__abc_16259_n8463), .B(AES_CORE_DATAPATH__abc_16259_n8464), .Y(AES_CORE_DATAPATH__abc_16259_n8465) );
  AND2X2 AND2X2_2932 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf8), .B(AES_CORE_DATAPATH__abc_16259_n8465), .Y(AES_CORE_DATAPATH__abc_16259_n8466) );
  AND2X2 AND2X2_2933 ( .A(AES_CORE_DATAPATH__abc_16259_n8467), .B(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n8468) );
  AND2X2 AND2X2_2934 ( .A(AES_CORE_DATAPATH__abc_16259_n8219_bF_buf1), .B(AES_CORE_DATAPATH_col_3__29_), .Y(AES_CORE_DATAPATH__abc_16259_n8470) );
  AND2X2 AND2X2_2935 ( .A(AES_CORE_DATAPATH__abc_16259_n8471), .B(AES_CORE_DATAPATH__abc_16259_n8472), .Y(AES_CORE_DATAPATH__abc_16259_n8473) );
  AND2X2 AND2X2_2936 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf7), .B(AES_CORE_DATAPATH__abc_16259_n8473), .Y(AES_CORE_DATAPATH__abc_16259_n8474) );
  AND2X2 AND2X2_2937 ( .A(AES_CORE_DATAPATH__abc_16259_n8475), .B(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n8476) );
  AND2X2 AND2X2_2938 ( .A(AES_CORE_DATAPATH__abc_16259_n8219_bF_buf0), .B(AES_CORE_DATAPATH_col_3__30_), .Y(AES_CORE_DATAPATH__abc_16259_n8478) );
  AND2X2 AND2X2_2939 ( .A(AES_CORE_DATAPATH__abc_16259_n8479), .B(AES_CORE_DATAPATH__abc_16259_n8480), .Y(AES_CORE_DATAPATH__abc_16259_n8481) );
  AND2X2 AND2X2_294 ( .A(AES_CORE_DATAPATH__abc_16259_n2836), .B(AES_CORE_DATAPATH__abc_16259_n2829_1), .Y(AES_CORE_DATAPATH__abc_16259_n2837_1) );
  AND2X2 AND2X2_2940 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf6), .B(AES_CORE_DATAPATH__abc_16259_n8481), .Y(AES_CORE_DATAPATH__abc_16259_n8482) );
  AND2X2 AND2X2_2941 ( .A(AES_CORE_DATAPATH__abc_16259_n8483), .B(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n8484) );
  AND2X2 AND2X2_2942 ( .A(AES_CORE_DATAPATH__abc_16259_n8219_bF_buf4), .B(AES_CORE_DATAPATH_col_3__31_), .Y(AES_CORE_DATAPATH__abc_16259_n8486) );
  AND2X2 AND2X2_2943 ( .A(AES_CORE_DATAPATH__abc_16259_n8487), .B(AES_CORE_DATAPATH__abc_16259_n8488), .Y(AES_CORE_DATAPATH__abc_16259_n8489) );
  AND2X2 AND2X2_2944 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf5), .B(AES_CORE_DATAPATH__abc_16259_n8489), .Y(AES_CORE_DATAPATH__abc_16259_n8490) );
  AND2X2 AND2X2_2945 ( .A(AES_CORE_DATAPATH__abc_16259_n8491), .B(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n8492) );
  AND2X2 AND2X2_2946 ( .A(AES_CORE_DATAPATH__abc_16259_n6595), .B(AES_CORE_DATAPATH__abc_16259_n6059_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n8494) );
  AND2X2 AND2X2_2947 ( .A(AES_CORE_DATAPATH__abc_16259_n8494), .B(AES_CORE_DATAPATH_col_en_host_3_), .Y(AES_CORE_DATAPATH__abc_16259_n8495) );
  AND2X2 AND2X2_2948 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf12), .B(AES_CORE_CONTROL_UNIT_mode_cbc_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n8496) );
  AND2X2 AND2X2_2949 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf11), .B(AES_CORE_CONTROL_UNIT_last_round_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n8497) );
  AND2X2 AND2X2_295 ( .A(AES_CORE_DATAPATH__abc_16259_n2837_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__0_), .Y(AES_CORE_DATAPATH__abc_16259_n2838) );
  AND2X2 AND2X2_2950 ( .A(AES_CORE_DATAPATH__abc_16259_n8497), .B(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_3_), .Y(AES_CORE_DATAPATH__abc_16259_n8498) );
  AND2X2 AND2X2_2951 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf6), .B(AES_CORE_DATAPATH_bkp_1_3__0_), .Y(AES_CORE_DATAPATH__abc_16259_n8501) );
  AND2X2 AND2X2_2952 ( .A(AES_CORE_DATAPATH__abc_16259_n6112), .B(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n8502) );
  AND2X2 AND2X2_2953 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf5), .B(AES_CORE_DATAPATH_bkp_1_3__1_), .Y(AES_CORE_DATAPATH__abc_16259_n8504) );
  AND2X2 AND2X2_2954 ( .A(AES_CORE_DATAPATH__abc_16259_n6161), .B(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n8505) );
  AND2X2 AND2X2_2955 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf4), .B(AES_CORE_DATAPATH_bkp_1_3__2_), .Y(AES_CORE_DATAPATH__abc_16259_n8507) );
  AND2X2 AND2X2_2956 ( .A(AES_CORE_DATAPATH__abc_16259_n6210), .B(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n8508) );
  AND2X2 AND2X2_2957 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1_3__3_), .Y(AES_CORE_DATAPATH__abc_16259_n8510) );
  AND2X2 AND2X2_2958 ( .A(AES_CORE_DATAPATH__abc_16259_n6259), .B(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n8511) );
  AND2X2 AND2X2_2959 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf2), .B(AES_CORE_DATAPATH_bkp_1_3__4_), .Y(AES_CORE_DATAPATH__abc_16259_n8513) );
  AND2X2 AND2X2_296 ( .A(AES_CORE_DATAPATH__abc_16259_n2840), .B(AES_CORE_DATAPATH__abc_16259_n2842), .Y(_auto_iopadmap_cc_313_execute_26949_0_) );
  AND2X2 AND2X2_2960 ( .A(AES_CORE_DATAPATH__abc_16259_n6308), .B(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n8514) );
  AND2X2 AND2X2_2961 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf1), .B(AES_CORE_DATAPATH_bkp_1_3__5_), .Y(AES_CORE_DATAPATH__abc_16259_n8516) );
  AND2X2 AND2X2_2962 ( .A(AES_CORE_DATAPATH__abc_16259_n6357), .B(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n8517) );
  AND2X2 AND2X2_2963 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf0), .B(AES_CORE_DATAPATH_bkp_1_3__6_), .Y(AES_CORE_DATAPATH__abc_16259_n8519) );
  AND2X2 AND2X2_2964 ( .A(AES_CORE_DATAPATH__abc_16259_n6406), .B(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n8520) );
  AND2X2 AND2X2_2965 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf6), .B(AES_CORE_DATAPATH_bkp_1_3__7_), .Y(AES_CORE_DATAPATH__abc_16259_n8522) );
  AND2X2 AND2X2_2966 ( .A(AES_CORE_DATAPATH__abc_16259_n6455), .B(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n8523) );
  AND2X2 AND2X2_2967 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf5), .B(AES_CORE_DATAPATH_bkp_1_3__8_), .Y(AES_CORE_DATAPATH__abc_16259_n8525) );
  AND2X2 AND2X2_2968 ( .A(AES_CORE_DATAPATH__abc_16259_n6504), .B(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n8526) );
  AND2X2 AND2X2_2969 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf4), .B(AES_CORE_DATAPATH_bkp_1_3__9_), .Y(AES_CORE_DATAPATH__abc_16259_n8528) );
  AND2X2 AND2X2_297 ( .A(AES_CORE_DATAPATH__abc_16259_n2457_1), .B(AES_CORE_DATAPATH_rk_sel_pp2_1_), .Y(AES_CORE_DATAPATH__abc_16259_n2844) );
  AND2X2 AND2X2_2970 ( .A(AES_CORE_DATAPATH__abc_16259_n6553), .B(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n8529) );
  AND2X2 AND2X2_2971 ( .A(AES_CORE_DATAPATH__abc_16259_n6610), .B(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n8531) );
  AND2X2 AND2X2_2972 ( .A(AES_CORE_DATAPATH__abc_16259_n8532), .B(AES_CORE_DATAPATH__abc_16259_n8533), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__10_) );
  AND2X2 AND2X2_2973 ( .A(AES_CORE_DATAPATH__abc_16259_n6664), .B(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n8535) );
  AND2X2 AND2X2_2974 ( .A(AES_CORE_DATAPATH__abc_16259_n8536), .B(AES_CORE_DATAPATH__abc_16259_n8537), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__11_) );
  AND2X2 AND2X2_2975 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1_3__12_), .Y(AES_CORE_DATAPATH__abc_16259_n8539) );
  AND2X2 AND2X2_2976 ( .A(AES_CORE_DATAPATH__abc_16259_n6715), .B(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n8540) );
  AND2X2 AND2X2_2977 ( .A(AES_CORE_DATAPATH__abc_16259_n6767), .B(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n8542) );
  AND2X2 AND2X2_2978 ( .A(AES_CORE_DATAPATH__abc_16259_n8543), .B(AES_CORE_DATAPATH__abc_16259_n8544), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__13_) );
  AND2X2 AND2X2_2979 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf2), .B(AES_CORE_DATAPATH_bkp_1_3__14_), .Y(AES_CORE_DATAPATH__abc_16259_n8546) );
  AND2X2 AND2X2_298 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk_bF_buf0), .B(AES_CORE_CONTROL_UNIT_rk_sel_1_), .Y(AES_CORE_DATAPATH__abc_16259_n2845) );
  AND2X2 AND2X2_2980 ( .A(AES_CORE_DATAPATH__abc_16259_n6818), .B(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n8547) );
  AND2X2 AND2X2_2981 ( .A(AES_CORE_DATAPATH__abc_16259_n6870), .B(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n8549) );
  AND2X2 AND2X2_2982 ( .A(AES_CORE_DATAPATH__abc_16259_n8550), .B(AES_CORE_DATAPATH__abc_16259_n8551), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__15_) );
  AND2X2 AND2X2_2983 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf1), .B(AES_CORE_DATAPATH_bkp_1_3__16_), .Y(AES_CORE_DATAPATH__abc_16259_n8553) );
  AND2X2 AND2X2_2984 ( .A(AES_CORE_DATAPATH__abc_16259_n6921), .B(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n8554) );
  AND2X2 AND2X2_2985 ( .A(AES_CORE_DATAPATH__abc_16259_n6973), .B(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n8556) );
  AND2X2 AND2X2_2986 ( .A(AES_CORE_DATAPATH__abc_16259_n8557), .B(AES_CORE_DATAPATH__abc_16259_n8558), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__17_) );
  AND2X2 AND2X2_2987 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf0), .B(AES_CORE_DATAPATH_bkp_1_3__18_), .Y(AES_CORE_DATAPATH__abc_16259_n8560) );
  AND2X2 AND2X2_2988 ( .A(AES_CORE_DATAPATH__abc_16259_n7024), .B(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n8561) );
  AND2X2 AND2X2_2989 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf6), .B(AES_CORE_DATAPATH_bkp_1_3__19_), .Y(AES_CORE_DATAPATH__abc_16259_n8563) );
  AND2X2 AND2X2_299 ( .A(AES_CORE_DATAPATH__abc_16259_n2457_1), .B(AES_CORE_DATAPATH_rk_sel_pp2_0_), .Y(AES_CORE_DATAPATH__abc_16259_n2848) );
  AND2X2 AND2X2_2990 ( .A(AES_CORE_DATAPATH__abc_16259_n7073), .B(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n8564) );
  AND2X2 AND2X2_2991 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf5), .B(AES_CORE_DATAPATH_bkp_1_3__20_), .Y(AES_CORE_DATAPATH__abc_16259_n8566) );
  AND2X2 AND2X2_2992 ( .A(AES_CORE_DATAPATH__abc_16259_n7122), .B(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n8567) );
  AND2X2 AND2X2_2993 ( .A(AES_CORE_DATAPATH__abc_16259_n7174), .B(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n8569) );
  AND2X2 AND2X2_2994 ( .A(AES_CORE_DATAPATH__abc_16259_n8570), .B(AES_CORE_DATAPATH__abc_16259_n8571), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__21_) );
  AND2X2 AND2X2_2995 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf4), .B(AES_CORE_DATAPATH_bkp_1_3__22_), .Y(AES_CORE_DATAPATH__abc_16259_n8573) );
  AND2X2 AND2X2_2996 ( .A(AES_CORE_DATAPATH__abc_16259_n7225), .B(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n8574) );
  AND2X2 AND2X2_2997 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1_3__23_), .Y(AES_CORE_DATAPATH__abc_16259_n8576) );
  AND2X2 AND2X2_2998 ( .A(AES_CORE_DATAPATH__abc_16259_n7274), .B(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n8577) );
  AND2X2 AND2X2_2999 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf2), .B(AES_CORE_DATAPATH_bkp_1_3__24_), .Y(AES_CORE_DATAPATH__abc_16259_n8579) );
  AND2X2 AND2X2_3 ( .A(\addr[0] ), .B(write_en), .Y(_abc_15830_n15) );
  AND2X2 AND2X2_30 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf13), .B(AES_CORE_CONTROL_UNIT_state_14_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n117_1) );
  AND2X2 AND2X2_300 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk_bF_buf3), .B(AES_CORE_CONTROL_UNIT_rk_sel_0_), .Y(AES_CORE_DATAPATH__abc_16259_n2849) );
  AND2X2 AND2X2_3000 ( .A(AES_CORE_DATAPATH__abc_16259_n7323), .B(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n8580) );
  AND2X2 AND2X2_3001 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf1), .B(AES_CORE_DATAPATH_bkp_1_3__25_), .Y(AES_CORE_DATAPATH__abc_16259_n8582) );
  AND2X2 AND2X2_3002 ( .A(AES_CORE_DATAPATH__abc_16259_n7372), .B(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n8583) );
  AND2X2 AND2X2_3003 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf0), .B(AES_CORE_DATAPATH_bkp_1_3__26_), .Y(AES_CORE_DATAPATH__abc_16259_n8585) );
  AND2X2 AND2X2_3004 ( .A(AES_CORE_DATAPATH__abc_16259_n7421), .B(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n8586) );
  AND2X2 AND2X2_3005 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf6), .B(AES_CORE_DATAPATH_bkp_1_3__27_), .Y(AES_CORE_DATAPATH__abc_16259_n8588) );
  AND2X2 AND2X2_3006 ( .A(AES_CORE_DATAPATH__abc_16259_n7470), .B(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n8589) );
  AND2X2 AND2X2_3007 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf5), .B(AES_CORE_DATAPATH_bkp_1_3__28_), .Y(AES_CORE_DATAPATH__abc_16259_n8591) );
  AND2X2 AND2X2_3008 ( .A(AES_CORE_DATAPATH__abc_16259_n7519), .B(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n8592) );
  AND2X2 AND2X2_3009 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf4), .B(AES_CORE_DATAPATH_bkp_1_3__29_), .Y(AES_CORE_DATAPATH__abc_16259_n8594) );
  AND2X2 AND2X2_301 ( .A(AES_CORE_DATAPATH__abc_16259_n2847), .B(AES_CORE_DATAPATH__abc_16259_n2851_1), .Y(AES_CORE_DATAPATH__abc_16259_n2852) );
  AND2X2 AND2X2_3010 ( .A(AES_CORE_DATAPATH__abc_16259_n7568), .B(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n8595) );
  AND2X2 AND2X2_3011 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1_3__30_), .Y(AES_CORE_DATAPATH__abc_16259_n8597) );
  AND2X2 AND2X2_3012 ( .A(AES_CORE_DATAPATH__abc_16259_n7617), .B(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n8598) );
  AND2X2 AND2X2_3013 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf2), .B(AES_CORE_DATAPATH_bkp_1_3__31_), .Y(AES_CORE_DATAPATH__abc_16259_n8600) );
  AND2X2 AND2X2_3014 ( .A(AES_CORE_DATAPATH__abc_16259_n7666), .B(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n8601) );
  AND2X2 AND2X2_3015 ( .A(AES_CORE_DATAPATH__abc_16259_n8605), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n8606) );
  AND2X2 AND2X2_3016 ( .A(AES_CORE_DATAPATH__abc_16259_n8604), .B(AES_CORE_DATAPATH__abc_16259_n8606), .Y(AES_CORE_DATAPATH__abc_16259_n8607) );
  AND2X2 AND2X2_3017 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf0), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_0_), .Y(AES_CORE_DATAPATH__abc_16259_n8608) );
  AND2X2 AND2X2_3018 ( .A(AES_CORE_DATAPATH__abc_16259_n8610), .B(AES_CORE_DATAPATH__abc_16259_n8611), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__0_) );
  AND2X2 AND2X2_3019 ( .A(AES_CORE_DATAPATH__abc_16259_n8614), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n8615) );
  AND2X2 AND2X2_302 ( .A(AES_CORE_DATAPATH__abc_16259_n2851_1), .B(AES_CORE_DATAPATH__abc_16259_n2846), .Y(AES_CORE_DATAPATH__abc_16259_n2855) );
  AND2X2 AND2X2_3020 ( .A(AES_CORE_DATAPATH__abc_16259_n8613), .B(AES_CORE_DATAPATH__abc_16259_n8615), .Y(AES_CORE_DATAPATH__abc_16259_n8616) );
  AND2X2 AND2X2_3021 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf5), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_1_), .Y(AES_CORE_DATAPATH__abc_16259_n8617) );
  AND2X2 AND2X2_3022 ( .A(AES_CORE_DATAPATH__abc_16259_n8619), .B(AES_CORE_DATAPATH__abc_16259_n8620), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__1_) );
  AND2X2 AND2X2_3023 ( .A(AES_CORE_DATAPATH__abc_16259_n8623), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n8624) );
  AND2X2 AND2X2_3024 ( .A(AES_CORE_DATAPATH__abc_16259_n8622), .B(AES_CORE_DATAPATH__abc_16259_n8624), .Y(AES_CORE_DATAPATH__abc_16259_n8625) );
  AND2X2 AND2X2_3025 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf4), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_2_), .Y(AES_CORE_DATAPATH__abc_16259_n8626) );
  AND2X2 AND2X2_3026 ( .A(AES_CORE_DATAPATH__abc_16259_n8628), .B(AES_CORE_DATAPATH__abc_16259_n8629), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__2_) );
  AND2X2 AND2X2_3027 ( .A(AES_CORE_DATAPATH__abc_16259_n8632), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n8633) );
  AND2X2 AND2X2_3028 ( .A(AES_CORE_DATAPATH__abc_16259_n8631), .B(AES_CORE_DATAPATH__abc_16259_n8633), .Y(AES_CORE_DATAPATH__abc_16259_n8634) );
  AND2X2 AND2X2_3029 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf3), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_3_), .Y(AES_CORE_DATAPATH__abc_16259_n8635) );
  AND2X2 AND2X2_303 ( .A(AES_CORE_DATAPATH__abc_16259_n2855_bF_buf4), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_0_), .Y(AES_CORE_DATAPATH__abc_16259_n2856) );
  AND2X2 AND2X2_3030 ( .A(AES_CORE_DATAPATH__abc_16259_n8637), .B(AES_CORE_DATAPATH__abc_16259_n8638), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__3_) );
  AND2X2 AND2X2_3031 ( .A(AES_CORE_DATAPATH__abc_16259_n8641), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n8642) );
  AND2X2 AND2X2_3032 ( .A(AES_CORE_DATAPATH__abc_16259_n8640), .B(AES_CORE_DATAPATH__abc_16259_n8642), .Y(AES_CORE_DATAPATH__abc_16259_n8643) );
  AND2X2 AND2X2_3033 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf2), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_4_), .Y(AES_CORE_DATAPATH__abc_16259_n8644) );
  AND2X2 AND2X2_3034 ( .A(AES_CORE_DATAPATH__abc_16259_n8646), .B(AES_CORE_DATAPATH__abc_16259_n8647), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__4_) );
  AND2X2 AND2X2_3035 ( .A(AES_CORE_DATAPATH__abc_16259_n8650), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n8651) );
  AND2X2 AND2X2_3036 ( .A(AES_CORE_DATAPATH__abc_16259_n8649), .B(AES_CORE_DATAPATH__abc_16259_n8651), .Y(AES_CORE_DATAPATH__abc_16259_n8652) );
  AND2X2 AND2X2_3037 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf1), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_5_), .Y(AES_CORE_DATAPATH__abc_16259_n8653) );
  AND2X2 AND2X2_3038 ( .A(AES_CORE_DATAPATH__abc_16259_n8655), .B(AES_CORE_DATAPATH__abc_16259_n8656), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__5_) );
  AND2X2 AND2X2_3039 ( .A(AES_CORE_DATAPATH__abc_16259_n8659), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n8660) );
  AND2X2 AND2X2_304 ( .A(AES_CORE_DATAPATH__abc_16259_n2847), .B(AES_CORE_DATAPATH__abc_16259_n2850), .Y(AES_CORE_DATAPATH__abc_16259_n2857) );
  AND2X2 AND2X2_3040 ( .A(AES_CORE_DATAPATH__abc_16259_n8658), .B(AES_CORE_DATAPATH__abc_16259_n8660), .Y(AES_CORE_DATAPATH__abc_16259_n8661) );
  AND2X2 AND2X2_3041 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf0), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_6_), .Y(AES_CORE_DATAPATH__abc_16259_n8662) );
  AND2X2 AND2X2_3042 ( .A(AES_CORE_DATAPATH__abc_16259_n8664), .B(AES_CORE_DATAPATH__abc_16259_n8665), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__6_) );
  AND2X2 AND2X2_3043 ( .A(AES_CORE_DATAPATH__abc_16259_n8668), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf10), .Y(AES_CORE_DATAPATH__abc_16259_n8669) );
  AND2X2 AND2X2_3044 ( .A(AES_CORE_DATAPATH__abc_16259_n8667), .B(AES_CORE_DATAPATH__abc_16259_n8669), .Y(AES_CORE_DATAPATH__abc_16259_n8670) );
  AND2X2 AND2X2_3045 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf5), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_7_), .Y(AES_CORE_DATAPATH__abc_16259_n8671) );
  AND2X2 AND2X2_3046 ( .A(AES_CORE_DATAPATH__abc_16259_n8673), .B(AES_CORE_DATAPATH__abc_16259_n8674), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__7_) );
  AND2X2 AND2X2_3047 ( .A(AES_CORE_DATAPATH__abc_16259_n8677), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf9), .Y(AES_CORE_DATAPATH__abc_16259_n8678) );
  AND2X2 AND2X2_3048 ( .A(AES_CORE_DATAPATH__abc_16259_n8676), .B(AES_CORE_DATAPATH__abc_16259_n8678), .Y(AES_CORE_DATAPATH__abc_16259_n8679) );
  AND2X2 AND2X2_3049 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf4), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_8_), .Y(AES_CORE_DATAPATH__abc_16259_n8680) );
  AND2X2 AND2X2_305 ( .A(AES_CORE_DATAPATH__abc_16259_n2857_bF_buf4), .B(AES_CORE_DATAPATH_MIX_COL_col_0__0_), .Y(AES_CORE_DATAPATH__abc_16259_n2858_1) );
  AND2X2 AND2X2_3050 ( .A(AES_CORE_DATAPATH__abc_16259_n8682), .B(AES_CORE_DATAPATH__abc_16259_n8683), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__8_) );
  AND2X2 AND2X2_3051 ( .A(AES_CORE_DATAPATH__abc_16259_n8686), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf8), .Y(AES_CORE_DATAPATH__abc_16259_n8687) );
  AND2X2 AND2X2_3052 ( .A(AES_CORE_DATAPATH__abc_16259_n8685), .B(AES_CORE_DATAPATH__abc_16259_n8687), .Y(AES_CORE_DATAPATH__abc_16259_n8688) );
  AND2X2 AND2X2_3053 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf3), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_9_), .Y(AES_CORE_DATAPATH__abc_16259_n8689) );
  AND2X2 AND2X2_3054 ( .A(AES_CORE_DATAPATH__abc_16259_n8691), .B(AES_CORE_DATAPATH__abc_16259_n8692), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__9_) );
  AND2X2 AND2X2_3055 ( .A(AES_CORE_DATAPATH__abc_16259_n6610), .B(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf11), .Y(AES_CORE_DATAPATH__abc_16259_n8694) );
  AND2X2 AND2X2_3056 ( .A(AES_CORE_DATAPATH__abc_16259_n8696), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n8697) );
  AND2X2 AND2X2_3057 ( .A(AES_CORE_DATAPATH__abc_16259_n8695), .B(AES_CORE_DATAPATH__abc_16259_n8697), .Y(AES_CORE_DATAPATH__abc_16259_n8698) );
  AND2X2 AND2X2_3058 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf2), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_10_), .Y(AES_CORE_DATAPATH__abc_16259_n8699) );
  AND2X2 AND2X2_3059 ( .A(AES_CORE_DATAPATH__abc_16259_n8701), .B(AES_CORE_DATAPATH__abc_16259_n8702), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__10_) );
  AND2X2 AND2X2_306 ( .A(AES_CORE_DATAPATH__abc_16259_n2854), .B(AES_CORE_DATAPATH__abc_16259_n2860), .Y(AES_CORE_DATAPATH__abc_16259_n2861) );
  AND2X2 AND2X2_3060 ( .A(AES_CORE_DATAPATH__abc_16259_n6664), .B(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf9), .Y(AES_CORE_DATAPATH__abc_16259_n8704) );
  AND2X2 AND2X2_3061 ( .A(AES_CORE_DATAPATH__abc_16259_n8706), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n8707) );
  AND2X2 AND2X2_3062 ( .A(AES_CORE_DATAPATH__abc_16259_n8705), .B(AES_CORE_DATAPATH__abc_16259_n8707), .Y(AES_CORE_DATAPATH__abc_16259_n8708) );
  AND2X2 AND2X2_3063 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf1), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_11_), .Y(AES_CORE_DATAPATH__abc_16259_n8709) );
  AND2X2 AND2X2_3064 ( .A(AES_CORE_DATAPATH__abc_16259_n8711), .B(AES_CORE_DATAPATH__abc_16259_n8712), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__11_) );
  AND2X2 AND2X2_3065 ( .A(AES_CORE_DATAPATH__abc_16259_n8715), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n8716) );
  AND2X2 AND2X2_3066 ( .A(AES_CORE_DATAPATH__abc_16259_n8714), .B(AES_CORE_DATAPATH__abc_16259_n8716), .Y(AES_CORE_DATAPATH__abc_16259_n8717) );
  AND2X2 AND2X2_3067 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf0), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_12_), .Y(AES_CORE_DATAPATH__abc_16259_n8718) );
  AND2X2 AND2X2_3068 ( .A(AES_CORE_DATAPATH__abc_16259_n8720), .B(AES_CORE_DATAPATH__abc_16259_n8721), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__12_) );
  AND2X2 AND2X2_3069 ( .A(AES_CORE_DATAPATH__abc_16259_n6767), .B(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n8723) );
  AND2X2 AND2X2_307 ( .A(_auto_iopadmap_cc_313_execute_26949_0_), .B(AES_CORE_DATAPATH__abc_16259_n2861), .Y(AES_CORE_DATAPATH__abc_16259_n2865) );
  AND2X2 AND2X2_3070 ( .A(AES_CORE_DATAPATH__abc_16259_n8725), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n8726) );
  AND2X2 AND2X2_3071 ( .A(AES_CORE_DATAPATH__abc_16259_n8724), .B(AES_CORE_DATAPATH__abc_16259_n8726), .Y(AES_CORE_DATAPATH__abc_16259_n8727) );
  AND2X2 AND2X2_3072 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf5), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_13_), .Y(AES_CORE_DATAPATH__abc_16259_n8728) );
  AND2X2 AND2X2_3073 ( .A(AES_CORE_DATAPATH__abc_16259_n8730), .B(AES_CORE_DATAPATH__abc_16259_n8731), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__13_) );
  AND2X2 AND2X2_3074 ( .A(AES_CORE_DATAPATH__abc_16259_n8734), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n8735) );
  AND2X2 AND2X2_3075 ( .A(AES_CORE_DATAPATH__abc_16259_n8733), .B(AES_CORE_DATAPATH__abc_16259_n8735), .Y(AES_CORE_DATAPATH__abc_16259_n8736) );
  AND2X2 AND2X2_3076 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf4), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_14_), .Y(AES_CORE_DATAPATH__abc_16259_n8737) );
  AND2X2 AND2X2_3077 ( .A(AES_CORE_DATAPATH__abc_16259_n8739), .B(AES_CORE_DATAPATH__abc_16259_n8740), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__14_) );
  AND2X2 AND2X2_3078 ( .A(AES_CORE_DATAPATH__abc_16259_n6870), .B(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n8742) );
  AND2X2 AND2X2_3079 ( .A(AES_CORE_DATAPATH__abc_16259_n8744), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n8745) );
  AND2X2 AND2X2_308 ( .A(AES_CORE_DATAPATH__abc_16259_n2867), .B(AES_CORE_DATAPATH__abc_16259_n2801_1), .Y(AES_CORE_DATAPATH__abc_16259_n2868_1) );
  AND2X2 AND2X2_3080 ( .A(AES_CORE_DATAPATH__abc_16259_n8743), .B(AES_CORE_DATAPATH__abc_16259_n8745), .Y(AES_CORE_DATAPATH__abc_16259_n8746) );
  AND2X2 AND2X2_3081 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf3), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_15_), .Y(AES_CORE_DATAPATH__abc_16259_n8747) );
  AND2X2 AND2X2_3082 ( .A(AES_CORE_DATAPATH__abc_16259_n8749), .B(AES_CORE_DATAPATH__abc_16259_n8750), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__15_) );
  AND2X2 AND2X2_3083 ( .A(AES_CORE_DATAPATH__abc_16259_n8753), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n8754) );
  AND2X2 AND2X2_3084 ( .A(AES_CORE_DATAPATH__abc_16259_n8752), .B(AES_CORE_DATAPATH__abc_16259_n8754), .Y(AES_CORE_DATAPATH__abc_16259_n8755) );
  AND2X2 AND2X2_3085 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf2), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_16_), .Y(AES_CORE_DATAPATH__abc_16259_n8756) );
  AND2X2 AND2X2_3086 ( .A(AES_CORE_DATAPATH__abc_16259_n8758), .B(AES_CORE_DATAPATH__abc_16259_n8759), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__16_) );
  AND2X2 AND2X2_3087 ( .A(AES_CORE_DATAPATH__abc_16259_n6973), .B(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n8761) );
  AND2X2 AND2X2_3088 ( .A(AES_CORE_DATAPATH__abc_16259_n8763), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n8764) );
  AND2X2 AND2X2_3089 ( .A(AES_CORE_DATAPATH__abc_16259_n8762), .B(AES_CORE_DATAPATH__abc_16259_n8764), .Y(AES_CORE_DATAPATH__abc_16259_n8765) );
  AND2X2 AND2X2_309 ( .A(AES_CORE_DATAPATH__abc_16259_n2868_1), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n2869) );
  AND2X2 AND2X2_3090 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf1), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_17_), .Y(AES_CORE_DATAPATH__abc_16259_n8766) );
  AND2X2 AND2X2_3091 ( .A(AES_CORE_DATAPATH__abc_16259_n8768), .B(AES_CORE_DATAPATH__abc_16259_n8769), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__17_) );
  AND2X2 AND2X2_3092 ( .A(AES_CORE_DATAPATH__abc_16259_n8772), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf10), .Y(AES_CORE_DATAPATH__abc_16259_n8773) );
  AND2X2 AND2X2_3093 ( .A(AES_CORE_DATAPATH__abc_16259_n8771), .B(AES_CORE_DATAPATH__abc_16259_n8773), .Y(AES_CORE_DATAPATH__abc_16259_n8774) );
  AND2X2 AND2X2_3094 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf0), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_18_), .Y(AES_CORE_DATAPATH__abc_16259_n8775) );
  AND2X2 AND2X2_3095 ( .A(AES_CORE_DATAPATH__abc_16259_n8777), .B(AES_CORE_DATAPATH__abc_16259_n8778), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__18_) );
  AND2X2 AND2X2_3096 ( .A(AES_CORE_DATAPATH__abc_16259_n8781), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf9), .Y(AES_CORE_DATAPATH__abc_16259_n8782) );
  AND2X2 AND2X2_3097 ( .A(AES_CORE_DATAPATH__abc_16259_n8780), .B(AES_CORE_DATAPATH__abc_16259_n8782), .Y(AES_CORE_DATAPATH__abc_16259_n8783) );
  AND2X2 AND2X2_3098 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf5), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_19_), .Y(AES_CORE_DATAPATH__abc_16259_n8784) );
  AND2X2 AND2X2_3099 ( .A(AES_CORE_DATAPATH__abc_16259_n8786), .B(AES_CORE_DATAPATH__abc_16259_n8787), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__19_) );
  AND2X2 AND2X2_31 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n106_1), .B(AES_CORE_CONTROL_UNIT_state_9_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n118) );
  AND2X2 AND2X2_310 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf11), .B(AES_CORE_DATAPATH_col_3__0_), .Y(AES_CORE_DATAPATH__abc_16259_n2870) );
  AND2X2 AND2X2_3100 ( .A(AES_CORE_DATAPATH__abc_16259_n8790), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf8), .Y(AES_CORE_DATAPATH__abc_16259_n8791) );
  AND2X2 AND2X2_3101 ( .A(AES_CORE_DATAPATH__abc_16259_n8789), .B(AES_CORE_DATAPATH__abc_16259_n8791), .Y(AES_CORE_DATAPATH__abc_16259_n8792) );
  AND2X2 AND2X2_3102 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf4), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_20_), .Y(AES_CORE_DATAPATH__abc_16259_n8793) );
  AND2X2 AND2X2_3103 ( .A(AES_CORE_DATAPATH__abc_16259_n8795), .B(AES_CORE_DATAPATH__abc_16259_n8796), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__20_) );
  AND2X2 AND2X2_3104 ( .A(AES_CORE_DATAPATH__abc_16259_n7174), .B(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n8798) );
  AND2X2 AND2X2_3105 ( .A(AES_CORE_DATAPATH__abc_16259_n8800), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n8801) );
  AND2X2 AND2X2_3106 ( .A(AES_CORE_DATAPATH__abc_16259_n8799), .B(AES_CORE_DATAPATH__abc_16259_n8801), .Y(AES_CORE_DATAPATH__abc_16259_n8802) );
  AND2X2 AND2X2_3107 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf3), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_21_), .Y(AES_CORE_DATAPATH__abc_16259_n8803) );
  AND2X2 AND2X2_3108 ( .A(AES_CORE_DATAPATH__abc_16259_n8805), .B(AES_CORE_DATAPATH__abc_16259_n8806), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__21_) );
  AND2X2 AND2X2_3109 ( .A(AES_CORE_DATAPATH__abc_16259_n8809), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n8810) );
  AND2X2 AND2X2_311 ( .A(AES_CORE_DATAPATH__abc_16259_n2873), .B(AES_CORE_DATAPATH__abc_16259_n2875), .Y(AES_CORE_DATAPATH__abc_16259_n2876) );
  AND2X2 AND2X2_3110 ( .A(AES_CORE_DATAPATH__abc_16259_n8808), .B(AES_CORE_DATAPATH__abc_16259_n8810), .Y(AES_CORE_DATAPATH__abc_16259_n8811) );
  AND2X2 AND2X2_3111 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf2), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_22_), .Y(AES_CORE_DATAPATH__abc_16259_n8812) );
  AND2X2 AND2X2_3112 ( .A(AES_CORE_DATAPATH__abc_16259_n8814), .B(AES_CORE_DATAPATH__abc_16259_n8815), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__22_) );
  AND2X2 AND2X2_3113 ( .A(AES_CORE_DATAPATH__abc_16259_n8818), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n8819) );
  AND2X2 AND2X2_3114 ( .A(AES_CORE_DATAPATH__abc_16259_n8817), .B(AES_CORE_DATAPATH__abc_16259_n8819), .Y(AES_CORE_DATAPATH__abc_16259_n8820) );
  AND2X2 AND2X2_3115 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf1), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_23_), .Y(AES_CORE_DATAPATH__abc_16259_n8821) );
  AND2X2 AND2X2_3116 ( .A(AES_CORE_DATAPATH__abc_16259_n8823), .B(AES_CORE_DATAPATH__abc_16259_n8824), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__23_) );
  AND2X2 AND2X2_3117 ( .A(AES_CORE_DATAPATH__abc_16259_n8827), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n8828) );
  AND2X2 AND2X2_3118 ( .A(AES_CORE_DATAPATH__abc_16259_n8826), .B(AES_CORE_DATAPATH__abc_16259_n8828), .Y(AES_CORE_DATAPATH__abc_16259_n8829) );
  AND2X2 AND2X2_3119 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf0), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_24_), .Y(AES_CORE_DATAPATH__abc_16259_n8830) );
  AND2X2 AND2X2_312 ( .A(AES_CORE_DATAPATH__abc_16259_n2782_bF_buf3), .B(AES_CORE_DATAPATH_col_3__1_), .Y(AES_CORE_DATAPATH__abc_16259_n2877) );
  AND2X2 AND2X2_3120 ( .A(AES_CORE_DATAPATH__abc_16259_n8832), .B(AES_CORE_DATAPATH__abc_16259_n8833), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__24_) );
  AND2X2 AND2X2_3121 ( .A(AES_CORE_DATAPATH__abc_16259_n8836), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n8837) );
  AND2X2 AND2X2_3122 ( .A(AES_CORE_DATAPATH__abc_16259_n8835), .B(AES_CORE_DATAPATH__abc_16259_n8837), .Y(AES_CORE_DATAPATH__abc_16259_n8838) );
  AND2X2 AND2X2_3123 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf5), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_25_), .Y(AES_CORE_DATAPATH__abc_16259_n8839) );
  AND2X2 AND2X2_3124 ( .A(AES_CORE_DATAPATH__abc_16259_n8841), .B(AES_CORE_DATAPATH__abc_16259_n8842), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__25_) );
  AND2X2 AND2X2_3125 ( .A(AES_CORE_DATAPATH__abc_16259_n8845), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n8846) );
  AND2X2 AND2X2_3126 ( .A(AES_CORE_DATAPATH__abc_16259_n8844), .B(AES_CORE_DATAPATH__abc_16259_n8846), .Y(AES_CORE_DATAPATH__abc_16259_n8847) );
  AND2X2 AND2X2_3127 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf4), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_26_), .Y(AES_CORE_DATAPATH__abc_16259_n8848) );
  AND2X2 AND2X2_3128 ( .A(AES_CORE_DATAPATH__abc_16259_n8850), .B(AES_CORE_DATAPATH__abc_16259_n8851), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__26_) );
  AND2X2 AND2X2_3129 ( .A(AES_CORE_DATAPATH__abc_16259_n8854), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n8855) );
  AND2X2 AND2X2_313 ( .A(AES_CORE_DATAPATH__abc_16259_n2786_bF_buf3), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_65_), .Y(AES_CORE_DATAPATH__abc_16259_n2878) );
  AND2X2 AND2X2_3130 ( .A(AES_CORE_DATAPATH__abc_16259_n8853), .B(AES_CORE_DATAPATH__abc_16259_n8855), .Y(AES_CORE_DATAPATH__abc_16259_n8856) );
  AND2X2 AND2X2_3131 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf3), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_27_), .Y(AES_CORE_DATAPATH__abc_16259_n8857) );
  AND2X2 AND2X2_3132 ( .A(AES_CORE_DATAPATH__abc_16259_n8859), .B(AES_CORE_DATAPATH__abc_16259_n8860), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__27_) );
  AND2X2 AND2X2_3133 ( .A(AES_CORE_DATAPATH__abc_16259_n8863), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n8864) );
  AND2X2 AND2X2_3134 ( .A(AES_CORE_DATAPATH__abc_16259_n8862), .B(AES_CORE_DATAPATH__abc_16259_n8864), .Y(AES_CORE_DATAPATH__abc_16259_n8865) );
  AND2X2 AND2X2_3135 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf2), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_28_), .Y(AES_CORE_DATAPATH__abc_16259_n8866) );
  AND2X2 AND2X2_3136 ( .A(AES_CORE_DATAPATH__abc_16259_n8868), .B(AES_CORE_DATAPATH__abc_16259_n8869), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__28_) );
  AND2X2 AND2X2_3137 ( .A(AES_CORE_DATAPATH__abc_16259_n8872), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf10), .Y(AES_CORE_DATAPATH__abc_16259_n8873) );
  AND2X2 AND2X2_3138 ( .A(AES_CORE_DATAPATH__abc_16259_n8871), .B(AES_CORE_DATAPATH__abc_16259_n8873), .Y(AES_CORE_DATAPATH__abc_16259_n8874) );
  AND2X2 AND2X2_3139 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf1), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_29_), .Y(AES_CORE_DATAPATH__abc_16259_n8875) );
  AND2X2 AND2X2_314 ( .A(AES_CORE_DATAPATH__abc_16259_n2789_bF_buf3), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_33_), .Y(AES_CORE_DATAPATH__abc_16259_n2879) );
  AND2X2 AND2X2_3140 ( .A(AES_CORE_DATAPATH__abc_16259_n8877), .B(AES_CORE_DATAPATH__abc_16259_n8878), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__29_) );
  AND2X2 AND2X2_3141 ( .A(AES_CORE_DATAPATH__abc_16259_n8881), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf9), .Y(AES_CORE_DATAPATH__abc_16259_n8882) );
  AND2X2 AND2X2_3142 ( .A(AES_CORE_DATAPATH__abc_16259_n8880), .B(AES_CORE_DATAPATH__abc_16259_n8882), .Y(AES_CORE_DATAPATH__abc_16259_n8883) );
  AND2X2 AND2X2_3143 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf0), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_30_), .Y(AES_CORE_DATAPATH__abc_16259_n8884) );
  AND2X2 AND2X2_3144 ( .A(AES_CORE_DATAPATH__abc_16259_n8886), .B(AES_CORE_DATAPATH__abc_16259_n8887), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__30_) );
  AND2X2 AND2X2_3145 ( .A(AES_CORE_DATAPATH__abc_16259_n8890), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf8), .Y(AES_CORE_DATAPATH__abc_16259_n8891) );
  AND2X2 AND2X2_3146 ( .A(AES_CORE_DATAPATH__abc_16259_n8889), .B(AES_CORE_DATAPATH__abc_16259_n8891), .Y(AES_CORE_DATAPATH__abc_16259_n8892) );
  AND2X2 AND2X2_3147 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf5), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_31_), .Y(AES_CORE_DATAPATH__abc_16259_n8893) );
  AND2X2 AND2X2_3148 ( .A(AES_CORE_DATAPATH__abc_16259_n8895), .B(AES_CORE_DATAPATH__abc_16259_n8896), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__31_) );
  AND2X2 AND2X2_3149 ( .A(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf7), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .Y(AES_CORE_DATAPATH__abc_16259_n8900) );
  AND2X2 AND2X2_315 ( .A(AES_CORE_DATAPATH__abc_16259_n2882_1), .B(AES_CORE_DATAPATH__abc_16259_n2876), .Y(AES_CORE_DATAPATH__abc_16259_n2883) );
  AND2X2 AND2X2_3150 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf4), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .Y(AES_CORE_DATAPATH__abc_16259_n8905) );
  AND2X2 AND2X2_3151 ( .A(AES_CORE_DATAPATH__abc_16259_n8905_bF_buf4), .B(AES_CORE_DATAPATH_iv_3__0_), .Y(AES_CORE_DATAPATH__abc_16259_n8906) );
  AND2X2 AND2X2_3152 ( .A(AES_CORE_DATAPATH__abc_16259_n8907), .B(AES_CORE_DATAPATH__abc_16259_n8904), .Y(AES_CORE_DATAPATH__abc_16259_n8908) );
  AND2X2 AND2X2_3153 ( .A(AES_CORE_DATAPATH__abc_16259_n8909), .B(AES_CORE_DATAPATH__abc_16259_n8903), .Y(AES_CORE_DATAPATH__0iv_3__31_0__0_) );
  AND2X2 AND2X2_3154 ( .A(AES_CORE_DATAPATH_iv_3__0_), .B(AES_CORE_DATAPATH_iv_3__1_), .Y(AES_CORE_DATAPATH__abc_16259_n8912) );
  AND2X2 AND2X2_3155 ( .A(AES_CORE_DATAPATH__abc_16259_n8912), .B(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n8913) );
  AND2X2 AND2X2_3156 ( .A(AES_CORE_DATAPATH__abc_16259_n8913), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .Y(AES_CORE_DATAPATH__abc_16259_n8914) );
  AND2X2 AND2X2_3157 ( .A(AES_CORE_DATAPATH__abc_16259_n8915), .B(AES_CORE_DATAPATH__abc_16259_n8911), .Y(AES_CORE_DATAPATH__abc_16259_n8916) );
  AND2X2 AND2X2_3158 ( .A(AES_CORE_DATAPATH_iv_3__0_), .B(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n8919) );
  AND2X2 AND2X2_3159 ( .A(AES_CORE_DATAPATH__abc_16259_n8920), .B(AES_CORE_DATAPATH__abc_16259_n8898_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n8921) );
  AND2X2 AND2X2_316 ( .A(AES_CORE_DATAPATH__abc_16259_n2837_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__1_), .Y(AES_CORE_DATAPATH__abc_16259_n2885) );
  AND2X2 AND2X2_3160 ( .A(AES_CORE_DATAPATH__abc_16259_n8917), .B(AES_CORE_DATAPATH__abc_16259_n8922), .Y(AES_CORE_DATAPATH__0iv_3__31_0__1_) );
  AND2X2 AND2X2_3161 ( .A(AES_CORE_DATAPATH__abc_16259_n8924), .B(AES_CORE_DATAPATH__abc_16259_n8898_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n8925) );
  AND2X2 AND2X2_3162 ( .A(AES_CORE_DATAPATH__abc_16259_n8913), .B(AES_CORE_DATAPATH_iv_3__2_), .Y(AES_CORE_DATAPATH__abc_16259_n8928) );
  AND2X2 AND2X2_3163 ( .A(AES_CORE_DATAPATH__abc_16259_n8928), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .Y(AES_CORE_DATAPATH__abc_16259_n8929) );
  AND2X2 AND2X2_3164 ( .A(AES_CORE_DATAPATH__abc_16259_n8930), .B(AES_CORE_DATAPATH__abc_16259_n8927), .Y(AES_CORE_DATAPATH__abc_16259_n8931) );
  AND2X2 AND2X2_3165 ( .A(AES_CORE_DATAPATH__abc_16259_n8932), .B(AES_CORE_DATAPATH__abc_16259_n8926), .Y(AES_CORE_DATAPATH__0iv_3__31_0__2_) );
  AND2X2 AND2X2_3166 ( .A(AES_CORE_DATAPATH__abc_16259_n8934), .B(AES_CORE_DATAPATH__abc_16259_n8898_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n8935) );
  AND2X2 AND2X2_3167 ( .A(AES_CORE_DATAPATH_iv_3__2_), .B(AES_CORE_DATAPATH_iv_3__3_), .Y(AES_CORE_DATAPATH__abc_16259_n8938) );
  AND2X2 AND2X2_3168 ( .A(AES_CORE_DATAPATH__abc_16259_n8912), .B(AES_CORE_DATAPATH__abc_16259_n8938), .Y(AES_CORE_DATAPATH__abc_16259_n8939) );
  AND2X2 AND2X2_3169 ( .A(AES_CORE_DATAPATH__abc_16259_n8939), .B(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n8940) );
  AND2X2 AND2X2_317 ( .A(AES_CORE_DATAPATH__abc_16259_n2815), .B(AES_CORE_DATAPATH__abc_16259_n2836), .Y(AES_CORE_DATAPATH__abc_16259_n2887_1) );
  AND2X2 AND2X2_3170 ( .A(AES_CORE_DATAPATH__abc_16259_n8940), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .Y(AES_CORE_DATAPATH__abc_16259_n8941) );
  AND2X2 AND2X2_3171 ( .A(AES_CORE_DATAPATH__abc_16259_n8942), .B(AES_CORE_DATAPATH__abc_16259_n8937), .Y(AES_CORE_DATAPATH__abc_16259_n8943) );
  AND2X2 AND2X2_3172 ( .A(AES_CORE_DATAPATH__abc_16259_n8944), .B(AES_CORE_DATAPATH__abc_16259_n8936), .Y(AES_CORE_DATAPATH__0iv_3__31_0__3_) );
  AND2X2 AND2X2_3173 ( .A(AES_CORE_DATAPATH__abc_16259_n8946), .B(AES_CORE_DATAPATH__abc_16259_n8898_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n8947) );
  AND2X2 AND2X2_3174 ( .A(AES_CORE_DATAPATH__abc_16259_n8940), .B(AES_CORE_DATAPATH_iv_3__4_), .Y(AES_CORE_DATAPATH__abc_16259_n8950) );
  AND2X2 AND2X2_3175 ( .A(AES_CORE_DATAPATH__abc_16259_n8950), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .Y(AES_CORE_DATAPATH__abc_16259_n8951) );
  AND2X2 AND2X2_3176 ( .A(AES_CORE_DATAPATH__abc_16259_n8952), .B(AES_CORE_DATAPATH__abc_16259_n8949), .Y(AES_CORE_DATAPATH__abc_16259_n8953) );
  AND2X2 AND2X2_3177 ( .A(AES_CORE_DATAPATH__abc_16259_n8954), .B(AES_CORE_DATAPATH__abc_16259_n8948), .Y(AES_CORE_DATAPATH__0iv_3__31_0__4_) );
  AND2X2 AND2X2_3178 ( .A(AES_CORE_DATAPATH__abc_16259_n8918_bF_buf0), .B(\bus_in[5] ), .Y(AES_CORE_DATAPATH__abc_16259_n8956) );
  AND2X2 AND2X2_3179 ( .A(AES_CORE_DATAPATH__abc_16259_n8957), .B(AES_CORE_DATAPATH__abc_16259_n8898_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n8958) );
  AND2X2 AND2X2_318 ( .A(AES_CORE_DATAPATH__abc_16259_n2887_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__1_), .Y(AES_CORE_DATAPATH__abc_16259_n2888_1) );
  AND2X2 AND2X2_3180 ( .A(AES_CORE_DATAPATH_iv_3__4_), .B(AES_CORE_DATAPATH_iv_3__5_), .Y(AES_CORE_DATAPATH__abc_16259_n8960) );
  AND2X2 AND2X2_3181 ( .A(AES_CORE_DATAPATH__abc_16259_n8940), .B(AES_CORE_DATAPATH__abc_16259_n8960), .Y(AES_CORE_DATAPATH__abc_16259_n8961) );
  AND2X2 AND2X2_3182 ( .A(AES_CORE_DATAPATH__abc_16259_n8962), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .Y(AES_CORE_DATAPATH__abc_16259_n8963) );
  AND2X2 AND2X2_3183 ( .A(AES_CORE_DATAPATH__abc_16259_n8959), .B(AES_CORE_DATAPATH__abc_16259_n8965), .Y(AES_CORE_DATAPATH__0iv_3__31_0__5_) );
  AND2X2 AND2X2_3184 ( .A(AES_CORE_DATAPATH__abc_16259_n8899_bF_buf2), .B(AES_CORE_DATAPATH_iv_3__6_), .Y(AES_CORE_DATAPATH__abc_16259_n8967) );
  AND2X2 AND2X2_3185 ( .A(AES_CORE_DATAPATH__abc_16259_n8898_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n8968), .Y(AES_CORE_DATAPATH__abc_16259_n8969) );
  AND2X2 AND2X2_3186 ( .A(AES_CORE_DATAPATH__abc_16259_n8962), .B(AES_CORE_DATAPATH_iv_3__6_), .Y(AES_CORE_DATAPATH__abc_16259_n8970) );
  AND2X2 AND2X2_3187 ( .A(AES_CORE_DATAPATH__abc_16259_n8961), .B(AES_CORE_DATAPATH__abc_16259_n8971), .Y(AES_CORE_DATAPATH__abc_16259_n8972) );
  AND2X2 AND2X2_3188 ( .A(AES_CORE_DATAPATH__abc_16259_n8974), .B(AES_CORE_DATAPATH__abc_16259_n8969), .Y(AES_CORE_DATAPATH__abc_16259_n8975) );
  AND2X2 AND2X2_3189 ( .A(AES_CORE_DATAPATH__abc_16259_n8918_bF_buf3), .B(\bus_in[7] ), .Y(AES_CORE_DATAPATH__abc_16259_n8977) );
  AND2X2 AND2X2_319 ( .A(AES_CORE_DATAPATH__abc_16259_n2830_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__1_), .Y(AES_CORE_DATAPATH__abc_16259_n2889) );
  AND2X2 AND2X2_3190 ( .A(AES_CORE_DATAPATH__abc_16259_n8960), .B(AES_CORE_DATAPATH_iv_3__6_), .Y(AES_CORE_DATAPATH__abc_16259_n8978) );
  AND2X2 AND2X2_3191 ( .A(AES_CORE_DATAPATH__abc_16259_n8939), .B(AES_CORE_DATAPATH__abc_16259_n8978), .Y(AES_CORE_DATAPATH__abc_16259_n8979) );
  AND2X2 AND2X2_3192 ( .A(AES_CORE_DATAPATH__abc_16259_n8979), .B(AES_CORE_DATAPATH_iv_3__7_), .Y(AES_CORE_DATAPATH__abc_16259_n8980) );
  AND2X2 AND2X2_3193 ( .A(AES_CORE_DATAPATH__abc_16259_n8981), .B(AES_CORE_DATAPATH__abc_16259_n8905_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n8982) );
  AND2X2 AND2X2_3194 ( .A(AES_CORE_DATAPATH__abc_16259_n8982), .B(AES_CORE_DATAPATH__abc_16259_n8979), .Y(AES_CORE_DATAPATH__abc_16259_n8983) );
  AND2X2 AND2X2_3195 ( .A(AES_CORE_DATAPATH__abc_16259_n8984), .B(AES_CORE_DATAPATH__abc_16259_n8898_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n8985) );
  AND2X2 AND2X2_3196 ( .A(AES_CORE_DATAPATH__abc_16259_n8986), .B(AES_CORE_DATAPATH_iv_3__7_), .Y(AES_CORE_DATAPATH__abc_16259_n8987) );
  AND2X2 AND2X2_3197 ( .A(AES_CORE_DATAPATH__abc_16259_n8918_bF_buf2), .B(\bus_in[8] ), .Y(AES_CORE_DATAPATH__abc_16259_n8989) );
  AND2X2 AND2X2_3198 ( .A(AES_CORE_DATAPATH__abc_16259_n8980), .B(AES_CORE_DATAPATH_iv_3__8_), .Y(AES_CORE_DATAPATH__abc_16259_n8990) );
  AND2X2 AND2X2_3199 ( .A(AES_CORE_DATAPATH__abc_16259_n8991), .B(AES_CORE_DATAPATH__abc_16259_n8905_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n8992) );
  AND2X2 AND2X2_32 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n119), .B(AES_CORE_CONTROL_UNIT__abc_15841_n84_1), .Y(AES_CORE_CONTROL_UNIT__abc_10818_n24) );
  AND2X2 AND2X2_320 ( .A(AES_CORE_DATAPATH__abc_16259_n2891_1), .B(AES_CORE_DATAPATH__abc_16259_n2892), .Y(_auto_iopadmap_cc_313_execute_26949_1_) );
  AND2X2 AND2X2_3200 ( .A(AES_CORE_DATAPATH__abc_16259_n8992), .B(AES_CORE_DATAPATH__abc_16259_n8980), .Y(AES_CORE_DATAPATH__abc_16259_n8993) );
  AND2X2 AND2X2_3201 ( .A(AES_CORE_DATAPATH__abc_16259_n8994), .B(AES_CORE_DATAPATH__abc_16259_n8898_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n8995) );
  AND2X2 AND2X2_3202 ( .A(AES_CORE_DATAPATH__abc_16259_n8996), .B(AES_CORE_DATAPATH_iv_3__8_), .Y(AES_CORE_DATAPATH__abc_16259_n8997) );
  AND2X2 AND2X2_3203 ( .A(AES_CORE_DATAPATH__abc_16259_n8900_bF_buf2), .B(AES_CORE_DATAPATH_iv_3__9_), .Y(AES_CORE_DATAPATH__abc_16259_n9001) );
  AND2X2 AND2X2_3204 ( .A(AES_CORE_DATAPATH_iv_3__8_), .B(AES_CORE_DATAPATH_iv_3__9_), .Y(AES_CORE_DATAPATH__abc_16259_n9002) );
  AND2X2 AND2X2_3205 ( .A(AES_CORE_DATAPATH__abc_16259_n8980), .B(AES_CORE_DATAPATH__abc_16259_n9002), .Y(AES_CORE_DATAPATH__abc_16259_n9003) );
  AND2X2 AND2X2_3206 ( .A(AES_CORE_DATAPATH__abc_16259_n9004), .B(AES_CORE_DATAPATH__abc_16259_n8905_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n9005) );
  AND2X2 AND2X2_3207 ( .A(AES_CORE_DATAPATH__abc_16259_n9006), .B(AES_CORE_DATAPATH__abc_16259_n9000), .Y(AES_CORE_DATAPATH__abc_16259_n9007) );
  AND2X2 AND2X2_3208 ( .A(AES_CORE_DATAPATH__abc_16259_n8918_bF_buf1), .B(\bus_in[9] ), .Y(AES_CORE_DATAPATH__abc_16259_n9008) );
  AND2X2 AND2X2_3209 ( .A(AES_CORE_DATAPATH__abc_16259_n9010), .B(AES_CORE_DATAPATH__abc_16259_n8999), .Y(AES_CORE_DATAPATH__0iv_3__31_0__9_) );
  AND2X2 AND2X2_321 ( .A(AES_CORE_DATAPATH__abc_16259_n2855_bF_buf3), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_1_), .Y(AES_CORE_DATAPATH__abc_16259_n2895_1) );
  AND2X2 AND2X2_3210 ( .A(AES_CORE_DATAPATH__abc_16259_n9003), .B(AES_CORE_DATAPATH_iv_3__10_), .Y(AES_CORE_DATAPATH__abc_16259_n9014) );
  AND2X2 AND2X2_3211 ( .A(AES_CORE_DATAPATH__abc_16259_n9015), .B(AES_CORE_DATAPATH__abc_16259_n9013), .Y(AES_CORE_DATAPATH__abc_16259_n9016) );
  AND2X2 AND2X2_3212 ( .A(AES_CORE_DATAPATH__abc_16259_n9016), .B(AES_CORE_DATAPATH__abc_16259_n8905_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n9017) );
  AND2X2 AND2X2_3213 ( .A(AES_CORE_DATAPATH__abc_16259_n8900_bF_buf1), .B(AES_CORE_DATAPATH_iv_3__10_), .Y(AES_CORE_DATAPATH__abc_16259_n9018) );
  AND2X2 AND2X2_3214 ( .A(AES_CORE_DATAPATH__abc_16259_n8918_bF_buf0), .B(\bus_in[10] ), .Y(AES_CORE_DATAPATH__abc_16259_n9019) );
  AND2X2 AND2X2_3215 ( .A(AES_CORE_DATAPATH__abc_16259_n9022), .B(AES_CORE_DATAPATH__abc_16259_n9012), .Y(AES_CORE_DATAPATH__0iv_3__31_0__10_) );
  AND2X2 AND2X2_3216 ( .A(AES_CORE_DATAPATH__abc_16259_n8900_bF_buf0), .B(AES_CORE_DATAPATH_iv_3__11_), .Y(AES_CORE_DATAPATH__abc_16259_n9026) );
  AND2X2 AND2X2_3217 ( .A(AES_CORE_DATAPATH__abc_16259_n9014), .B(AES_CORE_DATAPATH_iv_3__11_), .Y(AES_CORE_DATAPATH__abc_16259_n9027) );
  AND2X2 AND2X2_3218 ( .A(AES_CORE_DATAPATH__abc_16259_n9028), .B(AES_CORE_DATAPATH__abc_16259_n8905_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n9029) );
  AND2X2 AND2X2_3219 ( .A(AES_CORE_DATAPATH__abc_16259_n9030), .B(AES_CORE_DATAPATH__abc_16259_n9025), .Y(AES_CORE_DATAPATH__abc_16259_n9031) );
  AND2X2 AND2X2_322 ( .A(AES_CORE_DATAPATH__abc_16259_n2857_bF_buf3), .B(AES_CORE_DATAPATH_MIX_COL_col_0__1_), .Y(AES_CORE_DATAPATH__abc_16259_n2896) );
  AND2X2 AND2X2_3220 ( .A(AES_CORE_DATAPATH__abc_16259_n8918_bF_buf4), .B(\bus_in[11] ), .Y(AES_CORE_DATAPATH__abc_16259_n9032) );
  AND2X2 AND2X2_3221 ( .A(AES_CORE_DATAPATH__abc_16259_n9034), .B(AES_CORE_DATAPATH__abc_16259_n9024), .Y(AES_CORE_DATAPATH__0iv_3__31_0__11_) );
  AND2X2 AND2X2_3222 ( .A(AES_CORE_DATAPATH__abc_16259_n9027), .B(AES_CORE_DATAPATH_iv_3__12_), .Y(AES_CORE_DATAPATH__abc_16259_n9037) );
  AND2X2 AND2X2_3223 ( .A(AES_CORE_DATAPATH__abc_16259_n9039), .B(AES_CORE_DATAPATH__abc_16259_n8905_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n9040) );
  AND2X2 AND2X2_3224 ( .A(AES_CORE_DATAPATH__abc_16259_n9040), .B(AES_CORE_DATAPATH__abc_16259_n9038), .Y(AES_CORE_DATAPATH__abc_16259_n9041) );
  AND2X2 AND2X2_3225 ( .A(AES_CORE_DATAPATH__abc_16259_n8900_bF_buf3), .B(AES_CORE_DATAPATH_iv_3__12_), .Y(AES_CORE_DATAPATH__abc_16259_n9042) );
  AND2X2 AND2X2_3226 ( .A(AES_CORE_DATAPATH__abc_16259_n8918_bF_buf3), .B(\bus_in[12] ), .Y(AES_CORE_DATAPATH__abc_16259_n9043) );
  AND2X2 AND2X2_3227 ( .A(AES_CORE_DATAPATH__abc_16259_n9046), .B(AES_CORE_DATAPATH__abc_16259_n9036), .Y(AES_CORE_DATAPATH__0iv_3__31_0__12_) );
  AND2X2 AND2X2_3228 ( .A(AES_CORE_DATAPATH__abc_16259_n9037), .B(AES_CORE_DATAPATH_iv_3__13_), .Y(AES_CORE_DATAPATH__abc_16259_n9049) );
  AND2X2 AND2X2_3229 ( .A(AES_CORE_DATAPATH__abc_16259_n9051), .B(AES_CORE_DATAPATH__abc_16259_n8905_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n9052) );
  AND2X2 AND2X2_323 ( .A(AES_CORE_DATAPATH__abc_16259_n2894), .B(AES_CORE_DATAPATH__abc_16259_n2898), .Y(AES_CORE_DATAPATH__abc_16259_n2899) );
  AND2X2 AND2X2_3230 ( .A(AES_CORE_DATAPATH__abc_16259_n9052), .B(AES_CORE_DATAPATH__abc_16259_n9050), .Y(AES_CORE_DATAPATH__abc_16259_n9053) );
  AND2X2 AND2X2_3231 ( .A(AES_CORE_DATAPATH__abc_16259_n8900_bF_buf2), .B(AES_CORE_DATAPATH_iv_3__13_), .Y(AES_CORE_DATAPATH__abc_16259_n9054) );
  AND2X2 AND2X2_3232 ( .A(AES_CORE_DATAPATH__abc_16259_n8918_bF_buf2), .B(\bus_in[13] ), .Y(AES_CORE_DATAPATH__abc_16259_n9055) );
  AND2X2 AND2X2_3233 ( .A(AES_CORE_DATAPATH__abc_16259_n9058), .B(AES_CORE_DATAPATH__abc_16259_n9048), .Y(AES_CORE_DATAPATH__0iv_3__31_0__13_) );
  AND2X2 AND2X2_3234 ( .A(AES_CORE_DATAPATH__abc_16259_n9049), .B(AES_CORE_DATAPATH_iv_3__14_), .Y(AES_CORE_DATAPATH__abc_16259_n9061) );
  AND2X2 AND2X2_3235 ( .A(AES_CORE_DATAPATH__abc_16259_n9063), .B(AES_CORE_DATAPATH__abc_16259_n8905_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n9064) );
  AND2X2 AND2X2_3236 ( .A(AES_CORE_DATAPATH__abc_16259_n9064), .B(AES_CORE_DATAPATH__abc_16259_n9062), .Y(AES_CORE_DATAPATH__abc_16259_n9065) );
  AND2X2 AND2X2_3237 ( .A(AES_CORE_DATAPATH__abc_16259_n8900_bF_buf1), .B(AES_CORE_DATAPATH_iv_3__14_), .Y(AES_CORE_DATAPATH__abc_16259_n9066) );
  AND2X2 AND2X2_3238 ( .A(AES_CORE_DATAPATH__abc_16259_n8918_bF_buf1), .B(\bus_in[14] ), .Y(AES_CORE_DATAPATH__abc_16259_n9067) );
  AND2X2 AND2X2_3239 ( .A(AES_CORE_DATAPATH__abc_16259_n9070), .B(AES_CORE_DATAPATH__abc_16259_n9060), .Y(AES_CORE_DATAPATH__0iv_3__31_0__14_) );
  AND2X2 AND2X2_324 ( .A(_auto_iopadmap_cc_313_execute_26949_1_), .B(AES_CORE_DATAPATH__abc_16259_n2899), .Y(AES_CORE_DATAPATH__abc_16259_n2902) );
  AND2X2 AND2X2_3240 ( .A(AES_CORE_DATAPATH__abc_16259_n9061), .B(AES_CORE_DATAPATH_iv_3__15_), .Y(AES_CORE_DATAPATH__abc_16259_n9073) );
  AND2X2 AND2X2_3241 ( .A(AES_CORE_DATAPATH__abc_16259_n9075), .B(AES_CORE_DATAPATH__abc_16259_n8905_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n9076) );
  AND2X2 AND2X2_3242 ( .A(AES_CORE_DATAPATH__abc_16259_n9076), .B(AES_CORE_DATAPATH__abc_16259_n9074), .Y(AES_CORE_DATAPATH__abc_16259_n9077) );
  AND2X2 AND2X2_3243 ( .A(AES_CORE_DATAPATH__abc_16259_n8900_bF_buf0), .B(AES_CORE_DATAPATH_iv_3__15_), .Y(AES_CORE_DATAPATH__abc_16259_n9078) );
  AND2X2 AND2X2_3244 ( .A(AES_CORE_DATAPATH__abc_16259_n8918_bF_buf0), .B(\bus_in[15] ), .Y(AES_CORE_DATAPATH__abc_16259_n9079) );
  AND2X2 AND2X2_3245 ( .A(AES_CORE_DATAPATH__abc_16259_n9082), .B(AES_CORE_DATAPATH__abc_16259_n9072), .Y(AES_CORE_DATAPATH__0iv_3__31_0__15_) );
  AND2X2 AND2X2_3246 ( .A(AES_CORE_DATAPATH__abc_16259_n9073), .B(AES_CORE_DATAPATH_iv_3__16_), .Y(AES_CORE_DATAPATH__abc_16259_n9085) );
  AND2X2 AND2X2_3247 ( .A(AES_CORE_DATAPATH__abc_16259_n9087), .B(AES_CORE_DATAPATH__abc_16259_n8905_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n9088) );
  AND2X2 AND2X2_3248 ( .A(AES_CORE_DATAPATH__abc_16259_n9088), .B(AES_CORE_DATAPATH__abc_16259_n9086), .Y(AES_CORE_DATAPATH__abc_16259_n9089) );
  AND2X2 AND2X2_3249 ( .A(AES_CORE_DATAPATH__abc_16259_n8900_bF_buf3), .B(AES_CORE_DATAPATH_iv_3__16_), .Y(AES_CORE_DATAPATH__abc_16259_n9090) );
  AND2X2 AND2X2_325 ( .A(AES_CORE_DATAPATH_last_round_pp2_bF_buf2), .B(AES_CORE_DATAPATH_MIX_COL_col_0__1_), .Y(AES_CORE_DATAPATH__abc_16259_n2905) );
  AND2X2 AND2X2_3250 ( .A(AES_CORE_DATAPATH__abc_16259_n8918_bF_buf4), .B(\bus_in[16] ), .Y(AES_CORE_DATAPATH__abc_16259_n9091) );
  AND2X2 AND2X2_3251 ( .A(AES_CORE_DATAPATH__abc_16259_n9094), .B(AES_CORE_DATAPATH__abc_16259_n9084), .Y(AES_CORE_DATAPATH__0iv_3__31_0__16_) );
  AND2X2 AND2X2_3252 ( .A(AES_CORE_DATAPATH__abc_16259_n9085), .B(AES_CORE_DATAPATH_iv_3__17_), .Y(AES_CORE_DATAPATH__abc_16259_n9097) );
  AND2X2 AND2X2_3253 ( .A(AES_CORE_DATAPATH__abc_16259_n9099), .B(AES_CORE_DATAPATH__abc_16259_n8905_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n9100) );
  AND2X2 AND2X2_3254 ( .A(AES_CORE_DATAPATH__abc_16259_n9100), .B(AES_CORE_DATAPATH__abc_16259_n9098), .Y(AES_CORE_DATAPATH__abc_16259_n9101) );
  AND2X2 AND2X2_3255 ( .A(AES_CORE_DATAPATH__abc_16259_n8900_bF_buf2), .B(AES_CORE_DATAPATH_iv_3__17_), .Y(AES_CORE_DATAPATH__abc_16259_n9102) );
  AND2X2 AND2X2_3256 ( .A(AES_CORE_DATAPATH__abc_16259_n8918_bF_buf3), .B(\bus_in[17] ), .Y(AES_CORE_DATAPATH__abc_16259_n9103) );
  AND2X2 AND2X2_3257 ( .A(AES_CORE_DATAPATH__abc_16259_n9106), .B(AES_CORE_DATAPATH__abc_16259_n9096), .Y(AES_CORE_DATAPATH__0iv_3__31_0__17_) );
  AND2X2 AND2X2_3258 ( .A(AES_CORE_DATAPATH_iv_3__17_), .B(AES_CORE_DATAPATH_iv_3__18_), .Y(AES_CORE_DATAPATH__abc_16259_n9110) );
  AND2X2 AND2X2_3259 ( .A(AES_CORE_DATAPATH__abc_16259_n9085), .B(AES_CORE_DATAPATH__abc_16259_n9110), .Y(AES_CORE_DATAPATH__abc_16259_n9111) );
  AND2X2 AND2X2_326 ( .A(AES_CORE_DATAPATH__abc_16259_n2798_bF_buf3), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_1_), .Y(AES_CORE_DATAPATH__abc_16259_n2906) );
  AND2X2 AND2X2_3260 ( .A(AES_CORE_DATAPATH__abc_16259_n9112), .B(AES_CORE_DATAPATH__abc_16259_n8905_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n9113) );
  AND2X2 AND2X2_3261 ( .A(AES_CORE_DATAPATH__abc_16259_n9113), .B(AES_CORE_DATAPATH__abc_16259_n9109), .Y(AES_CORE_DATAPATH__abc_16259_n9114) );
  AND2X2 AND2X2_3262 ( .A(AES_CORE_DATAPATH__abc_16259_n8900_bF_buf1), .B(AES_CORE_DATAPATH_iv_3__18_), .Y(AES_CORE_DATAPATH__abc_16259_n9115) );
  AND2X2 AND2X2_3263 ( .A(AES_CORE_DATAPATH__abc_16259_n8918_bF_buf2), .B(\bus_in[18] ), .Y(AES_CORE_DATAPATH__abc_16259_n9116) );
  AND2X2 AND2X2_3264 ( .A(AES_CORE_DATAPATH__abc_16259_n9119), .B(AES_CORE_DATAPATH__abc_16259_n9108), .Y(AES_CORE_DATAPATH__0iv_3__31_0__18_) );
  AND2X2 AND2X2_3265 ( .A(AES_CORE_DATAPATH__abc_16259_n9111), .B(AES_CORE_DATAPATH_iv_3__19_), .Y(AES_CORE_DATAPATH__abc_16259_n9122) );
  AND2X2 AND2X2_3266 ( .A(AES_CORE_DATAPATH__abc_16259_n9124), .B(AES_CORE_DATAPATH__abc_16259_n8905_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n9125) );
  AND2X2 AND2X2_3267 ( .A(AES_CORE_DATAPATH__abc_16259_n9125), .B(AES_CORE_DATAPATH__abc_16259_n9123), .Y(AES_CORE_DATAPATH__abc_16259_n9126) );
  AND2X2 AND2X2_3268 ( .A(AES_CORE_DATAPATH__abc_16259_n8900_bF_buf0), .B(AES_CORE_DATAPATH_iv_3__19_), .Y(AES_CORE_DATAPATH__abc_16259_n9127) );
  AND2X2 AND2X2_3269 ( .A(AES_CORE_DATAPATH__abc_16259_n8918_bF_buf1), .B(\bus_in[19] ), .Y(AES_CORE_DATAPATH__abc_16259_n9128) );
  AND2X2 AND2X2_327 ( .A(AES_CORE_DATAPATH__abc_16259_n2904), .B(AES_CORE_DATAPATH__abc_16259_n2908), .Y(AES_CORE_DATAPATH__abc_16259_n2909_1) );
  AND2X2 AND2X2_3270 ( .A(AES_CORE_DATAPATH__abc_16259_n9131), .B(AES_CORE_DATAPATH__abc_16259_n9121), .Y(AES_CORE_DATAPATH__0iv_3__31_0__19_) );
  AND2X2 AND2X2_3271 ( .A(AES_CORE_DATAPATH__abc_16259_n9110), .B(AES_CORE_DATAPATH_iv_3__19_), .Y(AES_CORE_DATAPATH__abc_16259_n9134) );
  AND2X2 AND2X2_3272 ( .A(AES_CORE_DATAPATH__abc_16259_n9085), .B(AES_CORE_DATAPATH__abc_16259_n9134), .Y(AES_CORE_DATAPATH__abc_16259_n9135) );
  AND2X2 AND2X2_3273 ( .A(AES_CORE_DATAPATH__abc_16259_n9135), .B(AES_CORE_DATAPATH_iv_3__20_), .Y(AES_CORE_DATAPATH__abc_16259_n9137) );
  AND2X2 AND2X2_3274 ( .A(AES_CORE_DATAPATH__abc_16259_n9138), .B(AES_CORE_DATAPATH__abc_16259_n9136), .Y(AES_CORE_DATAPATH__abc_16259_n9139) );
  AND2X2 AND2X2_3275 ( .A(AES_CORE_DATAPATH__abc_16259_n9139), .B(AES_CORE_DATAPATH__abc_16259_n8905_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n9140) );
  AND2X2 AND2X2_3276 ( .A(AES_CORE_DATAPATH__abc_16259_n8900_bF_buf3), .B(AES_CORE_DATAPATH_iv_3__20_), .Y(AES_CORE_DATAPATH__abc_16259_n9141) );
  AND2X2 AND2X2_3277 ( .A(AES_CORE_DATAPATH__abc_16259_n8918_bF_buf0), .B(\bus_in[20] ), .Y(AES_CORE_DATAPATH__abc_16259_n9142) );
  AND2X2 AND2X2_3278 ( .A(AES_CORE_DATAPATH__abc_16259_n9145), .B(AES_CORE_DATAPATH__abc_16259_n9133), .Y(AES_CORE_DATAPATH__0iv_3__31_0__20_) );
  AND2X2 AND2X2_3279 ( .A(AES_CORE_DATAPATH__abc_16259_n9138), .B(AES_CORE_DATAPATH_iv_3__21_), .Y(AES_CORE_DATAPATH__abc_16259_n9148) );
  AND2X2 AND2X2_328 ( .A(AES_CORE_DATAPATH__abc_16259_n2909_1), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n2910) );
  AND2X2 AND2X2_3280 ( .A(AES_CORE_DATAPATH__abc_16259_n9137), .B(AES_CORE_DATAPATH__abc_16259_n9149), .Y(AES_CORE_DATAPATH__abc_16259_n9150) );
  AND2X2 AND2X2_3281 ( .A(AES_CORE_DATAPATH__abc_16259_n9151), .B(AES_CORE_DATAPATH__abc_16259_n8905_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n9152) );
  AND2X2 AND2X2_3282 ( .A(AES_CORE_DATAPATH__abc_16259_n8900_bF_buf2), .B(AES_CORE_DATAPATH_iv_3__21_), .Y(AES_CORE_DATAPATH__abc_16259_n9153) );
  AND2X2 AND2X2_3283 ( .A(AES_CORE_DATAPATH__abc_16259_n8918_bF_buf4), .B(\bus_in[21] ), .Y(AES_CORE_DATAPATH__abc_16259_n9154) );
  AND2X2 AND2X2_3284 ( .A(AES_CORE_DATAPATH__abc_16259_n9157), .B(AES_CORE_DATAPATH__abc_16259_n9147), .Y(AES_CORE_DATAPATH__0iv_3__31_0__21_) );
  AND2X2 AND2X2_3285 ( .A(AES_CORE_DATAPATH__abc_16259_n9137), .B(AES_CORE_DATAPATH_iv_3__21_), .Y(AES_CORE_DATAPATH__abc_16259_n9160) );
  AND2X2 AND2X2_3286 ( .A(AES_CORE_DATAPATH__abc_16259_n9122), .B(AES_CORE_DATAPATH_iv_3__20_), .Y(AES_CORE_DATAPATH__abc_16259_n9162) );
  AND2X2 AND2X2_3287 ( .A(AES_CORE_DATAPATH_iv_3__21_), .B(AES_CORE_DATAPATH_iv_3__22_), .Y(AES_CORE_DATAPATH__abc_16259_n9163) );
  AND2X2 AND2X2_3288 ( .A(AES_CORE_DATAPATH__abc_16259_n9162), .B(AES_CORE_DATAPATH__abc_16259_n9163), .Y(AES_CORE_DATAPATH__abc_16259_n9164) );
  AND2X2 AND2X2_3289 ( .A(AES_CORE_DATAPATH__abc_16259_n9165), .B(AES_CORE_DATAPATH__abc_16259_n8905_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n9166) );
  AND2X2 AND2X2_329 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf10), .B(AES_CORE_DATAPATH_col_3__1_), .Y(AES_CORE_DATAPATH__abc_16259_n2911_1) );
  AND2X2 AND2X2_3290 ( .A(AES_CORE_DATAPATH__abc_16259_n9166), .B(AES_CORE_DATAPATH__abc_16259_n9161), .Y(AES_CORE_DATAPATH__abc_16259_n9167) );
  AND2X2 AND2X2_3291 ( .A(AES_CORE_DATAPATH__abc_16259_n8900_bF_buf1), .B(AES_CORE_DATAPATH_iv_3__22_), .Y(AES_CORE_DATAPATH__abc_16259_n9168) );
  AND2X2 AND2X2_3292 ( .A(AES_CORE_DATAPATH__abc_16259_n8918_bF_buf3), .B(\bus_in[22] ), .Y(AES_CORE_DATAPATH__abc_16259_n9169) );
  AND2X2 AND2X2_3293 ( .A(AES_CORE_DATAPATH__abc_16259_n9172), .B(AES_CORE_DATAPATH__abc_16259_n9159), .Y(AES_CORE_DATAPATH__0iv_3__31_0__22_) );
  AND2X2 AND2X2_3294 ( .A(AES_CORE_DATAPATH__abc_16259_n9164), .B(AES_CORE_DATAPATH_iv_3__23_), .Y(AES_CORE_DATAPATH__abc_16259_n9175) );
  AND2X2 AND2X2_3295 ( .A(AES_CORE_DATAPATH__abc_16259_n9177), .B(AES_CORE_DATAPATH__abc_16259_n8905_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n9178) );
  AND2X2 AND2X2_3296 ( .A(AES_CORE_DATAPATH__abc_16259_n9178), .B(AES_CORE_DATAPATH__abc_16259_n9176), .Y(AES_CORE_DATAPATH__abc_16259_n9179) );
  AND2X2 AND2X2_3297 ( .A(AES_CORE_DATAPATH__abc_16259_n8900_bF_buf0), .B(AES_CORE_DATAPATH_iv_3__23_), .Y(AES_CORE_DATAPATH__abc_16259_n9180) );
  AND2X2 AND2X2_3298 ( .A(AES_CORE_DATAPATH__abc_16259_n8918_bF_buf2), .B(\bus_in[23] ), .Y(AES_CORE_DATAPATH__abc_16259_n9181) );
  AND2X2 AND2X2_3299 ( .A(AES_CORE_DATAPATH__abc_16259_n9184), .B(AES_CORE_DATAPATH__abc_16259_n9174), .Y(AES_CORE_DATAPATH__0iv_3__31_0__23_) );
  AND2X2 AND2X2_33 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n111), .B(AES_CORE_CONTROL_UNIT_key_gen), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n121) );
  AND2X2 AND2X2_330 ( .A(AES_CORE_DATAPATH__abc_16259_n2914), .B(AES_CORE_DATAPATH__abc_16259_n2916_1), .Y(AES_CORE_DATAPATH__abc_16259_n2917_1) );
  AND2X2 AND2X2_3300 ( .A(AES_CORE_DATAPATH__abc_16259_n9163), .B(AES_CORE_DATAPATH_iv_3__23_), .Y(AES_CORE_DATAPATH__abc_16259_n9187) );
  AND2X2 AND2X2_3301 ( .A(AES_CORE_DATAPATH__abc_16259_n9137), .B(AES_CORE_DATAPATH__abc_16259_n9187), .Y(AES_CORE_DATAPATH__abc_16259_n9188) );
  AND2X2 AND2X2_3302 ( .A(AES_CORE_DATAPATH__abc_16259_n9188), .B(AES_CORE_DATAPATH_iv_3__24_), .Y(AES_CORE_DATAPATH__abc_16259_n9190) );
  AND2X2 AND2X2_3303 ( .A(AES_CORE_DATAPATH__abc_16259_n9191), .B(AES_CORE_DATAPATH__abc_16259_n9189), .Y(AES_CORE_DATAPATH__abc_16259_n9192) );
  AND2X2 AND2X2_3304 ( .A(AES_CORE_DATAPATH__abc_16259_n9192), .B(AES_CORE_DATAPATH__abc_16259_n8905_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n9193) );
  AND2X2 AND2X2_3305 ( .A(AES_CORE_DATAPATH__abc_16259_n8900_bF_buf3), .B(AES_CORE_DATAPATH_iv_3__24_), .Y(AES_CORE_DATAPATH__abc_16259_n9194) );
  AND2X2 AND2X2_3306 ( .A(AES_CORE_DATAPATH__abc_16259_n8918_bF_buf1), .B(\bus_in[24] ), .Y(AES_CORE_DATAPATH__abc_16259_n9195) );
  AND2X2 AND2X2_3307 ( .A(AES_CORE_DATAPATH__abc_16259_n9198), .B(AES_CORE_DATAPATH__abc_16259_n9186), .Y(AES_CORE_DATAPATH__0iv_3__31_0__24_) );
  AND2X2 AND2X2_3308 ( .A(AES_CORE_DATAPATH__abc_16259_n9191), .B(AES_CORE_DATAPATH_iv_3__25_), .Y(AES_CORE_DATAPATH__abc_16259_n9201) );
  AND2X2 AND2X2_3309 ( .A(AES_CORE_DATAPATH__abc_16259_n9190), .B(AES_CORE_DATAPATH__abc_16259_n9202), .Y(AES_CORE_DATAPATH__abc_16259_n9203) );
  AND2X2 AND2X2_331 ( .A(AES_CORE_DATAPATH__abc_16259_n2782_bF_buf2), .B(AES_CORE_DATAPATH_col_3__2_), .Y(AES_CORE_DATAPATH__abc_16259_n2918) );
  AND2X2 AND2X2_3310 ( .A(AES_CORE_DATAPATH__abc_16259_n9204), .B(AES_CORE_DATAPATH__abc_16259_n8905_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n9205) );
  AND2X2 AND2X2_3311 ( .A(AES_CORE_DATAPATH__abc_16259_n8900_bF_buf2), .B(AES_CORE_DATAPATH_iv_3__25_), .Y(AES_CORE_DATAPATH__abc_16259_n9206) );
  AND2X2 AND2X2_3312 ( .A(AES_CORE_DATAPATH__abc_16259_n8918_bF_buf0), .B(\bus_in[25] ), .Y(AES_CORE_DATAPATH__abc_16259_n9207) );
  AND2X2 AND2X2_3313 ( .A(AES_CORE_DATAPATH__abc_16259_n9210), .B(AES_CORE_DATAPATH__abc_16259_n9200), .Y(AES_CORE_DATAPATH__0iv_3__31_0__25_) );
  AND2X2 AND2X2_3314 ( .A(AES_CORE_DATAPATH__abc_16259_n9190), .B(AES_CORE_DATAPATH_iv_3__25_), .Y(AES_CORE_DATAPATH__abc_16259_n9213) );
  AND2X2 AND2X2_3315 ( .A(AES_CORE_DATAPATH__abc_16259_n9213), .B(AES_CORE_DATAPATH_iv_3__26_), .Y(AES_CORE_DATAPATH__abc_16259_n9215) );
  AND2X2 AND2X2_3316 ( .A(AES_CORE_DATAPATH__abc_16259_n9216), .B(AES_CORE_DATAPATH__abc_16259_n9214), .Y(AES_CORE_DATAPATH__abc_16259_n9217) );
  AND2X2 AND2X2_3317 ( .A(AES_CORE_DATAPATH__abc_16259_n9217), .B(AES_CORE_DATAPATH__abc_16259_n8905_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n9218) );
  AND2X2 AND2X2_3318 ( .A(AES_CORE_DATAPATH__abc_16259_n8900_bF_buf1), .B(AES_CORE_DATAPATH_iv_3__26_), .Y(AES_CORE_DATAPATH__abc_16259_n9219) );
  AND2X2 AND2X2_3319 ( .A(AES_CORE_DATAPATH__abc_16259_n8918_bF_buf4), .B(\bus_in[26] ), .Y(AES_CORE_DATAPATH__abc_16259_n9220) );
  AND2X2 AND2X2_332 ( .A(AES_CORE_DATAPATH__abc_16259_n2786_bF_buf2), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_66_), .Y(AES_CORE_DATAPATH__abc_16259_n2919) );
  AND2X2 AND2X2_3320 ( .A(AES_CORE_DATAPATH__abc_16259_n9223), .B(AES_CORE_DATAPATH__abc_16259_n9212), .Y(AES_CORE_DATAPATH__0iv_3__31_0__26_) );
  AND2X2 AND2X2_3321 ( .A(AES_CORE_DATAPATH__abc_16259_n9215), .B(AES_CORE_DATAPATH_iv_3__27_), .Y(AES_CORE_DATAPATH__abc_16259_n9227) );
  AND2X2 AND2X2_3322 ( .A(AES_CORE_DATAPATH__abc_16259_n9228), .B(AES_CORE_DATAPATH__abc_16259_n9226), .Y(AES_CORE_DATAPATH__abc_16259_n9229) );
  AND2X2 AND2X2_3323 ( .A(AES_CORE_DATAPATH__abc_16259_n9229), .B(AES_CORE_DATAPATH__abc_16259_n8905_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n9230) );
  AND2X2 AND2X2_3324 ( .A(AES_CORE_DATAPATH__abc_16259_n8900_bF_buf0), .B(AES_CORE_DATAPATH_iv_3__27_), .Y(AES_CORE_DATAPATH__abc_16259_n9231) );
  AND2X2 AND2X2_3325 ( .A(AES_CORE_DATAPATH__abc_16259_n8918_bF_buf3), .B(\bus_in[27] ), .Y(AES_CORE_DATAPATH__abc_16259_n9232) );
  AND2X2 AND2X2_3326 ( .A(AES_CORE_DATAPATH__abc_16259_n9235), .B(AES_CORE_DATAPATH__abc_16259_n9225), .Y(AES_CORE_DATAPATH__0iv_3__31_0__27_) );
  AND2X2 AND2X2_3327 ( .A(AES_CORE_DATAPATH__abc_16259_n9227), .B(AES_CORE_DATAPATH_iv_3__28_), .Y(AES_CORE_DATAPATH__abc_16259_n9239) );
  AND2X2 AND2X2_3328 ( .A(AES_CORE_DATAPATH__abc_16259_n9240), .B(AES_CORE_DATAPATH__abc_16259_n9238), .Y(AES_CORE_DATAPATH__abc_16259_n9241) );
  AND2X2 AND2X2_3329 ( .A(AES_CORE_DATAPATH__abc_16259_n9241), .B(AES_CORE_DATAPATH__abc_16259_n8905_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n9242) );
  AND2X2 AND2X2_333 ( .A(AES_CORE_DATAPATH__abc_16259_n2789_bF_buf2), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_34_), .Y(AES_CORE_DATAPATH__abc_16259_n2920_1) );
  AND2X2 AND2X2_3330 ( .A(AES_CORE_DATAPATH__abc_16259_n8900_bF_buf3), .B(AES_CORE_DATAPATH_iv_3__28_), .Y(AES_CORE_DATAPATH__abc_16259_n9243) );
  AND2X2 AND2X2_3331 ( .A(AES_CORE_DATAPATH__abc_16259_n8918_bF_buf2), .B(\bus_in[28] ), .Y(AES_CORE_DATAPATH__abc_16259_n9244) );
  AND2X2 AND2X2_3332 ( .A(AES_CORE_DATAPATH__abc_16259_n9247), .B(AES_CORE_DATAPATH__abc_16259_n9237), .Y(AES_CORE_DATAPATH__0iv_3__31_0__28_) );
  AND2X2 AND2X2_3333 ( .A(AES_CORE_DATAPATH__abc_16259_n9239), .B(AES_CORE_DATAPATH_iv_3__29_), .Y(AES_CORE_DATAPATH__abc_16259_n9251) );
  AND2X2 AND2X2_3334 ( .A(AES_CORE_DATAPATH__abc_16259_n9252), .B(AES_CORE_DATAPATH__abc_16259_n9250), .Y(AES_CORE_DATAPATH__abc_16259_n9253) );
  AND2X2 AND2X2_3335 ( .A(AES_CORE_DATAPATH__abc_16259_n9253), .B(AES_CORE_DATAPATH__abc_16259_n8905_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n9254) );
  AND2X2 AND2X2_3336 ( .A(AES_CORE_DATAPATH__abc_16259_n8900_bF_buf2), .B(AES_CORE_DATAPATH_iv_3__29_), .Y(AES_CORE_DATAPATH__abc_16259_n9255) );
  AND2X2 AND2X2_3337 ( .A(AES_CORE_DATAPATH__abc_16259_n8918_bF_buf1), .B(\bus_in[29] ), .Y(AES_CORE_DATAPATH__abc_16259_n9256) );
  AND2X2 AND2X2_3338 ( .A(AES_CORE_DATAPATH__abc_16259_n9259), .B(AES_CORE_DATAPATH__abc_16259_n9249), .Y(AES_CORE_DATAPATH__0iv_3__31_0__29_) );
  AND2X2 AND2X2_3339 ( .A(AES_CORE_DATAPATH__abc_16259_n9251), .B(AES_CORE_DATAPATH_iv_3__30_), .Y(AES_CORE_DATAPATH__abc_16259_n9262) );
  AND2X2 AND2X2_334 ( .A(AES_CORE_DATAPATH__abc_16259_n2923), .B(AES_CORE_DATAPATH__abc_16259_n2917_1), .Y(AES_CORE_DATAPATH__abc_16259_n2924_1) );
  AND2X2 AND2X2_3340 ( .A(AES_CORE_DATAPATH__abc_16259_n9264), .B(AES_CORE_DATAPATH__abc_16259_n8905_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n9265) );
  AND2X2 AND2X2_3341 ( .A(AES_CORE_DATAPATH__abc_16259_n9265), .B(AES_CORE_DATAPATH__abc_16259_n9263), .Y(AES_CORE_DATAPATH__abc_16259_n9266) );
  AND2X2 AND2X2_3342 ( .A(AES_CORE_DATAPATH__abc_16259_n8900_bF_buf1), .B(AES_CORE_DATAPATH_iv_3__30_), .Y(AES_CORE_DATAPATH__abc_16259_n9267) );
  AND2X2 AND2X2_3343 ( .A(AES_CORE_DATAPATH__abc_16259_n8918_bF_buf0), .B(\bus_in[30] ), .Y(AES_CORE_DATAPATH__abc_16259_n9268) );
  AND2X2 AND2X2_3344 ( .A(AES_CORE_DATAPATH__abc_16259_n9271), .B(AES_CORE_DATAPATH__abc_16259_n9261), .Y(AES_CORE_DATAPATH__0iv_3__31_0__30_) );
  AND2X2 AND2X2_3345 ( .A(AES_CORE_DATAPATH__abc_16259_n9263), .B(AES_CORE_DATAPATH_iv_3__31_), .Y(AES_CORE_DATAPATH__abc_16259_n9274) );
  AND2X2 AND2X2_3346 ( .A(AES_CORE_DATAPATH__abc_16259_n9262), .B(AES_CORE_DATAPATH__abc_16259_n9275), .Y(AES_CORE_DATAPATH__abc_16259_n9276) );
  AND2X2 AND2X2_3347 ( .A(AES_CORE_DATAPATH__abc_16259_n9277), .B(AES_CORE_DATAPATH__abc_16259_n8905_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n9278) );
  AND2X2 AND2X2_3348 ( .A(AES_CORE_DATAPATH__abc_16259_n8900_bF_buf0), .B(AES_CORE_DATAPATH_iv_3__31_), .Y(AES_CORE_DATAPATH__abc_16259_n9279) );
  AND2X2 AND2X2_3349 ( .A(AES_CORE_DATAPATH__abc_16259_n8918_bF_buf4), .B(\bus_in[31] ), .Y(AES_CORE_DATAPATH__abc_16259_n9280) );
  AND2X2 AND2X2_335 ( .A(AES_CORE_DATAPATH__abc_16259_n2837_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__2_), .Y(AES_CORE_DATAPATH__abc_16259_n2926_1) );
  AND2X2 AND2X2_3350 ( .A(AES_CORE_DATAPATH__abc_16259_n9283), .B(AES_CORE_DATAPATH__abc_16259_n9273), .Y(AES_CORE_DATAPATH__0iv_3__31_0__31_) );
  AND2X2 AND2X2_3351 ( .A(AES_CORE_DATAPATH__abc_16259_n8494), .B(AES_CORE_DATAPATH_col_en_host_2_), .Y(AES_CORE_DATAPATH__abc_16259_n9285) );
  AND2X2 AND2X2_3352 ( .A(AES_CORE_DATAPATH__abc_16259_n8497), .B(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_2_), .Y(AES_CORE_DATAPATH__abc_16259_n9286) );
  AND2X2 AND2X2_3353 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf6), .B(AES_CORE_DATAPATH_bkp_1_2__0_), .Y(AES_CORE_DATAPATH__abc_16259_n9289) );
  AND2X2 AND2X2_3354 ( .A(AES_CORE_DATAPATH__abc_16259_n7675), .B(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n9290) );
  AND2X2 AND2X2_3355 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf5), .B(AES_CORE_DATAPATH_bkp_1_2__1_), .Y(AES_CORE_DATAPATH__abc_16259_n9292) );
  AND2X2 AND2X2_3356 ( .A(AES_CORE_DATAPATH__abc_16259_n7683), .B(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n9293) );
  AND2X2 AND2X2_3357 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf4), .B(AES_CORE_DATAPATH_bkp_1_2__2_), .Y(AES_CORE_DATAPATH__abc_16259_n9295) );
  AND2X2 AND2X2_3358 ( .A(AES_CORE_DATAPATH__abc_16259_n7691), .B(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n9296) );
  AND2X2 AND2X2_3359 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1_2__3_), .Y(AES_CORE_DATAPATH__abc_16259_n9298) );
  AND2X2 AND2X2_336 ( .A(AES_CORE_DATAPATH__abc_16259_n2887_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__2_), .Y(AES_CORE_DATAPATH__abc_16259_n2928) );
  AND2X2 AND2X2_3360 ( .A(AES_CORE_DATAPATH__abc_16259_n7699), .B(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n9299) );
  AND2X2 AND2X2_3361 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf2), .B(AES_CORE_DATAPATH_bkp_1_2__4_), .Y(AES_CORE_DATAPATH__abc_16259_n9301) );
  AND2X2 AND2X2_3362 ( .A(AES_CORE_DATAPATH__abc_16259_n7707), .B(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n9302) );
  AND2X2 AND2X2_3363 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf1), .B(AES_CORE_DATAPATH_bkp_1_2__5_), .Y(AES_CORE_DATAPATH__abc_16259_n9304) );
  AND2X2 AND2X2_3364 ( .A(AES_CORE_DATAPATH__abc_16259_n7715), .B(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n9305) );
  AND2X2 AND2X2_3365 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf0), .B(AES_CORE_DATAPATH_bkp_1_2__6_), .Y(AES_CORE_DATAPATH__abc_16259_n9307) );
  AND2X2 AND2X2_3366 ( .A(AES_CORE_DATAPATH__abc_16259_n7723), .B(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n9308) );
  AND2X2 AND2X2_3367 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf6), .B(AES_CORE_DATAPATH_bkp_1_2__7_), .Y(AES_CORE_DATAPATH__abc_16259_n9310) );
  AND2X2 AND2X2_3368 ( .A(AES_CORE_DATAPATH__abc_16259_n7731), .B(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n9311) );
  AND2X2 AND2X2_3369 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf5), .B(AES_CORE_DATAPATH_bkp_1_2__8_), .Y(AES_CORE_DATAPATH__abc_16259_n9313) );
  AND2X2 AND2X2_337 ( .A(AES_CORE_DATAPATH__abc_16259_n2830_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__2_), .Y(AES_CORE_DATAPATH__abc_16259_n2929) );
  AND2X2 AND2X2_3370 ( .A(AES_CORE_DATAPATH__abc_16259_n7739), .B(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n9314) );
  AND2X2 AND2X2_3371 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf4), .B(AES_CORE_DATAPATH_bkp_1_2__9_), .Y(AES_CORE_DATAPATH__abc_16259_n9316) );
  AND2X2 AND2X2_3372 ( .A(AES_CORE_DATAPATH__abc_16259_n7747), .B(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n9317) );
  AND2X2 AND2X2_3373 ( .A(AES_CORE_DATAPATH__abc_16259_n7757), .B(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n9319) );
  AND2X2 AND2X2_3374 ( .A(AES_CORE_DATAPATH__abc_16259_n9320), .B(AES_CORE_DATAPATH__abc_16259_n9321), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__10_) );
  AND2X2 AND2X2_3375 ( .A(AES_CORE_DATAPATH__abc_16259_n7767), .B(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n9323) );
  AND2X2 AND2X2_3376 ( .A(AES_CORE_DATAPATH__abc_16259_n9324), .B(AES_CORE_DATAPATH__abc_16259_n9325), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__11_) );
  AND2X2 AND2X2_3377 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1_2__12_), .Y(AES_CORE_DATAPATH__abc_16259_n9327) );
  AND2X2 AND2X2_3378 ( .A(AES_CORE_DATAPATH__abc_16259_n7777), .B(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n9328) );
  AND2X2 AND2X2_3379 ( .A(AES_CORE_DATAPATH__abc_16259_n7786), .B(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n9330) );
  AND2X2 AND2X2_338 ( .A(AES_CORE_DATAPATH__abc_16259_n2931), .B(AES_CORE_DATAPATH__abc_16259_n2932), .Y(_auto_iopadmap_cc_313_execute_26949_2_) );
  AND2X2 AND2X2_3380 ( .A(AES_CORE_DATAPATH__abc_16259_n9331), .B(AES_CORE_DATAPATH__abc_16259_n9332), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__13_) );
  AND2X2 AND2X2_3381 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf2), .B(AES_CORE_DATAPATH_bkp_1_2__14_), .Y(AES_CORE_DATAPATH__abc_16259_n9334) );
  AND2X2 AND2X2_3382 ( .A(AES_CORE_DATAPATH__abc_16259_n7796), .B(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n9335) );
  AND2X2 AND2X2_3383 ( .A(AES_CORE_DATAPATH__abc_16259_n7805), .B(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n9337) );
  AND2X2 AND2X2_3384 ( .A(AES_CORE_DATAPATH__abc_16259_n9338), .B(AES_CORE_DATAPATH__abc_16259_n9339), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__15_) );
  AND2X2 AND2X2_3385 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf1), .B(AES_CORE_DATAPATH_bkp_1_2__16_), .Y(AES_CORE_DATAPATH__abc_16259_n9341) );
  AND2X2 AND2X2_3386 ( .A(AES_CORE_DATAPATH__abc_16259_n7815), .B(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n9342) );
  AND2X2 AND2X2_3387 ( .A(AES_CORE_DATAPATH__abc_16259_n7824), .B(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n9344) );
  AND2X2 AND2X2_3388 ( .A(AES_CORE_DATAPATH__abc_16259_n9345), .B(AES_CORE_DATAPATH__abc_16259_n9346), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__17_) );
  AND2X2 AND2X2_3389 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf0), .B(AES_CORE_DATAPATH_bkp_1_2__18_), .Y(AES_CORE_DATAPATH__abc_16259_n9348) );
  AND2X2 AND2X2_339 ( .A(AES_CORE_DATAPATH__abc_16259_n2855_bF_buf2), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_2_), .Y(AES_CORE_DATAPATH__abc_16259_n2935) );
  AND2X2 AND2X2_3390 ( .A(AES_CORE_DATAPATH__abc_16259_n7834), .B(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n9349) );
  AND2X2 AND2X2_3391 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf6), .B(AES_CORE_DATAPATH_bkp_1_2__19_), .Y(AES_CORE_DATAPATH__abc_16259_n9351) );
  AND2X2 AND2X2_3392 ( .A(AES_CORE_DATAPATH__abc_16259_n7842), .B(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n9352) );
  AND2X2 AND2X2_3393 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf5), .B(AES_CORE_DATAPATH_bkp_1_2__20_), .Y(AES_CORE_DATAPATH__abc_16259_n9354) );
  AND2X2 AND2X2_3394 ( .A(AES_CORE_DATAPATH__abc_16259_n7850), .B(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n9355) );
  AND2X2 AND2X2_3395 ( .A(AES_CORE_DATAPATH__abc_16259_n7859), .B(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n9357) );
  AND2X2 AND2X2_3396 ( .A(AES_CORE_DATAPATH__abc_16259_n9358), .B(AES_CORE_DATAPATH__abc_16259_n9359), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__21_) );
  AND2X2 AND2X2_3397 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf4), .B(AES_CORE_DATAPATH_bkp_1_2__22_), .Y(AES_CORE_DATAPATH__abc_16259_n9361) );
  AND2X2 AND2X2_3398 ( .A(AES_CORE_DATAPATH__abc_16259_n7869), .B(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n9362) );
  AND2X2 AND2X2_3399 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1_2__23_), .Y(AES_CORE_DATAPATH__abc_16259_n9364) );
  AND2X2 AND2X2_34 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n91), .B(AES_CORE_CONTROL_UNIT_state_7_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n122) );
  AND2X2 AND2X2_340 ( .A(AES_CORE_DATAPATH__abc_16259_n2857_bF_buf2), .B(AES_CORE_DATAPATH_MIX_COL_col_0__2_), .Y(AES_CORE_DATAPATH__abc_16259_n2936) );
  AND2X2 AND2X2_3400 ( .A(AES_CORE_DATAPATH__abc_16259_n7877), .B(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n9365) );
  AND2X2 AND2X2_3401 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf2), .B(AES_CORE_DATAPATH_bkp_1_2__24_), .Y(AES_CORE_DATAPATH__abc_16259_n9367) );
  AND2X2 AND2X2_3402 ( .A(AES_CORE_DATAPATH__abc_16259_n7885), .B(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n9368) );
  AND2X2 AND2X2_3403 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf1), .B(AES_CORE_DATAPATH_bkp_1_2__25_), .Y(AES_CORE_DATAPATH__abc_16259_n9370) );
  AND2X2 AND2X2_3404 ( .A(AES_CORE_DATAPATH__abc_16259_n7893), .B(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n9371) );
  AND2X2 AND2X2_3405 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf0), .B(AES_CORE_DATAPATH_bkp_1_2__26_), .Y(AES_CORE_DATAPATH__abc_16259_n9373) );
  AND2X2 AND2X2_3406 ( .A(AES_CORE_DATAPATH__abc_16259_n7901), .B(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n9374) );
  AND2X2 AND2X2_3407 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf6), .B(AES_CORE_DATAPATH_bkp_1_2__27_), .Y(AES_CORE_DATAPATH__abc_16259_n9376) );
  AND2X2 AND2X2_3408 ( .A(AES_CORE_DATAPATH__abc_16259_n7909), .B(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n9377) );
  AND2X2 AND2X2_3409 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf5), .B(AES_CORE_DATAPATH_bkp_1_2__28_), .Y(AES_CORE_DATAPATH__abc_16259_n9379) );
  AND2X2 AND2X2_341 ( .A(AES_CORE_DATAPATH__abc_16259_n2934), .B(AES_CORE_DATAPATH__abc_16259_n2938_1), .Y(AES_CORE_DATAPATH__abc_16259_n2939) );
  AND2X2 AND2X2_3410 ( .A(AES_CORE_DATAPATH__abc_16259_n7917), .B(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n9380) );
  AND2X2 AND2X2_3411 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf4), .B(AES_CORE_DATAPATH_bkp_1_2__29_), .Y(AES_CORE_DATAPATH__abc_16259_n9382) );
  AND2X2 AND2X2_3412 ( .A(AES_CORE_DATAPATH__abc_16259_n7925), .B(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n9383) );
  AND2X2 AND2X2_3413 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1_2__30_), .Y(AES_CORE_DATAPATH__abc_16259_n9385) );
  AND2X2 AND2X2_3414 ( .A(AES_CORE_DATAPATH__abc_16259_n7933), .B(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n9386) );
  AND2X2 AND2X2_3415 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf2), .B(AES_CORE_DATAPATH_bkp_1_2__31_), .Y(AES_CORE_DATAPATH__abc_16259_n9388) );
  AND2X2 AND2X2_3416 ( .A(AES_CORE_DATAPATH__abc_16259_n7941), .B(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n9389) );
  AND2X2 AND2X2_3417 ( .A(AES_CORE_DATAPATH__abc_16259_n9392), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n9393) );
  AND2X2 AND2X2_3418 ( .A(AES_CORE_DATAPATH__abc_16259_n9391), .B(AES_CORE_DATAPATH__abc_16259_n9393), .Y(AES_CORE_DATAPATH__abc_16259_n9394) );
  AND2X2 AND2X2_3419 ( .A(AES_CORE_DATAPATH__abc_16259_n9396), .B(AES_CORE_DATAPATH__abc_16259_n9397), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__0_) );
  AND2X2 AND2X2_342 ( .A(_auto_iopadmap_cc_313_execute_26949_2_), .B(AES_CORE_DATAPATH__abc_16259_n2939), .Y(AES_CORE_DATAPATH__abc_16259_n2942) );
  AND2X2 AND2X2_3420 ( .A(AES_CORE_DATAPATH__abc_16259_n9400), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n9401) );
  AND2X2 AND2X2_3421 ( .A(AES_CORE_DATAPATH__abc_16259_n9399), .B(AES_CORE_DATAPATH__abc_16259_n9401), .Y(AES_CORE_DATAPATH__abc_16259_n9402) );
  AND2X2 AND2X2_3422 ( .A(AES_CORE_DATAPATH__abc_16259_n9404), .B(AES_CORE_DATAPATH__abc_16259_n9405), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__1_) );
  AND2X2 AND2X2_3423 ( .A(AES_CORE_DATAPATH__abc_16259_n9408), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n9409) );
  AND2X2 AND2X2_3424 ( .A(AES_CORE_DATAPATH__abc_16259_n9407), .B(AES_CORE_DATAPATH__abc_16259_n9409), .Y(AES_CORE_DATAPATH__abc_16259_n9410) );
  AND2X2 AND2X2_3425 ( .A(AES_CORE_DATAPATH__abc_16259_n9412), .B(AES_CORE_DATAPATH__abc_16259_n9413), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__2_) );
  AND2X2 AND2X2_3426 ( .A(AES_CORE_DATAPATH__abc_16259_n9416), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n9417) );
  AND2X2 AND2X2_3427 ( .A(AES_CORE_DATAPATH__abc_16259_n9415), .B(AES_CORE_DATAPATH__abc_16259_n9417), .Y(AES_CORE_DATAPATH__abc_16259_n9418) );
  AND2X2 AND2X2_3428 ( .A(AES_CORE_DATAPATH__abc_16259_n9420), .B(AES_CORE_DATAPATH__abc_16259_n9421), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__3_) );
  AND2X2 AND2X2_3429 ( .A(AES_CORE_DATAPATH__abc_16259_n9424), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n9425) );
  AND2X2 AND2X2_343 ( .A(AES_CORE_DATAPATH_last_round_pp2_bF_buf1), .B(AES_CORE_DATAPATH_MIX_COL_col_0__2_), .Y(AES_CORE_DATAPATH__abc_16259_n2945_1) );
  AND2X2 AND2X2_3430 ( .A(AES_CORE_DATAPATH__abc_16259_n9423), .B(AES_CORE_DATAPATH__abc_16259_n9425), .Y(AES_CORE_DATAPATH__abc_16259_n9426) );
  AND2X2 AND2X2_3431 ( .A(AES_CORE_DATAPATH__abc_16259_n9428), .B(AES_CORE_DATAPATH__abc_16259_n9429), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__4_) );
  AND2X2 AND2X2_3432 ( .A(AES_CORE_DATAPATH__abc_16259_n9432), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n9433) );
  AND2X2 AND2X2_3433 ( .A(AES_CORE_DATAPATH__abc_16259_n9431), .B(AES_CORE_DATAPATH__abc_16259_n9433), .Y(AES_CORE_DATAPATH__abc_16259_n9434) );
  AND2X2 AND2X2_3434 ( .A(AES_CORE_DATAPATH__abc_16259_n9436), .B(AES_CORE_DATAPATH__abc_16259_n9437), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__5_) );
  AND2X2 AND2X2_3435 ( .A(AES_CORE_DATAPATH__abc_16259_n9440), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n9441) );
  AND2X2 AND2X2_3436 ( .A(AES_CORE_DATAPATH__abc_16259_n9439), .B(AES_CORE_DATAPATH__abc_16259_n9441), .Y(AES_CORE_DATAPATH__abc_16259_n9442) );
  AND2X2 AND2X2_3437 ( .A(AES_CORE_DATAPATH__abc_16259_n9444), .B(AES_CORE_DATAPATH__abc_16259_n9445), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__6_) );
  AND2X2 AND2X2_3438 ( .A(AES_CORE_DATAPATH__abc_16259_n9448), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf10), .Y(AES_CORE_DATAPATH__abc_16259_n9449) );
  AND2X2 AND2X2_3439 ( .A(AES_CORE_DATAPATH__abc_16259_n9447), .B(AES_CORE_DATAPATH__abc_16259_n9449), .Y(AES_CORE_DATAPATH__abc_16259_n9450) );
  AND2X2 AND2X2_344 ( .A(AES_CORE_DATAPATH__abc_16259_n2798_bF_buf2), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_2_), .Y(AES_CORE_DATAPATH__abc_16259_n2946_1) );
  AND2X2 AND2X2_3440 ( .A(AES_CORE_DATAPATH__abc_16259_n9452), .B(AES_CORE_DATAPATH__abc_16259_n9453), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__7_) );
  AND2X2 AND2X2_3441 ( .A(AES_CORE_DATAPATH__abc_16259_n9456), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf9), .Y(AES_CORE_DATAPATH__abc_16259_n9457) );
  AND2X2 AND2X2_3442 ( .A(AES_CORE_DATAPATH__abc_16259_n9455), .B(AES_CORE_DATAPATH__abc_16259_n9457), .Y(AES_CORE_DATAPATH__abc_16259_n9458) );
  AND2X2 AND2X2_3443 ( .A(AES_CORE_DATAPATH__abc_16259_n9460), .B(AES_CORE_DATAPATH__abc_16259_n9461), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__8_) );
  AND2X2 AND2X2_3444 ( .A(AES_CORE_DATAPATH__abc_16259_n9464), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf8), .Y(AES_CORE_DATAPATH__abc_16259_n9465) );
  AND2X2 AND2X2_3445 ( .A(AES_CORE_DATAPATH__abc_16259_n9463), .B(AES_CORE_DATAPATH__abc_16259_n9465), .Y(AES_CORE_DATAPATH__abc_16259_n9466) );
  AND2X2 AND2X2_3446 ( .A(AES_CORE_DATAPATH__abc_16259_n9468), .B(AES_CORE_DATAPATH__abc_16259_n9469), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__9_) );
  AND2X2 AND2X2_3447 ( .A(AES_CORE_DATAPATH__abc_16259_n7757), .B(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf9), .Y(AES_CORE_DATAPATH__abc_16259_n9471) );
  AND2X2 AND2X2_3448 ( .A(AES_CORE_DATAPATH__abc_16259_n9473), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n9474) );
  AND2X2 AND2X2_3449 ( .A(AES_CORE_DATAPATH__abc_16259_n9472), .B(AES_CORE_DATAPATH__abc_16259_n9474), .Y(AES_CORE_DATAPATH__abc_16259_n9475) );
  AND2X2 AND2X2_345 ( .A(AES_CORE_DATAPATH__abc_16259_n2944), .B(AES_CORE_DATAPATH__abc_16259_n2948), .Y(AES_CORE_DATAPATH__abc_16259_n2949_1) );
  AND2X2 AND2X2_3450 ( .A(AES_CORE_DATAPATH__abc_16259_n9477), .B(AES_CORE_DATAPATH__abc_16259_n9478), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__10_) );
  AND2X2 AND2X2_3451 ( .A(AES_CORE_DATAPATH__abc_16259_n7767), .B(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n9480) );
  AND2X2 AND2X2_3452 ( .A(AES_CORE_DATAPATH__abc_16259_n9482), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n9483) );
  AND2X2 AND2X2_3453 ( .A(AES_CORE_DATAPATH__abc_16259_n9481), .B(AES_CORE_DATAPATH__abc_16259_n9483), .Y(AES_CORE_DATAPATH__abc_16259_n9484) );
  AND2X2 AND2X2_3454 ( .A(AES_CORE_DATAPATH__abc_16259_n9486), .B(AES_CORE_DATAPATH__abc_16259_n9487), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__11_) );
  AND2X2 AND2X2_3455 ( .A(AES_CORE_DATAPATH__abc_16259_n9490), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n9491) );
  AND2X2 AND2X2_3456 ( .A(AES_CORE_DATAPATH__abc_16259_n9489), .B(AES_CORE_DATAPATH__abc_16259_n9491), .Y(AES_CORE_DATAPATH__abc_16259_n9492) );
  AND2X2 AND2X2_3457 ( .A(AES_CORE_DATAPATH__abc_16259_n9494), .B(AES_CORE_DATAPATH__abc_16259_n9495), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__12_) );
  AND2X2 AND2X2_3458 ( .A(AES_CORE_DATAPATH__abc_16259_n7786), .B(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n9497) );
  AND2X2 AND2X2_3459 ( .A(AES_CORE_DATAPATH__abc_16259_n9499), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n9500) );
  AND2X2 AND2X2_346 ( .A(AES_CORE_DATAPATH__abc_16259_n2949_1), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n2950) );
  AND2X2 AND2X2_3460 ( .A(AES_CORE_DATAPATH__abc_16259_n9498), .B(AES_CORE_DATAPATH__abc_16259_n9500), .Y(AES_CORE_DATAPATH__abc_16259_n9501) );
  AND2X2 AND2X2_3461 ( .A(AES_CORE_DATAPATH__abc_16259_n9503), .B(AES_CORE_DATAPATH__abc_16259_n9504), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__13_) );
  AND2X2 AND2X2_3462 ( .A(AES_CORE_DATAPATH__abc_16259_n9507), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n9508) );
  AND2X2 AND2X2_3463 ( .A(AES_CORE_DATAPATH__abc_16259_n9506), .B(AES_CORE_DATAPATH__abc_16259_n9508), .Y(AES_CORE_DATAPATH__abc_16259_n9509) );
  AND2X2 AND2X2_3464 ( .A(AES_CORE_DATAPATH__abc_16259_n9511), .B(AES_CORE_DATAPATH__abc_16259_n9512), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__14_) );
  AND2X2 AND2X2_3465 ( .A(AES_CORE_DATAPATH__abc_16259_n7805), .B(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n9514) );
  AND2X2 AND2X2_3466 ( .A(AES_CORE_DATAPATH__abc_16259_n9516), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n9517) );
  AND2X2 AND2X2_3467 ( .A(AES_CORE_DATAPATH__abc_16259_n9515), .B(AES_CORE_DATAPATH__abc_16259_n9517), .Y(AES_CORE_DATAPATH__abc_16259_n9518) );
  AND2X2 AND2X2_3468 ( .A(AES_CORE_DATAPATH__abc_16259_n9520), .B(AES_CORE_DATAPATH__abc_16259_n9521), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__15_) );
  AND2X2 AND2X2_3469 ( .A(AES_CORE_DATAPATH__abc_16259_n9524), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n9525) );
  AND2X2 AND2X2_347 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf9), .B(AES_CORE_DATAPATH_col_3__2_), .Y(AES_CORE_DATAPATH__abc_16259_n2951_1) );
  AND2X2 AND2X2_3470 ( .A(AES_CORE_DATAPATH__abc_16259_n9523), .B(AES_CORE_DATAPATH__abc_16259_n9525), .Y(AES_CORE_DATAPATH__abc_16259_n9526) );
  AND2X2 AND2X2_3471 ( .A(AES_CORE_DATAPATH__abc_16259_n9528), .B(AES_CORE_DATAPATH__abc_16259_n9529), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__16_) );
  AND2X2 AND2X2_3472 ( .A(AES_CORE_DATAPATH__abc_16259_n7824), .B(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf10), .Y(AES_CORE_DATAPATH__abc_16259_n9531) );
  AND2X2 AND2X2_3473 ( .A(AES_CORE_DATAPATH__abc_16259_n9533), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n9534) );
  AND2X2 AND2X2_3474 ( .A(AES_CORE_DATAPATH__abc_16259_n9532), .B(AES_CORE_DATAPATH__abc_16259_n9534), .Y(AES_CORE_DATAPATH__abc_16259_n9535) );
  AND2X2 AND2X2_3475 ( .A(AES_CORE_DATAPATH__abc_16259_n9537), .B(AES_CORE_DATAPATH__abc_16259_n9538), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__17_) );
  AND2X2 AND2X2_3476 ( .A(AES_CORE_DATAPATH__abc_16259_n9541), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf10), .Y(AES_CORE_DATAPATH__abc_16259_n9542) );
  AND2X2 AND2X2_3477 ( .A(AES_CORE_DATAPATH__abc_16259_n9540), .B(AES_CORE_DATAPATH__abc_16259_n9542), .Y(AES_CORE_DATAPATH__abc_16259_n9543) );
  AND2X2 AND2X2_3478 ( .A(AES_CORE_DATAPATH__abc_16259_n9545), .B(AES_CORE_DATAPATH__abc_16259_n9546), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__18_) );
  AND2X2 AND2X2_3479 ( .A(AES_CORE_DATAPATH__abc_16259_n9549), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf9), .Y(AES_CORE_DATAPATH__abc_16259_n9550) );
  AND2X2 AND2X2_348 ( .A(AES_CORE_DATAPATH__abc_16259_n2954), .B(AES_CORE_DATAPATH__abc_16259_n2956), .Y(AES_CORE_DATAPATH__abc_16259_n2957) );
  AND2X2 AND2X2_3480 ( .A(AES_CORE_DATAPATH__abc_16259_n9548), .B(AES_CORE_DATAPATH__abc_16259_n9550), .Y(AES_CORE_DATAPATH__abc_16259_n9551) );
  AND2X2 AND2X2_3481 ( .A(AES_CORE_DATAPATH__abc_16259_n9553), .B(AES_CORE_DATAPATH__abc_16259_n9554), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__19_) );
  AND2X2 AND2X2_3482 ( .A(AES_CORE_DATAPATH__abc_16259_n9557), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf8), .Y(AES_CORE_DATAPATH__abc_16259_n9558) );
  AND2X2 AND2X2_3483 ( .A(AES_CORE_DATAPATH__abc_16259_n9556), .B(AES_CORE_DATAPATH__abc_16259_n9558), .Y(AES_CORE_DATAPATH__abc_16259_n9559) );
  AND2X2 AND2X2_3484 ( .A(AES_CORE_DATAPATH__abc_16259_n9561), .B(AES_CORE_DATAPATH__abc_16259_n9562), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__20_) );
  AND2X2 AND2X2_3485 ( .A(AES_CORE_DATAPATH__abc_16259_n7859), .B(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n9564) );
  AND2X2 AND2X2_3486 ( .A(AES_CORE_DATAPATH__abc_16259_n9566), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n9567) );
  AND2X2 AND2X2_3487 ( .A(AES_CORE_DATAPATH__abc_16259_n9565), .B(AES_CORE_DATAPATH__abc_16259_n9567), .Y(AES_CORE_DATAPATH__abc_16259_n9568) );
  AND2X2 AND2X2_3488 ( .A(AES_CORE_DATAPATH__abc_16259_n9570), .B(AES_CORE_DATAPATH__abc_16259_n9571), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__21_) );
  AND2X2 AND2X2_3489 ( .A(AES_CORE_DATAPATH__abc_16259_n9574), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n9575) );
  AND2X2 AND2X2_349 ( .A(AES_CORE_DATAPATH__abc_16259_n2782_bF_buf1), .B(AES_CORE_DATAPATH_col_3__3_), .Y(AES_CORE_DATAPATH__abc_16259_n2958) );
  AND2X2 AND2X2_3490 ( .A(AES_CORE_DATAPATH__abc_16259_n9573), .B(AES_CORE_DATAPATH__abc_16259_n9575), .Y(AES_CORE_DATAPATH__abc_16259_n9576) );
  AND2X2 AND2X2_3491 ( .A(AES_CORE_DATAPATH__abc_16259_n9578), .B(AES_CORE_DATAPATH__abc_16259_n9579), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__22_) );
  AND2X2 AND2X2_3492 ( .A(AES_CORE_DATAPATH__abc_16259_n9582), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n9583) );
  AND2X2 AND2X2_3493 ( .A(AES_CORE_DATAPATH__abc_16259_n9581), .B(AES_CORE_DATAPATH__abc_16259_n9583), .Y(AES_CORE_DATAPATH__abc_16259_n9584) );
  AND2X2 AND2X2_3494 ( .A(AES_CORE_DATAPATH__abc_16259_n9586), .B(AES_CORE_DATAPATH__abc_16259_n9587), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__23_) );
  AND2X2 AND2X2_3495 ( .A(AES_CORE_DATAPATH__abc_16259_n9590), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n9591) );
  AND2X2 AND2X2_3496 ( .A(AES_CORE_DATAPATH__abc_16259_n9589), .B(AES_CORE_DATAPATH__abc_16259_n9591), .Y(AES_CORE_DATAPATH__abc_16259_n9592) );
  AND2X2 AND2X2_3497 ( .A(AES_CORE_DATAPATH__abc_16259_n9594), .B(AES_CORE_DATAPATH__abc_16259_n9595), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__24_) );
  AND2X2 AND2X2_3498 ( .A(AES_CORE_DATAPATH__abc_16259_n9598), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n9599) );
  AND2X2 AND2X2_3499 ( .A(AES_CORE_DATAPATH__abc_16259_n9597), .B(AES_CORE_DATAPATH__abc_16259_n9599), .Y(AES_CORE_DATAPATH__abc_16259_n9600) );
  AND2X2 AND2X2_35 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf12), .B(AES_CORE_CONTROL_UNIT_state_9_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n124_1) );
  AND2X2 AND2X2_350 ( .A(AES_CORE_DATAPATH__abc_16259_n2786_bF_buf1), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_67_), .Y(AES_CORE_DATAPATH__abc_16259_n2959) );
  AND2X2 AND2X2_3500 ( .A(AES_CORE_DATAPATH__abc_16259_n9602), .B(AES_CORE_DATAPATH__abc_16259_n9603), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__25_) );
  AND2X2 AND2X2_3501 ( .A(AES_CORE_DATAPATH__abc_16259_n9606), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n9607) );
  AND2X2 AND2X2_3502 ( .A(AES_CORE_DATAPATH__abc_16259_n9605), .B(AES_CORE_DATAPATH__abc_16259_n9607), .Y(AES_CORE_DATAPATH__abc_16259_n9608) );
  AND2X2 AND2X2_3503 ( .A(AES_CORE_DATAPATH__abc_16259_n9610), .B(AES_CORE_DATAPATH__abc_16259_n9611), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__26_) );
  AND2X2 AND2X2_3504 ( .A(AES_CORE_DATAPATH__abc_16259_n9614), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n9615) );
  AND2X2 AND2X2_3505 ( .A(AES_CORE_DATAPATH__abc_16259_n9613), .B(AES_CORE_DATAPATH__abc_16259_n9615), .Y(AES_CORE_DATAPATH__abc_16259_n9616) );
  AND2X2 AND2X2_3506 ( .A(AES_CORE_DATAPATH__abc_16259_n9618), .B(AES_CORE_DATAPATH__abc_16259_n9619), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__27_) );
  AND2X2 AND2X2_3507 ( .A(AES_CORE_DATAPATH__abc_16259_n9622), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n9623) );
  AND2X2 AND2X2_3508 ( .A(AES_CORE_DATAPATH__abc_16259_n9621), .B(AES_CORE_DATAPATH__abc_16259_n9623), .Y(AES_CORE_DATAPATH__abc_16259_n9624) );
  AND2X2 AND2X2_3509 ( .A(AES_CORE_DATAPATH__abc_16259_n9626), .B(AES_CORE_DATAPATH__abc_16259_n9627), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__28_) );
  AND2X2 AND2X2_351 ( .A(AES_CORE_DATAPATH__abc_16259_n2789_bF_buf1), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_35_), .Y(AES_CORE_DATAPATH__abc_16259_n2960) );
  AND2X2 AND2X2_3510 ( .A(AES_CORE_DATAPATH__abc_16259_n9630), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf10), .Y(AES_CORE_DATAPATH__abc_16259_n9631) );
  AND2X2 AND2X2_3511 ( .A(AES_CORE_DATAPATH__abc_16259_n9629), .B(AES_CORE_DATAPATH__abc_16259_n9631), .Y(AES_CORE_DATAPATH__abc_16259_n9632) );
  AND2X2 AND2X2_3512 ( .A(AES_CORE_DATAPATH__abc_16259_n9634), .B(AES_CORE_DATAPATH__abc_16259_n9635), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__29_) );
  AND2X2 AND2X2_3513 ( .A(AES_CORE_DATAPATH__abc_16259_n9638), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf9), .Y(AES_CORE_DATAPATH__abc_16259_n9639) );
  AND2X2 AND2X2_3514 ( .A(AES_CORE_DATAPATH__abc_16259_n9637), .B(AES_CORE_DATAPATH__abc_16259_n9639), .Y(AES_CORE_DATAPATH__abc_16259_n9640) );
  AND2X2 AND2X2_3515 ( .A(AES_CORE_DATAPATH__abc_16259_n9642), .B(AES_CORE_DATAPATH__abc_16259_n9643), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__30_) );
  AND2X2 AND2X2_3516 ( .A(AES_CORE_DATAPATH__abc_16259_n9646), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf8), .Y(AES_CORE_DATAPATH__abc_16259_n9647) );
  AND2X2 AND2X2_3517 ( .A(AES_CORE_DATAPATH__abc_16259_n9645), .B(AES_CORE_DATAPATH__abc_16259_n9647), .Y(AES_CORE_DATAPATH__abc_16259_n9648) );
  AND2X2 AND2X2_3518 ( .A(AES_CORE_DATAPATH__abc_16259_n9650), .B(AES_CORE_DATAPATH__abc_16259_n9651), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__31_) );
  AND2X2 AND2X2_3519 ( .A(AES_CORE_DATAPATH__abc_16259_n9655), .B(AES_CORE_DATAPATH__abc_16259_n9653), .Y(AES_CORE_DATAPATH__0iv_2__31_0__0_) );
  AND2X2 AND2X2_352 ( .A(AES_CORE_DATAPATH__abc_16259_n2963), .B(AES_CORE_DATAPATH__abc_16259_n2957), .Y(AES_CORE_DATAPATH__abc_16259_n2964) );
  AND2X2 AND2X2_3520 ( .A(AES_CORE_DATAPATH__abc_16259_n9658), .B(AES_CORE_DATAPATH__abc_16259_n9657), .Y(AES_CORE_DATAPATH__0iv_2__31_0__1_) );
  AND2X2 AND2X2_3521 ( .A(AES_CORE_DATAPATH__abc_16259_n9661), .B(AES_CORE_DATAPATH__abc_16259_n9660), .Y(AES_CORE_DATAPATH__0iv_2__31_0__2_) );
  AND2X2 AND2X2_3522 ( .A(AES_CORE_DATAPATH__abc_16259_n9664), .B(AES_CORE_DATAPATH__abc_16259_n9663), .Y(AES_CORE_DATAPATH__0iv_2__31_0__3_) );
  AND2X2 AND2X2_3523 ( .A(AES_CORE_DATAPATH__abc_16259_n9667), .B(AES_CORE_DATAPATH__abc_16259_n9666), .Y(AES_CORE_DATAPATH__0iv_2__31_0__4_) );
  AND2X2 AND2X2_3524 ( .A(AES_CORE_DATAPATH__abc_16259_n9670), .B(AES_CORE_DATAPATH__abc_16259_n9669), .Y(AES_CORE_DATAPATH__0iv_2__31_0__5_) );
  AND2X2 AND2X2_3525 ( .A(AES_CORE_DATAPATH__abc_16259_n9673), .B(AES_CORE_DATAPATH__abc_16259_n9672), .Y(AES_CORE_DATAPATH__0iv_2__31_0__6_) );
  AND2X2 AND2X2_3526 ( .A(AES_CORE_DATAPATH__abc_16259_n9676), .B(AES_CORE_DATAPATH__abc_16259_n9675), .Y(AES_CORE_DATAPATH__0iv_2__31_0__7_) );
  AND2X2 AND2X2_3527 ( .A(AES_CORE_DATAPATH__abc_16259_n9679), .B(AES_CORE_DATAPATH__abc_16259_n9678), .Y(AES_CORE_DATAPATH__0iv_2__31_0__8_) );
  AND2X2 AND2X2_3528 ( .A(AES_CORE_DATAPATH__abc_16259_n9682), .B(AES_CORE_DATAPATH__abc_16259_n9681), .Y(AES_CORE_DATAPATH__0iv_2__31_0__9_) );
  AND2X2 AND2X2_3529 ( .A(AES_CORE_DATAPATH__abc_16259_n9685), .B(AES_CORE_DATAPATH__abc_16259_n9684), .Y(AES_CORE_DATAPATH__0iv_2__31_0__10_) );
  AND2X2 AND2X2_353 ( .A(AES_CORE_DATAPATH__abc_16259_n2837_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__3_), .Y(AES_CORE_DATAPATH__abc_16259_n2966) );
  AND2X2 AND2X2_3530 ( .A(AES_CORE_DATAPATH__abc_16259_n9688), .B(AES_CORE_DATAPATH__abc_16259_n9687), .Y(AES_CORE_DATAPATH__0iv_2__31_0__11_) );
  AND2X2 AND2X2_3531 ( .A(AES_CORE_DATAPATH__abc_16259_n9691), .B(AES_CORE_DATAPATH__abc_16259_n9690), .Y(AES_CORE_DATAPATH__0iv_2__31_0__12_) );
  AND2X2 AND2X2_3532 ( .A(AES_CORE_DATAPATH__abc_16259_n9694), .B(AES_CORE_DATAPATH__abc_16259_n9693), .Y(AES_CORE_DATAPATH__0iv_2__31_0__13_) );
  AND2X2 AND2X2_3533 ( .A(AES_CORE_DATAPATH__abc_16259_n9697), .B(AES_CORE_DATAPATH__abc_16259_n9696), .Y(AES_CORE_DATAPATH__0iv_2__31_0__14_) );
  AND2X2 AND2X2_3534 ( .A(AES_CORE_DATAPATH__abc_16259_n9700), .B(AES_CORE_DATAPATH__abc_16259_n9699), .Y(AES_CORE_DATAPATH__0iv_2__31_0__15_) );
  AND2X2 AND2X2_3535 ( .A(AES_CORE_DATAPATH__abc_16259_n9703), .B(AES_CORE_DATAPATH__abc_16259_n9702), .Y(AES_CORE_DATAPATH__0iv_2__31_0__16_) );
  AND2X2 AND2X2_3536 ( .A(AES_CORE_DATAPATH__abc_16259_n9706), .B(AES_CORE_DATAPATH__abc_16259_n9705), .Y(AES_CORE_DATAPATH__0iv_2__31_0__17_) );
  AND2X2 AND2X2_3537 ( .A(AES_CORE_DATAPATH__abc_16259_n9709), .B(AES_CORE_DATAPATH__abc_16259_n9708), .Y(AES_CORE_DATAPATH__0iv_2__31_0__18_) );
  AND2X2 AND2X2_3538 ( .A(AES_CORE_DATAPATH__abc_16259_n9712), .B(AES_CORE_DATAPATH__abc_16259_n9711), .Y(AES_CORE_DATAPATH__0iv_2__31_0__19_) );
  AND2X2 AND2X2_3539 ( .A(AES_CORE_DATAPATH__abc_16259_n9715), .B(AES_CORE_DATAPATH__abc_16259_n9714), .Y(AES_CORE_DATAPATH__0iv_2__31_0__20_) );
  AND2X2 AND2X2_354 ( .A(AES_CORE_DATAPATH__abc_16259_n2887_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__3_), .Y(AES_CORE_DATAPATH__abc_16259_n2968) );
  AND2X2 AND2X2_3540 ( .A(AES_CORE_DATAPATH__abc_16259_n9718), .B(AES_CORE_DATAPATH__abc_16259_n9717), .Y(AES_CORE_DATAPATH__0iv_2__31_0__21_) );
  AND2X2 AND2X2_3541 ( .A(AES_CORE_DATAPATH__abc_16259_n9721), .B(AES_CORE_DATAPATH__abc_16259_n9720), .Y(AES_CORE_DATAPATH__0iv_2__31_0__22_) );
  AND2X2 AND2X2_3542 ( .A(AES_CORE_DATAPATH__abc_16259_n9724), .B(AES_CORE_DATAPATH__abc_16259_n9723), .Y(AES_CORE_DATAPATH__0iv_2__31_0__23_) );
  AND2X2 AND2X2_3543 ( .A(AES_CORE_DATAPATH__abc_16259_n9727), .B(AES_CORE_DATAPATH__abc_16259_n9726), .Y(AES_CORE_DATAPATH__0iv_2__31_0__24_) );
  AND2X2 AND2X2_3544 ( .A(AES_CORE_DATAPATH__abc_16259_n9730), .B(AES_CORE_DATAPATH__abc_16259_n9729), .Y(AES_CORE_DATAPATH__0iv_2__31_0__25_) );
  AND2X2 AND2X2_3545 ( .A(AES_CORE_DATAPATH__abc_16259_n9733), .B(AES_CORE_DATAPATH__abc_16259_n9732), .Y(AES_CORE_DATAPATH__0iv_2__31_0__26_) );
  AND2X2 AND2X2_3546 ( .A(AES_CORE_DATAPATH__abc_16259_n9736), .B(AES_CORE_DATAPATH__abc_16259_n9735), .Y(AES_CORE_DATAPATH__0iv_2__31_0__27_) );
  AND2X2 AND2X2_3547 ( .A(AES_CORE_DATAPATH__abc_16259_n9739), .B(AES_CORE_DATAPATH__abc_16259_n9738), .Y(AES_CORE_DATAPATH__0iv_2__31_0__28_) );
  AND2X2 AND2X2_3548 ( .A(AES_CORE_DATAPATH__abc_16259_n9742), .B(AES_CORE_DATAPATH__abc_16259_n9741), .Y(AES_CORE_DATAPATH__0iv_2__31_0__29_) );
  AND2X2 AND2X2_3549 ( .A(AES_CORE_DATAPATH__abc_16259_n9745), .B(AES_CORE_DATAPATH__abc_16259_n9744), .Y(AES_CORE_DATAPATH__0iv_2__31_0__30_) );
  AND2X2 AND2X2_355 ( .A(AES_CORE_DATAPATH__abc_16259_n2830_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__3_), .Y(AES_CORE_DATAPATH__abc_16259_n2969_1) );
  AND2X2 AND2X2_3550 ( .A(AES_CORE_DATAPATH__abc_16259_n9748), .B(AES_CORE_DATAPATH__abc_16259_n9747), .Y(AES_CORE_DATAPATH__0iv_2__31_0__31_) );
  AND2X2 AND2X2_3551 ( .A(AES_CORE_DATAPATH__abc_16259_n8494), .B(AES_CORE_DATAPATH_col_en_host_1_), .Y(AES_CORE_DATAPATH__abc_16259_n9750) );
  AND2X2 AND2X2_3552 ( .A(AES_CORE_DATAPATH__abc_16259_n8497), .B(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_1_), .Y(AES_CORE_DATAPATH__abc_16259_n9751) );
  AND2X2 AND2X2_3553 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf6), .B(AES_CORE_DATAPATH_bkp_1_1__0_), .Y(AES_CORE_DATAPATH__abc_16259_n9754) );
  AND2X2 AND2X2_3554 ( .A(AES_CORE_DATAPATH__abc_16259_n7950), .B(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n9755) );
  AND2X2 AND2X2_3555 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf5), .B(AES_CORE_DATAPATH_bkp_1_1__1_), .Y(AES_CORE_DATAPATH__abc_16259_n9757) );
  AND2X2 AND2X2_3556 ( .A(AES_CORE_DATAPATH__abc_16259_n7958), .B(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n9758) );
  AND2X2 AND2X2_3557 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf4), .B(AES_CORE_DATAPATH_bkp_1_1__2_), .Y(AES_CORE_DATAPATH__abc_16259_n9760) );
  AND2X2 AND2X2_3558 ( .A(AES_CORE_DATAPATH__abc_16259_n7966), .B(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n9761) );
  AND2X2 AND2X2_3559 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1_1__3_), .Y(AES_CORE_DATAPATH__abc_16259_n9763) );
  AND2X2 AND2X2_356 ( .A(AES_CORE_DATAPATH__abc_16259_n2971), .B(AES_CORE_DATAPATH__abc_16259_n2972), .Y(_auto_iopadmap_cc_313_execute_26949_3_) );
  AND2X2 AND2X2_3560 ( .A(AES_CORE_DATAPATH__abc_16259_n7974), .B(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n9764) );
  AND2X2 AND2X2_3561 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf2), .B(AES_CORE_DATAPATH_bkp_1_1__4_), .Y(AES_CORE_DATAPATH__abc_16259_n9766) );
  AND2X2 AND2X2_3562 ( .A(AES_CORE_DATAPATH__abc_16259_n7982), .B(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n9767) );
  AND2X2 AND2X2_3563 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf1), .B(AES_CORE_DATAPATH_bkp_1_1__5_), .Y(AES_CORE_DATAPATH__abc_16259_n9769) );
  AND2X2 AND2X2_3564 ( .A(AES_CORE_DATAPATH__abc_16259_n7990), .B(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n9770) );
  AND2X2 AND2X2_3565 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf0), .B(AES_CORE_DATAPATH_bkp_1_1__6_), .Y(AES_CORE_DATAPATH__abc_16259_n9772) );
  AND2X2 AND2X2_3566 ( .A(AES_CORE_DATAPATH__abc_16259_n7998), .B(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n9773) );
  AND2X2 AND2X2_3567 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf6), .B(AES_CORE_DATAPATH_bkp_1_1__7_), .Y(AES_CORE_DATAPATH__abc_16259_n9775) );
  AND2X2 AND2X2_3568 ( .A(AES_CORE_DATAPATH__abc_16259_n8006), .B(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n9776) );
  AND2X2 AND2X2_3569 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf5), .B(AES_CORE_DATAPATH_bkp_1_1__8_), .Y(AES_CORE_DATAPATH__abc_16259_n9778) );
  AND2X2 AND2X2_357 ( .A(AES_CORE_DATAPATH__abc_16259_n2855_bF_buf1), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_3_), .Y(AES_CORE_DATAPATH__abc_16259_n2975_1) );
  AND2X2 AND2X2_3570 ( .A(AES_CORE_DATAPATH__abc_16259_n8014), .B(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n9779) );
  AND2X2 AND2X2_3571 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf4), .B(AES_CORE_DATAPATH_bkp_1_1__9_), .Y(AES_CORE_DATAPATH__abc_16259_n9781) );
  AND2X2 AND2X2_3572 ( .A(AES_CORE_DATAPATH__abc_16259_n8022), .B(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n9782) );
  AND2X2 AND2X2_3573 ( .A(AES_CORE_DATAPATH__abc_16259_n8031), .B(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n9784) );
  AND2X2 AND2X2_3574 ( .A(AES_CORE_DATAPATH__abc_16259_n9785), .B(AES_CORE_DATAPATH__abc_16259_n9786), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__10_) );
  AND2X2 AND2X2_3575 ( .A(AES_CORE_DATAPATH__abc_16259_n8043), .B(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n9788) );
  AND2X2 AND2X2_3576 ( .A(AES_CORE_DATAPATH__abc_16259_n9789), .B(AES_CORE_DATAPATH__abc_16259_n9790), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__11_) );
  AND2X2 AND2X2_3577 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1_1__12_), .Y(AES_CORE_DATAPATH__abc_16259_n9792) );
  AND2X2 AND2X2_3578 ( .A(AES_CORE_DATAPATH__abc_16259_n8052), .B(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n9793) );
  AND2X2 AND2X2_3579 ( .A(AES_CORE_DATAPATH__abc_16259_n8061), .B(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n9795) );
  AND2X2 AND2X2_358 ( .A(AES_CORE_DATAPATH__abc_16259_n2857_bF_buf1), .B(AES_CORE_DATAPATH_MIX_COL_col_0__3_), .Y(AES_CORE_DATAPATH__abc_16259_n2976) );
  AND2X2 AND2X2_3580 ( .A(AES_CORE_DATAPATH__abc_16259_n9796), .B(AES_CORE_DATAPATH__abc_16259_n9797), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__13_) );
  AND2X2 AND2X2_3581 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf2), .B(AES_CORE_DATAPATH_bkp_1_1__14_), .Y(AES_CORE_DATAPATH__abc_16259_n9799) );
  AND2X2 AND2X2_3582 ( .A(AES_CORE_DATAPATH__abc_16259_n8071), .B(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n9800) );
  AND2X2 AND2X2_3583 ( .A(AES_CORE_DATAPATH__abc_16259_n8080), .B(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n9802) );
  AND2X2 AND2X2_3584 ( .A(AES_CORE_DATAPATH__abc_16259_n9803), .B(AES_CORE_DATAPATH__abc_16259_n9804), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__15_) );
  AND2X2 AND2X2_3585 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf1), .B(AES_CORE_DATAPATH_bkp_1_1__16_), .Y(AES_CORE_DATAPATH__abc_16259_n9806) );
  AND2X2 AND2X2_3586 ( .A(AES_CORE_DATAPATH__abc_16259_n8090), .B(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n9807) );
  AND2X2 AND2X2_3587 ( .A(AES_CORE_DATAPATH__abc_16259_n8099), .B(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n9809) );
  AND2X2 AND2X2_3588 ( .A(AES_CORE_DATAPATH__abc_16259_n9810), .B(AES_CORE_DATAPATH__abc_16259_n9811), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__17_) );
  AND2X2 AND2X2_3589 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf0), .B(AES_CORE_DATAPATH_bkp_1_1__18_), .Y(AES_CORE_DATAPATH__abc_16259_n9813) );
  AND2X2 AND2X2_359 ( .A(AES_CORE_DATAPATH__abc_16259_n2974_1), .B(AES_CORE_DATAPATH__abc_16259_n2978_1), .Y(AES_CORE_DATAPATH__abc_16259_n2979) );
  AND2X2 AND2X2_3590 ( .A(AES_CORE_DATAPATH__abc_16259_n8109), .B(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n9814) );
  AND2X2 AND2X2_3591 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf6), .B(AES_CORE_DATAPATH_bkp_1_1__19_), .Y(AES_CORE_DATAPATH__abc_16259_n9816) );
  AND2X2 AND2X2_3592 ( .A(AES_CORE_DATAPATH__abc_16259_n8117), .B(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n9817) );
  AND2X2 AND2X2_3593 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf5), .B(AES_CORE_DATAPATH_bkp_1_1__20_), .Y(AES_CORE_DATAPATH__abc_16259_n9819) );
  AND2X2 AND2X2_3594 ( .A(AES_CORE_DATAPATH__abc_16259_n8125), .B(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n9820) );
  AND2X2 AND2X2_3595 ( .A(AES_CORE_DATAPATH__abc_16259_n8134), .B(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n9822) );
  AND2X2 AND2X2_3596 ( .A(AES_CORE_DATAPATH__abc_16259_n9823), .B(AES_CORE_DATAPATH__abc_16259_n9824), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__21_) );
  AND2X2 AND2X2_3597 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf4), .B(AES_CORE_DATAPATH_bkp_1_1__22_), .Y(AES_CORE_DATAPATH__abc_16259_n9826) );
  AND2X2 AND2X2_3598 ( .A(AES_CORE_DATAPATH__abc_16259_n8144), .B(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n9827) );
  AND2X2 AND2X2_3599 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1_1__23_), .Y(AES_CORE_DATAPATH__abc_16259_n9829) );
  AND2X2 AND2X2_36 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n125), .B(AES_CORE_CONTROL_UNIT__abc_15841_n87_1), .Y(AES_CORE_CONTROL_UNIT__abc_10818_n29) );
  AND2X2 AND2X2_360 ( .A(_auto_iopadmap_cc_313_execute_26949_3_), .B(AES_CORE_DATAPATH__abc_16259_n2979), .Y(AES_CORE_DATAPATH__abc_16259_n2982_1) );
  AND2X2 AND2X2_3600 ( .A(AES_CORE_DATAPATH__abc_16259_n8152), .B(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n9830) );
  AND2X2 AND2X2_3601 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf2), .B(AES_CORE_DATAPATH_bkp_1_1__24_), .Y(AES_CORE_DATAPATH__abc_16259_n9832) );
  AND2X2 AND2X2_3602 ( .A(AES_CORE_DATAPATH__abc_16259_n8160), .B(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n9833) );
  AND2X2 AND2X2_3603 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf1), .B(AES_CORE_DATAPATH_bkp_1_1__25_), .Y(AES_CORE_DATAPATH__abc_16259_n9835) );
  AND2X2 AND2X2_3604 ( .A(AES_CORE_DATAPATH__abc_16259_n8168), .B(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n9836) );
  AND2X2 AND2X2_3605 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf0), .B(AES_CORE_DATAPATH_bkp_1_1__26_), .Y(AES_CORE_DATAPATH__abc_16259_n9838) );
  AND2X2 AND2X2_3606 ( .A(AES_CORE_DATAPATH__abc_16259_n8176), .B(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n9839) );
  AND2X2 AND2X2_3607 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf6), .B(AES_CORE_DATAPATH_bkp_1_1__27_), .Y(AES_CORE_DATAPATH__abc_16259_n9841) );
  AND2X2 AND2X2_3608 ( .A(AES_CORE_DATAPATH__abc_16259_n8184), .B(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n9842) );
  AND2X2 AND2X2_3609 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf5), .B(AES_CORE_DATAPATH_bkp_1_1__28_), .Y(AES_CORE_DATAPATH__abc_16259_n9844) );
  AND2X2 AND2X2_361 ( .A(AES_CORE_DATAPATH_last_round_pp2_bF_buf0), .B(AES_CORE_DATAPATH_MIX_COL_col_0__3_), .Y(AES_CORE_DATAPATH__abc_16259_n2985) );
  AND2X2 AND2X2_3610 ( .A(AES_CORE_DATAPATH__abc_16259_n8192), .B(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n9845) );
  AND2X2 AND2X2_3611 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf4), .B(AES_CORE_DATAPATH_bkp_1_1__29_), .Y(AES_CORE_DATAPATH__abc_16259_n9847) );
  AND2X2 AND2X2_3612 ( .A(AES_CORE_DATAPATH__abc_16259_n8200), .B(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n9848) );
  AND2X2 AND2X2_3613 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1_1__30_), .Y(AES_CORE_DATAPATH__abc_16259_n9850) );
  AND2X2 AND2X2_3614 ( .A(AES_CORE_DATAPATH__abc_16259_n8208), .B(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n9851) );
  AND2X2 AND2X2_3615 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf2), .B(AES_CORE_DATAPATH_bkp_1_1__31_), .Y(AES_CORE_DATAPATH__abc_16259_n9853) );
  AND2X2 AND2X2_3616 ( .A(AES_CORE_DATAPATH__abc_16259_n8216), .B(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n9854) );
  AND2X2 AND2X2_3617 ( .A(AES_CORE_DATAPATH__abc_16259_n9857), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n9858) );
  AND2X2 AND2X2_3618 ( .A(AES_CORE_DATAPATH__abc_16259_n9856), .B(AES_CORE_DATAPATH__abc_16259_n9858), .Y(AES_CORE_DATAPATH__abc_16259_n9859) );
  AND2X2 AND2X2_3619 ( .A(AES_CORE_DATAPATH__abc_16259_n9861), .B(AES_CORE_DATAPATH__abc_16259_n9862), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__0_) );
  AND2X2 AND2X2_362 ( .A(AES_CORE_DATAPATH__abc_16259_n2798_bF_buf1), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_3_), .Y(AES_CORE_DATAPATH__abc_16259_n2986) );
  AND2X2 AND2X2_3620 ( .A(AES_CORE_DATAPATH__abc_16259_n9865), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n9866) );
  AND2X2 AND2X2_3621 ( .A(AES_CORE_DATAPATH__abc_16259_n9864), .B(AES_CORE_DATAPATH__abc_16259_n9866), .Y(AES_CORE_DATAPATH__abc_16259_n9867) );
  AND2X2 AND2X2_3622 ( .A(AES_CORE_DATAPATH__abc_16259_n9869), .B(AES_CORE_DATAPATH__abc_16259_n9870), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__1_) );
  AND2X2 AND2X2_3623 ( .A(AES_CORE_DATAPATH__abc_16259_n9873), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n9874) );
  AND2X2 AND2X2_3624 ( .A(AES_CORE_DATAPATH__abc_16259_n9872), .B(AES_CORE_DATAPATH__abc_16259_n9874), .Y(AES_CORE_DATAPATH__abc_16259_n9875) );
  AND2X2 AND2X2_3625 ( .A(AES_CORE_DATAPATH__abc_16259_n9877), .B(AES_CORE_DATAPATH__abc_16259_n9878), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__2_) );
  AND2X2 AND2X2_3626 ( .A(AES_CORE_DATAPATH__abc_16259_n9881), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n9882) );
  AND2X2 AND2X2_3627 ( .A(AES_CORE_DATAPATH__abc_16259_n9880), .B(AES_CORE_DATAPATH__abc_16259_n9882), .Y(AES_CORE_DATAPATH__abc_16259_n9883) );
  AND2X2 AND2X2_3628 ( .A(AES_CORE_DATAPATH__abc_16259_n9885), .B(AES_CORE_DATAPATH__abc_16259_n9886), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__3_) );
  AND2X2 AND2X2_3629 ( .A(AES_CORE_DATAPATH__abc_16259_n9889), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n9890) );
  AND2X2 AND2X2_363 ( .A(AES_CORE_DATAPATH__abc_16259_n2984_1), .B(AES_CORE_DATAPATH__abc_16259_n2988), .Y(AES_CORE_DATAPATH__abc_16259_n2989) );
  AND2X2 AND2X2_3630 ( .A(AES_CORE_DATAPATH__abc_16259_n9888), .B(AES_CORE_DATAPATH__abc_16259_n9890), .Y(AES_CORE_DATAPATH__abc_16259_n9891) );
  AND2X2 AND2X2_3631 ( .A(AES_CORE_DATAPATH__abc_16259_n9893), .B(AES_CORE_DATAPATH__abc_16259_n9894), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__4_) );
  AND2X2 AND2X2_3632 ( .A(AES_CORE_DATAPATH__abc_16259_n9897), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n9898) );
  AND2X2 AND2X2_3633 ( .A(AES_CORE_DATAPATH__abc_16259_n9896), .B(AES_CORE_DATAPATH__abc_16259_n9898), .Y(AES_CORE_DATAPATH__abc_16259_n9899) );
  AND2X2 AND2X2_3634 ( .A(AES_CORE_DATAPATH__abc_16259_n9901), .B(AES_CORE_DATAPATH__abc_16259_n9902), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__5_) );
  AND2X2 AND2X2_3635 ( .A(AES_CORE_DATAPATH__abc_16259_n9905), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n9906) );
  AND2X2 AND2X2_3636 ( .A(AES_CORE_DATAPATH__abc_16259_n9904), .B(AES_CORE_DATAPATH__abc_16259_n9906), .Y(AES_CORE_DATAPATH__abc_16259_n9907) );
  AND2X2 AND2X2_3637 ( .A(AES_CORE_DATAPATH__abc_16259_n9909), .B(AES_CORE_DATAPATH__abc_16259_n9910), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__6_) );
  AND2X2 AND2X2_3638 ( .A(AES_CORE_DATAPATH__abc_16259_n9913), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n9914) );
  AND2X2 AND2X2_3639 ( .A(AES_CORE_DATAPATH__abc_16259_n9912), .B(AES_CORE_DATAPATH__abc_16259_n9914), .Y(AES_CORE_DATAPATH__abc_16259_n9915) );
  AND2X2 AND2X2_364 ( .A(AES_CORE_DATAPATH__abc_16259_n2989), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n2990) );
  AND2X2 AND2X2_3640 ( .A(AES_CORE_DATAPATH__abc_16259_n9917), .B(AES_CORE_DATAPATH__abc_16259_n9918), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__7_) );
  AND2X2 AND2X2_3641 ( .A(AES_CORE_DATAPATH__abc_16259_n9921), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf10), .Y(AES_CORE_DATAPATH__abc_16259_n9922) );
  AND2X2 AND2X2_3642 ( .A(AES_CORE_DATAPATH__abc_16259_n9920), .B(AES_CORE_DATAPATH__abc_16259_n9922), .Y(AES_CORE_DATAPATH__abc_16259_n9923) );
  AND2X2 AND2X2_3643 ( .A(AES_CORE_DATAPATH__abc_16259_n9925), .B(AES_CORE_DATAPATH__abc_16259_n9926), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__8_) );
  AND2X2 AND2X2_3644 ( .A(AES_CORE_DATAPATH__abc_16259_n9929), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf9), .Y(AES_CORE_DATAPATH__abc_16259_n9930) );
  AND2X2 AND2X2_3645 ( .A(AES_CORE_DATAPATH__abc_16259_n9928), .B(AES_CORE_DATAPATH__abc_16259_n9930), .Y(AES_CORE_DATAPATH__abc_16259_n9931) );
  AND2X2 AND2X2_3646 ( .A(AES_CORE_DATAPATH__abc_16259_n9933), .B(AES_CORE_DATAPATH__abc_16259_n9934), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__9_) );
  AND2X2 AND2X2_3647 ( .A(AES_CORE_DATAPATH__abc_16259_n8031), .B(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n9936) );
  AND2X2 AND2X2_3648 ( .A(AES_CORE_DATAPATH__abc_16259_n9938), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf8), .Y(AES_CORE_DATAPATH__abc_16259_n9939) );
  AND2X2 AND2X2_3649 ( .A(AES_CORE_DATAPATH__abc_16259_n9937), .B(AES_CORE_DATAPATH__abc_16259_n9939), .Y(AES_CORE_DATAPATH__abc_16259_n9940) );
  AND2X2 AND2X2_365 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf8), .B(AES_CORE_DATAPATH_col_3__3_), .Y(AES_CORE_DATAPATH__abc_16259_n2991) );
  AND2X2 AND2X2_3650 ( .A(AES_CORE_DATAPATH__abc_16259_n9942), .B(AES_CORE_DATAPATH__abc_16259_n9943), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__10_) );
  AND2X2 AND2X2_3651 ( .A(AES_CORE_DATAPATH__abc_16259_n8043), .B(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n9945) );
  AND2X2 AND2X2_3652 ( .A(AES_CORE_DATAPATH__abc_16259_n9947), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n9948) );
  AND2X2 AND2X2_3653 ( .A(AES_CORE_DATAPATH__abc_16259_n9946), .B(AES_CORE_DATAPATH__abc_16259_n9948), .Y(AES_CORE_DATAPATH__abc_16259_n9949) );
  AND2X2 AND2X2_3654 ( .A(AES_CORE_DATAPATH__abc_16259_n9951), .B(AES_CORE_DATAPATH__abc_16259_n9952), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__11_) );
  AND2X2 AND2X2_3655 ( .A(AES_CORE_DATAPATH__abc_16259_n9955), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n9956) );
  AND2X2 AND2X2_3656 ( .A(AES_CORE_DATAPATH__abc_16259_n9954), .B(AES_CORE_DATAPATH__abc_16259_n9956), .Y(AES_CORE_DATAPATH__abc_16259_n9957) );
  AND2X2 AND2X2_3657 ( .A(AES_CORE_DATAPATH__abc_16259_n9959), .B(AES_CORE_DATAPATH__abc_16259_n9960), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__12_) );
  AND2X2 AND2X2_3658 ( .A(AES_CORE_DATAPATH__abc_16259_n8061), .B(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n9962) );
  AND2X2 AND2X2_3659 ( .A(AES_CORE_DATAPATH__abc_16259_n9964), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n9965) );
  AND2X2 AND2X2_366 ( .A(AES_CORE_DATAPATH__abc_16259_n2994), .B(AES_CORE_DATAPATH__abc_16259_n2996_1), .Y(AES_CORE_DATAPATH__abc_16259_n2997) );
  AND2X2 AND2X2_3660 ( .A(AES_CORE_DATAPATH__abc_16259_n9963), .B(AES_CORE_DATAPATH__abc_16259_n9965), .Y(AES_CORE_DATAPATH__abc_16259_n9966) );
  AND2X2 AND2X2_3661 ( .A(AES_CORE_DATAPATH__abc_16259_n9968), .B(AES_CORE_DATAPATH__abc_16259_n9969), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__13_) );
  AND2X2 AND2X2_3662 ( .A(AES_CORE_DATAPATH__abc_16259_n9972), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n9973) );
  AND2X2 AND2X2_3663 ( .A(AES_CORE_DATAPATH__abc_16259_n9971), .B(AES_CORE_DATAPATH__abc_16259_n9973), .Y(AES_CORE_DATAPATH__abc_16259_n9974) );
  AND2X2 AND2X2_3664 ( .A(AES_CORE_DATAPATH__abc_16259_n9976), .B(AES_CORE_DATAPATH__abc_16259_n9977), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__14_) );
  AND2X2 AND2X2_3665 ( .A(AES_CORE_DATAPATH__abc_16259_n8080), .B(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf11), .Y(AES_CORE_DATAPATH__abc_16259_n9979) );
  AND2X2 AND2X2_3666 ( .A(AES_CORE_DATAPATH__abc_16259_n9981), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n9982) );
  AND2X2 AND2X2_3667 ( .A(AES_CORE_DATAPATH__abc_16259_n9980), .B(AES_CORE_DATAPATH__abc_16259_n9982), .Y(AES_CORE_DATAPATH__abc_16259_n9983) );
  AND2X2 AND2X2_3668 ( .A(AES_CORE_DATAPATH__abc_16259_n9985), .B(AES_CORE_DATAPATH__abc_16259_n9986), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__15_) );
  AND2X2 AND2X2_3669 ( .A(AES_CORE_DATAPATH__abc_16259_n9989), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n9990) );
  AND2X2 AND2X2_367 ( .A(AES_CORE_DATAPATH__abc_16259_n2782_bF_buf0), .B(AES_CORE_DATAPATH_col_3__4_), .Y(AES_CORE_DATAPATH__abc_16259_n2998_1) );
  AND2X2 AND2X2_3670 ( .A(AES_CORE_DATAPATH__abc_16259_n9988), .B(AES_CORE_DATAPATH__abc_16259_n9990), .Y(AES_CORE_DATAPATH__abc_16259_n9991) );
  AND2X2 AND2X2_3671 ( .A(AES_CORE_DATAPATH__abc_16259_n9993), .B(AES_CORE_DATAPATH__abc_16259_n9994), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__16_) );
  AND2X2 AND2X2_3672 ( .A(AES_CORE_DATAPATH__abc_16259_n8099), .B(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf8), .Y(AES_CORE_DATAPATH__abc_16259_n9996) );
  AND2X2 AND2X2_3673 ( .A(AES_CORE_DATAPATH__abc_16259_n9998), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n9999) );
  AND2X2 AND2X2_3674 ( .A(AES_CORE_DATAPATH__abc_16259_n9997), .B(AES_CORE_DATAPATH__abc_16259_n9999), .Y(AES_CORE_DATAPATH__abc_16259_n10000) );
  AND2X2 AND2X2_3675 ( .A(AES_CORE_DATAPATH__abc_16259_n10002), .B(AES_CORE_DATAPATH__abc_16259_n10003), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__17_) );
  AND2X2 AND2X2_3676 ( .A(AES_CORE_DATAPATH__abc_16259_n10006), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n10007) );
  AND2X2 AND2X2_3677 ( .A(AES_CORE_DATAPATH__abc_16259_n10005), .B(AES_CORE_DATAPATH__abc_16259_n10007), .Y(AES_CORE_DATAPATH__abc_16259_n10008) );
  AND2X2 AND2X2_3678 ( .A(AES_CORE_DATAPATH__abc_16259_n10010), .B(AES_CORE_DATAPATH__abc_16259_n10011), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__18_) );
  AND2X2 AND2X2_3679 ( .A(AES_CORE_DATAPATH__abc_16259_n10014), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf10), .Y(AES_CORE_DATAPATH__abc_16259_n10015) );
  AND2X2 AND2X2_368 ( .A(AES_CORE_DATAPATH__abc_16259_n2786_bF_buf0), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_68_), .Y(AES_CORE_DATAPATH__abc_16259_n2999) );
  AND2X2 AND2X2_3680 ( .A(AES_CORE_DATAPATH__abc_16259_n10013), .B(AES_CORE_DATAPATH__abc_16259_n10015), .Y(AES_CORE_DATAPATH__abc_16259_n10016) );
  AND2X2 AND2X2_3681 ( .A(AES_CORE_DATAPATH__abc_16259_n10018), .B(AES_CORE_DATAPATH__abc_16259_n10019), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__19_) );
  AND2X2 AND2X2_3682 ( .A(AES_CORE_DATAPATH__abc_16259_n10022), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf9), .Y(AES_CORE_DATAPATH__abc_16259_n10023) );
  AND2X2 AND2X2_3683 ( .A(AES_CORE_DATAPATH__abc_16259_n10021), .B(AES_CORE_DATAPATH__abc_16259_n10023), .Y(AES_CORE_DATAPATH__abc_16259_n10024) );
  AND2X2 AND2X2_3684 ( .A(AES_CORE_DATAPATH__abc_16259_n10026), .B(AES_CORE_DATAPATH__abc_16259_n10027), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__20_) );
  AND2X2 AND2X2_3685 ( .A(AES_CORE_DATAPATH__abc_16259_n8134), .B(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n10029) );
  AND2X2 AND2X2_3686 ( .A(AES_CORE_DATAPATH__abc_16259_n10031), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf8), .Y(AES_CORE_DATAPATH__abc_16259_n10032) );
  AND2X2 AND2X2_3687 ( .A(AES_CORE_DATAPATH__abc_16259_n10030), .B(AES_CORE_DATAPATH__abc_16259_n10032), .Y(AES_CORE_DATAPATH__abc_16259_n10033) );
  AND2X2 AND2X2_3688 ( .A(AES_CORE_DATAPATH__abc_16259_n10035), .B(AES_CORE_DATAPATH__abc_16259_n10036), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__21_) );
  AND2X2 AND2X2_3689 ( .A(AES_CORE_DATAPATH__abc_16259_n10039), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n10040) );
  AND2X2 AND2X2_369 ( .A(AES_CORE_DATAPATH__abc_16259_n2789_bF_buf0), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_36_), .Y(AES_CORE_DATAPATH__abc_16259_n3000) );
  AND2X2 AND2X2_3690 ( .A(AES_CORE_DATAPATH__abc_16259_n10038), .B(AES_CORE_DATAPATH__abc_16259_n10040), .Y(AES_CORE_DATAPATH__abc_16259_n10041) );
  AND2X2 AND2X2_3691 ( .A(AES_CORE_DATAPATH__abc_16259_n10043), .B(AES_CORE_DATAPATH__abc_16259_n10044), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__22_) );
  AND2X2 AND2X2_3692 ( .A(AES_CORE_DATAPATH__abc_16259_n10047), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n10048) );
  AND2X2 AND2X2_3693 ( .A(AES_CORE_DATAPATH__abc_16259_n10046), .B(AES_CORE_DATAPATH__abc_16259_n10048), .Y(AES_CORE_DATAPATH__abc_16259_n10049) );
  AND2X2 AND2X2_3694 ( .A(AES_CORE_DATAPATH__abc_16259_n10051), .B(AES_CORE_DATAPATH__abc_16259_n10052), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__23_) );
  AND2X2 AND2X2_3695 ( .A(AES_CORE_DATAPATH__abc_16259_n10055), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n10056) );
  AND2X2 AND2X2_3696 ( .A(AES_CORE_DATAPATH__abc_16259_n10054), .B(AES_CORE_DATAPATH__abc_16259_n10056), .Y(AES_CORE_DATAPATH__abc_16259_n10057) );
  AND2X2 AND2X2_3697 ( .A(AES_CORE_DATAPATH__abc_16259_n10059), .B(AES_CORE_DATAPATH__abc_16259_n10060), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__24_) );
  AND2X2 AND2X2_3698 ( .A(AES_CORE_DATAPATH__abc_16259_n10063), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n10064) );
  AND2X2 AND2X2_3699 ( .A(AES_CORE_DATAPATH__abc_16259_n10062), .B(AES_CORE_DATAPATH__abc_16259_n10064), .Y(AES_CORE_DATAPATH__abc_16259_n10065) );
  AND2X2 AND2X2_37 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n99_1), .B(AES_CORE_CONTROL_UNIT__abc_15841_n78), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n127) );
  AND2X2 AND2X2_370 ( .A(AES_CORE_DATAPATH__abc_16259_n3003_1), .B(AES_CORE_DATAPATH__abc_16259_n2997), .Y(AES_CORE_DATAPATH__abc_16259_n3004_1) );
  AND2X2 AND2X2_3700 ( .A(AES_CORE_DATAPATH__abc_16259_n10067), .B(AES_CORE_DATAPATH__abc_16259_n10068), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__25_) );
  AND2X2 AND2X2_3701 ( .A(AES_CORE_DATAPATH__abc_16259_n10071), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n10072) );
  AND2X2 AND2X2_3702 ( .A(AES_CORE_DATAPATH__abc_16259_n10070), .B(AES_CORE_DATAPATH__abc_16259_n10072), .Y(AES_CORE_DATAPATH__abc_16259_n10073) );
  AND2X2 AND2X2_3703 ( .A(AES_CORE_DATAPATH__abc_16259_n10075), .B(AES_CORE_DATAPATH__abc_16259_n10076), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__26_) );
  AND2X2 AND2X2_3704 ( .A(AES_CORE_DATAPATH__abc_16259_n10079), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n10080) );
  AND2X2 AND2X2_3705 ( .A(AES_CORE_DATAPATH__abc_16259_n10078), .B(AES_CORE_DATAPATH__abc_16259_n10080), .Y(AES_CORE_DATAPATH__abc_16259_n10081) );
  AND2X2 AND2X2_3706 ( .A(AES_CORE_DATAPATH__abc_16259_n10083), .B(AES_CORE_DATAPATH__abc_16259_n10084), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__27_) );
  AND2X2 AND2X2_3707 ( .A(AES_CORE_DATAPATH__abc_16259_n10087), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n10088) );
  AND2X2 AND2X2_3708 ( .A(AES_CORE_DATAPATH__abc_16259_n10086), .B(AES_CORE_DATAPATH__abc_16259_n10088), .Y(AES_CORE_DATAPATH__abc_16259_n10089) );
  AND2X2 AND2X2_3709 ( .A(AES_CORE_DATAPATH__abc_16259_n10091), .B(AES_CORE_DATAPATH__abc_16259_n10092), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__28_) );
  AND2X2 AND2X2_371 ( .A(AES_CORE_DATAPATH__abc_16259_n2837_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__4_), .Y(AES_CORE_DATAPATH__abc_16259_n3006) );
  AND2X2 AND2X2_3710 ( .A(AES_CORE_DATAPATH__abc_16259_n10095), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n10096) );
  AND2X2 AND2X2_3711 ( .A(AES_CORE_DATAPATH__abc_16259_n10094), .B(AES_CORE_DATAPATH__abc_16259_n10096), .Y(AES_CORE_DATAPATH__abc_16259_n10097) );
  AND2X2 AND2X2_3712 ( .A(AES_CORE_DATAPATH__abc_16259_n10099), .B(AES_CORE_DATAPATH__abc_16259_n10100), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__29_) );
  AND2X2 AND2X2_3713 ( .A(AES_CORE_DATAPATH__abc_16259_n10103), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf10), .Y(AES_CORE_DATAPATH__abc_16259_n10104) );
  AND2X2 AND2X2_3714 ( .A(AES_CORE_DATAPATH__abc_16259_n10102), .B(AES_CORE_DATAPATH__abc_16259_n10104), .Y(AES_CORE_DATAPATH__abc_16259_n10105) );
  AND2X2 AND2X2_3715 ( .A(AES_CORE_DATAPATH__abc_16259_n10107), .B(AES_CORE_DATAPATH__abc_16259_n10108), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__30_) );
  AND2X2 AND2X2_3716 ( .A(AES_CORE_DATAPATH__abc_16259_n10111), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf9), .Y(AES_CORE_DATAPATH__abc_16259_n10112) );
  AND2X2 AND2X2_3717 ( .A(AES_CORE_DATAPATH__abc_16259_n10110), .B(AES_CORE_DATAPATH__abc_16259_n10112), .Y(AES_CORE_DATAPATH__abc_16259_n10113) );
  AND2X2 AND2X2_3718 ( .A(AES_CORE_DATAPATH__abc_16259_n10115), .B(AES_CORE_DATAPATH__abc_16259_n10116), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__31_) );
  AND2X2 AND2X2_3719 ( .A(AES_CORE_DATAPATH__abc_16259_n10120), .B(AES_CORE_DATAPATH__abc_16259_n10118), .Y(AES_CORE_DATAPATH__0iv_1__31_0__0_) );
  AND2X2 AND2X2_372 ( .A(AES_CORE_DATAPATH__abc_16259_n2887_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__4_), .Y(AES_CORE_DATAPATH__abc_16259_n3008) );
  AND2X2 AND2X2_3720 ( .A(AES_CORE_DATAPATH__abc_16259_n10123), .B(AES_CORE_DATAPATH__abc_16259_n10122), .Y(AES_CORE_DATAPATH__0iv_1__31_0__1_) );
  AND2X2 AND2X2_3721 ( .A(AES_CORE_DATAPATH__abc_16259_n10126), .B(AES_CORE_DATAPATH__abc_16259_n10125), .Y(AES_CORE_DATAPATH__0iv_1__31_0__2_) );
  AND2X2 AND2X2_3722 ( .A(AES_CORE_DATAPATH__abc_16259_n10129), .B(AES_CORE_DATAPATH__abc_16259_n10128), .Y(AES_CORE_DATAPATH__0iv_1__31_0__3_) );
  AND2X2 AND2X2_3723 ( .A(AES_CORE_DATAPATH__abc_16259_n10132), .B(AES_CORE_DATAPATH__abc_16259_n10131), .Y(AES_CORE_DATAPATH__0iv_1__31_0__4_) );
  AND2X2 AND2X2_3724 ( .A(AES_CORE_DATAPATH__abc_16259_n10135), .B(AES_CORE_DATAPATH__abc_16259_n10134), .Y(AES_CORE_DATAPATH__0iv_1__31_0__5_) );
  AND2X2 AND2X2_3725 ( .A(AES_CORE_DATAPATH__abc_16259_n10138), .B(AES_CORE_DATAPATH__abc_16259_n10137), .Y(AES_CORE_DATAPATH__0iv_1__31_0__6_) );
  AND2X2 AND2X2_3726 ( .A(AES_CORE_DATAPATH__abc_16259_n10141), .B(AES_CORE_DATAPATH__abc_16259_n10140), .Y(AES_CORE_DATAPATH__0iv_1__31_0__7_) );
  AND2X2 AND2X2_3727 ( .A(AES_CORE_DATAPATH__abc_16259_n10144), .B(AES_CORE_DATAPATH__abc_16259_n10143), .Y(AES_CORE_DATAPATH__0iv_1__31_0__8_) );
  AND2X2 AND2X2_3728 ( .A(AES_CORE_DATAPATH__abc_16259_n10147), .B(AES_CORE_DATAPATH__abc_16259_n10146), .Y(AES_CORE_DATAPATH__0iv_1__31_0__9_) );
  AND2X2 AND2X2_3729 ( .A(AES_CORE_DATAPATH__abc_16259_n10150), .B(AES_CORE_DATAPATH__abc_16259_n10149), .Y(AES_CORE_DATAPATH__0iv_1__31_0__10_) );
  AND2X2 AND2X2_373 ( .A(AES_CORE_DATAPATH__abc_16259_n2830_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__4_), .Y(AES_CORE_DATAPATH__abc_16259_n3009_1) );
  AND2X2 AND2X2_3730 ( .A(AES_CORE_DATAPATH__abc_16259_n10153), .B(AES_CORE_DATAPATH__abc_16259_n10152), .Y(AES_CORE_DATAPATH__0iv_1__31_0__11_) );
  AND2X2 AND2X2_3731 ( .A(AES_CORE_DATAPATH__abc_16259_n10156), .B(AES_CORE_DATAPATH__abc_16259_n10155), .Y(AES_CORE_DATAPATH__0iv_1__31_0__12_) );
  AND2X2 AND2X2_3732 ( .A(AES_CORE_DATAPATH__abc_16259_n10159), .B(AES_CORE_DATAPATH__abc_16259_n10158), .Y(AES_CORE_DATAPATH__0iv_1__31_0__13_) );
  AND2X2 AND2X2_3733 ( .A(AES_CORE_DATAPATH__abc_16259_n10162), .B(AES_CORE_DATAPATH__abc_16259_n10161), .Y(AES_CORE_DATAPATH__0iv_1__31_0__14_) );
  AND2X2 AND2X2_3734 ( .A(AES_CORE_DATAPATH__abc_16259_n10165), .B(AES_CORE_DATAPATH__abc_16259_n10164), .Y(AES_CORE_DATAPATH__0iv_1__31_0__15_) );
  AND2X2 AND2X2_3735 ( .A(AES_CORE_DATAPATH__abc_16259_n10168), .B(AES_CORE_DATAPATH__abc_16259_n10167), .Y(AES_CORE_DATAPATH__0iv_1__31_0__16_) );
  AND2X2 AND2X2_3736 ( .A(AES_CORE_DATAPATH__abc_16259_n10171), .B(AES_CORE_DATAPATH__abc_16259_n10170), .Y(AES_CORE_DATAPATH__0iv_1__31_0__17_) );
  AND2X2 AND2X2_3737 ( .A(AES_CORE_DATAPATH__abc_16259_n10174), .B(AES_CORE_DATAPATH__abc_16259_n10173), .Y(AES_CORE_DATAPATH__0iv_1__31_0__18_) );
  AND2X2 AND2X2_3738 ( .A(AES_CORE_DATAPATH__abc_16259_n10177), .B(AES_CORE_DATAPATH__abc_16259_n10176), .Y(AES_CORE_DATAPATH__0iv_1__31_0__19_) );
  AND2X2 AND2X2_3739 ( .A(AES_CORE_DATAPATH__abc_16259_n10180), .B(AES_CORE_DATAPATH__abc_16259_n10179), .Y(AES_CORE_DATAPATH__0iv_1__31_0__20_) );
  AND2X2 AND2X2_374 ( .A(AES_CORE_DATAPATH__abc_16259_n3011_1), .B(AES_CORE_DATAPATH__abc_16259_n3012), .Y(_auto_iopadmap_cc_313_execute_26949_4_) );
  AND2X2 AND2X2_3740 ( .A(AES_CORE_DATAPATH__abc_16259_n10183), .B(AES_CORE_DATAPATH__abc_16259_n10182), .Y(AES_CORE_DATAPATH__0iv_1__31_0__21_) );
  AND2X2 AND2X2_3741 ( .A(AES_CORE_DATAPATH__abc_16259_n10186), .B(AES_CORE_DATAPATH__abc_16259_n10185), .Y(AES_CORE_DATAPATH__0iv_1__31_0__22_) );
  AND2X2 AND2X2_3742 ( .A(AES_CORE_DATAPATH__abc_16259_n10189), .B(AES_CORE_DATAPATH__abc_16259_n10188), .Y(AES_CORE_DATAPATH__0iv_1__31_0__23_) );
  AND2X2 AND2X2_3743 ( .A(AES_CORE_DATAPATH__abc_16259_n10192), .B(AES_CORE_DATAPATH__abc_16259_n10191), .Y(AES_CORE_DATAPATH__0iv_1__31_0__24_) );
  AND2X2 AND2X2_3744 ( .A(AES_CORE_DATAPATH__abc_16259_n10195), .B(AES_CORE_DATAPATH__abc_16259_n10194), .Y(AES_CORE_DATAPATH__0iv_1__31_0__25_) );
  AND2X2 AND2X2_3745 ( .A(AES_CORE_DATAPATH__abc_16259_n10198), .B(AES_CORE_DATAPATH__abc_16259_n10197), .Y(AES_CORE_DATAPATH__0iv_1__31_0__26_) );
  AND2X2 AND2X2_3746 ( .A(AES_CORE_DATAPATH__abc_16259_n10201), .B(AES_CORE_DATAPATH__abc_16259_n10200), .Y(AES_CORE_DATAPATH__0iv_1__31_0__27_) );
  AND2X2 AND2X2_3747 ( .A(AES_CORE_DATAPATH__abc_16259_n10204), .B(AES_CORE_DATAPATH__abc_16259_n10203), .Y(AES_CORE_DATAPATH__0iv_1__31_0__28_) );
  AND2X2 AND2X2_3748 ( .A(AES_CORE_DATAPATH__abc_16259_n10207), .B(AES_CORE_DATAPATH__abc_16259_n10206), .Y(AES_CORE_DATAPATH__0iv_1__31_0__29_) );
  AND2X2 AND2X2_3749 ( .A(AES_CORE_DATAPATH__abc_16259_n10210), .B(AES_CORE_DATAPATH__abc_16259_n10209), .Y(AES_CORE_DATAPATH__0iv_1__31_0__30_) );
  AND2X2 AND2X2_375 ( .A(AES_CORE_DATAPATH__abc_16259_n2855_bF_buf0), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_4_), .Y(AES_CORE_DATAPATH__abc_16259_n3015) );
  AND2X2 AND2X2_3750 ( .A(AES_CORE_DATAPATH__abc_16259_n10213), .B(AES_CORE_DATAPATH__abc_16259_n10212), .Y(AES_CORE_DATAPATH__0iv_1__31_0__31_) );
  AND2X2 AND2X2_3751 ( .A(AES_CORE_DATAPATH__abc_16259_n8494), .B(AES_CORE_DATAPATH_col_en_host_0_), .Y(AES_CORE_DATAPATH__abc_16259_n10215) );
  AND2X2 AND2X2_3752 ( .A(AES_CORE_DATAPATH__abc_16259_n8497), .B(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_0_), .Y(AES_CORE_DATAPATH__abc_16259_n10216) );
  AND2X2 AND2X2_3753 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf6), .B(AES_CORE_DATAPATH_bkp_1_0__0_), .Y(AES_CORE_DATAPATH__abc_16259_n10219) );
  AND2X2 AND2X2_3754 ( .A(AES_CORE_DATAPATH__abc_16259_n8225), .B(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n10220) );
  AND2X2 AND2X2_3755 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf5), .B(AES_CORE_DATAPATH_bkp_1_0__1_), .Y(AES_CORE_DATAPATH__abc_16259_n10222) );
  AND2X2 AND2X2_3756 ( .A(AES_CORE_DATAPATH__abc_16259_n8233), .B(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n10223) );
  AND2X2 AND2X2_3757 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf4), .B(AES_CORE_DATAPATH_bkp_1_0__2_), .Y(AES_CORE_DATAPATH__abc_16259_n10225) );
  AND2X2 AND2X2_3758 ( .A(AES_CORE_DATAPATH__abc_16259_n8241), .B(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n10226) );
  AND2X2 AND2X2_3759 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1_0__3_), .Y(AES_CORE_DATAPATH__abc_16259_n10228) );
  AND2X2 AND2X2_376 ( .A(AES_CORE_DATAPATH__abc_16259_n2857_bF_buf0), .B(AES_CORE_DATAPATH_MIX_COL_col_0__4_), .Y(AES_CORE_DATAPATH__abc_16259_n3016) );
  AND2X2 AND2X2_3760 ( .A(AES_CORE_DATAPATH__abc_16259_n8249), .B(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n10229) );
  AND2X2 AND2X2_3761 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf2), .B(AES_CORE_DATAPATH_bkp_1_0__4_), .Y(AES_CORE_DATAPATH__abc_16259_n10231) );
  AND2X2 AND2X2_3762 ( .A(AES_CORE_DATAPATH__abc_16259_n8257), .B(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n10232) );
  AND2X2 AND2X2_3763 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf1), .B(AES_CORE_DATAPATH_bkp_1_0__5_), .Y(AES_CORE_DATAPATH__abc_16259_n10234) );
  AND2X2 AND2X2_3764 ( .A(AES_CORE_DATAPATH__abc_16259_n8265), .B(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n10235) );
  AND2X2 AND2X2_3765 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf0), .B(AES_CORE_DATAPATH_bkp_1_0__6_), .Y(AES_CORE_DATAPATH__abc_16259_n10237) );
  AND2X2 AND2X2_3766 ( .A(AES_CORE_DATAPATH__abc_16259_n8273), .B(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n10238) );
  AND2X2 AND2X2_3767 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf6), .B(AES_CORE_DATAPATH_bkp_1_0__7_), .Y(AES_CORE_DATAPATH__abc_16259_n10240) );
  AND2X2 AND2X2_3768 ( .A(AES_CORE_DATAPATH__abc_16259_n8281), .B(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n10241) );
  AND2X2 AND2X2_3769 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf5), .B(AES_CORE_DATAPATH_bkp_1_0__8_), .Y(AES_CORE_DATAPATH__abc_16259_n10243) );
  AND2X2 AND2X2_377 ( .A(AES_CORE_DATAPATH__abc_16259_n3014), .B(AES_CORE_DATAPATH__abc_16259_n3018), .Y(AES_CORE_DATAPATH__abc_16259_n3019) );
  AND2X2 AND2X2_3770 ( .A(AES_CORE_DATAPATH__abc_16259_n8289), .B(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n10244) );
  AND2X2 AND2X2_3771 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf4), .B(AES_CORE_DATAPATH_bkp_1_0__9_), .Y(AES_CORE_DATAPATH__abc_16259_n10246) );
  AND2X2 AND2X2_3772 ( .A(AES_CORE_DATAPATH__abc_16259_n8297), .B(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n10247) );
  AND2X2 AND2X2_3773 ( .A(AES_CORE_DATAPATH__abc_16259_n8306), .B(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n10249) );
  AND2X2 AND2X2_3774 ( .A(AES_CORE_DATAPATH__abc_16259_n10250), .B(AES_CORE_DATAPATH__abc_16259_n10251), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__10_) );
  AND2X2 AND2X2_3775 ( .A(AES_CORE_DATAPATH__abc_16259_n8317), .B(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n10253) );
  AND2X2 AND2X2_3776 ( .A(AES_CORE_DATAPATH__abc_16259_n10254), .B(AES_CORE_DATAPATH__abc_16259_n10255), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__11_) );
  AND2X2 AND2X2_3777 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1_0__12_), .Y(AES_CORE_DATAPATH__abc_16259_n10257) );
  AND2X2 AND2X2_3778 ( .A(AES_CORE_DATAPATH__abc_16259_n8327), .B(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n10258) );
  AND2X2 AND2X2_3779 ( .A(AES_CORE_DATAPATH__abc_16259_n8336), .B(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n10260) );
  AND2X2 AND2X2_378 ( .A(_auto_iopadmap_cc_313_execute_26949_4_), .B(AES_CORE_DATAPATH__abc_16259_n3019), .Y(AES_CORE_DATAPATH__abc_16259_n3022) );
  AND2X2 AND2X2_3780 ( .A(AES_CORE_DATAPATH__abc_16259_n10261), .B(AES_CORE_DATAPATH__abc_16259_n10262), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__13_) );
  AND2X2 AND2X2_3781 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf2), .B(AES_CORE_DATAPATH_bkp_1_0__14_), .Y(AES_CORE_DATAPATH__abc_16259_n10264) );
  AND2X2 AND2X2_3782 ( .A(AES_CORE_DATAPATH__abc_16259_n8346), .B(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n10265) );
  AND2X2 AND2X2_3783 ( .A(AES_CORE_DATAPATH__abc_16259_n8355), .B(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n10267) );
  AND2X2 AND2X2_3784 ( .A(AES_CORE_DATAPATH__abc_16259_n10268), .B(AES_CORE_DATAPATH__abc_16259_n10269), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__15_) );
  AND2X2 AND2X2_3785 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf1), .B(AES_CORE_DATAPATH_bkp_1_0__16_), .Y(AES_CORE_DATAPATH__abc_16259_n10271) );
  AND2X2 AND2X2_3786 ( .A(AES_CORE_DATAPATH__abc_16259_n8365), .B(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n10272) );
  AND2X2 AND2X2_3787 ( .A(AES_CORE_DATAPATH__abc_16259_n8374), .B(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n10274) );
  AND2X2 AND2X2_3788 ( .A(AES_CORE_DATAPATH__abc_16259_n10275), .B(AES_CORE_DATAPATH__abc_16259_n10276), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__17_) );
  AND2X2 AND2X2_3789 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf0), .B(AES_CORE_DATAPATH_bkp_1_0__18_), .Y(AES_CORE_DATAPATH__abc_16259_n10278) );
  AND2X2 AND2X2_379 ( .A(AES_CORE_DATAPATH_last_round_pp2_bF_buf4), .B(AES_CORE_DATAPATH_MIX_COL_col_0__4_), .Y(AES_CORE_DATAPATH__abc_16259_n3025_1) );
  AND2X2 AND2X2_3790 ( .A(AES_CORE_DATAPATH__abc_16259_n8384), .B(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n10279) );
  AND2X2 AND2X2_3791 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf6), .B(AES_CORE_DATAPATH_bkp_1_0__19_), .Y(AES_CORE_DATAPATH__abc_16259_n10281) );
  AND2X2 AND2X2_3792 ( .A(AES_CORE_DATAPATH__abc_16259_n8392), .B(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n10282) );
  AND2X2 AND2X2_3793 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf5), .B(AES_CORE_DATAPATH_bkp_1_0__20_), .Y(AES_CORE_DATAPATH__abc_16259_n10284) );
  AND2X2 AND2X2_3794 ( .A(AES_CORE_DATAPATH__abc_16259_n8400), .B(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n10285) );
  AND2X2 AND2X2_3795 ( .A(AES_CORE_DATAPATH__abc_16259_n8409), .B(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n10287) );
  AND2X2 AND2X2_3796 ( .A(AES_CORE_DATAPATH__abc_16259_n10288), .B(AES_CORE_DATAPATH__abc_16259_n10289), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__21_) );
  AND2X2 AND2X2_3797 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf4), .B(AES_CORE_DATAPATH_bkp_1_0__22_), .Y(AES_CORE_DATAPATH__abc_16259_n10291) );
  AND2X2 AND2X2_3798 ( .A(AES_CORE_DATAPATH__abc_16259_n8419), .B(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n10292) );
  AND2X2 AND2X2_3799 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1_0__23_), .Y(AES_CORE_DATAPATH__abc_16259_n10294) );
  AND2X2 AND2X2_38 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n107), .B(AES_CORE_CONTROL_UNIT_state_4_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n128) );
  AND2X2 AND2X2_380 ( .A(AES_CORE_DATAPATH__abc_16259_n2798_bF_buf0), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_4_), .Y(AES_CORE_DATAPATH__abc_16259_n3026) );
  AND2X2 AND2X2_3800 ( .A(AES_CORE_DATAPATH__abc_16259_n8427), .B(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n10295) );
  AND2X2 AND2X2_3801 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf2), .B(AES_CORE_DATAPATH_bkp_1_0__24_), .Y(AES_CORE_DATAPATH__abc_16259_n10297) );
  AND2X2 AND2X2_3802 ( .A(AES_CORE_DATAPATH__abc_16259_n8435), .B(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n10298) );
  AND2X2 AND2X2_3803 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf1), .B(AES_CORE_DATAPATH_bkp_1_0__25_), .Y(AES_CORE_DATAPATH__abc_16259_n10300) );
  AND2X2 AND2X2_3804 ( .A(AES_CORE_DATAPATH__abc_16259_n8443), .B(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n10301) );
  AND2X2 AND2X2_3805 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf0), .B(AES_CORE_DATAPATH_bkp_1_0__26_), .Y(AES_CORE_DATAPATH__abc_16259_n10303) );
  AND2X2 AND2X2_3806 ( .A(AES_CORE_DATAPATH__abc_16259_n8451), .B(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n10304) );
  AND2X2 AND2X2_3807 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf6), .B(AES_CORE_DATAPATH_bkp_1_0__27_), .Y(AES_CORE_DATAPATH__abc_16259_n10306) );
  AND2X2 AND2X2_3808 ( .A(AES_CORE_DATAPATH__abc_16259_n8459), .B(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n10307) );
  AND2X2 AND2X2_3809 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf5), .B(AES_CORE_DATAPATH_bkp_1_0__28_), .Y(AES_CORE_DATAPATH__abc_16259_n10309) );
  AND2X2 AND2X2_381 ( .A(AES_CORE_DATAPATH__abc_16259_n3024), .B(AES_CORE_DATAPATH__abc_16259_n3028), .Y(AES_CORE_DATAPATH__abc_16259_n3029) );
  AND2X2 AND2X2_3810 ( .A(AES_CORE_DATAPATH__abc_16259_n8467), .B(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n10310) );
  AND2X2 AND2X2_3811 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf4), .B(AES_CORE_DATAPATH_bkp_1_0__29_), .Y(AES_CORE_DATAPATH__abc_16259_n10312) );
  AND2X2 AND2X2_3812 ( .A(AES_CORE_DATAPATH__abc_16259_n8475), .B(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n10313) );
  AND2X2 AND2X2_3813 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1_0__30_), .Y(AES_CORE_DATAPATH__abc_16259_n10315) );
  AND2X2 AND2X2_3814 ( .A(AES_CORE_DATAPATH__abc_16259_n8483), .B(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n10316) );
  AND2X2 AND2X2_3815 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf2), .B(AES_CORE_DATAPATH_bkp_1_0__31_), .Y(AES_CORE_DATAPATH__abc_16259_n10318) );
  AND2X2 AND2X2_3816 ( .A(AES_CORE_DATAPATH__abc_16259_n8491), .B(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n10319) );
  AND2X2 AND2X2_3817 ( .A(AES_CORE_DATAPATH__abc_16259_n10322), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf8), .Y(AES_CORE_DATAPATH__abc_16259_n10323) );
  AND2X2 AND2X2_3818 ( .A(AES_CORE_DATAPATH__abc_16259_n10321), .B(AES_CORE_DATAPATH__abc_16259_n10323), .Y(AES_CORE_DATAPATH__abc_16259_n10324) );
  AND2X2 AND2X2_3819 ( .A(AES_CORE_DATAPATH__abc_16259_n10326), .B(AES_CORE_DATAPATH__abc_16259_n10327), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__0_) );
  AND2X2 AND2X2_382 ( .A(AES_CORE_DATAPATH__abc_16259_n3029), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n3030) );
  AND2X2 AND2X2_3820 ( .A(AES_CORE_DATAPATH__abc_16259_n10330), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n10331) );
  AND2X2 AND2X2_3821 ( .A(AES_CORE_DATAPATH__abc_16259_n10329), .B(AES_CORE_DATAPATH__abc_16259_n10331), .Y(AES_CORE_DATAPATH__abc_16259_n10332) );
  AND2X2 AND2X2_3822 ( .A(AES_CORE_DATAPATH__abc_16259_n10334), .B(AES_CORE_DATAPATH__abc_16259_n10335), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__1_) );
  AND2X2 AND2X2_3823 ( .A(AES_CORE_DATAPATH__abc_16259_n10338), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n10339) );
  AND2X2 AND2X2_3824 ( .A(AES_CORE_DATAPATH__abc_16259_n10337), .B(AES_CORE_DATAPATH__abc_16259_n10339), .Y(AES_CORE_DATAPATH__abc_16259_n10340) );
  AND2X2 AND2X2_3825 ( .A(AES_CORE_DATAPATH__abc_16259_n10342), .B(AES_CORE_DATAPATH__abc_16259_n10343), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__2_) );
  AND2X2 AND2X2_3826 ( .A(AES_CORE_DATAPATH__abc_16259_n10346), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n10347) );
  AND2X2 AND2X2_3827 ( .A(AES_CORE_DATAPATH__abc_16259_n10345), .B(AES_CORE_DATAPATH__abc_16259_n10347), .Y(AES_CORE_DATAPATH__abc_16259_n10348) );
  AND2X2 AND2X2_3828 ( .A(AES_CORE_DATAPATH__abc_16259_n10350), .B(AES_CORE_DATAPATH__abc_16259_n10351), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__3_) );
  AND2X2 AND2X2_3829 ( .A(AES_CORE_DATAPATH__abc_16259_n10354), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n10355) );
  AND2X2 AND2X2_383 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf7), .B(AES_CORE_DATAPATH_col_3__4_), .Y(AES_CORE_DATAPATH__abc_16259_n3031) );
  AND2X2 AND2X2_3830 ( .A(AES_CORE_DATAPATH__abc_16259_n10353), .B(AES_CORE_DATAPATH__abc_16259_n10355), .Y(AES_CORE_DATAPATH__abc_16259_n10356) );
  AND2X2 AND2X2_3831 ( .A(AES_CORE_DATAPATH__abc_16259_n10358), .B(AES_CORE_DATAPATH__abc_16259_n10359), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__4_) );
  AND2X2 AND2X2_3832 ( .A(AES_CORE_DATAPATH__abc_16259_n10362), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n10363) );
  AND2X2 AND2X2_3833 ( .A(AES_CORE_DATAPATH__abc_16259_n10361), .B(AES_CORE_DATAPATH__abc_16259_n10363), .Y(AES_CORE_DATAPATH__abc_16259_n10364) );
  AND2X2 AND2X2_3834 ( .A(AES_CORE_DATAPATH__abc_16259_n10366), .B(AES_CORE_DATAPATH__abc_16259_n10367), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__5_) );
  AND2X2 AND2X2_3835 ( .A(AES_CORE_DATAPATH__abc_16259_n10370), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n10371) );
  AND2X2 AND2X2_3836 ( .A(AES_CORE_DATAPATH__abc_16259_n10369), .B(AES_CORE_DATAPATH__abc_16259_n10371), .Y(AES_CORE_DATAPATH__abc_16259_n10372) );
  AND2X2 AND2X2_3837 ( .A(AES_CORE_DATAPATH__abc_16259_n10374), .B(AES_CORE_DATAPATH__abc_16259_n10375), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__6_) );
  AND2X2 AND2X2_3838 ( .A(AES_CORE_DATAPATH__abc_16259_n10378), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n10379) );
  AND2X2 AND2X2_3839 ( .A(AES_CORE_DATAPATH__abc_16259_n10377), .B(AES_CORE_DATAPATH__abc_16259_n10379), .Y(AES_CORE_DATAPATH__abc_16259_n10380) );
  AND2X2 AND2X2_384 ( .A(AES_CORE_DATAPATH__abc_16259_n3034), .B(AES_CORE_DATAPATH__abc_16259_n3036_1), .Y(AES_CORE_DATAPATH__abc_16259_n3037) );
  AND2X2 AND2X2_3840 ( .A(AES_CORE_DATAPATH__abc_16259_n10382), .B(AES_CORE_DATAPATH__abc_16259_n10383), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__7_) );
  AND2X2 AND2X2_3841 ( .A(AES_CORE_DATAPATH__abc_16259_n10386), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n10387) );
  AND2X2 AND2X2_3842 ( .A(AES_CORE_DATAPATH__abc_16259_n10385), .B(AES_CORE_DATAPATH__abc_16259_n10387), .Y(AES_CORE_DATAPATH__abc_16259_n10388) );
  AND2X2 AND2X2_3843 ( .A(AES_CORE_DATAPATH__abc_16259_n10390), .B(AES_CORE_DATAPATH__abc_16259_n10391), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__8_) );
  AND2X2 AND2X2_3844 ( .A(AES_CORE_DATAPATH__abc_16259_n10394), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf10), .Y(AES_CORE_DATAPATH__abc_16259_n10395) );
  AND2X2 AND2X2_3845 ( .A(AES_CORE_DATAPATH__abc_16259_n10393), .B(AES_CORE_DATAPATH__abc_16259_n10395), .Y(AES_CORE_DATAPATH__abc_16259_n10396) );
  AND2X2 AND2X2_3846 ( .A(AES_CORE_DATAPATH__abc_16259_n10398), .B(AES_CORE_DATAPATH__abc_16259_n10399), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__9_) );
  AND2X2 AND2X2_3847 ( .A(AES_CORE_DATAPATH__abc_16259_n8306), .B(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n10401) );
  AND2X2 AND2X2_3848 ( .A(AES_CORE_DATAPATH__abc_16259_n10403), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf9), .Y(AES_CORE_DATAPATH__abc_16259_n10404) );
  AND2X2 AND2X2_3849 ( .A(AES_CORE_DATAPATH__abc_16259_n10402), .B(AES_CORE_DATAPATH__abc_16259_n10404), .Y(AES_CORE_DATAPATH__abc_16259_n10405) );
  AND2X2 AND2X2_385 ( .A(AES_CORE_DATAPATH__abc_16259_n2782_bF_buf4), .B(AES_CORE_DATAPATH_col_3__5_), .Y(AES_CORE_DATAPATH__abc_16259_n3038_1) );
  AND2X2 AND2X2_3850 ( .A(AES_CORE_DATAPATH__abc_16259_n10407), .B(AES_CORE_DATAPATH__abc_16259_n10408), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__10_) );
  AND2X2 AND2X2_3851 ( .A(AES_CORE_DATAPATH__abc_16259_n8317), .B(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n10410) );
  AND2X2 AND2X2_3852 ( .A(AES_CORE_DATAPATH__abc_16259_n10412), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf8), .Y(AES_CORE_DATAPATH__abc_16259_n10413) );
  AND2X2 AND2X2_3853 ( .A(AES_CORE_DATAPATH__abc_16259_n10411), .B(AES_CORE_DATAPATH__abc_16259_n10413), .Y(AES_CORE_DATAPATH__abc_16259_n10414) );
  AND2X2 AND2X2_3854 ( .A(AES_CORE_DATAPATH__abc_16259_n10416), .B(AES_CORE_DATAPATH__abc_16259_n10417), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__11_) );
  AND2X2 AND2X2_3855 ( .A(AES_CORE_DATAPATH__abc_16259_n10420), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n10421) );
  AND2X2 AND2X2_3856 ( .A(AES_CORE_DATAPATH__abc_16259_n10419), .B(AES_CORE_DATAPATH__abc_16259_n10421), .Y(AES_CORE_DATAPATH__abc_16259_n10422) );
  AND2X2 AND2X2_3857 ( .A(AES_CORE_DATAPATH__abc_16259_n10424), .B(AES_CORE_DATAPATH__abc_16259_n10425), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__12_) );
  AND2X2 AND2X2_3858 ( .A(AES_CORE_DATAPATH__abc_16259_n8336), .B(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n10427) );
  AND2X2 AND2X2_3859 ( .A(AES_CORE_DATAPATH__abc_16259_n10429), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n10430) );
  AND2X2 AND2X2_386 ( .A(AES_CORE_DATAPATH__abc_16259_n2786_bF_buf4), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_69_), .Y(AES_CORE_DATAPATH__abc_16259_n3039) );
  AND2X2 AND2X2_3860 ( .A(AES_CORE_DATAPATH__abc_16259_n10428), .B(AES_CORE_DATAPATH__abc_16259_n10430), .Y(AES_CORE_DATAPATH__abc_16259_n10431) );
  AND2X2 AND2X2_3861 ( .A(AES_CORE_DATAPATH__abc_16259_n10433), .B(AES_CORE_DATAPATH__abc_16259_n10434), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__13_) );
  AND2X2 AND2X2_3862 ( .A(AES_CORE_DATAPATH__abc_16259_n10437), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n10438) );
  AND2X2 AND2X2_3863 ( .A(AES_CORE_DATAPATH__abc_16259_n10436), .B(AES_CORE_DATAPATH__abc_16259_n10438), .Y(AES_CORE_DATAPATH__abc_16259_n10439) );
  AND2X2 AND2X2_3864 ( .A(AES_CORE_DATAPATH__abc_16259_n10441), .B(AES_CORE_DATAPATH__abc_16259_n10442), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__14_) );
  AND2X2 AND2X2_3865 ( .A(AES_CORE_DATAPATH__abc_16259_n8355), .B(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf9), .Y(AES_CORE_DATAPATH__abc_16259_n10444) );
  AND2X2 AND2X2_3866 ( .A(AES_CORE_DATAPATH__abc_16259_n10446), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n10447) );
  AND2X2 AND2X2_3867 ( .A(AES_CORE_DATAPATH__abc_16259_n10445), .B(AES_CORE_DATAPATH__abc_16259_n10447), .Y(AES_CORE_DATAPATH__abc_16259_n10448) );
  AND2X2 AND2X2_3868 ( .A(AES_CORE_DATAPATH__abc_16259_n10450), .B(AES_CORE_DATAPATH__abc_16259_n10451), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__15_) );
  AND2X2 AND2X2_3869 ( .A(AES_CORE_DATAPATH__abc_16259_n10454), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n10455) );
  AND2X2 AND2X2_387 ( .A(AES_CORE_DATAPATH__abc_16259_n2789_bF_buf4), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_37_), .Y(AES_CORE_DATAPATH__abc_16259_n3040_1) );
  AND2X2 AND2X2_3870 ( .A(AES_CORE_DATAPATH__abc_16259_n10453), .B(AES_CORE_DATAPATH__abc_16259_n10455), .Y(AES_CORE_DATAPATH__abc_16259_n10456) );
  AND2X2 AND2X2_3871 ( .A(AES_CORE_DATAPATH__abc_16259_n10458), .B(AES_CORE_DATAPATH__abc_16259_n10459), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__16_) );
  AND2X2 AND2X2_3872 ( .A(AES_CORE_DATAPATH__abc_16259_n8374), .B(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n10461) );
  AND2X2 AND2X2_3873 ( .A(AES_CORE_DATAPATH__abc_16259_n10463), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n10464) );
  AND2X2 AND2X2_3874 ( .A(AES_CORE_DATAPATH__abc_16259_n10462), .B(AES_CORE_DATAPATH__abc_16259_n10464), .Y(AES_CORE_DATAPATH__abc_16259_n10465) );
  AND2X2 AND2X2_3875 ( .A(AES_CORE_DATAPATH__abc_16259_n10467), .B(AES_CORE_DATAPATH__abc_16259_n10468), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__17_) );
  AND2X2 AND2X2_3876 ( .A(AES_CORE_DATAPATH__abc_16259_n10471), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n10472) );
  AND2X2 AND2X2_3877 ( .A(AES_CORE_DATAPATH__abc_16259_n10470), .B(AES_CORE_DATAPATH__abc_16259_n10472), .Y(AES_CORE_DATAPATH__abc_16259_n10473) );
  AND2X2 AND2X2_3878 ( .A(AES_CORE_DATAPATH__abc_16259_n10475), .B(AES_CORE_DATAPATH__abc_16259_n10476), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__18_) );
  AND2X2 AND2X2_3879 ( .A(AES_CORE_DATAPATH__abc_16259_n10479), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n10480) );
  AND2X2 AND2X2_388 ( .A(AES_CORE_DATAPATH__abc_16259_n3043), .B(AES_CORE_DATAPATH__abc_16259_n3037), .Y(AES_CORE_DATAPATH__abc_16259_n3044) );
  AND2X2 AND2X2_3880 ( .A(AES_CORE_DATAPATH__abc_16259_n10478), .B(AES_CORE_DATAPATH__abc_16259_n10480), .Y(AES_CORE_DATAPATH__abc_16259_n10481) );
  AND2X2 AND2X2_3881 ( .A(AES_CORE_DATAPATH__abc_16259_n10483), .B(AES_CORE_DATAPATH__abc_16259_n10484), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__19_) );
  AND2X2 AND2X2_3882 ( .A(AES_CORE_DATAPATH__abc_16259_n10487), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf10), .Y(AES_CORE_DATAPATH__abc_16259_n10488) );
  AND2X2 AND2X2_3883 ( .A(AES_CORE_DATAPATH__abc_16259_n10486), .B(AES_CORE_DATAPATH__abc_16259_n10488), .Y(AES_CORE_DATAPATH__abc_16259_n10489) );
  AND2X2 AND2X2_3884 ( .A(AES_CORE_DATAPATH__abc_16259_n10491), .B(AES_CORE_DATAPATH__abc_16259_n10492), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__20_) );
  AND2X2 AND2X2_3885 ( .A(AES_CORE_DATAPATH__abc_16259_n8409), .B(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n10494) );
  AND2X2 AND2X2_3886 ( .A(AES_CORE_DATAPATH__abc_16259_n10496), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf9), .Y(AES_CORE_DATAPATH__abc_16259_n10497) );
  AND2X2 AND2X2_3887 ( .A(AES_CORE_DATAPATH__abc_16259_n10495), .B(AES_CORE_DATAPATH__abc_16259_n10497), .Y(AES_CORE_DATAPATH__abc_16259_n10498) );
  AND2X2 AND2X2_3888 ( .A(AES_CORE_DATAPATH__abc_16259_n10500), .B(AES_CORE_DATAPATH__abc_16259_n10501), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__21_) );
  AND2X2 AND2X2_3889 ( .A(AES_CORE_DATAPATH__abc_16259_n10504), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf8), .Y(AES_CORE_DATAPATH__abc_16259_n10505) );
  AND2X2 AND2X2_389 ( .A(AES_CORE_DATAPATH__abc_16259_n2837_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__5_), .Y(AES_CORE_DATAPATH__abc_16259_n3046) );
  AND2X2 AND2X2_3890 ( .A(AES_CORE_DATAPATH__abc_16259_n10503), .B(AES_CORE_DATAPATH__abc_16259_n10505), .Y(AES_CORE_DATAPATH__abc_16259_n10506) );
  AND2X2 AND2X2_3891 ( .A(AES_CORE_DATAPATH__abc_16259_n10508), .B(AES_CORE_DATAPATH__abc_16259_n10509), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__22_) );
  AND2X2 AND2X2_3892 ( .A(AES_CORE_DATAPATH__abc_16259_n10512), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n10513) );
  AND2X2 AND2X2_3893 ( .A(AES_CORE_DATAPATH__abc_16259_n10511), .B(AES_CORE_DATAPATH__abc_16259_n10513), .Y(AES_CORE_DATAPATH__abc_16259_n10514) );
  AND2X2 AND2X2_3894 ( .A(AES_CORE_DATAPATH__abc_16259_n10516), .B(AES_CORE_DATAPATH__abc_16259_n10517), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__23_) );
  AND2X2 AND2X2_3895 ( .A(AES_CORE_DATAPATH__abc_16259_n10520), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n10521) );
  AND2X2 AND2X2_3896 ( .A(AES_CORE_DATAPATH__abc_16259_n10519), .B(AES_CORE_DATAPATH__abc_16259_n10521), .Y(AES_CORE_DATAPATH__abc_16259_n10522) );
  AND2X2 AND2X2_3897 ( .A(AES_CORE_DATAPATH__abc_16259_n10524), .B(AES_CORE_DATAPATH__abc_16259_n10525), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__24_) );
  AND2X2 AND2X2_3898 ( .A(AES_CORE_DATAPATH__abc_16259_n10528), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n10529) );
  AND2X2 AND2X2_3899 ( .A(AES_CORE_DATAPATH__abc_16259_n10527), .B(AES_CORE_DATAPATH__abc_16259_n10529), .Y(AES_CORE_DATAPATH__abc_16259_n10530) );
  AND2X2 AND2X2_39 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n131), .B(AES_CORE_CONTROL_UNIT_state_0_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n132) );
  AND2X2 AND2X2_390 ( .A(AES_CORE_DATAPATH__abc_16259_n2887_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__5_), .Y(AES_CORE_DATAPATH__abc_16259_n3048) );
  AND2X2 AND2X2_3900 ( .A(AES_CORE_DATAPATH__abc_16259_n10532), .B(AES_CORE_DATAPATH__abc_16259_n10533), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__25_) );
  AND2X2 AND2X2_3901 ( .A(AES_CORE_DATAPATH__abc_16259_n10536), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n10537) );
  AND2X2 AND2X2_3902 ( .A(AES_CORE_DATAPATH__abc_16259_n10535), .B(AES_CORE_DATAPATH__abc_16259_n10537), .Y(AES_CORE_DATAPATH__abc_16259_n10538) );
  AND2X2 AND2X2_3903 ( .A(AES_CORE_DATAPATH__abc_16259_n10540), .B(AES_CORE_DATAPATH__abc_16259_n10541), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__26_) );
  AND2X2 AND2X2_3904 ( .A(AES_CORE_DATAPATH__abc_16259_n10544), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n10545) );
  AND2X2 AND2X2_3905 ( .A(AES_CORE_DATAPATH__abc_16259_n10543), .B(AES_CORE_DATAPATH__abc_16259_n10545), .Y(AES_CORE_DATAPATH__abc_16259_n10546) );
  AND2X2 AND2X2_3906 ( .A(AES_CORE_DATAPATH__abc_16259_n10548), .B(AES_CORE_DATAPATH__abc_16259_n10549), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__27_) );
  AND2X2 AND2X2_3907 ( .A(AES_CORE_DATAPATH__abc_16259_n10552), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n10553) );
  AND2X2 AND2X2_3908 ( .A(AES_CORE_DATAPATH__abc_16259_n10551), .B(AES_CORE_DATAPATH__abc_16259_n10553), .Y(AES_CORE_DATAPATH__abc_16259_n10554) );
  AND2X2 AND2X2_3909 ( .A(AES_CORE_DATAPATH__abc_16259_n10556), .B(AES_CORE_DATAPATH__abc_16259_n10557), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__28_) );
  AND2X2 AND2X2_391 ( .A(AES_CORE_DATAPATH__abc_16259_n2830_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__5_), .Y(AES_CORE_DATAPATH__abc_16259_n3049) );
  AND2X2 AND2X2_3910 ( .A(AES_CORE_DATAPATH__abc_16259_n10560), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n10561) );
  AND2X2 AND2X2_3911 ( .A(AES_CORE_DATAPATH__abc_16259_n10559), .B(AES_CORE_DATAPATH__abc_16259_n10561), .Y(AES_CORE_DATAPATH__abc_16259_n10562) );
  AND2X2 AND2X2_3912 ( .A(AES_CORE_DATAPATH__abc_16259_n10564), .B(AES_CORE_DATAPATH__abc_16259_n10565), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__29_) );
  AND2X2 AND2X2_3913 ( .A(AES_CORE_DATAPATH__abc_16259_n10568), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n10569) );
  AND2X2 AND2X2_3914 ( .A(AES_CORE_DATAPATH__abc_16259_n10567), .B(AES_CORE_DATAPATH__abc_16259_n10569), .Y(AES_CORE_DATAPATH__abc_16259_n10570) );
  AND2X2 AND2X2_3915 ( .A(AES_CORE_DATAPATH__abc_16259_n10572), .B(AES_CORE_DATAPATH__abc_16259_n10573), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__30_) );
  AND2X2 AND2X2_3916 ( .A(AES_CORE_DATAPATH__abc_16259_n10576), .B(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf10), .Y(AES_CORE_DATAPATH__abc_16259_n10577) );
  AND2X2 AND2X2_3917 ( .A(AES_CORE_DATAPATH__abc_16259_n10575), .B(AES_CORE_DATAPATH__abc_16259_n10577), .Y(AES_CORE_DATAPATH__abc_16259_n10578) );
  AND2X2 AND2X2_3918 ( .A(AES_CORE_DATAPATH__abc_16259_n10580), .B(AES_CORE_DATAPATH__abc_16259_n10581), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__31_) );
  AND2X2 AND2X2_3919 ( .A(AES_CORE_DATAPATH__abc_16259_n10585), .B(AES_CORE_DATAPATH__abc_16259_n10583), .Y(AES_CORE_DATAPATH__0iv_0__31_0__0_) );
  AND2X2 AND2X2_392 ( .A(AES_CORE_DATAPATH__abc_16259_n3051), .B(AES_CORE_DATAPATH__abc_16259_n3052), .Y(_auto_iopadmap_cc_313_execute_26949_5_) );
  AND2X2 AND2X2_3920 ( .A(AES_CORE_DATAPATH__abc_16259_n10588), .B(AES_CORE_DATAPATH__abc_16259_n10587), .Y(AES_CORE_DATAPATH__0iv_0__31_0__1_) );
  AND2X2 AND2X2_3921 ( .A(AES_CORE_DATAPATH__abc_16259_n10591), .B(AES_CORE_DATAPATH__abc_16259_n10590), .Y(AES_CORE_DATAPATH__0iv_0__31_0__2_) );
  AND2X2 AND2X2_3922 ( .A(AES_CORE_DATAPATH__abc_16259_n10594), .B(AES_CORE_DATAPATH__abc_16259_n10593), .Y(AES_CORE_DATAPATH__0iv_0__31_0__3_) );
  AND2X2 AND2X2_3923 ( .A(AES_CORE_DATAPATH__abc_16259_n10597), .B(AES_CORE_DATAPATH__abc_16259_n10596), .Y(AES_CORE_DATAPATH__0iv_0__31_0__4_) );
  AND2X2 AND2X2_3924 ( .A(AES_CORE_DATAPATH__abc_16259_n10600), .B(AES_CORE_DATAPATH__abc_16259_n10599), .Y(AES_CORE_DATAPATH__0iv_0__31_0__5_) );
  AND2X2 AND2X2_3925 ( .A(AES_CORE_DATAPATH__abc_16259_n10603), .B(AES_CORE_DATAPATH__abc_16259_n10602), .Y(AES_CORE_DATAPATH__0iv_0__31_0__6_) );
  AND2X2 AND2X2_3926 ( .A(AES_CORE_DATAPATH__abc_16259_n10606), .B(AES_CORE_DATAPATH__abc_16259_n10605), .Y(AES_CORE_DATAPATH__0iv_0__31_0__7_) );
  AND2X2 AND2X2_3927 ( .A(AES_CORE_DATAPATH__abc_16259_n10609), .B(AES_CORE_DATAPATH__abc_16259_n10608), .Y(AES_CORE_DATAPATH__0iv_0__31_0__8_) );
  AND2X2 AND2X2_3928 ( .A(AES_CORE_DATAPATH__abc_16259_n10612), .B(AES_CORE_DATAPATH__abc_16259_n10611), .Y(AES_CORE_DATAPATH__0iv_0__31_0__9_) );
  AND2X2 AND2X2_3929 ( .A(AES_CORE_DATAPATH__abc_16259_n10615), .B(AES_CORE_DATAPATH__abc_16259_n10614), .Y(AES_CORE_DATAPATH__0iv_0__31_0__10_) );
  AND2X2 AND2X2_393 ( .A(AES_CORE_DATAPATH__abc_16259_n2855_bF_buf4), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_5_), .Y(AES_CORE_DATAPATH__abc_16259_n3055) );
  AND2X2 AND2X2_3930 ( .A(AES_CORE_DATAPATH__abc_16259_n10618), .B(AES_CORE_DATAPATH__abc_16259_n10617), .Y(AES_CORE_DATAPATH__0iv_0__31_0__11_) );
  AND2X2 AND2X2_3931 ( .A(AES_CORE_DATAPATH__abc_16259_n10621), .B(AES_CORE_DATAPATH__abc_16259_n10620), .Y(AES_CORE_DATAPATH__0iv_0__31_0__12_) );
  AND2X2 AND2X2_3932 ( .A(AES_CORE_DATAPATH__abc_16259_n10624), .B(AES_CORE_DATAPATH__abc_16259_n10623), .Y(AES_CORE_DATAPATH__0iv_0__31_0__13_) );
  AND2X2 AND2X2_3933 ( .A(AES_CORE_DATAPATH__abc_16259_n10627), .B(AES_CORE_DATAPATH__abc_16259_n10626), .Y(AES_CORE_DATAPATH__0iv_0__31_0__14_) );
  AND2X2 AND2X2_3934 ( .A(AES_CORE_DATAPATH__abc_16259_n10630), .B(AES_CORE_DATAPATH__abc_16259_n10629), .Y(AES_CORE_DATAPATH__0iv_0__31_0__15_) );
  AND2X2 AND2X2_3935 ( .A(AES_CORE_DATAPATH__abc_16259_n10633), .B(AES_CORE_DATAPATH__abc_16259_n10632), .Y(AES_CORE_DATAPATH__0iv_0__31_0__16_) );
  AND2X2 AND2X2_3936 ( .A(AES_CORE_DATAPATH__abc_16259_n10636), .B(AES_CORE_DATAPATH__abc_16259_n10635), .Y(AES_CORE_DATAPATH__0iv_0__31_0__17_) );
  AND2X2 AND2X2_3937 ( .A(AES_CORE_DATAPATH__abc_16259_n10639), .B(AES_CORE_DATAPATH__abc_16259_n10638), .Y(AES_CORE_DATAPATH__0iv_0__31_0__18_) );
  AND2X2 AND2X2_3938 ( .A(AES_CORE_DATAPATH__abc_16259_n10642), .B(AES_CORE_DATAPATH__abc_16259_n10641), .Y(AES_CORE_DATAPATH__0iv_0__31_0__19_) );
  AND2X2 AND2X2_3939 ( .A(AES_CORE_DATAPATH__abc_16259_n10645), .B(AES_CORE_DATAPATH__abc_16259_n10644), .Y(AES_CORE_DATAPATH__0iv_0__31_0__20_) );
  AND2X2 AND2X2_394 ( .A(AES_CORE_DATAPATH__abc_16259_n2857_bF_buf4), .B(AES_CORE_DATAPATH_MIX_COL_col_0__5_), .Y(AES_CORE_DATAPATH__abc_16259_n3056_1) );
  AND2X2 AND2X2_3940 ( .A(AES_CORE_DATAPATH__abc_16259_n10648), .B(AES_CORE_DATAPATH__abc_16259_n10647), .Y(AES_CORE_DATAPATH__0iv_0__31_0__21_) );
  AND2X2 AND2X2_3941 ( .A(AES_CORE_DATAPATH__abc_16259_n10651), .B(AES_CORE_DATAPATH__abc_16259_n10650), .Y(AES_CORE_DATAPATH__0iv_0__31_0__22_) );
  AND2X2 AND2X2_3942 ( .A(AES_CORE_DATAPATH__abc_16259_n10654), .B(AES_CORE_DATAPATH__abc_16259_n10653), .Y(AES_CORE_DATAPATH__0iv_0__31_0__23_) );
  AND2X2 AND2X2_3943 ( .A(AES_CORE_DATAPATH__abc_16259_n10657), .B(AES_CORE_DATAPATH__abc_16259_n10656), .Y(AES_CORE_DATAPATH__0iv_0__31_0__24_) );
  AND2X2 AND2X2_3944 ( .A(AES_CORE_DATAPATH__abc_16259_n10660), .B(AES_CORE_DATAPATH__abc_16259_n10659), .Y(AES_CORE_DATAPATH__0iv_0__31_0__25_) );
  AND2X2 AND2X2_3945 ( .A(AES_CORE_DATAPATH__abc_16259_n10663), .B(AES_CORE_DATAPATH__abc_16259_n10662), .Y(AES_CORE_DATAPATH__0iv_0__31_0__26_) );
  AND2X2 AND2X2_3946 ( .A(AES_CORE_DATAPATH__abc_16259_n10666), .B(AES_CORE_DATAPATH__abc_16259_n10665), .Y(AES_CORE_DATAPATH__0iv_0__31_0__27_) );
  AND2X2 AND2X2_3947 ( .A(AES_CORE_DATAPATH__abc_16259_n10669), .B(AES_CORE_DATAPATH__abc_16259_n10668), .Y(AES_CORE_DATAPATH__0iv_0__31_0__28_) );
  AND2X2 AND2X2_3948 ( .A(AES_CORE_DATAPATH__abc_16259_n10672), .B(AES_CORE_DATAPATH__abc_16259_n10671), .Y(AES_CORE_DATAPATH__0iv_0__31_0__29_) );
  AND2X2 AND2X2_3949 ( .A(AES_CORE_DATAPATH__abc_16259_n10675), .B(AES_CORE_DATAPATH__abc_16259_n10674), .Y(AES_CORE_DATAPATH__0iv_0__31_0__30_) );
  AND2X2 AND2X2_395 ( .A(AES_CORE_DATAPATH__abc_16259_n3054_1), .B(AES_CORE_DATAPATH__abc_16259_n3058), .Y(AES_CORE_DATAPATH__abc_16259_n3059) );
  AND2X2 AND2X2_3950 ( .A(AES_CORE_DATAPATH__abc_16259_n10678), .B(AES_CORE_DATAPATH__abc_16259_n10677), .Y(AES_CORE_DATAPATH__0iv_0__31_0__31_) );
  AND2X2 AND2X2_3951 ( .A(AES_CORE_DATAPATH__abc_16259_n10681), .B(AES_CORE_DATAPATH__abc_16259_n10680), .Y(AES_CORE_DATAPATH_key_en_pp1_0__FF_INPUT) );
  AND2X2 AND2X2_3952 ( .A(AES_CORE_DATAPATH__abc_16259_n10684), .B(AES_CORE_DATAPATH__abc_16259_n10683), .Y(AES_CORE_DATAPATH_key_en_pp1_1__FF_INPUT) );
  AND2X2 AND2X2_3953 ( .A(AES_CORE_DATAPATH__abc_16259_n10687), .B(AES_CORE_DATAPATH__abc_16259_n10686), .Y(AES_CORE_DATAPATH_key_en_pp1_2__FF_INPUT) );
  AND2X2 AND2X2_3954 ( .A(AES_CORE_DATAPATH__abc_16259_n10690), .B(AES_CORE_DATAPATH__abc_16259_n10689), .Y(AES_CORE_DATAPATH_key_en_pp1_3__FF_INPUT) );
  AND2X2 AND2X2_3955 ( .A(AES_CORE_DATAPATH__abc_16259_n10693), .B(AES_CORE_DATAPATH__abc_16259_n10692), .Y(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_0__FF_INPUT) );
  AND2X2 AND2X2_3956 ( .A(AES_CORE_DATAPATH__abc_16259_n10696), .B(AES_CORE_DATAPATH__abc_16259_n10695), .Y(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_1__FF_INPUT) );
  AND2X2 AND2X2_3957 ( .A(AES_CORE_DATAPATH__abc_16259_n10699), .B(AES_CORE_DATAPATH__abc_16259_n10698), .Y(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_2__FF_INPUT) );
  AND2X2 AND2X2_3958 ( .A(AES_CORE_DATAPATH__abc_16259_n10702), .B(AES_CORE_DATAPATH__abc_16259_n10701), .Y(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_3__FF_INPUT) );
  AND2X2 AND2X2_3959 ( .A(AES_CORE_DATAPATH__abc_16259_n10705), .B(AES_CORE_DATAPATH__abc_16259_n10704), .Y(AES_CORE_DATAPATH_col_en_cnt_unit_pp1_0__FF_INPUT) );
  AND2X2 AND2X2_396 ( .A(_auto_iopadmap_cc_313_execute_26949_5_), .B(AES_CORE_DATAPATH__abc_16259_n3059), .Y(AES_CORE_DATAPATH__abc_16259_n3062_1) );
  AND2X2 AND2X2_3960 ( .A(AES_CORE_DATAPATH__abc_16259_n10708), .B(AES_CORE_DATAPATH__abc_16259_n10707), .Y(AES_CORE_DATAPATH_col_en_cnt_unit_pp1_1__FF_INPUT) );
  AND2X2 AND2X2_3961 ( .A(AES_CORE_DATAPATH__abc_16259_n10711), .B(AES_CORE_DATAPATH__abc_16259_n10710), .Y(AES_CORE_DATAPATH_col_en_cnt_unit_pp1_2__FF_INPUT) );
  AND2X2 AND2X2_3962 ( .A(AES_CORE_DATAPATH__abc_16259_n10714), .B(AES_CORE_DATAPATH__abc_16259_n10713), .Y(AES_CORE_DATAPATH_col_en_cnt_unit_pp1_3__FF_INPUT) );
  AND2X2 AND2X2_3963 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf10), .B(AES_CORE_CONTROL_UNIT_bypass_key_en), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out) );
  AND2X2 AND2X2_3964 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n328_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n330_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n331_1) );
  AND2X2 AND2X2_3965 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_0_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out_bF_buf4), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n333_1) );
  AND2X2 AND2X2_3966 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n334_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n336_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_64_) );
  AND2X2 AND2X2_3967 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n339_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n341_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n342_1) );
  AND2X2 AND2X2_3968 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_1_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n344_1) );
  AND2X2 AND2X2_3969 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n345_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n347_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_65_) );
  AND2X2 AND2X2_397 ( .A(AES_CORE_DATAPATH_last_round_pp2_bF_buf3), .B(AES_CORE_DATAPATH_MIX_COL_col_0__5_), .Y(AES_CORE_DATAPATH__abc_16259_n3065_1) );
  AND2X2 AND2X2_3970 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n350_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n352_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n353_1) );
  AND2X2 AND2X2_3971 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_2_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n355_1) );
  AND2X2 AND2X2_3972 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n356_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n358_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_66_) );
  AND2X2 AND2X2_3973 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n361_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n363_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n364_1) );
  AND2X2 AND2X2_3974 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_3_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n366_1) );
  AND2X2 AND2X2_3975 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n367_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n369_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_67_) );
  AND2X2 AND2X2_3976 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n372_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n374_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n375_1) );
  AND2X2 AND2X2_3977 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_4_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n377_1) );
  AND2X2 AND2X2_3978 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n378_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n380_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_68_) );
  AND2X2 AND2X2_3979 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n383_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n385_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n386_1) );
  AND2X2 AND2X2_398 ( .A(AES_CORE_DATAPATH__abc_16259_n2798_bF_buf4), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_5_), .Y(AES_CORE_DATAPATH__abc_16259_n3066) );
  AND2X2 AND2X2_3980 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_5_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n388_1) );
  AND2X2 AND2X2_3981 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n389_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n391_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_69_) );
  AND2X2 AND2X2_3982 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n394_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n396_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n397_1) );
  AND2X2 AND2X2_3983 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_6_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n399_1) );
  AND2X2 AND2X2_3984 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n400_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n402_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_70_) );
  AND2X2 AND2X2_3985 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n405_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n407_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n408_1) );
  AND2X2 AND2X2_3986 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_7_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n410_1) );
  AND2X2 AND2X2_3987 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n411_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n413_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_71_) );
  AND2X2 AND2X2_3988 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n416_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n418_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n419_1) );
  AND2X2 AND2X2_3989 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_8_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n421_1) );
  AND2X2 AND2X2_399 ( .A(AES_CORE_DATAPATH__abc_16259_n3064), .B(AES_CORE_DATAPATH__abc_16259_n3068), .Y(AES_CORE_DATAPATH__abc_16259_n3069_1) );
  AND2X2 AND2X2_3990 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n422_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n424_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_72_) );
  AND2X2 AND2X2_3991 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n427_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n429_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n430_1) );
  AND2X2 AND2X2_3992 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_9_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n432_1) );
  AND2X2 AND2X2_3993 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n433_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n435_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_73_) );
  AND2X2 AND2X2_3994 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n438_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n440_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n441_1) );
  AND2X2 AND2X2_3995 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_10_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n443_1) );
  AND2X2 AND2X2_3996 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n444_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n446_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_74_) );
  AND2X2 AND2X2_3997 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n449_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n451_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n452_1) );
  AND2X2 AND2X2_3998 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_11_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n454_1) );
  AND2X2 AND2X2_3999 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n455_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n457_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_75_) );
  AND2X2 AND2X2_4 ( .A(_abc_15830_n15), .B(_abc_15830_n11_1), .Y(AES_CORE_DATAPATH_col_en_host_1_) );
  AND2X2 AND2X2_40 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n85), .B(AES_CORE_CONTROL_UNIT_state_1_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n134) );
  AND2X2 AND2X2_400 ( .A(AES_CORE_DATAPATH__abc_16259_n3069_1), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf14), .Y(AES_CORE_DATAPATH__abc_16259_n3070) );
  AND2X2 AND2X2_4000 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n460_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n462_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n463_1) );
  AND2X2 AND2X2_4001 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_12_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n465_1) );
  AND2X2 AND2X2_4002 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n466_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n468_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_76_) );
  AND2X2 AND2X2_4003 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n471_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n473_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n474_1) );
  AND2X2 AND2X2_4004 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_13_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n476_1) );
  AND2X2 AND2X2_4005 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n477_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n479_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_77_) );
  AND2X2 AND2X2_4006 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n482_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n484_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n485_1) );
  AND2X2 AND2X2_4007 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_14_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n487_1) );
  AND2X2 AND2X2_4008 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n488_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n490_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_78_) );
  AND2X2 AND2X2_4009 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n493_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n495_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n496_1) );
  AND2X2 AND2X2_401 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf6), .B(AES_CORE_DATAPATH_col_3__5_), .Y(AES_CORE_DATAPATH__abc_16259_n3071_1) );
  AND2X2 AND2X2_4010 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_15_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n498_1) );
  AND2X2 AND2X2_4011 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n499_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n501_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_79_) );
  AND2X2 AND2X2_4012 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n504), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n506), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n507) );
  AND2X2 AND2X2_4013 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_16_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n509) );
  AND2X2 AND2X2_4014 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n510), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n512), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_80_) );
  AND2X2 AND2X2_4015 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n515), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n517), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n518) );
  AND2X2 AND2X2_4016 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_17_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n520) );
  AND2X2 AND2X2_4017 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n521), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n523), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_81_) );
  AND2X2 AND2X2_4018 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n526), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n528), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n529) );
  AND2X2 AND2X2_4019 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_18_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n531) );
  AND2X2 AND2X2_402 ( .A(AES_CORE_DATAPATH__abc_16259_n3074), .B(AES_CORE_DATAPATH__abc_16259_n3076), .Y(AES_CORE_DATAPATH__abc_16259_n3077) );
  AND2X2 AND2X2_4020 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n532), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n534), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_82_) );
  AND2X2 AND2X2_4021 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n537), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n539), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n540) );
  AND2X2 AND2X2_4022 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_19_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n542) );
  AND2X2 AND2X2_4023 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n543), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n545), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_83_) );
  AND2X2 AND2X2_4024 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n548), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n550), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n551) );
  AND2X2 AND2X2_4025 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_20_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n553) );
  AND2X2 AND2X2_4026 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n554), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n556), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_84_) );
  AND2X2 AND2X2_4027 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n559), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n561), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n562) );
  AND2X2 AND2X2_4028 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_21_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n564) );
  AND2X2 AND2X2_4029 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n565), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n567), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_85_) );
  AND2X2 AND2X2_403 ( .A(AES_CORE_DATAPATH__abc_16259_n2782_bF_buf3), .B(AES_CORE_DATAPATH_col_3__6_), .Y(AES_CORE_DATAPATH__abc_16259_n3078) );
  AND2X2 AND2X2_4030 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n570), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n572), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n573) );
  AND2X2 AND2X2_4031 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_22_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n575) );
  AND2X2 AND2X2_4032 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n576), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n578), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_86_) );
  AND2X2 AND2X2_4033 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n581), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n583), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n584) );
  AND2X2 AND2X2_4034 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_23_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n586) );
  AND2X2 AND2X2_4035 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n587), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n589), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_87_) );
  AND2X2 AND2X2_4036 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__24_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__24_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n592) );
  AND2X2 AND2X2_4037 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n593), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n591), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n594) );
  AND2X2 AND2X2_4038 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n599), .B(AES_CORE_DATAPATH_KEY_EXPANDER_round_0_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n600) );
  AND2X2 AND2X2_4039 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n600), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n598), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n601) );
  AND2X2 AND2X2_404 ( .A(AES_CORE_DATAPATH__abc_16259_n2786_bF_buf3), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_70_), .Y(AES_CORE_DATAPATH__abc_16259_n3079) );
  AND2X2 AND2X2_4040 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n602), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597_bF_buf4), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n603) );
  AND2X2 AND2X2_4041 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n605), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf6), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n606) );
  AND2X2 AND2X2_4042 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n607), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_24_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n608) );
  AND2X2 AND2X2_4043 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n609), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n610), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n611) );
  AND2X2 AND2X2_4044 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n613), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n595), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n614) );
  AND2X2 AND2X2_4045 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n612), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n594), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n615) );
  AND2X2 AND2X2_4046 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__25_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__25_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n618) );
  AND2X2 AND2X2_4047 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n619), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n617), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n620) );
  AND2X2 AND2X2_4048 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n626), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597_bF_buf3), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n627) );
  AND2X2 AND2X2_4049 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n627), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n605), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n628) );
  AND2X2 AND2X2_405 ( .A(AES_CORE_DATAPATH__abc_16259_n2789_bF_buf3), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_38_), .Y(AES_CORE_DATAPATH__abc_16259_n3080) );
  AND2X2 AND2X2_4050 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n599), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n623), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n629) );
  AND2X2 AND2X2_4051 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n598), .B(AES_CORE_DATAPATH_KEY_EXPANDER_round_3_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n630) );
  AND2X2 AND2X2_4052 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n629), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n630), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n631) );
  AND2X2 AND2X2_4053 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n633), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n602), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n634) );
  AND2X2 AND2X2_4054 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n635), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n622), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n637) );
  AND2X2 AND2X2_4055 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n638), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n636), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n639) );
  AND2X2 AND2X2_4056 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n639), .B(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out_bF_buf4), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n640) );
  AND2X2 AND2X2_4057 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n640), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n621), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n641) );
  AND2X2 AND2X2_4058 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n643), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n642), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n644) );
  AND2X2 AND2X2_4059 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n644), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_25_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n645) );
  AND2X2 AND2X2_406 ( .A(AES_CORE_DATAPATH__abc_16259_n3083_1), .B(AES_CORE_DATAPATH__abc_16259_n3077), .Y(AES_CORE_DATAPATH__abc_16259_n3084) );
  AND2X2 AND2X2_4060 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n647), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n620), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n648) );
  AND2X2 AND2X2_4061 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__26_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__26_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n651) );
  AND2X2 AND2X2_4062 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n652), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n650), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n653) );
  AND2X2 AND2X2_4063 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n656), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n598), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n659) );
  AND2X2 AND2X2_4064 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n623), .B(AES_CORE_DATAPATH_KEY_EXPANDER_round_1_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n660) );
  AND2X2 AND2X2_4065 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n659), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n660), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n661) );
  AND2X2 AND2X2_4066 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n658), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n662), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n663) );
  AND2X2 AND2X2_4067 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n659), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n629), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n665) );
  AND2X2 AND2X2_4068 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_round_1_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_round_0_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n666) );
  AND2X2 AND2X2_4069 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n656), .B(AES_CORE_DATAPATH_KEY_EXPANDER_round_2_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n667) );
  AND2X2 AND2X2_407 ( .A(AES_CORE_DATAPATH__abc_16259_n2837_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__6_), .Y(AES_CORE_DATAPATH__abc_16259_n3086) );
  AND2X2 AND2X2_4070 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n667), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n666), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n668) );
  AND2X2 AND2X2_4071 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n627), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n669), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n670) );
  AND2X2 AND2X2_4072 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n664), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n671), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n672) );
  AND2X2 AND2X2_4073 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n672), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n655), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n673) );
  AND2X2 AND2X2_4074 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n674), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n675), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n676) );
  AND2X2 AND2X2_4075 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n676), .B(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out_bF_buf3), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n677) );
  AND2X2 AND2X2_4076 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n677), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n654), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n678) );
  AND2X2 AND2X2_4077 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n679), .B(AES_CORE_DATAPATH_KEY_EXPANDER_round_3_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n680) );
  AND2X2 AND2X2_4078 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n680), .B(AES_CORE_DATAPATH_KEY_EXPANDER_round_0_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n681) );
  AND2X2 AND2X2_4079 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n682), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n633), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n683) );
  AND2X2 AND2X2_408 ( .A(AES_CORE_DATAPATH__abc_16259_n2887_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__6_), .Y(AES_CORE_DATAPATH__abc_16259_n3088) );
  AND2X2 AND2X2_4080 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n684), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_26_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n685) );
  AND2X2 AND2X2_4081 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n687), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n653), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n688) );
  AND2X2 AND2X2_4082 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__27_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__27_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n691) );
  AND2X2 AND2X2_4083 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n692), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n690), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n693) );
  AND2X2 AND2X2_4084 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n659), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n600), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n695) );
  AND2X2 AND2X2_4085 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n660), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n667), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n697) );
  AND2X2 AND2X2_4086 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n659), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n666), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n699) );
  AND2X2 AND2X2_4087 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n698), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n700), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n701) );
  AND2X2 AND2X2_4088 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n701), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_27_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n702) );
  AND2X2 AND2X2_4089 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n703), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n704), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n705) );
  AND2X2 AND2X2_409 ( .A(AES_CORE_DATAPATH__abc_16259_n2830_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__6_), .Y(AES_CORE_DATAPATH__abc_16259_n3089) );
  AND2X2 AND2X2_4090 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n705), .B(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out_bF_buf2), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n706) );
  AND2X2 AND2X2_4091 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n706), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n694), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n707) );
  AND2X2 AND2X2_4092 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n708), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n693), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n709) );
  AND2X2 AND2X2_4093 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__28_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__28_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n712) );
  AND2X2 AND2X2_4094 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n713), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n711), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n714) );
  AND2X2 AND2X2_4095 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n659), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n599), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n717) );
  AND2X2 AND2X2_4096 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n600), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n667), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n719) );
  AND2X2 AND2X2_4097 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n629), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n667), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n722) );
  AND2X2 AND2X2_4098 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n658), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n723), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n724) );
  AND2X2 AND2X2_4099 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n724), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n633), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n725) );
  AND2X2 AND2X2_41 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n107), .B(AES_CORE_CONTROL_UNIT__abc_15841_n114_1), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n135) );
  AND2X2 AND2X2_410 ( .A(AES_CORE_DATAPATH__abc_16259_n3091_1), .B(AES_CORE_DATAPATH__abc_16259_n3092), .Y(_auto_iopadmap_cc_313_execute_26949_6_) );
  AND2X2 AND2X2_4100 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n728), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n720), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n729) );
  AND2X2 AND2X2_4101 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n730), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n727), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n731) );
  AND2X2 AND2X2_4102 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n731), .B(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out_bF_buf1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n732) );
  AND2X2 AND2X2_4103 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n732), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n715), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n733) );
  AND2X2 AND2X2_4104 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n729), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_28_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n734) );
  AND2X2 AND2X2_4105 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n726), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n716), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n735) );
  AND2X2 AND2X2_4106 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n737), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n714), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n738) );
  AND2X2 AND2X2_4107 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__29_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__29_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n741) );
  AND2X2 AND2X2_4108 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n742), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n740), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n743) );
  AND2X2 AND2X2_4109 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n658), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n746), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n747) );
  AND2X2 AND2X2_411 ( .A(AES_CORE_DATAPATH__abc_16259_n2855_bF_buf3), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_6_), .Y(AES_CORE_DATAPATH__abc_16259_n3095) );
  AND2X2 AND2X2_4110 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n748), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n751), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n752) );
  AND2X2 AND2X2_4111 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n752), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n745), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n753) );
  AND2X2 AND2X2_4112 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n754), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n755), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n756) );
  AND2X2 AND2X2_4113 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n756), .B(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out_bF_buf0), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n757) );
  AND2X2 AND2X2_4114 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n757), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n744), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n758) );
  AND2X2 AND2X2_4115 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n759), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n633), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n760) );
  AND2X2 AND2X2_4116 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n762), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_29_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n763) );
  AND2X2 AND2X2_4117 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n765), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n743), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n766) );
  AND2X2 AND2X2_4118 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__30_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__30_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n769) );
  AND2X2 AND2X2_4119 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n770), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n768), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n771) );
  AND2X2 AND2X2_412 ( .A(AES_CORE_DATAPATH__abc_16259_n2857_bF_buf3), .B(AES_CORE_DATAPATH_MIX_COL_col_0__6_), .Y(AES_CORE_DATAPATH__abc_16259_n3096_1) );
  AND2X2 AND2X2_4120 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n604), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n656), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n775) );
  AND2X2 AND2X2_4121 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_round_2_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_round_1_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n776) );
  AND2X2 AND2X2_4122 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n775), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n777), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n778) );
  AND2X2 AND2X2_4123 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n667), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf3), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n782) );
  AND2X2 AND2X2_4124 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n782), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n660), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n783) );
  AND2X2 AND2X2_4125 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n781), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n784), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n785) );
  AND2X2 AND2X2_4126 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n627), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n778), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n787) );
  AND2X2 AND2X2_4127 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n787), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n666), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n788) );
  AND2X2 AND2X2_4128 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n786), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n790), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n791) );
  AND2X2 AND2X2_4129 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n791), .B(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out_bF_buf4), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n792) );
  AND2X2 AND2X2_413 ( .A(AES_CORE_DATAPATH__abc_16259_n3094_1), .B(AES_CORE_DATAPATH__abc_16259_n3098_1), .Y(AES_CORE_DATAPATH__abc_16259_n3099) );
  AND2X2 AND2X2_4130 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n792), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n772), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n793) );
  AND2X2 AND2X2_4131 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n789), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_30_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n794) );
  AND2X2 AND2X2_4132 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n785), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n773), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n795) );
  AND2X2 AND2X2_4133 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n797), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n771), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n798) );
  AND2X2 AND2X2_4134 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__31_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__31_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n801) );
  AND2X2 AND2X2_4135 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n802), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n800), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n803) );
  AND2X2 AND2X2_4136 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n782), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n666), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n808) );
  AND2X2 AND2X2_4137 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n807), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n809), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n810) );
  AND2X2 AND2X2_4138 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n787), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n660), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n812) );
  AND2X2 AND2X2_4139 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n811), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n814), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n815) );
  AND2X2 AND2X2_414 ( .A(_auto_iopadmap_cc_313_execute_26949_6_), .B(AES_CORE_DATAPATH__abc_16259_n3099), .Y(AES_CORE_DATAPATH__abc_16259_n3102) );
  AND2X2 AND2X2_4140 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n815), .B(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out_bF_buf3), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n816) );
  AND2X2 AND2X2_4141 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n816), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n804), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n817) );
  AND2X2 AND2X2_4142 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n813), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_31_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n818) );
  AND2X2 AND2X2_4143 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n810), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n805), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n819) );
  AND2X2 AND2X2_4144 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n821), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n803), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n822) );
  AND2X2 AND2X2_4145 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__0_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__0_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n825) );
  AND2X2 AND2X2_4146 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n826), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n824), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_0_) );
  AND2X2 AND2X2_4147 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n828), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n829), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_8_) );
  AND2X2 AND2X2_4148 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__1_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__1_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n832) );
  AND2X2 AND2X2_4149 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n833), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n831), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_1_) );
  AND2X2 AND2X2_415 ( .A(AES_CORE_DATAPATH_last_round_pp2_bF_buf2), .B(AES_CORE_DATAPATH_MIX_COL_col_0__6_), .Y(AES_CORE_DATAPATH__abc_16259_n3105) );
  AND2X2 AND2X2_4150 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n835), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n836), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_9_) );
  AND2X2 AND2X2_4151 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__2_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__2_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n839) );
  AND2X2 AND2X2_4152 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n840), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n838), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_2_) );
  AND2X2 AND2X2_4153 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n842), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n843), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_10_) );
  AND2X2 AND2X2_4154 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__3_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__3_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n846) );
  AND2X2 AND2X2_4155 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n847), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n845), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_3_) );
  AND2X2 AND2X2_4156 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n849), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n850), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_11_) );
  AND2X2 AND2X2_4157 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__4_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__4_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n853) );
  AND2X2 AND2X2_4158 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n854), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n852), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_4_) );
  AND2X2 AND2X2_4159 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n856), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n857), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_12_) );
  AND2X2 AND2X2_416 ( .A(AES_CORE_DATAPATH__abc_16259_n2798_bF_buf3), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_6_), .Y(AES_CORE_DATAPATH__abc_16259_n3106) );
  AND2X2 AND2X2_4160 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__5_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__5_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n860) );
  AND2X2 AND2X2_4161 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n861), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n859), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_5_) );
  AND2X2 AND2X2_4162 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n863), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n864), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_13_) );
  AND2X2 AND2X2_4163 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__6_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__6_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n867) );
  AND2X2 AND2X2_4164 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n868), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n866), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_6_) );
  AND2X2 AND2X2_4165 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n870), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n871), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_14_) );
  AND2X2 AND2X2_4166 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__7_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__7_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n874) );
  AND2X2 AND2X2_4167 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n875), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n873), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_7_) );
  AND2X2 AND2X2_4168 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n877), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n878), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_15_) );
  AND2X2 AND2X2_4169 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__8_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__8_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n881) );
  AND2X2 AND2X2_417 ( .A(AES_CORE_DATAPATH__abc_16259_n3104), .B(AES_CORE_DATAPATH__abc_16259_n3108), .Y(AES_CORE_DATAPATH__abc_16259_n3109) );
  AND2X2 AND2X2_4170 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n882), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n880), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_8_) );
  AND2X2 AND2X2_4171 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n884), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n885), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_16_) );
  AND2X2 AND2X2_4172 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__9_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__9_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n888) );
  AND2X2 AND2X2_4173 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n889), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n887), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_9_) );
  AND2X2 AND2X2_4174 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n891), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n892), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_17_) );
  AND2X2 AND2X2_4175 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__10_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__10_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n895) );
  AND2X2 AND2X2_4176 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n896), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n894), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_10_) );
  AND2X2 AND2X2_4177 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n898), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n899), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_18_) );
  AND2X2 AND2X2_4178 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__11_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__11_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n902) );
  AND2X2 AND2X2_4179 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n903), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n901), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_11_) );
  AND2X2 AND2X2_418 ( .A(AES_CORE_DATAPATH__abc_16259_n3109), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf13), .Y(AES_CORE_DATAPATH__abc_16259_n3110) );
  AND2X2 AND2X2_4180 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n905), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n906), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_19_) );
  AND2X2 AND2X2_4181 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__12_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__12_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n909) );
  AND2X2 AND2X2_4182 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n910), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n908), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_12_) );
  AND2X2 AND2X2_4183 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n912), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n913), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_20_) );
  AND2X2 AND2X2_4184 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__13_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__13_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n916) );
  AND2X2 AND2X2_4185 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n917), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n915), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_13_) );
  AND2X2 AND2X2_4186 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n919), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n920), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_21_) );
  AND2X2 AND2X2_4187 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__14_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__14_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n923) );
  AND2X2 AND2X2_4188 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n924), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n922), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_14_) );
  AND2X2 AND2X2_4189 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n926), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n927), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_22_) );
  AND2X2 AND2X2_419 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf5), .B(AES_CORE_DATAPATH_col_3__6_), .Y(AES_CORE_DATAPATH__abc_16259_n3111) );
  AND2X2 AND2X2_4190 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__15_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__15_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n930) );
  AND2X2 AND2X2_4191 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n931), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n929), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_15_) );
  AND2X2 AND2X2_4192 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n933), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n934), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_23_) );
  AND2X2 AND2X2_4193 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__16_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__16_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n937) );
  AND2X2 AND2X2_4194 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n938), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n936), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_16_) );
  AND2X2 AND2X2_4195 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n940), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n941), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_24_) );
  AND2X2 AND2X2_4196 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__17_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__17_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n944) );
  AND2X2 AND2X2_4197 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n945), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n943), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_17_) );
  AND2X2 AND2X2_4198 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n947), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n948), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_25_) );
  AND2X2 AND2X2_4199 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__18_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__18_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n951) );
  AND2X2 AND2X2_42 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n107), .B(AES_CORE_CONTROL_UNIT__abc_15841_n140), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n141_1) );
  AND2X2 AND2X2_420 ( .A(AES_CORE_DATAPATH__abc_16259_n3114_1), .B(AES_CORE_DATAPATH__abc_16259_n3116), .Y(AES_CORE_DATAPATH__abc_16259_n3117) );
  AND2X2 AND2X2_4200 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n952), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n950), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_18_) );
  AND2X2 AND2X2_4201 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n954), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n955), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_26_) );
  AND2X2 AND2X2_4202 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__19_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__19_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n958) );
  AND2X2 AND2X2_4203 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n959), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n957), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_19_) );
  AND2X2 AND2X2_4204 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n961), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n962), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_27_) );
  AND2X2 AND2X2_4205 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__20_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__20_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n965) );
  AND2X2 AND2X2_4206 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n966), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n964), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_20_) );
  AND2X2 AND2X2_4207 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n968), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n969), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_28_) );
  AND2X2 AND2X2_4208 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__21_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__21_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n972) );
  AND2X2 AND2X2_4209 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n973), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n971), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_21_) );
  AND2X2 AND2X2_421 ( .A(AES_CORE_DATAPATH__abc_16259_n2782_bF_buf2), .B(AES_CORE_DATAPATH_col_3__7_), .Y(AES_CORE_DATAPATH__abc_16259_n3118) );
  AND2X2 AND2X2_4210 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n975), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n976), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_29_) );
  AND2X2 AND2X2_4211 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__22_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__22_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n979) );
  AND2X2 AND2X2_4212 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n980), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n978), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_22_) );
  AND2X2 AND2X2_4213 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n982), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n983), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_30_) );
  AND2X2 AND2X2_4214 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__23_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__23_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n986) );
  AND2X2 AND2X2_4215 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n987), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n985), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_23_) );
  AND2X2 AND2X2_4216 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n989), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n990), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_31_) );
  AND2X2 AND2X2_4217 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__24_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__24_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n993) );
  AND2X2 AND2X2_4218 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n994), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n992), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_24_) );
  AND2X2 AND2X2_4219 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n996), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n997), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_0_) );
  AND2X2 AND2X2_422 ( .A(AES_CORE_DATAPATH__abc_16259_n2786_bF_buf2), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_71_), .Y(AES_CORE_DATAPATH__abc_16259_n3119_1) );
  AND2X2 AND2X2_4220 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__25_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__25_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1000) );
  AND2X2 AND2X2_4221 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1001), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n999), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_25_) );
  AND2X2 AND2X2_4222 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1003), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1004), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_1_) );
  AND2X2 AND2X2_4223 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__26_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__26_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1007) );
  AND2X2 AND2X2_4224 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1008), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1006), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_26_) );
  AND2X2 AND2X2_4225 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1010), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1011), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_2_) );
  AND2X2 AND2X2_4226 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__27_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__27_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1014) );
  AND2X2 AND2X2_4227 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1015), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1013), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_27_) );
  AND2X2 AND2X2_4228 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1017), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1018), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_3_) );
  AND2X2 AND2X2_4229 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__28_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__28_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1021) );
  AND2X2 AND2X2_423 ( .A(AES_CORE_DATAPATH__abc_16259_n2789_bF_buf2), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_39_), .Y(AES_CORE_DATAPATH__abc_16259_n3120_1) );
  AND2X2 AND2X2_4230 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1022), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1020), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_28_) );
  AND2X2 AND2X2_4231 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1024), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1025), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_4_) );
  AND2X2 AND2X2_4232 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__29_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__29_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1028) );
  AND2X2 AND2X2_4233 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1029), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1027), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_29_) );
  AND2X2 AND2X2_4234 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1031), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1032), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_5_) );
  AND2X2 AND2X2_4235 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__30_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__30_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1035) );
  AND2X2 AND2X2_4236 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1036), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1034), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_30_) );
  AND2X2 AND2X2_4237 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1038), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1039), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_6_) );
  AND2X2 AND2X2_4238 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__31_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__31_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1042) );
  AND2X2 AND2X2_4239 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1043), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1041), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_31_) );
  AND2X2 AND2X2_424 ( .A(AES_CORE_DATAPATH__abc_16259_n3123_1), .B(AES_CORE_DATAPATH__abc_16259_n3117), .Y(AES_CORE_DATAPATH__abc_16259_n3124) );
  AND2X2 AND2X2_4240 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1045), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1046), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_7_) );
  AND2X2 AND2X2_4241 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__0_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_0_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1049) );
  AND2X2 AND2X2_4242 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1050), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1048), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_96_) );
  AND2X2 AND2X2_4243 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__1_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_1_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1053) );
  AND2X2 AND2X2_4244 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1054), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1052), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_97_) );
  AND2X2 AND2X2_4245 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__2_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_2_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1057) );
  AND2X2 AND2X2_4246 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1058), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1056), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_98_) );
  AND2X2 AND2X2_4247 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__3_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_3_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1061) );
  AND2X2 AND2X2_4248 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1062), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1060), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_99_) );
  AND2X2 AND2X2_4249 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__4_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_4_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1065) );
  AND2X2 AND2X2_425 ( .A(AES_CORE_DATAPATH__abc_16259_n2837_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__7_), .Y(AES_CORE_DATAPATH__abc_16259_n3126) );
  AND2X2 AND2X2_4250 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1066), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1064), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_100_) );
  AND2X2 AND2X2_4251 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__5_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_5_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1069) );
  AND2X2 AND2X2_4252 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1070), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1068), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_101_) );
  AND2X2 AND2X2_4253 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__6_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_6_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1073) );
  AND2X2 AND2X2_4254 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1074), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1072), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_102_) );
  AND2X2 AND2X2_4255 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__7_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_7_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1077) );
  AND2X2 AND2X2_4256 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1078), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1076), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_103_) );
  AND2X2 AND2X2_4257 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__8_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_8_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1081) );
  AND2X2 AND2X2_4258 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1082), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1080), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_104_) );
  AND2X2 AND2X2_4259 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__9_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_9_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1085) );
  AND2X2 AND2X2_426 ( .A(AES_CORE_DATAPATH__abc_16259_n2887_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__7_), .Y(AES_CORE_DATAPATH__abc_16259_n3128) );
  AND2X2 AND2X2_4260 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1086), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1084), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_105_) );
  AND2X2 AND2X2_4261 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__10_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_10_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1089) );
  AND2X2 AND2X2_4262 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1090), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1088), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_106_) );
  AND2X2 AND2X2_4263 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__11_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_11_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1093) );
  AND2X2 AND2X2_4264 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1094), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1092), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_107_) );
  AND2X2 AND2X2_4265 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__12_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_12_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1097) );
  AND2X2 AND2X2_4266 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1098), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1096), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_108_) );
  AND2X2 AND2X2_4267 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__13_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_13_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1101) );
  AND2X2 AND2X2_4268 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1102), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1100), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_109_) );
  AND2X2 AND2X2_4269 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__14_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_14_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1105) );
  AND2X2 AND2X2_427 ( .A(AES_CORE_DATAPATH__abc_16259_n2830_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__7_), .Y(AES_CORE_DATAPATH__abc_16259_n3129_1) );
  AND2X2 AND2X2_4270 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1106), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1104), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_110_) );
  AND2X2 AND2X2_4271 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__15_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_15_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1109) );
  AND2X2 AND2X2_4272 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1110), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1108), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_111_) );
  AND2X2 AND2X2_4273 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__16_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_16_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1113) );
  AND2X2 AND2X2_4274 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1114), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1112), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_112_) );
  AND2X2 AND2X2_4275 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__17_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_17_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1117) );
  AND2X2 AND2X2_4276 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1118), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1116), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_113_) );
  AND2X2 AND2X2_4277 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__18_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_18_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1121) );
  AND2X2 AND2X2_4278 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1122), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1120), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_114_) );
  AND2X2 AND2X2_4279 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__19_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_19_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1125) );
  AND2X2 AND2X2_428 ( .A(AES_CORE_DATAPATH__abc_16259_n3131), .B(AES_CORE_DATAPATH__abc_16259_n3132), .Y(_auto_iopadmap_cc_313_execute_26949_7_) );
  AND2X2 AND2X2_4280 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1126), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1124), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_115_) );
  AND2X2 AND2X2_4281 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__20_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_20_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1129) );
  AND2X2 AND2X2_4282 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1130), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1128), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_116_) );
  AND2X2 AND2X2_4283 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__21_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_21_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1133) );
  AND2X2 AND2X2_4284 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1134), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1132), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_117_) );
  AND2X2 AND2X2_4285 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__22_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_22_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1137) );
  AND2X2 AND2X2_4286 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1138), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1136), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_118_) );
  AND2X2 AND2X2_4287 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__23_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_23_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1141) );
  AND2X2 AND2X2_4288 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1142), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1140), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_119_) );
  AND2X2 AND2X2_4289 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1145), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1144), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1146) );
  AND2X2 AND2X2_429 ( .A(AES_CORE_DATAPATH__abc_16259_n2855_bF_buf2), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_7_), .Y(AES_CORE_DATAPATH__abc_16259_n3135) );
  AND2X2 AND2X2_4290 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n611), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__24_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1147) );
  AND2X2 AND2X2_4291 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1150), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1151), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_121_) );
  AND2X2 AND2X2_4292 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n686), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__26_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1153) );
  AND2X2 AND2X2_4293 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n676), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1154), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1155) );
  AND2X2 AND2X2_4294 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1159), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1160), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_123_) );
  AND2X2 AND2X2_4295 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1163), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1164), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_124_) );
  AND2X2 AND2X2_4296 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n764), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__29_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1166) );
  AND2X2 AND2X2_4297 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n756), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1167), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1168) );
  AND2X2 AND2X2_4298 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1170), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1172), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_126_) );
  AND2X2 AND2X2_4299 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1174), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1176), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_127_) );
  AND2X2 AND2X2_43 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n142), .B(AES_CORE_CONTROL_UNIT_state_9_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n143) );
  AND2X2 AND2X2_430 ( .A(AES_CORE_DATAPATH__abc_16259_n2857_bF_buf2), .B(AES_CORE_DATAPATH_MIX_COL_col_0__7_), .Y(AES_CORE_DATAPATH__abc_16259_n3136) );
  AND2X2 AND2X2_4300 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__0_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__0_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1179) );
  AND2X2 AND2X2_4301 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1180), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1178), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_32_) );
  AND2X2 AND2X2_4302 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__1_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__1_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1183) );
  AND2X2 AND2X2_4303 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1184), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1182), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_33_) );
  AND2X2 AND2X2_4304 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__2_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__2_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1187) );
  AND2X2 AND2X2_4305 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1188), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1186), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_34_) );
  AND2X2 AND2X2_4306 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__3_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__3_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1191) );
  AND2X2 AND2X2_4307 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1192), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1190), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_35_) );
  AND2X2 AND2X2_4308 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__4_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__4_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1195) );
  AND2X2 AND2X2_4309 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1196), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1194), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_36_) );
  AND2X2 AND2X2_431 ( .A(AES_CORE_DATAPATH__abc_16259_n3134), .B(AES_CORE_DATAPATH__abc_16259_n3138), .Y(AES_CORE_DATAPATH__abc_16259_n3139) );
  AND2X2 AND2X2_4310 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__5_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__5_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1199) );
  AND2X2 AND2X2_4311 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1200), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1198), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_37_) );
  AND2X2 AND2X2_4312 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__6_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__6_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1203) );
  AND2X2 AND2X2_4313 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1204), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1202), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_38_) );
  AND2X2 AND2X2_4314 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__7_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__7_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1207) );
  AND2X2 AND2X2_4315 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1208), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1206), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_39_) );
  AND2X2 AND2X2_4316 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__8_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__8_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1211) );
  AND2X2 AND2X2_4317 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1212), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1210), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_40_) );
  AND2X2 AND2X2_4318 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__9_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__9_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1215) );
  AND2X2 AND2X2_4319 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1216), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1214), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_41_) );
  AND2X2 AND2X2_432 ( .A(_auto_iopadmap_cc_313_execute_26949_7_), .B(AES_CORE_DATAPATH__abc_16259_n3139), .Y(AES_CORE_DATAPATH__abc_16259_n3142) );
  AND2X2 AND2X2_4320 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__10_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__10_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1219) );
  AND2X2 AND2X2_4321 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1220), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1218), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_42_) );
  AND2X2 AND2X2_4322 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__11_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__11_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1223) );
  AND2X2 AND2X2_4323 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1224), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1222), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_43_) );
  AND2X2 AND2X2_4324 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__12_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__12_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1227) );
  AND2X2 AND2X2_4325 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1228), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1226), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_44_) );
  AND2X2 AND2X2_4326 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__13_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__13_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1231) );
  AND2X2 AND2X2_4327 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1232), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1230), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_45_) );
  AND2X2 AND2X2_4328 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__14_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__14_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1235) );
  AND2X2 AND2X2_4329 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1236), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1234), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_46_) );
  AND2X2 AND2X2_433 ( .A(AES_CORE_DATAPATH_last_round_pp2_bF_buf1), .B(AES_CORE_DATAPATH_MIX_COL_col_0__7_), .Y(AES_CORE_DATAPATH__abc_16259_n3145) );
  AND2X2 AND2X2_4330 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__15_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__15_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1239) );
  AND2X2 AND2X2_4331 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1240), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1238), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_47_) );
  AND2X2 AND2X2_4332 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__16_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__16_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1243) );
  AND2X2 AND2X2_4333 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1244), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1242), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_48_) );
  AND2X2 AND2X2_4334 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__17_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__17_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1247) );
  AND2X2 AND2X2_4335 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1248), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1246), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_49_) );
  AND2X2 AND2X2_4336 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__18_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__18_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1251) );
  AND2X2 AND2X2_4337 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1252), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1250), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_50_) );
  AND2X2 AND2X2_4338 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__19_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__19_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1255) );
  AND2X2 AND2X2_4339 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1256), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1254), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_51_) );
  AND2X2 AND2X2_434 ( .A(AES_CORE_DATAPATH__abc_16259_n2798_bF_buf2), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_7_), .Y(AES_CORE_DATAPATH__abc_16259_n3146) );
  AND2X2 AND2X2_4340 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__20_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__20_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1259) );
  AND2X2 AND2X2_4341 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1260), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1258), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_52_) );
  AND2X2 AND2X2_4342 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__21_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__21_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1263) );
  AND2X2 AND2X2_4343 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1264), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1262), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_53_) );
  AND2X2 AND2X2_4344 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__22_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__22_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1267) );
  AND2X2 AND2X2_4345 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1268), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1266), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_54_) );
  AND2X2 AND2X2_4346 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__23_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__23_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1271) );
  AND2X2 AND2X2_4347 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1272), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1270), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_55_) );
  AND2X2 AND2X2_4348 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__24_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__24_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1275) );
  AND2X2 AND2X2_4349 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1276), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1274), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_56_) );
  AND2X2 AND2X2_435 ( .A(AES_CORE_DATAPATH__abc_16259_n3144), .B(AES_CORE_DATAPATH__abc_16259_n3148_1), .Y(AES_CORE_DATAPATH__abc_16259_n3149_1) );
  AND2X2 AND2X2_4350 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__25_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__25_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1279) );
  AND2X2 AND2X2_4351 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1280), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1278), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_57_) );
  AND2X2 AND2X2_4352 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__26_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__26_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1283) );
  AND2X2 AND2X2_4353 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1284), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1282), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_58_) );
  AND2X2 AND2X2_4354 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__27_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__27_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1287) );
  AND2X2 AND2X2_4355 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1288), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1286), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_59_) );
  AND2X2 AND2X2_4356 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__28_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__28_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1291) );
  AND2X2 AND2X2_4357 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1292), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1290), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_60_) );
  AND2X2 AND2X2_4358 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__29_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__29_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1295) );
  AND2X2 AND2X2_4359 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1296), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1294), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_61_) );
  AND2X2 AND2X2_436 ( .A(AES_CORE_DATAPATH__abc_16259_n3149_1), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf12), .Y(AES_CORE_DATAPATH__abc_16259_n3150) );
  AND2X2 AND2X2_4360 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__30_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__30_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1299) );
  AND2X2 AND2X2_4361 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1300), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1298), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_62_) );
  AND2X2 AND2X2_4362 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__31_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__31_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1303) );
  AND2X2 AND2X2_4363 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1304), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1302), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_63_) );
  AND2X2 AND2X2_4364 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n97_1), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n98), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n99) );
  AND2X2 AND2X2_4365 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__0_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n100) );
  AND2X2 AND2X2_4366 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n103), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n105_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n106) );
  AND2X2 AND2X2_4367 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n107), .B(AES_CORE_DATAPATH_MIX_COL_col_2__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n108) );
  AND2X2 AND2X2_4368 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n106), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n109_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n110) );
  AND2X2 AND2X2_4369 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n114), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n113), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n115_1) );
  AND2X2 AND2X2_437 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf4), .B(AES_CORE_DATAPATH_col_3__7_), .Y(AES_CORE_DATAPATH__abc_16259_n3151) );
  AND2X2 AND2X2_4370 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n117), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n112), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_0_) );
  AND2X2 AND2X2_4371 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n120), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n121), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n122) );
  AND2X2 AND2X2_4372 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__6_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n123_1) );
  AND2X2 AND2X2_4373 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__5_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n126) );
  AND2X2 AND2X2_4374 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n127_1), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n125), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n128) );
  AND2X2 AND2X2_4375 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__5_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n130) );
  AND2X2 AND2X2_4376 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n131), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n129_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n132) );
  AND2X2 AND2X2_4377 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n134_1), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n135), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n136_1) );
  AND2X2 AND2X2_4378 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n138), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n139), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n140_1) );
  AND2X2 AND2X2_4379 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n142_1), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n133), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n143) );
  AND2X2 AND2X2_438 ( .A(AES_CORE_DATAPATH__abc_16259_n3154_1), .B(AES_CORE_DATAPATH__abc_16259_n3156_1), .Y(AES_CORE_DATAPATH__abc_16259_n3157) );
  AND2X2 AND2X2_4380 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n146), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n145), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n147_1) );
  AND2X2 AND2X2_4381 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n137), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n141), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n148) );
  AND2X2 AND2X2_4382 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n128), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n132), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n149_1) );
  AND2X2 AND2X2_4383 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n144), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n151), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n152) );
  AND2X2 AND2X2_4384 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n154_1), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n155), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n156_1) );
  AND2X2 AND2X2_4385 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n153), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n157), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_0_) );
  AND2X2 AND2X2_4386 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n159), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n161), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n162_1) );
  AND2X2 AND2X2_4387 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n107), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n162_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n163) );
  AND2X2 AND2X2_4388 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n164), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n165), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n166_1) );
  AND2X2 AND2X2_4389 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__1_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n169) );
  AND2X2 AND2X2_439 ( .A(AES_CORE_DATAPATH__abc_16259_n2782_bF_buf1), .B(AES_CORE_DATAPATH_col_3__8_), .Y(AES_CORE_DATAPATH__abc_16259_n3158_1) );
  AND2X2 AND2X2_4390 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n170), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n168_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n171) );
  AND2X2 AND2X2_4391 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n171), .B(AES_CORE_DATAPATH_MIX_COL_col_2__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n172_1) );
  AND2X2 AND2X2_4392 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n174_1), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n175), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n176_1) );
  AND2X2 AND2X2_4393 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n177_1), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n173), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n178) );
  AND2X2 AND2X2_4394 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n167), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n180_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n181_1) );
  AND2X2 AND2X2_4395 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n166_1), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n179), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n182) );
  AND2X2 AND2X2_4396 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__7_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n186) );
  AND2X2 AND2X2_4397 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n187_1), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n185), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n188_1) );
  AND2X2 AND2X2_4398 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n124), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n188_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n189) );
  AND2X2 AND2X2_4399 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n104), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n190), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n191_1) );
  AND2X2 AND2X2_44 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n85), .B(AES_CORE_CONTROL_UNIT__abc_15841_n144), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n145) );
  AND2X2 AND2X2_440 ( .A(AES_CORE_DATAPATH__abc_16259_n2786_bF_buf1), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_72_), .Y(AES_CORE_DATAPATH__abc_16259_n3159) );
  AND2X2 AND2X2_4400 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n192_1), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n147_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n193) );
  AND2X2 AND2X2_4401 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n195_1), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n196), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n197_1) );
  AND2X2 AND2X2_4402 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__6_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n198_1) );
  AND2X2 AND2X2_4403 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n202), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n201_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n203_1) );
  AND2X2 AND2X2_4404 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n200_1), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n204_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n205) );
  AND2X2 AND2X2_4405 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n207_1), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n208_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n209) );
  AND2X2 AND2X2_4406 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n156_1), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n203_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n210_1) );
  AND2X2 AND2X2_4407 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n152), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n199), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n211_1) );
  AND2X2 AND2X2_4408 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n213), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n206), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n214_1) );
  AND2X2 AND2X2_4409 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n216), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n217), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n218_1) );
  AND2X2 AND2X2_441 ( .A(AES_CORE_DATAPATH__abc_16259_n2789_bF_buf1), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_40_), .Y(AES_CORE_DATAPATH__abc_16259_n3160) );
  AND2X2 AND2X2_4410 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n215_1), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n219_1), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_1_) );
  AND2X2 AND2X2_4411 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n221_1), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n223), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n224_1) );
  AND2X2 AND2X2_4412 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n224_1), .B(AES_CORE_DATAPATH_MIX_COL_col_2__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n225_1) );
  AND2X2 AND2X2_4413 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n226), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n227_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n228_1) );
  AND2X2 AND2X2_4414 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n230), .B(AES_CORE_DATAPATH_MIX_COL_col_1__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n231) );
  AND2X2 AND2X2_4415 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n232), .B(AES_CORE_DATAPATH_MIX_COL_col_3__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n233) );
  AND2X2 AND2X2_4416 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n229), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n235), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n236) );
  AND2X2 AND2X2_4417 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n228_1), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n234), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n237) );
  AND2X2 AND2X2_4418 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__0_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n240) );
  AND2X2 AND2X2_4419 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n241), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n239), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n242) );
  AND2X2 AND2X2_442 ( .A(AES_CORE_DATAPATH__abc_16259_n3163), .B(AES_CORE_DATAPATH__abc_16259_n3157), .Y(AES_CORE_DATAPATH__abc_16259_n3164) );
  AND2X2 AND2X2_4420 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n109_1), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n160_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n244) );
  AND2X2 AND2X2_4421 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n243), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n246), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n247) );
  AND2X2 AND2X2_4422 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n102), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n248), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n249) );
  AND2X2 AND2X2_4423 ( .A(AES_CORE_DATAPATH_MIX_COL_col_3__7_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n250) );
  AND2X2 AND2X2_4424 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n251), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n203_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n252) );
  AND2X2 AND2X2_4425 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n254), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n253), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n255) );
  AND2X2 AND2X2_4426 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n199), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n255), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n256) );
  AND2X2 AND2X2_4427 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n194_1), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n257), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n258) );
  AND2X2 AND2X2_4428 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n259), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n260), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n261) );
  AND2X2 AND2X2_4429 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n209), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n261), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n262) );
  AND2X2 AND2X2_443 ( .A(AES_CORE_DATAPATH__abc_16259_n2837_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__8_), .Y(AES_CORE_DATAPATH__abc_16259_n3166) );
  AND2X2 AND2X2_4430 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n245), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n188_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n266) );
  AND2X2 AND2X2_4431 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n192_1), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n242), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n267) );
  AND2X2 AND2X2_4432 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n265), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n269), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n270) );
  AND2X2 AND2X2_4433 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n272), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n274), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_2_) );
  AND2X2 AND2X2_4434 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n276), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n278), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n279) );
  AND2X2 AND2X2_4435 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n107), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n279), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n280) );
  AND2X2 AND2X2_4436 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n281), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n282), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n283) );
  AND2X2 AND2X2_4437 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n285), .B(AES_CORE_DATAPATH_MIX_COL_col_1__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n286) );
  AND2X2 AND2X2_4438 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n287), .B(AES_CORE_DATAPATH_MIX_COL_col_3__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n288) );
  AND2X2 AND2X2_4439 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n289), .B(AES_CORE_DATAPATH_MIX_COL_col_2__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n290) );
  AND2X2 AND2X2_444 ( .A(AES_CORE_DATAPATH__abc_16259_n2887_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__8_), .Y(AES_CORE_DATAPATH__abc_16259_n3168) );
  AND2X2 AND2X2_4440 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n292), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n291), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n293) );
  AND2X2 AND2X2_4441 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n284), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n295), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n296) );
  AND2X2 AND2X2_4442 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n283), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n294), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n297) );
  AND2X2 AND2X2_4443 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n300), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n301), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n302) );
  AND2X2 AND2X2_4444 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n251), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n115_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n304) );
  AND2X2 AND2X2_4445 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n101), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n255), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n305) );
  AND2X2 AND2X2_4446 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n307), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n303), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n308) );
  AND2X2 AND2X2_4447 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n268), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n306), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n310) );
  AND2X2 AND2X2_4448 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n247), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n302), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n311) );
  AND2X2 AND2X2_4449 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n309), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n313), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n314) );
  AND2X2 AND2X2_445 ( .A(AES_CORE_DATAPATH__abc_16259_n2830_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__8_), .Y(AES_CORE_DATAPATH__abc_16259_n3169) );
  AND2X2 AND2X2_4450 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__1_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n316) );
  AND2X2 AND2X2_4451 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n317), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n315), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n318) );
  AND2X2 AND2X2_4452 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n173), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n222_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n320) );
  AND2X2 AND2X2_4453 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n322), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n319), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n323) );
  AND2X2 AND2X2_4454 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n326), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n325), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n327) );
  AND2X2 AND2X2_4455 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n124), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n321), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n328) );
  AND2X2 AND2X2_4456 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n147_1), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n318), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n329) );
  AND2X2 AND2X2_4457 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n324), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n331), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n332) );
  AND2X2 AND2X2_4458 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n334), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n335), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n336) );
  AND2X2 AND2X2_4459 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n333), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n337), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_3_) );
  AND2X2 AND2X2_446 ( .A(AES_CORE_DATAPATH__abc_16259_n3171), .B(AES_CORE_DATAPATH__abc_16259_n3172_1), .Y(_auto_iopadmap_cc_313_execute_26949_8_) );
  AND2X2 AND2X2_4460 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n339), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n341), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n342) );
  AND2X2 AND2X2_4461 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n107), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n342), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n343) );
  AND2X2 AND2X2_4462 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n344), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n345), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n346) );
  AND2X2 AND2X2_4463 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n349), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n351), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n352) );
  AND2X2 AND2X2_4464 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n353), .B(AES_CORE_DATAPATH_MIX_COL_col_2__4_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n354) );
  AND2X2 AND2X2_4465 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n352), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n355), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n356) );
  AND2X2 AND2X2_4466 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n347), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n358), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n359) );
  AND2X2 AND2X2_4467 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n346), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n357), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n360) );
  AND2X2 AND2X2_4468 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n277), .B(AES_CORE_DATAPATH_MIX_COL_col_2__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n363) );
  AND2X2 AND2X2_4469 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n364), .B(AES_CORE_DATAPATH_MIX_COL_col_0__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n365) );
  AND2X2 AND2X2_447 ( .A(AES_CORE_DATAPATH__abc_16259_n2855_bF_buf1), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_8_), .Y(AES_CORE_DATAPATH__abc_16259_n3175) );
  AND2X2 AND2X2_4470 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n369), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n367), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n370) );
  AND2X2 AND2X2_4471 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n171), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n203_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n371) );
  AND2X2 AND2X2_4472 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n177_1), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n199), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n372) );
  AND2X2 AND2X2_4473 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n330), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n373), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n374) );
  AND2X2 AND2X2_4474 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n375), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n376), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n377) );
  AND2X2 AND2X2_4475 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n323), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n377), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n378) );
  AND2X2 AND2X2_4476 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n381), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n382), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n383) );
  AND2X2 AND2X2_4477 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n384), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n380), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n385) );
  AND2X2 AND2X2_4478 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n388), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n387), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n389) );
  AND2X2 AND2X2_4479 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n390), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n391), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n392) );
  AND2X2 AND2X2_448 ( .A(AES_CORE_DATAPATH__abc_16259_n2857_bF_buf1), .B(AES_CORE_DATAPATH_MIX_COL_col_1__0_), .Y(AES_CORE_DATAPATH__abc_16259_n3176) );
  AND2X2 AND2X2_4480 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n386), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n393), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n394) );
  AND2X2 AND2X2_4481 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n396), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n397), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n398) );
  AND2X2 AND2X2_4482 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n395), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n399), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_4_) );
  AND2X2 AND2X2_4483 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n132), .B(AES_CORE_DATAPATH_MIX_COL_col_2__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n401) );
  AND2X2 AND2X2_4484 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n141), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n135), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n402) );
  AND2X2 AND2X2_4485 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n350), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n405), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n406) );
  AND2X2 AND2X2_4486 ( .A(AES_CORE_DATAPATH_MIX_COL_col_3__4_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__4_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n407) );
  AND2X2 AND2X2_4487 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n404), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n409), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n410) );
  AND2X2 AND2X2_4488 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n403), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n408), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n411) );
  AND2X2 AND2X2_4489 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__3_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n415) );
  AND2X2 AND2X2_449 ( .A(AES_CORE_DATAPATH__abc_16259_n3174), .B(AES_CORE_DATAPATH__abc_16259_n3178_1), .Y(AES_CORE_DATAPATH__abc_16259_n3179) );
  AND2X2 AND2X2_4490 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n416), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n414), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n417) );
  AND2X2 AND2X2_4491 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n418), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n188_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n419) );
  AND2X2 AND2X2_4492 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n192_1), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n417), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n420) );
  AND2X2 AND2X2_4493 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n423), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n422), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n424) );
  AND2X2 AND2X2_4494 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n257), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n234), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n426) );
  AND2X2 AND2X2_4495 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n261), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n235), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n427) );
  AND2X2 AND2X2_4496 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n425), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n429), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n430) );
  AND2X2 AND2X2_4497 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n428), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n370), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n433) );
  AND2X2 AND2X2_4498 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n389), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n424), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n434) );
  AND2X2 AND2X2_4499 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n431), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n436), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n437) );
  AND2X2 AND2X2_45 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n85), .B(AES_CORE_CONTROL_UNIT_state_8_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n148) );
  AND2X2 AND2X2_450 ( .A(_auto_iopadmap_cc_313_execute_26949_8_), .B(AES_CORE_DATAPATH__abc_16259_n3179), .Y(AES_CORE_DATAPATH__abc_16259_n3182) );
  AND2X2 AND2X2_4500 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n435), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n432), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n439) );
  AND2X2 AND2X2_4501 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n430), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n421), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n440) );
  AND2X2 AND2X2_4502 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n442), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n438), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_5_) );
  AND2X2 AND2X2_4503 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n444), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n445), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n446) );
  AND2X2 AND2X2_4504 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n446), .B(AES_CORE_DATAPATH_MIX_COL_col_1__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n447) );
  AND2X2 AND2X2_4505 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n448), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n449), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n450) );
  AND2X2 AND2X2_4506 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n451), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n452), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n453) );
  AND2X2 AND2X2_4507 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n457), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n454), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_6_) );
  AND2X2 AND2X2_4508 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n355), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n405), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n460) );
  AND2X2 AND2X2_4509 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__4_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__4_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n461) );
  AND2X2 AND2X2_451 ( .A(AES_CORE_DATAPATH_last_round_pp2_bF_buf0), .B(AES_CORE_DATAPATH_MIX_COL_col_1__0_), .Y(AES_CORE_DATAPATH__abc_16259_n3185_1) );
  AND2X2 AND2X2_4510 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n289), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n251), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n463) );
  AND2X2 AND2X2_4511 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n292), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n255), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n464) );
  AND2X2 AND2X2_4512 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n467), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n468), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n469) );
  AND2X2 AND2X2_4513 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n473), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n470), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n474) );
  AND2X2 AND2X2_4514 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n475), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n459), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n476) );
  AND2X2 AND2X2_4515 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n474), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n477) );
  AND2X2 AND2X2_4516 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n479), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n480), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n481) );
  AND2X2 AND2X2_4517 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n482), .B(AES_CORE_DATAPATH_MIX_COL_col_2__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n483) );
  AND2X2 AND2X2_4518 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n481), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n190), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n484) );
  AND2X2 AND2X2_4519 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n488), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n486), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_7_) );
  AND2X2 AND2X2_452 ( .A(AES_CORE_DATAPATH__abc_16259_n2798_bF_buf1), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_8_), .Y(AES_CORE_DATAPATH__abc_16259_n3186) );
  AND2X2 AND2X2_4520 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n353), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n462), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n491) );
  AND2X2 AND2X2_4521 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n471), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n352), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n492) );
  AND2X2 AND2X2_4522 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n495), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n496), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n497) );
  AND2X2 AND2X2_4523 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n500), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n498), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_7_) );
  AND2X2 AND2X2_4524 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n502), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n503), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n504) );
  AND2X2 AND2X2_4525 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n245), .B(AES_CORE_DATAPATH_MIX_COL_col_3__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n505) );
  AND2X2 AND2X2_4526 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n242), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n98), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n506) );
  AND2X2 AND2X2_4527 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n509), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n511), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_8_) );
  AND2X2 AND2X2_4528 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n514), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n515), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n516) );
  AND2X2 AND2X2_4529 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n513), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n517), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n518) );
  AND2X2 AND2X2_453 ( .A(AES_CORE_DATAPATH__abc_16259_n3184), .B(AES_CORE_DATAPATH__abc_16259_n3188), .Y(AES_CORE_DATAPATH__abc_16259_n3189) );
  AND2X2 AND2X2_4530 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_8_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n516), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n519) );
  AND2X2 AND2X2_4531 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n521), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n522), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n523) );
  AND2X2 AND2X2_4532 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n524), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n504), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n525) );
  AND2X2 AND2X2_4533 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n510), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n523), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n526) );
  AND2X2 AND2X2_4534 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n321), .B(AES_CORE_DATAPATH_MIX_COL_col_3__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n528) );
  AND2X2 AND2X2_4535 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n318), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n175), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n529) );
  AND2X2 AND2X2_4536 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n527), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n531), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n532) );
  AND2X2 AND2X2_4537 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n533), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n534), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n535) );
  AND2X2 AND2X2_4538 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n156_1), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n251), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n537) );
  AND2X2 AND2X2_4539 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n152), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n255), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n538) );
  AND2X2 AND2X2_454 ( .A(AES_CORE_DATAPATH__abc_16259_n3189), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf11), .Y(AES_CORE_DATAPATH__abc_16259_n3190) );
  AND2X2 AND2X2_4540 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n539), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n535), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n540) );
  AND2X2 AND2X2_4541 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n541), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_9_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n542) );
  AND2X2 AND2X2_4542 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n544), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n545), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n546) );
  AND2X2 AND2X2_4543 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n368), .B(AES_CORE_DATAPATH_MIX_COL_col_3__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n547) );
  AND2X2 AND2X2_4544 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n366), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n230), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n548) );
  AND2X2 AND2X2_4545 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n551), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n553), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_10_) );
  AND2X2 AND2X2_4546 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n556), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n557), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n558) );
  AND2X2 AND2X2_4547 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n561), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n559), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_10_) );
  AND2X2 AND2X2_4548 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n418), .B(AES_CORE_DATAPATH_MIX_COL_col_3__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n563) );
  AND2X2 AND2X2_4549 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n417), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n285), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n564) );
  AND2X2 AND2X2_455 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf3), .B(AES_CORE_DATAPATH_col_3__8_), .Y(AES_CORE_DATAPATH__abc_16259_n3191) );
  AND2X2 AND2X2_4550 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n567), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n568), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n569) );
  AND2X2 AND2X2_4551 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n510), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n570), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n571) );
  AND2X2 AND2X2_4552 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n504), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n569), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n572) );
  AND2X2 AND2X2_4553 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n574), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n566), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n575) );
  AND2X2 AND2X2_4554 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n573), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n565), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n576) );
  AND2X2 AND2X2_4555 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n327), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n373), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n578) );
  AND2X2 AND2X2_4556 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n314), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n377), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n579) );
  AND2X2 AND2X2_4557 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n580), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_11_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n581) );
  AND2X2 AND2X2_4558 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n583), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n584), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n585) );
  AND2X2 AND2X2_4559 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n585), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n582), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n586) );
  AND2X2 AND2X2_456 ( .A(AES_CORE_DATAPATH__abc_16259_n3194), .B(AES_CORE_DATAPATH__abc_16259_n3196), .Y(AES_CORE_DATAPATH__abc_16259_n3197) );
  AND2X2 AND2X2_4560 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n462), .B(AES_CORE_DATAPATH_MIX_COL_col_3__4_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n588) );
  AND2X2 AND2X2_4561 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n471), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n350), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n589) );
  AND2X2 AND2X2_4562 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n592), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n593), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n594) );
  AND2X2 AND2X2_4563 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n510), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n595), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n596) );
  AND2X2 AND2X2_4564 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n504), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n594), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n597) );
  AND2X2 AND2X2_4565 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n599), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n591), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n600) );
  AND2X2 AND2X2_4566 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n598), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n590), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n601) );
  AND2X2 AND2X2_4567 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n603), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n604), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n605) );
  AND2X2 AND2X2_4568 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n608), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n609), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n610) );
  AND2X2 AND2X2_4569 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n606), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n611), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_12_) );
  AND2X2 AND2X2_457 ( .A(AES_CORE_DATAPATH__abc_16259_n2782_bF_buf0), .B(AES_CORE_DATAPATH_col_3__9_), .Y(AES_CORE_DATAPATH__abc_16259_n3198) );
  AND2X2 AND2X2_4570 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n613), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n614), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n615) );
  AND2X2 AND2X2_4571 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n137), .B(AES_CORE_DATAPATH_MIX_COL_col_3__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n616) );
  AND2X2 AND2X2_4572 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n128), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n139), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n617) );
  AND2X2 AND2X2_4573 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n620), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n622), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_13_) );
  AND2X2 AND2X2_4574 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n625), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n626), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n627) );
  AND2X2 AND2X2_4575 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n629), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n630), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n631) );
  AND2X2 AND2X2_4576 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n628), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n632), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_13_) );
  AND2X2 AND2X2_4577 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n634), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n635), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n636) );
  AND2X2 AND2X2_4578 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n147_1), .B(AES_CORE_DATAPATH_MIX_COL_col_3__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n638) );
  AND2X2 AND2X2_4579 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n124), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n196), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n639) );
  AND2X2 AND2X2_458 ( .A(AES_CORE_DATAPATH__abc_16259_n2786_bF_buf0), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_73_), .Y(AES_CORE_DATAPATH__abc_16259_n3199_1) );
  AND2X2 AND2X2_4580 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n641), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n637), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n642) );
  AND2X2 AND2X2_4581 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n640), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n636), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n643) );
  AND2X2 AND2X2_4582 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n647), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n646), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n648) );
  AND2X2 AND2X2_4583 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n651), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n649), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_14_) );
  AND2X2 AND2X2_4584 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n653), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n654), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n655) );
  AND2X2 AND2X2_4585 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n656), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n657), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n658) );
  AND2X2 AND2X2_4586 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n659), .B(AES_CORE_DATAPATH_MIX_COL_col_0__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n660) );
  AND2X2 AND2X2_4587 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n658), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n104), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n661) );
  AND2X2 AND2X2_4588 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n664), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n666), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n667) );
  AND2X2 AND2X2_4589 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n669), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n670), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n671) );
  AND2X2 AND2X2_459 ( .A(AES_CORE_DATAPATH__abc_16259_n2789_bF_buf0), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_41_), .Y(AES_CORE_DATAPATH__abc_16259_n3200) );
  AND2X2 AND2X2_4590 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n674), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n672), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_15_) );
  AND2X2 AND2X2_4591 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n190), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n248), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n676) );
  AND2X2 AND2X2_4592 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__7_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n677) );
  AND2X2 AND2X2_4593 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n115_1), .B(AES_CORE_DATAPATH_MIX_COL_col_0__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n679) );
  AND2X2 AND2X2_4594 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n101), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n160_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n680) );
  AND2X2 AND2X2_4595 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n682), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n678), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n683) );
  AND2X2 AND2X2_4596 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n681), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n684), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n685) );
  AND2X2 AND2X2_4597 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n687), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n156_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n688) );
  AND2X2 AND2X2_4598 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_16_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n152), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n689) );
  AND2X2 AND2X2_4599 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n552), .B(AES_CORE_DATAPATH_MIX_COL_col_3__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n691) );
  AND2X2 AND2X2_46 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n107), .B(AES_CORE_CONTROL_UNIT_state_12_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n149) );
  AND2X2 AND2X2_460 ( .A(AES_CORE_DATAPATH__abc_16259_n3203), .B(AES_CORE_DATAPATH__abc_16259_n3197), .Y(AES_CORE_DATAPATH__abc_16259_n3204) );
  AND2X2 AND2X2_4600 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n546), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n175), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n692) );
  AND2X2 AND2X2_4601 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n97_1), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n109_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n695) );
  AND2X2 AND2X2_4602 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__0_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n696) );
  AND2X2 AND2X2_4603 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n698), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n684), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n699) );
  AND2X2 AND2X2_4604 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n697), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n678), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n700) );
  AND2X2 AND2X2_4605 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n702), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n694), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n703) );
  AND2X2 AND2X2_4606 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n701), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n693), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n704) );
  AND2X2 AND2X2_4607 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n707), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n708), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_17_) );
  AND2X2 AND2X2_4608 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n174_1), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n173), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n710) );
  AND2X2 AND2X2_4609 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__1_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n711) );
  AND2X2 AND2X2_461 ( .A(AES_CORE_DATAPATH__abc_16259_n2837_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__9_), .Y(AES_CORE_DATAPATH__abc_16259_n3206_1) );
  AND2X2 AND2X2_4610 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n570), .B(AES_CORE_DATAPATH_MIX_COL_col_3__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n713) );
  AND2X2 AND2X2_4611 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n569), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n230), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n714) );
  AND2X2 AND2X2_4612 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n719), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n716), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_18_) );
  AND2X2 AND2X2_4613 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n723), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n722), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_18_) );
  AND2X2 AND2X2_4614 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n232), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n364), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n725) );
  AND2X2 AND2X2_4615 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__2_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n726) );
  AND2X2 AND2X2_4616 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n684), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n727), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n728) );
  AND2X2 AND2X2_4617 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n729), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n678), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n730) );
  AND2X2 AND2X2_4618 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n733), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n732), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n734) );
  AND2X2 AND2X2_4619 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n731), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n734), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n735) );
  AND2X2 AND2X2_462 ( .A(AES_CORE_DATAPATH__abc_16259_n2887_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__9_), .Y(AES_CORE_DATAPATH__abc_16259_n3208) );
  AND2X2 AND2X2_4620 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n736), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n737), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_19_) );
  AND2X2 AND2X2_4621 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n739), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n741), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_19_) );
  AND2X2 AND2X2_4622 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n287), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n291), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n743) );
  AND2X2 AND2X2_4623 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__3_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n744) );
  AND2X2 AND2X2_4624 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n684), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n745), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n746) );
  AND2X2 AND2X2_4625 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n747), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n748), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n749) );
  AND2X2 AND2X2_4626 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n353), .B(AES_CORE_DATAPATH_MIX_COL_col_0__4_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n751) );
  AND2X2 AND2X2_4627 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n352), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n405), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n752) );
  AND2X2 AND2X2_4628 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n750), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n754), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n755) );
  AND2X2 AND2X2_4629 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n749), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n753), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n756) );
  AND2X2 AND2X2_463 ( .A(AES_CORE_DATAPATH__abc_16259_n2830_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__9_), .Y(AES_CORE_DATAPATH__abc_16259_n3209) );
  AND2X2 AND2X2_4630 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n759), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n760), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_20_) );
  AND2X2 AND2X2_4631 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n348), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n355), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n762) );
  AND2X2 AND2X2_4632 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__4_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__4_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n763) );
  AND2X2 AND2X2_4633 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n764), .B(AES_CORE_DATAPATH_MIX_COL_col_0__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n765) );
  AND2X2 AND2X2_4634 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n766), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n767), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n768) );
  AND2X2 AND2X2_4635 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n771), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n769), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n772) );
  AND2X2 AND2X2_4636 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n775), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n774), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_21_) );
  AND2X2 AND2X2_4637 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n777), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n778), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n779) );
  AND2X2 AND2X2_4638 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n780), .B(AES_CORE_DATAPATH_MIX_COL_col_1__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n781) );
  AND2X2 AND2X2_4639 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n779), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n195_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n782) );
  AND2X2 AND2X2_464 ( .A(AES_CORE_DATAPATH__abc_16259_n3211), .B(AES_CORE_DATAPATH__abc_16259_n3212_1), .Y(_auto_iopadmap_cc_313_execute_26949_9_) );
  AND2X2 AND2X2_4640 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n784), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n481), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n785) );
  AND2X2 AND2X2_4641 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n783), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n482), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n786) );
  AND2X2 AND2X2_4642 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n475), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n788), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n789) );
  AND2X2 AND2X2_4643 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n474), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_22_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n790) );
  AND2X2 AND2X2_4644 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n121), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n195_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n792) );
  AND2X2 AND2X2_4645 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__6_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n793) );
  AND2X2 AND2X2_4646 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n107), .B(AES_CORE_DATAPATH_MIX_COL_col_1__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n795) );
  AND2X2 AND2X2_4647 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n106), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n248), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n796) );
  AND2X2 AND2X2_4648 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n798), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n794), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n799) );
  AND2X2 AND2X2_4649 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n800), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n801), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n802) );
  AND2X2 AND2X2_465 ( .A(AES_CORE_DATAPATH__abc_16259_n2855_bF_buf0), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_9_), .Y(AES_CORE_DATAPATH__abc_16259_n3215) );
  AND2X2 AND2X2_4650 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n805), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n804), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_23_) );
  AND2X2 AND2X2_4651 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n698), .B(AES_CORE_DATAPATH_MIX_COL_col_0__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n807) );
  AND2X2 AND2X2_4652 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n697), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n160_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n808) );
  AND2X2 AND2X2_4653 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n810), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n658), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n811) );
  AND2X2 AND2X2_4654 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n809), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n659), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n812) );
  AND2X2 AND2X2_4655 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n814), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n517), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n815) );
  AND2X2 AND2X2_4656 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_24_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n516), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n816) );
  AND2X2 AND2X2_4657 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n109_1), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n98), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n818) );
  AND2X2 AND2X2_4658 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__0_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n819) );
  AND2X2 AND2X2_4659 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n659), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n820), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n821) );
  AND2X2 AND2X2_466 ( .A(AES_CORE_DATAPATH__abc_16259_n2857_bF_buf0), .B(AES_CORE_DATAPATH_MIX_COL_col_1__1_), .Y(AES_CORE_DATAPATH__abc_16259_n3216_1) );
  AND2X2 AND2X2_4660 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n822), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n823), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n824) );
  AND2X2 AND2X2_4661 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n827), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n826), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n828) );
  AND2X2 AND2X2_4662 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n825), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n828), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n829) );
  AND2X2 AND2X2_4663 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n830), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n831), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n832) );
  AND2X2 AND2X2_4664 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n834), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n835), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_25_) );
  AND2X2 AND2X2_4665 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n173), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n175), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n837) );
  AND2X2 AND2X2_4666 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__1_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n838) );
  AND2X2 AND2X2_4667 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n839), .B(AES_CORE_DATAPATH_MIX_COL_col_0__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n840) );
  AND2X2 AND2X2_4668 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n845), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n846), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n847) );
  AND2X2 AND2X2_4669 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n560), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n847), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n849) );
  AND2X2 AND2X2_467 ( .A(AES_CORE_DATAPATH__abc_16259_n3214_1), .B(AES_CORE_DATAPATH__abc_16259_n3218), .Y(AES_CORE_DATAPATH__abc_16259_n3219) );
  AND2X2 AND2X2_4670 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n558), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_26_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n850) );
  AND2X2 AND2X2_4671 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n364), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n230), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n852) );
  AND2X2 AND2X2_4672 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__2_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n853) );
  AND2X2 AND2X2_4673 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n659), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n854), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n855) );
  AND2X2 AND2X2_4674 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n856), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n857), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n858) );
  AND2X2 AND2X2_4675 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n418), .B(AES_CORE_DATAPATH_MIX_COL_col_1__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n860) );
  AND2X2 AND2X2_4676 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n417), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n287), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n861) );
  AND2X2 AND2X2_4677 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n859), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n863), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n864) );
  AND2X2 AND2X2_4678 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n858), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n862), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n865) );
  AND2X2 AND2X2_4679 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n869), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n867), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_27_) );
  AND2X2 AND2X2_468 ( .A(_auto_iopadmap_cc_313_execute_26949_9_), .B(AES_CORE_DATAPATH__abc_16259_n3219), .Y(AES_CORE_DATAPATH__abc_16259_n3222) );
  AND2X2 AND2X2_4680 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n471), .B(AES_CORE_DATAPATH_MIX_COL_col_1__4_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n871) );
  AND2X2 AND2X2_4681 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n462), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n348), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n872) );
  AND2X2 AND2X2_4682 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n291), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n285), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n875) );
  AND2X2 AND2X2_4683 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__3_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n876) );
  AND2X2 AND2X2_4684 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n659), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n877), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n878) );
  AND2X2 AND2X2_4685 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n879), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n880), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n881) );
  AND2X2 AND2X2_4686 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n882), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n874), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n883) );
  AND2X2 AND2X2_4687 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n881), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n873), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n884) );
  AND2X2 AND2X2_4688 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n887), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n888), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_28_) );
  AND2X2 AND2X2_4689 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n355), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n350), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n890) );
  AND2X2 AND2X2_469 ( .A(AES_CORE_DATAPATH_last_round_pp2_bF_buf4), .B(AES_CORE_DATAPATH_MIX_COL_col_1__1_), .Y(AES_CORE_DATAPATH__abc_16259_n3225) );
  AND2X2 AND2X2_4690 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__4_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__4_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n891) );
  AND2X2 AND2X2_4691 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n637), .B(AES_CORE_DATAPATH_MIX_COL_col_2__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n894) );
  AND2X2 AND2X2_4692 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n636), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n135), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n895) );
  AND2X2 AND2X2_4693 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n899), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n897), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n900) );
  AND2X2 AND2X2_4694 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n902), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n903), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_29_) );
  AND2X2 AND2X2_4695 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n139), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n135), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n905) );
  AND2X2 AND2X2_4696 ( .A(AES_CORE_DATAPATH_MIX_COL_col_3__5_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n906) );
  AND2X2 AND2X2_4697 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n907), .B(AES_CORE_DATAPATH_MIX_COL_col_1__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n908) );
  AND2X2 AND2X2_4698 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n909), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n195_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n910) );
  AND2X2 AND2X2_4699 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n913), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n914), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_30_) );
  AND2X2 AND2X2_47 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n85), .B(AES_CORE_CONTROL_UNIT_state_4_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n151) );
  AND2X2 AND2X2_470 ( .A(AES_CORE_DATAPATH__abc_16259_n2798_bF_buf0), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_9_), .Y(AES_CORE_DATAPATH__abc_16259_n3226) );
  AND2X2 AND2X2_4700 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n918), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n917), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_30_) );
  AND2X2 AND2X2_4701 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n504), .B(AES_CORE_DATAPATH_MIX_COL_col_2__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n920) );
  AND2X2 AND2X2_4702 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n510), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n190), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n921) );
  AND2X2 AND2X2_4703 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n924), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n925), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n926) );
  AND2X2 AND2X2_4704 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n673), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n926), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n928) );
  AND2X2 AND2X2_4705 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_31_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n671), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n929) );
  AND2X2 AND2X2_4706 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n50), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n51_1) );
  AND2X2 AND2X2_4707 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n52), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n53_1) );
  AND2X2 AND2X2_4708 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n57), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n59), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n60) );
  AND2X2 AND2X2_4709 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n55), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n61), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n62) );
  AND2X2 AND2X2_471 ( .A(AES_CORE_DATAPATH__abc_16259_n3224), .B(AES_CORE_DATAPATH__abc_16259_n3228_1), .Y(AES_CORE_DATAPATH__abc_16259_n3229) );
  AND2X2 AND2X2_4710 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n54_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n60), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n63) );
  AND2X2 AND2X2_4711 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n64), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf2), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n65) );
  AND2X2 AND2X2_4712 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n54_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n67), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n68) );
  AND2X2 AND2X2_4713 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n55), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n69) );
  AND2X2 AND2X2_4714 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n70), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n71_1) );
  AND2X2 AND2X2_4715 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n73), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n72), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n74) );
  AND2X2 AND2X2_4716 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n75), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n66_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n76) );
  AND2X2 AND2X2_4717 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n78), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n80), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n81) );
  AND2X2 AND2X2_4718 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n70), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n83) );
  AND2X2 AND2X2_4719 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n73), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n56), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n84_1) );
  AND2X2 AND2X2_472 ( .A(AES_CORE_DATAPATH__abc_16259_n3229), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf10), .Y(AES_CORE_DATAPATH__abc_16259_n3230_1) );
  AND2X2 AND2X2_4720 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n85), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf7), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n86_1) );
  AND2X2 AND2X2_4721 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n87), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n82), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_5_) );
  AND2X2 AND2X2_4722 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n54_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n89) );
  AND2X2 AND2X2_4723 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n55), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n56), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n90) );
  AND2X2 AND2X2_4724 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n73), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n66_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n94_1) );
  AND2X2 AND2X2_4725 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n96), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n97_1) );
  AND2X2 AND2X2_4726 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n95), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n79), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n98) );
  AND2X2 AND2X2_4727 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n100), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n101_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n102) );
  AND2X2 AND2X2_4728 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n102), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n66_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n103) );
  AND2X2 AND2X2_4729 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n61), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n104_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n105) );
  AND2X2 AND2X2_473 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf2), .B(AES_CORE_DATAPATH_col_3__9_), .Y(AES_CORE_DATAPATH__abc_16259_n3231) );
  AND2X2 AND2X2_4730 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n60), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n106) );
  AND2X2 AND2X2_4731 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n73), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n107), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n108) );
  AND2X2 AND2X2_4732 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n109), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n70), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n110) );
  AND2X2 AND2X2_4733 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n75), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n116) );
  AND2X2 AND2X2_4734 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n117), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n118), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n119) );
  AND2X2 AND2X2_4735 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n85), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n121_1) );
  AND2X2 AND2X2_4736 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n122), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n123), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n124) );
  AND2X2 AND2X2_4737 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n120), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n125), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n126_1) );
  AND2X2 AND2X2_4738 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n128), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n129), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n130) );
  AND2X2 AND2X2_4739 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n131), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n79), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n132) );
  AND2X2 AND2X2_474 ( .A(AES_CORE_DATAPATH__abc_16259_n3234), .B(AES_CORE_DATAPATH__abc_16259_n3236_1), .Y(AES_CORE_DATAPATH__abc_16259_n3237) );
  AND2X2 AND2X2_4740 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n130), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n133) );
  AND2X2 AND2X2_4741 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n92), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n135), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n136) );
  AND2X2 AND2X2_4742 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n107), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n66_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n138) );
  AND2X2 AND2X2_4743 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n50), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf4), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n139_1) );
  AND2X2 AND2X2_4744 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n142), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n143_1) );
  AND2X2 AND2X2_4745 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n102), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n52), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n144) );
  AND2X2 AND2X2_4746 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n142), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n147) );
  AND2X2 AND2X2_4747 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n102), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n67), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n148_1) );
  AND2X2 AND2X2_4748 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n150_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n130), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n151_1) );
  AND2X2 AND2X2_4749 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n149), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n131), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n152_1) );
  AND2X2 AND2X2_475 ( .A(AES_CORE_DATAPATH__abc_16259_n2782_bF_buf4), .B(AES_CORE_DATAPATH_col_3__10_), .Y(AES_CORE_DATAPATH__abc_16259_n3238) );
  AND2X2 AND2X2_4750 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n154), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n146_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_3_) );
  AND2X2 AND2X2_4751 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n156) );
  AND2X2 AND2X2_4752 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n157) );
  AND2X2 AND2X2_4753 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n159), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n160) );
  AND2X2 AND2X2_4754 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n161), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n162) );
  AND2X2 AND2X2_4755 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n164) );
  AND2X2 AND2X2_4756 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n165), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n164), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n167) );
  AND2X2 AND2X2_4757 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n168), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n166_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n169) );
  AND2X2 AND2X2_4758 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n169), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n163), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n170) );
  AND2X2 AND2X2_4759 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n170), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n158), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n171) );
  AND2X2 AND2X2_476 ( .A(AES_CORE_DATAPATH__abc_16259_n2786_bF_buf4), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_74_), .Y(AES_CORE_DATAPATH__abc_16259_n3239_1) );
  AND2X2 AND2X2_4760 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_1_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n173) );
  AND2X2 AND2X2_4761 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n161), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n176_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n177) );
  AND2X2 AND2X2_4762 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n175), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n177), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n178) );
  AND2X2 AND2X2_4763 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n183), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n174), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n184) );
  AND2X2 AND2X2_4764 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n189_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n186), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n190_1) );
  AND2X2 AND2X2_4765 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n169), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n180), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n191) );
  AND2X2 AND2X2_4766 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n191), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n158), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n192) );
  AND2X2 AND2X2_4767 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n185), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n194), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n195) );
  AND2X2 AND2X2_4768 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n197), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n199), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n200) );
  AND2X2 AND2X2_4769 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n195), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n201), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n202) );
  AND2X2 AND2X2_477 ( .A(AES_CORE_DATAPATH__abc_16259_n2789_bF_buf4), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_42_), .Y(AES_CORE_DATAPATH__abc_16259_n3240) );
  AND2X2 AND2X2_4770 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n173), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n159), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n203) );
  AND2X2 AND2X2_4771 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n163), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n176_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n205) );
  AND2X2 AND2X2_4772 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n169), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n162), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n207) );
  AND2X2 AND2X2_4773 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n214), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n208), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n215) );
  AND2X2 AND2X2_4774 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n211), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n216), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n217) );
  AND2X2 AND2X2_4775 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n219), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n221), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n222) );
  AND2X2 AND2X2_4776 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n217), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n222), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n223) );
  AND2X2 AND2X2_4777 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n202), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n223), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n224) );
  AND2X2 AND2X2_4778 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n190_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n193), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n225) );
  AND2X2 AND2X2_4779 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n184), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n172), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n226) );
  AND2X2 AND2X2_478 ( .A(AES_CORE_DATAPATH__abc_16259_n3243_1), .B(AES_CORE_DATAPATH__abc_16259_n3237), .Y(AES_CORE_DATAPATH__abc_16259_n3244) );
  AND2X2 AND2X2_4780 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n230), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n229), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n231) );
  AND2X2 AND2X2_4781 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n233), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n234), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n235) );
  AND2X2 AND2X2_4782 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n228), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n235), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n236) );
  AND2X2 AND2X2_4783 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n158), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n159), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n238) );
  AND2X2 AND2X2_4784 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n156), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n239) );
  AND2X2 AND2X2_4785 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n241), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n242), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n243) );
  AND2X2 AND2X2_4786 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n215), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n245) );
  AND2X2 AND2X2_4787 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n245), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n244), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n246) );
  AND2X2 AND2X2_4788 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n247), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n248), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n249) );
  AND2X2 AND2X2_4789 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n231), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n200), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n253) );
  AND2X2 AND2X2_479 ( .A(AES_CORE_DATAPATH__abc_16259_n2837_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__10_), .Y(AES_CORE_DATAPATH__abc_16259_n3246) );
  AND2X2 AND2X2_4790 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n252), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n255), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n256) );
  AND2X2 AND2X2_4791 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n251), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n257), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n258) );
  AND2X2 AND2X2_4792 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n260), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n262), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n263) );
  AND2X2 AND2X2_4793 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n217), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n264), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n265) );
  AND2X2 AND2X2_4794 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n268), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n270), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n271) );
  AND2X2 AND2X2_4795 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n227), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n272), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n273) );
  AND2X2 AND2X2_4796 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n276), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n274), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n277) );
  AND2X2 AND2X2_4797 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n193), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n212), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n278) );
  AND2X2 AND2X2_4798 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n267), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n259), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n280) );
  AND2X2 AND2X2_4799 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n281) );
  AND2X2 AND2X2_48 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n107), .B(AES_CORE_CONTROL_UNIT_state_2_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n152) );
  AND2X2 AND2X2_480 ( .A(AES_CORE_DATAPATH__abc_16259_n2887_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__10_), .Y(AES_CORE_DATAPATH__abc_16259_n3248) );
  AND2X2 AND2X2_4800 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n193), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n284) );
  AND2X2 AND2X2_4801 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n287), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n180), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n288) );
  AND2X2 AND2X2_4802 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n288), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n289), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n290) );
  AND2X2 AND2X2_4803 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n286), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n291), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n292) );
  AND2X2 AND2X2_4804 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n296), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n294), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n297) );
  AND2X2 AND2X2_4805 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n298), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n299), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n300) );
  AND2X2 AND2X2_4806 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n172), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n302) );
  AND2X2 AND2X2_4807 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n302), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n301), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n303) );
  AND2X2 AND2X2_4808 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n304), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n305), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n306) );
  AND2X2 AND2X2_4809 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n308), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n309), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n310) );
  AND2X2 AND2X2_481 ( .A(AES_CORE_DATAPATH__abc_16259_n2830_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__10_), .Y(AES_CORE_DATAPATH__abc_16259_n3249) );
  AND2X2 AND2X2_4810 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n311), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n297), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n312) );
  AND2X2 AND2X2_4811 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n313), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n310), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n314) );
  AND2X2 AND2X2_4812 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n315), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n258), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n316) );
  AND2X2 AND2X2_4813 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n318), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n317), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n319) );
  AND2X2 AND2X2_4814 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n227), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n232), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n321) );
  AND2X2 AND2X2_4815 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n217), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n201), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n323) );
  AND2X2 AND2X2_4816 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n325), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n326), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n327) );
  AND2X2 AND2X2_4817 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n172), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n329) );
  AND2X2 AND2X2_4818 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n329), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n244), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n330) );
  AND2X2 AND2X2_4819 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n331), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n332), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n333) );
  AND2X2 AND2X2_482 ( .A(AES_CORE_DATAPATH__abc_16259_n3251), .B(AES_CORE_DATAPATH__abc_16259_n3252), .Y(_auto_iopadmap_cc_313_execute_26949_10_) );
  AND2X2 AND2X2_4820 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n334), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n336), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n337) );
  AND2X2 AND2X2_4821 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n313), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n338), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n339) );
  AND2X2 AND2X2_4822 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n297), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n337), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n340) );
  AND2X2 AND2X2_4823 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n342), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n343), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n344) );
  AND2X2 AND2X2_4824 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n288), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n345), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n346) );
  AND2X2 AND2X2_4825 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n193), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n347) );
  AND2X2 AND2X2_4826 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n351), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n349), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n352) );
  AND2X2 AND2X2_4827 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n354), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n355), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n356) );
  AND2X2 AND2X2_4828 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n212), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n358) );
  AND2X2 AND2X2_4829 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n361), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n359), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n362) );
  AND2X2 AND2X2_483 ( .A(AES_CORE_DATAPATH__abc_16259_n2855_bF_buf4), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_10_), .Y(AES_CORE_DATAPATH__abc_16259_n3255) );
  AND2X2 AND2X2_4830 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n365), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n364), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n366) );
  AND2X2 AND2X2_4831 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n363), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n367), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n368) );
  AND2X2 AND2X2_4832 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n195), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n264), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n369) );
  AND2X2 AND2X2_4833 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n217), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n271), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n370) );
  AND2X2 AND2X2_4834 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n369), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n370), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n371) );
  AND2X2 AND2X2_4835 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n373), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n374), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n375) );
  AND2X2 AND2X2_4836 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n372), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n375), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n376) );
  AND2X2 AND2X2_4837 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n215), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n378) );
  AND2X2 AND2X2_4838 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n378), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n301), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n379) );
  AND2X2 AND2X2_4839 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n380), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n381), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n382) );
  AND2X2 AND2X2_484 ( .A(AES_CORE_DATAPATH__abc_16259_n2857_bF_buf4), .B(AES_CORE_DATAPATH_MIX_COL_col_1__2_), .Y(AES_CORE_DATAPATH__abc_16259_n3256) );
  AND2X2 AND2X2_4840 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n231), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n263), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n386) );
  AND2X2 AND2X2_4841 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n385), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n388), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n389) );
  AND2X2 AND2X2_4842 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n384), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n390), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n391) );
  AND2X2 AND2X2_4843 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n393), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n394), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n395) );
  AND2X2 AND2X2_4844 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n396), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n397), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n398) );
  AND2X2 AND2X2_4845 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n392), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n399), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_7_) );
  AND2X2 AND2X2_4846 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n395), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n398), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n403) );
  AND2X2 AND2X2_4847 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n368), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n391), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n404) );
  AND2X2 AND2X2_4848 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n402), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n406), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n407) );
  AND2X2 AND2X2_4849 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n410), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n408), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_2_) );
  AND2X2 AND2X2_485 ( .A(AES_CORE_DATAPATH__abc_16259_n3254), .B(AES_CORE_DATAPATH__abc_16259_n3258), .Y(AES_CORE_DATAPATH__abc_16259_n3259_1) );
  AND2X2 AND2X2_4850 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n212), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n412) );
  AND2X2 AND2X2_4851 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n415), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n414), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n416) );
  AND2X2 AND2X2_4852 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n419), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n418), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n420) );
  AND2X2 AND2X2_4853 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n417), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n421), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n422) );
  AND2X2 AND2X2_4854 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n395), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n422), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n423) );
  AND2X2 AND2X2_4855 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n424), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n425), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n426) );
  AND2X2 AND2X2_4856 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n368), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n426), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n427) );
  AND2X2 AND2X2_4857 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n429), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n430), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n431) );
  AND2X2 AND2X2_4858 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n434), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n435), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n436) );
  AND2X2 AND2X2_4859 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n433), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n437), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_4_) );
  AND2X2 AND2X2_486 ( .A(_auto_iopadmap_cc_313_execute_26949_10_), .B(AES_CORE_DATAPATH__abc_16259_n3259_1), .Y(AES_CORE_DATAPATH__abc_16259_n3262) );
  AND2X2 AND2X2_4860 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n432), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n439), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_3_) );
  AND2X2 AND2X2_4861 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n441), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n442), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n443) );
  AND2X2 AND2X2_4862 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n445), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n444), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_3_) );
  AND2X2 AND2X2_4863 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n447), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n448), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n449) );
  AND2X2 AND2X2_4864 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_4_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n451) );
  AND2X2 AND2X2_4865 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n431), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n401), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n452) );
  AND2X2 AND2X2_4866 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n454), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n450), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_5_) );
  AND2X2 AND2X2_4867 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n457), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n456), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_6_) );
  AND2X2 AND2X2_4868 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n317), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n398), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n459) );
  AND2X2 AND2X2_4869 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n258), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n391), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n460) );
  AND2X2 AND2X2_487 ( .A(AES_CORE_DATAPATH_last_round_pp2_bF_buf3), .B(AES_CORE_DATAPATH_MIX_COL_col_1__2_), .Y(AES_CORE_DATAPATH__abc_16259_n3265_1) );
  AND2X2 AND2X2_4870 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n463), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n464), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_1_) );
  AND2X2 AND2X2_4871 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n467), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n466), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n468) );
  AND2X2 AND2X2_4872 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n126_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n469), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n470) );
  AND2X2 AND2X2_4873 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n472), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n473) );
  AND2X2 AND2X2_4874 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n469), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n474) );
  AND2X2 AND2X2_4875 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n471), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n475), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n476) );
  AND2X2 AND2X2_4876 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n468), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n476), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n477) );
  AND2X2 AND2X2_4877 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n478) );
  AND2X2 AND2X2_4878 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n470), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n479), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n480) );
  AND2X2 AND2X2_4879 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n483), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n482), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n484) );
  AND2X2 AND2X2_488 ( .A(AES_CORE_DATAPATH__abc_16259_n2798_bF_buf4), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_10_), .Y(AES_CORE_DATAPATH__abc_16259_n3266) );
  AND2X2 AND2X2_4880 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n486), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n487) );
  AND2X2 AND2X2_4881 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n469), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n488) );
  AND2X2 AND2X2_4882 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n485), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n489), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n490) );
  AND2X2 AND2X2_4883 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n494), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n492), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n495) );
  AND2X2 AND2X2_4884 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n472), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n114), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n497) );
  AND2X2 AND2X2_4885 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n498), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n496), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n499) );
  AND2X2 AND2X2_4886 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n499), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n495), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n500) );
  AND2X2 AND2X2_4887 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n491), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n500), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n501) );
  AND2X2 AND2X2_4888 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n502), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n503), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n504) );
  AND2X2 AND2X2_4889 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n505), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n481), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n506) );
  AND2X2 AND2X2_489 ( .A(AES_CORE_DATAPATH__abc_16259_n3264_1), .B(AES_CORE_DATAPATH__abc_16259_n3268_1), .Y(AES_CORE_DATAPATH__abc_16259_n3269) );
  AND2X2 AND2X2_4890 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n504), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n507), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n508) );
  AND2X2 AND2X2_4891 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n114), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n512) );
  AND2X2 AND2X2_4892 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n513), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n511), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n514) );
  AND2X2 AND2X2_4893 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n515), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n510), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n516) );
  AND2X2 AND2X2_4894 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n514), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n475), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n517) );
  AND2X2 AND2X2_4895 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n519), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n520), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n521) );
  AND2X2 AND2X2_4896 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n522), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n523), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n524) );
  AND2X2 AND2X2_4897 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n521), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n525), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n526) );
  AND2X2 AND2X2_4898 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n468), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n524), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n527) );
  AND2X2 AND2X2_4899 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n528), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n518), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n529) );
  AND2X2 AND2X2_49 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n142), .B(AES_CORE_CONTROL_UNIT__abc_15841_n84_1), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n154) );
  AND2X2 AND2X2_490 ( .A(AES_CORE_DATAPATH__abc_16259_n3269), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf9), .Y(AES_CORE_DATAPATH__abc_16259_n3270_1) );
  AND2X2 AND2X2_4900 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n521), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n510), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n530) );
  AND2X2 AND2X2_4901 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n530), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n479), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n531) );
  AND2X2 AND2X2_4902 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n532), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n478), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n533) );
  AND2X2 AND2X2_4903 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n534), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n490), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n535) );
  AND2X2 AND2X2_4904 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n536), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n537), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n538) );
  AND2X2 AND2X2_4905 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n538), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n491), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n539) );
  AND2X2 AND2X2_4906 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n543), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n544), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n545) );
  AND2X2 AND2X2_4907 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n541), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n546), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_stage1_1_) );
  AND2X2 AND2X2_4908 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n515), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n525), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n548) );
  AND2X2 AND2X2_4909 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n549) );
  AND2X2 AND2X2_491 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf1), .B(AES_CORE_DATAPATH_col_3__10_), .Y(AES_CORE_DATAPATH__abc_16259_n3271) );
  AND2X2 AND2X2_4910 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n551), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n549), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n552) );
  AND2X2 AND2X2_4911 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n553), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n554), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n555) );
  AND2X2 AND2X2_4912 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n557), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n559), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n560) );
  AND2X2 AND2X2_4913 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n562), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n563), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n564) );
  AND2X2 AND2X2_4914 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n561), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n565), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_stage1_2_) );
  AND2X2 AND2X2_4915 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_7_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n569) );
  AND2X2 AND2X2_4916 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n558), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n570), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n571) );
  AND2X2 AND2X2_4917 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n548), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n569), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n572) );
  AND2X2 AND2X2_4918 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n576), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n574), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n577) );
  AND2X2 AND2X2_4919 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n579), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n580), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_stage1_3_) );
  AND2X2 AND2X2_492 ( .A(AES_CORE_DATAPATH__abc_16259_n3274_1), .B(AES_CORE_DATAPATH__abc_16259_n3276), .Y(AES_CORE_DATAPATH__abc_16259_n3277) );
  AND2X2 AND2X2_4920 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n584), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n582), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_2_) );
  AND2X2 AND2X2_4921 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n313), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n258), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n586) );
  AND2X2 AND2X2_4922 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n297), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n317), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n587) );
  AND2X2 AND2X2_4923 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n590), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n589), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_7_) );
  AND2X2 AND2X2_4924 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n50), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n51_1) );
  AND2X2 AND2X2_4925 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n52), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n53_1) );
  AND2X2 AND2X2_4926 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n57), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n59), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n60) );
  AND2X2 AND2X2_4927 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n55), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n61), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n62) );
  AND2X2 AND2X2_4928 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n54_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n60), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n63) );
  AND2X2 AND2X2_4929 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n64), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf2), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n65) );
  AND2X2 AND2X2_493 ( .A(AES_CORE_DATAPATH__abc_16259_n2782_bF_buf3), .B(AES_CORE_DATAPATH_col_3__11_), .Y(AES_CORE_DATAPATH__abc_16259_n3278) );
  AND2X2 AND2X2_4930 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n54_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n67), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n68) );
  AND2X2 AND2X2_4931 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n55), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n69) );
  AND2X2 AND2X2_4932 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n70), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n71_1) );
  AND2X2 AND2X2_4933 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n73), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n72), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n74) );
  AND2X2 AND2X2_4934 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n75), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n66_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n76) );
  AND2X2 AND2X2_4935 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n78), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n80), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n81) );
  AND2X2 AND2X2_4936 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n70), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n83) );
  AND2X2 AND2X2_4937 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n73), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n56), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n84_1) );
  AND2X2 AND2X2_4938 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n85), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf7), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n86_1) );
  AND2X2 AND2X2_4939 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n87), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n82), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_5_) );
  AND2X2 AND2X2_494 ( .A(AES_CORE_DATAPATH__abc_16259_n2786_bF_buf3), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_75_), .Y(AES_CORE_DATAPATH__abc_16259_n3279) );
  AND2X2 AND2X2_4940 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n54_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n89) );
  AND2X2 AND2X2_4941 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n55), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n56), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n90) );
  AND2X2 AND2X2_4942 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n73), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n66_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n94_1) );
  AND2X2 AND2X2_4943 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n96), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n97_1) );
  AND2X2 AND2X2_4944 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n95), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n79), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n98) );
  AND2X2 AND2X2_4945 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n100), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n101_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n102) );
  AND2X2 AND2X2_4946 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n102), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n66_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n103) );
  AND2X2 AND2X2_4947 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n61), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n104_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n105) );
  AND2X2 AND2X2_4948 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n60), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n106) );
  AND2X2 AND2X2_4949 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n73), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n107), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n108) );
  AND2X2 AND2X2_495 ( .A(AES_CORE_DATAPATH__abc_16259_n2789_bF_buf3), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_43_), .Y(AES_CORE_DATAPATH__abc_16259_n3280) );
  AND2X2 AND2X2_4950 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n109), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n70), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n110) );
  AND2X2 AND2X2_4951 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n75), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n116) );
  AND2X2 AND2X2_4952 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n117), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n118), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n119) );
  AND2X2 AND2X2_4953 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n85), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n121_1) );
  AND2X2 AND2X2_4954 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n122), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n123), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n124) );
  AND2X2 AND2X2_4955 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n120), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n125), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n126_1) );
  AND2X2 AND2X2_4956 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n128), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n129), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n130) );
  AND2X2 AND2X2_4957 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n131), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n79), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n132) );
  AND2X2 AND2X2_4958 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n130), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n133) );
  AND2X2 AND2X2_4959 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n92), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n135), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n136) );
  AND2X2 AND2X2_496 ( .A(AES_CORE_DATAPATH__abc_16259_n3283), .B(AES_CORE_DATAPATH__abc_16259_n3277), .Y(AES_CORE_DATAPATH__abc_16259_n3284) );
  AND2X2 AND2X2_4960 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n107), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n66_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n138) );
  AND2X2 AND2X2_4961 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n50), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf4), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n139_1) );
  AND2X2 AND2X2_4962 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n142), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n143_1) );
  AND2X2 AND2X2_4963 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n102), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n52), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n144) );
  AND2X2 AND2X2_4964 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n142), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n147) );
  AND2X2 AND2X2_4965 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n102), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n67), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n148_1) );
  AND2X2 AND2X2_4966 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n150_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n130), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n151_1) );
  AND2X2 AND2X2_4967 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n149), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n131), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n152_1) );
  AND2X2 AND2X2_4968 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n154), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n146_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_3_) );
  AND2X2 AND2X2_4969 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n156) );
  AND2X2 AND2X2_497 ( .A(AES_CORE_DATAPATH__abc_16259_n2837_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__11_), .Y(AES_CORE_DATAPATH__abc_16259_n3286_1) );
  AND2X2 AND2X2_4970 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n157) );
  AND2X2 AND2X2_4971 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n159), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n160) );
  AND2X2 AND2X2_4972 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n161), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n162) );
  AND2X2 AND2X2_4973 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n164) );
  AND2X2 AND2X2_4974 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n165), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n164), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n167) );
  AND2X2 AND2X2_4975 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n168), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n166_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n169) );
  AND2X2 AND2X2_4976 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n169), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n163), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n170) );
  AND2X2 AND2X2_4977 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n170), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n158), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n171) );
  AND2X2 AND2X2_4978 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_1_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n173) );
  AND2X2 AND2X2_4979 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n161), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n176_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n177) );
  AND2X2 AND2X2_498 ( .A(AES_CORE_DATAPATH__abc_16259_n2887_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__11_), .Y(AES_CORE_DATAPATH__abc_16259_n3288_1) );
  AND2X2 AND2X2_4980 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n175), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n177), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n178) );
  AND2X2 AND2X2_4981 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n183), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n174), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n184) );
  AND2X2 AND2X2_4982 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n189_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n186), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n190_1) );
  AND2X2 AND2X2_4983 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n169), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n180), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n191) );
  AND2X2 AND2X2_4984 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n191), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n158), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n192) );
  AND2X2 AND2X2_4985 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n185), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n194), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n195) );
  AND2X2 AND2X2_4986 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n197), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n199), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n200) );
  AND2X2 AND2X2_4987 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n195), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n201), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n202) );
  AND2X2 AND2X2_4988 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n173), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n159), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n203) );
  AND2X2 AND2X2_4989 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n163), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n176_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n205) );
  AND2X2 AND2X2_499 ( .A(AES_CORE_DATAPATH__abc_16259_n2830_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__11_), .Y(AES_CORE_DATAPATH__abc_16259_n3289) );
  AND2X2 AND2X2_4990 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n169), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n162), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n207) );
  AND2X2 AND2X2_4991 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n214), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n208), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n215) );
  AND2X2 AND2X2_4992 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n211), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n216), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n217) );
  AND2X2 AND2X2_4993 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n219), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n221), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n222) );
  AND2X2 AND2X2_4994 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n217), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n222), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n223) );
  AND2X2 AND2X2_4995 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n202), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n223), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n224) );
  AND2X2 AND2X2_4996 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n190_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n193), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n225) );
  AND2X2 AND2X2_4997 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n184), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n172), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n226) );
  AND2X2 AND2X2_4998 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n230), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n229), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n231) );
  AND2X2 AND2X2_4999 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n233), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n234), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n235) );
  AND2X2 AND2X2_5 ( .A(_abc_15830_n13_1), .B(\addr[1] ), .Y(AES_CORE_DATAPATH_col_en_host_2_) );
  AND2X2 AND2X2_50 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n154), .B(AES_CORE_CONTROL_UNIT_state_7_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n155_1) );
  AND2X2 AND2X2_500 ( .A(AES_CORE_DATAPATH__abc_16259_n3291), .B(AES_CORE_DATAPATH__abc_16259_n3292), .Y(_auto_iopadmap_cc_313_execute_26949_11_) );
  AND2X2 AND2X2_5000 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n228), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n235), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n236) );
  AND2X2 AND2X2_5001 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n158), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n159), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n238) );
  AND2X2 AND2X2_5002 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n156), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n239) );
  AND2X2 AND2X2_5003 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n241), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n242), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n243) );
  AND2X2 AND2X2_5004 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n215), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n245) );
  AND2X2 AND2X2_5005 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n245), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n244), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n246) );
  AND2X2 AND2X2_5006 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n247), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n248), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n249) );
  AND2X2 AND2X2_5007 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n231), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n200), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n253) );
  AND2X2 AND2X2_5008 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n252), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n255), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n256) );
  AND2X2 AND2X2_5009 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n251), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n257), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n258) );
  AND2X2 AND2X2_501 ( .A(AES_CORE_DATAPATH__abc_16259_n2855_bF_buf3), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_11_), .Y(AES_CORE_DATAPATH__abc_16259_n3295) );
  AND2X2 AND2X2_5010 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n260), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n262), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n263) );
  AND2X2 AND2X2_5011 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n217), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n264), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n265) );
  AND2X2 AND2X2_5012 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n268), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n270), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n271) );
  AND2X2 AND2X2_5013 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n227), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n272), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n273) );
  AND2X2 AND2X2_5014 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n276), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n274), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n277) );
  AND2X2 AND2X2_5015 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n193), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n212), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n278) );
  AND2X2 AND2X2_5016 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n267), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n259), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n280) );
  AND2X2 AND2X2_5017 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n281) );
  AND2X2 AND2X2_5018 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n193), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n284) );
  AND2X2 AND2X2_5019 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n287), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n180), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n288) );
  AND2X2 AND2X2_502 ( .A(AES_CORE_DATAPATH__abc_16259_n2857_bF_buf3), .B(AES_CORE_DATAPATH_MIX_COL_col_1__3_), .Y(AES_CORE_DATAPATH__abc_16259_n3296) );
  AND2X2 AND2X2_5020 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n288), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n289), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n290) );
  AND2X2 AND2X2_5021 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n286), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n291), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n292) );
  AND2X2 AND2X2_5022 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n296), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n294), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n297) );
  AND2X2 AND2X2_5023 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n298), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n299), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n300) );
  AND2X2 AND2X2_5024 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n172), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n302) );
  AND2X2 AND2X2_5025 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n302), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n301), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n303) );
  AND2X2 AND2X2_5026 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n304), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n305), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n306) );
  AND2X2 AND2X2_5027 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n308), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n309), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n310) );
  AND2X2 AND2X2_5028 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n311), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n297), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n312) );
  AND2X2 AND2X2_5029 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n313), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n310), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n314) );
  AND2X2 AND2X2_503 ( .A(AES_CORE_DATAPATH__abc_16259_n3294_1), .B(AES_CORE_DATAPATH__abc_16259_n3298), .Y(AES_CORE_DATAPATH__abc_16259_n3299_1) );
  AND2X2 AND2X2_5030 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n315), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n258), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n316) );
  AND2X2 AND2X2_5031 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n318), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n317), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n319) );
  AND2X2 AND2X2_5032 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n227), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n232), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n321) );
  AND2X2 AND2X2_5033 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n217), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n201), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n323) );
  AND2X2 AND2X2_5034 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n325), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n326), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n327) );
  AND2X2 AND2X2_5035 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n172), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n329) );
  AND2X2 AND2X2_5036 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n329), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n244), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n330) );
  AND2X2 AND2X2_5037 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n331), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n332), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n333) );
  AND2X2 AND2X2_5038 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n334), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n336), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n337) );
  AND2X2 AND2X2_5039 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n313), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n338), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n339) );
  AND2X2 AND2X2_504 ( .A(_auto_iopadmap_cc_313_execute_26949_11_), .B(AES_CORE_DATAPATH__abc_16259_n3299_1), .Y(AES_CORE_DATAPATH__abc_16259_n3302) );
  AND2X2 AND2X2_5040 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n297), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n337), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n340) );
  AND2X2 AND2X2_5041 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n342), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n343), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n344) );
  AND2X2 AND2X2_5042 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n288), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n345), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n346) );
  AND2X2 AND2X2_5043 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n193), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n347) );
  AND2X2 AND2X2_5044 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n351), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n349), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n352) );
  AND2X2 AND2X2_5045 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n354), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n355), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n356) );
  AND2X2 AND2X2_5046 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n212), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n358) );
  AND2X2 AND2X2_5047 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n361), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n359), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n362) );
  AND2X2 AND2X2_5048 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n365), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n364), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n366) );
  AND2X2 AND2X2_5049 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n363), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n367), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n368) );
  AND2X2 AND2X2_505 ( .A(AES_CORE_DATAPATH_last_round_pp2_bF_buf2), .B(AES_CORE_DATAPATH_MIX_COL_col_1__3_), .Y(AES_CORE_DATAPATH__abc_16259_n3305) );
  AND2X2 AND2X2_5050 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n195), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n264), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n369) );
  AND2X2 AND2X2_5051 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n217), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n271), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n370) );
  AND2X2 AND2X2_5052 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n369), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n370), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n371) );
  AND2X2 AND2X2_5053 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n373), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n374), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n375) );
  AND2X2 AND2X2_5054 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n372), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n375), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n376) );
  AND2X2 AND2X2_5055 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n215), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n378) );
  AND2X2 AND2X2_5056 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n378), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n301), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n379) );
  AND2X2 AND2X2_5057 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n380), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n381), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n382) );
  AND2X2 AND2X2_5058 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n231), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n263), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n386) );
  AND2X2 AND2X2_5059 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n385), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n388), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n389) );
  AND2X2 AND2X2_506 ( .A(AES_CORE_DATAPATH__abc_16259_n2798_bF_buf3), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_11_), .Y(AES_CORE_DATAPATH__abc_16259_n3306) );
  AND2X2 AND2X2_5060 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n384), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n390), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n391) );
  AND2X2 AND2X2_5061 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n393), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n394), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n395) );
  AND2X2 AND2X2_5062 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n396), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n397), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n398) );
  AND2X2 AND2X2_5063 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n392), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n399), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_15_) );
  AND2X2 AND2X2_5064 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n395), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n398), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n403) );
  AND2X2 AND2X2_5065 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n368), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n391), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n404) );
  AND2X2 AND2X2_5066 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n402), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n406), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n407) );
  AND2X2 AND2X2_5067 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n410), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n408), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_10_) );
  AND2X2 AND2X2_5068 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n212), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n412) );
  AND2X2 AND2X2_5069 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n415), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n414), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n416) );
  AND2X2 AND2X2_507 ( .A(AES_CORE_DATAPATH__abc_16259_n3304), .B(AES_CORE_DATAPATH__abc_16259_n3308), .Y(AES_CORE_DATAPATH__abc_16259_n3309) );
  AND2X2 AND2X2_5070 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n419), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n418), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n420) );
  AND2X2 AND2X2_5071 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n417), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n421), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n422) );
  AND2X2 AND2X2_5072 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n395), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n422), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n423) );
  AND2X2 AND2X2_5073 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n424), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n425), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n426) );
  AND2X2 AND2X2_5074 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n368), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n426), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n427) );
  AND2X2 AND2X2_5075 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n429), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n430), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n431) );
  AND2X2 AND2X2_5076 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n434), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n435), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n436) );
  AND2X2 AND2X2_5077 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n433), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n437), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_12_) );
  AND2X2 AND2X2_5078 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n432), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n439), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_11_) );
  AND2X2 AND2X2_5079 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n441), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n442), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n443) );
  AND2X2 AND2X2_508 ( .A(AES_CORE_DATAPATH__abc_16259_n3309), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf8), .Y(AES_CORE_DATAPATH__abc_16259_n3310) );
  AND2X2 AND2X2_5080 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n445), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n444), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_3_) );
  AND2X2 AND2X2_5081 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n447), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n448), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n449) );
  AND2X2 AND2X2_5082 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_12_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_13_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n451) );
  AND2X2 AND2X2_5083 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n431), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n401), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n452) );
  AND2X2 AND2X2_5084 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n454), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n450), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_5_) );
  AND2X2 AND2X2_5085 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n457), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n456), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_6_) );
  AND2X2 AND2X2_5086 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n317), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n398), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n459) );
  AND2X2 AND2X2_5087 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n258), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n391), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n460) );
  AND2X2 AND2X2_5088 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n463), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n464), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_9_) );
  AND2X2 AND2X2_5089 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n467), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n466), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n468) );
  AND2X2 AND2X2_509 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf0), .B(AES_CORE_DATAPATH_col_3__11_), .Y(AES_CORE_DATAPATH__abc_16259_n3311) );
  AND2X2 AND2X2_5090 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n126_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n469), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n470) );
  AND2X2 AND2X2_5091 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n472), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n473) );
  AND2X2 AND2X2_5092 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n469), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n474) );
  AND2X2 AND2X2_5093 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n471), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n475), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n476) );
  AND2X2 AND2X2_5094 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n468), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n476), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n477) );
  AND2X2 AND2X2_5095 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n478) );
  AND2X2 AND2X2_5096 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n470), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n479), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n480) );
  AND2X2 AND2X2_5097 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n483), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n482), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n484) );
  AND2X2 AND2X2_5098 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n486), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n487) );
  AND2X2 AND2X2_5099 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n469), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n488) );
  AND2X2 AND2X2_51 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n90), .B(AES_CORE_CONTROL_UNIT__abc_15841_n98), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n156) );
  AND2X2 AND2X2_510 ( .A(AES_CORE_DATAPATH__abc_16259_n3314), .B(AES_CORE_DATAPATH__abc_16259_n3316), .Y(AES_CORE_DATAPATH__abc_16259_n3317_1) );
  AND2X2 AND2X2_5100 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n485), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n489), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n490) );
  AND2X2 AND2X2_5101 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n494), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n492), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n495) );
  AND2X2 AND2X2_5102 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n472), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n114), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n497) );
  AND2X2 AND2X2_5103 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n498), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n496), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n499) );
  AND2X2 AND2X2_5104 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n499), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n495), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n500) );
  AND2X2 AND2X2_5105 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n491), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n500), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n501) );
  AND2X2 AND2X2_5106 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n502), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n503), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n504) );
  AND2X2 AND2X2_5107 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n505), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n481), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n506) );
  AND2X2 AND2X2_5108 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n504), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n507), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n508) );
  AND2X2 AND2X2_5109 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n114), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n512) );
  AND2X2 AND2X2_511 ( .A(AES_CORE_DATAPATH__abc_16259_n2782_bF_buf2), .B(AES_CORE_DATAPATH_col_3__12_), .Y(AES_CORE_DATAPATH__abc_16259_n3318) );
  AND2X2 AND2X2_5110 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n513), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n511), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n514) );
  AND2X2 AND2X2_5111 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n515), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n510), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n516) );
  AND2X2 AND2X2_5112 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n514), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n475), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n517) );
  AND2X2 AND2X2_5113 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n519), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n520), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n521) );
  AND2X2 AND2X2_5114 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n522), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n523), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n524) );
  AND2X2 AND2X2_5115 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n521), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n525), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n526) );
  AND2X2 AND2X2_5116 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n468), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n524), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n527) );
  AND2X2 AND2X2_5117 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n528), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n518), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n529) );
  AND2X2 AND2X2_5118 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n521), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n510), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n530) );
  AND2X2 AND2X2_5119 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n530), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n479), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n531) );
  AND2X2 AND2X2_512 ( .A(AES_CORE_DATAPATH__abc_16259_n2786_bF_buf2), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_76_), .Y(AES_CORE_DATAPATH__abc_16259_n3319) );
  AND2X2 AND2X2_5120 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n532), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n478), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n533) );
  AND2X2 AND2X2_5121 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n534), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n490), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n535) );
  AND2X2 AND2X2_5122 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n536), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n537), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n538) );
  AND2X2 AND2X2_5123 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n538), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n491), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n539) );
  AND2X2 AND2X2_5124 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n543), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n544), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n545) );
  AND2X2 AND2X2_5125 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n541), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n546), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_stage1_1_) );
  AND2X2 AND2X2_5126 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n515), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n525), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n548) );
  AND2X2 AND2X2_5127 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n549) );
  AND2X2 AND2X2_5128 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n551), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n549), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n552) );
  AND2X2 AND2X2_5129 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n553), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n554), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n555) );
  AND2X2 AND2X2_513 ( .A(AES_CORE_DATAPATH__abc_16259_n2789_bF_buf2), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_44_), .Y(AES_CORE_DATAPATH__abc_16259_n3320) );
  AND2X2 AND2X2_5130 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n557), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n559), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n560) );
  AND2X2 AND2X2_5131 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n562), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n563), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n564) );
  AND2X2 AND2X2_5132 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n561), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n565), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_stage1_2_) );
  AND2X2 AND2X2_5133 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_7_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n569) );
  AND2X2 AND2X2_5134 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n558), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n570), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n571) );
  AND2X2 AND2X2_5135 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n548), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n569), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n572) );
  AND2X2 AND2X2_5136 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n576), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n574), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n577) );
  AND2X2 AND2X2_5137 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n579), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n580), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_stage1_3_) );
  AND2X2 AND2X2_5138 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n584), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n582), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_2_) );
  AND2X2 AND2X2_5139 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n313), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n258), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n586) );
  AND2X2 AND2X2_514 ( .A(AES_CORE_DATAPATH__abc_16259_n3323_1), .B(AES_CORE_DATAPATH__abc_16259_n3317_1), .Y(AES_CORE_DATAPATH__abc_16259_n3324) );
  AND2X2 AND2X2_5140 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n297), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n317), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n587) );
  AND2X2 AND2X2_5141 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n590), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n589), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_7_) );
  AND2X2 AND2X2_5142 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n50), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n51_1) );
  AND2X2 AND2X2_5143 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n52), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n53_1) );
  AND2X2 AND2X2_5144 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n57), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n59), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n60) );
  AND2X2 AND2X2_5145 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n55), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n61), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n62) );
  AND2X2 AND2X2_5146 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n54_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n60), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n63) );
  AND2X2 AND2X2_5147 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n64), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf2), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n65) );
  AND2X2 AND2X2_5148 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n54_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n67), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n68) );
  AND2X2 AND2X2_5149 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n55), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n69) );
  AND2X2 AND2X2_515 ( .A(AES_CORE_DATAPATH__abc_16259_n2837_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__12_), .Y(AES_CORE_DATAPATH__abc_16259_n3326_1) );
  AND2X2 AND2X2_5150 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n70), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n71_1) );
  AND2X2 AND2X2_5151 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n73), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n72), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n74) );
  AND2X2 AND2X2_5152 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n75), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n66_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n76) );
  AND2X2 AND2X2_5153 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n78), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n80), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n81) );
  AND2X2 AND2X2_5154 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n70), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n83) );
  AND2X2 AND2X2_5155 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n73), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n56), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n84_1) );
  AND2X2 AND2X2_5156 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n85), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf7), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n86_1) );
  AND2X2 AND2X2_5157 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n87), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n82), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_5_) );
  AND2X2 AND2X2_5158 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n54_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n89) );
  AND2X2 AND2X2_5159 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n55), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n56), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n90) );
  AND2X2 AND2X2_516 ( .A(AES_CORE_DATAPATH__abc_16259_n2887_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__12_), .Y(AES_CORE_DATAPATH__abc_16259_n3328_1) );
  AND2X2 AND2X2_5160 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n73), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n66_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n94_1) );
  AND2X2 AND2X2_5161 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n96), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n97_1) );
  AND2X2 AND2X2_5162 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n95), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n79), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n98) );
  AND2X2 AND2X2_5163 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n100), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n101_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n102) );
  AND2X2 AND2X2_5164 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n102), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n66_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n103) );
  AND2X2 AND2X2_5165 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n61), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n104_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n105) );
  AND2X2 AND2X2_5166 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n60), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n106) );
  AND2X2 AND2X2_5167 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n73), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n107), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n108) );
  AND2X2 AND2X2_5168 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n109), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n70), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n110) );
  AND2X2 AND2X2_5169 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n75), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n116) );
  AND2X2 AND2X2_517 ( .A(AES_CORE_DATAPATH__abc_16259_n2830_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__12_), .Y(AES_CORE_DATAPATH__abc_16259_n3329) );
  AND2X2 AND2X2_5170 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n117), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n118), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n119) );
  AND2X2 AND2X2_5171 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n85), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n121_1) );
  AND2X2 AND2X2_5172 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n122), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n123), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n124) );
  AND2X2 AND2X2_5173 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n120), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n125), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n126_1) );
  AND2X2 AND2X2_5174 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n128), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n129), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n130) );
  AND2X2 AND2X2_5175 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n131), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n79), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n132) );
  AND2X2 AND2X2_5176 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n130), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n133) );
  AND2X2 AND2X2_5177 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n92), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n135), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n136) );
  AND2X2 AND2X2_5178 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n107), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n66_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n138) );
  AND2X2 AND2X2_5179 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n50), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf4), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n139_1) );
  AND2X2 AND2X2_518 ( .A(AES_CORE_DATAPATH__abc_16259_n3331), .B(AES_CORE_DATAPATH__abc_16259_n3332_1), .Y(_auto_iopadmap_cc_313_execute_26949_12_) );
  AND2X2 AND2X2_5180 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n142), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n143_1) );
  AND2X2 AND2X2_5181 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n102), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n52), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n144) );
  AND2X2 AND2X2_5182 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n142), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n147) );
  AND2X2 AND2X2_5183 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n102), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n67), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n148_1) );
  AND2X2 AND2X2_5184 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n150_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n130), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n151_1) );
  AND2X2 AND2X2_5185 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n149), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n131), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n152_1) );
  AND2X2 AND2X2_5186 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n154), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n146_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_3_) );
  AND2X2 AND2X2_5187 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n156) );
  AND2X2 AND2X2_5188 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n157) );
  AND2X2 AND2X2_5189 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n159), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n160) );
  AND2X2 AND2X2_519 ( .A(AES_CORE_DATAPATH__abc_16259_n2855_bF_buf2), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_12_), .Y(AES_CORE_DATAPATH__abc_16259_n3335) );
  AND2X2 AND2X2_5190 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n161), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n162) );
  AND2X2 AND2X2_5191 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n164) );
  AND2X2 AND2X2_5192 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n165), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n164), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n167) );
  AND2X2 AND2X2_5193 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n168), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n166_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n169) );
  AND2X2 AND2X2_5194 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n169), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n163), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n170) );
  AND2X2 AND2X2_5195 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n170), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n158), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n171) );
  AND2X2 AND2X2_5196 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_1_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n173) );
  AND2X2 AND2X2_5197 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n161), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n176_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n177) );
  AND2X2 AND2X2_5198 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n175), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n177), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n178) );
  AND2X2 AND2X2_5199 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n183), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n174), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n184) );
  AND2X2 AND2X2_52 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf11), .B(AES_CORE_CONTROL_UNIT_state_6_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n158) );
  AND2X2 AND2X2_520 ( .A(AES_CORE_DATAPATH__abc_16259_n2857_bF_buf2), .B(AES_CORE_DATAPATH_MIX_COL_col_1__4_), .Y(AES_CORE_DATAPATH__abc_16259_n3336) );
  AND2X2 AND2X2_5200 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n189_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n186), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n190_1) );
  AND2X2 AND2X2_5201 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n169), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n180), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n191) );
  AND2X2 AND2X2_5202 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n191), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n158), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n192) );
  AND2X2 AND2X2_5203 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n185), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n194), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n195) );
  AND2X2 AND2X2_5204 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n197), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n199), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n200) );
  AND2X2 AND2X2_5205 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n195), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n201), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n202) );
  AND2X2 AND2X2_5206 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n173), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n159), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n203) );
  AND2X2 AND2X2_5207 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n163), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n176_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n205) );
  AND2X2 AND2X2_5208 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n169), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n162), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n207) );
  AND2X2 AND2X2_5209 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n214), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n208), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n215) );
  AND2X2 AND2X2_521 ( .A(AES_CORE_DATAPATH__abc_16259_n3334), .B(AES_CORE_DATAPATH__abc_16259_n3338), .Y(AES_CORE_DATAPATH__abc_16259_n3339) );
  AND2X2 AND2X2_5210 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n211), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n216), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n217) );
  AND2X2 AND2X2_5211 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n219), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n221), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n222) );
  AND2X2 AND2X2_5212 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n217), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n222), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n223) );
  AND2X2 AND2X2_5213 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n202), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n223), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n224) );
  AND2X2 AND2X2_5214 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n190_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n193), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n225) );
  AND2X2 AND2X2_5215 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n184), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n172), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n226) );
  AND2X2 AND2X2_5216 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n230), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n229), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n231) );
  AND2X2 AND2X2_5217 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n233), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n234), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n235) );
  AND2X2 AND2X2_5218 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n228), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n235), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n236) );
  AND2X2 AND2X2_5219 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n158), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n159), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n238) );
  AND2X2 AND2X2_522 ( .A(_auto_iopadmap_cc_313_execute_26949_12_), .B(AES_CORE_DATAPATH__abc_16259_n3339), .Y(AES_CORE_DATAPATH__abc_16259_n3342) );
  AND2X2 AND2X2_5220 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n156), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n239) );
  AND2X2 AND2X2_5221 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n241), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n242), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n243) );
  AND2X2 AND2X2_5222 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n215), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n245) );
  AND2X2 AND2X2_5223 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n245), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n244), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n246) );
  AND2X2 AND2X2_5224 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n247), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n248), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n249) );
  AND2X2 AND2X2_5225 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n231), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n200), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n253) );
  AND2X2 AND2X2_5226 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n252), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n255), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n256) );
  AND2X2 AND2X2_5227 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n251), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n257), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n258) );
  AND2X2 AND2X2_5228 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n260), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n262), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n263) );
  AND2X2 AND2X2_5229 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n217), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n264), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n265) );
  AND2X2 AND2X2_523 ( .A(AES_CORE_DATAPATH_last_round_pp2_bF_buf1), .B(AES_CORE_DATAPATH_MIX_COL_col_1__4_), .Y(AES_CORE_DATAPATH__abc_16259_n3345) );
  AND2X2 AND2X2_5230 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n268), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n270), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n271) );
  AND2X2 AND2X2_5231 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n227), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n272), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n273) );
  AND2X2 AND2X2_5232 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n276), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n274), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n277) );
  AND2X2 AND2X2_5233 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n193), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n212), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n278) );
  AND2X2 AND2X2_5234 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n267), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n259), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n280) );
  AND2X2 AND2X2_5235 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n281) );
  AND2X2 AND2X2_5236 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n193), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n284) );
  AND2X2 AND2X2_5237 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n287), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n180), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n288) );
  AND2X2 AND2X2_5238 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n288), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n289), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n290) );
  AND2X2 AND2X2_5239 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n286), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n291), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n292) );
  AND2X2 AND2X2_524 ( .A(AES_CORE_DATAPATH__abc_16259_n2798_bF_buf2), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_12_), .Y(AES_CORE_DATAPATH__abc_16259_n3346_1) );
  AND2X2 AND2X2_5240 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n296), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n294), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n297) );
  AND2X2 AND2X2_5241 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n298), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n299), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n300) );
  AND2X2 AND2X2_5242 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n172), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n302) );
  AND2X2 AND2X2_5243 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n302), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n301), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n303) );
  AND2X2 AND2X2_5244 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n304), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n305), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n306) );
  AND2X2 AND2X2_5245 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n308), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n309), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n310) );
  AND2X2 AND2X2_5246 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n311), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n297), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n312) );
  AND2X2 AND2X2_5247 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n313), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n310), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n314) );
  AND2X2 AND2X2_5248 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n315), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n258), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n316) );
  AND2X2 AND2X2_5249 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n318), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n317), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n319) );
  AND2X2 AND2X2_525 ( .A(AES_CORE_DATAPATH__abc_16259_n3344_1), .B(AES_CORE_DATAPATH__abc_16259_n3348), .Y(AES_CORE_DATAPATH__abc_16259_n3349) );
  AND2X2 AND2X2_5250 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n227), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n232), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n321) );
  AND2X2 AND2X2_5251 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n217), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n201), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n323) );
  AND2X2 AND2X2_5252 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n325), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n326), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n327) );
  AND2X2 AND2X2_5253 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n172), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n329) );
  AND2X2 AND2X2_5254 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n329), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n244), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n330) );
  AND2X2 AND2X2_5255 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n331), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n332), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n333) );
  AND2X2 AND2X2_5256 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n334), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n336), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n337) );
  AND2X2 AND2X2_5257 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n313), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n338), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n339) );
  AND2X2 AND2X2_5258 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n297), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n337), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n340) );
  AND2X2 AND2X2_5259 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n342), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n343), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n344) );
  AND2X2 AND2X2_526 ( .A(AES_CORE_DATAPATH__abc_16259_n3349), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n3350) );
  AND2X2 AND2X2_5260 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n288), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n345), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n346) );
  AND2X2 AND2X2_5261 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n193), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n347) );
  AND2X2 AND2X2_5262 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n351), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n349), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n352) );
  AND2X2 AND2X2_5263 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n354), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n355), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n356) );
  AND2X2 AND2X2_5264 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n212), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n358) );
  AND2X2 AND2X2_5265 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n361), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n359), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n362) );
  AND2X2 AND2X2_5266 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n365), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n364), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n366) );
  AND2X2 AND2X2_5267 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n363), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n367), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n368) );
  AND2X2 AND2X2_5268 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n195), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n264), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n369) );
  AND2X2 AND2X2_5269 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n217), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n271), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n370) );
  AND2X2 AND2X2_527 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf12), .B(AES_CORE_DATAPATH_col_3__12_), .Y(AES_CORE_DATAPATH__abc_16259_n3351_1) );
  AND2X2 AND2X2_5270 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n369), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n370), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n371) );
  AND2X2 AND2X2_5271 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n373), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n374), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n375) );
  AND2X2 AND2X2_5272 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n372), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n375), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n376) );
  AND2X2 AND2X2_5273 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n215), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n378) );
  AND2X2 AND2X2_5274 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n378), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n301), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n379) );
  AND2X2 AND2X2_5275 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n380), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n381), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n382) );
  AND2X2 AND2X2_5276 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n231), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n263), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n386) );
  AND2X2 AND2X2_5277 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n385), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n388), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n389) );
  AND2X2 AND2X2_5278 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n384), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n390), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n391) );
  AND2X2 AND2X2_5279 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n393), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n394), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n395) );
  AND2X2 AND2X2_528 ( .A(AES_CORE_DATAPATH__abc_16259_n3354), .B(AES_CORE_DATAPATH__abc_16259_n3356), .Y(AES_CORE_DATAPATH__abc_16259_n3357_1) );
  AND2X2 AND2X2_5280 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n396), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n397), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n398) );
  AND2X2 AND2X2_5281 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n392), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n399), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_23_) );
  AND2X2 AND2X2_5282 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n395), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n398), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n403) );
  AND2X2 AND2X2_5283 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n368), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n391), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n404) );
  AND2X2 AND2X2_5284 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n402), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n406), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n407) );
  AND2X2 AND2X2_5285 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n410), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n408), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_18_) );
  AND2X2 AND2X2_5286 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n212), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n412) );
  AND2X2 AND2X2_5287 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n415), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n414), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n416) );
  AND2X2 AND2X2_5288 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n419), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n418), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n420) );
  AND2X2 AND2X2_5289 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n417), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n421), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n422) );
  AND2X2 AND2X2_529 ( .A(AES_CORE_DATAPATH__abc_16259_n2782_bF_buf1), .B(AES_CORE_DATAPATH_col_3__13_), .Y(AES_CORE_DATAPATH__abc_16259_n3358) );
  AND2X2 AND2X2_5290 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n395), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n422), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n423) );
  AND2X2 AND2X2_5291 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n424), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n425), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n426) );
  AND2X2 AND2X2_5292 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n368), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n426), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n427) );
  AND2X2 AND2X2_5293 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n429), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n430), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n431) );
  AND2X2 AND2X2_5294 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n434), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n435), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n436) );
  AND2X2 AND2X2_5295 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n433), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n437), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_20_) );
  AND2X2 AND2X2_5296 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n432), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n439), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_19_) );
  AND2X2 AND2X2_5297 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n441), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n442), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n443) );
  AND2X2 AND2X2_5298 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n445), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n444), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_3_) );
  AND2X2 AND2X2_5299 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n447), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n448), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n449) );
  AND2X2 AND2X2_53 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n106_1), .B(AES_CORE_CONTROL_UNIT_state_1_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n159) );
  AND2X2 AND2X2_530 ( .A(AES_CORE_DATAPATH__abc_16259_n2786_bF_buf1), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_77_), .Y(AES_CORE_DATAPATH__abc_16259_n3359_1) );
  AND2X2 AND2X2_5300 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_20_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_21_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n451) );
  AND2X2 AND2X2_5301 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n431), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n401), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n452) );
  AND2X2 AND2X2_5302 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n454), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n450), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_5_) );
  AND2X2 AND2X2_5303 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n457), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n456), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_6_) );
  AND2X2 AND2X2_5304 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n317), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n398), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n459) );
  AND2X2 AND2X2_5305 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n258), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n391), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n460) );
  AND2X2 AND2X2_5306 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n463), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n464), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_17_) );
  AND2X2 AND2X2_5307 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n467), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n466), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n468) );
  AND2X2 AND2X2_5308 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n126_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n469), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n470) );
  AND2X2 AND2X2_5309 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n472), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n473) );
  AND2X2 AND2X2_531 ( .A(AES_CORE_DATAPATH__abc_16259_n2789_bF_buf1), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_45_), .Y(AES_CORE_DATAPATH__abc_16259_n3360) );
  AND2X2 AND2X2_5310 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n469), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n474) );
  AND2X2 AND2X2_5311 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n471), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n475), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n476) );
  AND2X2 AND2X2_5312 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n468), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n476), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n477) );
  AND2X2 AND2X2_5313 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n478) );
  AND2X2 AND2X2_5314 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n470), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n479), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n480) );
  AND2X2 AND2X2_5315 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n483), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n482), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n484) );
  AND2X2 AND2X2_5316 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n486), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n487) );
  AND2X2 AND2X2_5317 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n469), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n488) );
  AND2X2 AND2X2_5318 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n485), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n489), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n490) );
  AND2X2 AND2X2_5319 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n494), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n492), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n495) );
  AND2X2 AND2X2_532 ( .A(AES_CORE_DATAPATH__abc_16259_n3363), .B(AES_CORE_DATAPATH__abc_16259_n3357_1), .Y(AES_CORE_DATAPATH__abc_16259_n3364) );
  AND2X2 AND2X2_5320 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n472), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n114), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n497) );
  AND2X2 AND2X2_5321 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n498), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n496), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n499) );
  AND2X2 AND2X2_5322 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n499), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n495), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n500) );
  AND2X2 AND2X2_5323 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n491), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n500), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n501) );
  AND2X2 AND2X2_5324 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n502), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n503), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n504) );
  AND2X2 AND2X2_5325 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n505), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n481), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n506) );
  AND2X2 AND2X2_5326 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n504), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n507), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n508) );
  AND2X2 AND2X2_5327 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n114), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n512) );
  AND2X2 AND2X2_5328 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n513), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n511), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n514) );
  AND2X2 AND2X2_5329 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n515), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n510), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n516) );
  AND2X2 AND2X2_533 ( .A(AES_CORE_DATAPATH__abc_16259_n2837_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__13_), .Y(AES_CORE_DATAPATH__abc_16259_n3366) );
  AND2X2 AND2X2_5330 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n514), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n475), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n517) );
  AND2X2 AND2X2_5331 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n519), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n520), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n521) );
  AND2X2 AND2X2_5332 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n522), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n523), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n524) );
  AND2X2 AND2X2_5333 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n521), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n525), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n526) );
  AND2X2 AND2X2_5334 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n468), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n524), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n527) );
  AND2X2 AND2X2_5335 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n528), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n518), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n529) );
  AND2X2 AND2X2_5336 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n521), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n510), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n530) );
  AND2X2 AND2X2_5337 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n530), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n479), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n531) );
  AND2X2 AND2X2_5338 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n532), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n478), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n533) );
  AND2X2 AND2X2_5339 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n534), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n490), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n535) );
  AND2X2 AND2X2_534 ( .A(AES_CORE_DATAPATH__abc_16259_n2887_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__13_), .Y(AES_CORE_DATAPATH__abc_16259_n3368) );
  AND2X2 AND2X2_5340 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n536), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n537), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n538) );
  AND2X2 AND2X2_5341 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n538), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n491), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n539) );
  AND2X2 AND2X2_5342 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n543), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n544), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n545) );
  AND2X2 AND2X2_5343 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n541), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n546), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_stage1_1_) );
  AND2X2 AND2X2_5344 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n515), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n525), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n548) );
  AND2X2 AND2X2_5345 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n549) );
  AND2X2 AND2X2_5346 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n551), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n549), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n552) );
  AND2X2 AND2X2_5347 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n553), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n554), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n555) );
  AND2X2 AND2X2_5348 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n557), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n559), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n560) );
  AND2X2 AND2X2_5349 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n562), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n563), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n564) );
  AND2X2 AND2X2_535 ( .A(AES_CORE_DATAPATH__abc_16259_n2830_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__13_), .Y(AES_CORE_DATAPATH__abc_16259_n3369) );
  AND2X2 AND2X2_5350 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n561), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n565), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_stage1_2_) );
  AND2X2 AND2X2_5351 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_7_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n569) );
  AND2X2 AND2X2_5352 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n558), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n570), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n571) );
  AND2X2 AND2X2_5353 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n548), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n569), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n572) );
  AND2X2 AND2X2_5354 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n576), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n574), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n577) );
  AND2X2 AND2X2_5355 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n579), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n580), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_stage1_3_) );
  AND2X2 AND2X2_5356 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n584), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n582), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_2_) );
  AND2X2 AND2X2_5357 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n313), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n258), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n586) );
  AND2X2 AND2X2_5358 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n297), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n317), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n587) );
  AND2X2 AND2X2_5359 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n590), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n589), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_7_) );
  AND2X2 AND2X2_536 ( .A(AES_CORE_DATAPATH__abc_16259_n3371), .B(AES_CORE_DATAPATH__abc_16259_n3372), .Y(_auto_iopadmap_cc_313_execute_26949_13_) );
  AND2X2 AND2X2_5360 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n50), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n51_1) );
  AND2X2 AND2X2_5361 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n52), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n53_1) );
  AND2X2 AND2X2_5362 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n57), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n59), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n60) );
  AND2X2 AND2X2_5363 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n55), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n61), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n62) );
  AND2X2 AND2X2_5364 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n54_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n60), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n63) );
  AND2X2 AND2X2_5365 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n64), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf2), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n65) );
  AND2X2 AND2X2_5366 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n54_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n67), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n68) );
  AND2X2 AND2X2_5367 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n55), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n69) );
  AND2X2 AND2X2_5368 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n70), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n71_1) );
  AND2X2 AND2X2_5369 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n73), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n72), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n74) );
  AND2X2 AND2X2_537 ( .A(AES_CORE_DATAPATH__abc_16259_n2855_bF_buf1), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_13_), .Y(AES_CORE_DATAPATH__abc_16259_n3375_1) );
  AND2X2 AND2X2_5370 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n75), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n66_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n76) );
  AND2X2 AND2X2_5371 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n78), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n80), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n81) );
  AND2X2 AND2X2_5372 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n70), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n83) );
  AND2X2 AND2X2_5373 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n73), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n56), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n84_1) );
  AND2X2 AND2X2_5374 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n85), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf7), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n86_1) );
  AND2X2 AND2X2_5375 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n87), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n82), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_5_) );
  AND2X2 AND2X2_5376 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n54_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n89) );
  AND2X2 AND2X2_5377 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n55), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n56), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n90) );
  AND2X2 AND2X2_5378 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n73), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n66_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n94_1) );
  AND2X2 AND2X2_5379 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n96), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n97_1) );
  AND2X2 AND2X2_538 ( .A(AES_CORE_DATAPATH__abc_16259_n2857_bF_buf1), .B(AES_CORE_DATAPATH_MIX_COL_col_1__5_), .Y(AES_CORE_DATAPATH__abc_16259_n3376) );
  AND2X2 AND2X2_5380 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n95), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n79), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n98) );
  AND2X2 AND2X2_5381 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n100), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n101_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n102) );
  AND2X2 AND2X2_5382 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n102), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n66_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n103) );
  AND2X2 AND2X2_5383 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n61), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n104_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n105) );
  AND2X2 AND2X2_5384 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n60), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n106) );
  AND2X2 AND2X2_5385 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n73), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n107), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n108) );
  AND2X2 AND2X2_5386 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n109), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n70), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n110) );
  AND2X2 AND2X2_5387 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n75), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n116) );
  AND2X2 AND2X2_5388 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n117), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n118), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n119) );
  AND2X2 AND2X2_5389 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n85), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n121_1) );
  AND2X2 AND2X2_539 ( .A(AES_CORE_DATAPATH__abc_16259_n3374), .B(AES_CORE_DATAPATH__abc_16259_n3378), .Y(AES_CORE_DATAPATH__abc_16259_n3379) );
  AND2X2 AND2X2_5390 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n122), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n123), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n124) );
  AND2X2 AND2X2_5391 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n120), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n125), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n126_1) );
  AND2X2 AND2X2_5392 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n128), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n129), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n130) );
  AND2X2 AND2X2_5393 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n131), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n79), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n132) );
  AND2X2 AND2X2_5394 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n130), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n133) );
  AND2X2 AND2X2_5395 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n92), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n135), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n136) );
  AND2X2 AND2X2_5396 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n107), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n66_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n138) );
  AND2X2 AND2X2_5397 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n50), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf4), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n139_1) );
  AND2X2 AND2X2_5398 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n142), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n143_1) );
  AND2X2 AND2X2_5399 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n102), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n52), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n144) );
  AND2X2 AND2X2_54 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n160), .B(AES_CORE_CONTROL_UNIT__abc_15841_n84_1), .Y(AES_CORE_CONTROL_UNIT__abc_10818_n122) );
  AND2X2 AND2X2_540 ( .A(_auto_iopadmap_cc_313_execute_26949_13_), .B(AES_CORE_DATAPATH__abc_16259_n3379), .Y(AES_CORE_DATAPATH__abc_16259_n3382) );
  AND2X2 AND2X2_5400 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n142), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n147) );
  AND2X2 AND2X2_5401 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n102), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n67), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n148_1) );
  AND2X2 AND2X2_5402 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n150_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n130), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n151_1) );
  AND2X2 AND2X2_5403 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n149), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n131), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n152_1) );
  AND2X2 AND2X2_5404 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n154), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n146_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_3_) );
  AND2X2 AND2X2_5405 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n156) );
  AND2X2 AND2X2_5406 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n157) );
  AND2X2 AND2X2_5407 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n159), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n160) );
  AND2X2 AND2X2_5408 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n161), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n162) );
  AND2X2 AND2X2_5409 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n164) );
  AND2X2 AND2X2_541 ( .A(AES_CORE_DATAPATH_last_round_pp2_bF_buf0), .B(AES_CORE_DATAPATH_MIX_COL_col_1__5_), .Y(AES_CORE_DATAPATH__abc_16259_n3385) );
  AND2X2 AND2X2_5410 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n165), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n164), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n167) );
  AND2X2 AND2X2_5411 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n168), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n166_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n169) );
  AND2X2 AND2X2_5412 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n169), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n163), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n170) );
  AND2X2 AND2X2_5413 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n170), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n158), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n171) );
  AND2X2 AND2X2_5414 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_1_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n173) );
  AND2X2 AND2X2_5415 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n161), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n176_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n177) );
  AND2X2 AND2X2_5416 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n175), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n177), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n178) );
  AND2X2 AND2X2_5417 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n183), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n174), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n184) );
  AND2X2 AND2X2_5418 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n189_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n186), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n190_1) );
  AND2X2 AND2X2_5419 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n169), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n180), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n191) );
  AND2X2 AND2X2_542 ( .A(AES_CORE_DATAPATH__abc_16259_n2798_bF_buf1), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_13_), .Y(AES_CORE_DATAPATH__abc_16259_n3386_1) );
  AND2X2 AND2X2_5420 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n191), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n158), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n192) );
  AND2X2 AND2X2_5421 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n185), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n194), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n195) );
  AND2X2 AND2X2_5422 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n197), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n199), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n200) );
  AND2X2 AND2X2_5423 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n195), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n201), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n202) );
  AND2X2 AND2X2_5424 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n173), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n159), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n203) );
  AND2X2 AND2X2_5425 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n163), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n176_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n205) );
  AND2X2 AND2X2_5426 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n169), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n162), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n207) );
  AND2X2 AND2X2_5427 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n214), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n208), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n215) );
  AND2X2 AND2X2_5428 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n211), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n216), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n217) );
  AND2X2 AND2X2_5429 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n219), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n221), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n222) );
  AND2X2 AND2X2_543 ( .A(AES_CORE_DATAPATH__abc_16259_n3384_1), .B(AES_CORE_DATAPATH__abc_16259_n3388_1), .Y(AES_CORE_DATAPATH__abc_16259_n3389) );
  AND2X2 AND2X2_5430 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n217), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n222), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n223) );
  AND2X2 AND2X2_5431 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n202), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n223), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n224) );
  AND2X2 AND2X2_5432 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n190_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n193), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n225) );
  AND2X2 AND2X2_5433 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n184), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n172), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n226) );
  AND2X2 AND2X2_5434 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n230), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n229), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n231) );
  AND2X2 AND2X2_5435 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n233), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n234), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n235) );
  AND2X2 AND2X2_5436 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n228), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n235), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n236) );
  AND2X2 AND2X2_5437 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n158), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n159), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n238) );
  AND2X2 AND2X2_5438 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n156), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n239) );
  AND2X2 AND2X2_5439 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n241), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n242), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n243) );
  AND2X2 AND2X2_544 ( .A(AES_CORE_DATAPATH__abc_16259_n3389), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n3390_1) );
  AND2X2 AND2X2_5440 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n215), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n245) );
  AND2X2 AND2X2_5441 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n245), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n244), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n246) );
  AND2X2 AND2X2_5442 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n247), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n248), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n249) );
  AND2X2 AND2X2_5443 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n231), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n200), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n253) );
  AND2X2 AND2X2_5444 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n252), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n255), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n256) );
  AND2X2 AND2X2_5445 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n251), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n257), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n258) );
  AND2X2 AND2X2_5446 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n260), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n262), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n263) );
  AND2X2 AND2X2_5447 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n217), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n264), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n265) );
  AND2X2 AND2X2_5448 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n268), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n270), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n271) );
  AND2X2 AND2X2_5449 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n227), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n272), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n273) );
  AND2X2 AND2X2_545 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf11), .B(AES_CORE_DATAPATH_col_3__13_), .Y(AES_CORE_DATAPATH__abc_16259_n3391) );
  AND2X2 AND2X2_5450 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n276), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n274), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n277) );
  AND2X2 AND2X2_5451 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n193), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n212), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n278) );
  AND2X2 AND2X2_5452 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n267), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n259), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n280) );
  AND2X2 AND2X2_5453 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n281) );
  AND2X2 AND2X2_5454 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n193), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n284) );
  AND2X2 AND2X2_5455 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n287), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n180), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n288) );
  AND2X2 AND2X2_5456 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n288), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n289), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n290) );
  AND2X2 AND2X2_5457 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n286), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n291), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n292) );
  AND2X2 AND2X2_5458 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n296), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n294), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n297) );
  AND2X2 AND2X2_5459 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n298), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n299), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n300) );
  AND2X2 AND2X2_546 ( .A(AES_CORE_DATAPATH__abc_16259_n3394), .B(AES_CORE_DATAPATH__abc_16259_n3396), .Y(AES_CORE_DATAPATH__abc_16259_n3397) );
  AND2X2 AND2X2_5460 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n172), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n302) );
  AND2X2 AND2X2_5461 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n302), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n301), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n303) );
  AND2X2 AND2X2_5462 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n304), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n305), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n306) );
  AND2X2 AND2X2_5463 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n308), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n309), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n310) );
  AND2X2 AND2X2_5464 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n311), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n297), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n312) );
  AND2X2 AND2X2_5465 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n313), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n310), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n314) );
  AND2X2 AND2X2_5466 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n315), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n258), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n316) );
  AND2X2 AND2X2_5467 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n318), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n317), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n319) );
  AND2X2 AND2X2_5468 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n227), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n232), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n321) );
  AND2X2 AND2X2_5469 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n217), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n201), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n323) );
  AND2X2 AND2X2_547 ( .A(AES_CORE_DATAPATH__abc_16259_n2782_bF_buf0), .B(AES_CORE_DATAPATH_col_3__14_), .Y(AES_CORE_DATAPATH__abc_16259_n3398) );
  AND2X2 AND2X2_5470 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n325), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n326), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n327) );
  AND2X2 AND2X2_5471 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n172), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n329) );
  AND2X2 AND2X2_5472 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n329), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n244), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n330) );
  AND2X2 AND2X2_5473 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n331), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n332), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n333) );
  AND2X2 AND2X2_5474 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n334), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n336), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n337) );
  AND2X2 AND2X2_5475 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n313), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n338), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n339) );
  AND2X2 AND2X2_5476 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n297), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n337), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n340) );
  AND2X2 AND2X2_5477 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n342), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n343), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n344) );
  AND2X2 AND2X2_5478 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n288), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n345), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n346) );
  AND2X2 AND2X2_5479 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n193), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n347) );
  AND2X2 AND2X2_548 ( .A(AES_CORE_DATAPATH__abc_16259_n2786_bF_buf0), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_78_), .Y(AES_CORE_DATAPATH__abc_16259_n3399) );
  AND2X2 AND2X2_5480 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n351), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n349), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n352) );
  AND2X2 AND2X2_5481 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n354), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n355), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n356) );
  AND2X2 AND2X2_5482 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n212), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n358) );
  AND2X2 AND2X2_5483 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n361), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n359), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n362) );
  AND2X2 AND2X2_5484 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n365), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n364), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n366) );
  AND2X2 AND2X2_5485 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n363), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n367), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n368) );
  AND2X2 AND2X2_5486 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n195), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n264), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n369) );
  AND2X2 AND2X2_5487 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n217), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n271), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n370) );
  AND2X2 AND2X2_5488 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n369), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n370), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n371) );
  AND2X2 AND2X2_5489 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n373), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n374), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n375) );
  AND2X2 AND2X2_549 ( .A(AES_CORE_DATAPATH__abc_16259_n2789_bF_buf0), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_46_), .Y(AES_CORE_DATAPATH__abc_16259_n3400) );
  AND2X2 AND2X2_5490 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n372), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n375), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n376) );
  AND2X2 AND2X2_5491 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n215), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n378) );
  AND2X2 AND2X2_5492 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n378), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n301), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n379) );
  AND2X2 AND2X2_5493 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n380), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n381), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n382) );
  AND2X2 AND2X2_5494 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n231), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n263), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n386) );
  AND2X2 AND2X2_5495 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n385), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n388), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n389) );
  AND2X2 AND2X2_5496 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n384), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n390), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n391) );
  AND2X2 AND2X2_5497 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n393), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n394), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n395) );
  AND2X2 AND2X2_5498 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n396), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n397), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n398) );
  AND2X2 AND2X2_5499 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n392), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n399), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_31_) );
  AND2X2 AND2X2_55 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n88), .B(\aes_mode[0] ), .Y(AES_CORE_CONTROL_UNIT_mode_cbc) );
  AND2X2 AND2X2_550 ( .A(AES_CORE_DATAPATH__abc_16259_n3403), .B(AES_CORE_DATAPATH__abc_16259_n3397), .Y(AES_CORE_DATAPATH__abc_16259_n3404_1) );
  AND2X2 AND2X2_5500 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n395), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n398), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n403) );
  AND2X2 AND2X2_5501 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n368), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n391), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n404) );
  AND2X2 AND2X2_5502 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n402), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n406), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n407) );
  AND2X2 AND2X2_5503 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n410), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n408), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_26_) );
  AND2X2 AND2X2_5504 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n212), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n412) );
  AND2X2 AND2X2_5505 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n415), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n414), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n416) );
  AND2X2 AND2X2_5506 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n419), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n418), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n420) );
  AND2X2 AND2X2_5507 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n417), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n421), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n422) );
  AND2X2 AND2X2_5508 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n395), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n422), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n423) );
  AND2X2 AND2X2_5509 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n424), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n425), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n426) );
  AND2X2 AND2X2_551 ( .A(AES_CORE_DATAPATH__abc_16259_n2837_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__14_), .Y(AES_CORE_DATAPATH__abc_16259_n3406) );
  AND2X2 AND2X2_5510 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n368), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n426), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n427) );
  AND2X2 AND2X2_5511 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n429), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n430), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n431) );
  AND2X2 AND2X2_5512 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n434), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n435), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n436) );
  AND2X2 AND2X2_5513 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n433), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n437), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_28_) );
  AND2X2 AND2X2_5514 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n432), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n439), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_27_) );
  AND2X2 AND2X2_5515 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n441), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n442), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n443) );
  AND2X2 AND2X2_5516 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n445), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n444), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_3_) );
  AND2X2 AND2X2_5517 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n447), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n448), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n449) );
  AND2X2 AND2X2_5518 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_28_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_29_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n451) );
  AND2X2 AND2X2_5519 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n431), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n401), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n452) );
  AND2X2 AND2X2_552 ( .A(AES_CORE_DATAPATH__abc_16259_n2887_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__14_), .Y(AES_CORE_DATAPATH__abc_16259_n3408) );
  AND2X2 AND2X2_5520 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n454), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n450), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_5_) );
  AND2X2 AND2X2_5521 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n457), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n456), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_6_) );
  AND2X2 AND2X2_5522 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n317), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n398), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n459) );
  AND2X2 AND2X2_5523 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n258), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n391), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n460) );
  AND2X2 AND2X2_5524 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n463), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n464), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_25_) );
  AND2X2 AND2X2_5525 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n467), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n466), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n468) );
  AND2X2 AND2X2_5526 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n126_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n469), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n470) );
  AND2X2 AND2X2_5527 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n472), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n473) );
  AND2X2 AND2X2_5528 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n469), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n474) );
  AND2X2 AND2X2_5529 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n471), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n475), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n476) );
  AND2X2 AND2X2_553 ( .A(AES_CORE_DATAPATH__abc_16259_n2830_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__14_), .Y(AES_CORE_DATAPATH__abc_16259_n3409_1) );
  AND2X2 AND2X2_5530 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n468), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n476), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n477) );
  AND2X2 AND2X2_5531 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n478) );
  AND2X2 AND2X2_5532 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n470), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n479), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n480) );
  AND2X2 AND2X2_5533 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n483), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n482), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n484) );
  AND2X2 AND2X2_5534 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n486), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n487) );
  AND2X2 AND2X2_5535 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n469), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n488) );
  AND2X2 AND2X2_5536 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n485), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n489), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n490) );
  AND2X2 AND2X2_5537 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n494), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n492), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n495) );
  AND2X2 AND2X2_5538 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n472), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n114), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n497) );
  AND2X2 AND2X2_5539 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n498), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n496), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n499) );
  AND2X2 AND2X2_554 ( .A(AES_CORE_DATAPATH__abc_16259_n3411), .B(AES_CORE_DATAPATH__abc_16259_n3412), .Y(_auto_iopadmap_cc_313_execute_26949_14_) );
  AND2X2 AND2X2_5540 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n499), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n495), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n500) );
  AND2X2 AND2X2_5541 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n491), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n500), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n501) );
  AND2X2 AND2X2_5542 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n502), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n503), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n504) );
  AND2X2 AND2X2_5543 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n505), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n481), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n506) );
  AND2X2 AND2X2_5544 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n504), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n507), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n508) );
  AND2X2 AND2X2_5545 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n114), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n512) );
  AND2X2 AND2X2_5546 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n513), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n511), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n514) );
  AND2X2 AND2X2_5547 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n515), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n510), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n516) );
  AND2X2 AND2X2_5548 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n514), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n475), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n517) );
  AND2X2 AND2X2_5549 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n519), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n520), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n521) );
  AND2X2 AND2X2_555 ( .A(AES_CORE_DATAPATH__abc_16259_n2855_bF_buf0), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_14_), .Y(AES_CORE_DATAPATH__abc_16259_n3415_1) );
  AND2X2 AND2X2_5550 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n522), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n523), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n524) );
  AND2X2 AND2X2_5551 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n521), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n525), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n526) );
  AND2X2 AND2X2_5552 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n468), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n524), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n527) );
  AND2X2 AND2X2_5553 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n528), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n518), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n529) );
  AND2X2 AND2X2_5554 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n521), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n510), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n530) );
  AND2X2 AND2X2_5555 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n530), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n479), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n531) );
  AND2X2 AND2X2_5556 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n532), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n478), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n533) );
  AND2X2 AND2X2_5557 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n534), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n490), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n535) );
  AND2X2 AND2X2_5558 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n536), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n537), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n538) );
  AND2X2 AND2X2_5559 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n538), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n491), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n539) );
  AND2X2 AND2X2_556 ( .A(AES_CORE_DATAPATH__abc_16259_n2857_bF_buf0), .B(AES_CORE_DATAPATH_MIX_COL_col_1__6_), .Y(AES_CORE_DATAPATH__abc_16259_n3416) );
  AND2X2 AND2X2_5560 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n543), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n544), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n545) );
  AND2X2 AND2X2_5561 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n541), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n546), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_stage1_1_) );
  AND2X2 AND2X2_5562 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n515), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n525), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n548) );
  AND2X2 AND2X2_5563 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n549) );
  AND2X2 AND2X2_5564 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n551), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n549), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n552) );
  AND2X2 AND2X2_5565 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n553), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n554), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n555) );
  AND2X2 AND2X2_5566 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n557), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n559), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n560) );
  AND2X2 AND2X2_5567 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n562), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n563), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n564) );
  AND2X2 AND2X2_5568 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n561), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n565), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_stage1_2_) );
  AND2X2 AND2X2_5569 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_7_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n569) );
  AND2X2 AND2X2_557 ( .A(AES_CORE_DATAPATH__abc_16259_n3414), .B(AES_CORE_DATAPATH__abc_16259_n3418), .Y(AES_CORE_DATAPATH__abc_16259_n3419_1) );
  AND2X2 AND2X2_5570 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n558), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n570), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n571) );
  AND2X2 AND2X2_5571 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n548), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n569), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n572) );
  AND2X2 AND2X2_5572 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n576), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n574), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n577) );
  AND2X2 AND2X2_5573 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n579), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n580), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_stage1_3_) );
  AND2X2 AND2X2_5574 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n584), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n582), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_2_) );
  AND2X2 AND2X2_5575 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n313), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n258), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n586) );
  AND2X2 AND2X2_5576 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n297), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n317), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n587) );
  AND2X2 AND2X2_5577 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n590), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n589), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_7_) );
  AND2X2 AND2X2_5578 ( .A(\data_type[1] ), .B(\data_type[0] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1) );
  AND2X2 AND2X2_5579 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1_bF_buf4), .B(\bus_in[31] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n68) );
  AND2X2 AND2X2_558 ( .A(_auto_iopadmap_cc_313_execute_26949_14_), .B(AES_CORE_DATAPATH__abc_16259_n3419_1), .Y(AES_CORE_DATAPATH__abc_16259_n3422) );
  AND2X2 AND2X2_5580 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n69), .B(\data_type[1] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70) );
  AND2X2 AND2X2_5581 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70_bF_buf4), .B(\bus_in[24] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n71_1) );
  AND2X2 AND2X2_5582 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n73), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n69), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74) );
  AND2X2 AND2X2_5583 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74_bF_buf4), .B(\bus_in[0] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n75) );
  AND2X2 AND2X2_5584 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n73), .B(\data_type[0] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1) );
  AND2X2 AND2X2_5585 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1_bF_buf4), .B(\bus_in[16] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n77_1) );
  AND2X2 AND2X2_5586 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1_bF_buf3), .B(\bus_in[30] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n80) );
  AND2X2 AND2X2_5587 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70_bF_buf3), .B(\bus_in[25] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n81_1) );
  AND2X2 AND2X2_5588 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74_bF_buf3), .B(\bus_in[1] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n83) );
  AND2X2 AND2X2_5589 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1_bF_buf3), .B(\bus_in[17] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n84) );
  AND2X2 AND2X2_559 ( .A(AES_CORE_DATAPATH_last_round_pp2_bF_buf4), .B(AES_CORE_DATAPATH_MIX_COL_col_1__6_), .Y(AES_CORE_DATAPATH__abc_16259_n3425) );
  AND2X2 AND2X2_5590 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1_bF_buf2), .B(\bus_in[29] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n87_1) );
  AND2X2 AND2X2_5591 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70_bF_buf2), .B(\bus_in[26] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n88) );
  AND2X2 AND2X2_5592 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74_bF_buf2), .B(\bus_in[2] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n90) );
  AND2X2 AND2X2_5593 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1_bF_buf2), .B(\bus_in[18] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n91_1) );
  AND2X2 AND2X2_5594 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1_bF_buf1), .B(\bus_in[28] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n94) );
  AND2X2 AND2X2_5595 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70_bF_buf1), .B(\bus_in[27] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n95) );
  AND2X2 AND2X2_5596 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74_bF_buf1), .B(\bus_in[3] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n97_1) );
  AND2X2 AND2X2_5597 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1_bF_buf1), .B(\bus_in[19] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n98) );
  AND2X2 AND2X2_5598 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1_bF_buf0), .B(\bus_in[27] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n101_1) );
  AND2X2 AND2X2_5599 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70_bF_buf0), .B(\bus_in[28] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n102_1) );
  AND2X2 AND2X2_56 ( .A(AES_CORE_CONTROL_UNIT_last_round_bF_buf3), .B(AES_CORE_CONTROL_UNIT_state_7_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n164) );
  AND2X2 AND2X2_560 ( .A(AES_CORE_DATAPATH__abc_16259_n2798_bF_buf0), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_14_), .Y(AES_CORE_DATAPATH__abc_16259_n3426) );
  AND2X2 AND2X2_5600 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74_bF_buf0), .B(\bus_in[4] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n104) );
  AND2X2 AND2X2_5601 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1_bF_buf0), .B(\bus_in[20] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n105) );
  AND2X2 AND2X2_5602 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1_bF_buf4), .B(\bus_in[26] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n108) );
  AND2X2 AND2X2_5603 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70_bF_buf4), .B(\bus_in[29] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n109) );
  AND2X2 AND2X2_5604 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74_bF_buf4), .B(\bus_in[5] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n111) );
  AND2X2 AND2X2_5605 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1_bF_buf4), .B(\bus_in[21] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n112) );
  AND2X2 AND2X2_5606 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1_bF_buf3), .B(\bus_in[25] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n115) );
  AND2X2 AND2X2_5607 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70_bF_buf3), .B(\bus_in[30] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n116) );
  AND2X2 AND2X2_5608 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74_bF_buf3), .B(\bus_in[6] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n118_1) );
  AND2X2 AND2X2_5609 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1_bF_buf3), .B(\bus_in[22] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n119) );
  AND2X2 AND2X2_561 ( .A(AES_CORE_DATAPATH__abc_16259_n3424), .B(AES_CORE_DATAPATH__abc_16259_n3428), .Y(AES_CORE_DATAPATH__abc_16259_n3429) );
  AND2X2 AND2X2_5610 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1_bF_buf2), .B(\bus_in[24] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n122_1) );
  AND2X2 AND2X2_5611 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70_bF_buf2), .B(\bus_in[31] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n123) );
  AND2X2 AND2X2_5612 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74_bF_buf2), .B(\bus_in[7] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n125) );
  AND2X2 AND2X2_5613 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1_bF_buf2), .B(\bus_in[23] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n126_1) );
  AND2X2 AND2X2_5614 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1_bF_buf1), .B(\bus_in[23] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n129) );
  AND2X2 AND2X2_5615 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70_bF_buf1), .B(\bus_in[16] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n130_1) );
  AND2X2 AND2X2_5616 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74_bF_buf1), .B(\bus_in[8] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n132) );
  AND2X2 AND2X2_5617 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1_bF_buf1), .B(\bus_in[24] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n133) );
  AND2X2 AND2X2_5618 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1_bF_buf0), .B(\bus_in[22] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n136) );
  AND2X2 AND2X2_5619 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70_bF_buf0), .B(\bus_in[17] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n137) );
  AND2X2 AND2X2_562 ( .A(AES_CORE_DATAPATH__abc_16259_n3429), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n3430) );
  AND2X2 AND2X2_5620 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74_bF_buf0), .B(\bus_in[9] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n139) );
  AND2X2 AND2X2_5621 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1_bF_buf0), .B(\bus_in[25] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n140) );
  AND2X2 AND2X2_5622 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1_bF_buf4), .B(\bus_in[21] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n143) );
  AND2X2 AND2X2_5623 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70_bF_buf4), .B(\bus_in[18] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n144) );
  AND2X2 AND2X2_5624 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74_bF_buf4), .B(\bus_in[10] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n146_1) );
  AND2X2 AND2X2_5625 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1_bF_buf4), .B(\bus_in[26] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n147) );
  AND2X2 AND2X2_5626 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1_bF_buf3), .B(\bus_in[20] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n150_1) );
  AND2X2 AND2X2_5627 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70_bF_buf3), .B(\bus_in[19] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n151) );
  AND2X2 AND2X2_5628 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74_bF_buf3), .B(\bus_in[11] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n153) );
  AND2X2 AND2X2_5629 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1_bF_buf3), .B(\bus_in[27] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n154_1) );
  AND2X2 AND2X2_563 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf10), .B(AES_CORE_DATAPATH_col_3__14_), .Y(AES_CORE_DATAPATH__abc_16259_n3431_1) );
  AND2X2 AND2X2_5630 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1_bF_buf2), .B(\bus_in[19] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n157) );
  AND2X2 AND2X2_5631 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70_bF_buf2), .B(\bus_in[20] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n158_1) );
  AND2X2 AND2X2_5632 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74_bF_buf2), .B(\bus_in[12] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n160) );
  AND2X2 AND2X2_5633 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1_bF_buf2), .B(\bus_in[28] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n161) );
  AND2X2 AND2X2_5634 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1_bF_buf1), .B(\bus_in[18] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n164) );
  AND2X2 AND2X2_5635 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70_bF_buf1), .B(\bus_in[21] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n165) );
  AND2X2 AND2X2_5636 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74_bF_buf1), .B(\bus_in[13] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n167) );
  AND2X2 AND2X2_5637 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1_bF_buf1), .B(\bus_in[29] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n168) );
  AND2X2 AND2X2_5638 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1_bF_buf0), .B(\bus_in[17] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n171) );
  AND2X2 AND2X2_5639 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70_bF_buf0), .B(\bus_in[22] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n172) );
  AND2X2 AND2X2_564 ( .A(AES_CORE_DATAPATH__abc_16259_n3434), .B(AES_CORE_DATAPATH__abc_16259_n3436), .Y(AES_CORE_DATAPATH__abc_16259_n3437) );
  AND2X2 AND2X2_5640 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74_bF_buf0), .B(\bus_in[14] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n174) );
  AND2X2 AND2X2_5641 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1_bF_buf0), .B(\bus_in[30] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n175) );
  AND2X2 AND2X2_5642 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1_bF_buf4), .B(\bus_in[16] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n178) );
  AND2X2 AND2X2_5643 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70_bF_buf4), .B(\bus_in[23] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n179) );
  AND2X2 AND2X2_5644 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74_bF_buf4), .B(\bus_in[15] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n181) );
  AND2X2 AND2X2_5645 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1_bF_buf4), .B(\bus_in[31] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n182) );
  AND2X2 AND2X2_5646 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1_bF_buf3), .B(\bus_in[15] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n185) );
  AND2X2 AND2X2_5647 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70_bF_buf3), .B(\bus_in[8] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n186) );
  AND2X2 AND2X2_5648 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74_bF_buf3), .B(\bus_in[16] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n188) );
  AND2X2 AND2X2_5649 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1_bF_buf3), .B(\bus_in[0] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n189) );
  AND2X2 AND2X2_565 ( .A(AES_CORE_DATAPATH__abc_16259_n2782_bF_buf4), .B(AES_CORE_DATAPATH_col_3__15_), .Y(AES_CORE_DATAPATH__abc_16259_n3438_1) );
  AND2X2 AND2X2_5650 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1_bF_buf2), .B(\bus_in[14] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n192) );
  AND2X2 AND2X2_5651 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70_bF_buf2), .B(\bus_in[9] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n193) );
  AND2X2 AND2X2_5652 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74_bF_buf2), .B(\bus_in[17] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n195) );
  AND2X2 AND2X2_5653 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1_bF_buf2), .B(\bus_in[1] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n196) );
  AND2X2 AND2X2_5654 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1_bF_buf1), .B(\bus_in[13] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n199) );
  AND2X2 AND2X2_5655 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70_bF_buf1), .B(\bus_in[10] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n200) );
  AND2X2 AND2X2_5656 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74_bF_buf1), .B(\bus_in[18] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n202) );
  AND2X2 AND2X2_5657 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1_bF_buf1), .B(\bus_in[2] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n203) );
  AND2X2 AND2X2_5658 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1_bF_buf0), .B(\bus_in[12] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n206) );
  AND2X2 AND2X2_5659 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70_bF_buf0), .B(\bus_in[11] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n207) );
  AND2X2 AND2X2_566 ( .A(AES_CORE_DATAPATH__abc_16259_n2786_bF_buf4), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_79_), .Y(AES_CORE_DATAPATH__abc_16259_n3439_1) );
  AND2X2 AND2X2_5660 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74_bF_buf0), .B(\bus_in[19] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n209) );
  AND2X2 AND2X2_5661 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1_bF_buf0), .B(\bus_in[3] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n210) );
  AND2X2 AND2X2_5662 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1_bF_buf4), .B(\bus_in[11] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n213) );
  AND2X2 AND2X2_5663 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70_bF_buf4), .B(\bus_in[12] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n214) );
  AND2X2 AND2X2_5664 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74_bF_buf4), .B(\bus_in[20] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n216) );
  AND2X2 AND2X2_5665 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1_bF_buf4), .B(\bus_in[4] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n217) );
  AND2X2 AND2X2_5666 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1_bF_buf3), .B(\bus_in[10] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n220) );
  AND2X2 AND2X2_5667 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70_bF_buf3), .B(\bus_in[13] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n221) );
  AND2X2 AND2X2_5668 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74_bF_buf3), .B(\bus_in[21] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n223) );
  AND2X2 AND2X2_5669 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1_bF_buf3), .B(\bus_in[5] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n224) );
  AND2X2 AND2X2_567 ( .A(AES_CORE_DATAPATH__abc_16259_n2789_bF_buf4), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_47_), .Y(AES_CORE_DATAPATH__abc_16259_n3440) );
  AND2X2 AND2X2_5670 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1_bF_buf2), .B(\bus_in[9] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n227) );
  AND2X2 AND2X2_5671 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70_bF_buf2), .B(\bus_in[14] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n228) );
  AND2X2 AND2X2_5672 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74_bF_buf2), .B(\bus_in[22] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n230) );
  AND2X2 AND2X2_5673 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1_bF_buf2), .B(\bus_in[6] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n231) );
  AND2X2 AND2X2_5674 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1_bF_buf1), .B(\bus_in[8] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n234) );
  AND2X2 AND2X2_5675 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70_bF_buf1), .B(\bus_in[15] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n235) );
  AND2X2 AND2X2_5676 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74_bF_buf1), .B(\bus_in[23] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n237) );
  AND2X2 AND2X2_5677 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1_bF_buf1), .B(\bus_in[7] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n238) );
  AND2X2 AND2X2_5678 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1_bF_buf0), .B(\bus_in[7] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n241) );
  AND2X2 AND2X2_5679 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70_bF_buf0), .B(\bus_in[0] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n242) );
  AND2X2 AND2X2_568 ( .A(AES_CORE_DATAPATH__abc_16259_n3443), .B(AES_CORE_DATAPATH__abc_16259_n3437), .Y(AES_CORE_DATAPATH__abc_16259_n3444_1) );
  AND2X2 AND2X2_5680 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74_bF_buf0), .B(\bus_in[24] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n244) );
  AND2X2 AND2X2_5681 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1_bF_buf0), .B(\bus_in[8] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n245) );
  AND2X2 AND2X2_5682 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1_bF_buf4), .B(\bus_in[6] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n248) );
  AND2X2 AND2X2_5683 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70_bF_buf4), .B(\bus_in[1] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n249) );
  AND2X2 AND2X2_5684 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74_bF_buf4), .B(\bus_in[25] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n251) );
  AND2X2 AND2X2_5685 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1_bF_buf4), .B(\bus_in[9] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n252) );
  AND2X2 AND2X2_5686 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1_bF_buf3), .B(\bus_in[5] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n255) );
  AND2X2 AND2X2_5687 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70_bF_buf3), .B(\bus_in[2] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n256) );
  AND2X2 AND2X2_5688 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74_bF_buf3), .B(\bus_in[26] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n258) );
  AND2X2 AND2X2_5689 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1_bF_buf3), .B(\bus_in[10] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n259) );
  AND2X2 AND2X2_569 ( .A(AES_CORE_DATAPATH__abc_16259_n2837_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__15_), .Y(AES_CORE_DATAPATH__abc_16259_n3446_1) );
  AND2X2 AND2X2_5690 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1_bF_buf2), .B(\bus_in[4] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n262) );
  AND2X2 AND2X2_5691 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70_bF_buf2), .B(\bus_in[3] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n263) );
  AND2X2 AND2X2_5692 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74_bF_buf2), .B(\bus_in[27] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n265) );
  AND2X2 AND2X2_5693 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1_bF_buf2), .B(\bus_in[11] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n266) );
  AND2X2 AND2X2_5694 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1_bF_buf1), .B(\bus_in[3] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n269) );
  AND2X2 AND2X2_5695 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70_bF_buf1), .B(\bus_in[4] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n270) );
  AND2X2 AND2X2_5696 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74_bF_buf1), .B(\bus_in[28] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n272) );
  AND2X2 AND2X2_5697 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1_bF_buf1), .B(\bus_in[12] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n273) );
  AND2X2 AND2X2_5698 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1_bF_buf0), .B(\bus_in[2] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n276) );
  AND2X2 AND2X2_5699 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70_bF_buf0), .B(\bus_in[5] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n277) );
  AND2X2 AND2X2_57 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n165), .B(AES_CORE_CONTROL_UNIT__abc_15841_n163), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n166) );
  AND2X2 AND2X2_570 ( .A(AES_CORE_DATAPATH__abc_16259_n2887_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__15_), .Y(AES_CORE_DATAPATH__abc_16259_n3448_1) );
  AND2X2 AND2X2_5700 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74_bF_buf0), .B(\bus_in[29] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n279) );
  AND2X2 AND2X2_5701 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1_bF_buf0), .B(\bus_in[13] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n280) );
  AND2X2 AND2X2_5702 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1_bF_buf4), .B(\bus_in[1] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n283) );
  AND2X2 AND2X2_5703 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70_bF_buf4), .B(\bus_in[6] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n284) );
  AND2X2 AND2X2_5704 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74_bF_buf4), .B(\bus_in[30] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n286) );
  AND2X2 AND2X2_5705 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1_bF_buf4), .B(\bus_in[14] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n287) );
  AND2X2 AND2X2_5706 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1_bF_buf3), .B(\bus_in[0] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n290) );
  AND2X2 AND2X2_5707 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70_bF_buf3), .B(\bus_in[7] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n291) );
  AND2X2 AND2X2_5708 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74_bF_buf3), .B(\bus_in[31] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n293) );
  AND2X2 AND2X2_5709 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1_bF_buf3), .B(\bus_in[15] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n294) );
  AND2X2 AND2X2_571 ( .A(AES_CORE_DATAPATH__abc_16259_n2830_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__15_), .Y(AES_CORE_DATAPATH__abc_16259_n3449) );
  AND2X2 AND2X2_5710 ( .A(\data_type[1] ), .B(\data_type[0] ), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1) );
  AND2X2 AND2X2_5711 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1_bF_buf4), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_7_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n68) );
  AND2X2 AND2X2_5712 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n69), .B(\data_type[1] ), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70) );
  AND2X2 AND2X2_5713 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70_bF_buf4), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_0_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n71_1) );
  AND2X2 AND2X2_5714 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n73), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n69), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74) );
  AND2X2 AND2X2_5715 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74_bF_buf4), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_0_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n75) );
  AND2X2 AND2X2_5716 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n73), .B(\data_type[0] ), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1) );
  AND2X2 AND2X2_5717 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1_bF_buf4), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_0_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n77_1) );
  AND2X2 AND2X2_5718 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1_bF_buf3), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_6_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n80) );
  AND2X2 AND2X2_5719 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70_bF_buf3), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_1_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n81_1) );
  AND2X2 AND2X2_572 ( .A(AES_CORE_DATAPATH__abc_16259_n3451), .B(AES_CORE_DATAPATH__abc_16259_n3452), .Y(_auto_iopadmap_cc_313_execute_26949_15_) );
  AND2X2 AND2X2_5720 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74_bF_buf3), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_1_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n83) );
  AND2X2 AND2X2_5721 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1_bF_buf3), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_1_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n84) );
  AND2X2 AND2X2_5722 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1_bF_buf2), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_5_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n87_1) );
  AND2X2 AND2X2_5723 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70_bF_buf2), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_2_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n88) );
  AND2X2 AND2X2_5724 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74_bF_buf2), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_2_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n90) );
  AND2X2 AND2X2_5725 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1_bF_buf2), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_2_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n91_1) );
  AND2X2 AND2X2_5726 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1_bF_buf1), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_4_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n94) );
  AND2X2 AND2X2_5727 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70_bF_buf1), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_3_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n95) );
  AND2X2 AND2X2_5728 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74_bF_buf1), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_3_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n97_1) );
  AND2X2 AND2X2_5729 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1_bF_buf1), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_3_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n98) );
  AND2X2 AND2X2_573 ( .A(AES_CORE_DATAPATH__abc_16259_n2855_bF_buf4), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_15_), .Y(AES_CORE_DATAPATH__abc_16259_n3455) );
  AND2X2 AND2X2_5730 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1_bF_buf0), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_3_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n101_1) );
  AND2X2 AND2X2_5731 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70_bF_buf0), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_4_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n102_1) );
  AND2X2 AND2X2_5732 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74_bF_buf0), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_4_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n104) );
  AND2X2 AND2X2_5733 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1_bF_buf0), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_4_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n105) );
  AND2X2 AND2X2_5734 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1_bF_buf4), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_2_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n108) );
  AND2X2 AND2X2_5735 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70_bF_buf4), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_5_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n109) );
  AND2X2 AND2X2_5736 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74_bF_buf4), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_5_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n111) );
  AND2X2 AND2X2_5737 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1_bF_buf4), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_5_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n112) );
  AND2X2 AND2X2_5738 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1_bF_buf3), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_1_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n115) );
  AND2X2 AND2X2_5739 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70_bF_buf3), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_6_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n116) );
  AND2X2 AND2X2_574 ( .A(AES_CORE_DATAPATH__abc_16259_n2857_bF_buf4), .B(AES_CORE_DATAPATH_MIX_COL_col_1__7_), .Y(AES_CORE_DATAPATH__abc_16259_n3456) );
  AND2X2 AND2X2_5740 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74_bF_buf3), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_6_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n118_1) );
  AND2X2 AND2X2_5741 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1_bF_buf3), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_6_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n119) );
  AND2X2 AND2X2_5742 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1_bF_buf2), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_0_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n122_1) );
  AND2X2 AND2X2_5743 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70_bF_buf2), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_7_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n123) );
  AND2X2 AND2X2_5744 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74_bF_buf2), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_7_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n125) );
  AND2X2 AND2X2_5745 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1_bF_buf2), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_7_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n126_1) );
  AND2X2 AND2X2_5746 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1_bF_buf1), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_7_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n129) );
  AND2X2 AND2X2_5747 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70_bF_buf1), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_0_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n130_1) );
  AND2X2 AND2X2_5748 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74_bF_buf1), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_0_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n132) );
  AND2X2 AND2X2_5749 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1_bF_buf1), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_0_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n133) );
  AND2X2 AND2X2_575 ( .A(AES_CORE_DATAPATH__abc_16259_n3454), .B(AES_CORE_DATAPATH__abc_16259_n3458), .Y(AES_CORE_DATAPATH__abc_16259_n3459) );
  AND2X2 AND2X2_5750 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1_bF_buf0), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_6_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n136) );
  AND2X2 AND2X2_5751 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70_bF_buf0), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_1_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n137) );
  AND2X2 AND2X2_5752 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74_bF_buf0), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_1_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n139) );
  AND2X2 AND2X2_5753 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1_bF_buf0), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_1_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n140) );
  AND2X2 AND2X2_5754 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1_bF_buf4), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_5_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n143) );
  AND2X2 AND2X2_5755 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70_bF_buf4), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_2_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n144) );
  AND2X2 AND2X2_5756 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74_bF_buf4), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_2_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n146_1) );
  AND2X2 AND2X2_5757 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1_bF_buf4), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_2_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n147) );
  AND2X2 AND2X2_5758 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1_bF_buf3), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_4_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n150_1) );
  AND2X2 AND2X2_5759 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70_bF_buf3), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_3_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n151) );
  AND2X2 AND2X2_576 ( .A(_auto_iopadmap_cc_313_execute_26949_15_), .B(AES_CORE_DATAPATH__abc_16259_n3459), .Y(AES_CORE_DATAPATH__abc_16259_n3462_1) );
  AND2X2 AND2X2_5760 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74_bF_buf3), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_3_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n153) );
  AND2X2 AND2X2_5761 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1_bF_buf3), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_3_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n154_1) );
  AND2X2 AND2X2_5762 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1_bF_buf2), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_3_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n157) );
  AND2X2 AND2X2_5763 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70_bF_buf2), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_4_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n158_1) );
  AND2X2 AND2X2_5764 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74_bF_buf2), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_4_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n160) );
  AND2X2 AND2X2_5765 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1_bF_buf2), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_4_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n161) );
  AND2X2 AND2X2_5766 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1_bF_buf1), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_2_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n164) );
  AND2X2 AND2X2_5767 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70_bF_buf1), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_5_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n165) );
  AND2X2 AND2X2_5768 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74_bF_buf1), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_5_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n167) );
  AND2X2 AND2X2_5769 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1_bF_buf1), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_5_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n168) );
  AND2X2 AND2X2_577 ( .A(AES_CORE_DATAPATH_last_round_pp2_bF_buf3), .B(AES_CORE_DATAPATH_MIX_COL_col_1__7_), .Y(AES_CORE_DATAPATH__abc_16259_n3465) );
  AND2X2 AND2X2_5770 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1_bF_buf0), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_1_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n171) );
  AND2X2 AND2X2_5771 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70_bF_buf0), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_6_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n172) );
  AND2X2 AND2X2_5772 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74_bF_buf0), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_6_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n174) );
  AND2X2 AND2X2_5773 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1_bF_buf0), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_6_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n175) );
  AND2X2 AND2X2_5774 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1_bF_buf4), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_0_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n178) );
  AND2X2 AND2X2_5775 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70_bF_buf4), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_7_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n179) );
  AND2X2 AND2X2_5776 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74_bF_buf4), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_7_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n181) );
  AND2X2 AND2X2_5777 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1_bF_buf4), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_7_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n182) );
  AND2X2 AND2X2_5778 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1_bF_buf3), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_7_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n185) );
  AND2X2 AND2X2_5779 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70_bF_buf3), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_0_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n186) );
  AND2X2 AND2X2_578 ( .A(AES_CORE_DATAPATH__abc_16259_n2798_bF_buf4), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_15_), .Y(AES_CORE_DATAPATH__abc_16259_n3466) );
  AND2X2 AND2X2_5780 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74_bF_buf3), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_0_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n188) );
  AND2X2 AND2X2_5781 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1_bF_buf3), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_0_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n189) );
  AND2X2 AND2X2_5782 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1_bF_buf2), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_6_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n192) );
  AND2X2 AND2X2_5783 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70_bF_buf2), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_1_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n193) );
  AND2X2 AND2X2_5784 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74_bF_buf2), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_1_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n195) );
  AND2X2 AND2X2_5785 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1_bF_buf2), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_1_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n196) );
  AND2X2 AND2X2_5786 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1_bF_buf1), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_5_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n199) );
  AND2X2 AND2X2_5787 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70_bF_buf1), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_2_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n200) );
  AND2X2 AND2X2_5788 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74_bF_buf1), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_2_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n202) );
  AND2X2 AND2X2_5789 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1_bF_buf1), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_2_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n203) );
  AND2X2 AND2X2_579 ( .A(AES_CORE_DATAPATH__abc_16259_n3464), .B(AES_CORE_DATAPATH__abc_16259_n3468_1), .Y(AES_CORE_DATAPATH__abc_16259_n3469) );
  AND2X2 AND2X2_5790 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1_bF_buf0), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_4_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n206) );
  AND2X2 AND2X2_5791 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70_bF_buf0), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_3_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n207) );
  AND2X2 AND2X2_5792 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74_bF_buf0), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_3_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n209) );
  AND2X2 AND2X2_5793 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1_bF_buf0), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_3_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n210) );
  AND2X2 AND2X2_5794 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1_bF_buf4), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_3_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n213) );
  AND2X2 AND2X2_5795 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70_bF_buf4), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_4_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n214) );
  AND2X2 AND2X2_5796 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74_bF_buf4), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_4_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n216) );
  AND2X2 AND2X2_5797 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1_bF_buf4), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_4_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n217) );
  AND2X2 AND2X2_5798 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1_bF_buf3), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_2_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n220) );
  AND2X2 AND2X2_5799 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70_bF_buf3), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_5_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n221) );
  AND2X2 AND2X2_58 ( .A(AES_CORE_CONTROL_UNIT_sbox_sel_2_), .B(AES_CORE_CONTROL_UNIT_rd_count_0_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n169) );
  AND2X2 AND2X2_580 ( .A(AES_CORE_DATAPATH__abc_16259_n3469), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n3470) );
  AND2X2 AND2X2_5800 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74_bF_buf3), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_5_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n223) );
  AND2X2 AND2X2_5801 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1_bF_buf3), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_5_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n224) );
  AND2X2 AND2X2_5802 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1_bF_buf2), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_1_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n227) );
  AND2X2 AND2X2_5803 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70_bF_buf2), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_6_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n228) );
  AND2X2 AND2X2_5804 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74_bF_buf2), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_6_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n230) );
  AND2X2 AND2X2_5805 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1_bF_buf2), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_6_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n231) );
  AND2X2 AND2X2_5806 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1_bF_buf1), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_0_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n234) );
  AND2X2 AND2X2_5807 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70_bF_buf1), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_7_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n235) );
  AND2X2 AND2X2_5808 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74_bF_buf1), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_7_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n237) );
  AND2X2 AND2X2_5809 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1_bF_buf1), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_7_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n238) );
  AND2X2 AND2X2_581 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf9), .B(AES_CORE_DATAPATH_col_3__15_), .Y(AES_CORE_DATAPATH__abc_16259_n3471_1) );
  AND2X2 AND2X2_5810 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1_bF_buf0), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_7_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n241) );
  AND2X2 AND2X2_5811 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70_bF_buf0), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_0_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n242) );
  AND2X2 AND2X2_5812 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74_bF_buf0), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_0_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n244) );
  AND2X2 AND2X2_5813 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1_bF_buf0), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_0_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n245) );
  AND2X2 AND2X2_5814 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1_bF_buf4), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_6_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n248) );
  AND2X2 AND2X2_5815 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70_bF_buf4), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_1_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n249) );
  AND2X2 AND2X2_5816 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74_bF_buf4), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_1_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n251) );
  AND2X2 AND2X2_5817 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1_bF_buf4), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_1_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n252) );
  AND2X2 AND2X2_5818 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1_bF_buf3), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_5_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n255) );
  AND2X2 AND2X2_5819 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70_bF_buf3), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_2_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n256) );
  AND2X2 AND2X2_582 ( .A(AES_CORE_DATAPATH__abc_16259_n3474), .B(AES_CORE_DATAPATH__abc_16259_n3476), .Y(AES_CORE_DATAPATH__abc_16259_n3477_1) );
  AND2X2 AND2X2_5820 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74_bF_buf3), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_2_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n258) );
  AND2X2 AND2X2_5821 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1_bF_buf3), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_2_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n259) );
  AND2X2 AND2X2_5822 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1_bF_buf2), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_4_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n262) );
  AND2X2 AND2X2_5823 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70_bF_buf2), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_3_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n263) );
  AND2X2 AND2X2_5824 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74_bF_buf2), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_3_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n265) );
  AND2X2 AND2X2_5825 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1_bF_buf2), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_3_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n266) );
  AND2X2 AND2X2_5826 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1_bF_buf1), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_3_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n269) );
  AND2X2 AND2X2_5827 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70_bF_buf1), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_4_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n270) );
  AND2X2 AND2X2_5828 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74_bF_buf1), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_4_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n272) );
  AND2X2 AND2X2_5829 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1_bF_buf1), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_4_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n273) );
  AND2X2 AND2X2_583 ( .A(AES_CORE_DATAPATH__abc_16259_n2782_bF_buf3), .B(AES_CORE_DATAPATH_col_3__16_), .Y(AES_CORE_DATAPATH__abc_16259_n3478) );
  AND2X2 AND2X2_5830 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1_bF_buf0), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_2_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n276) );
  AND2X2 AND2X2_5831 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70_bF_buf0), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_5_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n277) );
  AND2X2 AND2X2_5832 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74_bF_buf0), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_5_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n279) );
  AND2X2 AND2X2_5833 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1_bF_buf0), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_5_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n280) );
  AND2X2 AND2X2_5834 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1_bF_buf4), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_1_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n283) );
  AND2X2 AND2X2_5835 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70_bF_buf4), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_6_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n284) );
  AND2X2 AND2X2_5836 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74_bF_buf4), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_6_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n286) );
  AND2X2 AND2X2_5837 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1_bF_buf4), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_6_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n287) );
  AND2X2 AND2X2_5838 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1_bF_buf3), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_0_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n290) );
  AND2X2 AND2X2_5839 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70_bF_buf3), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_7_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n291) );
  AND2X2 AND2X2_584 ( .A(AES_CORE_DATAPATH__abc_16259_n2786_bF_buf3), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_80_), .Y(AES_CORE_DATAPATH__abc_16259_n3479) );
  AND2X2 AND2X2_5840 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74_bF_buf3), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_7_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n293) );
  AND2X2 AND2X2_5841 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1_bF_buf3), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_7_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n294) );
  AND2X2 AND2X2_585 ( .A(AES_CORE_DATAPATH__abc_16259_n2789_bF_buf3), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_48_), .Y(AES_CORE_DATAPATH__abc_16259_n3480) );
  AND2X2 AND2X2_586 ( .A(AES_CORE_DATAPATH__abc_16259_n3483), .B(AES_CORE_DATAPATH__abc_16259_n3477_1), .Y(AES_CORE_DATAPATH__abc_16259_n3484) );
  AND2X2 AND2X2_587 ( .A(AES_CORE_DATAPATH__abc_16259_n2837_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__16_), .Y(AES_CORE_DATAPATH__abc_16259_n3486) );
  AND2X2 AND2X2_588 ( .A(AES_CORE_DATAPATH__abc_16259_n2887_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__16_), .Y(AES_CORE_DATAPATH__abc_16259_n3488) );
  AND2X2 AND2X2_589 ( .A(AES_CORE_DATAPATH__abc_16259_n2830_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__16_), .Y(AES_CORE_DATAPATH__abc_16259_n3489_1) );
  AND2X2 AND2X2_59 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n170), .B(AES_CORE_CONTROL_UNIT__abc_15841_n168), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n171_1) );
  AND2X2 AND2X2_590 ( .A(AES_CORE_DATAPATH__abc_16259_n3491_1), .B(AES_CORE_DATAPATH__abc_16259_n3492), .Y(_auto_iopadmap_cc_313_execute_26949_16_) );
  AND2X2 AND2X2_591 ( .A(AES_CORE_DATAPATH__abc_16259_n2855_bF_buf3), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_16_), .Y(AES_CORE_DATAPATH__abc_16259_n3495) );
  AND2X2 AND2X2_592 ( .A(AES_CORE_DATAPATH__abc_16259_n2857_bF_buf3), .B(AES_CORE_DATAPATH_MIX_COL_col_2__0_), .Y(AES_CORE_DATAPATH__abc_16259_n3496_1) );
  AND2X2 AND2X2_593 ( .A(AES_CORE_DATAPATH__abc_16259_n3494), .B(AES_CORE_DATAPATH__abc_16259_n3498), .Y(AES_CORE_DATAPATH__abc_16259_n3499) );
  AND2X2 AND2X2_594 ( .A(_auto_iopadmap_cc_313_execute_26949_16_), .B(AES_CORE_DATAPATH__abc_16259_n3499), .Y(AES_CORE_DATAPATH__abc_16259_n3502_1) );
  AND2X2 AND2X2_595 ( .A(AES_CORE_DATAPATH_last_round_pp2_bF_buf2), .B(AES_CORE_DATAPATH_MIX_COL_col_2__0_), .Y(AES_CORE_DATAPATH__abc_16259_n3505) );
  AND2X2 AND2X2_596 ( .A(AES_CORE_DATAPATH__abc_16259_n2798_bF_buf3), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_16_), .Y(AES_CORE_DATAPATH__abc_16259_n3506_1) );
  AND2X2 AND2X2_597 ( .A(AES_CORE_DATAPATH__abc_16259_n3504_1), .B(AES_CORE_DATAPATH__abc_16259_n3508), .Y(AES_CORE_DATAPATH__abc_16259_n3509) );
  AND2X2 AND2X2_598 ( .A(AES_CORE_DATAPATH__abc_16259_n3509), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n3510) );
  AND2X2 AND2X2_599 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf8), .B(AES_CORE_DATAPATH_col_3__16_), .Y(AES_CORE_DATAPATH__abc_16259_n3511) );
  AND2X2 AND2X2_6 ( .A(_abc_15830_n15), .B(\addr[1] ), .Y(AES_CORE_DATAPATH_col_en_host_3_) );
  AND2X2 AND2X2_60 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n166), .B(AES_CORE_CONTROL_UNIT__abc_15841_n171_1), .Y(AES_CORE_CONTROL_UNIT_rd_count_0__FF_INPUT) );
  AND2X2 AND2X2_600 ( .A(AES_CORE_DATAPATH__abc_16259_n3514), .B(AES_CORE_DATAPATH__abc_16259_n3516), .Y(AES_CORE_DATAPATH__abc_16259_n3517) );
  AND2X2 AND2X2_601 ( .A(AES_CORE_DATAPATH__abc_16259_n2782_bF_buf2), .B(AES_CORE_DATAPATH_col_3__17_), .Y(AES_CORE_DATAPATH__abc_16259_n3518_1) );
  AND2X2 AND2X2_602 ( .A(AES_CORE_DATAPATH__abc_16259_n2786_bF_buf2), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_81_), .Y(AES_CORE_DATAPATH__abc_16259_n3519) );
  AND2X2 AND2X2_603 ( .A(AES_CORE_DATAPATH__abc_16259_n2789_bF_buf2), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_49_), .Y(AES_CORE_DATAPATH__abc_16259_n3520_1) );
  AND2X2 AND2X2_604 ( .A(AES_CORE_DATAPATH__abc_16259_n3523), .B(AES_CORE_DATAPATH__abc_16259_n3517), .Y(AES_CORE_DATAPATH__abc_16259_n3524) );
  AND2X2 AND2X2_605 ( .A(AES_CORE_DATAPATH__abc_16259_n2837_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__17_), .Y(AES_CORE_DATAPATH__abc_16259_n3526_1) );
  AND2X2 AND2X2_606 ( .A(AES_CORE_DATAPATH__abc_16259_n2887_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__17_), .Y(AES_CORE_DATAPATH__abc_16259_n3528) );
  AND2X2 AND2X2_607 ( .A(AES_CORE_DATAPATH__abc_16259_n2830_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__17_), .Y(AES_CORE_DATAPATH__abc_16259_n3529_1) );
  AND2X2 AND2X2_608 ( .A(AES_CORE_DATAPATH__abc_16259_n3531_1), .B(AES_CORE_DATAPATH__abc_16259_n3532), .Y(_auto_iopadmap_cc_313_execute_26949_17_) );
  AND2X2 AND2X2_609 ( .A(AES_CORE_DATAPATH__abc_16259_n2855_bF_buf2), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_17_), .Y(AES_CORE_DATAPATH__abc_16259_n3535_1) );
  AND2X2 AND2X2_61 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n169), .B(AES_CORE_CONTROL_UNIT_rd_count_1_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n173) );
  AND2X2 AND2X2_610 ( .A(AES_CORE_DATAPATH__abc_16259_n2857_bF_buf2), .B(AES_CORE_DATAPATH_MIX_COL_col_2__1_), .Y(AES_CORE_DATAPATH__abc_16259_n3536) );
  AND2X2 AND2X2_611 ( .A(AES_CORE_DATAPATH__abc_16259_n3534), .B(AES_CORE_DATAPATH__abc_16259_n3538), .Y(AES_CORE_DATAPATH__abc_16259_n3539) );
  AND2X2 AND2X2_612 ( .A(_auto_iopadmap_cc_313_execute_26949_17_), .B(AES_CORE_DATAPATH__abc_16259_n3539), .Y(AES_CORE_DATAPATH__abc_16259_n3542) );
  AND2X2 AND2X2_613 ( .A(AES_CORE_DATAPATH_last_round_pp2_bF_buf1), .B(AES_CORE_DATAPATH_MIX_COL_col_2__1_), .Y(AES_CORE_DATAPATH__abc_16259_n3545) );
  AND2X2 AND2X2_614 ( .A(AES_CORE_DATAPATH__abc_16259_n2798_bF_buf2), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_17_), .Y(AES_CORE_DATAPATH__abc_16259_n3546) );
  AND2X2 AND2X2_615 ( .A(AES_CORE_DATAPATH__abc_16259_n3544), .B(AES_CORE_DATAPATH__abc_16259_n3548), .Y(AES_CORE_DATAPATH__abc_16259_n3549_1) );
  AND2X2 AND2X2_616 ( .A(AES_CORE_DATAPATH__abc_16259_n3549_1), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n3550) );
  AND2X2 AND2X2_617 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf7), .B(AES_CORE_DATAPATH_col_3__17_), .Y(AES_CORE_DATAPATH__abc_16259_n3551) );
  AND2X2 AND2X2_618 ( .A(AES_CORE_DATAPATH__abc_16259_n3554_1), .B(AES_CORE_DATAPATH__abc_16259_n3556), .Y(AES_CORE_DATAPATH__abc_16259_n3557) );
  AND2X2 AND2X2_619 ( .A(AES_CORE_DATAPATH__abc_16259_n2782_bF_buf1), .B(AES_CORE_DATAPATH_col_3__18_), .Y(AES_CORE_DATAPATH__abc_16259_n3558_1) );
  AND2X2 AND2X2_62 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n174), .B(AES_CORE_CONTROL_UNIT__abc_15841_n175_1), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n176) );
  AND2X2 AND2X2_620 ( .A(AES_CORE_DATAPATH__abc_16259_n2786_bF_buf1), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_82_), .Y(AES_CORE_DATAPATH__abc_16259_n3559) );
  AND2X2 AND2X2_621 ( .A(AES_CORE_DATAPATH__abc_16259_n2789_bF_buf1), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_50_), .Y(AES_CORE_DATAPATH__abc_16259_n3560_1) );
  AND2X2 AND2X2_622 ( .A(AES_CORE_DATAPATH__abc_16259_n3563), .B(AES_CORE_DATAPATH__abc_16259_n3557), .Y(AES_CORE_DATAPATH__abc_16259_n3564_1) );
  AND2X2 AND2X2_623 ( .A(AES_CORE_DATAPATH__abc_16259_n2837_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__18_), .Y(AES_CORE_DATAPATH__abc_16259_n3566) );
  AND2X2 AND2X2_624 ( .A(AES_CORE_DATAPATH__abc_16259_n2887_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__18_), .Y(AES_CORE_DATAPATH__abc_16259_n3568) );
  AND2X2 AND2X2_625 ( .A(AES_CORE_DATAPATH__abc_16259_n2830_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__18_), .Y(AES_CORE_DATAPATH__abc_16259_n3569) );
  AND2X2 AND2X2_626 ( .A(AES_CORE_DATAPATH__abc_16259_n3571), .B(AES_CORE_DATAPATH__abc_16259_n3572), .Y(_auto_iopadmap_cc_313_execute_26949_18_) );
  AND2X2 AND2X2_627 ( .A(AES_CORE_DATAPATH__abc_16259_n2855_bF_buf1), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_18_), .Y(AES_CORE_DATAPATH__abc_16259_n3575) );
  AND2X2 AND2X2_628 ( .A(AES_CORE_DATAPATH__abc_16259_n2857_bF_buf1), .B(AES_CORE_DATAPATH_MIX_COL_col_2__2_), .Y(AES_CORE_DATAPATH__abc_16259_n3576_1) );
  AND2X2 AND2X2_629 ( .A(AES_CORE_DATAPATH__abc_16259_n3574), .B(AES_CORE_DATAPATH__abc_16259_n3578_1), .Y(AES_CORE_DATAPATH__abc_16259_n3579) );
  AND2X2 AND2X2_63 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n176), .B(AES_CORE_CONTROL_UNIT__abc_15841_n166), .Y(AES_CORE_CONTROL_UNIT_rd_count_1__FF_INPUT) );
  AND2X2 AND2X2_630 ( .A(_auto_iopadmap_cc_313_execute_26949_18_), .B(AES_CORE_DATAPATH__abc_16259_n3579), .Y(AES_CORE_DATAPATH__abc_16259_n3582) );
  AND2X2 AND2X2_631 ( .A(AES_CORE_DATAPATH_last_round_pp2_bF_buf0), .B(AES_CORE_DATAPATH_MIX_COL_col_2__2_), .Y(AES_CORE_DATAPATH__abc_16259_n3585) );
  AND2X2 AND2X2_632 ( .A(AES_CORE_DATAPATH__abc_16259_n2798_bF_buf1), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_18_), .Y(AES_CORE_DATAPATH__abc_16259_n3586) );
  AND2X2 AND2X2_633 ( .A(AES_CORE_DATAPATH__abc_16259_n3584_1), .B(AES_CORE_DATAPATH__abc_16259_n3588), .Y(AES_CORE_DATAPATH__abc_16259_n3589_1) );
  AND2X2 AND2X2_634 ( .A(AES_CORE_DATAPATH__abc_16259_n3589_1), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n3590) );
  AND2X2 AND2X2_635 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf6), .B(AES_CORE_DATAPATH_col_3__18_), .Y(AES_CORE_DATAPATH__abc_16259_n3591_1) );
  AND2X2 AND2X2_636 ( .A(AES_CORE_DATAPATH__abc_16259_n3594), .B(AES_CORE_DATAPATH__abc_16259_n3596), .Y(AES_CORE_DATAPATH__abc_16259_n3597) );
  AND2X2 AND2X2_637 ( .A(AES_CORE_DATAPATH__abc_16259_n2782_bF_buf0), .B(AES_CORE_DATAPATH_col_3__19_), .Y(AES_CORE_DATAPATH__abc_16259_n3598) );
  AND2X2 AND2X2_638 ( .A(AES_CORE_DATAPATH__abc_16259_n2786_bF_buf0), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_83_), .Y(AES_CORE_DATAPATH__abc_16259_n3599) );
  AND2X2 AND2X2_639 ( .A(AES_CORE_DATAPATH__abc_16259_n2789_bF_buf0), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_51_), .Y(AES_CORE_DATAPATH__abc_16259_n3600) );
  AND2X2 AND2X2_64 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n173), .B(AES_CORE_CONTROL_UNIT_rd_count_2_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n178) );
  AND2X2 AND2X2_640 ( .A(AES_CORE_DATAPATH__abc_16259_n3603), .B(AES_CORE_DATAPATH__abc_16259_n3597), .Y(AES_CORE_DATAPATH__abc_16259_n3604) );
  AND2X2 AND2X2_641 ( .A(AES_CORE_DATAPATH__abc_16259_n2837_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__19_), .Y(AES_CORE_DATAPATH__abc_16259_n3606) );
  AND2X2 AND2X2_642 ( .A(AES_CORE_DATAPATH__abc_16259_n2887_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__19_), .Y(AES_CORE_DATAPATH__abc_16259_n3608) );
  AND2X2 AND2X2_643 ( .A(AES_CORE_DATAPATH__abc_16259_n2830_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__19_), .Y(AES_CORE_DATAPATH__abc_16259_n3609) );
  AND2X2 AND2X2_644 ( .A(AES_CORE_DATAPATH__abc_16259_n3611), .B(AES_CORE_DATAPATH__abc_16259_n3612_1), .Y(_auto_iopadmap_cc_313_execute_26949_19_) );
  AND2X2 AND2X2_645 ( .A(AES_CORE_DATAPATH__abc_16259_n2855_bF_buf0), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_19_), .Y(AES_CORE_DATAPATH__abc_16259_n3615) );
  AND2X2 AND2X2_646 ( .A(AES_CORE_DATAPATH__abc_16259_n2857_bF_buf0), .B(AES_CORE_DATAPATH_MIX_COL_col_2__3_), .Y(AES_CORE_DATAPATH__abc_16259_n3616_1) );
  AND2X2 AND2X2_647 ( .A(AES_CORE_DATAPATH__abc_16259_n3614), .B(AES_CORE_DATAPATH__abc_16259_n3618_1), .Y(AES_CORE_DATAPATH__abc_16259_n3619) );
  AND2X2 AND2X2_648 ( .A(_auto_iopadmap_cc_313_execute_26949_19_), .B(AES_CORE_DATAPATH__abc_16259_n3619), .Y(AES_CORE_DATAPATH__abc_16259_n3622_1) );
  AND2X2 AND2X2_649 ( .A(AES_CORE_DATAPATH_last_round_pp2_bF_buf4), .B(AES_CORE_DATAPATH_MIX_COL_col_2__3_), .Y(AES_CORE_DATAPATH__abc_16259_n3625) );
  AND2X2 AND2X2_65 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n166), .B(AES_CORE_CONTROL_UNIT__abc_15841_n180), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n181_1) );
  AND2X2 AND2X2_650 ( .A(AES_CORE_DATAPATH__abc_16259_n2798_bF_buf0), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_19_), .Y(AES_CORE_DATAPATH__abc_16259_n3626) );
  AND2X2 AND2X2_651 ( .A(AES_CORE_DATAPATH__abc_16259_n3624), .B(AES_CORE_DATAPATH__abc_16259_n3628), .Y(AES_CORE_DATAPATH__abc_16259_n3629) );
  AND2X2 AND2X2_652 ( .A(AES_CORE_DATAPATH__abc_16259_n3629), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n3630) );
  AND2X2 AND2X2_653 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf5), .B(AES_CORE_DATAPATH_col_3__19_), .Y(AES_CORE_DATAPATH__abc_16259_n3631) );
  AND2X2 AND2X2_654 ( .A(AES_CORE_DATAPATH__abc_16259_n3634_1), .B(AES_CORE_DATAPATH__abc_16259_n3636_1), .Y(AES_CORE_DATAPATH__abc_16259_n3637) );
  AND2X2 AND2X2_655 ( .A(AES_CORE_DATAPATH__abc_16259_n2782_bF_buf4), .B(AES_CORE_DATAPATH_col_3__20_), .Y(AES_CORE_DATAPATH__abc_16259_n3638) );
  AND2X2 AND2X2_656 ( .A(AES_CORE_DATAPATH__abc_16259_n2786_bF_buf4), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_84_), .Y(AES_CORE_DATAPATH__abc_16259_n3639) );
  AND2X2 AND2X2_657 ( .A(AES_CORE_DATAPATH__abc_16259_n2789_bF_buf4), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_52_), .Y(AES_CORE_DATAPATH__abc_16259_n3640) );
  AND2X2 AND2X2_658 ( .A(AES_CORE_DATAPATH__abc_16259_n3643), .B(AES_CORE_DATAPATH__abc_16259_n3637), .Y(AES_CORE_DATAPATH__abc_16259_n3644) );
  AND2X2 AND2X2_659 ( .A(AES_CORE_DATAPATH__abc_16259_n2837_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__20_), .Y(AES_CORE_DATAPATH__abc_16259_n3646) );
  AND2X2 AND2X2_66 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n181_1), .B(AES_CORE_CONTROL_UNIT__abc_15841_n179_1), .Y(AES_CORE_CONTROL_UNIT_rd_count_2__FF_INPUT) );
  AND2X2 AND2X2_660 ( .A(AES_CORE_DATAPATH__abc_16259_n2887_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__20_), .Y(AES_CORE_DATAPATH__abc_16259_n3648) );
  AND2X2 AND2X2_661 ( .A(AES_CORE_DATAPATH__abc_16259_n2830_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__20_), .Y(AES_CORE_DATAPATH__abc_16259_n3649_1) );
  AND2X2 AND2X2_662 ( .A(AES_CORE_DATAPATH__abc_16259_n3651_1), .B(AES_CORE_DATAPATH__abc_16259_n3652), .Y(_auto_iopadmap_cc_313_execute_26949_20_) );
  AND2X2 AND2X2_663 ( .A(AES_CORE_DATAPATH__abc_16259_n2855_bF_buf4), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_20_), .Y(AES_CORE_DATAPATH__abc_16259_n3655) );
  AND2X2 AND2X2_664 ( .A(AES_CORE_DATAPATH__abc_16259_n2857_bF_buf4), .B(AES_CORE_DATAPATH_MIX_COL_col_2__4_), .Y(AES_CORE_DATAPATH__abc_16259_n3656) );
  AND2X2 AND2X2_665 ( .A(AES_CORE_DATAPATH__abc_16259_n3654), .B(AES_CORE_DATAPATH__abc_16259_n3658), .Y(AES_CORE_DATAPATH__abc_16259_n3659) );
  AND2X2 AND2X2_666 ( .A(_auto_iopadmap_cc_313_execute_26949_20_), .B(AES_CORE_DATAPATH__abc_16259_n3659), .Y(AES_CORE_DATAPATH__abc_16259_n3662) );
  AND2X2 AND2X2_667 ( .A(AES_CORE_DATAPATH_last_round_pp2_bF_buf3), .B(AES_CORE_DATAPATH_MIX_COL_col_2__4_), .Y(AES_CORE_DATAPATH__abc_16259_n3665_1) );
  AND2X2 AND2X2_668 ( .A(AES_CORE_DATAPATH__abc_16259_n2798_bF_buf4), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_20_), .Y(AES_CORE_DATAPATH__abc_16259_n3666) );
  AND2X2 AND2X2_669 ( .A(AES_CORE_DATAPATH__abc_16259_n3664), .B(AES_CORE_DATAPATH__abc_16259_n3668), .Y(AES_CORE_DATAPATH__abc_16259_n3669) );
  AND2X2 AND2X2_67 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n178), .B(AES_CORE_CONTROL_UNIT_rd_count_3_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n183_1) );
  AND2X2 AND2X2_670 ( .A(AES_CORE_DATAPATH__abc_16259_n3669), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf14), .Y(AES_CORE_DATAPATH__abc_16259_n3670_1) );
  AND2X2 AND2X2_671 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf4), .B(AES_CORE_DATAPATH_col_3__20_), .Y(AES_CORE_DATAPATH__abc_16259_n3671_1) );
  AND2X2 AND2X2_672 ( .A(AES_CORE_DATAPATH__abc_16259_n3674), .B(AES_CORE_DATAPATH__abc_16259_n3676), .Y(AES_CORE_DATAPATH__abc_16259_n3677) );
  AND2X2 AND2X2_673 ( .A(AES_CORE_DATAPATH__abc_16259_n2782_bF_buf3), .B(AES_CORE_DATAPATH_col_3__21_), .Y(AES_CORE_DATAPATH__abc_16259_n3678_1) );
  AND2X2 AND2X2_674 ( .A(AES_CORE_DATAPATH__abc_16259_n2786_bF_buf3), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_85_), .Y(AES_CORE_DATAPATH__abc_16259_n3679_1) );
  AND2X2 AND2X2_675 ( .A(AES_CORE_DATAPATH__abc_16259_n2789_bF_buf3), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_53_), .Y(AES_CORE_DATAPATH__abc_16259_n3680) );
  AND2X2 AND2X2_676 ( .A(AES_CORE_DATAPATH__abc_16259_n3683), .B(AES_CORE_DATAPATH__abc_16259_n3677), .Y(AES_CORE_DATAPATH__abc_16259_n3684) );
  AND2X2 AND2X2_677 ( .A(AES_CORE_DATAPATH__abc_16259_n2837_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__21_), .Y(AES_CORE_DATAPATH__abc_16259_n3686_1) );
  AND2X2 AND2X2_678 ( .A(AES_CORE_DATAPATH__abc_16259_n2887_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__21_), .Y(AES_CORE_DATAPATH__abc_16259_n3688) );
  AND2X2 AND2X2_679 ( .A(AES_CORE_DATAPATH__abc_16259_n2830_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__21_), .Y(AES_CORE_DATAPATH__abc_16259_n3689_1) );
  AND2X2 AND2X2_68 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n185), .B(AES_CORE_CONTROL_UNIT__abc_15841_n166), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n186) );
  AND2X2 AND2X2_680 ( .A(AES_CORE_DATAPATH__abc_16259_n3691), .B(AES_CORE_DATAPATH__abc_16259_n3692), .Y(_auto_iopadmap_cc_313_execute_26949_21_) );
  AND2X2 AND2X2_681 ( .A(AES_CORE_DATAPATH__abc_16259_n2855_bF_buf3), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_21_), .Y(AES_CORE_DATAPATH__abc_16259_n3695_1) );
  AND2X2 AND2X2_682 ( .A(AES_CORE_DATAPATH__abc_16259_n2857_bF_buf3), .B(AES_CORE_DATAPATH_MIX_COL_col_2__5_), .Y(AES_CORE_DATAPATH__abc_16259_n3696) );
  AND2X2 AND2X2_683 ( .A(AES_CORE_DATAPATH__abc_16259_n3694_1), .B(AES_CORE_DATAPATH__abc_16259_n3698), .Y(AES_CORE_DATAPATH__abc_16259_n3699) );
  AND2X2 AND2X2_684 ( .A(_auto_iopadmap_cc_313_execute_26949_21_), .B(AES_CORE_DATAPATH__abc_16259_n3699), .Y(AES_CORE_DATAPATH__abc_16259_n3702_1) );
  AND2X2 AND2X2_685 ( .A(AES_CORE_DATAPATH_last_round_pp2_bF_buf2), .B(AES_CORE_DATAPATH_MIX_COL_col_2__5_), .Y(AES_CORE_DATAPATH__abc_16259_n3705_1) );
  AND2X2 AND2X2_686 ( .A(AES_CORE_DATAPATH__abc_16259_n2798_bF_buf3), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_21_), .Y(AES_CORE_DATAPATH__abc_16259_n3706) );
  AND2X2 AND2X2_687 ( .A(AES_CORE_DATAPATH__abc_16259_n3704), .B(AES_CORE_DATAPATH__abc_16259_n3708), .Y(AES_CORE_DATAPATH__abc_16259_n3709) );
  AND2X2 AND2X2_688 ( .A(AES_CORE_DATAPATH__abc_16259_n3709), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf13), .Y(AES_CORE_DATAPATH__abc_16259_n3710_1) );
  AND2X2 AND2X2_689 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf3), .B(AES_CORE_DATAPATH_col_3__21_), .Y(AES_CORE_DATAPATH__abc_16259_n3711_1) );
  AND2X2 AND2X2_69 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n186), .B(AES_CORE_CONTROL_UNIT__abc_15841_n184_1), .Y(AES_CORE_CONTROL_UNIT_rd_count_3__FF_INPUT) );
  AND2X2 AND2X2_690 ( .A(AES_CORE_DATAPATH__abc_16259_n3714), .B(AES_CORE_DATAPATH__abc_16259_n3716), .Y(AES_CORE_DATAPATH__abc_16259_n3717) );
  AND2X2 AND2X2_691 ( .A(AES_CORE_DATAPATH__abc_16259_n2782_bF_buf2), .B(AES_CORE_DATAPATH_col_3__22_), .Y(AES_CORE_DATAPATH__abc_16259_n3718_1) );
  AND2X2 AND2X2_692 ( .A(AES_CORE_DATAPATH__abc_16259_n2786_bF_buf2), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_86_), .Y(AES_CORE_DATAPATH__abc_16259_n3719_1) );
  AND2X2 AND2X2_693 ( .A(AES_CORE_DATAPATH__abc_16259_n2789_bF_buf2), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_54_), .Y(AES_CORE_DATAPATH__abc_16259_n3720) );
  AND2X2 AND2X2_694 ( .A(AES_CORE_DATAPATH__abc_16259_n3723), .B(AES_CORE_DATAPATH__abc_16259_n3717), .Y(AES_CORE_DATAPATH__abc_16259_n3724) );
  AND2X2 AND2X2_695 ( .A(AES_CORE_DATAPATH__abc_16259_n2837_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__22_), .Y(AES_CORE_DATAPATH__abc_16259_n3726_1) );
  AND2X2 AND2X2_696 ( .A(AES_CORE_DATAPATH__abc_16259_n2887_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__22_), .Y(AES_CORE_DATAPATH__abc_16259_n3728) );
  AND2X2 AND2X2_697 ( .A(AES_CORE_DATAPATH__abc_16259_n2830_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__22_), .Y(AES_CORE_DATAPATH__abc_16259_n3729_1) );
  AND2X2 AND2X2_698 ( .A(AES_CORE_DATAPATH__abc_16259_n3731), .B(AES_CORE_DATAPATH__abc_16259_n3732), .Y(_auto_iopadmap_cc_313_execute_26949_22_) );
  AND2X2 AND2X2_699 ( .A(AES_CORE_DATAPATH__abc_16259_n2855_bF_buf2), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_22_), .Y(AES_CORE_DATAPATH__abc_16259_n3735_1) );
  AND2X2 AND2X2_7 ( .A(\addr[0] ), .B(read_en), .Y(AES_CORE_DATAPATH_col_sel_host_0_) );
  AND2X2 AND2X2_70 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n190), .B(AES_CORE_CONTROL_UNIT_last_round_bF_buf2), .Y(AES_CORE_CONTROL_UNIT_rk_sel_0_) );
  AND2X2 AND2X2_700 ( .A(AES_CORE_DATAPATH__abc_16259_n2857_bF_buf2), .B(AES_CORE_DATAPATH_MIX_COL_col_2__6_), .Y(AES_CORE_DATAPATH__abc_16259_n3736) );
  AND2X2 AND2X2_701 ( .A(AES_CORE_DATAPATH__abc_16259_n3734_1), .B(AES_CORE_DATAPATH__abc_16259_n3738), .Y(AES_CORE_DATAPATH__abc_16259_n3739) );
  AND2X2 AND2X2_702 ( .A(_auto_iopadmap_cc_313_execute_26949_22_), .B(AES_CORE_DATAPATH__abc_16259_n3739), .Y(AES_CORE_DATAPATH__abc_16259_n3742_1) );
  AND2X2 AND2X2_703 ( .A(AES_CORE_DATAPATH_last_round_pp2_bF_buf1), .B(AES_CORE_DATAPATH_MIX_COL_col_2__6_), .Y(AES_CORE_DATAPATH__abc_16259_n3745_1) );
  AND2X2 AND2X2_704 ( .A(AES_CORE_DATAPATH__abc_16259_n2798_bF_buf2), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_22_), .Y(AES_CORE_DATAPATH__abc_16259_n3746) );
  AND2X2 AND2X2_705 ( .A(AES_CORE_DATAPATH__abc_16259_n3744), .B(AES_CORE_DATAPATH__abc_16259_n3748), .Y(AES_CORE_DATAPATH__abc_16259_n3749) );
  AND2X2 AND2X2_706 ( .A(AES_CORE_DATAPATH__abc_16259_n3749), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf12), .Y(AES_CORE_DATAPATH__abc_16259_n3750_1) );
  AND2X2 AND2X2_707 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf2), .B(AES_CORE_DATAPATH_col_3__22_), .Y(AES_CORE_DATAPATH__abc_16259_n3751_1) );
  AND2X2 AND2X2_708 ( .A(AES_CORE_DATAPATH__abc_16259_n3754), .B(AES_CORE_DATAPATH__abc_16259_n3756), .Y(AES_CORE_DATAPATH__abc_16259_n3757) );
  AND2X2 AND2X2_709 ( .A(AES_CORE_DATAPATH__abc_16259_n2782_bF_buf1), .B(AES_CORE_DATAPATH_col_3__23_), .Y(AES_CORE_DATAPATH__abc_16259_n3758_1) );
  AND2X2 AND2X2_71 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n142), .B(AES_CORE_CONTROL_UNIT__abc_15841_n190), .Y(AES_CORE_CONTROL_UNIT_rk_sel_1_) );
  AND2X2 AND2X2_710 ( .A(AES_CORE_DATAPATH__abc_16259_n2786_bF_buf1), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_87_), .Y(AES_CORE_DATAPATH__abc_16259_n3759_1) );
  AND2X2 AND2X2_711 ( .A(AES_CORE_DATAPATH__abc_16259_n2789_bF_buf1), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_55_), .Y(AES_CORE_DATAPATH__abc_16259_n3760) );
  AND2X2 AND2X2_712 ( .A(AES_CORE_DATAPATH__abc_16259_n3763), .B(AES_CORE_DATAPATH__abc_16259_n3757), .Y(AES_CORE_DATAPATH__abc_16259_n3764) );
  AND2X2 AND2X2_713 ( .A(AES_CORE_DATAPATH__abc_16259_n2837_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__23_), .Y(AES_CORE_DATAPATH__abc_16259_n3766_1) );
  AND2X2 AND2X2_714 ( .A(AES_CORE_DATAPATH__abc_16259_n2887_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__23_), .Y(AES_CORE_DATAPATH__abc_16259_n3768) );
  AND2X2 AND2X2_715 ( .A(AES_CORE_DATAPATH__abc_16259_n2830_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__23_), .Y(AES_CORE_DATAPATH__abc_16259_n3769_1) );
  AND2X2 AND2X2_716 ( .A(AES_CORE_DATAPATH__abc_16259_n3771), .B(AES_CORE_DATAPATH__abc_16259_n3772), .Y(_auto_iopadmap_cc_313_execute_26949_23_) );
  AND2X2 AND2X2_717 ( .A(AES_CORE_DATAPATH__abc_16259_n2855_bF_buf1), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_23_), .Y(AES_CORE_DATAPATH__abc_16259_n3775_1) );
  AND2X2 AND2X2_718 ( .A(AES_CORE_DATAPATH__abc_16259_n2857_bF_buf1), .B(AES_CORE_DATAPATH_MIX_COL_col_2__7_), .Y(AES_CORE_DATAPATH__abc_16259_n3776) );
  AND2X2 AND2X2_719 ( .A(AES_CORE_DATAPATH__abc_16259_n3774_1), .B(AES_CORE_DATAPATH__abc_16259_n3778), .Y(AES_CORE_DATAPATH__abc_16259_n3779) );
  AND2X2 AND2X2_72 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf10), .B(AES_CORE_CONTROL_UNIT__abc_15841_n144), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n193) );
  AND2X2 AND2X2_720 ( .A(_auto_iopadmap_cc_313_execute_26949_23_), .B(AES_CORE_DATAPATH__abc_16259_n3779), .Y(AES_CORE_DATAPATH__abc_16259_n3782_1) );
  AND2X2 AND2X2_721 ( .A(AES_CORE_DATAPATH_last_round_pp2_bF_buf0), .B(AES_CORE_DATAPATH_MIX_COL_col_2__7_), .Y(AES_CORE_DATAPATH__abc_16259_n3785_1) );
  AND2X2 AND2X2_722 ( .A(AES_CORE_DATAPATH__abc_16259_n2798_bF_buf1), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_23_), .Y(AES_CORE_DATAPATH__abc_16259_n3786) );
  AND2X2 AND2X2_723 ( .A(AES_CORE_DATAPATH__abc_16259_n3784), .B(AES_CORE_DATAPATH__abc_16259_n3788), .Y(AES_CORE_DATAPATH__abc_16259_n3789) );
  AND2X2 AND2X2_724 ( .A(AES_CORE_DATAPATH__abc_16259_n3789), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf11), .Y(AES_CORE_DATAPATH__abc_16259_n3790_1) );
  AND2X2 AND2X2_725 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf1), .B(AES_CORE_DATAPATH_col_3__23_), .Y(AES_CORE_DATAPATH__abc_16259_n3791_1) );
  AND2X2 AND2X2_726 ( .A(AES_CORE_DATAPATH__abc_16259_n3794), .B(AES_CORE_DATAPATH__abc_16259_n3796), .Y(AES_CORE_DATAPATH__abc_16259_n3797) );
  AND2X2 AND2X2_727 ( .A(AES_CORE_DATAPATH__abc_16259_n2782_bF_buf0), .B(AES_CORE_DATAPATH_col_3__24_), .Y(AES_CORE_DATAPATH__abc_16259_n3798_1) );
  AND2X2 AND2X2_728 ( .A(AES_CORE_DATAPATH__abc_16259_n2786_bF_buf0), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_88_), .Y(AES_CORE_DATAPATH__abc_16259_n3799_1) );
  AND2X2 AND2X2_729 ( .A(AES_CORE_DATAPATH__abc_16259_n2789_bF_buf0), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_56_), .Y(AES_CORE_DATAPATH__abc_16259_n3800) );
  AND2X2 AND2X2_73 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n196), .B(AES_CORE_CONTROL_UNIT_state_6_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n197_1) );
  AND2X2 AND2X2_730 ( .A(AES_CORE_DATAPATH__abc_16259_n3803), .B(AES_CORE_DATAPATH__abc_16259_n3797), .Y(AES_CORE_DATAPATH__abc_16259_n3804) );
  AND2X2 AND2X2_731 ( .A(AES_CORE_DATAPATH__abc_16259_n2837_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__24_), .Y(AES_CORE_DATAPATH__abc_16259_n3806_1) );
  AND2X2 AND2X2_732 ( .A(AES_CORE_DATAPATH__abc_16259_n2887_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__24_), .Y(AES_CORE_DATAPATH__abc_16259_n3808) );
  AND2X2 AND2X2_733 ( .A(AES_CORE_DATAPATH__abc_16259_n2830_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__24_), .Y(AES_CORE_DATAPATH__abc_16259_n3809_1) );
  AND2X2 AND2X2_734 ( .A(AES_CORE_DATAPATH__abc_16259_n3811), .B(AES_CORE_DATAPATH__abc_16259_n3812), .Y(_auto_iopadmap_cc_313_execute_26949_24_) );
  AND2X2 AND2X2_735 ( .A(AES_CORE_DATAPATH__abc_16259_n2855_bF_buf0), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_24_), .Y(AES_CORE_DATAPATH__abc_16259_n3815_1) );
  AND2X2 AND2X2_736 ( .A(AES_CORE_DATAPATH__abc_16259_n2857_bF_buf0), .B(AES_CORE_DATAPATH_MIX_COL_col_3__0_), .Y(AES_CORE_DATAPATH__abc_16259_n3816) );
  AND2X2 AND2X2_737 ( .A(AES_CORE_DATAPATH__abc_16259_n3814_1), .B(AES_CORE_DATAPATH__abc_16259_n3818), .Y(AES_CORE_DATAPATH__abc_16259_n3819) );
  AND2X2 AND2X2_738 ( .A(_auto_iopadmap_cc_313_execute_26949_24_), .B(AES_CORE_DATAPATH__abc_16259_n3819), .Y(AES_CORE_DATAPATH__abc_16259_n3822_1) );
  AND2X2 AND2X2_739 ( .A(AES_CORE_DATAPATH_last_round_pp2_bF_buf4), .B(AES_CORE_DATAPATH_MIX_COL_col_3__0_), .Y(AES_CORE_DATAPATH__abc_16259_n3825_1) );
  AND2X2 AND2X2_74 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n106_1), .B(AES_CORE_CONTROL_UNIT_state_8_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n199) );
  AND2X2 AND2X2_740 ( .A(AES_CORE_DATAPATH__abc_16259_n2798_bF_buf0), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_24_), .Y(AES_CORE_DATAPATH__abc_16259_n3826) );
  AND2X2 AND2X2_741 ( .A(AES_CORE_DATAPATH__abc_16259_n3824), .B(AES_CORE_DATAPATH__abc_16259_n3828), .Y(AES_CORE_DATAPATH__abc_16259_n3829) );
  AND2X2 AND2X2_742 ( .A(AES_CORE_DATAPATH__abc_16259_n3829), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf10), .Y(AES_CORE_DATAPATH__abc_16259_n3830_1) );
  AND2X2 AND2X2_743 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf0), .B(AES_CORE_DATAPATH_col_3__24_), .Y(AES_CORE_DATAPATH__abc_16259_n3831_1) );
  AND2X2 AND2X2_744 ( .A(AES_CORE_DATAPATH__abc_16259_n3834), .B(AES_CORE_DATAPATH__abc_16259_n3836), .Y(AES_CORE_DATAPATH__abc_16259_n3837) );
  AND2X2 AND2X2_745 ( .A(AES_CORE_DATAPATH__abc_16259_n2782_bF_buf4), .B(AES_CORE_DATAPATH_col_3__25_), .Y(AES_CORE_DATAPATH__abc_16259_n3838_1) );
  AND2X2 AND2X2_746 ( .A(AES_CORE_DATAPATH__abc_16259_n2786_bF_buf4), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_89_), .Y(AES_CORE_DATAPATH__abc_16259_n3839_1) );
  AND2X2 AND2X2_747 ( .A(AES_CORE_DATAPATH__abc_16259_n2789_bF_buf4), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_57_), .Y(AES_CORE_DATAPATH__abc_16259_n3840) );
  AND2X2 AND2X2_748 ( .A(AES_CORE_DATAPATH__abc_16259_n3843), .B(AES_CORE_DATAPATH__abc_16259_n3837), .Y(AES_CORE_DATAPATH__abc_16259_n3844) );
  AND2X2 AND2X2_749 ( .A(AES_CORE_DATAPATH__abc_16259_n2837_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__25_), .Y(AES_CORE_DATAPATH__abc_16259_n3846_1) );
  AND2X2 AND2X2_75 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf8), .B(AES_CORE_CONTROL_UNIT_state_8_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n209_1) );
  AND2X2 AND2X2_750 ( .A(AES_CORE_DATAPATH__abc_16259_n2887_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__25_), .Y(AES_CORE_DATAPATH__abc_16259_n3848) );
  AND2X2 AND2X2_751 ( .A(AES_CORE_DATAPATH__abc_16259_n2830_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__25_), .Y(AES_CORE_DATAPATH__abc_16259_n3849_1) );
  AND2X2 AND2X2_752 ( .A(AES_CORE_DATAPATH__abc_16259_n3851), .B(AES_CORE_DATAPATH__abc_16259_n3852), .Y(_auto_iopadmap_cc_313_execute_26949_25_) );
  AND2X2 AND2X2_753 ( .A(AES_CORE_DATAPATH__abc_16259_n2855_bF_buf4), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_25_), .Y(AES_CORE_DATAPATH__abc_16259_n3855_1) );
  AND2X2 AND2X2_754 ( .A(AES_CORE_DATAPATH__abc_16259_n2857_bF_buf4), .B(AES_CORE_DATAPATH_MIX_COL_col_3__1_), .Y(AES_CORE_DATAPATH__abc_16259_n3856) );
  AND2X2 AND2X2_755 ( .A(AES_CORE_DATAPATH__abc_16259_n3854_1), .B(AES_CORE_DATAPATH__abc_16259_n3858), .Y(AES_CORE_DATAPATH__abc_16259_n3859) );
  AND2X2 AND2X2_756 ( .A(_auto_iopadmap_cc_313_execute_26949_25_), .B(AES_CORE_DATAPATH__abc_16259_n3859), .Y(AES_CORE_DATAPATH__abc_16259_n3862_1) );
  AND2X2 AND2X2_757 ( .A(AES_CORE_DATAPATH_last_round_pp2_bF_buf3), .B(AES_CORE_DATAPATH_MIX_COL_col_3__1_), .Y(AES_CORE_DATAPATH__abc_16259_n3865_1) );
  AND2X2 AND2X2_758 ( .A(AES_CORE_DATAPATH__abc_16259_n2798_bF_buf4), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_25_), .Y(AES_CORE_DATAPATH__abc_16259_n3866) );
  AND2X2 AND2X2_759 ( .A(AES_CORE_DATAPATH__abc_16259_n3864), .B(AES_CORE_DATAPATH__abc_16259_n3868), .Y(AES_CORE_DATAPATH__abc_16259_n3869) );
  AND2X2 AND2X2_76 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n106_1), .B(AES_CORE_CONTROL_UNIT_state_2_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n210_1) );
  AND2X2 AND2X2_760 ( .A(AES_CORE_DATAPATH__abc_16259_n3869), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf9), .Y(AES_CORE_DATAPATH__abc_16259_n3870_1) );
  AND2X2 AND2X2_761 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf12), .B(AES_CORE_DATAPATH_col_3__25_), .Y(AES_CORE_DATAPATH__abc_16259_n3871_1) );
  AND2X2 AND2X2_762 ( .A(AES_CORE_DATAPATH__abc_16259_n3874), .B(AES_CORE_DATAPATH__abc_16259_n3876), .Y(AES_CORE_DATAPATH__abc_16259_n3877) );
  AND2X2 AND2X2_763 ( .A(AES_CORE_DATAPATH__abc_16259_n2782_bF_buf3), .B(AES_CORE_DATAPATH_col_3__26_), .Y(AES_CORE_DATAPATH__abc_16259_n3878_1) );
  AND2X2 AND2X2_764 ( .A(AES_CORE_DATAPATH__abc_16259_n2786_bF_buf3), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_90_), .Y(AES_CORE_DATAPATH__abc_16259_n3879_1) );
  AND2X2 AND2X2_765 ( .A(AES_CORE_DATAPATH__abc_16259_n2789_bF_buf3), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_58_), .Y(AES_CORE_DATAPATH__abc_16259_n3880) );
  AND2X2 AND2X2_766 ( .A(AES_CORE_DATAPATH__abc_16259_n3883), .B(AES_CORE_DATAPATH__abc_16259_n3877), .Y(AES_CORE_DATAPATH__abc_16259_n3884) );
  AND2X2 AND2X2_767 ( .A(AES_CORE_DATAPATH__abc_16259_n2837_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__26_), .Y(AES_CORE_DATAPATH__abc_16259_n3886_1) );
  AND2X2 AND2X2_768 ( .A(AES_CORE_DATAPATH__abc_16259_n2887_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__26_), .Y(AES_CORE_DATAPATH__abc_16259_n3888) );
  AND2X2 AND2X2_769 ( .A(AES_CORE_DATAPATH__abc_16259_n2830_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__26_), .Y(AES_CORE_DATAPATH__abc_16259_n3889_1) );
  AND2X2 AND2X2_77 ( .A(AES_CORE_CONTROL_UNIT_last_round_bF_buf0), .B(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf4), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n213) );
  AND2X2 AND2X2_770 ( .A(AES_CORE_DATAPATH__abc_16259_n3891), .B(AES_CORE_DATAPATH__abc_16259_n3892), .Y(_auto_iopadmap_cc_313_execute_26949_26_) );
  AND2X2 AND2X2_771 ( .A(AES_CORE_DATAPATH__abc_16259_n2855_bF_buf3), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_26_), .Y(AES_CORE_DATAPATH__abc_16259_n3895_1) );
  AND2X2 AND2X2_772 ( .A(AES_CORE_DATAPATH__abc_16259_n2857_bF_buf3), .B(AES_CORE_DATAPATH_MIX_COL_col_3__2_), .Y(AES_CORE_DATAPATH__abc_16259_n3896) );
  AND2X2 AND2X2_773 ( .A(AES_CORE_DATAPATH__abc_16259_n3894_1), .B(AES_CORE_DATAPATH__abc_16259_n3898), .Y(AES_CORE_DATAPATH__abc_16259_n3899) );
  AND2X2 AND2X2_774 ( .A(_auto_iopadmap_cc_313_execute_26949_26_), .B(AES_CORE_DATAPATH__abc_16259_n3899), .Y(AES_CORE_DATAPATH__abc_16259_n3902_1) );
  AND2X2 AND2X2_775 ( .A(AES_CORE_DATAPATH_last_round_pp2_bF_buf2), .B(AES_CORE_DATAPATH_MIX_COL_col_3__2_), .Y(AES_CORE_DATAPATH__abc_16259_n3905_1) );
  AND2X2 AND2X2_776 ( .A(AES_CORE_DATAPATH__abc_16259_n2798_bF_buf3), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_26_), .Y(AES_CORE_DATAPATH__abc_16259_n3906) );
  AND2X2 AND2X2_777 ( .A(AES_CORE_DATAPATH__abc_16259_n3904), .B(AES_CORE_DATAPATH__abc_16259_n3908), .Y(AES_CORE_DATAPATH__abc_16259_n3909) );
  AND2X2 AND2X2_778 ( .A(AES_CORE_DATAPATH__abc_16259_n3909), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf8), .Y(AES_CORE_DATAPATH__abc_16259_n3910_1) );
  AND2X2 AND2X2_779 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf11), .B(AES_CORE_DATAPATH_col_3__26_), .Y(AES_CORE_DATAPATH__abc_16259_n3911_1) );
  AND2X2 AND2X2_78 ( .A(AES_CORE_CONTROL_UNIT_last_round_bF_buf5), .B(AES_CORE_CONTROL_UNIT_mode_cbc_bF_buf4), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n214) );
  AND2X2 AND2X2_780 ( .A(AES_CORE_DATAPATH__abc_16259_n3914), .B(AES_CORE_DATAPATH__abc_16259_n3916), .Y(AES_CORE_DATAPATH__abc_16259_n3917) );
  AND2X2 AND2X2_781 ( .A(AES_CORE_DATAPATH__abc_16259_n2782_bF_buf2), .B(AES_CORE_DATAPATH_col_3__27_), .Y(AES_CORE_DATAPATH__abc_16259_n3918_1) );
  AND2X2 AND2X2_782 ( .A(AES_CORE_DATAPATH__abc_16259_n2786_bF_buf2), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_91_), .Y(AES_CORE_DATAPATH__abc_16259_n3919_1) );
  AND2X2 AND2X2_783 ( .A(AES_CORE_DATAPATH__abc_16259_n2789_bF_buf2), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_59_), .Y(AES_CORE_DATAPATH__abc_16259_n3920) );
  AND2X2 AND2X2_784 ( .A(AES_CORE_DATAPATH__abc_16259_n3923), .B(AES_CORE_DATAPATH__abc_16259_n3917), .Y(AES_CORE_DATAPATH__abc_16259_n3924) );
  AND2X2 AND2X2_785 ( .A(AES_CORE_DATAPATH__abc_16259_n2837_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__27_), .Y(AES_CORE_DATAPATH__abc_16259_n3926_1) );
  AND2X2 AND2X2_786 ( .A(AES_CORE_DATAPATH__abc_16259_n2887_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__27_), .Y(AES_CORE_DATAPATH__abc_16259_n3928) );
  AND2X2 AND2X2_787 ( .A(AES_CORE_DATAPATH__abc_16259_n2830_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__27_), .Y(AES_CORE_DATAPATH__abc_16259_n3929_1) );
  AND2X2 AND2X2_788 ( .A(AES_CORE_DATAPATH__abc_16259_n3931), .B(AES_CORE_DATAPATH__abc_16259_n3932), .Y(_auto_iopadmap_cc_313_execute_26949_27_) );
  AND2X2 AND2X2_789 ( .A(AES_CORE_DATAPATH__abc_16259_n2855_bF_buf2), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_27_), .Y(AES_CORE_DATAPATH__abc_16259_n3935_1) );
  AND2X2 AND2X2_79 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n106_1), .B(AES_CORE_CONTROL_UNIT__abc_15841_n214), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n215) );
  AND2X2 AND2X2_790 ( .A(AES_CORE_DATAPATH__abc_16259_n2857_bF_buf2), .B(AES_CORE_DATAPATH_MIX_COL_col_3__3_), .Y(AES_CORE_DATAPATH__abc_16259_n3936) );
  AND2X2 AND2X2_791 ( .A(AES_CORE_DATAPATH__abc_16259_n3934_1), .B(AES_CORE_DATAPATH__abc_16259_n3938), .Y(AES_CORE_DATAPATH__abc_16259_n3939) );
  AND2X2 AND2X2_792 ( .A(_auto_iopadmap_cc_313_execute_26949_27_), .B(AES_CORE_DATAPATH__abc_16259_n3939), .Y(AES_CORE_DATAPATH__abc_16259_n3942_1) );
  AND2X2 AND2X2_793 ( .A(AES_CORE_DATAPATH_last_round_pp2_bF_buf1), .B(AES_CORE_DATAPATH_MIX_COL_col_3__3_), .Y(AES_CORE_DATAPATH__abc_16259_n3945_1) );
  AND2X2 AND2X2_794 ( .A(AES_CORE_DATAPATH__abc_16259_n2798_bF_buf2), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_27_), .Y(AES_CORE_DATAPATH__abc_16259_n3946) );
  AND2X2 AND2X2_795 ( .A(AES_CORE_DATAPATH__abc_16259_n3944), .B(AES_CORE_DATAPATH__abc_16259_n3948), .Y(AES_CORE_DATAPATH__abc_16259_n3949) );
  AND2X2 AND2X2_796 ( .A(AES_CORE_DATAPATH__abc_16259_n3949), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n3950_1) );
  AND2X2 AND2X2_797 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf10), .B(AES_CORE_DATAPATH_col_3__27_), .Y(AES_CORE_DATAPATH__abc_16259_n3951_1) );
  AND2X2 AND2X2_798 ( .A(AES_CORE_DATAPATH__abc_16259_n3954), .B(AES_CORE_DATAPATH__abc_16259_n3956), .Y(AES_CORE_DATAPATH__abc_16259_n3957) );
  AND2X2 AND2X2_799 ( .A(AES_CORE_DATAPATH__abc_16259_n2782_bF_buf1), .B(AES_CORE_DATAPATH_col_3__28_), .Y(AES_CORE_DATAPATH__abc_16259_n3958_1) );
  AND2X2 AND2X2_8 ( .A(\addr[1] ), .B(read_en), .Y(AES_CORE_DATAPATH_col_sel_host_1_) );
  AND2X2 AND2X2_80 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n195), .B(AES_CORE_CONTROL_UNIT_state_6_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n218) );
  AND2X2 AND2X2_800 ( .A(AES_CORE_DATAPATH__abc_16259_n2786_bF_buf1), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_92_), .Y(AES_CORE_DATAPATH__abc_16259_n3959_1) );
  AND2X2 AND2X2_801 ( .A(AES_CORE_DATAPATH__abc_16259_n2789_bF_buf1), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_60_), .Y(AES_CORE_DATAPATH__abc_16259_n3960) );
  AND2X2 AND2X2_802 ( .A(AES_CORE_DATAPATH__abc_16259_n3963), .B(AES_CORE_DATAPATH__abc_16259_n3957), .Y(AES_CORE_DATAPATH__abc_16259_n3964) );
  AND2X2 AND2X2_803 ( .A(AES_CORE_DATAPATH__abc_16259_n2837_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__28_), .Y(AES_CORE_DATAPATH__abc_16259_n3966_1) );
  AND2X2 AND2X2_804 ( .A(AES_CORE_DATAPATH__abc_16259_n2887_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__28_), .Y(AES_CORE_DATAPATH__abc_16259_n3968) );
  AND2X2 AND2X2_805 ( .A(AES_CORE_DATAPATH__abc_16259_n2830_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__28_), .Y(AES_CORE_DATAPATH__abc_16259_n3969_1) );
  AND2X2 AND2X2_806 ( .A(AES_CORE_DATAPATH__abc_16259_n3971), .B(AES_CORE_DATAPATH__abc_16259_n3972), .Y(_auto_iopadmap_cc_313_execute_26949_28_) );
  AND2X2 AND2X2_807 ( .A(AES_CORE_DATAPATH__abc_16259_n2855_bF_buf1), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_28_), .Y(AES_CORE_DATAPATH__abc_16259_n3975_1) );
  AND2X2 AND2X2_808 ( .A(AES_CORE_DATAPATH__abc_16259_n2857_bF_buf1), .B(AES_CORE_DATAPATH_MIX_COL_col_3__4_), .Y(AES_CORE_DATAPATH__abc_16259_n3976) );
  AND2X2 AND2X2_809 ( .A(AES_CORE_DATAPATH__abc_16259_n3974_1), .B(AES_CORE_DATAPATH__abc_16259_n3978), .Y(AES_CORE_DATAPATH__abc_16259_n3979) );
  AND2X2 AND2X2_81 ( .A(AES_CORE_CONTROL_UNIT_last_round_bF_buf4), .B(AES_CORE_CONTROL_UNIT_state_9_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n219) );
  AND2X2 AND2X2_810 ( .A(_auto_iopadmap_cc_313_execute_26949_28_), .B(AES_CORE_DATAPATH__abc_16259_n3979), .Y(AES_CORE_DATAPATH__abc_16259_n3982_1) );
  AND2X2 AND2X2_811 ( .A(AES_CORE_DATAPATH_last_round_pp2_bF_buf0), .B(AES_CORE_DATAPATH_MIX_COL_col_3__4_), .Y(AES_CORE_DATAPATH__abc_16259_n3985_1) );
  AND2X2 AND2X2_812 ( .A(AES_CORE_DATAPATH__abc_16259_n2798_bF_buf1), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_28_), .Y(AES_CORE_DATAPATH__abc_16259_n3986) );
  AND2X2 AND2X2_813 ( .A(AES_CORE_DATAPATH__abc_16259_n3984), .B(AES_CORE_DATAPATH__abc_16259_n3988), .Y(AES_CORE_DATAPATH__abc_16259_n3989) );
  AND2X2 AND2X2_814 ( .A(AES_CORE_DATAPATH__abc_16259_n3989), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n3990_1) );
  AND2X2 AND2X2_815 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf9), .B(AES_CORE_DATAPATH_col_3__28_), .Y(AES_CORE_DATAPATH__abc_16259_n3991_1) );
  AND2X2 AND2X2_816 ( .A(AES_CORE_DATAPATH__abc_16259_n3994), .B(AES_CORE_DATAPATH__abc_16259_n3996), .Y(AES_CORE_DATAPATH__abc_16259_n3997) );
  AND2X2 AND2X2_817 ( .A(AES_CORE_DATAPATH__abc_16259_n2782_bF_buf0), .B(AES_CORE_DATAPATH_col_3__29_), .Y(AES_CORE_DATAPATH__abc_16259_n3998_1) );
  AND2X2 AND2X2_818 ( .A(AES_CORE_DATAPATH__abc_16259_n2786_bF_buf0), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_93_), .Y(AES_CORE_DATAPATH__abc_16259_n3999_1) );
  AND2X2 AND2X2_819 ( .A(AES_CORE_DATAPATH__abc_16259_n2789_bF_buf0), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_61_), .Y(AES_CORE_DATAPATH__abc_16259_n4000) );
  AND2X2 AND2X2_82 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n222), .B(AES_CORE_CONTROL_UNIT__abc_15841_n217), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n223) );
  AND2X2 AND2X2_820 ( .A(AES_CORE_DATAPATH__abc_16259_n4003), .B(AES_CORE_DATAPATH__abc_16259_n3997), .Y(AES_CORE_DATAPATH__abc_16259_n4004) );
  AND2X2 AND2X2_821 ( .A(AES_CORE_DATAPATH__abc_16259_n2837_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__29_), .Y(AES_CORE_DATAPATH__abc_16259_n4006_1) );
  AND2X2 AND2X2_822 ( .A(AES_CORE_DATAPATH__abc_16259_n2887_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__29_), .Y(AES_CORE_DATAPATH__abc_16259_n4008) );
  AND2X2 AND2X2_823 ( .A(AES_CORE_DATAPATH__abc_16259_n2830_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__29_), .Y(AES_CORE_DATAPATH__abc_16259_n4009_1) );
  AND2X2 AND2X2_824 ( .A(AES_CORE_DATAPATH__abc_16259_n4011), .B(AES_CORE_DATAPATH__abc_16259_n4012), .Y(_auto_iopadmap_cc_313_execute_26949_29_) );
  AND2X2 AND2X2_825 ( .A(AES_CORE_DATAPATH__abc_16259_n2855_bF_buf0), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_29_), .Y(AES_CORE_DATAPATH__abc_16259_n4015_1) );
  AND2X2 AND2X2_826 ( .A(AES_CORE_DATAPATH__abc_16259_n2857_bF_buf0), .B(AES_CORE_DATAPATH_MIX_COL_col_3__5_), .Y(AES_CORE_DATAPATH__abc_16259_n4016) );
  AND2X2 AND2X2_827 ( .A(AES_CORE_DATAPATH__abc_16259_n4014_1), .B(AES_CORE_DATAPATH__abc_16259_n4018), .Y(AES_CORE_DATAPATH__abc_16259_n4019) );
  AND2X2 AND2X2_828 ( .A(_auto_iopadmap_cc_313_execute_26949_29_), .B(AES_CORE_DATAPATH__abc_16259_n4019), .Y(AES_CORE_DATAPATH__abc_16259_n4022_1) );
  AND2X2 AND2X2_829 ( .A(AES_CORE_DATAPATH_last_round_pp2_bF_buf4), .B(AES_CORE_DATAPATH_MIX_COL_col_3__5_), .Y(AES_CORE_DATAPATH__abc_16259_n4025_1) );
  AND2X2 AND2X2_83 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n216), .B(AES_CORE_CONTROL_UNIT__abc_15841_n190), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n225) );
  AND2X2 AND2X2_830 ( .A(AES_CORE_DATAPATH__abc_16259_n2798_bF_buf0), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_29_), .Y(AES_CORE_DATAPATH__abc_16259_n4026) );
  AND2X2 AND2X2_831 ( .A(AES_CORE_DATAPATH__abc_16259_n4024), .B(AES_CORE_DATAPATH__abc_16259_n4028), .Y(AES_CORE_DATAPATH__abc_16259_n4029) );
  AND2X2 AND2X2_832 ( .A(AES_CORE_DATAPATH__abc_16259_n4029), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n4030_1) );
  AND2X2 AND2X2_833 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf8), .B(AES_CORE_DATAPATH_col_3__29_), .Y(AES_CORE_DATAPATH__abc_16259_n4031_1) );
  AND2X2 AND2X2_834 ( .A(AES_CORE_DATAPATH__abc_16259_n4034), .B(AES_CORE_DATAPATH__abc_16259_n4036), .Y(AES_CORE_DATAPATH__abc_16259_n4037) );
  AND2X2 AND2X2_835 ( .A(AES_CORE_DATAPATH__abc_16259_n2782_bF_buf4), .B(AES_CORE_DATAPATH_col_3__30_), .Y(AES_CORE_DATAPATH__abc_16259_n4038_1) );
  AND2X2 AND2X2_836 ( .A(AES_CORE_DATAPATH__abc_16259_n2786_bF_buf4), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_94_), .Y(AES_CORE_DATAPATH__abc_16259_n4039_1) );
  AND2X2 AND2X2_837 ( .A(AES_CORE_DATAPATH__abc_16259_n2789_bF_buf4), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_62_), .Y(AES_CORE_DATAPATH__abc_16259_n4040) );
  AND2X2 AND2X2_838 ( .A(AES_CORE_DATAPATH__abc_16259_n4043), .B(AES_CORE_DATAPATH__abc_16259_n4037), .Y(AES_CORE_DATAPATH__abc_16259_n4044) );
  AND2X2 AND2X2_839 ( .A(AES_CORE_DATAPATH__abc_16259_n2837_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__30_), .Y(AES_CORE_DATAPATH__abc_16259_n4046_1) );
  AND2X2 AND2X2_84 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n226), .B(AES_CORE_CONTROL_UNIT__abc_15841_n227), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n228) );
  AND2X2 AND2X2_840 ( .A(AES_CORE_DATAPATH__abc_16259_n2887_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__30_), .Y(AES_CORE_DATAPATH__abc_16259_n4048) );
  AND2X2 AND2X2_841 ( .A(AES_CORE_DATAPATH__abc_16259_n2830_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__30_), .Y(AES_CORE_DATAPATH__abc_16259_n4049_1) );
  AND2X2 AND2X2_842 ( .A(AES_CORE_DATAPATH__abc_16259_n4051), .B(AES_CORE_DATAPATH__abc_16259_n4052), .Y(_auto_iopadmap_cc_313_execute_26949_30_) );
  AND2X2 AND2X2_843 ( .A(AES_CORE_DATAPATH__abc_16259_n2855_bF_buf4), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_30_), .Y(AES_CORE_DATAPATH__abc_16259_n4055_1) );
  AND2X2 AND2X2_844 ( .A(AES_CORE_DATAPATH__abc_16259_n2857_bF_buf4), .B(AES_CORE_DATAPATH_MIX_COL_col_3__6_), .Y(AES_CORE_DATAPATH__abc_16259_n4056) );
  AND2X2 AND2X2_845 ( .A(AES_CORE_DATAPATH__abc_16259_n4054_1), .B(AES_CORE_DATAPATH__abc_16259_n4058), .Y(AES_CORE_DATAPATH__abc_16259_n4059) );
  AND2X2 AND2X2_846 ( .A(_auto_iopadmap_cc_313_execute_26949_30_), .B(AES_CORE_DATAPATH__abc_16259_n4059), .Y(AES_CORE_DATAPATH__abc_16259_n4062_1) );
  AND2X2 AND2X2_847 ( .A(AES_CORE_DATAPATH_last_round_pp2_bF_buf3), .B(AES_CORE_DATAPATH_MIX_COL_col_3__6_), .Y(AES_CORE_DATAPATH__abc_16259_n4065_1) );
  AND2X2 AND2X2_848 ( .A(AES_CORE_DATAPATH__abc_16259_n2798_bF_buf4), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_30_), .Y(AES_CORE_DATAPATH__abc_16259_n4066) );
  AND2X2 AND2X2_849 ( .A(AES_CORE_DATAPATH__abc_16259_n4064), .B(AES_CORE_DATAPATH__abc_16259_n4068), .Y(AES_CORE_DATAPATH__abc_16259_n4069) );
  AND2X2 AND2X2_85 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n229), .B(AES_CORE_CONTROL_UNIT__abc_15841_n230), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n231) );
  AND2X2 AND2X2_850 ( .A(AES_CORE_DATAPATH__abc_16259_n4069), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n4070_1) );
  AND2X2 AND2X2_851 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf7), .B(AES_CORE_DATAPATH_col_3__30_), .Y(AES_CORE_DATAPATH__abc_16259_n4071_1) );
  AND2X2 AND2X2_852 ( .A(AES_CORE_DATAPATH__abc_16259_n4074), .B(AES_CORE_DATAPATH__abc_16259_n4076), .Y(AES_CORE_DATAPATH__abc_16259_n4077) );
  AND2X2 AND2X2_853 ( .A(AES_CORE_DATAPATH__abc_16259_n2782_bF_buf3), .B(AES_CORE_DATAPATH_col_3__31_), .Y(AES_CORE_DATAPATH__abc_16259_n4078_1) );
  AND2X2 AND2X2_854 ( .A(AES_CORE_DATAPATH__abc_16259_n2786_bF_buf3), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_95_), .Y(AES_CORE_DATAPATH__abc_16259_n4079_1) );
  AND2X2 AND2X2_855 ( .A(AES_CORE_DATAPATH__abc_16259_n2789_bF_buf3), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_63_), .Y(AES_CORE_DATAPATH__abc_16259_n4080) );
  AND2X2 AND2X2_856 ( .A(AES_CORE_DATAPATH__abc_16259_n4083), .B(AES_CORE_DATAPATH__abc_16259_n4077), .Y(AES_CORE_DATAPATH__abc_16259_n4084) );
  AND2X2 AND2X2_857 ( .A(AES_CORE_DATAPATH__abc_16259_n2837_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__31_), .Y(AES_CORE_DATAPATH__abc_16259_n4086_1) );
  AND2X2 AND2X2_858 ( .A(AES_CORE_DATAPATH__abc_16259_n2887_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__31_), .Y(AES_CORE_DATAPATH__abc_16259_n4088) );
  AND2X2 AND2X2_859 ( .A(AES_CORE_DATAPATH__abc_16259_n2830_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__31_), .Y(AES_CORE_DATAPATH__abc_16259_n4089_1) );
  AND2X2 AND2X2_86 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n228), .B(AES_CORE_CONTROL_UNIT__abc_15841_n231), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n232) );
  AND2X2 AND2X2_860 ( .A(AES_CORE_DATAPATH__abc_16259_n4091), .B(AES_CORE_DATAPATH__abc_16259_n4092), .Y(_auto_iopadmap_cc_313_execute_26949_31_) );
  AND2X2 AND2X2_861 ( .A(AES_CORE_DATAPATH__abc_16259_n2855_bF_buf3), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_31_), .Y(AES_CORE_DATAPATH__abc_16259_n4095_1) );
  AND2X2 AND2X2_862 ( .A(AES_CORE_DATAPATH__abc_16259_n2857_bF_buf3), .B(AES_CORE_DATAPATH_MIX_COL_col_3__7_), .Y(AES_CORE_DATAPATH__abc_16259_n4096) );
  AND2X2 AND2X2_863 ( .A(AES_CORE_DATAPATH__abc_16259_n4094_1), .B(AES_CORE_DATAPATH__abc_16259_n4098), .Y(AES_CORE_DATAPATH__abc_16259_n4099) );
  AND2X2 AND2X2_864 ( .A(_auto_iopadmap_cc_313_execute_26949_31_), .B(AES_CORE_DATAPATH__abc_16259_n4099), .Y(AES_CORE_DATAPATH__abc_16259_n4102_1) );
  AND2X2 AND2X2_865 ( .A(AES_CORE_DATAPATH_last_round_pp2_bF_buf2), .B(AES_CORE_DATAPATH_MIX_COL_col_3__7_), .Y(AES_CORE_DATAPATH__abc_16259_n4105_1) );
  AND2X2 AND2X2_866 ( .A(AES_CORE_DATAPATH__abc_16259_n2798_bF_buf3), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_31_), .Y(AES_CORE_DATAPATH__abc_16259_n4106) );
  AND2X2 AND2X2_867 ( .A(AES_CORE_DATAPATH__abc_16259_n4104), .B(AES_CORE_DATAPATH__abc_16259_n4108), .Y(AES_CORE_DATAPATH__abc_16259_n4109) );
  AND2X2 AND2X2_868 ( .A(AES_CORE_DATAPATH__abc_16259_n4109), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n4110_1) );
  AND2X2 AND2X2_869 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf6), .B(AES_CORE_DATAPATH_col_3__31_), .Y(AES_CORE_DATAPATH__abc_16259_n4111_1) );
  AND2X2 AND2X2_87 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n106_1), .B(AES_CORE_CONTROL_UNIT__abc_15841_n138), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n236) );
  AND2X2 AND2X2_870 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf2), .B(AES_CORE_DATAPATH_col_0__0_), .Y(AES_CORE_DATAPATH__abc_16259_n4113_1) );
  AND2X2 AND2X2_871 ( .A(AES_CORE_DATAPATH__abc_16259_n2868_1), .B(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n4114) );
  AND2X2 AND2X2_872 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf1), .B(AES_CORE_DATAPATH_col_0__1_), .Y(AES_CORE_DATAPATH__abc_16259_n4116) );
  AND2X2 AND2X2_873 ( .A(AES_CORE_DATAPATH__abc_16259_n2909_1), .B(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n4117) );
  AND2X2 AND2X2_874 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf0), .B(AES_CORE_DATAPATH_col_0__2_), .Y(AES_CORE_DATAPATH__abc_16259_n4119_1) );
  AND2X2 AND2X2_875 ( .A(AES_CORE_DATAPATH__abc_16259_n2949_1), .B(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n4120) );
  AND2X2 AND2X2_876 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf14), .B(AES_CORE_DATAPATH_col_0__3_), .Y(AES_CORE_DATAPATH__abc_16259_n4122) );
  AND2X2 AND2X2_877 ( .A(AES_CORE_DATAPATH__abc_16259_n2989), .B(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n4123) );
  AND2X2 AND2X2_878 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf13), .B(AES_CORE_DATAPATH_col_0__4_), .Y(AES_CORE_DATAPATH__abc_16259_n4125) );
  AND2X2 AND2X2_879 ( .A(AES_CORE_DATAPATH__abc_16259_n3029), .B(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n4126_1) );
  AND2X2 AND2X2_88 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n106_1), .B(AES_CORE_CONTROL_UNIT__abc_15841_n198), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n241) );
  AND2X2 AND2X2_880 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf12), .B(AES_CORE_DATAPATH_col_0__5_), .Y(AES_CORE_DATAPATH__abc_16259_n4128) );
  AND2X2 AND2X2_881 ( .A(AES_CORE_DATAPATH__abc_16259_n3069_1), .B(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n4129_1) );
  AND2X2 AND2X2_882 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf11), .B(AES_CORE_DATAPATH_col_0__6_), .Y(AES_CORE_DATAPATH__abc_16259_n4131) );
  AND2X2 AND2X2_883 ( .A(AES_CORE_DATAPATH__abc_16259_n3109), .B(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf12), .Y(AES_CORE_DATAPATH__abc_16259_n4132) );
  AND2X2 AND2X2_884 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf10), .B(AES_CORE_DATAPATH_col_0__7_), .Y(AES_CORE_DATAPATH__abc_16259_n4134_1) );
  AND2X2 AND2X2_885 ( .A(AES_CORE_DATAPATH__abc_16259_n3149_1), .B(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf11), .Y(AES_CORE_DATAPATH__abc_16259_n4135_1) );
  AND2X2 AND2X2_886 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf9), .B(AES_CORE_DATAPATH_col_0__8_), .Y(AES_CORE_DATAPATH__abc_16259_n4137_1) );
  AND2X2 AND2X2_887 ( .A(AES_CORE_DATAPATH__abc_16259_n3189), .B(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf10), .Y(AES_CORE_DATAPATH__abc_16259_n4138) );
  AND2X2 AND2X2_888 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf8), .B(AES_CORE_DATAPATH_col_0__9_), .Y(AES_CORE_DATAPATH__abc_16259_n4140) );
  AND2X2 AND2X2_889 ( .A(AES_CORE_DATAPATH__abc_16259_n3229), .B(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf9), .Y(AES_CORE_DATAPATH__abc_16259_n4141) );
  AND2X2 AND2X2_89 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n106_1), .B(AES_CORE_CONTROL_UNIT__abc_15841_n203_1), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n244) );
  AND2X2 AND2X2_890 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf7), .B(AES_CORE_DATAPATH_col_0__10_), .Y(AES_CORE_DATAPATH__abc_16259_n4143_1) );
  AND2X2 AND2X2_891 ( .A(AES_CORE_DATAPATH__abc_16259_n3269), .B(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf8), .Y(AES_CORE_DATAPATH__abc_16259_n4144) );
  AND2X2 AND2X2_892 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf6), .B(AES_CORE_DATAPATH_col_0__11_), .Y(AES_CORE_DATAPATH__abc_16259_n4146) );
  AND2X2 AND2X2_893 ( .A(AES_CORE_DATAPATH__abc_16259_n3309), .B(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n4147) );
  AND2X2 AND2X2_894 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf5), .B(AES_CORE_DATAPATH_col_0__12_), .Y(AES_CORE_DATAPATH__abc_16259_n4149) );
  AND2X2 AND2X2_895 ( .A(AES_CORE_DATAPATH__abc_16259_n3349), .B(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n4150_1) );
  AND2X2 AND2X2_896 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf4), .B(AES_CORE_DATAPATH_col_0__13_), .Y(AES_CORE_DATAPATH__abc_16259_n4152) );
  AND2X2 AND2X2_897 ( .A(AES_CORE_DATAPATH__abc_16259_n3389), .B(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n4153_1) );
  AND2X2 AND2X2_898 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf3), .B(AES_CORE_DATAPATH_col_0__14_), .Y(AES_CORE_DATAPATH__abc_16259_n4155) );
  AND2X2 AND2X2_899 ( .A(AES_CORE_DATAPATH__abc_16259_n3429), .B(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n4156) );
  AND2X2 AND2X2_9 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n73), .B(\aes_mode[1] ), .Y(AES_CORE_CONTROL_UNIT_mode_ctr) );
  AND2X2 AND2X2_90 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf7), .B(AES_CORE_CONTROL_UNIT_state_1_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n247) );
  AND2X2 AND2X2_900 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf2), .B(AES_CORE_DATAPATH_col_0__15_), .Y(AES_CORE_DATAPATH__abc_16259_n4158_1) );
  AND2X2 AND2X2_901 ( .A(AES_CORE_DATAPATH__abc_16259_n3469), .B(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n4159_1) );
  AND2X2 AND2X2_902 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf1), .B(AES_CORE_DATAPATH_col_0__16_), .Y(AES_CORE_DATAPATH__abc_16259_n4161_1) );
  AND2X2 AND2X2_903 ( .A(AES_CORE_DATAPATH__abc_16259_n3509), .B(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n4162) );
  AND2X2 AND2X2_904 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf0), .B(AES_CORE_DATAPATH_col_0__17_), .Y(AES_CORE_DATAPATH__abc_16259_n4164) );
  AND2X2 AND2X2_905 ( .A(AES_CORE_DATAPATH__abc_16259_n3549_1), .B(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n4165) );
  AND2X2 AND2X2_906 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf14), .B(AES_CORE_DATAPATH_col_0__18_), .Y(AES_CORE_DATAPATH__abc_16259_n4167_1) );
  AND2X2 AND2X2_907 ( .A(AES_CORE_DATAPATH__abc_16259_n3589_1), .B(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n4168) );
  AND2X2 AND2X2_908 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf13), .B(AES_CORE_DATAPATH_col_0__19_), .Y(AES_CORE_DATAPATH__abc_16259_n4170) );
  AND2X2 AND2X2_909 ( .A(AES_CORE_DATAPATH__abc_16259_n3629), .B(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf12), .Y(AES_CORE_DATAPATH__abc_16259_n4171) );
  AND2X2 AND2X2_91 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n106_1), .B(AES_CORE_CONTROL_UNIT__abc_15841_n206_1), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n248) );
  AND2X2 AND2X2_910 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf12), .B(AES_CORE_DATAPATH_col_0__20_), .Y(AES_CORE_DATAPATH__abc_16259_n4173) );
  AND2X2 AND2X2_911 ( .A(AES_CORE_DATAPATH__abc_16259_n3669), .B(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf11), .Y(AES_CORE_DATAPATH__abc_16259_n4174_1) );
  AND2X2 AND2X2_912 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf11), .B(AES_CORE_DATAPATH_col_0__21_), .Y(AES_CORE_DATAPATH__abc_16259_n4176) );
  AND2X2 AND2X2_913 ( .A(AES_CORE_DATAPATH__abc_16259_n3709), .B(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf10), .Y(AES_CORE_DATAPATH__abc_16259_n4177_1) );
  AND2X2 AND2X2_914 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf10), .B(AES_CORE_DATAPATH_col_0__22_), .Y(AES_CORE_DATAPATH__abc_16259_n4179) );
  AND2X2 AND2X2_915 ( .A(AES_CORE_DATAPATH__abc_16259_n3749), .B(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf9), .Y(AES_CORE_DATAPATH__abc_16259_n4180) );
  AND2X2 AND2X2_916 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf9), .B(AES_CORE_DATAPATH_col_0__23_), .Y(AES_CORE_DATAPATH__abc_16259_n4182_1) );
  AND2X2 AND2X2_917 ( .A(AES_CORE_DATAPATH__abc_16259_n3789), .B(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf8), .Y(AES_CORE_DATAPATH__abc_16259_n4183_1) );
  AND2X2 AND2X2_918 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf8), .B(AES_CORE_DATAPATH_col_0__24_), .Y(AES_CORE_DATAPATH__abc_16259_n4185_1) );
  AND2X2 AND2X2_919 ( .A(AES_CORE_DATAPATH__abc_16259_n3829), .B(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n4186) );
  AND2X2 AND2X2_92 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n84_1), .B(AES_CORE_CONTROL_UNIT_state_11_), .Y(AES_CORE_CONTROL_UNIT__abc_10818_n303) );
  AND2X2 AND2X2_920 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf7), .B(AES_CORE_DATAPATH_col_0__25_), .Y(AES_CORE_DATAPATH__abc_16259_n4188) );
  AND2X2 AND2X2_921 ( .A(AES_CORE_DATAPATH__abc_16259_n3869), .B(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n4189) );
  AND2X2 AND2X2_922 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf6), .B(AES_CORE_DATAPATH_col_0__26_), .Y(AES_CORE_DATAPATH__abc_16259_n4191_1) );
  AND2X2 AND2X2_923 ( .A(AES_CORE_DATAPATH__abc_16259_n3909), .B(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n4192) );
  AND2X2 AND2X2_924 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf5), .B(AES_CORE_DATAPATH_col_0__27_), .Y(AES_CORE_DATAPATH__abc_16259_n4194) );
  AND2X2 AND2X2_925 ( .A(AES_CORE_DATAPATH__abc_16259_n3949), .B(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n4195) );
  AND2X2 AND2X2_926 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf4), .B(AES_CORE_DATAPATH_col_0__28_), .Y(AES_CORE_DATAPATH__abc_16259_n4197) );
  AND2X2 AND2X2_927 ( .A(AES_CORE_DATAPATH__abc_16259_n3989), .B(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n4198_1) );
  AND2X2 AND2X2_928 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf3), .B(AES_CORE_DATAPATH_col_0__29_), .Y(AES_CORE_DATAPATH__abc_16259_n4200) );
  AND2X2 AND2X2_929 ( .A(AES_CORE_DATAPATH__abc_16259_n4029), .B(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n4201_1) );
  AND2X2 AND2X2_93 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n84_1), .B(AES_CORE_CONTROL_UNIT_state_3_), .Y(AES_CORE_CONTROL_UNIT__abc_10818_n306) );
  AND2X2 AND2X2_930 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf2), .B(AES_CORE_DATAPATH_col_0__30_), .Y(AES_CORE_DATAPATH__abc_16259_n4203) );
  AND2X2 AND2X2_931 ( .A(AES_CORE_DATAPATH__abc_16259_n4069), .B(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n4204) );
  AND2X2 AND2X2_932 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf1), .B(AES_CORE_DATAPATH_col_0__31_), .Y(AES_CORE_DATAPATH__abc_16259_n4206_1) );
  AND2X2 AND2X2_933 ( .A(AES_CORE_DATAPATH__abc_16259_n4109), .B(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n4207_1) );
  AND2X2 AND2X2_934 ( .A(_auto_iopadmap_cc_313_execute_26949_0_), .B(AES_CORE_DATAPATH__abc_16259_n4210), .Y(AES_CORE_DATAPATH__abc_16259_n4211) );
  AND2X2 AND2X2_935 ( .A(AES_CORE_DATAPATH__abc_16259_n4212), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_1_2_), .Y(AES_CORE_DATAPATH__abc_16259_n4213) );
  AND2X2 AND2X2_936 ( .A(AES_CORE_DATAPATH__abc_16259_n4215_1), .B(AES_CORE_DATAPATH__abc_16259_n4209_1), .Y(AES_CORE_DATAPATH_sbox_pp2_0__FF_INPUT) );
  AND2X2 AND2X2_937 ( .A(_auto_iopadmap_cc_313_execute_26949_1_), .B(AES_CORE_DATAPATH__abc_16259_n4218), .Y(AES_CORE_DATAPATH__abc_16259_n4219) );
  AND2X2 AND2X2_938 ( .A(AES_CORE_DATAPATH__abc_16259_n4220), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_1_), .Y(AES_CORE_DATAPATH__abc_16259_n4221) );
  AND2X2 AND2X2_939 ( .A(AES_CORE_DATAPATH__abc_16259_n4223_1), .B(AES_CORE_DATAPATH__abc_16259_n4217_1), .Y(AES_CORE_DATAPATH_sbox_pp2_1__FF_INPUT) );
  AND2X2 AND2X2_94 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n154), .B(AES_CORE_CONTROL_UNIT__abc_15841_n121), .Y(AES_CORE_CONTROL_UNIT__abc_10818_n307) );
  AND2X2 AND2X2_940 ( .A(_auto_iopadmap_cc_313_execute_26949_2_), .B(AES_CORE_DATAPATH__abc_16259_n4226), .Y(AES_CORE_DATAPATH__abc_16259_n4227) );
  AND2X2 AND2X2_941 ( .A(AES_CORE_DATAPATH__abc_16259_n4228), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_2_), .Y(AES_CORE_DATAPATH__abc_16259_n4229) );
  AND2X2 AND2X2_942 ( .A(AES_CORE_DATAPATH__abc_16259_n4231_1), .B(AES_CORE_DATAPATH__abc_16259_n4225_1), .Y(AES_CORE_DATAPATH_sbox_pp2_2__FF_INPUT) );
  AND2X2 AND2X2_943 ( .A(_auto_iopadmap_cc_313_execute_26949_3_), .B(AES_CORE_DATAPATH__abc_16259_n4234), .Y(AES_CORE_DATAPATH__abc_16259_n4235) );
  AND2X2 AND2X2_944 ( .A(AES_CORE_DATAPATH__abc_16259_n4236), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_3_), .Y(AES_CORE_DATAPATH__abc_16259_n4237) );
  AND2X2 AND2X2_945 ( .A(AES_CORE_DATAPATH__abc_16259_n4239_1), .B(AES_CORE_DATAPATH__abc_16259_n4233_1), .Y(AES_CORE_DATAPATH_sbox_pp2_3__FF_INPUT) );
  AND2X2 AND2X2_946 ( .A(_auto_iopadmap_cc_313_execute_26949_4_), .B(AES_CORE_DATAPATH__abc_16259_n4242), .Y(AES_CORE_DATAPATH__abc_16259_n4243) );
  AND2X2 AND2X2_947 ( .A(AES_CORE_DATAPATH__abc_16259_n4244), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_4_), .Y(AES_CORE_DATAPATH__abc_16259_n4245) );
  AND2X2 AND2X2_948 ( .A(AES_CORE_DATAPATH__abc_16259_n4247_1), .B(AES_CORE_DATAPATH__abc_16259_n4241_1), .Y(AES_CORE_DATAPATH_sbox_pp2_4__FF_INPUT) );
  AND2X2 AND2X2_949 ( .A(_auto_iopadmap_cc_313_execute_26949_5_), .B(AES_CORE_DATAPATH__abc_16259_n4250), .Y(AES_CORE_DATAPATH__abc_16259_n4251) );
  AND2X2 AND2X2_95 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n91), .B(_auto_iopadmap_cc_313_execute_26914), .Y(AES_CORE_CONTROL_UNIT_key_derivation_en) );
  AND2X2 AND2X2_950 ( .A(AES_CORE_DATAPATH__abc_16259_n4252), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_5_), .Y(AES_CORE_DATAPATH__abc_16259_n4253) );
  AND2X2 AND2X2_951 ( .A(AES_CORE_DATAPATH__abc_16259_n4255_1), .B(AES_CORE_DATAPATH__abc_16259_n4249_1), .Y(AES_CORE_DATAPATH_sbox_pp2_5__FF_INPUT) );
  AND2X2 AND2X2_952 ( .A(_auto_iopadmap_cc_313_execute_26949_6_), .B(AES_CORE_DATAPATH__abc_16259_n4258), .Y(AES_CORE_DATAPATH__abc_16259_n4259) );
  AND2X2 AND2X2_953 ( .A(AES_CORE_DATAPATH__abc_16259_n4260), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_6_), .Y(AES_CORE_DATAPATH__abc_16259_n4261) );
  AND2X2 AND2X2_954 ( .A(AES_CORE_DATAPATH__abc_16259_n4263_1), .B(AES_CORE_DATAPATH__abc_16259_n4257_1), .Y(AES_CORE_DATAPATH_sbox_pp2_6__FF_INPUT) );
  AND2X2 AND2X2_955 ( .A(_auto_iopadmap_cc_313_execute_26949_7_), .B(AES_CORE_DATAPATH__abc_16259_n4266), .Y(AES_CORE_DATAPATH__abc_16259_n4267) );
  AND2X2 AND2X2_956 ( .A(AES_CORE_DATAPATH__abc_16259_n4268), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_7_), .Y(AES_CORE_DATAPATH__abc_16259_n4269) );
  AND2X2 AND2X2_957 ( .A(AES_CORE_DATAPATH__abc_16259_n4271_1), .B(AES_CORE_DATAPATH__abc_16259_n4265_1), .Y(AES_CORE_DATAPATH_sbox_pp2_7__FF_INPUT) );
  AND2X2 AND2X2_958 ( .A(_auto_iopadmap_cc_313_execute_26949_8_), .B(AES_CORE_DATAPATH__abc_16259_n4274), .Y(AES_CORE_DATAPATH__abc_16259_n4275) );
  AND2X2 AND2X2_959 ( .A(AES_CORE_DATAPATH__abc_16259_n4276), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_1_2_), .Y(AES_CORE_DATAPATH__abc_16259_n4277) );
  AND2X2 AND2X2_96 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n213), .B(AES_CORE_CONTROL_UNIT_state_9_), .Y(AES_CORE_CONTROL_UNIT_iv_cnt_en) );
  AND2X2 AND2X2_960 ( .A(AES_CORE_DATAPATH__abc_16259_n4279_1), .B(AES_CORE_DATAPATH__abc_16259_n4273_1), .Y(AES_CORE_DATAPATH_sbox_pp2_8__FF_INPUT) );
  AND2X2 AND2X2_961 ( .A(_auto_iopadmap_cc_313_execute_26949_9_), .B(AES_CORE_DATAPATH__abc_16259_n4282), .Y(AES_CORE_DATAPATH__abc_16259_n4283) );
  AND2X2 AND2X2_962 ( .A(AES_CORE_DATAPATH__abc_16259_n4284), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_1_), .Y(AES_CORE_DATAPATH__abc_16259_n4285) );
  AND2X2 AND2X2_963 ( .A(AES_CORE_DATAPATH__abc_16259_n4287_1), .B(AES_CORE_DATAPATH__abc_16259_n4281_1), .Y(AES_CORE_DATAPATH_sbox_pp2_9__FF_INPUT) );
  AND2X2 AND2X2_964 ( .A(_auto_iopadmap_cc_313_execute_26949_10_), .B(AES_CORE_DATAPATH__abc_16259_n4290), .Y(AES_CORE_DATAPATH__abc_16259_n4291) );
  AND2X2 AND2X2_965 ( .A(AES_CORE_DATAPATH__abc_16259_n4292), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_2_), .Y(AES_CORE_DATAPATH__abc_16259_n4293) );
  AND2X2 AND2X2_966 ( .A(AES_CORE_DATAPATH__abc_16259_n4295_1), .B(AES_CORE_DATAPATH__abc_16259_n4289_1), .Y(AES_CORE_DATAPATH_sbox_pp2_10__FF_INPUT) );
  AND2X2 AND2X2_967 ( .A(_auto_iopadmap_cc_313_execute_26949_11_), .B(AES_CORE_DATAPATH__abc_16259_n4298), .Y(AES_CORE_DATAPATH__abc_16259_n4299) );
  AND2X2 AND2X2_968 ( .A(AES_CORE_DATAPATH__abc_16259_n4300), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_3_), .Y(AES_CORE_DATAPATH__abc_16259_n4301) );
  AND2X2 AND2X2_969 ( .A(AES_CORE_DATAPATH__abc_16259_n4303_1), .B(AES_CORE_DATAPATH__abc_16259_n4297_1), .Y(AES_CORE_DATAPATH_sbox_pp2_11__FF_INPUT) );
  AND2X2 AND2X2_97 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n84_1), .B(AES_CORE_CONTROL_UNIT_state_13_), .Y(AES_CORE_CONTROL_UNIT__abc_10818_n310) );
  AND2X2 AND2X2_970 ( .A(_auto_iopadmap_cc_313_execute_26949_12_), .B(AES_CORE_DATAPATH__abc_16259_n4306), .Y(AES_CORE_DATAPATH__abc_16259_n4307) );
  AND2X2 AND2X2_971 ( .A(AES_CORE_DATAPATH__abc_16259_n4308), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_4_), .Y(AES_CORE_DATAPATH__abc_16259_n4309) );
  AND2X2 AND2X2_972 ( .A(AES_CORE_DATAPATH__abc_16259_n4311_1), .B(AES_CORE_DATAPATH__abc_16259_n4305_1), .Y(AES_CORE_DATAPATH_sbox_pp2_12__FF_INPUT) );
  AND2X2 AND2X2_973 ( .A(AES_CORE_DATAPATH__abc_16259_n2807_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_13_), .Y(AES_CORE_DATAPATH__abc_16259_n4313_1) );
  AND2X2 AND2X2_974 ( .A(AES_CORE_DATAPATH__abc_16259_n4317), .B(AES_CORE_DATAPATH__abc_16259_n2804_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n4318_1) );
  AND2X2 AND2X2_975 ( .A(AES_CORE_DATAPATH__abc_16259_n4318_1), .B(AES_CORE_DATAPATH__abc_16259_n4316), .Y(AES_CORE_DATAPATH__abc_16259_n4319_1) );
  AND2X2 AND2X2_976 ( .A(_auto_iopadmap_cc_313_execute_26949_14_), .B(AES_CORE_DATAPATH__abc_16259_n4322), .Y(AES_CORE_DATAPATH__abc_16259_n4323) );
  AND2X2 AND2X2_977 ( .A(AES_CORE_DATAPATH__abc_16259_n4324), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_6_), .Y(AES_CORE_DATAPATH__abc_16259_n4325) );
  AND2X2 AND2X2_978 ( .A(AES_CORE_DATAPATH__abc_16259_n4327_1), .B(AES_CORE_DATAPATH__abc_16259_n4321_1), .Y(AES_CORE_DATAPATH_sbox_pp2_14__FF_INPUT) );
  AND2X2 AND2X2_979 ( .A(_auto_iopadmap_cc_313_execute_26949_15_), .B(AES_CORE_DATAPATH__abc_16259_n4330), .Y(AES_CORE_DATAPATH__abc_16259_n4331) );
  AND2X2 AND2X2_98 ( .A(AES_CORE_DATAPATH__abc_16259_n2457_1), .B(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_1_), .Y(AES_CORE_DATAPATH__abc_16259_n2458) );
  AND2X2 AND2X2_980 ( .A(AES_CORE_DATAPATH__abc_16259_n4332), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_7_), .Y(AES_CORE_DATAPATH__abc_16259_n4333) );
  AND2X2 AND2X2_981 ( .A(AES_CORE_DATAPATH__abc_16259_n4335_1), .B(AES_CORE_DATAPATH__abc_16259_n4329_1), .Y(AES_CORE_DATAPATH_sbox_pp2_15__FF_INPUT) );
  AND2X2 AND2X2_982 ( .A(_auto_iopadmap_cc_313_execute_26949_16_), .B(AES_CORE_DATAPATH__abc_16259_n4338), .Y(AES_CORE_DATAPATH__abc_16259_n4339) );
  AND2X2 AND2X2_983 ( .A(AES_CORE_DATAPATH__abc_16259_n4340), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_1_2_), .Y(AES_CORE_DATAPATH__abc_16259_n4341) );
  AND2X2 AND2X2_984 ( .A(AES_CORE_DATAPATH__abc_16259_n4343_1), .B(AES_CORE_DATAPATH__abc_16259_n4337_1), .Y(AES_CORE_DATAPATH_sbox_pp2_16__FF_INPUT) );
  AND2X2 AND2X2_985 ( .A(_auto_iopadmap_cc_313_execute_26949_17_), .B(AES_CORE_DATAPATH__abc_16259_n4346), .Y(AES_CORE_DATAPATH__abc_16259_n4347) );
  AND2X2 AND2X2_986 ( .A(AES_CORE_DATAPATH__abc_16259_n4348), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_1_), .Y(AES_CORE_DATAPATH__abc_16259_n4349) );
  AND2X2 AND2X2_987 ( .A(AES_CORE_DATAPATH__abc_16259_n4351_1), .B(AES_CORE_DATAPATH__abc_16259_n4345_1), .Y(AES_CORE_DATAPATH_sbox_pp2_17__FF_INPUT) );
  AND2X2 AND2X2_988 ( .A(_auto_iopadmap_cc_313_execute_26949_18_), .B(AES_CORE_DATAPATH__abc_16259_n4354), .Y(AES_CORE_DATAPATH__abc_16259_n4355) );
  AND2X2 AND2X2_989 ( .A(AES_CORE_DATAPATH__abc_16259_n4356), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_2_), .Y(AES_CORE_DATAPATH__abc_16259_n4357) );
  AND2X2 AND2X2_99 ( .A(AES_CORE_CONTROL_UNIT_col_en_1_), .B(AES_CORE_CONTROL_UNIT_bypass_rk_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n2459_1) );
  AND2X2 AND2X2_990 ( .A(AES_CORE_DATAPATH__abc_16259_n4359_1), .B(AES_CORE_DATAPATH__abc_16259_n4353_1), .Y(AES_CORE_DATAPATH_sbox_pp2_18__FF_INPUT) );
  AND2X2 AND2X2_991 ( .A(_auto_iopadmap_cc_313_execute_26949_19_), .B(AES_CORE_DATAPATH__abc_16259_n4362), .Y(AES_CORE_DATAPATH__abc_16259_n4363) );
  AND2X2 AND2X2_992 ( .A(AES_CORE_DATAPATH__abc_16259_n4364), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_3_), .Y(AES_CORE_DATAPATH__abc_16259_n4365) );
  AND2X2 AND2X2_993 ( .A(AES_CORE_DATAPATH__abc_16259_n4367_1), .B(AES_CORE_DATAPATH__abc_16259_n4361_1), .Y(AES_CORE_DATAPATH_sbox_pp2_19__FF_INPUT) );
  AND2X2 AND2X2_994 ( .A(_auto_iopadmap_cc_313_execute_26949_20_), .B(AES_CORE_DATAPATH__abc_16259_n4370), .Y(AES_CORE_DATAPATH__abc_16259_n4371) );
  AND2X2 AND2X2_995 ( .A(AES_CORE_DATAPATH__abc_16259_n4372), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_4_), .Y(AES_CORE_DATAPATH__abc_16259_n4373) );
  AND2X2 AND2X2_996 ( .A(AES_CORE_DATAPATH__abc_16259_n4375_1), .B(AES_CORE_DATAPATH__abc_16259_n4369_1), .Y(AES_CORE_DATAPATH_sbox_pp2_20__FF_INPUT) );
  AND2X2 AND2X2_997 ( .A(_auto_iopadmap_cc_313_execute_26949_21_), .B(AES_CORE_DATAPATH__abc_16259_n4378), .Y(AES_CORE_DATAPATH__abc_16259_n4379) );
  AND2X2 AND2X2_998 ( .A(AES_CORE_DATAPATH__abc_16259_n4380), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_5_), .Y(AES_CORE_DATAPATH__abc_16259_n4381) );
  AND2X2 AND2X2_999 ( .A(AES_CORE_DATAPATH__abc_16259_n4383_1), .B(AES_CORE_DATAPATH__abc_16259_n4377_1), .Y(AES_CORE_DATAPATH_sbox_pp2_21__FF_INPUT) );
  BUFX2 BUFX2_1 ( .A(rst_n), .Y(rst_n_hier0_bF_buf8) );
  BUFX2 BUFX2_10 ( .A(clk), .Y(clk_hier0_bF_buf8) );
  BUFX2 BUFX2_100 ( .A(rst_n_hier0_bF_buf2), .Y(rst_n_bF_buf44) );
  BUFX2 BUFX2_101 ( .A(rst_n_hier0_bF_buf1), .Y(rst_n_bF_buf43) );
  BUFX2 BUFX2_102 ( .A(rst_n_hier0_bF_buf0), .Y(rst_n_bF_buf42) );
  BUFX2 BUFX2_103 ( .A(rst_n_hier0_bF_buf8), .Y(rst_n_bF_buf41) );
  BUFX2 BUFX2_104 ( .A(rst_n_hier0_bF_buf7), .Y(rst_n_bF_buf40) );
  BUFX2 BUFX2_105 ( .A(rst_n_hier0_bF_buf6), .Y(rst_n_bF_buf39) );
  BUFX2 BUFX2_106 ( .A(rst_n_hier0_bF_buf5), .Y(rst_n_bF_buf38) );
  BUFX2 BUFX2_107 ( .A(rst_n_hier0_bF_buf4), .Y(rst_n_bF_buf37) );
  BUFX2 BUFX2_108 ( .A(rst_n_hier0_bF_buf3), .Y(rst_n_bF_buf36) );
  BUFX2 BUFX2_109 ( .A(rst_n_hier0_bF_buf2), .Y(rst_n_bF_buf35) );
  BUFX2 BUFX2_11 ( .A(clk), .Y(clk_hier0_bF_buf7) );
  BUFX2 BUFX2_110 ( .A(rst_n_hier0_bF_buf1), .Y(rst_n_bF_buf34) );
  BUFX2 BUFX2_111 ( .A(rst_n_hier0_bF_buf0), .Y(rst_n_bF_buf33) );
  BUFX2 BUFX2_112 ( .A(rst_n_hier0_bF_buf8), .Y(rst_n_bF_buf32) );
  BUFX2 BUFX2_113 ( .A(rst_n_hier0_bF_buf7), .Y(rst_n_bF_buf31) );
  BUFX2 BUFX2_114 ( .A(rst_n_hier0_bF_buf6), .Y(rst_n_bF_buf30) );
  BUFX2 BUFX2_115 ( .A(rst_n_hier0_bF_buf5), .Y(rst_n_bF_buf29) );
  BUFX2 BUFX2_116 ( .A(rst_n_hier0_bF_buf4), .Y(rst_n_bF_buf28) );
  BUFX2 BUFX2_117 ( .A(rst_n_hier0_bF_buf3), .Y(rst_n_bF_buf27) );
  BUFX2 BUFX2_118 ( .A(rst_n_hier0_bF_buf2), .Y(rst_n_bF_buf26) );
  BUFX2 BUFX2_119 ( .A(rst_n_hier0_bF_buf1), .Y(rst_n_bF_buf25) );
  BUFX2 BUFX2_12 ( .A(clk), .Y(clk_hier0_bF_buf6) );
  BUFX2 BUFX2_120 ( .A(rst_n_hier0_bF_buf0), .Y(rst_n_bF_buf24) );
  BUFX2 BUFX2_121 ( .A(rst_n_hier0_bF_buf8), .Y(rst_n_bF_buf23) );
  BUFX2 BUFX2_122 ( .A(rst_n_hier0_bF_buf7), .Y(rst_n_bF_buf22) );
  BUFX2 BUFX2_123 ( .A(rst_n_hier0_bF_buf6), .Y(rst_n_bF_buf21) );
  BUFX2 BUFX2_124 ( .A(rst_n_hier0_bF_buf5), .Y(rst_n_bF_buf20) );
  BUFX2 BUFX2_125 ( .A(rst_n_hier0_bF_buf4), .Y(rst_n_bF_buf19) );
  BUFX2 BUFX2_126 ( .A(rst_n_hier0_bF_buf3), .Y(rst_n_bF_buf18) );
  BUFX2 BUFX2_127 ( .A(rst_n_hier0_bF_buf2), .Y(rst_n_bF_buf17) );
  BUFX2 BUFX2_128 ( .A(rst_n_hier0_bF_buf1), .Y(rst_n_bF_buf16) );
  BUFX2 BUFX2_129 ( .A(rst_n_hier0_bF_buf0), .Y(rst_n_bF_buf15) );
  BUFX2 BUFX2_13 ( .A(clk), .Y(clk_hier0_bF_buf5) );
  BUFX2 BUFX2_130 ( .A(rst_n_hier0_bF_buf8), .Y(rst_n_bF_buf14) );
  BUFX2 BUFX2_131 ( .A(rst_n_hier0_bF_buf7), .Y(rst_n_bF_buf13) );
  BUFX2 BUFX2_132 ( .A(rst_n_hier0_bF_buf6), .Y(rst_n_bF_buf12) );
  BUFX2 BUFX2_133 ( .A(rst_n_hier0_bF_buf5), .Y(rst_n_bF_buf11) );
  BUFX2 BUFX2_134 ( .A(rst_n_hier0_bF_buf4), .Y(rst_n_bF_buf10) );
  BUFX2 BUFX2_135 ( .A(rst_n_hier0_bF_buf3), .Y(rst_n_bF_buf9) );
  BUFX2 BUFX2_136 ( .A(rst_n_hier0_bF_buf2), .Y(rst_n_bF_buf8) );
  BUFX2 BUFX2_137 ( .A(rst_n_hier0_bF_buf1), .Y(rst_n_bF_buf7) );
  BUFX2 BUFX2_138 ( .A(rst_n_hier0_bF_buf0), .Y(rst_n_bF_buf6) );
  BUFX2 BUFX2_139 ( .A(rst_n_hier0_bF_buf8), .Y(rst_n_bF_buf5) );
  BUFX2 BUFX2_14 ( .A(clk), .Y(clk_hier0_bF_buf4) );
  BUFX2 BUFX2_140 ( .A(rst_n_hier0_bF_buf7), .Y(rst_n_bF_buf4) );
  BUFX2 BUFX2_141 ( .A(rst_n_hier0_bF_buf6), .Y(rst_n_bF_buf3) );
  BUFX2 BUFX2_142 ( .A(rst_n_hier0_bF_buf5), .Y(rst_n_bF_buf2) );
  BUFX2 BUFX2_143 ( .A(rst_n_hier0_bF_buf4), .Y(rst_n_bF_buf1) );
  BUFX2 BUFX2_144 ( .A(rst_n_hier0_bF_buf3), .Y(rst_n_bF_buf0) );
  BUFX2 BUFX2_145 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1), .Y(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf7) );
  BUFX2 BUFX2_146 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1), .Y(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf6) );
  BUFX2 BUFX2_147 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1), .Y(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf5) );
  BUFX2 BUFX2_148 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1), .Y(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf4) );
  BUFX2 BUFX2_149 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1), .Y(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf3) );
  BUFX2 BUFX2_15 ( .A(clk), .Y(clk_hier0_bF_buf3) );
  BUFX2 BUFX2_150 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1), .Y(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf2) );
  BUFX2 BUFX2_151 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1), .Y(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf1) );
  BUFX2 BUFX2_152 ( .A(AES_CORE_DATAPATH__abc_16259_n2469_1), .Y(AES_CORE_DATAPATH__abc_16259_n2469_1_bF_buf0) );
  BUFX2 BUFX2_153 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf5) );
  BUFX2 BUFX2_154 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf4) );
  BUFX2 BUFX2_155 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf3) );
  BUFX2 BUFX2_156 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf2) );
  BUFX2 BUFX2_157 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf1) );
  BUFX2 BUFX2_158 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf0) );
  BUFX2 BUFX2_159 ( .A(AES_CORE_DATAPATH__abc_16259_n5266_1), .Y(AES_CORE_DATAPATH__abc_16259_n5266_1_bF_buf4) );
  BUFX2 BUFX2_16 ( .A(clk), .Y(clk_hier0_bF_buf2) );
  BUFX2 BUFX2_160 ( .A(AES_CORE_DATAPATH__abc_16259_n5266_1), .Y(AES_CORE_DATAPATH__abc_16259_n5266_1_bF_buf3) );
  BUFX2 BUFX2_161 ( .A(AES_CORE_DATAPATH__abc_16259_n5266_1), .Y(AES_CORE_DATAPATH__abc_16259_n5266_1_bF_buf2) );
  BUFX2 BUFX2_162 ( .A(AES_CORE_DATAPATH__abc_16259_n5266_1), .Y(AES_CORE_DATAPATH__abc_16259_n5266_1_bF_buf1) );
  BUFX2 BUFX2_163 ( .A(AES_CORE_DATAPATH__abc_16259_n5266_1), .Y(AES_CORE_DATAPATH__abc_16259_n5266_1_bF_buf0) );
  BUFX2 BUFX2_164 ( .A(AES_CORE_DATAPATH__abc_16259_n8918), .Y(AES_CORE_DATAPATH__abc_16259_n8918_bF_buf4) );
  BUFX2 BUFX2_165 ( .A(AES_CORE_DATAPATH__abc_16259_n8918), .Y(AES_CORE_DATAPATH__abc_16259_n8918_bF_buf3) );
  BUFX2 BUFX2_166 ( .A(AES_CORE_DATAPATH__abc_16259_n8918), .Y(AES_CORE_DATAPATH__abc_16259_n8918_bF_buf2) );
  BUFX2 BUFX2_167 ( .A(AES_CORE_DATAPATH__abc_16259_n8918), .Y(AES_CORE_DATAPATH__abc_16259_n8918_bF_buf1) );
  BUFX2 BUFX2_168 ( .A(AES_CORE_DATAPATH__abc_16259_n8918), .Y(AES_CORE_DATAPATH__abc_16259_n8918_bF_buf0) );
  BUFX2 BUFX2_169 ( .A(AES_CORE_DATAPATH__abc_16259_n2802), .Y(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf12) );
  BUFX2 BUFX2_17 ( .A(clk), .Y(clk_hier0_bF_buf1) );
  BUFX2 BUFX2_170 ( .A(AES_CORE_DATAPATH__abc_16259_n2802), .Y(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf11) );
  BUFX2 BUFX2_171 ( .A(AES_CORE_DATAPATH__abc_16259_n2802), .Y(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf10) );
  BUFX2 BUFX2_172 ( .A(AES_CORE_DATAPATH__abc_16259_n2802), .Y(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf9) );
  BUFX2 BUFX2_173 ( .A(AES_CORE_DATAPATH__abc_16259_n2802), .Y(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf8) );
  BUFX2 BUFX2_174 ( .A(AES_CORE_DATAPATH__abc_16259_n2802), .Y(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf7) );
  BUFX2 BUFX2_175 ( .A(AES_CORE_DATAPATH__abc_16259_n2802), .Y(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf6) );
  BUFX2 BUFX2_176 ( .A(AES_CORE_DATAPATH__abc_16259_n2802), .Y(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf5) );
  BUFX2 BUFX2_177 ( .A(AES_CORE_DATAPATH__abc_16259_n2802), .Y(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf4) );
  BUFX2 BUFX2_178 ( .A(AES_CORE_DATAPATH__abc_16259_n2802), .Y(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf3) );
  BUFX2 BUFX2_179 ( .A(AES_CORE_DATAPATH__abc_16259_n2802), .Y(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf2) );
  BUFX2 BUFX2_18 ( .A(clk), .Y(clk_hier0_bF_buf0) );
  BUFX2 BUFX2_180 ( .A(AES_CORE_DATAPATH__abc_16259_n2802), .Y(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf1) );
  BUFX2 BUFX2_181 ( .A(AES_CORE_DATAPATH__abc_16259_n2802), .Y(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf0) );
  BUFX2 BUFX2_182 ( .A(AES_CORE_DATAPATH__abc_16259_n2803), .Y(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf10) );
  BUFX2 BUFX2_183 ( .A(AES_CORE_DATAPATH__abc_16259_n2803), .Y(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf9) );
  BUFX2 BUFX2_184 ( .A(AES_CORE_DATAPATH__abc_16259_n2803), .Y(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf8) );
  BUFX2 BUFX2_185 ( .A(AES_CORE_DATAPATH__abc_16259_n2803), .Y(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf7) );
  BUFX2 BUFX2_186 ( .A(AES_CORE_DATAPATH__abc_16259_n2803), .Y(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf6) );
  BUFX2 BUFX2_187 ( .A(AES_CORE_DATAPATH__abc_16259_n2803), .Y(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf5) );
  BUFX2 BUFX2_188 ( .A(AES_CORE_DATAPATH__abc_16259_n2803), .Y(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf4) );
  BUFX2 BUFX2_189 ( .A(AES_CORE_DATAPATH__abc_16259_n2803), .Y(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf3) );
  BUFX2 BUFX2_19 ( .A(AES_CORE_DATAPATH__abc_16259_n2887_1), .Y(AES_CORE_DATAPATH__abc_16259_n2887_1_bF_buf4) );
  BUFX2 BUFX2_190 ( .A(AES_CORE_DATAPATH__abc_16259_n2803), .Y(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf2) );
  BUFX2 BUFX2_191 ( .A(AES_CORE_DATAPATH__abc_16259_n2803), .Y(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf1) );
  BUFX2 BUFX2_192 ( .A(AES_CORE_DATAPATH__abc_16259_n2803), .Y(AES_CORE_DATAPATH__abc_16259_n2803_bF_buf0) );
  BUFX2 BUFX2_193 ( .A(AES_CORE_DATAPATH__abc_16259_n2807), .Y(AES_CORE_DATAPATH__abc_16259_n2807_bF_buf5) );
  BUFX2 BUFX2_194 ( .A(AES_CORE_DATAPATH__abc_16259_n2807), .Y(AES_CORE_DATAPATH__abc_16259_n2807_bF_buf4) );
  BUFX2 BUFX2_195 ( .A(AES_CORE_DATAPATH__abc_16259_n2807), .Y(AES_CORE_DATAPATH__abc_16259_n2807_bF_buf3) );
  BUFX2 BUFX2_196 ( .A(AES_CORE_DATAPATH__abc_16259_n2807), .Y(AES_CORE_DATAPATH__abc_16259_n2807_bF_buf2) );
  BUFX2 BUFX2_197 ( .A(AES_CORE_DATAPATH__abc_16259_n2807), .Y(AES_CORE_DATAPATH__abc_16259_n2807_bF_buf1) );
  BUFX2 BUFX2_198 ( .A(AES_CORE_DATAPATH__abc_16259_n2807), .Y(AES_CORE_DATAPATH__abc_16259_n2807_bF_buf0) );
  BUFX2 BUFX2_199 ( .A(AES_CORE_DATAPATH__abc_16259_n5653), .Y(AES_CORE_DATAPATH__abc_16259_n5653_bF_buf4) );
  BUFX2 BUFX2_2 ( .A(rst_n), .Y(rst_n_hier0_bF_buf7) );
  BUFX2 BUFX2_20 ( .A(AES_CORE_DATAPATH__abc_16259_n2887_1), .Y(AES_CORE_DATAPATH__abc_16259_n2887_1_bF_buf3) );
  BUFX2 BUFX2_200 ( .A(AES_CORE_DATAPATH__abc_16259_n5653), .Y(AES_CORE_DATAPATH__abc_16259_n5653_bF_buf3) );
  BUFX2 BUFX2_201 ( .A(AES_CORE_DATAPATH__abc_16259_n5653), .Y(AES_CORE_DATAPATH__abc_16259_n5653_bF_buf2) );
  BUFX2 BUFX2_202 ( .A(AES_CORE_DATAPATH__abc_16259_n5653), .Y(AES_CORE_DATAPATH__abc_16259_n5653_bF_buf1) );
  BUFX2 BUFX2_203 ( .A(AES_CORE_DATAPATH__abc_16259_n5653), .Y(AES_CORE_DATAPATH__abc_16259_n5653_bF_buf0) );
  BUFX2 BUFX2_204 ( .A(AES_CORE_DATAPATH__abc_16259_n5658), .Y(AES_CORE_DATAPATH__abc_16259_n5658_bF_buf4) );
  BUFX2 BUFX2_205 ( .A(AES_CORE_DATAPATH__abc_16259_n5658), .Y(AES_CORE_DATAPATH__abc_16259_n5658_bF_buf3) );
  BUFX2 BUFX2_206 ( .A(AES_CORE_DATAPATH__abc_16259_n5658), .Y(AES_CORE_DATAPATH__abc_16259_n5658_bF_buf2) );
  BUFX2 BUFX2_207 ( .A(AES_CORE_DATAPATH__abc_16259_n5658), .Y(AES_CORE_DATAPATH__abc_16259_n5658_bF_buf1) );
  BUFX2 BUFX2_208 ( .A(AES_CORE_DATAPATH__abc_16259_n5658), .Y(AES_CORE_DATAPATH__abc_16259_n5658_bF_buf0) );
  BUFX2 BUFX2_209 ( .A(AES_CORE_DATAPATH__abc_16259_n5659), .Y(AES_CORE_DATAPATH__abc_16259_n5659_bF_buf4) );
  BUFX2 BUFX2_21 ( .A(AES_CORE_DATAPATH__abc_16259_n2887_1), .Y(AES_CORE_DATAPATH__abc_16259_n2887_1_bF_buf2) );
  BUFX2 BUFX2_210 ( .A(AES_CORE_DATAPATH__abc_16259_n5659), .Y(AES_CORE_DATAPATH__abc_16259_n5659_bF_buf3) );
  BUFX2 BUFX2_211 ( .A(AES_CORE_DATAPATH__abc_16259_n5659), .Y(AES_CORE_DATAPATH__abc_16259_n5659_bF_buf2) );
  BUFX2 BUFX2_212 ( .A(AES_CORE_DATAPATH__abc_16259_n5659), .Y(AES_CORE_DATAPATH__abc_16259_n5659_bF_buf1) );
  BUFX2 BUFX2_213 ( .A(AES_CORE_DATAPATH__abc_16259_n5659), .Y(AES_CORE_DATAPATH__abc_16259_n5659_bF_buf0) );
  BUFX2 BUFX2_214 ( .A(AES_CORE_DATAPATH__abc_16259_n7944), .Y(AES_CORE_DATAPATH__abc_16259_n7944_bF_buf4) );
  BUFX2 BUFX2_215 ( .A(AES_CORE_DATAPATH__abc_16259_n7944), .Y(AES_CORE_DATAPATH__abc_16259_n7944_bF_buf3) );
  BUFX2 BUFX2_216 ( .A(AES_CORE_DATAPATH__abc_16259_n7944), .Y(AES_CORE_DATAPATH__abc_16259_n7944_bF_buf2) );
  BUFX2 BUFX2_217 ( .A(AES_CORE_DATAPATH__abc_16259_n7944), .Y(AES_CORE_DATAPATH__abc_16259_n7944_bF_buf1) );
  BUFX2 BUFX2_218 ( .A(AES_CORE_DATAPATH__abc_16259_n7944), .Y(AES_CORE_DATAPATH__abc_16259_n7944_bF_buf0) );
  BUFX2 BUFX2_219 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1_bF_buf4) );
  BUFX2 BUFX2_22 ( .A(AES_CORE_DATAPATH__abc_16259_n2887_1), .Y(AES_CORE_DATAPATH__abc_16259_n2887_1_bF_buf1) );
  BUFX2 BUFX2_220 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1_bF_buf3) );
  BUFX2 BUFX2_221 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1_bF_buf2) );
  BUFX2 BUFX2_222 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1_bF_buf1) );
  BUFX2 BUFX2_223 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n67_1_bF_buf0) );
  BUFX2 BUFX2_224 ( .A(AES_CORE_DATAPATH__abc_16259_n4867_1), .Y(AES_CORE_DATAPATH__abc_16259_n4867_1_bF_buf4) );
  BUFX2 BUFX2_225 ( .A(AES_CORE_DATAPATH__abc_16259_n4867_1), .Y(AES_CORE_DATAPATH__abc_16259_n4867_1_bF_buf3) );
  BUFX2 BUFX2_226 ( .A(AES_CORE_DATAPATH__abc_16259_n4867_1), .Y(AES_CORE_DATAPATH__abc_16259_n4867_1_bF_buf2) );
  BUFX2 BUFX2_227 ( .A(AES_CORE_DATAPATH__abc_16259_n4867_1), .Y(AES_CORE_DATAPATH__abc_16259_n4867_1_bF_buf1) );
  BUFX2 BUFX2_228 ( .A(AES_CORE_DATAPATH__abc_16259_n4867_1), .Y(AES_CORE_DATAPATH__abc_16259_n4867_1_bF_buf0) );
  BUFX2 BUFX2_229 ( .A(AES_CORE_DATAPATH__abc_16259_n2774), .Y(AES_CORE_DATAPATH__abc_16259_n2774_bF_buf4) );
  BUFX2 BUFX2_23 ( .A(AES_CORE_DATAPATH__abc_16259_n2887_1), .Y(AES_CORE_DATAPATH__abc_16259_n2887_1_bF_buf0) );
  BUFX2 BUFX2_230 ( .A(AES_CORE_DATAPATH__abc_16259_n2774), .Y(AES_CORE_DATAPATH__abc_16259_n2774_bF_buf3) );
  BUFX2 BUFX2_231 ( .A(AES_CORE_DATAPATH__abc_16259_n2774), .Y(AES_CORE_DATAPATH__abc_16259_n2774_bF_buf2) );
  BUFX2 BUFX2_232 ( .A(AES_CORE_DATAPATH__abc_16259_n2774), .Y(AES_CORE_DATAPATH__abc_16259_n2774_bF_buf1) );
  BUFX2 BUFX2_233 ( .A(AES_CORE_DATAPATH__abc_16259_n2774), .Y(AES_CORE_DATAPATH__abc_16259_n2774_bF_buf0) );
  BUFX2 BUFX2_234 ( .A(AES_CORE_DATAPATH__abc_16259_n2778), .Y(AES_CORE_DATAPATH__abc_16259_n2778_bF_buf4) );
  BUFX2 BUFX2_235 ( .A(AES_CORE_DATAPATH__abc_16259_n2778), .Y(AES_CORE_DATAPATH__abc_16259_n2778_bF_buf3) );
  BUFX2 BUFX2_236 ( .A(AES_CORE_DATAPATH__abc_16259_n2778), .Y(AES_CORE_DATAPATH__abc_16259_n2778_bF_buf2) );
  BUFX2 BUFX2_237 ( .A(AES_CORE_DATAPATH__abc_16259_n2778), .Y(AES_CORE_DATAPATH__abc_16259_n2778_bF_buf1) );
  BUFX2 BUFX2_238 ( .A(AES_CORE_DATAPATH__abc_16259_n2778), .Y(AES_CORE_DATAPATH__abc_16259_n2778_bF_buf0) );
  BUFX2 BUFX2_239 ( .A(AES_CORE_DATAPATH__abc_16259_n8500), .Y(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf6) );
  BUFX2 BUFX2_24 ( .A(AES_CORE_DATAPATH__abc_16259_n10217), .Y(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf7) );
  BUFX2 BUFX2_240 ( .A(AES_CORE_DATAPATH__abc_16259_n8500), .Y(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf5) );
  BUFX2 BUFX2_241 ( .A(AES_CORE_DATAPATH__abc_16259_n8500), .Y(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf4) );
  BUFX2 BUFX2_242 ( .A(AES_CORE_DATAPATH__abc_16259_n8500), .Y(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf3) );
  BUFX2 BUFX2_243 ( .A(AES_CORE_DATAPATH__abc_16259_n8500), .Y(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf2) );
  BUFX2 BUFX2_244 ( .A(AES_CORE_DATAPATH__abc_16259_n8500), .Y(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf1) );
  BUFX2 BUFX2_245 ( .A(AES_CORE_DATAPATH__abc_16259_n8500), .Y(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf0) );
  BUFX2 BUFX2_246 ( .A(AES_CORE_DATAPATH__abc_16259_n4474_1), .Y(AES_CORE_DATAPATH__abc_16259_n4474_1_bF_buf4) );
  BUFX2 BUFX2_247 ( .A(AES_CORE_DATAPATH__abc_16259_n4474_1), .Y(AES_CORE_DATAPATH__abc_16259_n4474_1_bF_buf3) );
  BUFX2 BUFX2_248 ( .A(AES_CORE_DATAPATH__abc_16259_n4474_1), .Y(AES_CORE_DATAPATH__abc_16259_n4474_1_bF_buf2) );
  BUFX2 BUFX2_249 ( .A(AES_CORE_DATAPATH__abc_16259_n4474_1), .Y(AES_CORE_DATAPATH__abc_16259_n4474_1_bF_buf1) );
  BUFX2 BUFX2_25 ( .A(AES_CORE_DATAPATH__abc_16259_n10217), .Y(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf6) );
  BUFX2 BUFX2_250 ( .A(AES_CORE_DATAPATH__abc_16259_n4474_1), .Y(AES_CORE_DATAPATH__abc_16259_n4474_1_bF_buf0) );
  BUFX2 BUFX2_251 ( .A(\iv_en[0] ), .Y(iv_en_0_bF_buf4) );
  BUFX2 BUFX2_252 ( .A(\iv_en[0] ), .Y(iv_en_0_bF_buf3) );
  BUFX2 BUFX2_253 ( .A(\iv_en[0] ), .Y(iv_en_0_bF_buf2) );
  BUFX2 BUFX2_254 ( .A(\iv_en[0] ), .Y(iv_en_0_bF_buf1) );
  BUFX2 BUFX2_255 ( .A(\iv_en[0] ), .Y(iv_en_0_bF_buf0) );
  BUFX2 BUFX2_256 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf92) );
  BUFX2 BUFX2_257 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf91) );
  BUFX2 BUFX2_258 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf90) );
  BUFX2 BUFX2_259 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf89) );
  BUFX2 BUFX2_26 ( .A(AES_CORE_DATAPATH__abc_16259_n10217), .Y(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf5) );
  BUFX2 BUFX2_260 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf88) );
  BUFX2 BUFX2_261 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf87) );
  BUFX2 BUFX2_262 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf86) );
  BUFX2 BUFX2_263 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf85) );
  BUFX2 BUFX2_264 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf84) );
  BUFX2 BUFX2_265 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf83) );
  BUFX2 BUFX2_266 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf82) );
  BUFX2 BUFX2_267 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf81) );
  BUFX2 BUFX2_268 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf80) );
  BUFX2 BUFX2_269 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf79) );
  BUFX2 BUFX2_27 ( .A(AES_CORE_DATAPATH__abc_16259_n10217), .Y(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf4) );
  BUFX2 BUFX2_270 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf78) );
  BUFX2 BUFX2_271 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf77) );
  BUFX2 BUFX2_272 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf76) );
  BUFX2 BUFX2_273 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf75) );
  BUFX2 BUFX2_274 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf74) );
  BUFX2 BUFX2_275 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf73) );
  BUFX2 BUFX2_276 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf72) );
  BUFX2 BUFX2_277 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf71) );
  BUFX2 BUFX2_278 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf70) );
  BUFX2 BUFX2_279 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf69) );
  BUFX2 BUFX2_28 ( .A(AES_CORE_DATAPATH__abc_16259_n10217), .Y(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf3) );
  BUFX2 BUFX2_280 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf68) );
  BUFX2 BUFX2_281 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf67) );
  BUFX2 BUFX2_282 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf66) );
  BUFX2 BUFX2_283 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf65) );
  BUFX2 BUFX2_284 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf64) );
  BUFX2 BUFX2_285 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf63) );
  BUFX2 BUFX2_286 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf62) );
  BUFX2 BUFX2_287 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf61) );
  BUFX2 BUFX2_288 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf60) );
  BUFX2 BUFX2_289 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf59) );
  BUFX2 BUFX2_29 ( .A(AES_CORE_DATAPATH__abc_16259_n10217), .Y(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf2) );
  BUFX2 BUFX2_290 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf58) );
  BUFX2 BUFX2_291 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf57) );
  BUFX2 BUFX2_292 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf56) );
  BUFX2 BUFX2_293 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf55) );
  BUFX2 BUFX2_294 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf54) );
  BUFX2 BUFX2_295 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf53) );
  BUFX2 BUFX2_296 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf52) );
  BUFX2 BUFX2_297 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf51) );
  BUFX2 BUFX2_298 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf50) );
  BUFX2 BUFX2_299 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf49) );
  BUFX2 BUFX2_3 ( .A(rst_n), .Y(rst_n_hier0_bF_buf6) );
  BUFX2 BUFX2_30 ( .A(AES_CORE_DATAPATH__abc_16259_n10217), .Y(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf1) );
  BUFX2 BUFX2_300 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf48) );
  BUFX2 BUFX2_301 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf47) );
  BUFX2 BUFX2_302 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf46) );
  BUFX2 BUFX2_303 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf45) );
  BUFX2 BUFX2_304 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf44) );
  BUFX2 BUFX2_305 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf43) );
  BUFX2 BUFX2_306 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf42) );
  BUFX2 BUFX2_307 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf41) );
  BUFX2 BUFX2_308 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf40) );
  BUFX2 BUFX2_309 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf39) );
  BUFX2 BUFX2_31 ( .A(AES_CORE_DATAPATH__abc_16259_n10217), .Y(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf0) );
  BUFX2 BUFX2_310 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf38) );
  BUFX2 BUFX2_311 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf37) );
  BUFX2 BUFX2_312 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf36) );
  BUFX2 BUFX2_313 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf35) );
  BUFX2 BUFX2_314 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf34) );
  BUFX2 BUFX2_315 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf33) );
  BUFX2 BUFX2_316 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf32) );
  BUFX2 BUFX2_317 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf31) );
  BUFX2 BUFX2_318 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf30) );
  BUFX2 BUFX2_319 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf29) );
  BUFX2 BUFX2_32 ( .A(AES_CORE_DATAPATH__abc_16259_n10218), .Y(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf6) );
  BUFX2 BUFX2_320 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf28) );
  BUFX2 BUFX2_321 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf27) );
  BUFX2 BUFX2_322 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf26) );
  BUFX2 BUFX2_323 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf25) );
  BUFX2 BUFX2_324 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf24) );
  BUFX2 BUFX2_325 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf23) );
  BUFX2 BUFX2_326 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf22) );
  BUFX2 BUFX2_327 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf21) );
  BUFX2 BUFX2_328 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf20) );
  BUFX2 BUFX2_329 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf19) );
  BUFX2 BUFX2_33 ( .A(AES_CORE_DATAPATH__abc_16259_n10218), .Y(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf5) );
  BUFX2 BUFX2_330 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf18) );
  BUFX2 BUFX2_331 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf17) );
  BUFX2 BUFX2_332 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf16) );
  BUFX2 BUFX2_333 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf15) );
  BUFX2 BUFX2_334 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf14) );
  BUFX2 BUFX2_335 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf13) );
  BUFX2 BUFX2_336 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf12) );
  BUFX2 BUFX2_337 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf11) );
  BUFX2 BUFX2_338 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf10) );
  BUFX2 BUFX2_339 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf9) );
  BUFX2 BUFX2_34 ( .A(AES_CORE_DATAPATH__abc_16259_n10218), .Y(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf4) );
  BUFX2 BUFX2_340 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf8) );
  BUFX2 BUFX2_341 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf7) );
  BUFX2 BUFX2_342 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf6) );
  BUFX2 BUFX2_343 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf5) );
  BUFX2 BUFX2_344 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf4) );
  BUFX2 BUFX2_345 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf3) );
  BUFX2 BUFX2_346 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf2) );
  BUFX2 BUFX2_347 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf1) );
  BUFX2 BUFX2_348 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf0) );
  BUFX2 BUFX2_349 ( .A(AES_CORE_DATAPATH__abc_16259_n2830_1), .Y(AES_CORE_DATAPATH__abc_16259_n2830_1_bF_buf4) );
  BUFX2 BUFX2_35 ( .A(AES_CORE_DATAPATH__abc_16259_n10218), .Y(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf3) );
  BUFX2 BUFX2_350 ( .A(AES_CORE_DATAPATH__abc_16259_n2830_1), .Y(AES_CORE_DATAPATH__abc_16259_n2830_1_bF_buf3) );
  BUFX2 BUFX2_351 ( .A(AES_CORE_DATAPATH__abc_16259_n2830_1), .Y(AES_CORE_DATAPATH__abc_16259_n2830_1_bF_buf2) );
  BUFX2 BUFX2_352 ( .A(AES_CORE_DATAPATH__abc_16259_n2830_1), .Y(AES_CORE_DATAPATH__abc_16259_n2830_1_bF_buf1) );
  BUFX2 BUFX2_353 ( .A(AES_CORE_DATAPATH__abc_16259_n2830_1), .Y(AES_CORE_DATAPATH__abc_16259_n2830_1_bF_buf0) );
  BUFX2 BUFX2_354 ( .A(AES_CORE_DATAPATH__abc_16259_n4872_1), .Y(AES_CORE_DATAPATH__abc_16259_n4872_1_bF_buf4) );
  BUFX2 BUFX2_355 ( .A(AES_CORE_DATAPATH__abc_16259_n4872_1), .Y(AES_CORE_DATAPATH__abc_16259_n4872_1_bF_buf3) );
  BUFX2 BUFX2_356 ( .A(AES_CORE_DATAPATH__abc_16259_n4872_1), .Y(AES_CORE_DATAPATH__abc_16259_n4872_1_bF_buf2) );
  BUFX2 BUFX2_357 ( .A(AES_CORE_DATAPATH__abc_16259_n4872_1), .Y(AES_CORE_DATAPATH__abc_16259_n4872_1_bF_buf1) );
  BUFX2 BUFX2_358 ( .A(AES_CORE_DATAPATH__abc_16259_n4872_1), .Y(AES_CORE_DATAPATH__abc_16259_n4872_1_bF_buf0) );
  BUFX2 BUFX2_359 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70_bF_buf4) );
  BUFX2 BUFX2_36 ( .A(AES_CORE_DATAPATH__abc_16259_n10218), .Y(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf2) );
  BUFX2 BUFX2_360 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70_bF_buf3) );
  BUFX2 BUFX2_361 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70_bF_buf2) );
  BUFX2 BUFX2_362 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70_bF_buf1) );
  BUFX2 BUFX2_363 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n70_bF_buf0) );
  BUFX2 BUFX2_364 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74_bF_buf4) );
  BUFX2 BUFX2_365 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74_bF_buf3) );
  BUFX2 BUFX2_366 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74_bF_buf2) );
  BUFX2 BUFX2_367 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74_bF_buf1) );
  BUFX2 BUFX2_368 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n74_bF_buf0) );
  BUFX2 BUFX2_369 ( .A(AES_CORE_DATAPATH__abc_16259_n6092), .Y(AES_CORE_DATAPATH__abc_16259_n6092_bF_buf4) );
  BUFX2 BUFX2_37 ( .A(AES_CORE_DATAPATH__abc_16259_n10218), .Y(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf1) );
  BUFX2 BUFX2_370 ( .A(AES_CORE_DATAPATH__abc_16259_n6092), .Y(AES_CORE_DATAPATH__abc_16259_n6092_bF_buf3) );
  BUFX2 BUFX2_371 ( .A(AES_CORE_DATAPATH__abc_16259_n6092), .Y(AES_CORE_DATAPATH__abc_16259_n6092_bF_buf2) );
  BUFX2 BUFX2_372 ( .A(AES_CORE_DATAPATH__abc_16259_n6092), .Y(AES_CORE_DATAPATH__abc_16259_n6092_bF_buf1) );
  BUFX2 BUFX2_373 ( .A(AES_CORE_DATAPATH__abc_16259_n6092), .Y(AES_CORE_DATAPATH__abc_16259_n6092_bF_buf0) );
  BUFX2 BUFX2_374 ( .A(AES_CORE_DATAPATH__abc_16259_n6095), .Y(AES_CORE_DATAPATH__abc_16259_n6095_bF_buf4) );
  BUFX2 BUFX2_375 ( .A(AES_CORE_DATAPATH__abc_16259_n6095), .Y(AES_CORE_DATAPATH__abc_16259_n6095_bF_buf3) );
  BUFX2 BUFX2_376 ( .A(AES_CORE_DATAPATH__abc_16259_n6095), .Y(AES_CORE_DATAPATH__abc_16259_n6095_bF_buf2) );
  BUFX2 BUFX2_377 ( .A(AES_CORE_DATAPATH__abc_16259_n6095), .Y(AES_CORE_DATAPATH__abc_16259_n6095_bF_buf1) );
  BUFX2 BUFX2_378 ( .A(AES_CORE_DATAPATH__abc_16259_n6095), .Y(AES_CORE_DATAPATH__abc_16259_n6095_bF_buf0) );
  BUFX2 BUFX2_379 ( .A(AES_CORE_DATAPATH__abc_16259_n6097), .Y(AES_CORE_DATAPATH__abc_16259_n6097_bF_buf4) );
  BUFX2 BUFX2_38 ( .A(AES_CORE_DATAPATH__abc_16259_n10218), .Y(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf0) );
  BUFX2 BUFX2_380 ( .A(AES_CORE_DATAPATH__abc_16259_n6097), .Y(AES_CORE_DATAPATH__abc_16259_n6097_bF_buf3) );
  BUFX2 BUFX2_381 ( .A(AES_CORE_DATAPATH__abc_16259_n6097), .Y(AES_CORE_DATAPATH__abc_16259_n6097_bF_buf2) );
  BUFX2 BUFX2_382 ( .A(AES_CORE_DATAPATH__abc_16259_n6097), .Y(AES_CORE_DATAPATH__abc_16259_n6097_bF_buf1) );
  BUFX2 BUFX2_383 ( .A(AES_CORE_DATAPATH__abc_16259_n6097), .Y(AES_CORE_DATAPATH__abc_16259_n6097_bF_buf0) );
  BUFX2 BUFX2_384 ( .A(AES_CORE_DATAPATH__abc_16259_n2837_1), .Y(AES_CORE_DATAPATH__abc_16259_n2837_1_bF_buf4) );
  BUFX2 BUFX2_385 ( .A(AES_CORE_DATAPATH__abc_16259_n2837_1), .Y(AES_CORE_DATAPATH__abc_16259_n2837_1_bF_buf3) );
  BUFX2 BUFX2_386 ( .A(AES_CORE_DATAPATH__abc_16259_n2837_1), .Y(AES_CORE_DATAPATH__abc_16259_n2837_1_bF_buf2) );
  BUFX2 BUFX2_387 ( .A(AES_CORE_DATAPATH__abc_16259_n2837_1), .Y(AES_CORE_DATAPATH__abc_16259_n2837_1_bF_buf1) );
  BUFX2 BUFX2_388 ( .A(AES_CORE_DATAPATH__abc_16259_n2837_1), .Y(AES_CORE_DATAPATH__abc_16259_n2837_1_bF_buf0) );
  BUFX2 BUFX2_389 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out_bF_buf4) );
  BUFX2 BUFX2_39 ( .A(AES_CORE_DATAPATH__abc_16259_n2482), .Y(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf5) );
  BUFX2 BUFX2_390 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out_bF_buf3) );
  BUFX2 BUFX2_391 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out_bF_buf2) );
  BUFX2 BUFX2_392 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out_bF_buf1) );
  BUFX2 BUFX2_393 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out_bF_buf0) );
  BUFX2 BUFX2_394 ( .A(AES_CORE_DATAPATH__abc_16259_n6063), .Y(AES_CORE_DATAPATH__abc_16259_n6063_bF_buf4) );
  BUFX2 BUFX2_395 ( .A(AES_CORE_DATAPATH__abc_16259_n6063), .Y(AES_CORE_DATAPATH__abc_16259_n6063_bF_buf3) );
  BUFX2 BUFX2_396 ( .A(AES_CORE_DATAPATH__abc_16259_n6063), .Y(AES_CORE_DATAPATH__abc_16259_n6063_bF_buf2) );
  BUFX2 BUFX2_397 ( .A(AES_CORE_DATAPATH__abc_16259_n6063), .Y(AES_CORE_DATAPATH__abc_16259_n6063_bF_buf1) );
  BUFX2 BUFX2_398 ( .A(AES_CORE_DATAPATH__abc_16259_n6063), .Y(AES_CORE_DATAPATH__abc_16259_n6063_bF_buf0) );
  BUFX2 BUFX2_399 ( .A(\key_en[1] ), .Y(key_en_1_bF_buf4) );
  BUFX2 BUFX2_4 ( .A(rst_n), .Y(rst_n_hier0_bF_buf5) );
  BUFX2 BUFX2_40 ( .A(AES_CORE_DATAPATH__abc_16259_n2482), .Y(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf4) );
  BUFX2 BUFX2_400 ( .A(\key_en[1] ), .Y(key_en_1_bF_buf3) );
  BUFX2 BUFX2_401 ( .A(\key_en[1] ), .Y(key_en_1_bF_buf2) );
  BUFX2 BUFX2_402 ( .A(\key_en[1] ), .Y(key_en_1_bF_buf1) );
  BUFX2 BUFX2_403 ( .A(\key_en[1] ), .Y(key_en_1_bF_buf0) );
  BUFX2 BUFX2_404 ( .A(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_CONTROL_UNIT_mode_cbc_bF_buf4) );
  BUFX2 BUFX2_405 ( .A(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_CONTROL_UNIT_mode_cbc_bF_buf3) );
  BUFX2 BUFX2_406 ( .A(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_CONTROL_UNIT_mode_cbc_bF_buf2) );
  BUFX2 BUFX2_407 ( .A(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_CONTROL_UNIT_mode_cbc_bF_buf1) );
  BUFX2 BUFX2_408 ( .A(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_CONTROL_UNIT_mode_cbc_bF_buf0) );
  BUFX2 BUFX2_409 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1_bF_buf4) );
  BUFX2 BUFX2_41 ( .A(AES_CORE_DATAPATH__abc_16259_n2482), .Y(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf3) );
  BUFX2 BUFX2_410 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1_bF_buf3) );
  BUFX2 BUFX2_411 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1_bF_buf2) );
  BUFX2 BUFX2_412 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1_bF_buf1) );
  BUFX2 BUFX2_413 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n76_1_bF_buf0) );
  BUFX2 BUFX2_414 ( .A(AES_CORE_DATAPATH__abc_16259_n10584), .Y(AES_CORE_DATAPATH__abc_16259_n10584_bF_buf4) );
  BUFX2 BUFX2_415 ( .A(AES_CORE_DATAPATH__abc_16259_n10584), .Y(AES_CORE_DATAPATH__abc_16259_n10584_bF_buf3) );
  BUFX2 BUFX2_416 ( .A(AES_CORE_DATAPATH__abc_16259_n10584), .Y(AES_CORE_DATAPATH__abc_16259_n10584_bF_buf2) );
  BUFX2 BUFX2_417 ( .A(AES_CORE_DATAPATH__abc_16259_n10584), .Y(AES_CORE_DATAPATH__abc_16259_n10584_bF_buf1) );
  BUFX2 BUFX2_418 ( .A(AES_CORE_DATAPATH__abc_16259_n10584), .Y(AES_CORE_DATAPATH__abc_16259_n10584_bF_buf0) );
  BUFX2 BUFX2_419 ( .A(AES_CORE_DATAPATH__abc_16259_n2864_1), .Y(AES_CORE_DATAPATH__abc_16259_n2864_1_bF_buf4) );
  BUFX2 BUFX2_42 ( .A(AES_CORE_DATAPATH__abc_16259_n2482), .Y(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf2) );
  BUFX2 BUFX2_420 ( .A(AES_CORE_DATAPATH__abc_16259_n2864_1), .Y(AES_CORE_DATAPATH__abc_16259_n2864_1_bF_buf3) );
  BUFX2 BUFX2_421 ( .A(AES_CORE_DATAPATH__abc_16259_n2864_1), .Y(AES_CORE_DATAPATH__abc_16259_n2864_1_bF_buf2) );
  BUFX2 BUFX2_422 ( .A(AES_CORE_DATAPATH__abc_16259_n2864_1), .Y(AES_CORE_DATAPATH__abc_16259_n2864_1_bF_buf1) );
  BUFX2 BUFX2_423 ( .A(AES_CORE_DATAPATH__abc_16259_n2864_1), .Y(AES_CORE_DATAPATH__abc_16259_n2864_1_bF_buf0) );
  BUFX2 BUFX2_424 ( .A(AES_CORE_DATAPATH__abc_16259_n2474), .Y(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf5) );
  BUFX2 BUFX2_425 ( .A(AES_CORE_DATAPATH__abc_16259_n2474), .Y(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf4) );
  BUFX2 BUFX2_426 ( .A(AES_CORE_DATAPATH__abc_16259_n2474), .Y(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf3) );
  BUFX2 BUFX2_427 ( .A(AES_CORE_DATAPATH__abc_16259_n2474), .Y(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf2) );
  BUFX2 BUFX2_428 ( .A(AES_CORE_DATAPATH__abc_16259_n2474), .Y(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf1) );
  BUFX2 BUFX2_429 ( .A(AES_CORE_DATAPATH__abc_16259_n2474), .Y(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf0) );
  BUFX2 BUFX2_43 ( .A(AES_CORE_DATAPATH__abc_16259_n2482), .Y(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf1) );
  BUFX2 BUFX2_430 ( .A(AES_CORE_DATAPATH__abc_16259_n4769), .Y(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf10) );
  BUFX2 BUFX2_431 ( .A(AES_CORE_DATAPATH__abc_16259_n4769), .Y(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf9) );
  BUFX2 BUFX2_432 ( .A(AES_CORE_DATAPATH__abc_16259_n4769), .Y(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf8) );
  BUFX2 BUFX2_433 ( .A(AES_CORE_DATAPATH__abc_16259_n4769), .Y(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf7) );
  BUFX2 BUFX2_434 ( .A(AES_CORE_DATAPATH__abc_16259_n4769), .Y(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf6) );
  BUFX2 BUFX2_435 ( .A(AES_CORE_DATAPATH__abc_16259_n4769), .Y(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf5) );
  BUFX2 BUFX2_436 ( .A(AES_CORE_DATAPATH__abc_16259_n4769), .Y(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf4) );
  BUFX2 BUFX2_437 ( .A(AES_CORE_DATAPATH__abc_16259_n4769), .Y(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf3) );
  BUFX2 BUFX2_438 ( .A(AES_CORE_DATAPATH__abc_16259_n4769), .Y(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf2) );
  BUFX2 BUFX2_439 ( .A(AES_CORE_DATAPATH__abc_16259_n4769), .Y(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf1) );
  BUFX2 BUFX2_44 ( .A(AES_CORE_DATAPATH__abc_16259_n2482), .Y(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf0) );
  BUFX2 BUFX2_440 ( .A(AES_CORE_DATAPATH__abc_16259_n4769), .Y(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf0) );
  BUFX2 BUFX2_441 ( .A(AES_CORE_DATAPATH__abc_16259_n2855), .Y(AES_CORE_DATAPATH__abc_16259_n2855_bF_buf4) );
  BUFX2 BUFX2_442 ( .A(AES_CORE_DATAPATH__abc_16259_n2855), .Y(AES_CORE_DATAPATH__abc_16259_n2855_bF_buf3) );
  BUFX2 BUFX2_443 ( .A(AES_CORE_DATAPATH__abc_16259_n2855), .Y(AES_CORE_DATAPATH__abc_16259_n2855_bF_buf2) );
  BUFX2 BUFX2_444 ( .A(AES_CORE_DATAPATH__abc_16259_n2855), .Y(AES_CORE_DATAPATH__abc_16259_n2855_bF_buf1) );
  BUFX2 BUFX2_445 ( .A(AES_CORE_DATAPATH__abc_16259_n2855), .Y(AES_CORE_DATAPATH__abc_16259_n2855_bF_buf0) );
  BUFX2 BUFX2_446 ( .A(AES_CORE_DATAPATH__abc_16259_n2857), .Y(AES_CORE_DATAPATH__abc_16259_n2857_bF_buf4) );
  BUFX2 BUFX2_447 ( .A(AES_CORE_DATAPATH__abc_16259_n2857), .Y(AES_CORE_DATAPATH__abc_16259_n2857_bF_buf3) );
  BUFX2 BUFX2_448 ( .A(AES_CORE_DATAPATH__abc_16259_n2857), .Y(AES_CORE_DATAPATH__abc_16259_n2857_bF_buf2) );
  BUFX2 BUFX2_449 ( .A(AES_CORE_DATAPATH__abc_16259_n2857), .Y(AES_CORE_DATAPATH__abc_16259_n2857_bF_buf1) );
  BUFX2 BUFX2_45 ( .A(AES_CORE_DATAPATH__abc_16259_n2484), .Y(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf7) );
  BUFX2 BUFX2_450 ( .A(AES_CORE_DATAPATH__abc_16259_n2857), .Y(AES_CORE_DATAPATH__abc_16259_n2857_bF_buf0) );
  BUFX2 BUFX2_451 ( .A(AES_CORE_DATAPATH__abc_16259_n2826), .Y(AES_CORE_DATAPATH__abc_16259_n2826_bF_buf4) );
  BUFX2 BUFX2_452 ( .A(AES_CORE_DATAPATH__abc_16259_n2826), .Y(AES_CORE_DATAPATH__abc_16259_n2826_bF_buf3) );
  BUFX2 BUFX2_453 ( .A(AES_CORE_DATAPATH__abc_16259_n2826), .Y(AES_CORE_DATAPATH__abc_16259_n2826_bF_buf2) );
  BUFX2 BUFX2_454 ( .A(AES_CORE_DATAPATH__abc_16259_n2826), .Y(AES_CORE_DATAPATH__abc_16259_n2826_bF_buf1) );
  BUFX2 BUFX2_455 ( .A(AES_CORE_DATAPATH__abc_16259_n2826), .Y(AES_CORE_DATAPATH__abc_16259_n2826_bF_buf0) );
  BUFX2 BUFX2_456 ( .A(AES_CORE_DATAPATH__abc_16259_n2796), .Y(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf7) );
  BUFX2 BUFX2_457 ( .A(AES_CORE_DATAPATH__abc_16259_n2796), .Y(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf6) );
  BUFX2 BUFX2_458 ( .A(AES_CORE_DATAPATH__abc_16259_n2796), .Y(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf5) );
  BUFX2 BUFX2_459 ( .A(AES_CORE_DATAPATH__abc_16259_n2796), .Y(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf4) );
  BUFX2 BUFX2_46 ( .A(AES_CORE_DATAPATH__abc_16259_n2484), .Y(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf6) );
  BUFX2 BUFX2_460 ( .A(AES_CORE_DATAPATH__abc_16259_n2796), .Y(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf3) );
  BUFX2 BUFX2_461 ( .A(AES_CORE_DATAPATH__abc_16259_n2796), .Y(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf2) );
  BUFX2 BUFX2_462 ( .A(AES_CORE_DATAPATH__abc_16259_n2796), .Y(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf1) );
  BUFX2 BUFX2_463 ( .A(AES_CORE_DATAPATH__abc_16259_n2796), .Y(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf0) );
  BUFX2 BUFX2_464 ( .A(AES_CORE_DATAPATH__abc_16259_n2798), .Y(AES_CORE_DATAPATH__abc_16259_n2798_bF_buf4) );
  BUFX2 BUFX2_465 ( .A(AES_CORE_DATAPATH__abc_16259_n2798), .Y(AES_CORE_DATAPATH__abc_16259_n2798_bF_buf3) );
  BUFX2 BUFX2_466 ( .A(AES_CORE_DATAPATH__abc_16259_n2798), .Y(AES_CORE_DATAPATH__abc_16259_n2798_bF_buf2) );
  BUFX2 BUFX2_467 ( .A(AES_CORE_DATAPATH__abc_16259_n2798), .Y(AES_CORE_DATAPATH__abc_16259_n2798_bF_buf1) );
  BUFX2 BUFX2_468 ( .A(AES_CORE_DATAPATH__abc_16259_n2798), .Y(AES_CORE_DATAPATH__abc_16259_n2798_bF_buf0) );
  BUFX2 BUFX2_469 ( .A(AES_CORE_DATAPATH__abc_16259_n2461_1), .Y(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf5) );
  BUFX2 BUFX2_47 ( .A(AES_CORE_DATAPATH__abc_16259_n2484), .Y(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf5) );
  BUFX2 BUFX2_470 ( .A(AES_CORE_DATAPATH__abc_16259_n2461_1), .Y(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf4) );
  BUFX2 BUFX2_471 ( .A(AES_CORE_DATAPATH__abc_16259_n2461_1), .Y(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf3) );
  BUFX2 BUFX2_472 ( .A(AES_CORE_DATAPATH__abc_16259_n2461_1), .Y(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf2) );
  BUFX2 BUFX2_473 ( .A(AES_CORE_DATAPATH__abc_16259_n2461_1), .Y(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf1) );
  BUFX2 BUFX2_474 ( .A(AES_CORE_DATAPATH__abc_16259_n2461_1), .Y(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf0) );
  BUFX2 BUFX2_475 ( .A(AES_CORE_DATAPATH__abc_16259_n8900), .Y(AES_CORE_DATAPATH__abc_16259_n8900_bF_buf3) );
  BUFX2 BUFX2_476 ( .A(AES_CORE_DATAPATH__abc_16259_n8900), .Y(AES_CORE_DATAPATH__abc_16259_n8900_bF_buf2) );
  BUFX2 BUFX2_477 ( .A(AES_CORE_DATAPATH__abc_16259_n8900), .Y(AES_CORE_DATAPATH__abc_16259_n8900_bF_buf1) );
  BUFX2 BUFX2_478 ( .A(AES_CORE_DATAPATH__abc_16259_n8900), .Y(AES_CORE_DATAPATH__abc_16259_n8900_bF_buf0) );
  BUFX2 BUFX2_479 ( .A(AES_CORE_DATAPATH__abc_16259_n8905), .Y(AES_CORE_DATAPATH__abc_16259_n8905_bF_buf4) );
  BUFX2 BUFX2_48 ( .A(AES_CORE_DATAPATH__abc_16259_n2484), .Y(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf4) );
  BUFX2 BUFX2_480 ( .A(AES_CORE_DATAPATH__abc_16259_n8905), .Y(AES_CORE_DATAPATH__abc_16259_n8905_bF_buf3) );
  BUFX2 BUFX2_481 ( .A(AES_CORE_DATAPATH__abc_16259_n8905), .Y(AES_CORE_DATAPATH__abc_16259_n8905_bF_buf2) );
  BUFX2 BUFX2_482 ( .A(AES_CORE_DATAPATH__abc_16259_n8905), .Y(AES_CORE_DATAPATH__abc_16259_n8905_bF_buf1) );
  BUFX2 BUFX2_483 ( .A(AES_CORE_DATAPATH__abc_16259_n8905), .Y(AES_CORE_DATAPATH__abc_16259_n8905_bF_buf0) );
  BUFX2 BUFX2_484 ( .A(AES_CORE_DATAPATH__abc_16259_n10119), .Y(AES_CORE_DATAPATH__abc_16259_n10119_bF_buf4) );
  BUFX2 BUFX2_485 ( .A(AES_CORE_DATAPATH__abc_16259_n10119), .Y(AES_CORE_DATAPATH__abc_16259_n10119_bF_buf3) );
  BUFX2 BUFX2_486 ( .A(AES_CORE_DATAPATH__abc_16259_n10119), .Y(AES_CORE_DATAPATH__abc_16259_n10119_bF_buf2) );
  BUFX2 BUFX2_487 ( .A(AES_CORE_DATAPATH__abc_16259_n10119), .Y(AES_CORE_DATAPATH__abc_16259_n10119_bF_buf1) );
  BUFX2 BUFX2_488 ( .A(AES_CORE_DATAPATH__abc_16259_n10119), .Y(AES_CORE_DATAPATH__abc_16259_n10119_bF_buf0) );
  BUFX2 BUFX2_489 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf7) );
  BUFX2 BUFX2_49 ( .A(AES_CORE_DATAPATH__abc_16259_n2484), .Y(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf3) );
  BUFX2 BUFX2_490 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf6) );
  BUFX2 BUFX2_491 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf5) );
  BUFX2 BUFX2_492 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf4) );
  BUFX2 BUFX2_493 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf3) );
  BUFX2 BUFX2_494 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf2) );
  BUFX2 BUFX2_495 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf1) );
  BUFX2 BUFX2_496 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf0) );
  BUFX2 BUFX2_497 ( .A(AES_CORE_DATAPATH__abc_16259_n8496), .Y(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf11) );
  BUFX2 BUFX2_498 ( .A(AES_CORE_DATAPATH__abc_16259_n8496), .Y(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf10) );
  BUFX2 BUFX2_499 ( .A(AES_CORE_DATAPATH__abc_16259_n8496), .Y(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf9) );
  BUFX2 BUFX2_5 ( .A(rst_n), .Y(rst_n_hier0_bF_buf4) );
  BUFX2 BUFX2_50 ( .A(AES_CORE_DATAPATH__abc_16259_n2484), .Y(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf2) );
  BUFX2 BUFX2_500 ( .A(AES_CORE_DATAPATH__abc_16259_n8496), .Y(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf8) );
  BUFX2 BUFX2_501 ( .A(AES_CORE_DATAPATH__abc_16259_n8496), .Y(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf7) );
  BUFX2 BUFX2_502 ( .A(AES_CORE_DATAPATH__abc_16259_n8496), .Y(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf6) );
  BUFX2 BUFX2_503 ( .A(AES_CORE_DATAPATH__abc_16259_n8496), .Y(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf5) );
  BUFX2 BUFX2_504 ( .A(AES_CORE_DATAPATH__abc_16259_n8496), .Y(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf4) );
  BUFX2 BUFX2_505 ( .A(AES_CORE_DATAPATH__abc_16259_n8496), .Y(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf3) );
  BUFX2 BUFX2_506 ( .A(AES_CORE_DATAPATH__abc_16259_n8496), .Y(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf2) );
  BUFX2 BUFX2_507 ( .A(AES_CORE_DATAPATH__abc_16259_n8496), .Y(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf1) );
  BUFX2 BUFX2_508 ( .A(AES_CORE_DATAPATH__abc_16259_n8496), .Y(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf0) );
  BUFX2 BUFX2_509 ( .A(AES_CORE_DATAPATH__abc_16259_n8499), .Y(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf7) );
  BUFX2 BUFX2_51 ( .A(AES_CORE_DATAPATH__abc_16259_n2484), .Y(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf1) );
  BUFX2 BUFX2_510 ( .A(AES_CORE_DATAPATH__abc_16259_n8499), .Y(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf6) );
  BUFX2 BUFX2_511 ( .A(AES_CORE_DATAPATH__abc_16259_n8499), .Y(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf5) );
  BUFX2 BUFX2_512 ( .A(AES_CORE_DATAPATH__abc_16259_n8499), .Y(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf4) );
  BUFX2 BUFX2_513 ( .A(AES_CORE_DATAPATH__abc_16259_n8499), .Y(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf3) );
  BUFX2 BUFX2_514 ( .A(AES_CORE_DATAPATH__abc_16259_n8499), .Y(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf2) );
  BUFX2 BUFX2_515 ( .A(AES_CORE_DATAPATH__abc_16259_n8499), .Y(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf1) );
  BUFX2 BUFX2_516 ( .A(AES_CORE_DATAPATH__abc_16259_n8499), .Y(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf0) );
  BUFX2 BUFX2_517 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1), .Y(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf10) );
  BUFX2 BUFX2_518 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1), .Y(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf9) );
  BUFX2 BUFX2_519 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1), .Y(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf8) );
  BUFX2 BUFX2_52 ( .A(AES_CORE_DATAPATH__abc_16259_n2484), .Y(AES_CORE_DATAPATH__abc_16259_n2484_bF_buf0) );
  BUFX2 BUFX2_520 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1), .Y(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf7) );
  BUFX2 BUFX2_521 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1), .Y(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf6) );
  BUFX2 BUFX2_522 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1), .Y(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf5) );
  BUFX2 BUFX2_523 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1), .Y(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf4) );
  BUFX2 BUFX2_524 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1), .Y(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf3) );
  BUFX2 BUFX2_525 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1), .Y(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf2) );
  BUFX2 BUFX2_526 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1), .Y(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf1) );
  BUFX2 BUFX2_527 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1), .Y(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf0) );
  BUFX2 BUFX2_528 ( .A(\iv_en[2] ), .Y(iv_en_2_bF_buf4) );
  BUFX2 BUFX2_529 ( .A(\iv_en[2] ), .Y(iv_en_2_bF_buf3) );
  BUFX2 BUFX2_53 ( .A(AES_CORE_DATAPATH__abc_16259_n8219), .Y(AES_CORE_DATAPATH__abc_16259_n8219_bF_buf4) );
  BUFX2 BUFX2_530 ( .A(\iv_en[2] ), .Y(iv_en_2_bF_buf2) );
  BUFX2 BUFX2_531 ( .A(\iv_en[2] ), .Y(iv_en_2_bF_buf1) );
  BUFX2 BUFX2_532 ( .A(\iv_en[2] ), .Y(iv_en_2_bF_buf0) );
  BUFX2 BUFX2_533 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1_bF_buf4) );
  BUFX2 BUFX2_534 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1_bF_buf3) );
  BUFX2 BUFX2_535 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1_bF_buf2) );
  BUFX2 BUFX2_536 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1_bF_buf1) );
  BUFX2 BUFX2_537 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n76_1_bF_buf0) );
  BUFX2 BUFX2_538 ( .A(AES_CORE_DATAPATH__abc_16259_n4468_1), .Y(AES_CORE_DATAPATH__abc_16259_n4468_1_bF_buf4) );
  BUFX2 BUFX2_539 ( .A(AES_CORE_DATAPATH__abc_16259_n4468_1), .Y(AES_CORE_DATAPATH__abc_16259_n4468_1_bF_buf3) );
  BUFX2 BUFX2_54 ( .A(AES_CORE_DATAPATH__abc_16259_n8219), .Y(AES_CORE_DATAPATH__abc_16259_n8219_bF_buf3) );
  BUFX2 BUFX2_540 ( .A(AES_CORE_DATAPATH__abc_16259_n4468_1), .Y(AES_CORE_DATAPATH__abc_16259_n4468_1_bF_buf2) );
  BUFX2 BUFX2_541 ( .A(AES_CORE_DATAPATH__abc_16259_n4468_1), .Y(AES_CORE_DATAPATH__abc_16259_n4468_1_bF_buf1) );
  BUFX2 BUFX2_542 ( .A(AES_CORE_DATAPATH__abc_16259_n4468_1), .Y(AES_CORE_DATAPATH__abc_16259_n4468_1_bF_buf0) );
  BUFX2 BUFX2_543 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf14) );
  BUFX2 BUFX2_544 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf13) );
  BUFX2 BUFX2_545 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf12) );
  BUFX2 BUFX2_546 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf11) );
  BUFX2 BUFX2_547 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf10) );
  BUFX2 BUFX2_548 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf9) );
  BUFX2 BUFX2_549 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf8) );
  BUFX2 BUFX2_55 ( .A(AES_CORE_DATAPATH__abc_16259_n8219), .Y(AES_CORE_DATAPATH__abc_16259_n8219_bF_buf2) );
  BUFX2 BUFX2_550 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf7) );
  BUFX2 BUFX2_551 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf6) );
  BUFX2 BUFX2_552 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf5) );
  BUFX2 BUFX2_553 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf4) );
  BUFX2 BUFX2_554 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf3) );
  BUFX2 BUFX2_555 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf2) );
  BUFX2 BUFX2_556 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf1) );
  BUFX2 BUFX2_557 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf0) );
  BUFX2 BUFX2_558 ( .A(AES_CORE_DATAPATH__abc_16259_n5265_1), .Y(AES_CORE_DATAPATH__abc_16259_n5265_1_bF_buf4) );
  BUFX2 BUFX2_559 ( .A(AES_CORE_DATAPATH__abc_16259_n5265_1), .Y(AES_CORE_DATAPATH__abc_16259_n5265_1_bF_buf3) );
  BUFX2 BUFX2_56 ( .A(AES_CORE_DATAPATH__abc_16259_n8219), .Y(AES_CORE_DATAPATH__abc_16259_n8219_bF_buf1) );
  BUFX2 BUFX2_560 ( .A(AES_CORE_DATAPATH__abc_16259_n5265_1), .Y(AES_CORE_DATAPATH__abc_16259_n5265_1_bF_buf2) );
  BUFX2 BUFX2_561 ( .A(AES_CORE_DATAPATH__abc_16259_n5265_1), .Y(AES_CORE_DATAPATH__abc_16259_n5265_1_bF_buf1) );
  BUFX2 BUFX2_562 ( .A(AES_CORE_DATAPATH__abc_16259_n5265_1), .Y(AES_CORE_DATAPATH__abc_16259_n5265_1_bF_buf0) );
  BUFX2 BUFX2_563 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1), .Y(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf7) );
  BUFX2 BUFX2_564 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1), .Y(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf6) );
  BUFX2 BUFX2_565 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1), .Y(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf5) );
  BUFX2 BUFX2_566 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1), .Y(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf4) );
  BUFX2 BUFX2_567 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1), .Y(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf3) );
  BUFX2 BUFX2_568 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1), .Y(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf2) );
  BUFX2 BUFX2_569 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1), .Y(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf1) );
  BUFX2 BUFX2_57 ( .A(AES_CORE_DATAPATH__abc_16259_n8219), .Y(AES_CORE_DATAPATH__abc_16259_n8219_bF_buf0) );
  BUFX2 BUFX2_570 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1), .Y(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf0) );
  BUFX2 BUFX2_571 ( .A(AES_CORE_DATAPATH__abc_16259_n9752), .Y(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf7) );
  BUFX2 BUFX2_572 ( .A(AES_CORE_DATAPATH__abc_16259_n9752), .Y(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf6) );
  BUFX2 BUFX2_573 ( .A(AES_CORE_DATAPATH__abc_16259_n9752), .Y(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf5) );
  BUFX2 BUFX2_574 ( .A(AES_CORE_DATAPATH__abc_16259_n9752), .Y(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf4) );
  BUFX2 BUFX2_575 ( .A(AES_CORE_DATAPATH__abc_16259_n9752), .Y(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf3) );
  BUFX2 BUFX2_576 ( .A(AES_CORE_DATAPATH__abc_16259_n9752), .Y(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf2) );
  BUFX2 BUFX2_577 ( .A(AES_CORE_DATAPATH__abc_16259_n9752), .Y(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf1) );
  BUFX2 BUFX2_578 ( .A(AES_CORE_DATAPATH__abc_16259_n9752), .Y(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf0) );
  BUFX2 BUFX2_579 ( .A(AES_CORE_DATAPATH__abc_16259_n9753), .Y(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf6) );
  BUFX2 BUFX2_58 ( .A(rst_n_hier0_bF_buf8), .Y(rst_n_bF_buf86) );
  BUFX2 BUFX2_580 ( .A(AES_CORE_DATAPATH__abc_16259_n9753), .Y(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf5) );
  BUFX2 BUFX2_581 ( .A(AES_CORE_DATAPATH__abc_16259_n9753), .Y(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf4) );
  BUFX2 BUFX2_582 ( .A(AES_CORE_DATAPATH__abc_16259_n9753), .Y(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf3) );
  BUFX2 BUFX2_583 ( .A(AES_CORE_DATAPATH__abc_16259_n9753), .Y(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf2) );
  BUFX2 BUFX2_584 ( .A(AES_CORE_DATAPATH__abc_16259_n9753), .Y(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf1) );
  BUFX2 BUFX2_585 ( .A(AES_CORE_DATAPATH__abc_16259_n9753), .Y(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf0) );
  BUFX2 BUFX2_586 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk), .Y(AES_CORE_CONTROL_UNIT_bypass_rk_bF_buf3) );
  BUFX2 BUFX2_587 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk), .Y(AES_CORE_CONTROL_UNIT_bypass_rk_bF_buf2) );
  BUFX2 BUFX2_588 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk), .Y(AES_CORE_CONTROL_UNIT_bypass_rk_bF_buf1) );
  BUFX2 BUFX2_589 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk), .Y(AES_CORE_CONTROL_UNIT_bypass_rk_bF_buf0) );
  BUFX2 BUFX2_59 ( .A(rst_n_hier0_bF_buf7), .Y(rst_n_bF_buf85) );
  BUFX2 BUFX2_590 ( .A(\key_en[3] ), .Y(key_en_3_bF_buf4) );
  BUFX2 BUFX2_591 ( .A(\key_en[3] ), .Y(key_en_3_bF_buf3) );
  BUFX2 BUFX2_592 ( .A(\key_en[3] ), .Y(key_en_3_bF_buf2) );
  BUFX2 BUFX2_593 ( .A(\key_en[3] ), .Y(key_en_3_bF_buf1) );
  BUFX2 BUFX2_594 ( .A(\key_en[3] ), .Y(key_en_3_bF_buf0) );
  BUFX2 BUFX2_595 ( .A(AES_CORE_DATAPATH__abc_16259_n6053), .Y(AES_CORE_DATAPATH__abc_16259_n6053_bF_buf4) );
  BUFX2 BUFX2_596 ( .A(AES_CORE_DATAPATH__abc_16259_n6053), .Y(AES_CORE_DATAPATH__abc_16259_n6053_bF_buf3) );
  BUFX2 BUFX2_597 ( .A(AES_CORE_DATAPATH__abc_16259_n6053), .Y(AES_CORE_DATAPATH__abc_16259_n6053_bF_buf2) );
  BUFX2 BUFX2_598 ( .A(AES_CORE_DATAPATH__abc_16259_n6053), .Y(AES_CORE_DATAPATH__abc_16259_n6053_bF_buf1) );
  BUFX2 BUFX2_599 ( .A(AES_CORE_DATAPATH__abc_16259_n6053), .Y(AES_CORE_DATAPATH__abc_16259_n6053_bF_buf0) );
  BUFX2 BUFX2_6 ( .A(rst_n), .Y(rst_n_hier0_bF_buf3) );
  BUFX2 BUFX2_60 ( .A(rst_n_hier0_bF_buf6), .Y(rst_n_bF_buf84) );
  BUFX2 BUFX2_600 ( .A(AES_CORE_DATAPATH__abc_16259_n6056), .Y(AES_CORE_DATAPATH__abc_16259_n6056_bF_buf4) );
  BUFX2 BUFX2_601 ( .A(AES_CORE_DATAPATH__abc_16259_n6056), .Y(AES_CORE_DATAPATH__abc_16259_n6056_bF_buf3) );
  BUFX2 BUFX2_602 ( .A(AES_CORE_DATAPATH__abc_16259_n6056), .Y(AES_CORE_DATAPATH__abc_16259_n6056_bF_buf2) );
  BUFX2 BUFX2_603 ( .A(AES_CORE_DATAPATH__abc_16259_n6056), .Y(AES_CORE_DATAPATH__abc_16259_n6056_bF_buf1) );
  BUFX2 BUFX2_604 ( .A(AES_CORE_DATAPATH__abc_16259_n6056), .Y(AES_CORE_DATAPATH__abc_16259_n6056_bF_buf0) );
  BUFX2 BUFX2_605 ( .A(AES_CORE_DATAPATH__abc_16259_n6057), .Y(AES_CORE_DATAPATH__abc_16259_n6057_bF_buf4) );
  BUFX2 BUFX2_606 ( .A(AES_CORE_DATAPATH__abc_16259_n6057), .Y(AES_CORE_DATAPATH__abc_16259_n6057_bF_buf3) );
  BUFX2 BUFX2_607 ( .A(AES_CORE_DATAPATH__abc_16259_n6057), .Y(AES_CORE_DATAPATH__abc_16259_n6057_bF_buf2) );
  BUFX2 BUFX2_608 ( .A(AES_CORE_DATAPATH__abc_16259_n6057), .Y(AES_CORE_DATAPATH__abc_16259_n6057_bF_buf1) );
  BUFX2 BUFX2_609 ( .A(AES_CORE_DATAPATH__abc_16259_n6057), .Y(AES_CORE_DATAPATH__abc_16259_n6057_bF_buf0) );
  BUFX2 BUFX2_61 ( .A(rst_n_hier0_bF_buf5), .Y(rst_n_bF_buf83) );
  BUFX2 BUFX2_610 ( .A(AES_CORE_DATAPATH__abc_16259_n6058), .Y(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf6) );
  BUFX2 BUFX2_611 ( .A(AES_CORE_DATAPATH__abc_16259_n6058), .Y(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf5) );
  BUFX2 BUFX2_612 ( .A(AES_CORE_DATAPATH__abc_16259_n6058), .Y(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf4) );
  BUFX2 BUFX2_613 ( .A(AES_CORE_DATAPATH__abc_16259_n6058), .Y(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf3) );
  BUFX2 BUFX2_614 ( .A(AES_CORE_DATAPATH__abc_16259_n6058), .Y(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf2) );
  BUFX2 BUFX2_615 ( .A(AES_CORE_DATAPATH__abc_16259_n6058), .Y(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf1) );
  BUFX2 BUFX2_616 ( .A(AES_CORE_DATAPATH__abc_16259_n6058), .Y(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf0) );
  BUFX2 BUFX2_617 ( .A(AES_CORE_DATAPATH__abc_16259_n6059), .Y(AES_CORE_DATAPATH__abc_16259_n6059_bF_buf5) );
  BUFX2 BUFX2_618 ( .A(AES_CORE_DATAPATH__abc_16259_n6059), .Y(AES_CORE_DATAPATH__abc_16259_n6059_bF_buf4) );
  BUFX2 BUFX2_619 ( .A(AES_CORE_DATAPATH__abc_16259_n6059), .Y(AES_CORE_DATAPATH__abc_16259_n6059_bF_buf3) );
  BUFX2 BUFX2_62 ( .A(rst_n_hier0_bF_buf4), .Y(rst_n_bF_buf82) );
  BUFX2 BUFX2_620 ( .A(AES_CORE_DATAPATH__abc_16259_n6059), .Y(AES_CORE_DATAPATH__abc_16259_n6059_bF_buf2) );
  BUFX2 BUFX2_621 ( .A(AES_CORE_DATAPATH__abc_16259_n6059), .Y(AES_CORE_DATAPATH__abc_16259_n6059_bF_buf1) );
  BUFX2 BUFX2_622 ( .A(AES_CORE_DATAPATH__abc_16259_n6059), .Y(AES_CORE_DATAPATH__abc_16259_n6059_bF_buf0) );
  BUFX2 BUFX2_623 ( .A(AES_CORE_DATAPATH__abc_16259_n9287), .Y(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf7) );
  BUFX2 BUFX2_624 ( .A(AES_CORE_DATAPATH__abc_16259_n9287), .Y(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf6) );
  BUFX2 BUFX2_625 ( .A(AES_CORE_DATAPATH__abc_16259_n9287), .Y(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf5) );
  BUFX2 BUFX2_626 ( .A(AES_CORE_DATAPATH__abc_16259_n9287), .Y(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf4) );
  BUFX2 BUFX2_627 ( .A(AES_CORE_DATAPATH__abc_16259_n9287), .Y(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf3) );
  BUFX2 BUFX2_628 ( .A(AES_CORE_DATAPATH__abc_16259_n9287), .Y(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf2) );
  BUFX2 BUFX2_629 ( .A(AES_CORE_DATAPATH__abc_16259_n9287), .Y(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf1) );
  BUFX2 BUFX2_63 ( .A(rst_n_hier0_bF_buf3), .Y(rst_n_bF_buf81) );
  BUFX2 BUFX2_630 ( .A(AES_CORE_DATAPATH__abc_16259_n9287), .Y(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf0) );
  BUFX2 BUFX2_631 ( .A(AES_CORE_DATAPATH__abc_16259_n9288), .Y(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf6) );
  BUFX2 BUFX2_632 ( .A(AES_CORE_DATAPATH__abc_16259_n9288), .Y(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf5) );
  BUFX2 BUFX2_633 ( .A(AES_CORE_DATAPATH__abc_16259_n9288), .Y(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf4) );
  BUFX2 BUFX2_634 ( .A(AES_CORE_DATAPATH__abc_16259_n9288), .Y(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf3) );
  BUFX2 BUFX2_635 ( .A(AES_CORE_DATAPATH__abc_16259_n9288), .Y(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf2) );
  BUFX2 BUFX2_636 ( .A(AES_CORE_DATAPATH__abc_16259_n9288), .Y(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf1) );
  BUFX2 BUFX2_637 ( .A(AES_CORE_DATAPATH__abc_16259_n9288), .Y(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf0) );
  BUFX2 BUFX2_638 ( .A(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf10) );
  BUFX2 BUFX2_639 ( .A(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf9) );
  BUFX2 BUFX2_64 ( .A(rst_n_hier0_bF_buf2), .Y(rst_n_bF_buf80) );
  BUFX2 BUFX2_640 ( .A(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf8) );
  BUFX2 BUFX2_641 ( .A(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf7) );
  BUFX2 BUFX2_642 ( .A(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf6) );
  BUFX2 BUFX2_643 ( .A(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf5) );
  BUFX2 BUFX2_644 ( .A(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf4) );
  BUFX2 BUFX2_645 ( .A(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf3) );
  BUFX2 BUFX2_646 ( .A(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf2) );
  BUFX2 BUFX2_647 ( .A(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf1) );
  BUFX2 BUFX2_648 ( .A(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf0) );
  BUFX2 BUFX2_649 ( .A(AES_CORE_DATAPATH__abc_16259_n2804_1), .Y(AES_CORE_DATAPATH__abc_16259_n2804_1_bF_buf4) );
  BUFX2 BUFX2_65 ( .A(rst_n_hier0_bF_buf1), .Y(rst_n_bF_buf79) );
  BUFX2 BUFX2_650 ( .A(AES_CORE_DATAPATH__abc_16259_n2804_1), .Y(AES_CORE_DATAPATH__abc_16259_n2804_1_bF_buf3) );
  BUFX2 BUFX2_651 ( .A(AES_CORE_DATAPATH__abc_16259_n2804_1), .Y(AES_CORE_DATAPATH__abc_16259_n2804_1_bF_buf2) );
  BUFX2 BUFX2_652 ( .A(AES_CORE_DATAPATH__abc_16259_n2804_1), .Y(AES_CORE_DATAPATH__abc_16259_n2804_1_bF_buf1) );
  BUFX2 BUFX2_653 ( .A(AES_CORE_DATAPATH__abc_16259_n2804_1), .Y(AES_CORE_DATAPATH__abc_16259_n2804_1_bF_buf0) );
  BUFX2 BUFX2_654 ( .A(AES_CORE_DATAPATH__abc_16259_n5260_1), .Y(AES_CORE_DATAPATH__abc_16259_n5260_1_bF_buf4) );
  BUFX2 BUFX2_655 ( .A(AES_CORE_DATAPATH__abc_16259_n5260_1), .Y(AES_CORE_DATAPATH__abc_16259_n5260_1_bF_buf3) );
  BUFX2 BUFX2_656 ( .A(AES_CORE_DATAPATH__abc_16259_n5260_1), .Y(AES_CORE_DATAPATH__abc_16259_n5260_1_bF_buf2) );
  BUFX2 BUFX2_657 ( .A(AES_CORE_DATAPATH__abc_16259_n5260_1), .Y(AES_CORE_DATAPATH__abc_16259_n5260_1_bF_buf1) );
  BUFX2 BUFX2_658 ( .A(AES_CORE_DATAPATH__abc_16259_n5260_1), .Y(AES_CORE_DATAPATH__abc_16259_n5260_1_bF_buf0) );
  BUFX2 BUFX2_659 ( .A(\key_en[0] ), .Y(key_en_0_bF_buf4) );
  BUFX2 BUFX2_66 ( .A(rst_n_hier0_bF_buf0), .Y(rst_n_bF_buf78) );
  BUFX2 BUFX2_660 ( .A(\key_en[0] ), .Y(key_en_0_bF_buf3) );
  BUFX2 BUFX2_661 ( .A(\key_en[0] ), .Y(key_en_0_bF_buf2) );
  BUFX2 BUFX2_662 ( .A(\key_en[0] ), .Y(key_en_0_bF_buf1) );
  BUFX2 BUFX2_663 ( .A(\key_en[0] ), .Y(key_en_0_bF_buf0) );
  BUFX2 BUFX2_664 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597_bF_buf4) );
  BUFX2 BUFX2_665 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597_bF_buf3) );
  BUFX2 BUFX2_666 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597_bF_buf2) );
  BUFX2 BUFX2_667 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597_bF_buf1) );
  BUFX2 BUFX2_668 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597_bF_buf0) );
  BUFX2 BUFX2_669 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1), .Y(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf7) );
  BUFX2 BUFX2_67 ( .A(rst_n_hier0_bF_buf8), .Y(rst_n_bF_buf77) );
  BUFX2 BUFX2_670 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1), .Y(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf6) );
  BUFX2 BUFX2_671 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1), .Y(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf5) );
  BUFX2 BUFX2_672 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1), .Y(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf4) );
  BUFX2 BUFX2_673 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1), .Y(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf3) );
  BUFX2 BUFX2_674 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1), .Y(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf2) );
  BUFX2 BUFX2_675 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1), .Y(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf1) );
  BUFX2 BUFX2_676 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1), .Y(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf0) );
  BUFX2 BUFX2_677 ( .A(AES_CORE_DATAPATH__abc_16259_n7669), .Y(AES_CORE_DATAPATH__abc_16259_n7669_bF_buf4) );
  BUFX2 BUFX2_678 ( .A(AES_CORE_DATAPATH__abc_16259_n7669), .Y(AES_CORE_DATAPATH__abc_16259_n7669_bF_buf3) );
  BUFX2 BUFX2_679 ( .A(AES_CORE_DATAPATH__abc_16259_n7669), .Y(AES_CORE_DATAPATH__abc_16259_n7669_bF_buf2) );
  BUFX2 BUFX2_68 ( .A(rst_n_hier0_bF_buf7), .Y(rst_n_bF_buf76) );
  BUFX2 BUFX2_680 ( .A(AES_CORE_DATAPATH__abc_16259_n7669), .Y(AES_CORE_DATAPATH__abc_16259_n7669_bF_buf1) );
  BUFX2 BUFX2_681 ( .A(AES_CORE_DATAPATH__abc_16259_n7669), .Y(AES_CORE_DATAPATH__abc_16259_n7669_bF_buf0) );
  BUFX2 BUFX2_682 ( .A(AES_CORE_DATAPATH__abc_16259_n8603), .Y(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf9) );
  BUFX2 BUFX2_683 ( .A(AES_CORE_DATAPATH__abc_16259_n8603), .Y(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf8) );
  BUFX2 BUFX2_684 ( .A(AES_CORE_DATAPATH__abc_16259_n8603), .Y(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf7) );
  BUFX2 BUFX2_685 ( .A(AES_CORE_DATAPATH__abc_16259_n8603), .Y(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf6) );
  BUFX2 BUFX2_686 ( .A(AES_CORE_DATAPATH__abc_16259_n8603), .Y(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf5) );
  BUFX2 BUFX2_687 ( .A(AES_CORE_DATAPATH__abc_16259_n8603), .Y(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf4) );
  BUFX2 BUFX2_688 ( .A(AES_CORE_DATAPATH__abc_16259_n8603), .Y(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf3) );
  BUFX2 BUFX2_689 ( .A(AES_CORE_DATAPATH__abc_16259_n8603), .Y(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf2) );
  BUFX2 BUFX2_69 ( .A(rst_n_hier0_bF_buf6), .Y(rst_n_bF_buf75) );
  BUFX2 BUFX2_690 ( .A(AES_CORE_DATAPATH__abc_16259_n8603), .Y(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf1) );
  BUFX2 BUFX2_691 ( .A(AES_CORE_DATAPATH__abc_16259_n8603), .Y(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf0) );
  BUFX2 BUFX2_692 ( .A(AES_CORE_DATAPATH__abc_16259_n2475_1), .Y(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf7) );
  BUFX2 BUFX2_693 ( .A(AES_CORE_DATAPATH__abc_16259_n2475_1), .Y(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf6) );
  BUFX2 BUFX2_694 ( .A(AES_CORE_DATAPATH__abc_16259_n2475_1), .Y(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf5) );
  BUFX2 BUFX2_695 ( .A(AES_CORE_DATAPATH__abc_16259_n2475_1), .Y(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf4) );
  BUFX2 BUFX2_696 ( .A(AES_CORE_DATAPATH__abc_16259_n2475_1), .Y(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf3) );
  BUFX2 BUFX2_697 ( .A(AES_CORE_DATAPATH__abc_16259_n2475_1), .Y(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf2) );
  BUFX2 BUFX2_698 ( .A(AES_CORE_DATAPATH__abc_16259_n2475_1), .Y(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf1) );
  BUFX2 BUFX2_699 ( .A(AES_CORE_DATAPATH__abc_16259_n2475_1), .Y(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf0) );
  BUFX2 BUFX2_7 ( .A(rst_n), .Y(rst_n_hier0_bF_buf2) );
  BUFX2 BUFX2_70 ( .A(rst_n_hier0_bF_buf5), .Y(rst_n_bF_buf74) );
  BUFX2 BUFX2_700 ( .A(AES_CORE_DATAPATH__abc_16259_n4475_1), .Y(AES_CORE_DATAPATH__abc_16259_n4475_1_bF_buf4) );
  BUFX2 BUFX2_701 ( .A(AES_CORE_DATAPATH__abc_16259_n4475_1), .Y(AES_CORE_DATAPATH__abc_16259_n4475_1_bF_buf3) );
  BUFX2 BUFX2_702 ( .A(AES_CORE_DATAPATH__abc_16259_n4475_1), .Y(AES_CORE_DATAPATH__abc_16259_n4475_1_bF_buf2) );
  BUFX2 BUFX2_703 ( .A(AES_CORE_DATAPATH__abc_16259_n4475_1), .Y(AES_CORE_DATAPATH__abc_16259_n4475_1_bF_buf1) );
  BUFX2 BUFX2_704 ( .A(AES_CORE_DATAPATH__abc_16259_n4475_1), .Y(AES_CORE_DATAPATH__abc_16259_n4475_1_bF_buf0) );
  BUFX2 BUFX2_705 ( .A(AES_CORE_DATAPATH__abc_16259_n2462), .Y(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf7) );
  BUFX2 BUFX2_706 ( .A(AES_CORE_DATAPATH__abc_16259_n2462), .Y(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf6) );
  BUFX2 BUFX2_707 ( .A(AES_CORE_DATAPATH__abc_16259_n2462), .Y(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf5) );
  BUFX2 BUFX2_708 ( .A(AES_CORE_DATAPATH__abc_16259_n2462), .Y(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf4) );
  BUFX2 BUFX2_709 ( .A(AES_CORE_DATAPATH__abc_16259_n2462), .Y(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf3) );
  BUFX2 BUFX2_71 ( .A(rst_n_hier0_bF_buf4), .Y(rst_n_bF_buf73) );
  BUFX2 BUFX2_710 ( .A(AES_CORE_DATAPATH__abc_16259_n2462), .Y(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf2) );
  BUFX2 BUFX2_711 ( .A(AES_CORE_DATAPATH__abc_16259_n2462), .Y(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf1) );
  BUFX2 BUFX2_712 ( .A(AES_CORE_DATAPATH__abc_16259_n2462), .Y(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf0) );
  BUFX2 BUFX2_713 ( .A(AES_CORE_DATAPATH__abc_16259_n2841), .Y(AES_CORE_DATAPATH__abc_16259_n2841_bF_buf4) );
  BUFX2 BUFX2_714 ( .A(AES_CORE_DATAPATH__abc_16259_n2841), .Y(AES_CORE_DATAPATH__abc_16259_n2841_bF_buf3) );
  BUFX2 BUFX2_715 ( .A(AES_CORE_DATAPATH__abc_16259_n2841), .Y(AES_CORE_DATAPATH__abc_16259_n2841_bF_buf2) );
  BUFX2 BUFX2_716 ( .A(AES_CORE_DATAPATH__abc_16259_n2841), .Y(AES_CORE_DATAPATH__abc_16259_n2841_bF_buf1) );
  BUFX2 BUFX2_717 ( .A(AES_CORE_DATAPATH__abc_16259_n2841), .Y(AES_CORE_DATAPATH__abc_16259_n2841_bF_buf0) );
  BUFX2 BUFX2_718 ( .A(AES_CORE_DATAPATH__abc_16259_n4873_1), .Y(AES_CORE_DATAPATH__abc_16259_n4873_1_bF_buf4) );
  BUFX2 BUFX2_719 ( .A(AES_CORE_DATAPATH__abc_16259_n4873_1), .Y(AES_CORE_DATAPATH__abc_16259_n4873_1_bF_buf3) );
  BUFX2 BUFX2_72 ( .A(rst_n_hier0_bF_buf3), .Y(rst_n_bF_buf72) );
  BUFX2 BUFX2_720 ( .A(AES_CORE_DATAPATH__abc_16259_n4873_1), .Y(AES_CORE_DATAPATH__abc_16259_n4873_1_bF_buf2) );
  BUFX2 BUFX2_721 ( .A(AES_CORE_DATAPATH__abc_16259_n4873_1), .Y(AES_CORE_DATAPATH__abc_16259_n4873_1_bF_buf1) );
  BUFX2 BUFX2_722 ( .A(AES_CORE_DATAPATH__abc_16259_n4873_1), .Y(AES_CORE_DATAPATH__abc_16259_n4873_1_bF_buf0) );
  BUFX2 BUFX2_723 ( .A(AES_CORE_DATAPATH__abc_16259_n8898), .Y(AES_CORE_DATAPATH__abc_16259_n8898_bF_buf4) );
  BUFX2 BUFX2_724 ( .A(AES_CORE_DATAPATH__abc_16259_n8898), .Y(AES_CORE_DATAPATH__abc_16259_n8898_bF_buf3) );
  BUFX2 BUFX2_725 ( .A(AES_CORE_DATAPATH__abc_16259_n8898), .Y(AES_CORE_DATAPATH__abc_16259_n8898_bF_buf2) );
  BUFX2 BUFX2_726 ( .A(AES_CORE_DATAPATH__abc_16259_n8898), .Y(AES_CORE_DATAPATH__abc_16259_n8898_bF_buf1) );
  BUFX2 BUFX2_727 ( .A(AES_CORE_DATAPATH__abc_16259_n8898), .Y(AES_CORE_DATAPATH__abc_16259_n8898_bF_buf0) );
  BUFX2 BUFX2_728 ( .A(AES_CORE_DATAPATH__abc_16259_n8899), .Y(AES_CORE_DATAPATH__abc_16259_n8899_bF_buf4) );
  BUFX2 BUFX2_729 ( .A(AES_CORE_DATAPATH__abc_16259_n8899), .Y(AES_CORE_DATAPATH__abc_16259_n8899_bF_buf3) );
  BUFX2 BUFX2_73 ( .A(rst_n_hier0_bF_buf2), .Y(rst_n_bF_buf71) );
  BUFX2 BUFX2_730 ( .A(AES_CORE_DATAPATH__abc_16259_n8899), .Y(AES_CORE_DATAPATH__abc_16259_n8899_bF_buf2) );
  BUFX2 BUFX2_731 ( .A(AES_CORE_DATAPATH__abc_16259_n8899), .Y(AES_CORE_DATAPATH__abc_16259_n8899_bF_buf1) );
  BUFX2 BUFX2_732 ( .A(AES_CORE_DATAPATH__abc_16259_n8899), .Y(AES_CORE_DATAPATH__abc_16259_n8899_bF_buf0) );
  BUFX2 BUFX2_733 ( .A(AES_CORE_DATAPATH__abc_16259_n2782), .Y(AES_CORE_DATAPATH__abc_16259_n2782_bF_buf4) );
  BUFX2 BUFX2_734 ( .A(AES_CORE_DATAPATH__abc_16259_n2782), .Y(AES_CORE_DATAPATH__abc_16259_n2782_bF_buf3) );
  BUFX2 BUFX2_735 ( .A(AES_CORE_DATAPATH__abc_16259_n2782), .Y(AES_CORE_DATAPATH__abc_16259_n2782_bF_buf2) );
  BUFX2 BUFX2_736 ( .A(AES_CORE_DATAPATH__abc_16259_n2782), .Y(AES_CORE_DATAPATH__abc_16259_n2782_bF_buf1) );
  BUFX2 BUFX2_737 ( .A(AES_CORE_DATAPATH__abc_16259_n2782), .Y(AES_CORE_DATAPATH__abc_16259_n2782_bF_buf0) );
  BUFX2 BUFX2_738 ( .A(AES_CORE_DATAPATH__abc_16259_n2786), .Y(AES_CORE_DATAPATH__abc_16259_n2786_bF_buf4) );
  BUFX2 BUFX2_739 ( .A(AES_CORE_DATAPATH__abc_16259_n2786), .Y(AES_CORE_DATAPATH__abc_16259_n2786_bF_buf3) );
  BUFX2 BUFX2_74 ( .A(rst_n_hier0_bF_buf1), .Y(rst_n_bF_buf70) );
  BUFX2 BUFX2_740 ( .A(AES_CORE_DATAPATH__abc_16259_n2786), .Y(AES_CORE_DATAPATH__abc_16259_n2786_bF_buf2) );
  BUFX2 BUFX2_741 ( .A(AES_CORE_DATAPATH__abc_16259_n2786), .Y(AES_CORE_DATAPATH__abc_16259_n2786_bF_buf1) );
  BUFX2 BUFX2_742 ( .A(AES_CORE_DATAPATH__abc_16259_n2786), .Y(AES_CORE_DATAPATH__abc_16259_n2786_bF_buf0) );
  BUFX2 BUFX2_743 ( .A(AES_CORE_DATAPATH__abc_16259_n2789), .Y(AES_CORE_DATAPATH__abc_16259_n2789_bF_buf4) );
  BUFX2 BUFX2_744 ( .A(AES_CORE_DATAPATH__abc_16259_n2789), .Y(AES_CORE_DATAPATH__abc_16259_n2789_bF_buf3) );
  BUFX2 BUFX2_745 ( .A(AES_CORE_DATAPATH__abc_16259_n2789), .Y(AES_CORE_DATAPATH__abc_16259_n2789_bF_buf2) );
  BUFX2 BUFX2_746 ( .A(AES_CORE_DATAPATH__abc_16259_n2789), .Y(AES_CORE_DATAPATH__abc_16259_n2789_bF_buf1) );
  BUFX2 BUFX2_747 ( .A(AES_CORE_DATAPATH__abc_16259_n2789), .Y(AES_CORE_DATAPATH__abc_16259_n2789_bF_buf0) );
  BUFX2 BUFX2_748 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1), .Y(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf10) );
  BUFX2 BUFX2_749 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1), .Y(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf9) );
  BUFX2 BUFX2_75 ( .A(rst_n_hier0_bF_buf0), .Y(rst_n_bF_buf69) );
  BUFX2 BUFX2_750 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1), .Y(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf8) );
  BUFX2 BUFX2_751 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1), .Y(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf7) );
  BUFX2 BUFX2_752 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1), .Y(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf6) );
  BUFX2 BUFX2_753 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1), .Y(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf5) );
  BUFX2 BUFX2_754 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1), .Y(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf4) );
  BUFX2 BUFX2_755 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1), .Y(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf3) );
  BUFX2 BUFX2_756 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1), .Y(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf2) );
  BUFX2 BUFX2_757 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1), .Y(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf1) );
  BUFX2 BUFX2_758 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1), .Y(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf0) );
  BUFX2 BUFX2_759 ( .A(AES_CORE_DATAPATH__abc_16259_n6603), .Y(AES_CORE_DATAPATH__abc_16259_n6603_bF_buf3) );
  BUFX2 BUFX2_76 ( .A(rst_n_hier0_bF_buf8), .Y(rst_n_bF_buf68) );
  BUFX2 BUFX2_760 ( .A(AES_CORE_DATAPATH__abc_16259_n6603), .Y(AES_CORE_DATAPATH__abc_16259_n6603_bF_buf2) );
  BUFX2 BUFX2_761 ( .A(AES_CORE_DATAPATH__abc_16259_n6603), .Y(AES_CORE_DATAPATH__abc_16259_n6603_bF_buf1) );
  BUFX2 BUFX2_762 ( .A(AES_CORE_DATAPATH__abc_16259_n6603), .Y(AES_CORE_DATAPATH__abc_16259_n6603_bF_buf0) );
  BUFX2 BUFX2_763 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70_bF_buf4) );
  BUFX2 BUFX2_764 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70_bF_buf3) );
  BUFX2 BUFX2_765 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70_bF_buf2) );
  BUFX2 BUFX2_766 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70_bF_buf1) );
  BUFX2 BUFX2_767 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n70_bF_buf0) );
  BUFX2 BUFX2_768 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74_bF_buf4) );
  BUFX2 BUFX2_769 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74_bF_buf3) );
  BUFX2 BUFX2_77 ( .A(rst_n_hier0_bF_buf7), .Y(rst_n_bF_buf67) );
  BUFX2 BUFX2_770 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74_bF_buf2) );
  BUFX2 BUFX2_771 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74_bF_buf1) );
  BUFX2 BUFX2_772 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n74_bF_buf0) );
  BUFX2 BUFX2_773 ( .A(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_CONTROL_UNIT_last_round_bF_buf5) );
  BUFX2 BUFX2_774 ( .A(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_CONTROL_UNIT_last_round_bF_buf4) );
  BUFX2 BUFX2_775 ( .A(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_CONTROL_UNIT_last_round_bF_buf3) );
  BUFX2 BUFX2_776 ( .A(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_CONTROL_UNIT_last_round_bF_buf2) );
  BUFX2 BUFX2_777 ( .A(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_CONTROL_UNIT_last_round_bF_buf1) );
  BUFX2 BUFX2_778 ( .A(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_CONTROL_UNIT_last_round_bF_buf0) );
  BUFX2 BUFX2_779 ( .A(\iv_en[1] ), .Y(iv_en_1_bF_buf4) );
  BUFX2 BUFX2_78 ( .A(rst_n_hier0_bF_buf6), .Y(rst_n_bF_buf66) );
  BUFX2 BUFX2_780 ( .A(\iv_en[1] ), .Y(iv_en_1_bF_buf3) );
  BUFX2 BUFX2_781 ( .A(\iv_en[1] ), .Y(iv_en_1_bF_buf2) );
  BUFX2 BUFX2_782 ( .A(\iv_en[1] ), .Y(iv_en_1_bF_buf1) );
  BUFX2 BUFX2_783 ( .A(\iv_en[1] ), .Y(iv_en_1_bF_buf0) );
  BUFX2 BUFX2_784 ( .A(AES_CORE_DATAPATH__abc_16259_n2853_1), .Y(AES_CORE_DATAPATH__abc_16259_n2853_1_bF_buf4) );
  BUFX2 BUFX2_785 ( .A(AES_CORE_DATAPATH__abc_16259_n2853_1), .Y(AES_CORE_DATAPATH__abc_16259_n2853_1_bF_buf3) );
  BUFX2 BUFX2_786 ( .A(AES_CORE_DATAPATH__abc_16259_n2853_1), .Y(AES_CORE_DATAPATH__abc_16259_n2853_1_bF_buf2) );
  BUFX2 BUFX2_787 ( .A(AES_CORE_DATAPATH__abc_16259_n2853_1), .Y(AES_CORE_DATAPATH__abc_16259_n2853_1_bF_buf1) );
  BUFX2 BUFX2_788 ( .A(AES_CORE_DATAPATH__abc_16259_n2853_1), .Y(AES_CORE_DATAPATH__abc_16259_n2853_1_bF_buf0) );
  BUFX2 BUFX2_789 ( .A(AES_CORE_DATAPATH__abc_16259_n6101), .Y(AES_CORE_DATAPATH__abc_16259_n6101_bF_buf4) );
  BUFX2 BUFX2_79 ( .A(rst_n_hier0_bF_buf5), .Y(rst_n_bF_buf65) );
  BUFX2 BUFX2_790 ( .A(AES_CORE_DATAPATH__abc_16259_n6101), .Y(AES_CORE_DATAPATH__abc_16259_n6101_bF_buf3) );
  BUFX2 BUFX2_791 ( .A(AES_CORE_DATAPATH__abc_16259_n6101), .Y(AES_CORE_DATAPATH__abc_16259_n6101_bF_buf2) );
  BUFX2 BUFX2_792 ( .A(AES_CORE_DATAPATH__abc_16259_n6101), .Y(AES_CORE_DATAPATH__abc_16259_n6101_bF_buf1) );
  BUFX2 BUFX2_793 ( .A(AES_CORE_DATAPATH__abc_16259_n6101), .Y(AES_CORE_DATAPATH__abc_16259_n6101_bF_buf0) );
  BUFX2 BUFX2_794 ( .A(AES_CORE_DATAPATH__abc_16259_n6107), .Y(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf9) );
  BUFX2 BUFX2_795 ( .A(AES_CORE_DATAPATH__abc_16259_n6107), .Y(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf8) );
  BUFX2 BUFX2_796 ( .A(AES_CORE_DATAPATH__abc_16259_n6107), .Y(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf7) );
  BUFX2 BUFX2_797 ( .A(AES_CORE_DATAPATH__abc_16259_n6107), .Y(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf6) );
  BUFX2 BUFX2_798 ( .A(AES_CORE_DATAPATH__abc_16259_n6107), .Y(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf5) );
  BUFX2 BUFX2_799 ( .A(AES_CORE_DATAPATH__abc_16259_n6107), .Y(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf4) );
  BUFX2 BUFX2_8 ( .A(rst_n), .Y(rst_n_hier0_bF_buf1) );
  BUFX2 BUFX2_80 ( .A(rst_n_hier0_bF_buf4), .Y(rst_n_bF_buf64) );
  BUFX2 BUFX2_800 ( .A(AES_CORE_DATAPATH__abc_16259_n6107), .Y(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf3) );
  BUFX2 BUFX2_801 ( .A(AES_CORE_DATAPATH__abc_16259_n6107), .Y(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf2) );
  BUFX2 BUFX2_802 ( .A(AES_CORE_DATAPATH__abc_16259_n6107), .Y(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf1) );
  BUFX2 BUFX2_803 ( .A(AES_CORE_DATAPATH__abc_16259_n6107), .Y(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf0) );
  BUFX2 BUFX2_804 ( .A(AES_CORE_DATAPATH_last_round_pp2), .Y(AES_CORE_DATAPATH_last_round_pp2_bF_buf4) );
  BUFX2 BUFX2_805 ( .A(AES_CORE_DATAPATH_last_round_pp2), .Y(AES_CORE_DATAPATH_last_round_pp2_bF_buf3) );
  BUFX2 BUFX2_806 ( .A(AES_CORE_DATAPATH_last_round_pp2), .Y(AES_CORE_DATAPATH_last_round_pp2_bF_buf2) );
  BUFX2 BUFX2_807 ( .A(AES_CORE_DATAPATH_last_round_pp2), .Y(AES_CORE_DATAPATH_last_round_pp2_bF_buf1) );
  BUFX2 BUFX2_808 ( .A(AES_CORE_DATAPATH_last_round_pp2), .Y(AES_CORE_DATAPATH_last_round_pp2_bF_buf0) );
  BUFX2 BUFX2_809 ( .A(AES_CORE_DATAPATH__abc_16259_n6074), .Y(AES_CORE_DATAPATH__abc_16259_n6074_bF_buf4) );
  BUFX2 BUFX2_81 ( .A(rst_n_hier0_bF_buf3), .Y(rst_n_bF_buf63) );
  BUFX2 BUFX2_810 ( .A(AES_CORE_DATAPATH__abc_16259_n6074), .Y(AES_CORE_DATAPATH__abc_16259_n6074_bF_buf3) );
  BUFX2 BUFX2_811 ( .A(AES_CORE_DATAPATH__abc_16259_n6074), .Y(AES_CORE_DATAPATH__abc_16259_n6074_bF_buf2) );
  BUFX2 BUFX2_812 ( .A(AES_CORE_DATAPATH__abc_16259_n6074), .Y(AES_CORE_DATAPATH__abc_16259_n6074_bF_buf1) );
  BUFX2 BUFX2_813 ( .A(AES_CORE_DATAPATH__abc_16259_n6074), .Y(AES_CORE_DATAPATH__abc_16259_n6074_bF_buf0) );
  BUFX2 BUFX2_814 ( .A(AES_CORE_DATAPATH__abc_16259_n2467_1), .Y(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf5) );
  BUFX2 BUFX2_815 ( .A(AES_CORE_DATAPATH__abc_16259_n2467_1), .Y(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf4) );
  BUFX2 BUFX2_816 ( .A(AES_CORE_DATAPATH__abc_16259_n2467_1), .Y(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf3) );
  BUFX2 BUFX2_817 ( .A(AES_CORE_DATAPATH__abc_16259_n2467_1), .Y(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf2) );
  BUFX2 BUFX2_818 ( .A(AES_CORE_DATAPATH__abc_16259_n2467_1), .Y(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf1) );
  BUFX2 BUFX2_819 ( .A(AES_CORE_DATAPATH__abc_16259_n2467_1), .Y(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf0) );
  BUFX2 BUFX2_82 ( .A(rst_n_hier0_bF_buf2), .Y(rst_n_bF_buf62) );
  BUFX2 BUFX2_820 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1_bF_buf4) );
  BUFX2 BUFX2_821 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1_bF_buf3) );
  BUFX2 BUFX2_822 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1_bF_buf2) );
  BUFX2 BUFX2_823 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1_bF_buf1) );
  BUFX2 BUFX2_824 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n67_1_bF_buf0) );
  BUFX2 BUFX2_825 ( .A(\key_en[2] ), .Y(key_en_2_bF_buf4) );
  BUFX2 BUFX2_826 ( .A(\key_en[2] ), .Y(key_en_2_bF_buf3) );
  BUFX2 BUFX2_827 ( .A(\key_en[2] ), .Y(key_en_2_bF_buf2) );
  BUFX2 BUFX2_828 ( .A(\key_en[2] ), .Y(key_en_2_bF_buf1) );
  BUFX2 BUFX2_829 ( .A(\key_en[2] ), .Y(key_en_2_bF_buf0) );
  BUFX2 BUFX2_83 ( .A(rst_n_hier0_bF_buf1), .Y(rst_n_bF_buf61) );
  BUFX2 BUFX2_830 ( .A(AES_CORE_DATAPATH__abc_16259_n6044), .Y(AES_CORE_DATAPATH__abc_16259_n6044_bF_buf4) );
  BUFX2 BUFX2_831 ( .A(AES_CORE_DATAPATH__abc_16259_n6044), .Y(AES_CORE_DATAPATH__abc_16259_n6044_bF_buf3) );
  BUFX2 BUFX2_832 ( .A(AES_CORE_DATAPATH__abc_16259_n6044), .Y(AES_CORE_DATAPATH__abc_16259_n6044_bF_buf2) );
  BUFX2 BUFX2_833 ( .A(AES_CORE_DATAPATH__abc_16259_n6044), .Y(AES_CORE_DATAPATH__abc_16259_n6044_bF_buf1) );
  BUFX2 BUFX2_834 ( .A(AES_CORE_DATAPATH__abc_16259_n6044), .Y(AES_CORE_DATAPATH__abc_16259_n6044_bF_buf0) );
  BUFX2 BUFX2_835 ( .A(AES_CORE_DATAPATH__abc_16259_n9654), .Y(AES_CORE_DATAPATH__abc_16259_n9654_bF_buf4) );
  BUFX2 BUFX2_836 ( .A(AES_CORE_DATAPATH__abc_16259_n9654), .Y(AES_CORE_DATAPATH__abc_16259_n9654_bF_buf3) );
  BUFX2 BUFX2_837 ( .A(AES_CORE_DATAPATH__abc_16259_n9654), .Y(AES_CORE_DATAPATH__abc_16259_n9654_bF_buf2) );
  BUFX2 BUFX2_838 ( .A(AES_CORE_DATAPATH__abc_16259_n9654), .Y(AES_CORE_DATAPATH__abc_16259_n9654_bF_buf1) );
  BUFX2 BUFX2_839 ( .A(AES_CORE_DATAPATH__abc_16259_n9654), .Y(AES_CORE_DATAPATH__abc_16259_n9654_bF_buf0) );
  BUFX2 BUFX2_84 ( .A(rst_n_hier0_bF_buf0), .Y(rst_n_bF_buf60) );
  BUFX2 BUFX2_840 ( .A(_auto_iopadmap_cc_313_execute_26881_0_), .Y(\col_out[0] ) );
  BUFX2 BUFX2_841 ( .A(_auto_iopadmap_cc_313_execute_26881_1_), .Y(\col_out[1] ) );
  BUFX2 BUFX2_842 ( .A(_auto_iopadmap_cc_313_execute_26881_2_), .Y(\col_out[2] ) );
  BUFX2 BUFX2_843 ( .A(_auto_iopadmap_cc_313_execute_26881_3_), .Y(\col_out[3] ) );
  BUFX2 BUFX2_844 ( .A(_auto_iopadmap_cc_313_execute_26881_4_), .Y(\col_out[4] ) );
  BUFX2 BUFX2_845 ( .A(_auto_iopadmap_cc_313_execute_26881_5_), .Y(\col_out[5] ) );
  BUFX2 BUFX2_846 ( .A(_auto_iopadmap_cc_313_execute_26881_6_), .Y(\col_out[6] ) );
  BUFX2 BUFX2_847 ( .A(_auto_iopadmap_cc_313_execute_26881_7_), .Y(\col_out[7] ) );
  BUFX2 BUFX2_848 ( .A(_auto_iopadmap_cc_313_execute_26881_8_), .Y(\col_out[8] ) );
  BUFX2 BUFX2_849 ( .A(_auto_iopadmap_cc_313_execute_26881_9_), .Y(\col_out[9] ) );
  BUFX2 BUFX2_85 ( .A(rst_n_hier0_bF_buf8), .Y(rst_n_bF_buf59) );
  BUFX2 BUFX2_850 ( .A(_auto_iopadmap_cc_313_execute_26881_10_), .Y(\col_out[10] ) );
  BUFX2 BUFX2_851 ( .A(_auto_iopadmap_cc_313_execute_26881_11_), .Y(\col_out[11] ) );
  BUFX2 BUFX2_852 ( .A(_auto_iopadmap_cc_313_execute_26881_12_), .Y(\col_out[12] ) );
  BUFX2 BUFX2_853 ( .A(_auto_iopadmap_cc_313_execute_26881_13_), .Y(\col_out[13] ) );
  BUFX2 BUFX2_854 ( .A(_auto_iopadmap_cc_313_execute_26881_14_), .Y(\col_out[14] ) );
  BUFX2 BUFX2_855 ( .A(_auto_iopadmap_cc_313_execute_26881_15_), .Y(\col_out[15] ) );
  BUFX2 BUFX2_856 ( .A(_auto_iopadmap_cc_313_execute_26881_16_), .Y(\col_out[16] ) );
  BUFX2 BUFX2_857 ( .A(_auto_iopadmap_cc_313_execute_26881_17_), .Y(\col_out[17] ) );
  BUFX2 BUFX2_858 ( .A(_auto_iopadmap_cc_313_execute_26881_18_), .Y(\col_out[18] ) );
  BUFX2 BUFX2_859 ( .A(_auto_iopadmap_cc_313_execute_26881_19_), .Y(\col_out[19] ) );
  BUFX2 BUFX2_86 ( .A(rst_n_hier0_bF_buf7), .Y(rst_n_bF_buf58) );
  BUFX2 BUFX2_860 ( .A(_auto_iopadmap_cc_313_execute_26881_20_), .Y(\col_out[20] ) );
  BUFX2 BUFX2_861 ( .A(_auto_iopadmap_cc_313_execute_26881_21_), .Y(\col_out[21] ) );
  BUFX2 BUFX2_862 ( .A(_auto_iopadmap_cc_313_execute_26881_22_), .Y(\col_out[22] ) );
  BUFX2 BUFX2_863 ( .A(_auto_iopadmap_cc_313_execute_26881_23_), .Y(\col_out[23] ) );
  BUFX2 BUFX2_864 ( .A(_auto_iopadmap_cc_313_execute_26881_24_), .Y(\col_out[24] ) );
  BUFX2 BUFX2_865 ( .A(_auto_iopadmap_cc_313_execute_26881_25_), .Y(\col_out[25] ) );
  BUFX2 BUFX2_866 ( .A(_auto_iopadmap_cc_313_execute_26881_26_), .Y(\col_out[26] ) );
  BUFX2 BUFX2_867 ( .A(_auto_iopadmap_cc_313_execute_26881_27_), .Y(\col_out[27] ) );
  BUFX2 BUFX2_868 ( .A(_auto_iopadmap_cc_313_execute_26881_28_), .Y(\col_out[28] ) );
  BUFX2 BUFX2_869 ( .A(_auto_iopadmap_cc_313_execute_26881_29_), .Y(\col_out[29] ) );
  BUFX2 BUFX2_87 ( .A(rst_n_hier0_bF_buf6), .Y(rst_n_bF_buf57) );
  BUFX2 BUFX2_870 ( .A(_auto_iopadmap_cc_313_execute_26881_30_), .Y(\col_out[30] ) );
  BUFX2 BUFX2_871 ( .A(_auto_iopadmap_cc_313_execute_26881_31_), .Y(\col_out[31] ) );
  BUFX2 BUFX2_872 ( .A(_auto_iopadmap_cc_313_execute_26914), .Y(end_aes) );
  BUFX2 BUFX2_873 ( .A(_auto_iopadmap_cc_313_execute_26916_0_), .Y(\iv_out[0] ) );
  BUFX2 BUFX2_874 ( .A(_auto_iopadmap_cc_313_execute_26916_1_), .Y(\iv_out[1] ) );
  BUFX2 BUFX2_875 ( .A(_auto_iopadmap_cc_313_execute_26916_2_), .Y(\iv_out[2] ) );
  BUFX2 BUFX2_876 ( .A(_auto_iopadmap_cc_313_execute_26916_3_), .Y(\iv_out[3] ) );
  BUFX2 BUFX2_877 ( .A(_auto_iopadmap_cc_313_execute_26916_4_), .Y(\iv_out[4] ) );
  BUFX2 BUFX2_878 ( .A(_auto_iopadmap_cc_313_execute_26916_5_), .Y(\iv_out[5] ) );
  BUFX2 BUFX2_879 ( .A(_auto_iopadmap_cc_313_execute_26916_6_), .Y(\iv_out[6] ) );
  BUFX2 BUFX2_88 ( .A(rst_n_hier0_bF_buf5), .Y(rst_n_bF_buf56) );
  BUFX2 BUFX2_880 ( .A(_auto_iopadmap_cc_313_execute_26916_7_), .Y(\iv_out[7] ) );
  BUFX2 BUFX2_881 ( .A(_auto_iopadmap_cc_313_execute_26916_8_), .Y(\iv_out[8] ) );
  BUFX2 BUFX2_882 ( .A(_auto_iopadmap_cc_313_execute_26916_9_), .Y(\iv_out[9] ) );
  BUFX2 BUFX2_883 ( .A(_auto_iopadmap_cc_313_execute_26916_10_), .Y(\iv_out[10] ) );
  BUFX2 BUFX2_884 ( .A(_auto_iopadmap_cc_313_execute_26916_11_), .Y(\iv_out[11] ) );
  BUFX2 BUFX2_885 ( .A(_auto_iopadmap_cc_313_execute_26916_12_), .Y(\iv_out[12] ) );
  BUFX2 BUFX2_886 ( .A(_auto_iopadmap_cc_313_execute_26916_13_), .Y(\iv_out[13] ) );
  BUFX2 BUFX2_887 ( .A(_auto_iopadmap_cc_313_execute_26916_14_), .Y(\iv_out[14] ) );
  BUFX2 BUFX2_888 ( .A(_auto_iopadmap_cc_313_execute_26916_15_), .Y(\iv_out[15] ) );
  BUFX2 BUFX2_889 ( .A(_auto_iopadmap_cc_313_execute_26916_16_), .Y(\iv_out[16] ) );
  BUFX2 BUFX2_89 ( .A(rst_n_hier0_bF_buf4), .Y(rst_n_bF_buf55) );
  BUFX2 BUFX2_890 ( .A(_auto_iopadmap_cc_313_execute_26916_17_), .Y(\iv_out[17] ) );
  BUFX2 BUFX2_891 ( .A(_auto_iopadmap_cc_313_execute_26916_18_), .Y(\iv_out[18] ) );
  BUFX2 BUFX2_892 ( .A(_auto_iopadmap_cc_313_execute_26916_19_), .Y(\iv_out[19] ) );
  BUFX2 BUFX2_893 ( .A(_auto_iopadmap_cc_313_execute_26916_20_), .Y(\iv_out[20] ) );
  BUFX2 BUFX2_894 ( .A(_auto_iopadmap_cc_313_execute_26916_21_), .Y(\iv_out[21] ) );
  BUFX2 BUFX2_895 ( .A(_auto_iopadmap_cc_313_execute_26916_22_), .Y(\iv_out[22] ) );
  BUFX2 BUFX2_896 ( .A(_auto_iopadmap_cc_313_execute_26916_23_), .Y(\iv_out[23] ) );
  BUFX2 BUFX2_897 ( .A(_auto_iopadmap_cc_313_execute_26916_24_), .Y(\iv_out[24] ) );
  BUFX2 BUFX2_898 ( .A(_auto_iopadmap_cc_313_execute_26916_25_), .Y(\iv_out[25] ) );
  BUFX2 BUFX2_899 ( .A(_auto_iopadmap_cc_313_execute_26916_26_), .Y(\iv_out[26] ) );
  BUFX2 BUFX2_9 ( .A(rst_n), .Y(rst_n_hier0_bF_buf0) );
  BUFX2 BUFX2_90 ( .A(rst_n_hier0_bF_buf3), .Y(rst_n_bF_buf54) );
  BUFX2 BUFX2_900 ( .A(_auto_iopadmap_cc_313_execute_26916_27_), .Y(\iv_out[27] ) );
  BUFX2 BUFX2_901 ( .A(_auto_iopadmap_cc_313_execute_26916_28_), .Y(\iv_out[28] ) );
  BUFX2 BUFX2_902 ( .A(_auto_iopadmap_cc_313_execute_26916_29_), .Y(\iv_out[29] ) );
  BUFX2 BUFX2_903 ( .A(_auto_iopadmap_cc_313_execute_26916_30_), .Y(\iv_out[30] ) );
  BUFX2 BUFX2_904 ( .A(_auto_iopadmap_cc_313_execute_26916_31_), .Y(\iv_out[31] ) );
  BUFX2 BUFX2_905 ( .A(_auto_iopadmap_cc_313_execute_26949_0_), .Y(\key_out[0] ) );
  BUFX2 BUFX2_906 ( .A(_auto_iopadmap_cc_313_execute_26949_1_), .Y(\key_out[1] ) );
  BUFX2 BUFX2_907 ( .A(_auto_iopadmap_cc_313_execute_26949_2_), .Y(\key_out[2] ) );
  BUFX2 BUFX2_908 ( .A(_auto_iopadmap_cc_313_execute_26949_3_), .Y(\key_out[3] ) );
  BUFX2 BUFX2_909 ( .A(_auto_iopadmap_cc_313_execute_26949_4_), .Y(\key_out[4] ) );
  BUFX2 BUFX2_91 ( .A(rst_n_hier0_bF_buf2), .Y(rst_n_bF_buf53) );
  BUFX2 BUFX2_910 ( .A(_auto_iopadmap_cc_313_execute_26949_5_), .Y(\key_out[5] ) );
  BUFX2 BUFX2_911 ( .A(_auto_iopadmap_cc_313_execute_26949_6_), .Y(\key_out[6] ) );
  BUFX2 BUFX2_912 ( .A(_auto_iopadmap_cc_313_execute_26949_7_), .Y(\key_out[7] ) );
  BUFX2 BUFX2_913 ( .A(_auto_iopadmap_cc_313_execute_26949_8_), .Y(\key_out[8] ) );
  BUFX2 BUFX2_914 ( .A(_auto_iopadmap_cc_313_execute_26949_9_), .Y(\key_out[9] ) );
  BUFX2 BUFX2_915 ( .A(_auto_iopadmap_cc_313_execute_26949_10_), .Y(\key_out[10] ) );
  BUFX2 BUFX2_916 ( .A(_auto_iopadmap_cc_313_execute_26949_11_), .Y(\key_out[11] ) );
  BUFX2 BUFX2_917 ( .A(_auto_iopadmap_cc_313_execute_26949_12_), .Y(\key_out[12] ) );
  BUFX2 BUFX2_918 ( .A(_auto_iopadmap_cc_313_execute_26949_13_), .Y(\key_out[13] ) );
  BUFX2 BUFX2_919 ( .A(_auto_iopadmap_cc_313_execute_26949_14_), .Y(\key_out[14] ) );
  BUFX2 BUFX2_92 ( .A(rst_n_hier0_bF_buf1), .Y(rst_n_bF_buf52) );
  BUFX2 BUFX2_920 ( .A(_auto_iopadmap_cc_313_execute_26949_15_), .Y(\key_out[15] ) );
  BUFX2 BUFX2_921 ( .A(_auto_iopadmap_cc_313_execute_26949_16_), .Y(\key_out[16] ) );
  BUFX2 BUFX2_922 ( .A(_auto_iopadmap_cc_313_execute_26949_17_), .Y(\key_out[17] ) );
  BUFX2 BUFX2_923 ( .A(_auto_iopadmap_cc_313_execute_26949_18_), .Y(\key_out[18] ) );
  BUFX2 BUFX2_924 ( .A(_auto_iopadmap_cc_313_execute_26949_19_), .Y(\key_out[19] ) );
  BUFX2 BUFX2_925 ( .A(_auto_iopadmap_cc_313_execute_26949_20_), .Y(\key_out[20] ) );
  BUFX2 BUFX2_926 ( .A(_auto_iopadmap_cc_313_execute_26949_21_), .Y(\key_out[21] ) );
  BUFX2 BUFX2_927 ( .A(_auto_iopadmap_cc_313_execute_26949_22_), .Y(\key_out[22] ) );
  BUFX2 BUFX2_928 ( .A(_auto_iopadmap_cc_313_execute_26949_23_), .Y(\key_out[23] ) );
  BUFX2 BUFX2_929 ( .A(_auto_iopadmap_cc_313_execute_26949_24_), .Y(\key_out[24] ) );
  BUFX2 BUFX2_93 ( .A(rst_n_hier0_bF_buf0), .Y(rst_n_bF_buf51) );
  BUFX2 BUFX2_930 ( .A(_auto_iopadmap_cc_313_execute_26949_25_), .Y(\key_out[25] ) );
  BUFX2 BUFX2_931 ( .A(_auto_iopadmap_cc_313_execute_26949_26_), .Y(\key_out[26] ) );
  BUFX2 BUFX2_932 ( .A(_auto_iopadmap_cc_313_execute_26949_27_), .Y(\key_out[27] ) );
  BUFX2 BUFX2_933 ( .A(_auto_iopadmap_cc_313_execute_26949_28_), .Y(\key_out[28] ) );
  BUFX2 BUFX2_934 ( .A(_auto_iopadmap_cc_313_execute_26949_29_), .Y(\key_out[29] ) );
  BUFX2 BUFX2_935 ( .A(_auto_iopadmap_cc_313_execute_26949_30_), .Y(\key_out[30] ) );
  BUFX2 BUFX2_936 ( .A(_auto_iopadmap_cc_313_execute_26949_31_), .Y(\key_out[31] ) );
  BUFX2 BUFX2_94 ( .A(rst_n_hier0_bF_buf8), .Y(rst_n_bF_buf50) );
  BUFX2 BUFX2_95 ( .A(rst_n_hier0_bF_buf7), .Y(rst_n_bF_buf49) );
  BUFX2 BUFX2_96 ( .A(rst_n_hier0_bF_buf6), .Y(rst_n_bF_buf48) );
  BUFX2 BUFX2_97 ( .A(rst_n_hier0_bF_buf5), .Y(rst_n_bF_buf47) );
  BUFX2 BUFX2_98 ( .A(rst_n_hier0_bF_buf4), .Y(rst_n_bF_buf46) );
  BUFX2 BUFX2_99 ( .A(rst_n_hier0_bF_buf3), .Y(rst_n_bF_buf45) );
  DFFPOSX1 DFFPOSX1_1 ( .CLK(clk_bF_buf72), .D(AES_CORE_DATAPATH_sbox_pp2_0__FF_INPUT), .Q(AES_CORE_DATAPATH_MIX_COL_col_0__0_) );
  DFFPOSX1 DFFPOSX1_10 ( .CLK(clk_bF_buf63), .D(AES_CORE_DATAPATH_sbox_pp2_9__FF_INPUT), .Q(AES_CORE_DATAPATH_MIX_COL_col_1__1_) );
  DFFPOSX1 DFFPOSX1_11 ( .CLK(clk_bF_buf62), .D(AES_CORE_DATAPATH_sbox_pp2_10__FF_INPUT), .Q(AES_CORE_DATAPATH_MIX_COL_col_1__2_) );
  DFFPOSX1 DFFPOSX1_12 ( .CLK(clk_bF_buf61), .D(AES_CORE_DATAPATH_sbox_pp2_11__FF_INPUT), .Q(AES_CORE_DATAPATH_MIX_COL_col_1__3_) );
  DFFPOSX1 DFFPOSX1_13 ( .CLK(clk_bF_buf60), .D(AES_CORE_DATAPATH_sbox_pp2_12__FF_INPUT), .Q(AES_CORE_DATAPATH_MIX_COL_col_1__4_) );
  DFFPOSX1 DFFPOSX1_14 ( .CLK(clk_bF_buf59), .D(AES_CORE_DATAPATH_sbox_pp2_13__FF_INPUT), .Q(AES_CORE_DATAPATH_MIX_COL_col_1__5_) );
  DFFPOSX1 DFFPOSX1_15 ( .CLK(clk_bF_buf58), .D(AES_CORE_DATAPATH_sbox_pp2_14__FF_INPUT), .Q(AES_CORE_DATAPATH_MIX_COL_col_1__6_) );
  DFFPOSX1 DFFPOSX1_16 ( .CLK(clk_bF_buf57), .D(AES_CORE_DATAPATH_sbox_pp2_15__FF_INPUT), .Q(AES_CORE_DATAPATH_MIX_COL_col_1__7_) );
  DFFPOSX1 DFFPOSX1_17 ( .CLK(clk_bF_buf56), .D(AES_CORE_DATAPATH_sbox_pp2_16__FF_INPUT), .Q(AES_CORE_DATAPATH_MIX_COL_col_2__0_) );
  DFFPOSX1 DFFPOSX1_18 ( .CLK(clk_bF_buf55), .D(AES_CORE_DATAPATH_sbox_pp2_17__FF_INPUT), .Q(AES_CORE_DATAPATH_MIX_COL_col_2__1_) );
  DFFPOSX1 DFFPOSX1_19 ( .CLK(clk_bF_buf54), .D(AES_CORE_DATAPATH_sbox_pp2_18__FF_INPUT), .Q(AES_CORE_DATAPATH_MIX_COL_col_2__2_) );
  DFFPOSX1 DFFPOSX1_2 ( .CLK(clk_bF_buf71), .D(AES_CORE_DATAPATH_sbox_pp2_1__FF_INPUT), .Q(AES_CORE_DATAPATH_MIX_COL_col_0__1_) );
  DFFPOSX1 DFFPOSX1_20 ( .CLK(clk_bF_buf53), .D(AES_CORE_DATAPATH_sbox_pp2_19__FF_INPUT), .Q(AES_CORE_DATAPATH_MIX_COL_col_2__3_) );
  DFFPOSX1 DFFPOSX1_21 ( .CLK(clk_bF_buf52), .D(AES_CORE_DATAPATH_sbox_pp2_20__FF_INPUT), .Q(AES_CORE_DATAPATH_MIX_COL_col_2__4_) );
  DFFPOSX1 DFFPOSX1_22 ( .CLK(clk_bF_buf51), .D(AES_CORE_DATAPATH_sbox_pp2_21__FF_INPUT), .Q(AES_CORE_DATAPATH_MIX_COL_col_2__5_) );
  DFFPOSX1 DFFPOSX1_23 ( .CLK(clk_bF_buf50), .D(AES_CORE_DATAPATH_sbox_pp2_22__FF_INPUT), .Q(AES_CORE_DATAPATH_MIX_COL_col_2__6_) );
  DFFPOSX1 DFFPOSX1_24 ( .CLK(clk_bF_buf49), .D(AES_CORE_DATAPATH_sbox_pp2_23__FF_INPUT), .Q(AES_CORE_DATAPATH_MIX_COL_col_2__7_) );
  DFFPOSX1 DFFPOSX1_25 ( .CLK(clk_bF_buf48), .D(AES_CORE_DATAPATH_sbox_pp2_24__FF_INPUT), .Q(AES_CORE_DATAPATH_MIX_COL_col_3__0_) );
  DFFPOSX1 DFFPOSX1_26 ( .CLK(clk_bF_buf47), .D(AES_CORE_DATAPATH_sbox_pp2_25__FF_INPUT), .Q(AES_CORE_DATAPATH_MIX_COL_col_3__1_) );
  DFFPOSX1 DFFPOSX1_27 ( .CLK(clk_bF_buf46), .D(AES_CORE_DATAPATH_sbox_pp2_26__FF_INPUT), .Q(AES_CORE_DATAPATH_MIX_COL_col_3__2_) );
  DFFPOSX1 DFFPOSX1_28 ( .CLK(clk_bF_buf45), .D(AES_CORE_DATAPATH_sbox_pp2_27__FF_INPUT), .Q(AES_CORE_DATAPATH_MIX_COL_col_3__3_) );
  DFFPOSX1 DFFPOSX1_29 ( .CLK(clk_bF_buf44), .D(AES_CORE_DATAPATH_sbox_pp2_28__FF_INPUT), .Q(AES_CORE_DATAPATH_MIX_COL_col_3__4_) );
  DFFPOSX1 DFFPOSX1_3 ( .CLK(clk_bF_buf70), .D(AES_CORE_DATAPATH_sbox_pp2_2__FF_INPUT), .Q(AES_CORE_DATAPATH_MIX_COL_col_0__2_) );
  DFFPOSX1 DFFPOSX1_30 ( .CLK(clk_bF_buf43), .D(AES_CORE_DATAPATH_sbox_pp2_29__FF_INPUT), .Q(AES_CORE_DATAPATH_MIX_COL_col_3__5_) );
  DFFPOSX1 DFFPOSX1_31 ( .CLK(clk_bF_buf42), .D(AES_CORE_DATAPATH_sbox_pp2_30__FF_INPUT), .Q(AES_CORE_DATAPATH_MIX_COL_col_3__6_) );
  DFFPOSX1 DFFPOSX1_32 ( .CLK(clk_bF_buf41), .D(AES_CORE_DATAPATH_sbox_pp2_31__FF_INPUT), .Q(AES_CORE_DATAPATH_MIX_COL_col_3__7_) );
  DFFPOSX1 DFFPOSX1_33 ( .CLK(clk_bF_buf76), .D(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_stage1_0_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_0_) );
  DFFPOSX1 DFFPOSX1_34 ( .CLK(clk_bF_buf75), .D(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_stage1_1_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_1_) );
  DFFPOSX1 DFFPOSX1_35 ( .CLK(clk_bF_buf74), .D(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_stage1_2_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_2_) );
  DFFPOSX1 DFFPOSX1_36 ( .CLK(clk_bF_buf73), .D(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_stage1_3_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_3_) );
  DFFPOSX1 DFFPOSX1_37 ( .CLK(clk_bF_buf72), .D(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_0_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_0_) );
  DFFPOSX1 DFFPOSX1_38 ( .CLK(clk_bF_buf71), .D(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_1_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_1_) );
  DFFPOSX1 DFFPOSX1_39 ( .CLK(clk_bF_buf70), .D(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_2_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_2_) );
  DFFPOSX1 DFFPOSX1_4 ( .CLK(clk_bF_buf69), .D(AES_CORE_DATAPATH_sbox_pp2_3__FF_INPUT), .Q(AES_CORE_DATAPATH_MIX_COL_col_0__3_) );
  DFFPOSX1 DFFPOSX1_40 ( .CLK(clk_bF_buf69), .D(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_3_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_3_) );
  DFFPOSX1 DFFPOSX1_41 ( .CLK(clk_bF_buf68), .D(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_4_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_4_) );
  DFFPOSX1 DFFPOSX1_42 ( .CLK(clk_bF_buf67), .D(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_5_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_5_) );
  DFFPOSX1 DFFPOSX1_43 ( .CLK(clk_bF_buf66), .D(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_6_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_6_) );
  DFFPOSX1 DFFPOSX1_44 ( .CLK(clk_bF_buf65), .D(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_7_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_7_) );
  DFFPOSX1 DFFPOSX1_45 ( .CLK(clk_bF_buf64), .D(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_stage1_0_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_0_) );
  DFFPOSX1 DFFPOSX1_46 ( .CLK(clk_bF_buf63), .D(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_stage1_1_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_1_) );
  DFFPOSX1 DFFPOSX1_47 ( .CLK(clk_bF_buf62), .D(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_stage1_2_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_2_) );
  DFFPOSX1 DFFPOSX1_48 ( .CLK(clk_bF_buf61), .D(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_stage1_3_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_3_) );
  DFFPOSX1 DFFPOSX1_49 ( .CLK(clk_bF_buf60), .D(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_0_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_0_) );
  DFFPOSX1 DFFPOSX1_5 ( .CLK(clk_bF_buf68), .D(AES_CORE_DATAPATH_sbox_pp2_4__FF_INPUT), .Q(AES_CORE_DATAPATH_MIX_COL_col_0__4_) );
  DFFPOSX1 DFFPOSX1_50 ( .CLK(clk_bF_buf59), .D(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_1_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_1_) );
  DFFPOSX1 DFFPOSX1_51 ( .CLK(clk_bF_buf58), .D(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_2_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_2_) );
  DFFPOSX1 DFFPOSX1_52 ( .CLK(clk_bF_buf57), .D(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_3_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_3_) );
  DFFPOSX1 DFFPOSX1_53 ( .CLK(clk_bF_buf56), .D(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_4_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_4_) );
  DFFPOSX1 DFFPOSX1_54 ( .CLK(clk_bF_buf55), .D(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_5_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_5_) );
  DFFPOSX1 DFFPOSX1_55 ( .CLK(clk_bF_buf54), .D(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_6_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_6_) );
  DFFPOSX1 DFFPOSX1_56 ( .CLK(clk_bF_buf53), .D(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_7_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_7_) );
  DFFPOSX1 DFFPOSX1_57 ( .CLK(clk_bF_buf52), .D(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_stage1_0_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_0_) );
  DFFPOSX1 DFFPOSX1_58 ( .CLK(clk_bF_buf51), .D(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_stage1_1_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_1_) );
  DFFPOSX1 DFFPOSX1_59 ( .CLK(clk_bF_buf50), .D(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_stage1_2_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_2_) );
  DFFPOSX1 DFFPOSX1_6 ( .CLK(clk_bF_buf67), .D(AES_CORE_DATAPATH_sbox_pp2_5__FF_INPUT), .Q(AES_CORE_DATAPATH_MIX_COL_col_0__5_) );
  DFFPOSX1 DFFPOSX1_60 ( .CLK(clk_bF_buf49), .D(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_stage1_3_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_3_) );
  DFFPOSX1 DFFPOSX1_61 ( .CLK(clk_bF_buf48), .D(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_0_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_0_) );
  DFFPOSX1 DFFPOSX1_62 ( .CLK(clk_bF_buf47), .D(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_1_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_1_) );
  DFFPOSX1 DFFPOSX1_63 ( .CLK(clk_bF_buf46), .D(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_2_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_2_) );
  DFFPOSX1 DFFPOSX1_64 ( .CLK(clk_bF_buf45), .D(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_3_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_3_) );
  DFFPOSX1 DFFPOSX1_65 ( .CLK(clk_bF_buf44), .D(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_4_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_4_) );
  DFFPOSX1 DFFPOSX1_66 ( .CLK(clk_bF_buf43), .D(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_5_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_5_) );
  DFFPOSX1 DFFPOSX1_67 ( .CLK(clk_bF_buf42), .D(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_6_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_6_) );
  DFFPOSX1 DFFPOSX1_68 ( .CLK(clk_bF_buf41), .D(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_7_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_7_) );
  DFFPOSX1 DFFPOSX1_69 ( .CLK(clk_bF_buf40), .D(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_stage1_0_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_0_) );
  DFFPOSX1 DFFPOSX1_7 ( .CLK(clk_bF_buf66), .D(AES_CORE_DATAPATH_sbox_pp2_6__FF_INPUT), .Q(AES_CORE_DATAPATH_MIX_COL_col_0__6_) );
  DFFPOSX1 DFFPOSX1_70 ( .CLK(clk_bF_buf39), .D(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_stage1_1_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_1_) );
  DFFPOSX1 DFFPOSX1_71 ( .CLK(clk_bF_buf38), .D(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_stage1_2_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_2_) );
  DFFPOSX1 DFFPOSX1_72 ( .CLK(clk_bF_buf37), .D(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_stage1_3_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_3_) );
  DFFPOSX1 DFFPOSX1_73 ( .CLK(clk_bF_buf36), .D(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_0_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_0_) );
  DFFPOSX1 DFFPOSX1_74 ( .CLK(clk_bF_buf35), .D(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_1_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_1_) );
  DFFPOSX1 DFFPOSX1_75 ( .CLK(clk_bF_buf34), .D(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_2_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_2_) );
  DFFPOSX1 DFFPOSX1_76 ( .CLK(clk_bF_buf33), .D(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_3_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_3_) );
  DFFPOSX1 DFFPOSX1_77 ( .CLK(clk_bF_buf32), .D(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_4_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_4_) );
  DFFPOSX1 DFFPOSX1_78 ( .CLK(clk_bF_buf31), .D(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_5_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_5_) );
  DFFPOSX1 DFFPOSX1_79 ( .CLK(clk_bF_buf30), .D(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_6_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_6_) );
  DFFPOSX1 DFFPOSX1_8 ( .CLK(clk_bF_buf65), .D(AES_CORE_DATAPATH_sbox_pp2_7__FF_INPUT), .Q(AES_CORE_DATAPATH_MIX_COL_col_0__7_) );
  DFFPOSX1 DFFPOSX1_80 ( .CLK(clk_bF_buf29), .D(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_7_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_7_) );
  DFFPOSX1 DFFPOSX1_9 ( .CLK(clk_bF_buf64), .D(AES_CORE_DATAPATH_sbox_pp2_8__FF_INPUT), .Q(AES_CORE_DATAPATH_MIX_COL_col_1__0_) );
  DFFSR DFFSR_1 ( .CLK(clk_bF_buf92), .D(AES_CORE_CONTROL_UNIT_rd_count_0__FF_INPUT), .Q(AES_CORE_CONTROL_UNIT_rd_count_0_), .R(rst_n_bF_buf86), .S(1'b1) );
  DFFSR DFFSR_10 ( .CLK(clk_bF_buf83), .D(AES_CORE_CONTROL_UNIT__abc_10818_n29), .Q(_auto_iopadmap_cc_313_execute_26914), .R(rst_n_bF_buf77), .S(1'b1) );
  DFFSR DFFSR_100 ( .CLK(clk_bF_buf54), .D(AES_CORE_DATAPATH__0key_host_1__31_0__15_), .Q(AES_CORE_DATAPATH_key_host_1__15_), .R(rst_n_bF_buf74), .S(1'b1) );
  DFFSR DFFSR_101 ( .CLK(clk_bF_buf53), .D(AES_CORE_DATAPATH__0key_host_1__31_0__16_), .Q(AES_CORE_DATAPATH_key_host_1__16_), .R(rst_n_bF_buf73), .S(1'b1) );
  DFFSR DFFSR_102 ( .CLK(clk_bF_buf52), .D(AES_CORE_DATAPATH__0key_host_1__31_0__17_), .Q(AES_CORE_DATAPATH_key_host_1__17_), .R(rst_n_bF_buf72), .S(1'b1) );
  DFFSR DFFSR_103 ( .CLK(clk_bF_buf51), .D(AES_CORE_DATAPATH__0key_host_1__31_0__18_), .Q(AES_CORE_DATAPATH_key_host_1__18_), .R(rst_n_bF_buf71), .S(1'b1) );
  DFFSR DFFSR_104 ( .CLK(clk_bF_buf50), .D(AES_CORE_DATAPATH__0key_host_1__31_0__19_), .Q(AES_CORE_DATAPATH_key_host_1__19_), .R(rst_n_bF_buf70), .S(1'b1) );
  DFFSR DFFSR_105 ( .CLK(clk_bF_buf49), .D(AES_CORE_DATAPATH__0key_host_1__31_0__20_), .Q(AES_CORE_DATAPATH_key_host_1__20_), .R(rst_n_bF_buf69), .S(1'b1) );
  DFFSR DFFSR_106 ( .CLK(clk_bF_buf48), .D(AES_CORE_DATAPATH__0key_host_1__31_0__21_), .Q(AES_CORE_DATAPATH_key_host_1__21_), .R(rst_n_bF_buf68), .S(1'b1) );
  DFFSR DFFSR_107 ( .CLK(clk_bF_buf47), .D(AES_CORE_DATAPATH__0key_host_1__31_0__22_), .Q(AES_CORE_DATAPATH_key_host_1__22_), .R(rst_n_bF_buf67), .S(1'b1) );
  DFFSR DFFSR_108 ( .CLK(clk_bF_buf46), .D(AES_CORE_DATAPATH__0key_host_1__31_0__23_), .Q(AES_CORE_DATAPATH_key_host_1__23_), .R(rst_n_bF_buf66), .S(1'b1) );
  DFFSR DFFSR_109 ( .CLK(clk_bF_buf45), .D(AES_CORE_DATAPATH__0key_host_1__31_0__24_), .Q(AES_CORE_DATAPATH_key_host_1__24_), .R(rst_n_bF_buf65), .S(1'b1) );
  DFFSR DFFSR_11 ( .CLK(clk_bF_buf82), .D(AES_CORE_CONTROL_UNIT__abc_10818_n12), .Q(AES_CORE_CONTROL_UNIT_state_6_), .R(rst_n_bF_buf76), .S(1'b1) );
  DFFSR DFFSR_110 ( .CLK(clk_bF_buf44), .D(AES_CORE_DATAPATH__0key_host_1__31_0__25_), .Q(AES_CORE_DATAPATH_key_host_1__25_), .R(rst_n_bF_buf64), .S(1'b1) );
  DFFSR DFFSR_111 ( .CLK(clk_bF_buf43), .D(AES_CORE_DATAPATH__0key_host_1__31_0__26_), .Q(AES_CORE_DATAPATH_key_host_1__26_), .R(rst_n_bF_buf63), .S(1'b1) );
  DFFSR DFFSR_112 ( .CLK(clk_bF_buf42), .D(AES_CORE_DATAPATH__0key_host_1__31_0__27_), .Q(AES_CORE_DATAPATH_key_host_1__27_), .R(rst_n_bF_buf62), .S(1'b1) );
  DFFSR DFFSR_113 ( .CLK(clk_bF_buf41), .D(AES_CORE_DATAPATH__0key_host_1__31_0__28_), .Q(AES_CORE_DATAPATH_key_host_1__28_), .R(rst_n_bF_buf61), .S(1'b1) );
  DFFSR DFFSR_114 ( .CLK(clk_bF_buf40), .D(AES_CORE_DATAPATH__0key_host_1__31_0__29_), .Q(AES_CORE_DATAPATH_key_host_1__29_), .R(rst_n_bF_buf60), .S(1'b1) );
  DFFSR DFFSR_115 ( .CLK(clk_bF_buf39), .D(AES_CORE_DATAPATH__0key_host_1__31_0__30_), .Q(AES_CORE_DATAPATH_key_host_1__30_), .R(rst_n_bF_buf59), .S(1'b1) );
  DFFSR DFFSR_116 ( .CLK(clk_bF_buf38), .D(AES_CORE_DATAPATH__0key_host_1__31_0__31_), .Q(AES_CORE_DATAPATH_key_host_1__31_), .R(rst_n_bF_buf58), .S(1'b1) );
  DFFSR DFFSR_117 ( .CLK(clk_bF_buf37), .D(AES_CORE_DATAPATH__0key_1__31_0__0_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__0_), .R(rst_n_bF_buf57), .S(1'b1) );
  DFFSR DFFSR_118 ( .CLK(clk_bF_buf36), .D(AES_CORE_DATAPATH__0key_1__31_0__1_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__1_), .R(rst_n_bF_buf56), .S(1'b1) );
  DFFSR DFFSR_119 ( .CLK(clk_bF_buf35), .D(AES_CORE_DATAPATH__0key_1__31_0__2_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__2_), .R(rst_n_bF_buf55), .S(1'b1) );
  DFFSR DFFSR_12 ( .CLK(clk_bF_buf81), .D(AES_CORE_CONTROL_UNIT__abc_10818_n303), .Q(AES_CORE_CONTROL_UNIT_state_7_), .R(rst_n_bF_buf75), .S(1'b1) );
  DFFSR DFFSR_120 ( .CLK(clk_bF_buf34), .D(AES_CORE_DATAPATH__0key_1__31_0__3_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__3_), .R(rst_n_bF_buf54), .S(1'b1) );
  DFFSR DFFSR_121 ( .CLK(clk_bF_buf33), .D(AES_CORE_DATAPATH__0key_1__31_0__4_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__4_), .R(rst_n_bF_buf53), .S(1'b1) );
  DFFSR DFFSR_122 ( .CLK(clk_bF_buf32), .D(AES_CORE_DATAPATH__0key_1__31_0__5_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__5_), .R(rst_n_bF_buf52), .S(1'b1) );
  DFFSR DFFSR_123 ( .CLK(clk_bF_buf31), .D(AES_CORE_DATAPATH__0key_1__31_0__6_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__6_), .R(rst_n_bF_buf51), .S(1'b1) );
  DFFSR DFFSR_124 ( .CLK(clk_bF_buf30), .D(AES_CORE_DATAPATH__0key_1__31_0__7_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__7_), .R(rst_n_bF_buf50), .S(1'b1) );
  DFFSR DFFSR_125 ( .CLK(clk_bF_buf29), .D(AES_CORE_DATAPATH__0key_1__31_0__8_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__8_), .R(rst_n_bF_buf49), .S(1'b1) );
  DFFSR DFFSR_126 ( .CLK(clk_bF_buf28), .D(AES_CORE_DATAPATH__0key_1__31_0__9_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__9_), .R(rst_n_bF_buf48), .S(1'b1) );
  DFFSR DFFSR_127 ( .CLK(clk_bF_buf27), .D(AES_CORE_DATAPATH__0key_1__31_0__10_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__10_), .R(rst_n_bF_buf47), .S(1'b1) );
  DFFSR DFFSR_128 ( .CLK(clk_bF_buf26), .D(AES_CORE_DATAPATH__0key_1__31_0__11_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__11_), .R(rst_n_bF_buf46), .S(1'b1) );
  DFFSR DFFSR_129 ( .CLK(clk_bF_buf25), .D(AES_CORE_DATAPATH__0key_1__31_0__12_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__12_), .R(rst_n_bF_buf45), .S(1'b1) );
  DFFSR DFFSR_13 ( .CLK(clk_bF_buf80), .D(AES_CORE_CONTROL_UNIT__abc_10818_n41), .Q(AES_CORE_CONTROL_UNIT_state_8_), .R(rst_n_bF_buf74), .S(1'b1) );
  DFFSR DFFSR_130 ( .CLK(clk_bF_buf24), .D(AES_CORE_DATAPATH__0key_1__31_0__13_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__13_), .R(rst_n_bF_buf44), .S(1'b1) );
  DFFSR DFFSR_131 ( .CLK(clk_bF_buf23), .D(AES_CORE_DATAPATH__0key_1__31_0__14_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__14_), .R(rst_n_bF_buf43), .S(1'b1) );
  DFFSR DFFSR_132 ( .CLK(clk_bF_buf22), .D(AES_CORE_DATAPATH__0key_1__31_0__15_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__15_), .R(rst_n_bF_buf42), .S(1'b1) );
  DFFSR DFFSR_133 ( .CLK(clk_bF_buf21), .D(AES_CORE_DATAPATH__0key_1__31_0__16_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__16_), .R(rst_n_bF_buf41), .S(1'b1) );
  DFFSR DFFSR_134 ( .CLK(clk_bF_buf20), .D(AES_CORE_DATAPATH__0key_1__31_0__17_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__17_), .R(rst_n_bF_buf40), .S(1'b1) );
  DFFSR DFFSR_135 ( .CLK(clk_bF_buf19), .D(AES_CORE_DATAPATH__0key_1__31_0__18_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__18_), .R(rst_n_bF_buf39), .S(1'b1) );
  DFFSR DFFSR_136 ( .CLK(clk_bF_buf18), .D(AES_CORE_DATAPATH__0key_1__31_0__19_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__19_), .R(rst_n_bF_buf38), .S(1'b1) );
  DFFSR DFFSR_137 ( .CLK(clk_bF_buf17), .D(AES_CORE_DATAPATH__0key_1__31_0__20_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__20_), .R(rst_n_bF_buf37), .S(1'b1) );
  DFFSR DFFSR_138 ( .CLK(clk_bF_buf16), .D(AES_CORE_DATAPATH__0key_1__31_0__21_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__21_), .R(rst_n_bF_buf36), .S(1'b1) );
  DFFSR DFFSR_139 ( .CLK(clk_bF_buf15), .D(AES_CORE_DATAPATH__0key_1__31_0__22_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__22_), .R(rst_n_bF_buf35), .S(1'b1) );
  DFFSR DFFSR_14 ( .CLK(clk_bF_buf79), .D(AES_CORE_CONTROL_UNIT__abc_10818_n79), .Q(AES_CORE_CONTROL_UNIT_state_9_), .R(rst_n_bF_buf73), .S(1'b1) );
  DFFSR DFFSR_140 ( .CLK(clk_bF_buf14), .D(AES_CORE_DATAPATH__0key_1__31_0__23_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__23_), .R(rst_n_bF_buf34), .S(1'b1) );
  DFFSR DFFSR_141 ( .CLK(clk_bF_buf13), .D(AES_CORE_DATAPATH__0key_1__31_0__24_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__24_), .R(rst_n_bF_buf33), .S(1'b1) );
  DFFSR DFFSR_142 ( .CLK(clk_bF_buf12), .D(AES_CORE_DATAPATH__0key_1__31_0__25_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__25_), .R(rst_n_bF_buf32), .S(1'b1) );
  DFFSR DFFSR_143 ( .CLK(clk_bF_buf11), .D(AES_CORE_DATAPATH__0key_1__31_0__26_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__26_), .R(rst_n_bF_buf31), .S(1'b1) );
  DFFSR DFFSR_144 ( .CLK(clk_bF_buf10), .D(AES_CORE_DATAPATH__0key_1__31_0__27_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__27_), .R(rst_n_bF_buf30), .S(1'b1) );
  DFFSR DFFSR_145 ( .CLK(clk_bF_buf9), .D(AES_CORE_DATAPATH__0key_1__31_0__28_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__28_), .R(rst_n_bF_buf29), .S(1'b1) );
  DFFSR DFFSR_146 ( .CLK(clk_bF_buf8), .D(AES_CORE_DATAPATH__0key_1__31_0__29_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__29_), .R(rst_n_bF_buf28), .S(1'b1) );
  DFFSR DFFSR_147 ( .CLK(clk_bF_buf7), .D(AES_CORE_DATAPATH__0key_1__31_0__30_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__30_), .R(rst_n_bF_buf27), .S(1'b1) );
  DFFSR DFFSR_148 ( .CLK(clk_bF_buf6), .D(AES_CORE_DATAPATH__0key_1__31_0__31_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__31_), .R(rst_n_bF_buf26), .S(1'b1) );
  DFFSR DFFSR_149 ( .CLK(clk_bF_buf5), .D(AES_CORE_DATAPATH__0key_host_2__31_0__0_), .Q(AES_CORE_DATAPATH_key_host_2__0_), .R(rst_n_bF_buf25), .S(1'b1) );
  DFFSR DFFSR_15 ( .CLK(clk_bF_buf78), .D(AES_CORE_CONTROL_UNIT__abc_10818_n97), .Q(AES_CORE_CONTROL_UNIT_key_gen), .R(rst_n_bF_buf72), .S(1'b1) );
  DFFSR DFFSR_150 ( .CLK(clk_bF_buf4), .D(AES_CORE_DATAPATH__0key_host_2__31_0__1_), .Q(AES_CORE_DATAPATH_key_host_2__1_), .R(rst_n_bF_buf24), .S(1'b1) );
  DFFSR DFFSR_151 ( .CLK(clk_bF_buf3), .D(AES_CORE_DATAPATH__0key_host_2__31_0__2_), .Q(AES_CORE_DATAPATH_key_host_2__2_), .R(rst_n_bF_buf23), .S(1'b1) );
  DFFSR DFFSR_152 ( .CLK(clk_bF_buf2), .D(AES_CORE_DATAPATH__0key_host_2__31_0__3_), .Q(AES_CORE_DATAPATH_key_host_2__3_), .R(rst_n_bF_buf22), .S(1'b1) );
  DFFSR DFFSR_153 ( .CLK(clk_bF_buf1), .D(AES_CORE_DATAPATH__0key_host_2__31_0__4_), .Q(AES_CORE_DATAPATH_key_host_2__4_), .R(rst_n_bF_buf21), .S(1'b1) );
  DFFSR DFFSR_154 ( .CLK(clk_bF_buf0), .D(AES_CORE_DATAPATH__0key_host_2__31_0__5_), .Q(AES_CORE_DATAPATH_key_host_2__5_), .R(rst_n_bF_buf20), .S(1'b1) );
  DFFSR DFFSR_155 ( .CLK(clk_bF_buf92), .D(AES_CORE_DATAPATH__0key_host_2__31_0__6_), .Q(AES_CORE_DATAPATH_key_host_2__6_), .R(rst_n_bF_buf19), .S(1'b1) );
  DFFSR DFFSR_156 ( .CLK(clk_bF_buf91), .D(AES_CORE_DATAPATH__0key_host_2__31_0__7_), .Q(AES_CORE_DATAPATH_key_host_2__7_), .R(rst_n_bF_buf18), .S(1'b1) );
  DFFSR DFFSR_157 ( .CLK(clk_bF_buf90), .D(AES_CORE_DATAPATH__0key_host_2__31_0__8_), .Q(AES_CORE_DATAPATH_key_host_2__8_), .R(rst_n_bF_buf17), .S(1'b1) );
  DFFSR DFFSR_158 ( .CLK(clk_bF_buf89), .D(AES_CORE_DATAPATH__0key_host_2__31_0__9_), .Q(AES_CORE_DATAPATH_key_host_2__9_), .R(rst_n_bF_buf16), .S(1'b1) );
  DFFSR DFFSR_159 ( .CLK(clk_bF_buf88), .D(AES_CORE_DATAPATH__0key_host_2__31_0__10_), .Q(AES_CORE_DATAPATH_key_host_2__10_), .R(rst_n_bF_buf15), .S(1'b1) );
  DFFSR DFFSR_16 ( .CLK(clk_bF_buf77), .D(AES_CORE_CONTROL_UNIT__abc_10818_n306), .Q(AES_CORE_CONTROL_UNIT_state_11_), .R(rst_n_bF_buf71), .S(1'b1) );
  DFFSR DFFSR_160 ( .CLK(clk_bF_buf87), .D(AES_CORE_DATAPATH__0key_host_2__31_0__11_), .Q(AES_CORE_DATAPATH_key_host_2__11_), .R(rst_n_bF_buf14), .S(1'b1) );
  DFFSR DFFSR_161 ( .CLK(clk_bF_buf86), .D(AES_CORE_DATAPATH__0key_host_2__31_0__12_), .Q(AES_CORE_DATAPATH_key_host_2__12_), .R(rst_n_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_162 ( .CLK(clk_bF_buf85), .D(AES_CORE_DATAPATH__0key_host_2__31_0__13_), .Q(AES_CORE_DATAPATH_key_host_2__13_), .R(rst_n_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_163 ( .CLK(clk_bF_buf84), .D(AES_CORE_DATAPATH__0key_host_2__31_0__14_), .Q(AES_CORE_DATAPATH_key_host_2__14_), .R(rst_n_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_164 ( .CLK(clk_bF_buf83), .D(AES_CORE_DATAPATH__0key_host_2__31_0__15_), .Q(AES_CORE_DATAPATH_key_host_2__15_), .R(rst_n_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_165 ( .CLK(clk_bF_buf82), .D(AES_CORE_DATAPATH__0key_host_2__31_0__16_), .Q(AES_CORE_DATAPATH_key_host_2__16_), .R(rst_n_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_166 ( .CLK(clk_bF_buf81), .D(AES_CORE_DATAPATH__0key_host_2__31_0__17_), .Q(AES_CORE_DATAPATH_key_host_2__17_), .R(rst_n_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_167 ( .CLK(clk_bF_buf80), .D(AES_CORE_DATAPATH__0key_host_2__31_0__18_), .Q(AES_CORE_DATAPATH_key_host_2__18_), .R(rst_n_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_168 ( .CLK(clk_bF_buf79), .D(AES_CORE_DATAPATH__0key_host_2__31_0__19_), .Q(AES_CORE_DATAPATH_key_host_2__19_), .R(rst_n_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_169 ( .CLK(clk_bF_buf78), .D(AES_CORE_DATAPATH__0key_host_2__31_0__20_), .Q(AES_CORE_DATAPATH_key_host_2__20_), .R(rst_n_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_17 ( .CLK(clk_bF_buf76), .D(AES_CORE_CONTROL_UNIT__abc_10818_n112), .Q(AES_CORE_CONTROL_UNIT_state_12_), .R(rst_n_bF_buf70), .S(1'b1) );
  DFFSR DFFSR_170 ( .CLK(clk_bF_buf77), .D(AES_CORE_DATAPATH__0key_host_2__31_0__21_), .Q(AES_CORE_DATAPATH_key_host_2__21_), .R(rst_n_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_171 ( .CLK(clk_bF_buf76), .D(AES_CORE_DATAPATH__0key_host_2__31_0__22_), .Q(AES_CORE_DATAPATH_key_host_2__22_), .R(rst_n_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_172 ( .CLK(clk_bF_buf75), .D(AES_CORE_DATAPATH__0key_host_2__31_0__23_), .Q(AES_CORE_DATAPATH_key_host_2__23_), .R(rst_n_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_173 ( .CLK(clk_bF_buf74), .D(AES_CORE_DATAPATH__0key_host_2__31_0__24_), .Q(AES_CORE_DATAPATH_key_host_2__24_), .R(rst_n_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_174 ( .CLK(clk_bF_buf73), .D(AES_CORE_DATAPATH__0key_host_2__31_0__25_), .Q(AES_CORE_DATAPATH_key_host_2__25_), .R(rst_n_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_175 ( .CLK(clk_bF_buf72), .D(AES_CORE_DATAPATH__0key_host_2__31_0__26_), .Q(AES_CORE_DATAPATH_key_host_2__26_), .R(rst_n_bF_buf86), .S(1'b1) );
  DFFSR DFFSR_176 ( .CLK(clk_bF_buf71), .D(AES_CORE_DATAPATH__0key_host_2__31_0__27_), .Q(AES_CORE_DATAPATH_key_host_2__27_), .R(rst_n_bF_buf85), .S(1'b1) );
  DFFSR DFFSR_177 ( .CLK(clk_bF_buf70), .D(AES_CORE_DATAPATH__0key_host_2__31_0__28_), .Q(AES_CORE_DATAPATH_key_host_2__28_), .R(rst_n_bF_buf84), .S(1'b1) );
  DFFSR DFFSR_178 ( .CLK(clk_bF_buf69), .D(AES_CORE_DATAPATH__0key_host_2__31_0__29_), .Q(AES_CORE_DATAPATH_key_host_2__29_), .R(rst_n_bF_buf83), .S(1'b1) );
  DFFSR DFFSR_179 ( .CLK(clk_bF_buf68), .D(AES_CORE_DATAPATH__0key_host_2__31_0__30_), .Q(AES_CORE_DATAPATH_key_host_2__30_), .R(rst_n_bF_buf82), .S(1'b1) );
  DFFSR DFFSR_18 ( .CLK(clk_bF_buf75), .D(AES_CORE_CONTROL_UNIT__abc_10818_n118), .Q(AES_CORE_CONTROL_UNIT_state_13_), .R(rst_n_bF_buf69), .S(1'b1) );
  DFFSR DFFSR_180 ( .CLK(clk_bF_buf67), .D(AES_CORE_DATAPATH__0key_host_2__31_0__31_), .Q(AES_CORE_DATAPATH_key_host_2__31_), .R(rst_n_bF_buf81), .S(1'b1) );
  DFFSR DFFSR_181 ( .CLK(clk_bF_buf66), .D(AES_CORE_DATAPATH__0key_2__31_0__0_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__0_), .R(rst_n_bF_buf80), .S(1'b1) );
  DFFSR DFFSR_182 ( .CLK(clk_bF_buf65), .D(AES_CORE_DATAPATH__0key_2__31_0__1_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__1_), .R(rst_n_bF_buf79), .S(1'b1) );
  DFFSR DFFSR_183 ( .CLK(clk_bF_buf64), .D(AES_CORE_DATAPATH__0key_2__31_0__2_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__2_), .R(rst_n_bF_buf78), .S(1'b1) );
  DFFSR DFFSR_184 ( .CLK(clk_bF_buf63), .D(AES_CORE_DATAPATH__0key_2__31_0__3_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__3_), .R(rst_n_bF_buf77), .S(1'b1) );
  DFFSR DFFSR_185 ( .CLK(clk_bF_buf62), .D(AES_CORE_DATAPATH__0key_2__31_0__4_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__4_), .R(rst_n_bF_buf76), .S(1'b1) );
  DFFSR DFFSR_186 ( .CLK(clk_bF_buf61), .D(AES_CORE_DATAPATH__0key_2__31_0__5_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__5_), .R(rst_n_bF_buf75), .S(1'b1) );
  DFFSR DFFSR_187 ( .CLK(clk_bF_buf60), .D(AES_CORE_DATAPATH__0key_2__31_0__6_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__6_), .R(rst_n_bF_buf74), .S(1'b1) );
  DFFSR DFFSR_188 ( .CLK(clk_bF_buf59), .D(AES_CORE_DATAPATH__0key_2__31_0__7_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__7_), .R(rst_n_bF_buf73), .S(1'b1) );
  DFFSR DFFSR_189 ( .CLK(clk_bF_buf58), .D(AES_CORE_DATAPATH__0key_2__31_0__8_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__8_), .R(rst_n_bF_buf72), .S(1'b1) );
  DFFSR DFFSR_19 ( .CLK(clk_bF_buf74), .D(AES_CORE_CONTROL_UNIT__abc_10818_n122), .Q(AES_CORE_CONTROL_UNIT_state_14_), .R(rst_n_bF_buf68), .S(1'b1) );
  DFFSR DFFSR_190 ( .CLK(clk_bF_buf57), .D(AES_CORE_DATAPATH__0key_2__31_0__9_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__9_), .R(rst_n_bF_buf71), .S(1'b1) );
  DFFSR DFFSR_191 ( .CLK(clk_bF_buf56), .D(AES_CORE_DATAPATH__0key_2__31_0__10_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__10_), .R(rst_n_bF_buf70), .S(1'b1) );
  DFFSR DFFSR_192 ( .CLK(clk_bF_buf55), .D(AES_CORE_DATAPATH__0key_2__31_0__11_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__11_), .R(rst_n_bF_buf69), .S(1'b1) );
  DFFSR DFFSR_193 ( .CLK(clk_bF_buf54), .D(AES_CORE_DATAPATH__0key_2__31_0__12_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__12_), .R(rst_n_bF_buf68), .S(1'b1) );
  DFFSR DFFSR_194 ( .CLK(clk_bF_buf53), .D(AES_CORE_DATAPATH__0key_2__31_0__13_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__13_), .R(rst_n_bF_buf67), .S(1'b1) );
  DFFSR DFFSR_195 ( .CLK(clk_bF_buf52), .D(AES_CORE_DATAPATH__0key_2__31_0__14_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__14_), .R(rst_n_bF_buf66), .S(1'b1) );
  DFFSR DFFSR_196 ( .CLK(clk_bF_buf51), .D(AES_CORE_DATAPATH__0key_2__31_0__15_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__15_), .R(rst_n_bF_buf65), .S(1'b1) );
  DFFSR DFFSR_197 ( .CLK(clk_bF_buf50), .D(AES_CORE_DATAPATH__0key_2__31_0__16_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__16_), .R(rst_n_bF_buf64), .S(1'b1) );
  DFFSR DFFSR_198 ( .CLK(clk_bF_buf49), .D(AES_CORE_DATAPATH__0key_2__31_0__17_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__17_), .R(rst_n_bF_buf63), .S(1'b1) );
  DFFSR DFFSR_199 ( .CLK(clk_bF_buf48), .D(AES_CORE_DATAPATH__0key_2__31_0__18_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__18_), .R(rst_n_bF_buf62), .S(1'b1) );
  DFFSR DFFSR_2 ( .CLK(clk_bF_buf91), .D(AES_CORE_CONTROL_UNIT_rd_count_1__FF_INPUT), .Q(AES_CORE_CONTROL_UNIT_rd_count_1_), .R(rst_n_bF_buf85), .S(1'b1) );
  DFFSR DFFSR_20 ( .CLK(clk_bF_buf73), .D(AES_CORE_CONTROL_UNIT__abc_10818_n307), .Q(AES_CORE_CONTROL_UNIT_state_15_), .R(rst_n_bF_buf67), .S(1'b1) );
  DFFSR DFFSR_200 ( .CLK(clk_bF_buf47), .D(AES_CORE_DATAPATH__0key_2__31_0__19_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__19_), .R(rst_n_bF_buf61), .S(1'b1) );
  DFFSR DFFSR_201 ( .CLK(clk_bF_buf46), .D(AES_CORE_DATAPATH__0key_2__31_0__20_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__20_), .R(rst_n_bF_buf60), .S(1'b1) );
  DFFSR DFFSR_202 ( .CLK(clk_bF_buf45), .D(AES_CORE_DATAPATH__0key_2__31_0__21_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__21_), .R(rst_n_bF_buf59), .S(1'b1) );
  DFFSR DFFSR_203 ( .CLK(clk_bF_buf44), .D(AES_CORE_DATAPATH__0key_2__31_0__22_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__22_), .R(rst_n_bF_buf58), .S(1'b1) );
  DFFSR DFFSR_204 ( .CLK(clk_bF_buf43), .D(AES_CORE_DATAPATH__0key_2__31_0__23_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__23_), .R(rst_n_bF_buf57), .S(1'b1) );
  DFFSR DFFSR_205 ( .CLK(clk_bF_buf42), .D(AES_CORE_DATAPATH__0key_2__31_0__24_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__24_), .R(rst_n_bF_buf56), .S(1'b1) );
  DFFSR DFFSR_206 ( .CLK(clk_bF_buf41), .D(AES_CORE_DATAPATH__0key_2__31_0__25_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__25_), .R(rst_n_bF_buf55), .S(1'b1) );
  DFFSR DFFSR_207 ( .CLK(clk_bF_buf40), .D(AES_CORE_DATAPATH__0key_2__31_0__26_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__26_), .R(rst_n_bF_buf54), .S(1'b1) );
  DFFSR DFFSR_208 ( .CLK(clk_bF_buf39), .D(AES_CORE_DATAPATH__0key_2__31_0__27_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__27_), .R(rst_n_bF_buf53), .S(1'b1) );
  DFFSR DFFSR_209 ( .CLK(clk_bF_buf38), .D(AES_CORE_DATAPATH__0key_2__31_0__28_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__28_), .R(rst_n_bF_buf52), .S(1'b1) );
  DFFSR DFFSR_21 ( .CLK(clk_bF_buf40), .D(AES_CORE_DATAPATH__0key_host_0__31_0__0_), .Q(AES_CORE_DATAPATH_key_host_0__0_), .R(rst_n_bF_buf66), .S(1'b1) );
  DFFSR DFFSR_210 ( .CLK(clk_bF_buf37), .D(AES_CORE_DATAPATH__0key_2__31_0__29_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__29_), .R(rst_n_bF_buf51), .S(1'b1) );
  DFFSR DFFSR_211 ( .CLK(clk_bF_buf36), .D(AES_CORE_DATAPATH__0key_2__31_0__30_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__30_), .R(rst_n_bF_buf50), .S(1'b1) );
  DFFSR DFFSR_212 ( .CLK(clk_bF_buf35), .D(AES_CORE_DATAPATH__0key_2__31_0__31_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__31_), .R(rst_n_bF_buf49), .S(1'b1) );
  DFFSR DFFSR_213 ( .CLK(clk_bF_buf34), .D(AES_CORE_DATAPATH__0key_host_3__31_0__0_), .Q(AES_CORE_DATAPATH_key_host_3__0_), .R(rst_n_bF_buf48), .S(1'b1) );
  DFFSR DFFSR_214 ( .CLK(clk_bF_buf33), .D(AES_CORE_DATAPATH__0key_host_3__31_0__1_), .Q(AES_CORE_DATAPATH_key_host_3__1_), .R(rst_n_bF_buf47), .S(1'b1) );
  DFFSR DFFSR_215 ( .CLK(clk_bF_buf32), .D(AES_CORE_DATAPATH__0key_host_3__31_0__2_), .Q(AES_CORE_DATAPATH_key_host_3__2_), .R(rst_n_bF_buf46), .S(1'b1) );
  DFFSR DFFSR_216 ( .CLK(clk_bF_buf31), .D(AES_CORE_DATAPATH__0key_host_3__31_0__3_), .Q(AES_CORE_DATAPATH_key_host_3__3_), .R(rst_n_bF_buf45), .S(1'b1) );
  DFFSR DFFSR_217 ( .CLK(clk_bF_buf30), .D(AES_CORE_DATAPATH__0key_host_3__31_0__4_), .Q(AES_CORE_DATAPATH_key_host_3__4_), .R(rst_n_bF_buf44), .S(1'b1) );
  DFFSR DFFSR_218 ( .CLK(clk_bF_buf29), .D(AES_CORE_DATAPATH__0key_host_3__31_0__5_), .Q(AES_CORE_DATAPATH_key_host_3__5_), .R(rst_n_bF_buf43), .S(1'b1) );
  DFFSR DFFSR_219 ( .CLK(clk_bF_buf28), .D(AES_CORE_DATAPATH__0key_host_3__31_0__6_), .Q(AES_CORE_DATAPATH_key_host_3__6_), .R(rst_n_bF_buf42), .S(1'b1) );
  DFFSR DFFSR_22 ( .CLK(clk_bF_buf39), .D(AES_CORE_DATAPATH__0key_host_0__31_0__1_), .Q(AES_CORE_DATAPATH_key_host_0__1_), .R(rst_n_bF_buf65), .S(1'b1) );
  DFFSR DFFSR_220 ( .CLK(clk_bF_buf27), .D(AES_CORE_DATAPATH__0key_host_3__31_0__7_), .Q(AES_CORE_DATAPATH_key_host_3__7_), .R(rst_n_bF_buf41), .S(1'b1) );
  DFFSR DFFSR_221 ( .CLK(clk_bF_buf26), .D(AES_CORE_DATAPATH__0key_host_3__31_0__8_), .Q(AES_CORE_DATAPATH_key_host_3__8_), .R(rst_n_bF_buf40), .S(1'b1) );
  DFFSR DFFSR_222 ( .CLK(clk_bF_buf25), .D(AES_CORE_DATAPATH__0key_host_3__31_0__9_), .Q(AES_CORE_DATAPATH_key_host_3__9_), .R(rst_n_bF_buf39), .S(1'b1) );
  DFFSR DFFSR_223 ( .CLK(clk_bF_buf24), .D(AES_CORE_DATAPATH__0key_host_3__31_0__10_), .Q(AES_CORE_DATAPATH_key_host_3__10_), .R(rst_n_bF_buf38), .S(1'b1) );
  DFFSR DFFSR_224 ( .CLK(clk_bF_buf23), .D(AES_CORE_DATAPATH__0key_host_3__31_0__11_), .Q(AES_CORE_DATAPATH_key_host_3__11_), .R(rst_n_bF_buf37), .S(1'b1) );
  DFFSR DFFSR_225 ( .CLK(clk_bF_buf22), .D(AES_CORE_DATAPATH__0key_host_3__31_0__12_), .Q(AES_CORE_DATAPATH_key_host_3__12_), .R(rst_n_bF_buf36), .S(1'b1) );
  DFFSR DFFSR_226 ( .CLK(clk_bF_buf21), .D(AES_CORE_DATAPATH__0key_host_3__31_0__13_), .Q(AES_CORE_DATAPATH_key_host_3__13_), .R(rst_n_bF_buf35), .S(1'b1) );
  DFFSR DFFSR_227 ( .CLK(clk_bF_buf20), .D(AES_CORE_DATAPATH__0key_host_3__31_0__14_), .Q(AES_CORE_DATAPATH_key_host_3__14_), .R(rst_n_bF_buf34), .S(1'b1) );
  DFFSR DFFSR_228 ( .CLK(clk_bF_buf19), .D(AES_CORE_DATAPATH__0key_host_3__31_0__15_), .Q(AES_CORE_DATAPATH_key_host_3__15_), .R(rst_n_bF_buf33), .S(1'b1) );
  DFFSR DFFSR_229 ( .CLK(clk_bF_buf18), .D(AES_CORE_DATAPATH__0key_host_3__31_0__16_), .Q(AES_CORE_DATAPATH_key_host_3__16_), .R(rst_n_bF_buf32), .S(1'b1) );
  DFFSR DFFSR_23 ( .CLK(clk_bF_buf38), .D(AES_CORE_DATAPATH__0key_host_0__31_0__2_), .Q(AES_CORE_DATAPATH_key_host_0__2_), .R(rst_n_bF_buf64), .S(1'b1) );
  DFFSR DFFSR_230 ( .CLK(clk_bF_buf17), .D(AES_CORE_DATAPATH__0key_host_3__31_0__17_), .Q(AES_CORE_DATAPATH_key_host_3__17_), .R(rst_n_bF_buf31), .S(1'b1) );
  DFFSR DFFSR_231 ( .CLK(clk_bF_buf16), .D(AES_CORE_DATAPATH__0key_host_3__31_0__18_), .Q(AES_CORE_DATAPATH_key_host_3__18_), .R(rst_n_bF_buf30), .S(1'b1) );
  DFFSR DFFSR_232 ( .CLK(clk_bF_buf15), .D(AES_CORE_DATAPATH__0key_host_3__31_0__19_), .Q(AES_CORE_DATAPATH_key_host_3__19_), .R(rst_n_bF_buf29), .S(1'b1) );
  DFFSR DFFSR_233 ( .CLK(clk_bF_buf14), .D(AES_CORE_DATAPATH__0key_host_3__31_0__20_), .Q(AES_CORE_DATAPATH_key_host_3__20_), .R(rst_n_bF_buf28), .S(1'b1) );
  DFFSR DFFSR_234 ( .CLK(clk_bF_buf13), .D(AES_CORE_DATAPATH__0key_host_3__31_0__21_), .Q(AES_CORE_DATAPATH_key_host_3__21_), .R(rst_n_bF_buf27), .S(1'b1) );
  DFFSR DFFSR_235 ( .CLK(clk_bF_buf12), .D(AES_CORE_DATAPATH__0key_host_3__31_0__22_), .Q(AES_CORE_DATAPATH_key_host_3__22_), .R(rst_n_bF_buf26), .S(1'b1) );
  DFFSR DFFSR_236 ( .CLK(clk_bF_buf11), .D(AES_CORE_DATAPATH__0key_host_3__31_0__23_), .Q(AES_CORE_DATAPATH_key_host_3__23_), .R(rst_n_bF_buf25), .S(1'b1) );
  DFFSR DFFSR_237 ( .CLK(clk_bF_buf10), .D(AES_CORE_DATAPATH__0key_host_3__31_0__24_), .Q(AES_CORE_DATAPATH_key_host_3__24_), .R(rst_n_bF_buf24), .S(1'b1) );
  DFFSR DFFSR_238 ( .CLK(clk_bF_buf9), .D(AES_CORE_DATAPATH__0key_host_3__31_0__25_), .Q(AES_CORE_DATAPATH_key_host_3__25_), .R(rst_n_bF_buf23), .S(1'b1) );
  DFFSR DFFSR_239 ( .CLK(clk_bF_buf8), .D(AES_CORE_DATAPATH__0key_host_3__31_0__26_), .Q(AES_CORE_DATAPATH_key_host_3__26_), .R(rst_n_bF_buf22), .S(1'b1) );
  DFFSR DFFSR_24 ( .CLK(clk_bF_buf37), .D(AES_CORE_DATAPATH__0key_host_0__31_0__3_), .Q(AES_CORE_DATAPATH_key_host_0__3_), .R(rst_n_bF_buf63), .S(1'b1) );
  DFFSR DFFSR_240 ( .CLK(clk_bF_buf7), .D(AES_CORE_DATAPATH__0key_host_3__31_0__27_), .Q(AES_CORE_DATAPATH_key_host_3__27_), .R(rst_n_bF_buf21), .S(1'b1) );
  DFFSR DFFSR_241 ( .CLK(clk_bF_buf6), .D(AES_CORE_DATAPATH__0key_host_3__31_0__28_), .Q(AES_CORE_DATAPATH_key_host_3__28_), .R(rst_n_bF_buf20), .S(1'b1) );
  DFFSR DFFSR_242 ( .CLK(clk_bF_buf5), .D(AES_CORE_DATAPATH__0key_host_3__31_0__29_), .Q(AES_CORE_DATAPATH_key_host_3__29_), .R(rst_n_bF_buf19), .S(1'b1) );
  DFFSR DFFSR_243 ( .CLK(clk_bF_buf4), .D(AES_CORE_DATAPATH__0key_host_3__31_0__30_), .Q(AES_CORE_DATAPATH_key_host_3__30_), .R(rst_n_bF_buf18), .S(1'b1) );
  DFFSR DFFSR_244 ( .CLK(clk_bF_buf3), .D(AES_CORE_DATAPATH__0key_host_3__31_0__31_), .Q(AES_CORE_DATAPATH_key_host_3__31_), .R(rst_n_bF_buf17), .S(1'b1) );
  DFFSR DFFSR_245 ( .CLK(clk_bF_buf2), .D(AES_CORE_DATAPATH__0key_3__31_0__0_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__0_), .R(rst_n_bF_buf16), .S(1'b1) );
  DFFSR DFFSR_246 ( .CLK(clk_bF_buf1), .D(AES_CORE_DATAPATH__0key_3__31_0__1_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__1_), .R(rst_n_bF_buf15), .S(1'b1) );
  DFFSR DFFSR_247 ( .CLK(clk_bF_buf0), .D(AES_CORE_DATAPATH__0key_3__31_0__2_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__2_), .R(rst_n_bF_buf14), .S(1'b1) );
  DFFSR DFFSR_248 ( .CLK(clk_bF_buf92), .D(AES_CORE_DATAPATH__0key_3__31_0__3_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__3_), .R(rst_n_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_249 ( .CLK(clk_bF_buf91), .D(AES_CORE_DATAPATH__0key_3__31_0__4_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__4_), .R(rst_n_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_25 ( .CLK(clk_bF_buf36), .D(AES_CORE_DATAPATH__0key_host_0__31_0__4_), .Q(AES_CORE_DATAPATH_key_host_0__4_), .R(rst_n_bF_buf62), .S(1'b1) );
  DFFSR DFFSR_250 ( .CLK(clk_bF_buf90), .D(AES_CORE_DATAPATH__0key_3__31_0__5_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__5_), .R(rst_n_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_251 ( .CLK(clk_bF_buf89), .D(AES_CORE_DATAPATH__0key_3__31_0__6_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__6_), .R(rst_n_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_252 ( .CLK(clk_bF_buf88), .D(AES_CORE_DATAPATH__0key_3__31_0__7_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__7_), .R(rst_n_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_253 ( .CLK(clk_bF_buf87), .D(AES_CORE_DATAPATH__0key_3__31_0__8_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__8_), .R(rst_n_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_254 ( .CLK(clk_bF_buf86), .D(AES_CORE_DATAPATH__0key_3__31_0__9_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__9_), .R(rst_n_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_255 ( .CLK(clk_bF_buf85), .D(AES_CORE_DATAPATH__0key_3__31_0__10_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__10_), .R(rst_n_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_256 ( .CLK(clk_bF_buf84), .D(AES_CORE_DATAPATH__0key_3__31_0__11_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__11_), .R(rst_n_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_257 ( .CLK(clk_bF_buf83), .D(AES_CORE_DATAPATH__0key_3__31_0__12_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__12_), .R(rst_n_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_258 ( .CLK(clk_bF_buf82), .D(AES_CORE_DATAPATH__0key_3__31_0__13_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__13_), .R(rst_n_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_259 ( .CLK(clk_bF_buf81), .D(AES_CORE_DATAPATH__0key_3__31_0__14_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__14_), .R(rst_n_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_26 ( .CLK(clk_bF_buf35), .D(AES_CORE_DATAPATH__0key_host_0__31_0__5_), .Q(AES_CORE_DATAPATH_key_host_0__5_), .R(rst_n_bF_buf61), .S(1'b1) );
  DFFSR DFFSR_260 ( .CLK(clk_bF_buf80), .D(AES_CORE_DATAPATH__0key_3__31_0__15_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__15_), .R(rst_n_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_261 ( .CLK(clk_bF_buf79), .D(AES_CORE_DATAPATH__0key_3__31_0__16_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__16_), .R(rst_n_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_262 ( .CLK(clk_bF_buf78), .D(AES_CORE_DATAPATH__0key_3__31_0__17_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__17_), .R(rst_n_bF_buf86), .S(1'b1) );
  DFFSR DFFSR_263 ( .CLK(clk_bF_buf77), .D(AES_CORE_DATAPATH__0key_3__31_0__18_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__18_), .R(rst_n_bF_buf85), .S(1'b1) );
  DFFSR DFFSR_264 ( .CLK(clk_bF_buf76), .D(AES_CORE_DATAPATH__0key_3__31_0__19_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__19_), .R(rst_n_bF_buf84), .S(1'b1) );
  DFFSR DFFSR_265 ( .CLK(clk_bF_buf75), .D(AES_CORE_DATAPATH__0key_3__31_0__20_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__20_), .R(rst_n_bF_buf83), .S(1'b1) );
  DFFSR DFFSR_266 ( .CLK(clk_bF_buf74), .D(AES_CORE_DATAPATH__0key_3__31_0__21_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__21_), .R(rst_n_bF_buf82), .S(1'b1) );
  DFFSR DFFSR_267 ( .CLK(clk_bF_buf73), .D(AES_CORE_DATAPATH__0key_3__31_0__22_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__22_), .R(rst_n_bF_buf81), .S(1'b1) );
  DFFSR DFFSR_268 ( .CLK(clk_bF_buf72), .D(AES_CORE_DATAPATH__0key_3__31_0__23_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__23_), .R(rst_n_bF_buf80), .S(1'b1) );
  DFFSR DFFSR_269 ( .CLK(clk_bF_buf71), .D(AES_CORE_DATAPATH__0key_3__31_0__24_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__24_), .R(rst_n_bF_buf79), .S(1'b1) );
  DFFSR DFFSR_27 ( .CLK(clk_bF_buf34), .D(AES_CORE_DATAPATH__0key_host_0__31_0__6_), .Q(AES_CORE_DATAPATH_key_host_0__6_), .R(rst_n_bF_buf60), .S(1'b1) );
  DFFSR DFFSR_270 ( .CLK(clk_bF_buf70), .D(AES_CORE_DATAPATH__0key_3__31_0__25_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__25_), .R(rst_n_bF_buf78), .S(1'b1) );
  DFFSR DFFSR_271 ( .CLK(clk_bF_buf69), .D(AES_CORE_DATAPATH__0key_3__31_0__26_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__26_), .R(rst_n_bF_buf77), .S(1'b1) );
  DFFSR DFFSR_272 ( .CLK(clk_bF_buf68), .D(AES_CORE_DATAPATH__0key_3__31_0__27_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__27_), .R(rst_n_bF_buf76), .S(1'b1) );
  DFFSR DFFSR_273 ( .CLK(clk_bF_buf67), .D(AES_CORE_DATAPATH__0key_3__31_0__28_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__28_), .R(rst_n_bF_buf75), .S(1'b1) );
  DFFSR DFFSR_274 ( .CLK(clk_bF_buf66), .D(AES_CORE_DATAPATH__0key_3__31_0__29_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__29_), .R(rst_n_bF_buf74), .S(1'b1) );
  DFFSR DFFSR_275 ( .CLK(clk_bF_buf65), .D(AES_CORE_DATAPATH__0key_3__31_0__30_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__30_), .R(rst_n_bF_buf73), .S(1'b1) );
  DFFSR DFFSR_276 ( .CLK(clk_bF_buf64), .D(AES_CORE_DATAPATH__0key_3__31_0__31_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__31_), .R(rst_n_bF_buf72), .S(1'b1) );
  DFFSR DFFSR_277 ( .CLK(clk_bF_buf63), .D(AES_CORE_DATAPATH__0col_0__31_0__0_), .Q(AES_CORE_DATAPATH_col_0__0_), .R(rst_n_bF_buf71), .S(1'b1) );
  DFFSR DFFSR_278 ( .CLK(clk_bF_buf62), .D(AES_CORE_DATAPATH__0col_0__31_0__1_), .Q(AES_CORE_DATAPATH_col_0__1_), .R(rst_n_bF_buf70), .S(1'b1) );
  DFFSR DFFSR_279 ( .CLK(clk_bF_buf61), .D(AES_CORE_DATAPATH__0col_0__31_0__2_), .Q(AES_CORE_DATAPATH_col_0__2_), .R(rst_n_bF_buf69), .S(1'b1) );
  DFFSR DFFSR_28 ( .CLK(clk_bF_buf33), .D(AES_CORE_DATAPATH__0key_host_0__31_0__7_), .Q(AES_CORE_DATAPATH_key_host_0__7_), .R(rst_n_bF_buf59), .S(1'b1) );
  DFFSR DFFSR_280 ( .CLK(clk_bF_buf60), .D(AES_CORE_DATAPATH__0col_0__31_0__3_), .Q(AES_CORE_DATAPATH_col_0__3_), .R(rst_n_bF_buf68), .S(1'b1) );
  DFFSR DFFSR_281 ( .CLK(clk_bF_buf59), .D(AES_CORE_DATAPATH__0col_0__31_0__4_), .Q(AES_CORE_DATAPATH_col_0__4_), .R(rst_n_bF_buf67), .S(1'b1) );
  DFFSR DFFSR_282 ( .CLK(clk_bF_buf58), .D(AES_CORE_DATAPATH__0col_0__31_0__5_), .Q(AES_CORE_DATAPATH_col_0__5_), .R(rst_n_bF_buf66), .S(1'b1) );
  DFFSR DFFSR_283 ( .CLK(clk_bF_buf57), .D(AES_CORE_DATAPATH__0col_0__31_0__6_), .Q(AES_CORE_DATAPATH_col_0__6_), .R(rst_n_bF_buf65), .S(1'b1) );
  DFFSR DFFSR_284 ( .CLK(clk_bF_buf56), .D(AES_CORE_DATAPATH__0col_0__31_0__7_), .Q(AES_CORE_DATAPATH_col_0__7_), .R(rst_n_bF_buf64), .S(1'b1) );
  DFFSR DFFSR_285 ( .CLK(clk_bF_buf55), .D(AES_CORE_DATAPATH__0col_0__31_0__8_), .Q(AES_CORE_DATAPATH_col_0__8_), .R(rst_n_bF_buf63), .S(1'b1) );
  DFFSR DFFSR_286 ( .CLK(clk_bF_buf54), .D(AES_CORE_DATAPATH__0col_0__31_0__9_), .Q(AES_CORE_DATAPATH_col_0__9_), .R(rst_n_bF_buf62), .S(1'b1) );
  DFFSR DFFSR_287 ( .CLK(clk_bF_buf53), .D(AES_CORE_DATAPATH__0col_0__31_0__10_), .Q(AES_CORE_DATAPATH_col_0__10_), .R(rst_n_bF_buf61), .S(1'b1) );
  DFFSR DFFSR_288 ( .CLK(clk_bF_buf52), .D(AES_CORE_DATAPATH__0col_0__31_0__11_), .Q(AES_CORE_DATAPATH_col_0__11_), .R(rst_n_bF_buf60), .S(1'b1) );
  DFFSR DFFSR_289 ( .CLK(clk_bF_buf51), .D(AES_CORE_DATAPATH__0col_0__31_0__12_), .Q(AES_CORE_DATAPATH_col_0__12_), .R(rst_n_bF_buf59), .S(1'b1) );
  DFFSR DFFSR_29 ( .CLK(clk_bF_buf32), .D(AES_CORE_DATAPATH__0key_host_0__31_0__8_), .Q(AES_CORE_DATAPATH_key_host_0__8_), .R(rst_n_bF_buf58), .S(1'b1) );
  DFFSR DFFSR_290 ( .CLK(clk_bF_buf50), .D(AES_CORE_DATAPATH__0col_0__31_0__13_), .Q(AES_CORE_DATAPATH_col_0__13_), .R(rst_n_bF_buf58), .S(1'b1) );
  DFFSR DFFSR_291 ( .CLK(clk_bF_buf49), .D(AES_CORE_DATAPATH__0col_0__31_0__14_), .Q(AES_CORE_DATAPATH_col_0__14_), .R(rst_n_bF_buf57), .S(1'b1) );
  DFFSR DFFSR_292 ( .CLK(clk_bF_buf48), .D(AES_CORE_DATAPATH__0col_0__31_0__15_), .Q(AES_CORE_DATAPATH_col_0__15_), .R(rst_n_bF_buf56), .S(1'b1) );
  DFFSR DFFSR_293 ( .CLK(clk_bF_buf47), .D(AES_CORE_DATAPATH__0col_0__31_0__16_), .Q(AES_CORE_DATAPATH_col_0__16_), .R(rst_n_bF_buf55), .S(1'b1) );
  DFFSR DFFSR_294 ( .CLK(clk_bF_buf46), .D(AES_CORE_DATAPATH__0col_0__31_0__17_), .Q(AES_CORE_DATAPATH_col_0__17_), .R(rst_n_bF_buf54), .S(1'b1) );
  DFFSR DFFSR_295 ( .CLK(clk_bF_buf45), .D(AES_CORE_DATAPATH__0col_0__31_0__18_), .Q(AES_CORE_DATAPATH_col_0__18_), .R(rst_n_bF_buf53), .S(1'b1) );
  DFFSR DFFSR_296 ( .CLK(clk_bF_buf44), .D(AES_CORE_DATAPATH__0col_0__31_0__19_), .Q(AES_CORE_DATAPATH_col_0__19_), .R(rst_n_bF_buf52), .S(1'b1) );
  DFFSR DFFSR_297 ( .CLK(clk_bF_buf43), .D(AES_CORE_DATAPATH__0col_0__31_0__20_), .Q(AES_CORE_DATAPATH_col_0__20_), .R(rst_n_bF_buf51), .S(1'b1) );
  DFFSR DFFSR_298 ( .CLK(clk_bF_buf42), .D(AES_CORE_DATAPATH__0col_0__31_0__21_), .Q(AES_CORE_DATAPATH_col_0__21_), .R(rst_n_bF_buf50), .S(1'b1) );
  DFFSR DFFSR_299 ( .CLK(clk_bF_buf41), .D(AES_CORE_DATAPATH__0col_0__31_0__22_), .Q(AES_CORE_DATAPATH_col_0__22_), .R(rst_n_bF_buf49), .S(1'b1) );
  DFFSR DFFSR_3 ( .CLK(clk_bF_buf90), .D(AES_CORE_CONTROL_UNIT_rd_count_2__FF_INPUT), .Q(AES_CORE_CONTROL_UNIT_rd_count_2_), .R(rst_n_bF_buf84), .S(1'b1) );
  DFFSR DFFSR_30 ( .CLK(clk_bF_buf31), .D(AES_CORE_DATAPATH__0key_host_0__31_0__9_), .Q(AES_CORE_DATAPATH_key_host_0__9_), .R(rst_n_bF_buf57), .S(1'b1) );
  DFFSR DFFSR_300 ( .CLK(clk_bF_buf40), .D(AES_CORE_DATAPATH__0col_0__31_0__23_), .Q(AES_CORE_DATAPATH_col_0__23_), .R(rst_n_bF_buf48), .S(1'b1) );
  DFFSR DFFSR_301 ( .CLK(clk_bF_buf39), .D(AES_CORE_DATAPATH__0col_0__31_0__24_), .Q(AES_CORE_DATAPATH_col_0__24_), .R(rst_n_bF_buf47), .S(1'b1) );
  DFFSR DFFSR_302 ( .CLK(clk_bF_buf38), .D(AES_CORE_DATAPATH__0col_0__31_0__25_), .Q(AES_CORE_DATAPATH_col_0__25_), .R(rst_n_bF_buf46), .S(1'b1) );
  DFFSR DFFSR_303 ( .CLK(clk_bF_buf37), .D(AES_CORE_DATAPATH__0col_0__31_0__26_), .Q(AES_CORE_DATAPATH_col_0__26_), .R(rst_n_bF_buf45), .S(1'b1) );
  DFFSR DFFSR_304 ( .CLK(clk_bF_buf36), .D(AES_CORE_DATAPATH__0col_0__31_0__27_), .Q(AES_CORE_DATAPATH_col_0__27_), .R(rst_n_bF_buf44), .S(1'b1) );
  DFFSR DFFSR_305 ( .CLK(clk_bF_buf35), .D(AES_CORE_DATAPATH__0col_0__31_0__28_), .Q(AES_CORE_DATAPATH_col_0__28_), .R(rst_n_bF_buf43), .S(1'b1) );
  DFFSR DFFSR_306 ( .CLK(clk_bF_buf34), .D(AES_CORE_DATAPATH__0col_0__31_0__29_), .Q(AES_CORE_DATAPATH_col_0__29_), .R(rst_n_bF_buf42), .S(1'b1) );
  DFFSR DFFSR_307 ( .CLK(clk_bF_buf33), .D(AES_CORE_DATAPATH__0col_0__31_0__30_), .Q(AES_CORE_DATAPATH_col_0__30_), .R(rst_n_bF_buf41), .S(1'b1) );
  DFFSR DFFSR_308 ( .CLK(clk_bF_buf32), .D(AES_CORE_DATAPATH__0col_0__31_0__31_), .Q(AES_CORE_DATAPATH_col_0__31_), .R(rst_n_bF_buf40), .S(1'b1) );
  DFFSR DFFSR_309 ( .CLK(clk_bF_buf31), .D(AES_CORE_DATAPATH__0col_1__31_0__0_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_64_), .R(rst_n_bF_buf39), .S(1'b1) );
  DFFSR DFFSR_31 ( .CLK(clk_bF_buf30), .D(AES_CORE_DATAPATH__0key_host_0__31_0__10_), .Q(AES_CORE_DATAPATH_key_host_0__10_), .R(rst_n_bF_buf56), .S(1'b1) );
  DFFSR DFFSR_310 ( .CLK(clk_bF_buf30), .D(AES_CORE_DATAPATH__0col_1__31_0__1_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_65_), .R(rst_n_bF_buf38), .S(1'b1) );
  DFFSR DFFSR_311 ( .CLK(clk_bF_buf29), .D(AES_CORE_DATAPATH__0col_1__31_0__2_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_66_), .R(rst_n_bF_buf37), .S(1'b1) );
  DFFSR DFFSR_312 ( .CLK(clk_bF_buf28), .D(AES_CORE_DATAPATH__0col_1__31_0__3_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_67_), .R(rst_n_bF_buf36), .S(1'b1) );
  DFFSR DFFSR_313 ( .CLK(clk_bF_buf27), .D(AES_CORE_DATAPATH__0col_1__31_0__4_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_68_), .R(rst_n_bF_buf35), .S(1'b1) );
  DFFSR DFFSR_314 ( .CLK(clk_bF_buf26), .D(AES_CORE_DATAPATH__0col_1__31_0__5_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_69_), .R(rst_n_bF_buf34), .S(1'b1) );
  DFFSR DFFSR_315 ( .CLK(clk_bF_buf25), .D(AES_CORE_DATAPATH__0col_1__31_0__6_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_70_), .R(rst_n_bF_buf33), .S(1'b1) );
  DFFSR DFFSR_316 ( .CLK(clk_bF_buf24), .D(AES_CORE_DATAPATH__0col_1__31_0__7_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_71_), .R(rst_n_bF_buf32), .S(1'b1) );
  DFFSR DFFSR_317 ( .CLK(clk_bF_buf23), .D(AES_CORE_DATAPATH__0col_1__31_0__8_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_72_), .R(rst_n_bF_buf31), .S(1'b1) );
  DFFSR DFFSR_318 ( .CLK(clk_bF_buf22), .D(AES_CORE_DATAPATH__0col_1__31_0__9_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_73_), .R(rst_n_bF_buf30), .S(1'b1) );
  DFFSR DFFSR_319 ( .CLK(clk_bF_buf21), .D(AES_CORE_DATAPATH__0col_1__31_0__10_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_74_), .R(rst_n_bF_buf29), .S(1'b1) );
  DFFSR DFFSR_32 ( .CLK(clk_bF_buf29), .D(AES_CORE_DATAPATH__0key_host_0__31_0__11_), .Q(AES_CORE_DATAPATH_key_host_0__11_), .R(rst_n_bF_buf55), .S(1'b1) );
  DFFSR DFFSR_320 ( .CLK(clk_bF_buf20), .D(AES_CORE_DATAPATH__0col_1__31_0__11_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_75_), .R(rst_n_bF_buf28), .S(1'b1) );
  DFFSR DFFSR_321 ( .CLK(clk_bF_buf19), .D(AES_CORE_DATAPATH__0col_1__31_0__12_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_76_), .R(rst_n_bF_buf27), .S(1'b1) );
  DFFSR DFFSR_322 ( .CLK(clk_bF_buf18), .D(AES_CORE_DATAPATH__0col_1__31_0__13_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_77_), .R(rst_n_bF_buf26), .S(1'b1) );
  DFFSR DFFSR_323 ( .CLK(clk_bF_buf17), .D(AES_CORE_DATAPATH__0col_1__31_0__14_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_78_), .R(rst_n_bF_buf25), .S(1'b1) );
  DFFSR DFFSR_324 ( .CLK(clk_bF_buf16), .D(AES_CORE_DATAPATH__0col_1__31_0__15_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_79_), .R(rst_n_bF_buf24), .S(1'b1) );
  DFFSR DFFSR_325 ( .CLK(clk_bF_buf15), .D(AES_CORE_DATAPATH__0col_1__31_0__16_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_80_), .R(rst_n_bF_buf23), .S(1'b1) );
  DFFSR DFFSR_326 ( .CLK(clk_bF_buf14), .D(AES_CORE_DATAPATH__0col_1__31_0__17_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_81_), .R(rst_n_bF_buf22), .S(1'b1) );
  DFFSR DFFSR_327 ( .CLK(clk_bF_buf13), .D(AES_CORE_DATAPATH__0col_1__31_0__18_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_82_), .R(rst_n_bF_buf21), .S(1'b1) );
  DFFSR DFFSR_328 ( .CLK(clk_bF_buf12), .D(AES_CORE_DATAPATH__0col_1__31_0__19_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_83_), .R(rst_n_bF_buf20), .S(1'b1) );
  DFFSR DFFSR_329 ( .CLK(clk_bF_buf11), .D(AES_CORE_DATAPATH__0col_1__31_0__20_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_84_), .R(rst_n_bF_buf19), .S(1'b1) );
  DFFSR DFFSR_33 ( .CLK(clk_bF_buf28), .D(AES_CORE_DATAPATH__0key_host_0__31_0__12_), .Q(AES_CORE_DATAPATH_key_host_0__12_), .R(rst_n_bF_buf54), .S(1'b1) );
  DFFSR DFFSR_330 ( .CLK(clk_bF_buf10), .D(AES_CORE_DATAPATH__0col_1__31_0__21_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_85_), .R(rst_n_bF_buf18), .S(1'b1) );
  DFFSR DFFSR_331 ( .CLK(clk_bF_buf9), .D(AES_CORE_DATAPATH__0col_1__31_0__22_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_86_), .R(rst_n_bF_buf17), .S(1'b1) );
  DFFSR DFFSR_332 ( .CLK(clk_bF_buf8), .D(AES_CORE_DATAPATH__0col_1__31_0__23_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_87_), .R(rst_n_bF_buf16), .S(1'b1) );
  DFFSR DFFSR_333 ( .CLK(clk_bF_buf7), .D(AES_CORE_DATAPATH__0col_1__31_0__24_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_88_), .R(rst_n_bF_buf15), .S(1'b1) );
  DFFSR DFFSR_334 ( .CLK(clk_bF_buf6), .D(AES_CORE_DATAPATH__0col_1__31_0__25_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_89_), .R(rst_n_bF_buf14), .S(1'b1) );
  DFFSR DFFSR_335 ( .CLK(clk_bF_buf5), .D(AES_CORE_DATAPATH__0col_1__31_0__26_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_90_), .R(rst_n_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_336 ( .CLK(clk_bF_buf4), .D(AES_CORE_DATAPATH__0col_1__31_0__27_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_91_), .R(rst_n_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_337 ( .CLK(clk_bF_buf3), .D(AES_CORE_DATAPATH__0col_1__31_0__28_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_92_), .R(rst_n_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_338 ( .CLK(clk_bF_buf2), .D(AES_CORE_DATAPATH__0col_1__31_0__29_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_93_), .R(rst_n_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_339 ( .CLK(clk_bF_buf1), .D(AES_CORE_DATAPATH__0col_1__31_0__30_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_94_), .R(rst_n_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_34 ( .CLK(clk_bF_buf27), .D(AES_CORE_DATAPATH__0key_host_0__31_0__13_), .Q(AES_CORE_DATAPATH_key_host_0__13_), .R(rst_n_bF_buf53), .S(1'b1) );
  DFFSR DFFSR_340 ( .CLK(clk_bF_buf0), .D(AES_CORE_DATAPATH__0col_1__31_0__31_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_95_), .R(rst_n_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_341 ( .CLK(clk_bF_buf92), .D(AES_CORE_DATAPATH__0col_2__31_0__0_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_32_), .R(rst_n_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_342 ( .CLK(clk_bF_buf91), .D(AES_CORE_DATAPATH__0col_2__31_0__1_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_33_), .R(rst_n_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_343 ( .CLK(clk_bF_buf90), .D(AES_CORE_DATAPATH__0col_2__31_0__2_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_34_), .R(rst_n_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_344 ( .CLK(clk_bF_buf89), .D(AES_CORE_DATAPATH__0col_2__31_0__3_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_35_), .R(rst_n_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_345 ( .CLK(clk_bF_buf88), .D(AES_CORE_DATAPATH__0col_2__31_0__4_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_36_), .R(rst_n_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_346 ( .CLK(clk_bF_buf87), .D(AES_CORE_DATAPATH__0col_2__31_0__5_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_37_), .R(rst_n_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_347 ( .CLK(clk_bF_buf86), .D(AES_CORE_DATAPATH__0col_2__31_0__6_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_38_), .R(rst_n_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_348 ( .CLK(clk_bF_buf85), .D(AES_CORE_DATAPATH__0col_2__31_0__7_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_39_), .R(rst_n_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_349 ( .CLK(clk_bF_buf84), .D(AES_CORE_DATAPATH__0col_2__31_0__8_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_40_), .R(rst_n_bF_buf86), .S(1'b1) );
  DFFSR DFFSR_35 ( .CLK(clk_bF_buf26), .D(AES_CORE_DATAPATH__0key_host_0__31_0__14_), .Q(AES_CORE_DATAPATH_key_host_0__14_), .R(rst_n_bF_buf52), .S(1'b1) );
  DFFSR DFFSR_350 ( .CLK(clk_bF_buf83), .D(AES_CORE_DATAPATH__0col_2__31_0__9_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_41_), .R(rst_n_bF_buf85), .S(1'b1) );
  DFFSR DFFSR_351 ( .CLK(clk_bF_buf82), .D(AES_CORE_DATAPATH__0col_2__31_0__10_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_42_), .R(rst_n_bF_buf84), .S(1'b1) );
  DFFSR DFFSR_352 ( .CLK(clk_bF_buf81), .D(AES_CORE_DATAPATH__0col_2__31_0__11_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_43_), .R(rst_n_bF_buf83), .S(1'b1) );
  DFFSR DFFSR_353 ( .CLK(clk_bF_buf80), .D(AES_CORE_DATAPATH__0col_2__31_0__12_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_44_), .R(rst_n_bF_buf82), .S(1'b1) );
  DFFSR DFFSR_354 ( .CLK(clk_bF_buf79), .D(AES_CORE_DATAPATH__0col_2__31_0__13_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_45_), .R(rst_n_bF_buf81), .S(1'b1) );
  DFFSR DFFSR_355 ( .CLK(clk_bF_buf78), .D(AES_CORE_DATAPATH__0col_2__31_0__14_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_46_), .R(rst_n_bF_buf80), .S(1'b1) );
  DFFSR DFFSR_356 ( .CLK(clk_bF_buf77), .D(AES_CORE_DATAPATH__0col_2__31_0__15_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_47_), .R(rst_n_bF_buf79), .S(1'b1) );
  DFFSR DFFSR_357 ( .CLK(clk_bF_buf76), .D(AES_CORE_DATAPATH__0col_2__31_0__16_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_48_), .R(rst_n_bF_buf78), .S(1'b1) );
  DFFSR DFFSR_358 ( .CLK(clk_bF_buf75), .D(AES_CORE_DATAPATH__0col_2__31_0__17_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_49_), .R(rst_n_bF_buf77), .S(1'b1) );
  DFFSR DFFSR_359 ( .CLK(clk_bF_buf74), .D(AES_CORE_DATAPATH__0col_2__31_0__18_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_50_), .R(rst_n_bF_buf76), .S(1'b1) );
  DFFSR DFFSR_36 ( .CLK(clk_bF_buf25), .D(AES_CORE_DATAPATH__0key_host_0__31_0__15_), .Q(AES_CORE_DATAPATH_key_host_0__15_), .R(rst_n_bF_buf51), .S(1'b1) );
  DFFSR DFFSR_360 ( .CLK(clk_bF_buf73), .D(AES_CORE_DATAPATH__0col_2__31_0__19_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_51_), .R(rst_n_bF_buf75), .S(1'b1) );
  DFFSR DFFSR_361 ( .CLK(clk_bF_buf72), .D(AES_CORE_DATAPATH__0col_2__31_0__20_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_52_), .R(rst_n_bF_buf74), .S(1'b1) );
  DFFSR DFFSR_362 ( .CLK(clk_bF_buf71), .D(AES_CORE_DATAPATH__0col_2__31_0__21_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_53_), .R(rst_n_bF_buf73), .S(1'b1) );
  DFFSR DFFSR_363 ( .CLK(clk_bF_buf70), .D(AES_CORE_DATAPATH__0col_2__31_0__22_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_54_), .R(rst_n_bF_buf72), .S(1'b1) );
  DFFSR DFFSR_364 ( .CLK(clk_bF_buf69), .D(AES_CORE_DATAPATH__0col_2__31_0__23_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_55_), .R(rst_n_bF_buf71), .S(1'b1) );
  DFFSR DFFSR_365 ( .CLK(clk_bF_buf68), .D(AES_CORE_DATAPATH__0col_2__31_0__24_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_56_), .R(rst_n_bF_buf70), .S(1'b1) );
  DFFSR DFFSR_366 ( .CLK(clk_bF_buf67), .D(AES_CORE_DATAPATH__0col_2__31_0__25_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_57_), .R(rst_n_bF_buf69), .S(1'b1) );
  DFFSR DFFSR_367 ( .CLK(clk_bF_buf66), .D(AES_CORE_DATAPATH__0col_2__31_0__26_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_58_), .R(rst_n_bF_buf68), .S(1'b1) );
  DFFSR DFFSR_368 ( .CLK(clk_bF_buf65), .D(AES_CORE_DATAPATH__0col_2__31_0__27_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_59_), .R(rst_n_bF_buf67), .S(1'b1) );
  DFFSR DFFSR_369 ( .CLK(clk_bF_buf64), .D(AES_CORE_DATAPATH__0col_2__31_0__28_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_60_), .R(rst_n_bF_buf66), .S(1'b1) );
  DFFSR DFFSR_37 ( .CLK(clk_bF_buf24), .D(AES_CORE_DATAPATH__0key_host_0__31_0__16_), .Q(AES_CORE_DATAPATH_key_host_0__16_), .R(rst_n_bF_buf50), .S(1'b1) );
  DFFSR DFFSR_370 ( .CLK(clk_bF_buf63), .D(AES_CORE_DATAPATH__0col_2__31_0__29_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_61_), .R(rst_n_bF_buf65), .S(1'b1) );
  DFFSR DFFSR_371 ( .CLK(clk_bF_buf62), .D(AES_CORE_DATAPATH__0col_2__31_0__30_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_62_), .R(rst_n_bF_buf64), .S(1'b1) );
  DFFSR DFFSR_372 ( .CLK(clk_bF_buf61), .D(AES_CORE_DATAPATH__0col_2__31_0__31_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_63_), .R(rst_n_bF_buf63), .S(1'b1) );
  DFFSR DFFSR_373 ( .CLK(clk_bF_buf60), .D(AES_CORE_DATAPATH__0col_3__31_0__0_), .Q(AES_CORE_DATAPATH_col_3__0_), .R(rst_n_bF_buf62), .S(1'b1) );
  DFFSR DFFSR_374 ( .CLK(clk_bF_buf59), .D(AES_CORE_DATAPATH__0col_3__31_0__1_), .Q(AES_CORE_DATAPATH_col_3__1_), .R(rst_n_bF_buf61), .S(1'b1) );
  DFFSR DFFSR_375 ( .CLK(clk_bF_buf58), .D(AES_CORE_DATAPATH__0col_3__31_0__2_), .Q(AES_CORE_DATAPATH_col_3__2_), .R(rst_n_bF_buf60), .S(1'b1) );
  DFFSR DFFSR_376 ( .CLK(clk_bF_buf57), .D(AES_CORE_DATAPATH__0col_3__31_0__3_), .Q(AES_CORE_DATAPATH_col_3__3_), .R(rst_n_bF_buf59), .S(1'b1) );
  DFFSR DFFSR_377 ( .CLK(clk_bF_buf56), .D(AES_CORE_DATAPATH__0col_3__31_0__4_), .Q(AES_CORE_DATAPATH_col_3__4_), .R(rst_n_bF_buf58), .S(1'b1) );
  DFFSR DFFSR_378 ( .CLK(clk_bF_buf55), .D(AES_CORE_DATAPATH__0col_3__31_0__5_), .Q(AES_CORE_DATAPATH_col_3__5_), .R(rst_n_bF_buf57), .S(1'b1) );
  DFFSR DFFSR_379 ( .CLK(clk_bF_buf54), .D(AES_CORE_DATAPATH__0col_3__31_0__6_), .Q(AES_CORE_DATAPATH_col_3__6_), .R(rst_n_bF_buf56), .S(1'b1) );
  DFFSR DFFSR_38 ( .CLK(clk_bF_buf23), .D(AES_CORE_DATAPATH__0key_host_0__31_0__17_), .Q(AES_CORE_DATAPATH_key_host_0__17_), .R(rst_n_bF_buf49), .S(1'b1) );
  DFFSR DFFSR_380 ( .CLK(clk_bF_buf53), .D(AES_CORE_DATAPATH__0col_3__31_0__7_), .Q(AES_CORE_DATAPATH_col_3__7_), .R(rst_n_bF_buf55), .S(1'b1) );
  DFFSR DFFSR_381 ( .CLK(clk_bF_buf52), .D(AES_CORE_DATAPATH__0col_3__31_0__8_), .Q(AES_CORE_DATAPATH_col_3__8_), .R(rst_n_bF_buf54), .S(1'b1) );
  DFFSR DFFSR_382 ( .CLK(clk_bF_buf51), .D(AES_CORE_DATAPATH__0col_3__31_0__9_), .Q(AES_CORE_DATAPATH_col_3__9_), .R(rst_n_bF_buf53), .S(1'b1) );
  DFFSR DFFSR_383 ( .CLK(clk_bF_buf50), .D(AES_CORE_DATAPATH__0col_3__31_0__10_), .Q(AES_CORE_DATAPATH_col_3__10_), .R(rst_n_bF_buf52), .S(1'b1) );
  DFFSR DFFSR_384 ( .CLK(clk_bF_buf49), .D(AES_CORE_DATAPATH__0col_3__31_0__11_), .Q(AES_CORE_DATAPATH_col_3__11_), .R(rst_n_bF_buf51), .S(1'b1) );
  DFFSR DFFSR_385 ( .CLK(clk_bF_buf48), .D(AES_CORE_DATAPATH__0col_3__31_0__12_), .Q(AES_CORE_DATAPATH_col_3__12_), .R(rst_n_bF_buf50), .S(1'b1) );
  DFFSR DFFSR_386 ( .CLK(clk_bF_buf47), .D(AES_CORE_DATAPATH__0col_3__31_0__13_), .Q(AES_CORE_DATAPATH_col_3__13_), .R(rst_n_bF_buf49), .S(1'b1) );
  DFFSR DFFSR_387 ( .CLK(clk_bF_buf46), .D(AES_CORE_DATAPATH__0col_3__31_0__14_), .Q(AES_CORE_DATAPATH_col_3__14_), .R(rst_n_bF_buf48), .S(1'b1) );
  DFFSR DFFSR_388 ( .CLK(clk_bF_buf45), .D(AES_CORE_DATAPATH__0col_3__31_0__15_), .Q(AES_CORE_DATAPATH_col_3__15_), .R(rst_n_bF_buf47), .S(1'b1) );
  DFFSR DFFSR_389 ( .CLK(clk_bF_buf44), .D(AES_CORE_DATAPATH__0col_3__31_0__16_), .Q(AES_CORE_DATAPATH_col_3__16_), .R(rst_n_bF_buf46), .S(1'b1) );
  DFFSR DFFSR_39 ( .CLK(clk_bF_buf22), .D(AES_CORE_DATAPATH__0key_host_0__31_0__18_), .Q(AES_CORE_DATAPATH_key_host_0__18_), .R(rst_n_bF_buf48), .S(1'b1) );
  DFFSR DFFSR_390 ( .CLK(clk_bF_buf43), .D(AES_CORE_DATAPATH__0col_3__31_0__17_), .Q(AES_CORE_DATAPATH_col_3__17_), .R(rst_n_bF_buf45), .S(1'b1) );
  DFFSR DFFSR_391 ( .CLK(clk_bF_buf42), .D(AES_CORE_DATAPATH__0col_3__31_0__18_), .Q(AES_CORE_DATAPATH_col_3__18_), .R(rst_n_bF_buf44), .S(1'b1) );
  DFFSR DFFSR_392 ( .CLK(clk_bF_buf41), .D(AES_CORE_DATAPATH__0col_3__31_0__19_), .Q(AES_CORE_DATAPATH_col_3__19_), .R(rst_n_bF_buf43), .S(1'b1) );
  DFFSR DFFSR_393 ( .CLK(clk_bF_buf40), .D(AES_CORE_DATAPATH__0col_3__31_0__20_), .Q(AES_CORE_DATAPATH_col_3__20_), .R(rst_n_bF_buf42), .S(1'b1) );
  DFFSR DFFSR_394 ( .CLK(clk_bF_buf39), .D(AES_CORE_DATAPATH__0col_3__31_0__21_), .Q(AES_CORE_DATAPATH_col_3__21_), .R(rst_n_bF_buf41), .S(1'b1) );
  DFFSR DFFSR_395 ( .CLK(clk_bF_buf38), .D(AES_CORE_DATAPATH__0col_3__31_0__22_), .Q(AES_CORE_DATAPATH_col_3__22_), .R(rst_n_bF_buf40), .S(1'b1) );
  DFFSR DFFSR_396 ( .CLK(clk_bF_buf37), .D(AES_CORE_DATAPATH__0col_3__31_0__23_), .Q(AES_CORE_DATAPATH_col_3__23_), .R(rst_n_bF_buf39), .S(1'b1) );
  DFFSR DFFSR_397 ( .CLK(clk_bF_buf36), .D(AES_CORE_DATAPATH__0col_3__31_0__24_), .Q(AES_CORE_DATAPATH_col_3__24_), .R(rst_n_bF_buf38), .S(1'b1) );
  DFFSR DFFSR_398 ( .CLK(clk_bF_buf35), .D(AES_CORE_DATAPATH__0col_3__31_0__25_), .Q(AES_CORE_DATAPATH_col_3__25_), .R(rst_n_bF_buf37), .S(1'b1) );
  DFFSR DFFSR_399 ( .CLK(clk_bF_buf34), .D(AES_CORE_DATAPATH__0col_3__31_0__26_), .Q(AES_CORE_DATAPATH_col_3__26_), .R(rst_n_bF_buf36), .S(1'b1) );
  DFFSR DFFSR_4 ( .CLK(clk_bF_buf89), .D(AES_CORE_CONTROL_UNIT_rd_count_3__FF_INPUT), .Q(AES_CORE_CONTROL_UNIT_rd_count_3_), .R(rst_n_bF_buf83), .S(1'b1) );
  DFFSR DFFSR_40 ( .CLK(clk_bF_buf21), .D(AES_CORE_DATAPATH__0key_host_0__31_0__19_), .Q(AES_CORE_DATAPATH_key_host_0__19_), .R(rst_n_bF_buf47), .S(1'b1) );
  DFFSR DFFSR_400 ( .CLK(clk_bF_buf33), .D(AES_CORE_DATAPATH__0col_3__31_0__27_), .Q(AES_CORE_DATAPATH_col_3__27_), .R(rst_n_bF_buf35), .S(1'b1) );
  DFFSR DFFSR_401 ( .CLK(clk_bF_buf32), .D(AES_CORE_DATAPATH__0col_3__31_0__28_), .Q(AES_CORE_DATAPATH_col_3__28_), .R(rst_n_bF_buf34), .S(1'b1) );
  DFFSR DFFSR_402 ( .CLK(clk_bF_buf31), .D(AES_CORE_DATAPATH__0col_3__31_0__29_), .Q(AES_CORE_DATAPATH_col_3__29_), .R(rst_n_bF_buf33), .S(1'b1) );
  DFFSR DFFSR_403 ( .CLK(clk_bF_buf30), .D(AES_CORE_DATAPATH__0col_3__31_0__30_), .Q(AES_CORE_DATAPATH_col_3__30_), .R(rst_n_bF_buf32), .S(1'b1) );
  DFFSR DFFSR_404 ( .CLK(clk_bF_buf29), .D(AES_CORE_DATAPATH__0col_3__31_0__31_), .Q(AES_CORE_DATAPATH_col_3__31_), .R(rst_n_bF_buf31), .S(1'b1) );
  DFFSR DFFSR_405 ( .CLK(clk_bF_buf28), .D(AES_CORE_DATAPATH__0iv_3__31_0__0_), .Q(AES_CORE_DATAPATH_iv_3__0_), .R(rst_n_bF_buf30), .S(1'b1) );
  DFFSR DFFSR_406 ( .CLK(clk_bF_buf27), .D(AES_CORE_DATAPATH__0iv_3__31_0__1_), .Q(AES_CORE_DATAPATH_iv_3__1_), .R(rst_n_bF_buf29), .S(1'b1) );
  DFFSR DFFSR_407 ( .CLK(clk_bF_buf26), .D(AES_CORE_DATAPATH__0iv_3__31_0__2_), .Q(AES_CORE_DATAPATH_iv_3__2_), .R(rst_n_bF_buf28), .S(1'b1) );
  DFFSR DFFSR_408 ( .CLK(clk_bF_buf25), .D(AES_CORE_DATAPATH__0iv_3__31_0__3_), .Q(AES_CORE_DATAPATH_iv_3__3_), .R(rst_n_bF_buf27), .S(1'b1) );
  DFFSR DFFSR_409 ( .CLK(clk_bF_buf24), .D(AES_CORE_DATAPATH__0iv_3__31_0__4_), .Q(AES_CORE_DATAPATH_iv_3__4_), .R(rst_n_bF_buf26), .S(1'b1) );
  DFFSR DFFSR_41 ( .CLK(clk_bF_buf20), .D(AES_CORE_DATAPATH__0key_host_0__31_0__20_), .Q(AES_CORE_DATAPATH_key_host_0__20_), .R(rst_n_bF_buf46), .S(1'b1) );
  DFFSR DFFSR_410 ( .CLK(clk_bF_buf23), .D(AES_CORE_DATAPATH__0iv_3__31_0__5_), .Q(AES_CORE_DATAPATH_iv_3__5_), .R(rst_n_bF_buf25), .S(1'b1) );
  DFFSR DFFSR_411 ( .CLK(clk_bF_buf22), .D(AES_CORE_DATAPATH__0iv_3__31_0__6_), .Q(AES_CORE_DATAPATH_iv_3__6_), .R(rst_n_bF_buf24), .S(1'b1) );
  DFFSR DFFSR_412 ( .CLK(clk_bF_buf21), .D(AES_CORE_DATAPATH__0iv_3__31_0__7_), .Q(AES_CORE_DATAPATH_iv_3__7_), .R(rst_n_bF_buf23), .S(1'b1) );
  DFFSR DFFSR_413 ( .CLK(clk_bF_buf20), .D(AES_CORE_DATAPATH__0iv_3__31_0__8_), .Q(AES_CORE_DATAPATH_iv_3__8_), .R(rst_n_bF_buf22), .S(1'b1) );
  DFFSR DFFSR_414 ( .CLK(clk_bF_buf19), .D(AES_CORE_DATAPATH__0iv_3__31_0__9_), .Q(AES_CORE_DATAPATH_iv_3__9_), .R(rst_n_bF_buf21), .S(1'b1) );
  DFFSR DFFSR_415 ( .CLK(clk_bF_buf18), .D(AES_CORE_DATAPATH__0iv_3__31_0__10_), .Q(AES_CORE_DATAPATH_iv_3__10_), .R(rst_n_bF_buf20), .S(1'b1) );
  DFFSR DFFSR_416 ( .CLK(clk_bF_buf17), .D(AES_CORE_DATAPATH__0iv_3__31_0__11_), .Q(AES_CORE_DATAPATH_iv_3__11_), .R(rst_n_bF_buf19), .S(1'b1) );
  DFFSR DFFSR_417 ( .CLK(clk_bF_buf16), .D(AES_CORE_DATAPATH__0iv_3__31_0__12_), .Q(AES_CORE_DATAPATH_iv_3__12_), .R(rst_n_bF_buf18), .S(1'b1) );
  DFFSR DFFSR_418 ( .CLK(clk_bF_buf15), .D(AES_CORE_DATAPATH__0iv_3__31_0__13_), .Q(AES_CORE_DATAPATH_iv_3__13_), .R(rst_n_bF_buf17), .S(1'b1) );
  DFFSR DFFSR_419 ( .CLK(clk_bF_buf14), .D(AES_CORE_DATAPATH__0iv_3__31_0__14_), .Q(AES_CORE_DATAPATH_iv_3__14_), .R(rst_n_bF_buf16), .S(1'b1) );
  DFFSR DFFSR_42 ( .CLK(clk_bF_buf19), .D(AES_CORE_DATAPATH__0key_host_0__31_0__21_), .Q(AES_CORE_DATAPATH_key_host_0__21_), .R(rst_n_bF_buf45), .S(1'b1) );
  DFFSR DFFSR_420 ( .CLK(clk_bF_buf13), .D(AES_CORE_DATAPATH__0iv_3__31_0__15_), .Q(AES_CORE_DATAPATH_iv_3__15_), .R(rst_n_bF_buf15), .S(1'b1) );
  DFFSR DFFSR_421 ( .CLK(clk_bF_buf12), .D(AES_CORE_DATAPATH__0iv_3__31_0__16_), .Q(AES_CORE_DATAPATH_iv_3__16_), .R(rst_n_bF_buf14), .S(1'b1) );
  DFFSR DFFSR_422 ( .CLK(clk_bF_buf11), .D(AES_CORE_DATAPATH__0iv_3__31_0__17_), .Q(AES_CORE_DATAPATH_iv_3__17_), .R(rst_n_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_423 ( .CLK(clk_bF_buf10), .D(AES_CORE_DATAPATH__0iv_3__31_0__18_), .Q(AES_CORE_DATAPATH_iv_3__18_), .R(rst_n_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_424 ( .CLK(clk_bF_buf9), .D(AES_CORE_DATAPATH__0iv_3__31_0__19_), .Q(AES_CORE_DATAPATH_iv_3__19_), .R(rst_n_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_425 ( .CLK(clk_bF_buf8), .D(AES_CORE_DATAPATH__0iv_3__31_0__20_), .Q(AES_CORE_DATAPATH_iv_3__20_), .R(rst_n_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_426 ( .CLK(clk_bF_buf7), .D(AES_CORE_DATAPATH__0iv_3__31_0__21_), .Q(AES_CORE_DATAPATH_iv_3__21_), .R(rst_n_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_427 ( .CLK(clk_bF_buf6), .D(AES_CORE_DATAPATH__0iv_3__31_0__22_), .Q(AES_CORE_DATAPATH_iv_3__22_), .R(rst_n_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_428 ( .CLK(clk_bF_buf5), .D(AES_CORE_DATAPATH__0iv_3__31_0__23_), .Q(AES_CORE_DATAPATH_iv_3__23_), .R(rst_n_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_429 ( .CLK(clk_bF_buf4), .D(AES_CORE_DATAPATH__0iv_3__31_0__24_), .Q(AES_CORE_DATAPATH_iv_3__24_), .R(rst_n_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_43 ( .CLK(clk_bF_buf18), .D(AES_CORE_DATAPATH__0key_host_0__31_0__22_), .Q(AES_CORE_DATAPATH_key_host_0__22_), .R(rst_n_bF_buf44), .S(1'b1) );
  DFFSR DFFSR_430 ( .CLK(clk_bF_buf3), .D(AES_CORE_DATAPATH__0iv_3__31_0__25_), .Q(AES_CORE_DATAPATH_iv_3__25_), .R(rst_n_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_431 ( .CLK(clk_bF_buf2), .D(AES_CORE_DATAPATH__0iv_3__31_0__26_), .Q(AES_CORE_DATAPATH_iv_3__26_), .R(rst_n_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_432 ( .CLK(clk_bF_buf1), .D(AES_CORE_DATAPATH__0iv_3__31_0__27_), .Q(AES_CORE_DATAPATH_iv_3__27_), .R(rst_n_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_433 ( .CLK(clk_bF_buf0), .D(AES_CORE_DATAPATH__0iv_3__31_0__28_), .Q(AES_CORE_DATAPATH_iv_3__28_), .R(rst_n_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_434 ( .CLK(clk_bF_buf92), .D(AES_CORE_DATAPATH__0iv_3__31_0__29_), .Q(AES_CORE_DATAPATH_iv_3__29_), .R(rst_n_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_435 ( .CLK(clk_bF_buf91), .D(AES_CORE_DATAPATH__0iv_3__31_0__30_), .Q(AES_CORE_DATAPATH_iv_3__30_), .R(rst_n_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_436 ( .CLK(clk_bF_buf90), .D(AES_CORE_DATAPATH__0iv_3__31_0__31_), .Q(AES_CORE_DATAPATH_iv_3__31_), .R(rst_n_bF_buf86), .S(1'b1) );
  DFFSR DFFSR_437 ( .CLK(clk_bF_buf89), .D(AES_CORE_DATAPATH__0bkp_3__31_0__0_), .Q(AES_CORE_DATAPATH_bkp_3__0_), .R(rst_n_bF_buf85), .S(1'b1) );
  DFFSR DFFSR_438 ( .CLK(clk_bF_buf88), .D(AES_CORE_DATAPATH__0bkp_3__31_0__1_), .Q(AES_CORE_DATAPATH_bkp_3__1_), .R(rst_n_bF_buf84), .S(1'b1) );
  DFFSR DFFSR_439 ( .CLK(clk_bF_buf87), .D(AES_CORE_DATAPATH__0bkp_3__31_0__2_), .Q(AES_CORE_DATAPATH_bkp_3__2_), .R(rst_n_bF_buf83), .S(1'b1) );
  DFFSR DFFSR_44 ( .CLK(clk_bF_buf17), .D(AES_CORE_DATAPATH__0key_host_0__31_0__23_), .Q(AES_CORE_DATAPATH_key_host_0__23_), .R(rst_n_bF_buf43), .S(1'b1) );
  DFFSR DFFSR_440 ( .CLK(clk_bF_buf86), .D(AES_CORE_DATAPATH__0bkp_3__31_0__3_), .Q(AES_CORE_DATAPATH_bkp_3__3_), .R(rst_n_bF_buf82), .S(1'b1) );
  DFFSR DFFSR_441 ( .CLK(clk_bF_buf85), .D(AES_CORE_DATAPATH__0bkp_3__31_0__4_), .Q(AES_CORE_DATAPATH_bkp_3__4_), .R(rst_n_bF_buf81), .S(1'b1) );
  DFFSR DFFSR_442 ( .CLK(clk_bF_buf84), .D(AES_CORE_DATAPATH__0bkp_3__31_0__5_), .Q(AES_CORE_DATAPATH_bkp_3__5_), .R(rst_n_bF_buf80), .S(1'b1) );
  DFFSR DFFSR_443 ( .CLK(clk_bF_buf83), .D(AES_CORE_DATAPATH__0bkp_3__31_0__6_), .Q(AES_CORE_DATAPATH_bkp_3__6_), .R(rst_n_bF_buf79), .S(1'b1) );
  DFFSR DFFSR_444 ( .CLK(clk_bF_buf82), .D(AES_CORE_DATAPATH__0bkp_3__31_0__7_), .Q(AES_CORE_DATAPATH_bkp_3__7_), .R(rst_n_bF_buf78), .S(1'b1) );
  DFFSR DFFSR_445 ( .CLK(clk_bF_buf81), .D(AES_CORE_DATAPATH__0bkp_3__31_0__8_), .Q(AES_CORE_DATAPATH_bkp_3__8_), .R(rst_n_bF_buf77), .S(1'b1) );
  DFFSR DFFSR_446 ( .CLK(clk_bF_buf80), .D(AES_CORE_DATAPATH__0bkp_3__31_0__9_), .Q(AES_CORE_DATAPATH_bkp_3__9_), .R(rst_n_bF_buf76), .S(1'b1) );
  DFFSR DFFSR_447 ( .CLK(clk_bF_buf79), .D(AES_CORE_DATAPATH__0bkp_3__31_0__10_), .Q(AES_CORE_DATAPATH_bkp_3__10_), .R(rst_n_bF_buf75), .S(1'b1) );
  DFFSR DFFSR_448 ( .CLK(clk_bF_buf78), .D(AES_CORE_DATAPATH__0bkp_3__31_0__11_), .Q(AES_CORE_DATAPATH_bkp_3__11_), .R(rst_n_bF_buf74), .S(1'b1) );
  DFFSR DFFSR_449 ( .CLK(clk_bF_buf77), .D(AES_CORE_DATAPATH__0bkp_3__31_0__12_), .Q(AES_CORE_DATAPATH_bkp_3__12_), .R(rst_n_bF_buf73), .S(1'b1) );
  DFFSR DFFSR_45 ( .CLK(clk_bF_buf16), .D(AES_CORE_DATAPATH__0key_host_0__31_0__24_), .Q(AES_CORE_DATAPATH_key_host_0__24_), .R(rst_n_bF_buf42), .S(1'b1) );
  DFFSR DFFSR_450 ( .CLK(clk_bF_buf76), .D(AES_CORE_DATAPATH__0bkp_3__31_0__13_), .Q(AES_CORE_DATAPATH_bkp_3__13_), .R(rst_n_bF_buf72), .S(1'b1) );
  DFFSR DFFSR_451 ( .CLK(clk_bF_buf75), .D(AES_CORE_DATAPATH__0bkp_3__31_0__14_), .Q(AES_CORE_DATAPATH_bkp_3__14_), .R(rst_n_bF_buf71), .S(1'b1) );
  DFFSR DFFSR_452 ( .CLK(clk_bF_buf74), .D(AES_CORE_DATAPATH__0bkp_3__31_0__15_), .Q(AES_CORE_DATAPATH_bkp_3__15_), .R(rst_n_bF_buf70), .S(1'b1) );
  DFFSR DFFSR_453 ( .CLK(clk_bF_buf73), .D(AES_CORE_DATAPATH__0bkp_3__31_0__16_), .Q(AES_CORE_DATAPATH_bkp_3__16_), .R(rst_n_bF_buf69), .S(1'b1) );
  DFFSR DFFSR_454 ( .CLK(clk_bF_buf72), .D(AES_CORE_DATAPATH__0bkp_3__31_0__17_), .Q(AES_CORE_DATAPATH_bkp_3__17_), .R(rst_n_bF_buf68), .S(1'b1) );
  DFFSR DFFSR_455 ( .CLK(clk_bF_buf71), .D(AES_CORE_DATAPATH__0bkp_3__31_0__18_), .Q(AES_CORE_DATAPATH_bkp_3__18_), .R(rst_n_bF_buf67), .S(1'b1) );
  DFFSR DFFSR_456 ( .CLK(clk_bF_buf70), .D(AES_CORE_DATAPATH__0bkp_3__31_0__19_), .Q(AES_CORE_DATAPATH_bkp_3__19_), .R(rst_n_bF_buf66), .S(1'b1) );
  DFFSR DFFSR_457 ( .CLK(clk_bF_buf69), .D(AES_CORE_DATAPATH__0bkp_3__31_0__20_), .Q(AES_CORE_DATAPATH_bkp_3__20_), .R(rst_n_bF_buf65), .S(1'b1) );
  DFFSR DFFSR_458 ( .CLK(clk_bF_buf68), .D(AES_CORE_DATAPATH__0bkp_3__31_0__21_), .Q(AES_CORE_DATAPATH_bkp_3__21_), .R(rst_n_bF_buf64), .S(1'b1) );
  DFFSR DFFSR_459 ( .CLK(clk_bF_buf67), .D(AES_CORE_DATAPATH__0bkp_3__31_0__22_), .Q(AES_CORE_DATAPATH_bkp_3__22_), .R(rst_n_bF_buf63), .S(1'b1) );
  DFFSR DFFSR_46 ( .CLK(clk_bF_buf15), .D(AES_CORE_DATAPATH__0key_host_0__31_0__25_), .Q(AES_CORE_DATAPATH_key_host_0__25_), .R(rst_n_bF_buf41), .S(1'b1) );
  DFFSR DFFSR_460 ( .CLK(clk_bF_buf66), .D(AES_CORE_DATAPATH__0bkp_3__31_0__23_), .Q(AES_CORE_DATAPATH_bkp_3__23_), .R(rst_n_bF_buf62), .S(1'b1) );
  DFFSR DFFSR_461 ( .CLK(clk_bF_buf65), .D(AES_CORE_DATAPATH__0bkp_3__31_0__24_), .Q(AES_CORE_DATAPATH_bkp_3__24_), .R(rst_n_bF_buf61), .S(1'b1) );
  DFFSR DFFSR_462 ( .CLK(clk_bF_buf64), .D(AES_CORE_DATAPATH__0bkp_3__31_0__25_), .Q(AES_CORE_DATAPATH_bkp_3__25_), .R(rst_n_bF_buf60), .S(1'b1) );
  DFFSR DFFSR_463 ( .CLK(clk_bF_buf63), .D(AES_CORE_DATAPATH__0bkp_3__31_0__26_), .Q(AES_CORE_DATAPATH_bkp_3__26_), .R(rst_n_bF_buf59), .S(1'b1) );
  DFFSR DFFSR_464 ( .CLK(clk_bF_buf62), .D(AES_CORE_DATAPATH__0bkp_3__31_0__27_), .Q(AES_CORE_DATAPATH_bkp_3__27_), .R(rst_n_bF_buf58), .S(1'b1) );
  DFFSR DFFSR_465 ( .CLK(clk_bF_buf61), .D(AES_CORE_DATAPATH__0bkp_3__31_0__28_), .Q(AES_CORE_DATAPATH_bkp_3__28_), .R(rst_n_bF_buf57), .S(1'b1) );
  DFFSR DFFSR_466 ( .CLK(clk_bF_buf60), .D(AES_CORE_DATAPATH__0bkp_3__31_0__29_), .Q(AES_CORE_DATAPATH_bkp_3__29_), .R(rst_n_bF_buf56), .S(1'b1) );
  DFFSR DFFSR_467 ( .CLK(clk_bF_buf59), .D(AES_CORE_DATAPATH__0bkp_3__31_0__30_), .Q(AES_CORE_DATAPATH_bkp_3__30_), .R(rst_n_bF_buf55), .S(1'b1) );
  DFFSR DFFSR_468 ( .CLK(clk_bF_buf58), .D(AES_CORE_DATAPATH__0bkp_3__31_0__31_), .Q(AES_CORE_DATAPATH_bkp_3__31_), .R(rst_n_bF_buf54), .S(1'b1) );
  DFFSR DFFSR_469 ( .CLK(clk_bF_buf57), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__0_), .Q(AES_CORE_DATAPATH_bkp_1_3__0_), .R(rst_n_bF_buf53), .S(1'b1) );
  DFFSR DFFSR_47 ( .CLK(clk_bF_buf14), .D(AES_CORE_DATAPATH__0key_host_0__31_0__26_), .Q(AES_CORE_DATAPATH_key_host_0__26_), .R(rst_n_bF_buf40), .S(1'b1) );
  DFFSR DFFSR_470 ( .CLK(clk_bF_buf56), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__1_), .Q(AES_CORE_DATAPATH_bkp_1_3__1_), .R(rst_n_bF_buf52), .S(1'b1) );
  DFFSR DFFSR_471 ( .CLK(clk_bF_buf55), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__2_), .Q(AES_CORE_DATAPATH_bkp_1_3__2_), .R(rst_n_bF_buf51), .S(1'b1) );
  DFFSR DFFSR_472 ( .CLK(clk_bF_buf54), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__3_), .Q(AES_CORE_DATAPATH_bkp_1_3__3_), .R(rst_n_bF_buf50), .S(1'b1) );
  DFFSR DFFSR_473 ( .CLK(clk_bF_buf53), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__4_), .Q(AES_CORE_DATAPATH_bkp_1_3__4_), .R(rst_n_bF_buf49), .S(1'b1) );
  DFFSR DFFSR_474 ( .CLK(clk_bF_buf52), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__5_), .Q(AES_CORE_DATAPATH_bkp_1_3__5_), .R(rst_n_bF_buf48), .S(1'b1) );
  DFFSR DFFSR_475 ( .CLK(clk_bF_buf51), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__6_), .Q(AES_CORE_DATAPATH_bkp_1_3__6_), .R(rst_n_bF_buf47), .S(1'b1) );
  DFFSR DFFSR_476 ( .CLK(clk_bF_buf50), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__7_), .Q(AES_CORE_DATAPATH_bkp_1_3__7_), .R(rst_n_bF_buf46), .S(1'b1) );
  DFFSR DFFSR_477 ( .CLK(clk_bF_buf49), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__8_), .Q(AES_CORE_DATAPATH_bkp_1_3__8_), .R(rst_n_bF_buf45), .S(1'b1) );
  DFFSR DFFSR_478 ( .CLK(clk_bF_buf48), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__9_), .Q(AES_CORE_DATAPATH_bkp_1_3__9_), .R(rst_n_bF_buf44), .S(1'b1) );
  DFFSR DFFSR_479 ( .CLK(clk_bF_buf47), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__10_), .Q(AES_CORE_DATAPATH_bkp_1_3__10_), .R(rst_n_bF_buf43), .S(1'b1) );
  DFFSR DFFSR_48 ( .CLK(clk_bF_buf13), .D(AES_CORE_DATAPATH__0key_host_0__31_0__27_), .Q(AES_CORE_DATAPATH_key_host_0__27_), .R(rst_n_bF_buf39), .S(1'b1) );
  DFFSR DFFSR_480 ( .CLK(clk_bF_buf46), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__11_), .Q(AES_CORE_DATAPATH_bkp_1_3__11_), .R(rst_n_bF_buf42), .S(1'b1) );
  DFFSR DFFSR_481 ( .CLK(clk_bF_buf45), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__12_), .Q(AES_CORE_DATAPATH_bkp_1_3__12_), .R(rst_n_bF_buf41), .S(1'b1) );
  DFFSR DFFSR_482 ( .CLK(clk_bF_buf44), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__13_), .Q(AES_CORE_DATAPATH_bkp_1_3__13_), .R(rst_n_bF_buf40), .S(1'b1) );
  DFFSR DFFSR_483 ( .CLK(clk_bF_buf43), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__14_), .Q(AES_CORE_DATAPATH_bkp_1_3__14_), .R(rst_n_bF_buf39), .S(1'b1) );
  DFFSR DFFSR_484 ( .CLK(clk_bF_buf42), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__15_), .Q(AES_CORE_DATAPATH_bkp_1_3__15_), .R(rst_n_bF_buf38), .S(1'b1) );
  DFFSR DFFSR_485 ( .CLK(clk_bF_buf41), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__16_), .Q(AES_CORE_DATAPATH_bkp_1_3__16_), .R(rst_n_bF_buf37), .S(1'b1) );
  DFFSR DFFSR_486 ( .CLK(clk_bF_buf40), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__17_), .Q(AES_CORE_DATAPATH_bkp_1_3__17_), .R(rst_n_bF_buf36), .S(1'b1) );
  DFFSR DFFSR_487 ( .CLK(clk_bF_buf39), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__18_), .Q(AES_CORE_DATAPATH_bkp_1_3__18_), .R(rst_n_bF_buf35), .S(1'b1) );
  DFFSR DFFSR_488 ( .CLK(clk_bF_buf38), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__19_), .Q(AES_CORE_DATAPATH_bkp_1_3__19_), .R(rst_n_bF_buf34), .S(1'b1) );
  DFFSR DFFSR_489 ( .CLK(clk_bF_buf37), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__20_), .Q(AES_CORE_DATAPATH_bkp_1_3__20_), .R(rst_n_bF_buf33), .S(1'b1) );
  DFFSR DFFSR_49 ( .CLK(clk_bF_buf12), .D(AES_CORE_DATAPATH__0key_host_0__31_0__28_), .Q(AES_CORE_DATAPATH_key_host_0__28_), .R(rst_n_bF_buf38), .S(1'b1) );
  DFFSR DFFSR_490 ( .CLK(clk_bF_buf36), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__21_), .Q(AES_CORE_DATAPATH_bkp_1_3__21_), .R(rst_n_bF_buf32), .S(1'b1) );
  DFFSR DFFSR_491 ( .CLK(clk_bF_buf35), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__22_), .Q(AES_CORE_DATAPATH_bkp_1_3__22_), .R(rst_n_bF_buf31), .S(1'b1) );
  DFFSR DFFSR_492 ( .CLK(clk_bF_buf34), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__23_), .Q(AES_CORE_DATAPATH_bkp_1_3__23_), .R(rst_n_bF_buf30), .S(1'b1) );
  DFFSR DFFSR_493 ( .CLK(clk_bF_buf33), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__24_), .Q(AES_CORE_DATAPATH_bkp_1_3__24_), .R(rst_n_bF_buf29), .S(1'b1) );
  DFFSR DFFSR_494 ( .CLK(clk_bF_buf32), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__25_), .Q(AES_CORE_DATAPATH_bkp_1_3__25_), .R(rst_n_bF_buf28), .S(1'b1) );
  DFFSR DFFSR_495 ( .CLK(clk_bF_buf31), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__26_), .Q(AES_CORE_DATAPATH_bkp_1_3__26_), .R(rst_n_bF_buf27), .S(1'b1) );
  DFFSR DFFSR_496 ( .CLK(clk_bF_buf30), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__27_), .Q(AES_CORE_DATAPATH_bkp_1_3__27_), .R(rst_n_bF_buf26), .S(1'b1) );
  DFFSR DFFSR_497 ( .CLK(clk_bF_buf29), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__28_), .Q(AES_CORE_DATAPATH_bkp_1_3__28_), .R(rst_n_bF_buf25), .S(1'b1) );
  DFFSR DFFSR_498 ( .CLK(clk_bF_buf28), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__29_), .Q(AES_CORE_DATAPATH_bkp_1_3__29_), .R(rst_n_bF_buf24), .S(1'b1) );
  DFFSR DFFSR_499 ( .CLK(clk_bF_buf27), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__30_), .Q(AES_CORE_DATAPATH_bkp_1_3__30_), .R(rst_n_bF_buf23), .S(1'b1) );
  DFFSR DFFSR_5 ( .CLK(clk_bF_buf88), .D(AES_CORE_CONTROL_UNIT__abc_10818_n59), .Q(AES_CORE_CONTROL_UNIT_state_0_), .R(1'b1), .S(rst_n_bF_buf82) );
  DFFSR DFFSR_50 ( .CLK(clk_bF_buf11), .D(AES_CORE_DATAPATH__0key_host_0__31_0__29_), .Q(AES_CORE_DATAPATH_key_host_0__29_), .R(rst_n_bF_buf37), .S(1'b1) );
  DFFSR DFFSR_500 ( .CLK(clk_bF_buf26), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__31_), .Q(AES_CORE_DATAPATH_bkp_1_3__31_), .R(rst_n_bF_buf22), .S(1'b1) );
  DFFSR DFFSR_501 ( .CLK(clk_bF_buf25), .D(AES_CORE_DATAPATH__0iv_2__31_0__0_), .Q(AES_CORE_DATAPATH_iv_2__0_), .R(rst_n_bF_buf21), .S(1'b1) );
  DFFSR DFFSR_502 ( .CLK(clk_bF_buf24), .D(AES_CORE_DATAPATH__0iv_2__31_0__1_), .Q(AES_CORE_DATAPATH_iv_2__1_), .R(rst_n_bF_buf20), .S(1'b1) );
  DFFSR DFFSR_503 ( .CLK(clk_bF_buf23), .D(AES_CORE_DATAPATH__0iv_2__31_0__2_), .Q(AES_CORE_DATAPATH_iv_2__2_), .R(rst_n_bF_buf19), .S(1'b1) );
  DFFSR DFFSR_504 ( .CLK(clk_bF_buf22), .D(AES_CORE_DATAPATH__0iv_2__31_0__3_), .Q(AES_CORE_DATAPATH_iv_2__3_), .R(rst_n_bF_buf18), .S(1'b1) );
  DFFSR DFFSR_505 ( .CLK(clk_bF_buf21), .D(AES_CORE_DATAPATH__0iv_2__31_0__4_), .Q(AES_CORE_DATAPATH_iv_2__4_), .R(rst_n_bF_buf17), .S(1'b1) );
  DFFSR DFFSR_506 ( .CLK(clk_bF_buf20), .D(AES_CORE_DATAPATH__0iv_2__31_0__5_), .Q(AES_CORE_DATAPATH_iv_2__5_), .R(rst_n_bF_buf16), .S(1'b1) );
  DFFSR DFFSR_507 ( .CLK(clk_bF_buf19), .D(AES_CORE_DATAPATH__0iv_2__31_0__6_), .Q(AES_CORE_DATAPATH_iv_2__6_), .R(rst_n_bF_buf15), .S(1'b1) );
  DFFSR DFFSR_508 ( .CLK(clk_bF_buf18), .D(AES_CORE_DATAPATH__0iv_2__31_0__7_), .Q(AES_CORE_DATAPATH_iv_2__7_), .R(rst_n_bF_buf14), .S(1'b1) );
  DFFSR DFFSR_509 ( .CLK(clk_bF_buf17), .D(AES_CORE_DATAPATH__0iv_2__31_0__8_), .Q(AES_CORE_DATAPATH_iv_2__8_), .R(rst_n_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_51 ( .CLK(clk_bF_buf10), .D(AES_CORE_DATAPATH__0key_host_0__31_0__30_), .Q(AES_CORE_DATAPATH_key_host_0__30_), .R(rst_n_bF_buf36), .S(1'b1) );
  DFFSR DFFSR_510 ( .CLK(clk_bF_buf16), .D(AES_CORE_DATAPATH__0iv_2__31_0__9_), .Q(AES_CORE_DATAPATH_iv_2__9_), .R(rst_n_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_511 ( .CLK(clk_bF_buf15), .D(AES_CORE_DATAPATH__0iv_2__31_0__10_), .Q(AES_CORE_DATAPATH_iv_2__10_), .R(rst_n_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_512 ( .CLK(clk_bF_buf14), .D(AES_CORE_DATAPATH__0iv_2__31_0__11_), .Q(AES_CORE_DATAPATH_iv_2__11_), .R(rst_n_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_513 ( .CLK(clk_bF_buf13), .D(AES_CORE_DATAPATH__0iv_2__31_0__12_), .Q(AES_CORE_DATAPATH_iv_2__12_), .R(rst_n_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_514 ( .CLK(clk_bF_buf12), .D(AES_CORE_DATAPATH__0iv_2__31_0__13_), .Q(AES_CORE_DATAPATH_iv_2__13_), .R(rst_n_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_515 ( .CLK(clk_bF_buf11), .D(AES_CORE_DATAPATH__0iv_2__31_0__14_), .Q(AES_CORE_DATAPATH_iv_2__14_), .R(rst_n_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_516 ( .CLK(clk_bF_buf10), .D(AES_CORE_DATAPATH__0iv_2__31_0__15_), .Q(AES_CORE_DATAPATH_iv_2__15_), .R(rst_n_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_517 ( .CLK(clk_bF_buf9), .D(AES_CORE_DATAPATH__0iv_2__31_0__16_), .Q(AES_CORE_DATAPATH_iv_2__16_), .R(rst_n_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_518 ( .CLK(clk_bF_buf8), .D(AES_CORE_DATAPATH__0iv_2__31_0__17_), .Q(AES_CORE_DATAPATH_iv_2__17_), .R(rst_n_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_519 ( .CLK(clk_bF_buf7), .D(AES_CORE_DATAPATH__0iv_2__31_0__18_), .Q(AES_CORE_DATAPATH_iv_2__18_), .R(rst_n_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_52 ( .CLK(clk_bF_buf9), .D(AES_CORE_DATAPATH__0key_host_0__31_0__31_), .Q(AES_CORE_DATAPATH_key_host_0__31_), .R(rst_n_bF_buf35), .S(1'b1) );
  DFFSR DFFSR_520 ( .CLK(clk_bF_buf6), .D(AES_CORE_DATAPATH__0iv_2__31_0__19_), .Q(AES_CORE_DATAPATH_iv_2__19_), .R(rst_n_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_521 ( .CLK(clk_bF_buf5), .D(AES_CORE_DATAPATH__0iv_2__31_0__20_), .Q(AES_CORE_DATAPATH_iv_2__20_), .R(rst_n_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_522 ( .CLK(clk_bF_buf4), .D(AES_CORE_DATAPATH__0iv_2__31_0__21_), .Q(AES_CORE_DATAPATH_iv_2__21_), .R(rst_n_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_523 ( .CLK(clk_bF_buf3), .D(AES_CORE_DATAPATH__0iv_2__31_0__22_), .Q(AES_CORE_DATAPATH_iv_2__22_), .R(rst_n_bF_buf86), .S(1'b1) );
  DFFSR DFFSR_524 ( .CLK(clk_bF_buf2), .D(AES_CORE_DATAPATH__0iv_2__31_0__23_), .Q(AES_CORE_DATAPATH_iv_2__23_), .R(rst_n_bF_buf85), .S(1'b1) );
  DFFSR DFFSR_525 ( .CLK(clk_bF_buf1), .D(AES_CORE_DATAPATH__0iv_2__31_0__24_), .Q(AES_CORE_DATAPATH_iv_2__24_), .R(rst_n_bF_buf84), .S(1'b1) );
  DFFSR DFFSR_526 ( .CLK(clk_bF_buf0), .D(AES_CORE_DATAPATH__0iv_2__31_0__25_), .Q(AES_CORE_DATAPATH_iv_2__25_), .R(rst_n_bF_buf83), .S(1'b1) );
  DFFSR DFFSR_527 ( .CLK(clk_bF_buf92), .D(AES_CORE_DATAPATH__0iv_2__31_0__26_), .Q(AES_CORE_DATAPATH_iv_2__26_), .R(rst_n_bF_buf82), .S(1'b1) );
  DFFSR DFFSR_528 ( .CLK(clk_bF_buf91), .D(AES_CORE_DATAPATH__0iv_2__31_0__27_), .Q(AES_CORE_DATAPATH_iv_2__27_), .R(rst_n_bF_buf81), .S(1'b1) );
  DFFSR DFFSR_529 ( .CLK(clk_bF_buf90), .D(AES_CORE_DATAPATH__0iv_2__31_0__28_), .Q(AES_CORE_DATAPATH_iv_2__28_), .R(rst_n_bF_buf80), .S(1'b1) );
  DFFSR DFFSR_53 ( .CLK(clk_bF_buf8), .D(AES_CORE_DATAPATH__0key_0__31_0__0_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__0_), .R(rst_n_bF_buf34), .S(1'b1) );
  DFFSR DFFSR_530 ( .CLK(clk_bF_buf89), .D(AES_CORE_DATAPATH__0iv_2__31_0__29_), .Q(AES_CORE_DATAPATH_iv_2__29_), .R(rst_n_bF_buf79), .S(1'b1) );
  DFFSR DFFSR_531 ( .CLK(clk_bF_buf88), .D(AES_CORE_DATAPATH__0iv_2__31_0__30_), .Q(AES_CORE_DATAPATH_iv_2__30_), .R(rst_n_bF_buf78), .S(1'b1) );
  DFFSR DFFSR_532 ( .CLK(clk_bF_buf87), .D(AES_CORE_DATAPATH__0iv_2__31_0__31_), .Q(AES_CORE_DATAPATH_iv_2__31_), .R(rst_n_bF_buf77), .S(1'b1) );
  DFFSR DFFSR_533 ( .CLK(clk_bF_buf86), .D(AES_CORE_DATAPATH__0bkp_2__31_0__0_), .Q(AES_CORE_DATAPATH_bkp_2__0_), .R(rst_n_bF_buf76), .S(1'b1) );
  DFFSR DFFSR_534 ( .CLK(clk_bF_buf85), .D(AES_CORE_DATAPATH__0bkp_2__31_0__1_), .Q(AES_CORE_DATAPATH_bkp_2__1_), .R(rst_n_bF_buf75), .S(1'b1) );
  DFFSR DFFSR_535 ( .CLK(clk_bF_buf84), .D(AES_CORE_DATAPATH__0bkp_2__31_0__2_), .Q(AES_CORE_DATAPATH_bkp_2__2_), .R(rst_n_bF_buf74), .S(1'b1) );
  DFFSR DFFSR_536 ( .CLK(clk_bF_buf83), .D(AES_CORE_DATAPATH__0bkp_2__31_0__3_), .Q(AES_CORE_DATAPATH_bkp_2__3_), .R(rst_n_bF_buf73), .S(1'b1) );
  DFFSR DFFSR_537 ( .CLK(clk_bF_buf82), .D(AES_CORE_DATAPATH__0bkp_2__31_0__4_), .Q(AES_CORE_DATAPATH_bkp_2__4_), .R(rst_n_bF_buf72), .S(1'b1) );
  DFFSR DFFSR_538 ( .CLK(clk_bF_buf81), .D(AES_CORE_DATAPATH__0bkp_2__31_0__5_), .Q(AES_CORE_DATAPATH_bkp_2__5_), .R(rst_n_bF_buf71), .S(1'b1) );
  DFFSR DFFSR_539 ( .CLK(clk_bF_buf80), .D(AES_CORE_DATAPATH__0bkp_2__31_0__6_), .Q(AES_CORE_DATAPATH_bkp_2__6_), .R(rst_n_bF_buf70), .S(1'b1) );
  DFFSR DFFSR_54 ( .CLK(clk_bF_buf7), .D(AES_CORE_DATAPATH__0key_0__31_0__1_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__1_), .R(rst_n_bF_buf33), .S(1'b1) );
  DFFSR DFFSR_540 ( .CLK(clk_bF_buf79), .D(AES_CORE_DATAPATH__0bkp_2__31_0__7_), .Q(AES_CORE_DATAPATH_bkp_2__7_), .R(rst_n_bF_buf69), .S(1'b1) );
  DFFSR DFFSR_541 ( .CLK(clk_bF_buf78), .D(AES_CORE_DATAPATH__0bkp_2__31_0__8_), .Q(AES_CORE_DATAPATH_bkp_2__8_), .R(rst_n_bF_buf68), .S(1'b1) );
  DFFSR DFFSR_542 ( .CLK(clk_bF_buf77), .D(AES_CORE_DATAPATH__0bkp_2__31_0__9_), .Q(AES_CORE_DATAPATH_bkp_2__9_), .R(rst_n_bF_buf67), .S(1'b1) );
  DFFSR DFFSR_543 ( .CLK(clk_bF_buf76), .D(AES_CORE_DATAPATH__0bkp_2__31_0__10_), .Q(AES_CORE_DATAPATH_bkp_2__10_), .R(rst_n_bF_buf66), .S(1'b1) );
  DFFSR DFFSR_544 ( .CLK(clk_bF_buf75), .D(AES_CORE_DATAPATH__0bkp_2__31_0__11_), .Q(AES_CORE_DATAPATH_bkp_2__11_), .R(rst_n_bF_buf65), .S(1'b1) );
  DFFSR DFFSR_545 ( .CLK(clk_bF_buf74), .D(AES_CORE_DATAPATH__0bkp_2__31_0__12_), .Q(AES_CORE_DATAPATH_bkp_2__12_), .R(rst_n_bF_buf64), .S(1'b1) );
  DFFSR DFFSR_546 ( .CLK(clk_bF_buf73), .D(AES_CORE_DATAPATH__0bkp_2__31_0__13_), .Q(AES_CORE_DATAPATH_bkp_2__13_), .R(rst_n_bF_buf63), .S(1'b1) );
  DFFSR DFFSR_547 ( .CLK(clk_bF_buf72), .D(AES_CORE_DATAPATH__0bkp_2__31_0__14_), .Q(AES_CORE_DATAPATH_bkp_2__14_), .R(rst_n_bF_buf62), .S(1'b1) );
  DFFSR DFFSR_548 ( .CLK(clk_bF_buf71), .D(AES_CORE_DATAPATH__0bkp_2__31_0__15_), .Q(AES_CORE_DATAPATH_bkp_2__15_), .R(rst_n_bF_buf61), .S(1'b1) );
  DFFSR DFFSR_549 ( .CLK(clk_bF_buf70), .D(AES_CORE_DATAPATH__0bkp_2__31_0__16_), .Q(AES_CORE_DATAPATH_bkp_2__16_), .R(rst_n_bF_buf60), .S(1'b1) );
  DFFSR DFFSR_55 ( .CLK(clk_bF_buf6), .D(AES_CORE_DATAPATH__0key_0__31_0__2_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__2_), .R(rst_n_bF_buf32), .S(1'b1) );
  DFFSR DFFSR_550 ( .CLK(clk_bF_buf69), .D(AES_CORE_DATAPATH__0bkp_2__31_0__17_), .Q(AES_CORE_DATAPATH_bkp_2__17_), .R(rst_n_bF_buf59), .S(1'b1) );
  DFFSR DFFSR_551 ( .CLK(clk_bF_buf68), .D(AES_CORE_DATAPATH__0bkp_2__31_0__18_), .Q(AES_CORE_DATAPATH_bkp_2__18_), .R(rst_n_bF_buf58), .S(1'b1) );
  DFFSR DFFSR_552 ( .CLK(clk_bF_buf67), .D(AES_CORE_DATAPATH__0bkp_2__31_0__19_), .Q(AES_CORE_DATAPATH_bkp_2__19_), .R(rst_n_bF_buf57), .S(1'b1) );
  DFFSR DFFSR_553 ( .CLK(clk_bF_buf66), .D(AES_CORE_DATAPATH__0bkp_2__31_0__20_), .Q(AES_CORE_DATAPATH_bkp_2__20_), .R(rst_n_bF_buf56), .S(1'b1) );
  DFFSR DFFSR_554 ( .CLK(clk_bF_buf65), .D(AES_CORE_DATAPATH__0bkp_2__31_0__21_), .Q(AES_CORE_DATAPATH_bkp_2__21_), .R(rst_n_bF_buf55), .S(1'b1) );
  DFFSR DFFSR_555 ( .CLK(clk_bF_buf64), .D(AES_CORE_DATAPATH__0bkp_2__31_0__22_), .Q(AES_CORE_DATAPATH_bkp_2__22_), .R(rst_n_bF_buf54), .S(1'b1) );
  DFFSR DFFSR_556 ( .CLK(clk_bF_buf63), .D(AES_CORE_DATAPATH__0bkp_2__31_0__23_), .Q(AES_CORE_DATAPATH_bkp_2__23_), .R(rst_n_bF_buf53), .S(1'b1) );
  DFFSR DFFSR_557 ( .CLK(clk_bF_buf62), .D(AES_CORE_DATAPATH__0bkp_2__31_0__24_), .Q(AES_CORE_DATAPATH_bkp_2__24_), .R(rst_n_bF_buf52), .S(1'b1) );
  DFFSR DFFSR_558 ( .CLK(clk_bF_buf61), .D(AES_CORE_DATAPATH__0bkp_2__31_0__25_), .Q(AES_CORE_DATAPATH_bkp_2__25_), .R(rst_n_bF_buf51), .S(1'b1) );
  DFFSR DFFSR_559 ( .CLK(clk_bF_buf60), .D(AES_CORE_DATAPATH__0bkp_2__31_0__26_), .Q(AES_CORE_DATAPATH_bkp_2__26_), .R(rst_n_bF_buf50), .S(1'b1) );
  DFFSR DFFSR_56 ( .CLK(clk_bF_buf5), .D(AES_CORE_DATAPATH__0key_0__31_0__3_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__3_), .R(rst_n_bF_buf31), .S(1'b1) );
  DFFSR DFFSR_560 ( .CLK(clk_bF_buf59), .D(AES_CORE_DATAPATH__0bkp_2__31_0__27_), .Q(AES_CORE_DATAPATH_bkp_2__27_), .R(rst_n_bF_buf49), .S(1'b1) );
  DFFSR DFFSR_561 ( .CLK(clk_bF_buf58), .D(AES_CORE_DATAPATH__0bkp_2__31_0__28_), .Q(AES_CORE_DATAPATH_bkp_2__28_), .R(rst_n_bF_buf48), .S(1'b1) );
  DFFSR DFFSR_562 ( .CLK(clk_bF_buf57), .D(AES_CORE_DATAPATH__0bkp_2__31_0__29_), .Q(AES_CORE_DATAPATH_bkp_2__29_), .R(rst_n_bF_buf47), .S(1'b1) );
  DFFSR DFFSR_563 ( .CLK(clk_bF_buf56), .D(AES_CORE_DATAPATH__0bkp_2__31_0__30_), .Q(AES_CORE_DATAPATH_bkp_2__30_), .R(rst_n_bF_buf46), .S(1'b1) );
  DFFSR DFFSR_564 ( .CLK(clk_bF_buf55), .D(AES_CORE_DATAPATH__0bkp_2__31_0__31_), .Q(AES_CORE_DATAPATH_bkp_2__31_), .R(rst_n_bF_buf45), .S(1'b1) );
  DFFSR DFFSR_565 ( .CLK(clk_bF_buf54), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__0_), .Q(AES_CORE_DATAPATH_bkp_1_2__0_), .R(rst_n_bF_buf44), .S(1'b1) );
  DFFSR DFFSR_566 ( .CLK(clk_bF_buf53), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__1_), .Q(AES_CORE_DATAPATH_bkp_1_2__1_), .R(rst_n_bF_buf43), .S(1'b1) );
  DFFSR DFFSR_567 ( .CLK(clk_bF_buf52), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__2_), .Q(AES_CORE_DATAPATH_bkp_1_2__2_), .R(rst_n_bF_buf42), .S(1'b1) );
  DFFSR DFFSR_568 ( .CLK(clk_bF_buf51), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__3_), .Q(AES_CORE_DATAPATH_bkp_1_2__3_), .R(rst_n_bF_buf41), .S(1'b1) );
  DFFSR DFFSR_569 ( .CLK(clk_bF_buf50), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__4_), .Q(AES_CORE_DATAPATH_bkp_1_2__4_), .R(rst_n_bF_buf40), .S(1'b1) );
  DFFSR DFFSR_57 ( .CLK(clk_bF_buf4), .D(AES_CORE_DATAPATH__0key_0__31_0__4_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__4_), .R(rst_n_bF_buf30), .S(1'b1) );
  DFFSR DFFSR_570 ( .CLK(clk_bF_buf49), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__5_), .Q(AES_CORE_DATAPATH_bkp_1_2__5_), .R(rst_n_bF_buf39), .S(1'b1) );
  DFFSR DFFSR_571 ( .CLK(clk_bF_buf48), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__6_), .Q(AES_CORE_DATAPATH_bkp_1_2__6_), .R(rst_n_bF_buf38), .S(1'b1) );
  DFFSR DFFSR_572 ( .CLK(clk_bF_buf47), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__7_), .Q(AES_CORE_DATAPATH_bkp_1_2__7_), .R(rst_n_bF_buf37), .S(1'b1) );
  DFFSR DFFSR_573 ( .CLK(clk_bF_buf46), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__8_), .Q(AES_CORE_DATAPATH_bkp_1_2__8_), .R(rst_n_bF_buf36), .S(1'b1) );
  DFFSR DFFSR_574 ( .CLK(clk_bF_buf45), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__9_), .Q(AES_CORE_DATAPATH_bkp_1_2__9_), .R(rst_n_bF_buf35), .S(1'b1) );
  DFFSR DFFSR_575 ( .CLK(clk_bF_buf44), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__10_), .Q(AES_CORE_DATAPATH_bkp_1_2__10_), .R(rst_n_bF_buf34), .S(1'b1) );
  DFFSR DFFSR_576 ( .CLK(clk_bF_buf43), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__11_), .Q(AES_CORE_DATAPATH_bkp_1_2__11_), .R(rst_n_bF_buf33), .S(1'b1) );
  DFFSR DFFSR_577 ( .CLK(clk_bF_buf42), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__12_), .Q(AES_CORE_DATAPATH_bkp_1_2__12_), .R(rst_n_bF_buf32), .S(1'b1) );
  DFFSR DFFSR_578 ( .CLK(clk_bF_buf41), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__13_), .Q(AES_CORE_DATAPATH_bkp_1_2__13_), .R(rst_n_bF_buf31), .S(1'b1) );
  DFFSR DFFSR_579 ( .CLK(clk_bF_buf40), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__14_), .Q(AES_CORE_DATAPATH_bkp_1_2__14_), .R(rst_n_bF_buf30), .S(1'b1) );
  DFFSR DFFSR_58 ( .CLK(clk_bF_buf3), .D(AES_CORE_DATAPATH__0key_0__31_0__5_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__5_), .R(rst_n_bF_buf29), .S(1'b1) );
  DFFSR DFFSR_580 ( .CLK(clk_bF_buf39), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__15_), .Q(AES_CORE_DATAPATH_bkp_1_2__15_), .R(rst_n_bF_buf29), .S(1'b1) );
  DFFSR DFFSR_581 ( .CLK(clk_bF_buf38), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__16_), .Q(AES_CORE_DATAPATH_bkp_1_2__16_), .R(rst_n_bF_buf28), .S(1'b1) );
  DFFSR DFFSR_582 ( .CLK(clk_bF_buf37), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__17_), .Q(AES_CORE_DATAPATH_bkp_1_2__17_), .R(rst_n_bF_buf27), .S(1'b1) );
  DFFSR DFFSR_583 ( .CLK(clk_bF_buf36), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__18_), .Q(AES_CORE_DATAPATH_bkp_1_2__18_), .R(rst_n_bF_buf26), .S(1'b1) );
  DFFSR DFFSR_584 ( .CLK(clk_bF_buf35), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__19_), .Q(AES_CORE_DATAPATH_bkp_1_2__19_), .R(rst_n_bF_buf25), .S(1'b1) );
  DFFSR DFFSR_585 ( .CLK(clk_bF_buf34), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__20_), .Q(AES_CORE_DATAPATH_bkp_1_2__20_), .R(rst_n_bF_buf24), .S(1'b1) );
  DFFSR DFFSR_586 ( .CLK(clk_bF_buf33), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__21_), .Q(AES_CORE_DATAPATH_bkp_1_2__21_), .R(rst_n_bF_buf23), .S(1'b1) );
  DFFSR DFFSR_587 ( .CLK(clk_bF_buf32), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__22_), .Q(AES_CORE_DATAPATH_bkp_1_2__22_), .R(rst_n_bF_buf22), .S(1'b1) );
  DFFSR DFFSR_588 ( .CLK(clk_bF_buf31), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__23_), .Q(AES_CORE_DATAPATH_bkp_1_2__23_), .R(rst_n_bF_buf21), .S(1'b1) );
  DFFSR DFFSR_589 ( .CLK(clk_bF_buf30), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__24_), .Q(AES_CORE_DATAPATH_bkp_1_2__24_), .R(rst_n_bF_buf20), .S(1'b1) );
  DFFSR DFFSR_59 ( .CLK(clk_bF_buf2), .D(AES_CORE_DATAPATH__0key_0__31_0__6_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__6_), .R(rst_n_bF_buf28), .S(1'b1) );
  DFFSR DFFSR_590 ( .CLK(clk_bF_buf29), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__25_), .Q(AES_CORE_DATAPATH_bkp_1_2__25_), .R(rst_n_bF_buf19), .S(1'b1) );
  DFFSR DFFSR_591 ( .CLK(clk_bF_buf28), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__26_), .Q(AES_CORE_DATAPATH_bkp_1_2__26_), .R(rst_n_bF_buf18), .S(1'b1) );
  DFFSR DFFSR_592 ( .CLK(clk_bF_buf27), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__27_), .Q(AES_CORE_DATAPATH_bkp_1_2__27_), .R(rst_n_bF_buf17), .S(1'b1) );
  DFFSR DFFSR_593 ( .CLK(clk_bF_buf26), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__28_), .Q(AES_CORE_DATAPATH_bkp_1_2__28_), .R(rst_n_bF_buf16), .S(1'b1) );
  DFFSR DFFSR_594 ( .CLK(clk_bF_buf25), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__29_), .Q(AES_CORE_DATAPATH_bkp_1_2__29_), .R(rst_n_bF_buf15), .S(1'b1) );
  DFFSR DFFSR_595 ( .CLK(clk_bF_buf24), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__30_), .Q(AES_CORE_DATAPATH_bkp_1_2__30_), .R(rst_n_bF_buf14), .S(1'b1) );
  DFFSR DFFSR_596 ( .CLK(clk_bF_buf23), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__31_), .Q(AES_CORE_DATAPATH_bkp_1_2__31_), .R(rst_n_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_597 ( .CLK(clk_bF_buf22), .D(AES_CORE_DATAPATH__0iv_1__31_0__0_), .Q(AES_CORE_DATAPATH_iv_1__0_), .R(rst_n_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_598 ( .CLK(clk_bF_buf21), .D(AES_CORE_DATAPATH__0iv_1__31_0__1_), .Q(AES_CORE_DATAPATH_iv_1__1_), .R(rst_n_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_599 ( .CLK(clk_bF_buf20), .D(AES_CORE_DATAPATH__0iv_1__31_0__2_), .Q(AES_CORE_DATAPATH_iv_1__2_), .R(rst_n_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_6 ( .CLK(clk_bF_buf87), .D(AES_CORE_CONTROL_UNIT__abc_10818_n24), .Q(AES_CORE_CONTROL_UNIT_state_1_), .R(rst_n_bF_buf81), .S(1'b1) );
  DFFSR DFFSR_60 ( .CLK(clk_bF_buf1), .D(AES_CORE_DATAPATH__0key_0__31_0__7_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__7_), .R(rst_n_bF_buf27), .S(1'b1) );
  DFFSR DFFSR_600 ( .CLK(clk_bF_buf19), .D(AES_CORE_DATAPATH__0iv_1__31_0__3_), .Q(AES_CORE_DATAPATH_iv_1__3_), .R(rst_n_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_601 ( .CLK(clk_bF_buf18), .D(AES_CORE_DATAPATH__0iv_1__31_0__4_), .Q(AES_CORE_DATAPATH_iv_1__4_), .R(rst_n_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_602 ( .CLK(clk_bF_buf17), .D(AES_CORE_DATAPATH__0iv_1__31_0__5_), .Q(AES_CORE_DATAPATH_iv_1__5_), .R(rst_n_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_603 ( .CLK(clk_bF_buf16), .D(AES_CORE_DATAPATH__0iv_1__31_0__6_), .Q(AES_CORE_DATAPATH_iv_1__6_), .R(rst_n_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_604 ( .CLK(clk_bF_buf15), .D(AES_CORE_DATAPATH__0iv_1__31_0__7_), .Q(AES_CORE_DATAPATH_iv_1__7_), .R(rst_n_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_605 ( .CLK(clk_bF_buf14), .D(AES_CORE_DATAPATH__0iv_1__31_0__8_), .Q(AES_CORE_DATAPATH_iv_1__8_), .R(rst_n_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_606 ( .CLK(clk_bF_buf13), .D(AES_CORE_DATAPATH__0iv_1__31_0__9_), .Q(AES_CORE_DATAPATH_iv_1__9_), .R(rst_n_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_607 ( .CLK(clk_bF_buf12), .D(AES_CORE_DATAPATH__0iv_1__31_0__10_), .Q(AES_CORE_DATAPATH_iv_1__10_), .R(rst_n_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_608 ( .CLK(clk_bF_buf11), .D(AES_CORE_DATAPATH__0iv_1__31_0__11_), .Q(AES_CORE_DATAPATH_iv_1__11_), .R(rst_n_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_609 ( .CLK(clk_bF_buf10), .D(AES_CORE_DATAPATH__0iv_1__31_0__12_), .Q(AES_CORE_DATAPATH_iv_1__12_), .R(rst_n_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_61 ( .CLK(clk_bF_buf0), .D(AES_CORE_DATAPATH__0key_0__31_0__8_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__8_), .R(rst_n_bF_buf26), .S(1'b1) );
  DFFSR DFFSR_610 ( .CLK(clk_bF_buf9), .D(AES_CORE_DATAPATH__0iv_1__31_0__13_), .Q(AES_CORE_DATAPATH_iv_1__13_), .R(rst_n_bF_buf86), .S(1'b1) );
  DFFSR DFFSR_611 ( .CLK(clk_bF_buf8), .D(AES_CORE_DATAPATH__0iv_1__31_0__14_), .Q(AES_CORE_DATAPATH_iv_1__14_), .R(rst_n_bF_buf85), .S(1'b1) );
  DFFSR DFFSR_612 ( .CLK(clk_bF_buf7), .D(AES_CORE_DATAPATH__0iv_1__31_0__15_), .Q(AES_CORE_DATAPATH_iv_1__15_), .R(rst_n_bF_buf84), .S(1'b1) );
  DFFSR DFFSR_613 ( .CLK(clk_bF_buf6), .D(AES_CORE_DATAPATH__0iv_1__31_0__16_), .Q(AES_CORE_DATAPATH_iv_1__16_), .R(rst_n_bF_buf83), .S(1'b1) );
  DFFSR DFFSR_614 ( .CLK(clk_bF_buf5), .D(AES_CORE_DATAPATH__0iv_1__31_0__17_), .Q(AES_CORE_DATAPATH_iv_1__17_), .R(rst_n_bF_buf82), .S(1'b1) );
  DFFSR DFFSR_615 ( .CLK(clk_bF_buf4), .D(AES_CORE_DATAPATH__0iv_1__31_0__18_), .Q(AES_CORE_DATAPATH_iv_1__18_), .R(rst_n_bF_buf81), .S(1'b1) );
  DFFSR DFFSR_616 ( .CLK(clk_bF_buf3), .D(AES_CORE_DATAPATH__0iv_1__31_0__19_), .Q(AES_CORE_DATAPATH_iv_1__19_), .R(rst_n_bF_buf80), .S(1'b1) );
  DFFSR DFFSR_617 ( .CLK(clk_bF_buf2), .D(AES_CORE_DATAPATH__0iv_1__31_0__20_), .Q(AES_CORE_DATAPATH_iv_1__20_), .R(rst_n_bF_buf79), .S(1'b1) );
  DFFSR DFFSR_618 ( .CLK(clk_bF_buf1), .D(AES_CORE_DATAPATH__0iv_1__31_0__21_), .Q(AES_CORE_DATAPATH_iv_1__21_), .R(rst_n_bF_buf78), .S(1'b1) );
  DFFSR DFFSR_619 ( .CLK(clk_bF_buf0), .D(AES_CORE_DATAPATH__0iv_1__31_0__22_), .Q(AES_CORE_DATAPATH_iv_1__22_), .R(rst_n_bF_buf77), .S(1'b1) );
  DFFSR DFFSR_62 ( .CLK(clk_bF_buf92), .D(AES_CORE_DATAPATH__0key_0__31_0__9_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__9_), .R(rst_n_bF_buf25), .S(1'b1) );
  DFFSR DFFSR_620 ( .CLK(clk_bF_buf92), .D(AES_CORE_DATAPATH__0iv_1__31_0__23_), .Q(AES_CORE_DATAPATH_iv_1__23_), .R(rst_n_bF_buf76), .S(1'b1) );
  DFFSR DFFSR_621 ( .CLK(clk_bF_buf91), .D(AES_CORE_DATAPATH__0iv_1__31_0__24_), .Q(AES_CORE_DATAPATH_iv_1__24_), .R(rst_n_bF_buf75), .S(1'b1) );
  DFFSR DFFSR_622 ( .CLK(clk_bF_buf90), .D(AES_CORE_DATAPATH__0iv_1__31_0__25_), .Q(AES_CORE_DATAPATH_iv_1__25_), .R(rst_n_bF_buf74), .S(1'b1) );
  DFFSR DFFSR_623 ( .CLK(clk_bF_buf89), .D(AES_CORE_DATAPATH__0iv_1__31_0__26_), .Q(AES_CORE_DATAPATH_iv_1__26_), .R(rst_n_bF_buf73), .S(1'b1) );
  DFFSR DFFSR_624 ( .CLK(clk_bF_buf88), .D(AES_CORE_DATAPATH__0iv_1__31_0__27_), .Q(AES_CORE_DATAPATH_iv_1__27_), .R(rst_n_bF_buf72), .S(1'b1) );
  DFFSR DFFSR_625 ( .CLK(clk_bF_buf87), .D(AES_CORE_DATAPATH__0iv_1__31_0__28_), .Q(AES_CORE_DATAPATH_iv_1__28_), .R(rst_n_bF_buf71), .S(1'b1) );
  DFFSR DFFSR_626 ( .CLK(clk_bF_buf86), .D(AES_CORE_DATAPATH__0iv_1__31_0__29_), .Q(AES_CORE_DATAPATH_iv_1__29_), .R(rst_n_bF_buf70), .S(1'b1) );
  DFFSR DFFSR_627 ( .CLK(clk_bF_buf85), .D(AES_CORE_DATAPATH__0iv_1__31_0__30_), .Q(AES_CORE_DATAPATH_iv_1__30_), .R(rst_n_bF_buf69), .S(1'b1) );
  DFFSR DFFSR_628 ( .CLK(clk_bF_buf84), .D(AES_CORE_DATAPATH__0iv_1__31_0__31_), .Q(AES_CORE_DATAPATH_iv_1__31_), .R(rst_n_bF_buf68), .S(1'b1) );
  DFFSR DFFSR_629 ( .CLK(clk_bF_buf83), .D(AES_CORE_DATAPATH__0bkp_1__31_0__0_), .Q(AES_CORE_DATAPATH_bkp_1__0_), .R(rst_n_bF_buf67), .S(1'b1) );
  DFFSR DFFSR_63 ( .CLK(clk_bF_buf91), .D(AES_CORE_DATAPATH__0key_0__31_0__10_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__10_), .R(rst_n_bF_buf24), .S(1'b1) );
  DFFSR DFFSR_630 ( .CLK(clk_bF_buf82), .D(AES_CORE_DATAPATH__0bkp_1__31_0__1_), .Q(AES_CORE_DATAPATH_bkp_1__1_), .R(rst_n_bF_buf66), .S(1'b1) );
  DFFSR DFFSR_631 ( .CLK(clk_bF_buf81), .D(AES_CORE_DATAPATH__0bkp_1__31_0__2_), .Q(AES_CORE_DATAPATH_bkp_1__2_), .R(rst_n_bF_buf65), .S(1'b1) );
  DFFSR DFFSR_632 ( .CLK(clk_bF_buf80), .D(AES_CORE_DATAPATH__0bkp_1__31_0__3_), .Q(AES_CORE_DATAPATH_bkp_1__3_), .R(rst_n_bF_buf64), .S(1'b1) );
  DFFSR DFFSR_633 ( .CLK(clk_bF_buf79), .D(AES_CORE_DATAPATH__0bkp_1__31_0__4_), .Q(AES_CORE_DATAPATH_bkp_1__4_), .R(rst_n_bF_buf63), .S(1'b1) );
  DFFSR DFFSR_634 ( .CLK(clk_bF_buf78), .D(AES_CORE_DATAPATH__0bkp_1__31_0__5_), .Q(AES_CORE_DATAPATH_bkp_1__5_), .R(rst_n_bF_buf62), .S(1'b1) );
  DFFSR DFFSR_635 ( .CLK(clk_bF_buf77), .D(AES_CORE_DATAPATH__0bkp_1__31_0__6_), .Q(AES_CORE_DATAPATH_bkp_1__6_), .R(rst_n_bF_buf61), .S(1'b1) );
  DFFSR DFFSR_636 ( .CLK(clk_bF_buf76), .D(AES_CORE_DATAPATH__0bkp_1__31_0__7_), .Q(AES_CORE_DATAPATH_bkp_1__7_), .R(rst_n_bF_buf60), .S(1'b1) );
  DFFSR DFFSR_637 ( .CLK(clk_bF_buf75), .D(AES_CORE_DATAPATH__0bkp_1__31_0__8_), .Q(AES_CORE_DATAPATH_bkp_1__8_), .R(rst_n_bF_buf59), .S(1'b1) );
  DFFSR DFFSR_638 ( .CLK(clk_bF_buf74), .D(AES_CORE_DATAPATH__0bkp_1__31_0__9_), .Q(AES_CORE_DATAPATH_bkp_1__9_), .R(rst_n_bF_buf58), .S(1'b1) );
  DFFSR DFFSR_639 ( .CLK(clk_bF_buf73), .D(AES_CORE_DATAPATH__0bkp_1__31_0__10_), .Q(AES_CORE_DATAPATH_bkp_1__10_), .R(rst_n_bF_buf57), .S(1'b1) );
  DFFSR DFFSR_64 ( .CLK(clk_bF_buf90), .D(AES_CORE_DATAPATH__0key_0__31_0__11_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__11_), .R(rst_n_bF_buf23), .S(1'b1) );
  DFFSR DFFSR_640 ( .CLK(clk_bF_buf72), .D(AES_CORE_DATAPATH__0bkp_1__31_0__11_), .Q(AES_CORE_DATAPATH_bkp_1__11_), .R(rst_n_bF_buf56), .S(1'b1) );
  DFFSR DFFSR_641 ( .CLK(clk_bF_buf71), .D(AES_CORE_DATAPATH__0bkp_1__31_0__12_), .Q(AES_CORE_DATAPATH_bkp_1__12_), .R(rst_n_bF_buf55), .S(1'b1) );
  DFFSR DFFSR_642 ( .CLK(clk_bF_buf70), .D(AES_CORE_DATAPATH__0bkp_1__31_0__13_), .Q(AES_CORE_DATAPATH_bkp_1__13_), .R(rst_n_bF_buf54), .S(1'b1) );
  DFFSR DFFSR_643 ( .CLK(clk_bF_buf69), .D(AES_CORE_DATAPATH__0bkp_1__31_0__14_), .Q(AES_CORE_DATAPATH_bkp_1__14_), .R(rst_n_bF_buf53), .S(1'b1) );
  DFFSR DFFSR_644 ( .CLK(clk_bF_buf68), .D(AES_CORE_DATAPATH__0bkp_1__31_0__15_), .Q(AES_CORE_DATAPATH_bkp_1__15_), .R(rst_n_bF_buf52), .S(1'b1) );
  DFFSR DFFSR_645 ( .CLK(clk_bF_buf67), .D(AES_CORE_DATAPATH__0bkp_1__31_0__16_), .Q(AES_CORE_DATAPATH_bkp_1__16_), .R(rst_n_bF_buf51), .S(1'b1) );
  DFFSR DFFSR_646 ( .CLK(clk_bF_buf66), .D(AES_CORE_DATAPATH__0bkp_1__31_0__17_), .Q(AES_CORE_DATAPATH_bkp_1__17_), .R(rst_n_bF_buf50), .S(1'b1) );
  DFFSR DFFSR_647 ( .CLK(clk_bF_buf65), .D(AES_CORE_DATAPATH__0bkp_1__31_0__18_), .Q(AES_CORE_DATAPATH_bkp_1__18_), .R(rst_n_bF_buf49), .S(1'b1) );
  DFFSR DFFSR_648 ( .CLK(clk_bF_buf64), .D(AES_CORE_DATAPATH__0bkp_1__31_0__19_), .Q(AES_CORE_DATAPATH_bkp_1__19_), .R(rst_n_bF_buf48), .S(1'b1) );
  DFFSR DFFSR_649 ( .CLK(clk_bF_buf63), .D(AES_CORE_DATAPATH__0bkp_1__31_0__20_), .Q(AES_CORE_DATAPATH_bkp_1__20_), .R(rst_n_bF_buf47), .S(1'b1) );
  DFFSR DFFSR_65 ( .CLK(clk_bF_buf89), .D(AES_CORE_DATAPATH__0key_0__31_0__12_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__12_), .R(rst_n_bF_buf22), .S(1'b1) );
  DFFSR DFFSR_650 ( .CLK(clk_bF_buf62), .D(AES_CORE_DATAPATH__0bkp_1__31_0__21_), .Q(AES_CORE_DATAPATH_bkp_1__21_), .R(rst_n_bF_buf46), .S(1'b1) );
  DFFSR DFFSR_651 ( .CLK(clk_bF_buf61), .D(AES_CORE_DATAPATH__0bkp_1__31_0__22_), .Q(AES_CORE_DATAPATH_bkp_1__22_), .R(rst_n_bF_buf45), .S(1'b1) );
  DFFSR DFFSR_652 ( .CLK(clk_bF_buf60), .D(AES_CORE_DATAPATH__0bkp_1__31_0__23_), .Q(AES_CORE_DATAPATH_bkp_1__23_), .R(rst_n_bF_buf44), .S(1'b1) );
  DFFSR DFFSR_653 ( .CLK(clk_bF_buf59), .D(AES_CORE_DATAPATH__0bkp_1__31_0__24_), .Q(AES_CORE_DATAPATH_bkp_1__24_), .R(rst_n_bF_buf43), .S(1'b1) );
  DFFSR DFFSR_654 ( .CLK(clk_bF_buf58), .D(AES_CORE_DATAPATH__0bkp_1__31_0__25_), .Q(AES_CORE_DATAPATH_bkp_1__25_), .R(rst_n_bF_buf42), .S(1'b1) );
  DFFSR DFFSR_655 ( .CLK(clk_bF_buf57), .D(AES_CORE_DATAPATH__0bkp_1__31_0__26_), .Q(AES_CORE_DATAPATH_bkp_1__26_), .R(rst_n_bF_buf41), .S(1'b1) );
  DFFSR DFFSR_656 ( .CLK(clk_bF_buf56), .D(AES_CORE_DATAPATH__0bkp_1__31_0__27_), .Q(AES_CORE_DATAPATH_bkp_1__27_), .R(rst_n_bF_buf40), .S(1'b1) );
  DFFSR DFFSR_657 ( .CLK(clk_bF_buf55), .D(AES_CORE_DATAPATH__0bkp_1__31_0__28_), .Q(AES_CORE_DATAPATH_bkp_1__28_), .R(rst_n_bF_buf39), .S(1'b1) );
  DFFSR DFFSR_658 ( .CLK(clk_bF_buf54), .D(AES_CORE_DATAPATH__0bkp_1__31_0__29_), .Q(AES_CORE_DATAPATH_bkp_1__29_), .R(rst_n_bF_buf38), .S(1'b1) );
  DFFSR DFFSR_659 ( .CLK(clk_bF_buf53), .D(AES_CORE_DATAPATH__0bkp_1__31_0__30_), .Q(AES_CORE_DATAPATH_bkp_1__30_), .R(rst_n_bF_buf37), .S(1'b1) );
  DFFSR DFFSR_66 ( .CLK(clk_bF_buf88), .D(AES_CORE_DATAPATH__0key_0__31_0__13_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__13_), .R(rst_n_bF_buf21), .S(1'b1) );
  DFFSR DFFSR_660 ( .CLK(clk_bF_buf52), .D(AES_CORE_DATAPATH__0bkp_1__31_0__31_), .Q(AES_CORE_DATAPATH_bkp_1__31_), .R(rst_n_bF_buf36), .S(1'b1) );
  DFFSR DFFSR_661 ( .CLK(clk_bF_buf51), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__0_), .Q(AES_CORE_DATAPATH_bkp_1_1__0_), .R(rst_n_bF_buf35), .S(1'b1) );
  DFFSR DFFSR_662 ( .CLK(clk_bF_buf50), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__1_), .Q(AES_CORE_DATAPATH_bkp_1_1__1_), .R(rst_n_bF_buf34), .S(1'b1) );
  DFFSR DFFSR_663 ( .CLK(clk_bF_buf49), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__2_), .Q(AES_CORE_DATAPATH_bkp_1_1__2_), .R(rst_n_bF_buf33), .S(1'b1) );
  DFFSR DFFSR_664 ( .CLK(clk_bF_buf48), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__3_), .Q(AES_CORE_DATAPATH_bkp_1_1__3_), .R(rst_n_bF_buf32), .S(1'b1) );
  DFFSR DFFSR_665 ( .CLK(clk_bF_buf47), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__4_), .Q(AES_CORE_DATAPATH_bkp_1_1__4_), .R(rst_n_bF_buf31), .S(1'b1) );
  DFFSR DFFSR_666 ( .CLK(clk_bF_buf46), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__5_), .Q(AES_CORE_DATAPATH_bkp_1_1__5_), .R(rst_n_bF_buf30), .S(1'b1) );
  DFFSR DFFSR_667 ( .CLK(clk_bF_buf45), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__6_), .Q(AES_CORE_DATAPATH_bkp_1_1__6_), .R(rst_n_bF_buf29), .S(1'b1) );
  DFFSR DFFSR_668 ( .CLK(clk_bF_buf44), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__7_), .Q(AES_CORE_DATAPATH_bkp_1_1__7_), .R(rst_n_bF_buf28), .S(1'b1) );
  DFFSR DFFSR_669 ( .CLK(clk_bF_buf43), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__8_), .Q(AES_CORE_DATAPATH_bkp_1_1__8_), .R(rst_n_bF_buf27), .S(1'b1) );
  DFFSR DFFSR_67 ( .CLK(clk_bF_buf87), .D(AES_CORE_DATAPATH__0key_0__31_0__14_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__14_), .R(rst_n_bF_buf20), .S(1'b1) );
  DFFSR DFFSR_670 ( .CLK(clk_bF_buf42), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__9_), .Q(AES_CORE_DATAPATH_bkp_1_1__9_), .R(rst_n_bF_buf26), .S(1'b1) );
  DFFSR DFFSR_671 ( .CLK(clk_bF_buf41), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__10_), .Q(AES_CORE_DATAPATH_bkp_1_1__10_), .R(rst_n_bF_buf25), .S(1'b1) );
  DFFSR DFFSR_672 ( .CLK(clk_bF_buf40), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__11_), .Q(AES_CORE_DATAPATH_bkp_1_1__11_), .R(rst_n_bF_buf24), .S(1'b1) );
  DFFSR DFFSR_673 ( .CLK(clk_bF_buf39), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__12_), .Q(AES_CORE_DATAPATH_bkp_1_1__12_), .R(rst_n_bF_buf23), .S(1'b1) );
  DFFSR DFFSR_674 ( .CLK(clk_bF_buf38), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__13_), .Q(AES_CORE_DATAPATH_bkp_1_1__13_), .R(rst_n_bF_buf22), .S(1'b1) );
  DFFSR DFFSR_675 ( .CLK(clk_bF_buf37), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__14_), .Q(AES_CORE_DATAPATH_bkp_1_1__14_), .R(rst_n_bF_buf21), .S(1'b1) );
  DFFSR DFFSR_676 ( .CLK(clk_bF_buf36), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__15_), .Q(AES_CORE_DATAPATH_bkp_1_1__15_), .R(rst_n_bF_buf20), .S(1'b1) );
  DFFSR DFFSR_677 ( .CLK(clk_bF_buf35), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__16_), .Q(AES_CORE_DATAPATH_bkp_1_1__16_), .R(rst_n_bF_buf19), .S(1'b1) );
  DFFSR DFFSR_678 ( .CLK(clk_bF_buf34), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__17_), .Q(AES_CORE_DATAPATH_bkp_1_1__17_), .R(rst_n_bF_buf18), .S(1'b1) );
  DFFSR DFFSR_679 ( .CLK(clk_bF_buf33), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__18_), .Q(AES_CORE_DATAPATH_bkp_1_1__18_), .R(rst_n_bF_buf17), .S(1'b1) );
  DFFSR DFFSR_68 ( .CLK(clk_bF_buf86), .D(AES_CORE_DATAPATH__0key_0__31_0__15_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__15_), .R(rst_n_bF_buf19), .S(1'b1) );
  DFFSR DFFSR_680 ( .CLK(clk_bF_buf32), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__19_), .Q(AES_CORE_DATAPATH_bkp_1_1__19_), .R(rst_n_bF_buf16), .S(1'b1) );
  DFFSR DFFSR_681 ( .CLK(clk_bF_buf31), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__20_), .Q(AES_CORE_DATAPATH_bkp_1_1__20_), .R(rst_n_bF_buf15), .S(1'b1) );
  DFFSR DFFSR_682 ( .CLK(clk_bF_buf30), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__21_), .Q(AES_CORE_DATAPATH_bkp_1_1__21_), .R(rst_n_bF_buf14), .S(1'b1) );
  DFFSR DFFSR_683 ( .CLK(clk_bF_buf29), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__22_), .Q(AES_CORE_DATAPATH_bkp_1_1__22_), .R(rst_n_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_684 ( .CLK(clk_bF_buf28), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__23_), .Q(AES_CORE_DATAPATH_bkp_1_1__23_), .R(rst_n_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_685 ( .CLK(clk_bF_buf27), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__24_), .Q(AES_CORE_DATAPATH_bkp_1_1__24_), .R(rst_n_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_686 ( .CLK(clk_bF_buf26), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__25_), .Q(AES_CORE_DATAPATH_bkp_1_1__25_), .R(rst_n_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_687 ( .CLK(clk_bF_buf25), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__26_), .Q(AES_CORE_DATAPATH_bkp_1_1__26_), .R(rst_n_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_688 ( .CLK(clk_bF_buf24), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__27_), .Q(AES_CORE_DATAPATH_bkp_1_1__27_), .R(rst_n_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_689 ( .CLK(clk_bF_buf23), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__28_), .Q(AES_CORE_DATAPATH_bkp_1_1__28_), .R(rst_n_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_69 ( .CLK(clk_bF_buf85), .D(AES_CORE_DATAPATH__0key_0__31_0__16_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__16_), .R(rst_n_bF_buf18), .S(1'b1) );
  DFFSR DFFSR_690 ( .CLK(clk_bF_buf22), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__29_), .Q(AES_CORE_DATAPATH_bkp_1_1__29_), .R(rst_n_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_691 ( .CLK(clk_bF_buf21), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__30_), .Q(AES_CORE_DATAPATH_bkp_1_1__30_), .R(rst_n_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_692 ( .CLK(clk_bF_buf20), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__31_), .Q(AES_CORE_DATAPATH_bkp_1_1__31_), .R(rst_n_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_693 ( .CLK(clk_bF_buf19), .D(AES_CORE_DATAPATH__0iv_0__31_0__0_), .Q(AES_CORE_DATAPATH_iv_0__0_), .R(rst_n_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_694 ( .CLK(clk_bF_buf18), .D(AES_CORE_DATAPATH__0iv_0__31_0__1_), .Q(AES_CORE_DATAPATH_iv_0__1_), .R(rst_n_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_695 ( .CLK(clk_bF_buf17), .D(AES_CORE_DATAPATH__0iv_0__31_0__2_), .Q(AES_CORE_DATAPATH_iv_0__2_), .R(rst_n_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_696 ( .CLK(clk_bF_buf16), .D(AES_CORE_DATAPATH__0iv_0__31_0__3_), .Q(AES_CORE_DATAPATH_iv_0__3_), .R(rst_n_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_697 ( .CLK(clk_bF_buf15), .D(AES_CORE_DATAPATH__0iv_0__31_0__4_), .Q(AES_CORE_DATAPATH_iv_0__4_), .R(rst_n_bF_buf86), .S(1'b1) );
  DFFSR DFFSR_698 ( .CLK(clk_bF_buf14), .D(AES_CORE_DATAPATH__0iv_0__31_0__5_), .Q(AES_CORE_DATAPATH_iv_0__5_), .R(rst_n_bF_buf85), .S(1'b1) );
  DFFSR DFFSR_699 ( .CLK(clk_bF_buf13), .D(AES_CORE_DATAPATH__0iv_0__31_0__6_), .Q(AES_CORE_DATAPATH_iv_0__6_), .R(rst_n_bF_buf84), .S(1'b1) );
  DFFSR DFFSR_7 ( .CLK(clk_bF_buf86), .D(AES_CORE_CONTROL_UNIT__abc_10818_n4), .Q(AES_CORE_CONTROL_UNIT_state_2_), .R(rst_n_bF_buf80), .S(1'b1) );
  DFFSR DFFSR_70 ( .CLK(clk_bF_buf84), .D(AES_CORE_DATAPATH__0key_0__31_0__17_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__17_), .R(rst_n_bF_buf17), .S(1'b1) );
  DFFSR DFFSR_700 ( .CLK(clk_bF_buf12), .D(AES_CORE_DATAPATH__0iv_0__31_0__7_), .Q(AES_CORE_DATAPATH_iv_0__7_), .R(rst_n_bF_buf83), .S(1'b1) );
  DFFSR DFFSR_701 ( .CLK(clk_bF_buf11), .D(AES_CORE_DATAPATH__0iv_0__31_0__8_), .Q(AES_CORE_DATAPATH_iv_0__8_), .R(rst_n_bF_buf82), .S(1'b1) );
  DFFSR DFFSR_702 ( .CLK(clk_bF_buf10), .D(AES_CORE_DATAPATH__0iv_0__31_0__9_), .Q(AES_CORE_DATAPATH_iv_0__9_), .R(rst_n_bF_buf81), .S(1'b1) );
  DFFSR DFFSR_703 ( .CLK(clk_bF_buf9), .D(AES_CORE_DATAPATH__0iv_0__31_0__10_), .Q(AES_CORE_DATAPATH_iv_0__10_), .R(rst_n_bF_buf80), .S(1'b1) );
  DFFSR DFFSR_704 ( .CLK(clk_bF_buf8), .D(AES_CORE_DATAPATH__0iv_0__31_0__11_), .Q(AES_CORE_DATAPATH_iv_0__11_), .R(rst_n_bF_buf79), .S(1'b1) );
  DFFSR DFFSR_705 ( .CLK(clk_bF_buf7), .D(AES_CORE_DATAPATH__0iv_0__31_0__12_), .Q(AES_CORE_DATAPATH_iv_0__12_), .R(rst_n_bF_buf78), .S(1'b1) );
  DFFSR DFFSR_706 ( .CLK(clk_bF_buf6), .D(AES_CORE_DATAPATH__0iv_0__31_0__13_), .Q(AES_CORE_DATAPATH_iv_0__13_), .R(rst_n_bF_buf77), .S(1'b1) );
  DFFSR DFFSR_707 ( .CLK(clk_bF_buf5), .D(AES_CORE_DATAPATH__0iv_0__31_0__14_), .Q(AES_CORE_DATAPATH_iv_0__14_), .R(rst_n_bF_buf76), .S(1'b1) );
  DFFSR DFFSR_708 ( .CLK(clk_bF_buf4), .D(AES_CORE_DATAPATH__0iv_0__31_0__15_), .Q(AES_CORE_DATAPATH_iv_0__15_), .R(rst_n_bF_buf75), .S(1'b1) );
  DFFSR DFFSR_709 ( .CLK(clk_bF_buf3), .D(AES_CORE_DATAPATH__0iv_0__31_0__16_), .Q(AES_CORE_DATAPATH_iv_0__16_), .R(rst_n_bF_buf74), .S(1'b1) );
  DFFSR DFFSR_71 ( .CLK(clk_bF_buf83), .D(AES_CORE_DATAPATH__0key_0__31_0__18_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__18_), .R(rst_n_bF_buf16), .S(1'b1) );
  DFFSR DFFSR_710 ( .CLK(clk_bF_buf2), .D(AES_CORE_DATAPATH__0iv_0__31_0__17_), .Q(AES_CORE_DATAPATH_iv_0__17_), .R(rst_n_bF_buf73), .S(1'b1) );
  DFFSR DFFSR_711 ( .CLK(clk_bF_buf1), .D(AES_CORE_DATAPATH__0iv_0__31_0__18_), .Q(AES_CORE_DATAPATH_iv_0__18_), .R(rst_n_bF_buf72), .S(1'b1) );
  DFFSR DFFSR_712 ( .CLK(clk_bF_buf0), .D(AES_CORE_DATAPATH__0iv_0__31_0__19_), .Q(AES_CORE_DATAPATH_iv_0__19_), .R(rst_n_bF_buf71), .S(1'b1) );
  DFFSR DFFSR_713 ( .CLK(clk_bF_buf92), .D(AES_CORE_DATAPATH__0iv_0__31_0__20_), .Q(AES_CORE_DATAPATH_iv_0__20_), .R(rst_n_bF_buf70), .S(1'b1) );
  DFFSR DFFSR_714 ( .CLK(clk_bF_buf91), .D(AES_CORE_DATAPATH__0iv_0__31_0__21_), .Q(AES_CORE_DATAPATH_iv_0__21_), .R(rst_n_bF_buf69), .S(1'b1) );
  DFFSR DFFSR_715 ( .CLK(clk_bF_buf90), .D(AES_CORE_DATAPATH__0iv_0__31_0__22_), .Q(AES_CORE_DATAPATH_iv_0__22_), .R(rst_n_bF_buf68), .S(1'b1) );
  DFFSR DFFSR_716 ( .CLK(clk_bF_buf89), .D(AES_CORE_DATAPATH__0iv_0__31_0__23_), .Q(AES_CORE_DATAPATH_iv_0__23_), .R(rst_n_bF_buf67), .S(1'b1) );
  DFFSR DFFSR_717 ( .CLK(clk_bF_buf88), .D(AES_CORE_DATAPATH__0iv_0__31_0__24_), .Q(AES_CORE_DATAPATH_iv_0__24_), .R(rst_n_bF_buf66), .S(1'b1) );
  DFFSR DFFSR_718 ( .CLK(clk_bF_buf87), .D(AES_CORE_DATAPATH__0iv_0__31_0__25_), .Q(AES_CORE_DATAPATH_iv_0__25_), .R(rst_n_bF_buf65), .S(1'b1) );
  DFFSR DFFSR_719 ( .CLK(clk_bF_buf86), .D(AES_CORE_DATAPATH__0iv_0__31_0__26_), .Q(AES_CORE_DATAPATH_iv_0__26_), .R(rst_n_bF_buf64), .S(1'b1) );
  DFFSR DFFSR_72 ( .CLK(clk_bF_buf82), .D(AES_CORE_DATAPATH__0key_0__31_0__19_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__19_), .R(rst_n_bF_buf15), .S(1'b1) );
  DFFSR DFFSR_720 ( .CLK(clk_bF_buf85), .D(AES_CORE_DATAPATH__0iv_0__31_0__27_), .Q(AES_CORE_DATAPATH_iv_0__27_), .R(rst_n_bF_buf63), .S(1'b1) );
  DFFSR DFFSR_721 ( .CLK(clk_bF_buf84), .D(AES_CORE_DATAPATH__0iv_0__31_0__28_), .Q(AES_CORE_DATAPATH_iv_0__28_), .R(rst_n_bF_buf62), .S(1'b1) );
  DFFSR DFFSR_722 ( .CLK(clk_bF_buf83), .D(AES_CORE_DATAPATH__0iv_0__31_0__29_), .Q(AES_CORE_DATAPATH_iv_0__29_), .R(rst_n_bF_buf61), .S(1'b1) );
  DFFSR DFFSR_723 ( .CLK(clk_bF_buf82), .D(AES_CORE_DATAPATH__0iv_0__31_0__30_), .Q(AES_CORE_DATAPATH_iv_0__30_), .R(rst_n_bF_buf60), .S(1'b1) );
  DFFSR DFFSR_724 ( .CLK(clk_bF_buf81), .D(AES_CORE_DATAPATH__0iv_0__31_0__31_), .Q(AES_CORE_DATAPATH_iv_0__31_), .R(rst_n_bF_buf59), .S(1'b1) );
  DFFSR DFFSR_725 ( .CLK(clk_bF_buf80), .D(AES_CORE_DATAPATH__0bkp_0__31_0__0_), .Q(AES_CORE_DATAPATH_bkp_0__0_), .R(rst_n_bF_buf58), .S(1'b1) );
  DFFSR DFFSR_726 ( .CLK(clk_bF_buf79), .D(AES_CORE_DATAPATH__0bkp_0__31_0__1_), .Q(AES_CORE_DATAPATH_bkp_0__1_), .R(rst_n_bF_buf57), .S(1'b1) );
  DFFSR DFFSR_727 ( .CLK(clk_bF_buf78), .D(AES_CORE_DATAPATH__0bkp_0__31_0__2_), .Q(AES_CORE_DATAPATH_bkp_0__2_), .R(rst_n_bF_buf56), .S(1'b1) );
  DFFSR DFFSR_728 ( .CLK(clk_bF_buf77), .D(AES_CORE_DATAPATH__0bkp_0__31_0__3_), .Q(AES_CORE_DATAPATH_bkp_0__3_), .R(rst_n_bF_buf55), .S(1'b1) );
  DFFSR DFFSR_729 ( .CLK(clk_bF_buf76), .D(AES_CORE_DATAPATH__0bkp_0__31_0__4_), .Q(AES_CORE_DATAPATH_bkp_0__4_), .R(rst_n_bF_buf54), .S(1'b1) );
  DFFSR DFFSR_73 ( .CLK(clk_bF_buf81), .D(AES_CORE_DATAPATH__0key_0__31_0__20_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__20_), .R(rst_n_bF_buf14), .S(1'b1) );
  DFFSR DFFSR_730 ( .CLK(clk_bF_buf75), .D(AES_CORE_DATAPATH__0bkp_0__31_0__5_), .Q(AES_CORE_DATAPATH_bkp_0__5_), .R(rst_n_bF_buf53), .S(1'b1) );
  DFFSR DFFSR_731 ( .CLK(clk_bF_buf74), .D(AES_CORE_DATAPATH__0bkp_0__31_0__6_), .Q(AES_CORE_DATAPATH_bkp_0__6_), .R(rst_n_bF_buf52), .S(1'b1) );
  DFFSR DFFSR_732 ( .CLK(clk_bF_buf73), .D(AES_CORE_DATAPATH__0bkp_0__31_0__7_), .Q(AES_CORE_DATAPATH_bkp_0__7_), .R(rst_n_bF_buf51), .S(1'b1) );
  DFFSR DFFSR_733 ( .CLK(clk_bF_buf72), .D(AES_CORE_DATAPATH__0bkp_0__31_0__8_), .Q(AES_CORE_DATAPATH_bkp_0__8_), .R(rst_n_bF_buf50), .S(1'b1) );
  DFFSR DFFSR_734 ( .CLK(clk_bF_buf71), .D(AES_CORE_DATAPATH__0bkp_0__31_0__9_), .Q(AES_CORE_DATAPATH_bkp_0__9_), .R(rst_n_bF_buf49), .S(1'b1) );
  DFFSR DFFSR_735 ( .CLK(clk_bF_buf70), .D(AES_CORE_DATAPATH__0bkp_0__31_0__10_), .Q(AES_CORE_DATAPATH_bkp_0__10_), .R(rst_n_bF_buf48), .S(1'b1) );
  DFFSR DFFSR_736 ( .CLK(clk_bF_buf69), .D(AES_CORE_DATAPATH__0bkp_0__31_0__11_), .Q(AES_CORE_DATAPATH_bkp_0__11_), .R(rst_n_bF_buf47), .S(1'b1) );
  DFFSR DFFSR_737 ( .CLK(clk_bF_buf68), .D(AES_CORE_DATAPATH__0bkp_0__31_0__12_), .Q(AES_CORE_DATAPATH_bkp_0__12_), .R(rst_n_bF_buf46), .S(1'b1) );
  DFFSR DFFSR_738 ( .CLK(clk_bF_buf67), .D(AES_CORE_DATAPATH__0bkp_0__31_0__13_), .Q(AES_CORE_DATAPATH_bkp_0__13_), .R(rst_n_bF_buf45), .S(1'b1) );
  DFFSR DFFSR_739 ( .CLK(clk_bF_buf66), .D(AES_CORE_DATAPATH__0bkp_0__31_0__14_), .Q(AES_CORE_DATAPATH_bkp_0__14_), .R(rst_n_bF_buf44), .S(1'b1) );
  DFFSR DFFSR_74 ( .CLK(clk_bF_buf80), .D(AES_CORE_DATAPATH__0key_0__31_0__21_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__21_), .R(rst_n_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_740 ( .CLK(clk_bF_buf65), .D(AES_CORE_DATAPATH__0bkp_0__31_0__15_), .Q(AES_CORE_DATAPATH_bkp_0__15_), .R(rst_n_bF_buf43), .S(1'b1) );
  DFFSR DFFSR_741 ( .CLK(clk_bF_buf64), .D(AES_CORE_DATAPATH__0bkp_0__31_0__16_), .Q(AES_CORE_DATAPATH_bkp_0__16_), .R(rst_n_bF_buf42), .S(1'b1) );
  DFFSR DFFSR_742 ( .CLK(clk_bF_buf63), .D(AES_CORE_DATAPATH__0bkp_0__31_0__17_), .Q(AES_CORE_DATAPATH_bkp_0__17_), .R(rst_n_bF_buf41), .S(1'b1) );
  DFFSR DFFSR_743 ( .CLK(clk_bF_buf62), .D(AES_CORE_DATAPATH__0bkp_0__31_0__18_), .Q(AES_CORE_DATAPATH_bkp_0__18_), .R(rst_n_bF_buf40), .S(1'b1) );
  DFFSR DFFSR_744 ( .CLK(clk_bF_buf61), .D(AES_CORE_DATAPATH__0bkp_0__31_0__19_), .Q(AES_CORE_DATAPATH_bkp_0__19_), .R(rst_n_bF_buf39), .S(1'b1) );
  DFFSR DFFSR_745 ( .CLK(clk_bF_buf60), .D(AES_CORE_DATAPATH__0bkp_0__31_0__20_), .Q(AES_CORE_DATAPATH_bkp_0__20_), .R(rst_n_bF_buf38), .S(1'b1) );
  DFFSR DFFSR_746 ( .CLK(clk_bF_buf59), .D(AES_CORE_DATAPATH__0bkp_0__31_0__21_), .Q(AES_CORE_DATAPATH_bkp_0__21_), .R(rst_n_bF_buf37), .S(1'b1) );
  DFFSR DFFSR_747 ( .CLK(clk_bF_buf58), .D(AES_CORE_DATAPATH__0bkp_0__31_0__22_), .Q(AES_CORE_DATAPATH_bkp_0__22_), .R(rst_n_bF_buf36), .S(1'b1) );
  DFFSR DFFSR_748 ( .CLK(clk_bF_buf57), .D(AES_CORE_DATAPATH__0bkp_0__31_0__23_), .Q(AES_CORE_DATAPATH_bkp_0__23_), .R(rst_n_bF_buf35), .S(1'b1) );
  DFFSR DFFSR_749 ( .CLK(clk_bF_buf56), .D(AES_CORE_DATAPATH__0bkp_0__31_0__24_), .Q(AES_CORE_DATAPATH_bkp_0__24_), .R(rst_n_bF_buf34), .S(1'b1) );
  DFFSR DFFSR_75 ( .CLK(clk_bF_buf79), .D(AES_CORE_DATAPATH__0key_0__31_0__22_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__22_), .R(rst_n_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_750 ( .CLK(clk_bF_buf55), .D(AES_CORE_DATAPATH__0bkp_0__31_0__25_), .Q(AES_CORE_DATAPATH_bkp_0__25_), .R(rst_n_bF_buf33), .S(1'b1) );
  DFFSR DFFSR_751 ( .CLK(clk_bF_buf54), .D(AES_CORE_DATAPATH__0bkp_0__31_0__26_), .Q(AES_CORE_DATAPATH_bkp_0__26_), .R(rst_n_bF_buf32), .S(1'b1) );
  DFFSR DFFSR_752 ( .CLK(clk_bF_buf53), .D(AES_CORE_DATAPATH__0bkp_0__31_0__27_), .Q(AES_CORE_DATAPATH_bkp_0__27_), .R(rst_n_bF_buf31), .S(1'b1) );
  DFFSR DFFSR_753 ( .CLK(clk_bF_buf52), .D(AES_CORE_DATAPATH__0bkp_0__31_0__28_), .Q(AES_CORE_DATAPATH_bkp_0__28_), .R(rst_n_bF_buf30), .S(1'b1) );
  DFFSR DFFSR_754 ( .CLK(clk_bF_buf51), .D(AES_CORE_DATAPATH__0bkp_0__31_0__29_), .Q(AES_CORE_DATAPATH_bkp_0__29_), .R(rst_n_bF_buf29), .S(1'b1) );
  DFFSR DFFSR_755 ( .CLK(clk_bF_buf50), .D(AES_CORE_DATAPATH__0bkp_0__31_0__30_), .Q(AES_CORE_DATAPATH_bkp_0__30_), .R(rst_n_bF_buf28), .S(1'b1) );
  DFFSR DFFSR_756 ( .CLK(clk_bF_buf49), .D(AES_CORE_DATAPATH__0bkp_0__31_0__31_), .Q(AES_CORE_DATAPATH_bkp_0__31_), .R(rst_n_bF_buf27), .S(1'b1) );
  DFFSR DFFSR_757 ( .CLK(clk_bF_buf48), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__0_), .Q(AES_CORE_DATAPATH_bkp_1_0__0_), .R(rst_n_bF_buf26), .S(1'b1) );
  DFFSR DFFSR_758 ( .CLK(clk_bF_buf47), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__1_), .Q(AES_CORE_DATAPATH_bkp_1_0__1_), .R(rst_n_bF_buf25), .S(1'b1) );
  DFFSR DFFSR_759 ( .CLK(clk_bF_buf46), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__2_), .Q(AES_CORE_DATAPATH_bkp_1_0__2_), .R(rst_n_bF_buf24), .S(1'b1) );
  DFFSR DFFSR_76 ( .CLK(clk_bF_buf78), .D(AES_CORE_DATAPATH__0key_0__31_0__23_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__23_), .R(rst_n_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_760 ( .CLK(clk_bF_buf45), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__3_), .Q(AES_CORE_DATAPATH_bkp_1_0__3_), .R(rst_n_bF_buf23), .S(1'b1) );
  DFFSR DFFSR_761 ( .CLK(clk_bF_buf44), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__4_), .Q(AES_CORE_DATAPATH_bkp_1_0__4_), .R(rst_n_bF_buf22), .S(1'b1) );
  DFFSR DFFSR_762 ( .CLK(clk_bF_buf43), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__5_), .Q(AES_CORE_DATAPATH_bkp_1_0__5_), .R(rst_n_bF_buf21), .S(1'b1) );
  DFFSR DFFSR_763 ( .CLK(clk_bF_buf42), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__6_), .Q(AES_CORE_DATAPATH_bkp_1_0__6_), .R(rst_n_bF_buf20), .S(1'b1) );
  DFFSR DFFSR_764 ( .CLK(clk_bF_buf41), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__7_), .Q(AES_CORE_DATAPATH_bkp_1_0__7_), .R(rst_n_bF_buf19), .S(1'b1) );
  DFFSR DFFSR_765 ( .CLK(clk_bF_buf40), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__8_), .Q(AES_CORE_DATAPATH_bkp_1_0__8_), .R(rst_n_bF_buf18), .S(1'b1) );
  DFFSR DFFSR_766 ( .CLK(clk_bF_buf39), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__9_), .Q(AES_CORE_DATAPATH_bkp_1_0__9_), .R(rst_n_bF_buf17), .S(1'b1) );
  DFFSR DFFSR_767 ( .CLK(clk_bF_buf38), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__10_), .Q(AES_CORE_DATAPATH_bkp_1_0__10_), .R(rst_n_bF_buf16), .S(1'b1) );
  DFFSR DFFSR_768 ( .CLK(clk_bF_buf37), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__11_), .Q(AES_CORE_DATAPATH_bkp_1_0__11_), .R(rst_n_bF_buf15), .S(1'b1) );
  DFFSR DFFSR_769 ( .CLK(clk_bF_buf36), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__12_), .Q(AES_CORE_DATAPATH_bkp_1_0__12_), .R(rst_n_bF_buf14), .S(1'b1) );
  DFFSR DFFSR_77 ( .CLK(clk_bF_buf77), .D(AES_CORE_DATAPATH__0key_0__31_0__24_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__24_), .R(rst_n_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_770 ( .CLK(clk_bF_buf35), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__13_), .Q(AES_CORE_DATAPATH_bkp_1_0__13_), .R(rst_n_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_771 ( .CLK(clk_bF_buf34), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__14_), .Q(AES_CORE_DATAPATH_bkp_1_0__14_), .R(rst_n_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_772 ( .CLK(clk_bF_buf33), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__15_), .Q(AES_CORE_DATAPATH_bkp_1_0__15_), .R(rst_n_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_773 ( .CLK(clk_bF_buf32), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__16_), .Q(AES_CORE_DATAPATH_bkp_1_0__16_), .R(rst_n_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_774 ( .CLK(clk_bF_buf31), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__17_), .Q(AES_CORE_DATAPATH_bkp_1_0__17_), .R(rst_n_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_775 ( .CLK(clk_bF_buf30), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__18_), .Q(AES_CORE_DATAPATH_bkp_1_0__18_), .R(rst_n_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_776 ( .CLK(clk_bF_buf29), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__19_), .Q(AES_CORE_DATAPATH_bkp_1_0__19_), .R(rst_n_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_777 ( .CLK(clk_bF_buf28), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__20_), .Q(AES_CORE_DATAPATH_bkp_1_0__20_), .R(rst_n_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_778 ( .CLK(clk_bF_buf27), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__21_), .Q(AES_CORE_DATAPATH_bkp_1_0__21_), .R(rst_n_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_779 ( .CLK(clk_bF_buf26), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__22_), .Q(AES_CORE_DATAPATH_bkp_1_0__22_), .R(rst_n_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_78 ( .CLK(clk_bF_buf76), .D(AES_CORE_DATAPATH__0key_0__31_0__25_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__25_), .R(rst_n_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_780 ( .CLK(clk_bF_buf25), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__23_), .Q(AES_CORE_DATAPATH_bkp_1_0__23_), .R(rst_n_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_781 ( .CLK(clk_bF_buf24), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__24_), .Q(AES_CORE_DATAPATH_bkp_1_0__24_), .R(rst_n_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_782 ( .CLK(clk_bF_buf23), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__25_), .Q(AES_CORE_DATAPATH_bkp_1_0__25_), .R(rst_n_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_783 ( .CLK(clk_bF_buf22), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__26_), .Q(AES_CORE_DATAPATH_bkp_1_0__26_), .R(rst_n_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_784 ( .CLK(clk_bF_buf21), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__27_), .Q(AES_CORE_DATAPATH_bkp_1_0__27_), .R(rst_n_bF_buf86), .S(1'b1) );
  DFFSR DFFSR_785 ( .CLK(clk_bF_buf20), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__28_), .Q(AES_CORE_DATAPATH_bkp_1_0__28_), .R(rst_n_bF_buf85), .S(1'b1) );
  DFFSR DFFSR_786 ( .CLK(clk_bF_buf19), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__29_), .Q(AES_CORE_DATAPATH_bkp_1_0__29_), .R(rst_n_bF_buf84), .S(1'b1) );
  DFFSR DFFSR_787 ( .CLK(clk_bF_buf18), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__30_), .Q(AES_CORE_DATAPATH_bkp_1_0__30_), .R(rst_n_bF_buf83), .S(1'b1) );
  DFFSR DFFSR_788 ( .CLK(clk_bF_buf17), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__31_), .Q(AES_CORE_DATAPATH_bkp_1_0__31_), .R(rst_n_bF_buf82), .S(1'b1) );
  DFFSR DFFSR_789 ( .CLK(clk_bF_buf16), .D(AES_CORE_DATAPATH_col_en_cnt_unit_pp1_0__FF_INPUT), .Q(AES_CORE_DATAPATH_col_en_cnt_unit_pp1_0_), .R(rst_n_bF_buf81), .S(1'b1) );
  DFFSR DFFSR_79 ( .CLK(clk_bF_buf75), .D(AES_CORE_DATAPATH__0key_0__31_0__26_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__26_), .R(rst_n_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_790 ( .CLK(clk_bF_buf15), .D(AES_CORE_DATAPATH_col_en_cnt_unit_pp1_1__FF_INPUT), .Q(AES_CORE_DATAPATH_col_en_cnt_unit_pp1_1_), .R(rst_n_bF_buf80), .S(1'b1) );
  DFFSR DFFSR_791 ( .CLK(clk_bF_buf14), .D(AES_CORE_DATAPATH_col_en_cnt_unit_pp1_2__FF_INPUT), .Q(AES_CORE_DATAPATH_col_en_cnt_unit_pp1_2_), .R(rst_n_bF_buf79), .S(1'b1) );
  DFFSR DFFSR_792 ( .CLK(clk_bF_buf13), .D(AES_CORE_DATAPATH_col_en_cnt_unit_pp1_3__FF_INPUT), .Q(AES_CORE_DATAPATH_col_en_cnt_unit_pp1_3_), .R(rst_n_bF_buf78), .S(1'b1) );
  DFFSR DFFSR_793 ( .CLK(clk_bF_buf12), .D(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_0__FF_INPUT), .Q(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_0_), .R(rst_n_bF_buf77), .S(1'b1) );
  DFFSR DFFSR_794 ( .CLK(clk_bF_buf11), .D(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_1__FF_INPUT), .Q(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_1_), .R(rst_n_bF_buf76), .S(1'b1) );
  DFFSR DFFSR_795 ( .CLK(clk_bF_buf10), .D(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_2__FF_INPUT), .Q(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_2_), .R(rst_n_bF_buf75), .S(1'b1) );
  DFFSR DFFSR_796 ( .CLK(clk_bF_buf9), .D(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_3__FF_INPUT), .Q(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_3_), .R(rst_n_bF_buf74), .S(1'b1) );
  DFFSR DFFSR_797 ( .CLK(clk_bF_buf8), .D(AES_CORE_DATAPATH_key_en_pp1_0__FF_INPUT), .Q(AES_CORE_DATAPATH_key_en_pp1_0_), .R(rst_n_bF_buf73), .S(1'b1) );
  DFFSR DFFSR_798 ( .CLK(clk_bF_buf7), .D(AES_CORE_DATAPATH_key_en_pp1_1__FF_INPUT), .Q(AES_CORE_DATAPATH_key_en_pp1_1_), .R(rst_n_bF_buf72), .S(1'b1) );
  DFFSR DFFSR_799 ( .CLK(clk_bF_buf6), .D(AES_CORE_DATAPATH_key_en_pp1_2__FF_INPUT), .Q(AES_CORE_DATAPATH_key_en_pp1_2_), .R(rst_n_bF_buf71), .S(1'b1) );
  DFFSR DFFSR_8 ( .CLK(clk_bF_buf85), .D(AES_CORE_CONTROL_UNIT__abc_10818_n310), .Q(AES_CORE_CONTROL_UNIT_state_3_), .R(rst_n_bF_buf79), .S(1'b1) );
  DFFSR DFFSR_80 ( .CLK(clk_bF_buf74), .D(AES_CORE_DATAPATH__0key_0__31_0__27_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__27_), .R(rst_n_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_800 ( .CLK(clk_bF_buf5), .D(AES_CORE_DATAPATH_key_en_pp1_3__FF_INPUT), .Q(AES_CORE_DATAPATH_key_en_pp1_3_), .R(rst_n_bF_buf70), .S(1'b1) );
  DFFSR DFFSR_801 ( .CLK(clk_bF_buf4), .D(AES_CORE_CONTROL_UNIT_rd_count_0_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_round_0_), .R(rst_n_bF_buf69), .S(1'b1) );
  DFFSR DFFSR_802 ( .CLK(clk_bF_buf3), .D(AES_CORE_CONTROL_UNIT_rd_count_1_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_round_1_), .R(rst_n_bF_buf68), .S(1'b1) );
  DFFSR DFFSR_803 ( .CLK(clk_bF_buf2), .D(AES_CORE_CONTROL_UNIT_rd_count_2_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_round_2_), .R(rst_n_bF_buf67), .S(1'b1) );
  DFFSR DFFSR_804 ( .CLK(clk_bF_buf1), .D(AES_CORE_CONTROL_UNIT_rd_count_3_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_round_3_), .R(rst_n_bF_buf66), .S(1'b1) );
  DFFSR DFFSR_805 ( .CLK(clk_bF_buf0), .D(AES_CORE_CONTROL_UNIT_col_sel_0_), .Q(AES_CORE_DATAPATH_col_sel_pp1_0_), .R(rst_n_bF_buf65), .S(1'b1) );
  DFFSR DFFSR_806 ( .CLK(clk_bF_buf92), .D(AES_CORE_CONTROL_UNIT_col_sel_1_), .Q(AES_CORE_DATAPATH_col_sel_pp1_1_), .R(1'b1), .S(rst_n_bF_buf64) );
  DFFSR DFFSR_807 ( .CLK(clk_bF_buf91), .D(AES_CORE_DATAPATH_col_sel_pp1_0_), .Q(AES_CORE_DATAPATH_col_sel_pp2_0_), .R(rst_n_bF_buf63), .S(1'b1) );
  DFFSR DFFSR_808 ( .CLK(clk_bF_buf90), .D(AES_CORE_DATAPATH_col_sel_pp1_1_), .Q(AES_CORE_DATAPATH_col_sel_pp2_1_), .R(1'b1), .S(rst_n_bF_buf62) );
  DFFSR DFFSR_809 ( .CLK(clk_bF_buf89), .D(AES_CORE_CONTROL_UNIT_key_out_sel_0_), .Q(AES_CORE_DATAPATH_key_out_sel_pp1_0_), .R(rst_n_bF_buf61), .S(1'b1) );
  DFFSR DFFSR_81 ( .CLK(clk_bF_buf73), .D(AES_CORE_DATAPATH__0key_0__31_0__28_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__28_), .R(rst_n_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_810 ( .CLK(clk_bF_buf88), .D(AES_CORE_CONTROL_UNIT_key_out_sel_1_), .Q(AES_CORE_DATAPATH_key_out_sel_pp1_1_), .R(rst_n_bF_buf60), .S(1'b1) );
  DFFSR DFFSR_811 ( .CLK(clk_bF_buf87), .D(AES_CORE_DATAPATH_key_out_sel_pp1_0_), .Q(AES_CORE_DATAPATH_key_out_sel_pp2_0_), .R(rst_n_bF_buf59), .S(1'b1) );
  DFFSR DFFSR_812 ( .CLK(clk_bF_buf86), .D(AES_CORE_DATAPATH_key_out_sel_pp1_1_), .Q(AES_CORE_DATAPATH_key_out_sel_pp2_1_), .R(rst_n_bF_buf58), .S(1'b1) );
  DFFSR DFFSR_813 ( .CLK(clk_bF_buf85), .D(AES_CORE_CONTROL_UNIT_rk_sel_0_), .Q(AES_CORE_DATAPATH_rk_sel_pp1_0_), .R(rst_n_bF_buf57), .S(1'b1) );
  DFFSR DFFSR_814 ( .CLK(clk_bF_buf84), .D(AES_CORE_CONTROL_UNIT_rk_sel_1_), .Q(AES_CORE_DATAPATH_rk_sel_pp1_1_), .R(rst_n_bF_buf56), .S(1'b1) );
  DFFSR DFFSR_815 ( .CLK(clk_bF_buf83), .D(AES_CORE_DATAPATH_rk_sel_pp1_0_), .Q(AES_CORE_DATAPATH_rk_sel_pp2_0_), .R(rst_n_bF_buf55), .S(1'b1) );
  DFFSR DFFSR_816 ( .CLK(clk_bF_buf82), .D(AES_CORE_DATAPATH_rk_sel_pp1_1_), .Q(AES_CORE_DATAPATH_rk_sel_pp2_1_), .R(rst_n_bF_buf54), .S(1'b1) );
  DFFSR DFFSR_817 ( .CLK(clk_bF_buf81), .D(AES_CORE_CONTROL_UNIT_key_sel), .Q(AES_CORE_DATAPATH_key_sel_pp1), .R(rst_n_bF_buf53), .S(1'b1) );
  DFFSR DFFSR_818 ( .CLK(clk_bF_buf80), .D(AES_CORE_DATAPATH_rk_out_sel), .Q(AES_CORE_DATAPATH_rk_out_sel_pp1), .R(1'b1), .S(rst_n_bF_buf52) );
  DFFSR DFFSR_819 ( .CLK(clk_bF_buf79), .D(AES_CORE_DATAPATH_rk_out_sel_pp1), .Q(AES_CORE_DATAPATH_rk_out_sel_pp2), .R(1'b1), .S(rst_n_bF_buf51) );
  DFFSR DFFSR_82 ( .CLK(clk_bF_buf72), .D(AES_CORE_DATAPATH__0key_0__31_0__29_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__29_), .R(rst_n_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_820 ( .CLK(clk_bF_buf78), .D(AES_CORE_CONTROL_UNIT_last_round_bF_buf5), .Q(AES_CORE_DATAPATH_last_round_pp1), .R(1'b1), .S(rst_n_bF_buf50) );
  DFFSR DFFSR_821 ( .CLK(clk_bF_buf77), .D(AES_CORE_DATAPATH_last_round_pp1), .Q(AES_CORE_DATAPATH_last_round_pp2), .R(rst_n_bF_buf49), .S(1'b1) );
  DFFSR DFFSR_83 ( .CLK(clk_bF_buf71), .D(AES_CORE_DATAPATH__0key_0__31_0__30_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__30_), .R(rst_n_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_84 ( .CLK(clk_bF_buf70), .D(AES_CORE_DATAPATH__0key_0__31_0__31_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__31_), .R(rst_n_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_85 ( .CLK(clk_bF_buf69), .D(AES_CORE_DATAPATH__0key_host_1__31_0__0_), .Q(AES_CORE_DATAPATH_key_host_1__0_), .R(rst_n_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_86 ( .CLK(clk_bF_buf68), .D(AES_CORE_DATAPATH__0key_host_1__31_0__1_), .Q(AES_CORE_DATAPATH_key_host_1__1_), .R(rst_n_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_87 ( .CLK(clk_bF_buf67), .D(AES_CORE_DATAPATH__0key_host_1__31_0__2_), .Q(AES_CORE_DATAPATH_key_host_1__2_), .R(rst_n_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_88 ( .CLK(clk_bF_buf66), .D(AES_CORE_DATAPATH__0key_host_1__31_0__3_), .Q(AES_CORE_DATAPATH_key_host_1__3_), .R(rst_n_bF_buf86), .S(1'b1) );
  DFFSR DFFSR_89 ( .CLK(clk_bF_buf65), .D(AES_CORE_DATAPATH__0key_host_1__31_0__4_), .Q(AES_CORE_DATAPATH_key_host_1__4_), .R(rst_n_bF_buf85), .S(1'b1) );
  DFFSR DFFSR_9 ( .CLK(clk_bF_buf84), .D(AES_CORE_CONTROL_UNIT__abc_10818_n109), .Q(AES_CORE_CONTROL_UNIT_state_4_), .R(rst_n_bF_buf78), .S(1'b1) );
  DFFSR DFFSR_90 ( .CLK(clk_bF_buf64), .D(AES_CORE_DATAPATH__0key_host_1__31_0__5_), .Q(AES_CORE_DATAPATH_key_host_1__5_), .R(rst_n_bF_buf84), .S(1'b1) );
  DFFSR DFFSR_91 ( .CLK(clk_bF_buf63), .D(AES_CORE_DATAPATH__0key_host_1__31_0__6_), .Q(AES_CORE_DATAPATH_key_host_1__6_), .R(rst_n_bF_buf83), .S(1'b1) );
  DFFSR DFFSR_92 ( .CLK(clk_bF_buf62), .D(AES_CORE_DATAPATH__0key_host_1__31_0__7_), .Q(AES_CORE_DATAPATH_key_host_1__7_), .R(rst_n_bF_buf82), .S(1'b1) );
  DFFSR DFFSR_93 ( .CLK(clk_bF_buf61), .D(AES_CORE_DATAPATH__0key_host_1__31_0__8_), .Q(AES_CORE_DATAPATH_key_host_1__8_), .R(rst_n_bF_buf81), .S(1'b1) );
  DFFSR DFFSR_94 ( .CLK(clk_bF_buf60), .D(AES_CORE_DATAPATH__0key_host_1__31_0__9_), .Q(AES_CORE_DATAPATH_key_host_1__9_), .R(rst_n_bF_buf80), .S(1'b1) );
  DFFSR DFFSR_95 ( .CLK(clk_bF_buf59), .D(AES_CORE_DATAPATH__0key_host_1__31_0__10_), .Q(AES_CORE_DATAPATH_key_host_1__10_), .R(rst_n_bF_buf79), .S(1'b1) );
  DFFSR DFFSR_96 ( .CLK(clk_bF_buf58), .D(AES_CORE_DATAPATH__0key_host_1__31_0__11_), .Q(AES_CORE_DATAPATH_key_host_1__11_), .R(rst_n_bF_buf78), .S(1'b1) );
  DFFSR DFFSR_97 ( .CLK(clk_bF_buf57), .D(AES_CORE_DATAPATH__0key_host_1__31_0__12_), .Q(AES_CORE_DATAPATH_key_host_1__12_), .R(rst_n_bF_buf77), .S(1'b1) );
  DFFSR DFFSR_98 ( .CLK(clk_bF_buf56), .D(AES_CORE_DATAPATH__0key_host_1__31_0__13_), .Q(AES_CORE_DATAPATH_key_host_1__13_), .R(rst_n_bF_buf76), .S(1'b1) );
  DFFSR DFFSR_99 ( .CLK(clk_bF_buf55), .D(AES_CORE_DATAPATH__0key_host_1__31_0__14_), .Q(AES_CORE_DATAPATH_key_host_1__14_), .R(rst_n_bF_buf75), .S(1'b1) );
  INVX1 INVX1_1 ( .A(\addr[1] ), .Y(_abc_15830_n11_1) );
  INVX1 INVX1_10 ( .A(AES_CORE_CONTROL_UNIT_state_13_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n104) );
  INVX1 INVX1_100 ( .A(AES_CORE_DATAPATH__abc_16259_n3337), .Y(AES_CORE_DATAPATH__abc_16259_n3338) );
  INVX1 INVX1_1000 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n180), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n181) );
  INVX1 INVX1_1001 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n156), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n186) );
  INVX1 INVX1_1002 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n163), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n187_1) );
  INVX1 INVX1_1003 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n196) );
  INVX1 INVX1_1004 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n198) );
  INVX1 INVX1_1005 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n200), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n201) );
  INVX1 INVX1_1006 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n208), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n209) );
  INVX1 INVX1_1007 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n162), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n213) );
  INVX1 INVX1_1008 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n218) );
  INVX1 INVX1_1009 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n220) );
  INVX1 INVX1_101 ( .A(AES_CORE_DATAPATH__abc_16259_n3340), .Y(AES_CORE_DATAPATH__abc_16259_n3341) );
  INVX1 INVX1_1010 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n222), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n232) );
  INVX1 INVX1_1011 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n246), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n247) );
  INVX1 INVX1_1012 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n249), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n250) );
  INVX1 INVX1_1013 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n259) );
  INVX1 INVX1_1014 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n261) );
  INVX1 INVX1_1015 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n263), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n264) );
  INVX1 INVX1_1016 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n265), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n266) );
  INVX1 INVX1_1017 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n267) );
  INVX1 INVX1_1018 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n269) );
  INVX1 INVX1_1019 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n271), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n272) );
  INVX1 INVX1_102 ( .A(AES_CORE_DATAPATH_col_0__13_), .Y(AES_CORE_DATAPATH__abc_16259_n3353) );
  INVX1 INVX1_1020 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n273), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n275) );
  INVX1 INVX1_1021 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n284), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n285) );
  INVX1 INVX1_1022 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n282), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n289) );
  INVX1 INVX1_1023 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n292), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n293) );
  INVX1 INVX1_1024 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n277), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n295) );
  INVX1 INVX1_1025 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n303), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n304) );
  INVX1 INVX1_1026 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n306), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n307) );
  INVX1 INVX1_1027 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n310), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n311) );
  INVX1 INVX1_1028 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n297), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n313) );
  INVX1 INVX1_1029 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n315), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n318) );
  INVX1 INVX1_103 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_13_), .Y(AES_CORE_DATAPATH__abc_16259_n3355_1) );
  INVX1 INVX1_1030 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n321), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n322) );
  INVX1 INVX1_1031 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n323), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n324) );
  INVX1 INVX1_1032 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n327), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n328) );
  INVX1 INVX1_1033 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n330), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n331) );
  INVX1 INVX1_1034 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n333), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n335) );
  INVX1 INVX1_1035 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n337), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n338) );
  INVX1 INVX1_1036 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n344), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n345) );
  INVX1 INVX1_1037 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n347), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n348) );
  INVX1 INVX1_1038 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n352), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n353) );
  INVX1 INVX1_1039 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n356), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_1_2_) );
  INVX1 INVX1_104 ( .A(AES_CORE_DATAPATH__abc_16259_n3362), .Y(AES_CORE_DATAPATH__abc_16259_n3363) );
  INVX1 INVX1_1040 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n358), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n360) );
  INVX1 INVX1_1041 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n379), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n380) );
  INVX1 INVX1_1042 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n382), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n383) );
  INVX1 INVX1_1043 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n401) );
  INVX1 INVX1_1044 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n407), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n409) );
  INVX1 INVX1_1045 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n412), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n413) );
  INVX1 INVX1_1046 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n316), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n441) );
  INVX1 INVX1_1047 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n461), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_1_) );
  INVX1 INVX1_1048 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n469) );
  INVX1 INVX1_1049 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n470), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n471) );
  INVX1 INVX1_105 ( .A(AES_CORE_DATAPATH__abc_16259_n3377), .Y(AES_CORE_DATAPATH__abc_16259_n3378) );
  INVX1 INVX1_1050 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n472) );
  INVX1 INVX1_1051 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n478), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n479) );
  INVX1 INVX1_1052 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n484), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n485) );
  INVX1 INVX1_1053 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n486) );
  INVX1 INVX1_1054 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n493) );
  INVX1 INVX1_1055 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n497), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n498) );
  INVX1 INVX1_1056 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n501), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n502) );
  INVX1 INVX1_1057 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n504), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n505) );
  INVX1 INVX1_1058 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n481), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n507) );
  INVX1 INVX1_1059 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n475), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n510) );
  INVX1 INVX1_106 ( .A(AES_CORE_DATAPATH__abc_16259_n3380_1), .Y(AES_CORE_DATAPATH__abc_16259_n3381_1) );
  INVX1 INVX1_1060 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n512), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n513) );
  INVX1 INVX1_1061 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n514), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n515) );
  INVX1 INVX1_1062 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n524), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n525) );
  INVX1 INVX1_1063 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n529), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n542) );
  INVX1 INVX1_1064 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n550), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n551) );
  INVX1 INVX1_1065 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n552), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n553) );
  INVX1 INVX1_1066 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n555), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n556) );
  INVX1 INVX1_1067 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n548), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n558) );
  INVX1 INVX1_1068 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n567), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n568) );
  INVX1 INVX1_1069 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n569), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n570) );
  INVX1 INVX1_107 ( .A(AES_CORE_DATAPATH_col_0__14_), .Y(AES_CORE_DATAPATH__abc_16259_n3393) );
  INVX1 INVX1_1070 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n573), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n575) );
  INVX1 INVX1_1071 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n577), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n578) );
  INVX1 INVX1_1072 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n583) );
  INVX1 INVX1_1073 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n50) );
  INVX1 INVX1_1074 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n52) );
  INVX1 INVX1_1075 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n54_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n55) );
  INVX1 INVX1_1076 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n56) );
  INVX1 INVX1_1077 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n58) );
  INVX1 INVX1_1078 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n60), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n61) );
  INVX1 INVX1_1079 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n67) );
  INVX1 INVX1_108 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_14_), .Y(AES_CORE_DATAPATH__abc_16259_n3395) );
  INVX1 INVX1_1080 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n72) );
  INVX1 INVX1_1081 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n70), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n73) );
  INVX1 INVX1_1082 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n79) );
  INVX1 INVX1_1083 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n86_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n87) );
  INVX1 INVX1_1084 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n92), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n93) );
  INVX1 INVX1_1085 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n95), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n96) );
  INVX1 INVX1_1086 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n104_1) );
  INVX1 INVX1_1087 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n107), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n109) );
  INVX1 INVX1_1088 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n112), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n113) );
  INVX1 INVX1_1089 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n114), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_7_) );
  INVX1 INVX1_109 ( .A(AES_CORE_DATAPATH__abc_16259_n3402_1), .Y(AES_CORE_DATAPATH__abc_16259_n3403) );
  INVX1 INVX1_1090 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n116), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n117) );
  INVX1 INVX1_1091 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n121_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n122) );
  INVX1 INVX1_1092 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n126_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_0_) );
  INVX1 INVX1_1093 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n130), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n131) );
  INVX1 INVX1_1094 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n140), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_2_) );
  INVX1 INVX1_1095 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n102), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n142) );
  INVX1 INVX1_1096 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n149), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n150_1) );
  INVX1 INVX1_1097 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n157), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n158) );
  INVX1 INVX1_1098 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n159) );
  INVX1 INVX1_1099 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n161) );
  INVX1 INVX1_11 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n111), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n112) );
  INVX1 INVX1_110 ( .A(AES_CORE_DATAPATH__abc_16259_n3417_1), .Y(AES_CORE_DATAPATH__abc_16259_n3418) );
  INVX1 INVX1_1100 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n167), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n168) );
  INVX1 INVX1_1101 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n173), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n174) );
  INVX1 INVX1_1102 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n164), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n175) );
  INVX1 INVX1_1103 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n176_1) );
  INVX1 INVX1_1104 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n180), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n181) );
  INVX1 INVX1_1105 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n156), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n186) );
  INVX1 INVX1_1106 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n163), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n187_1) );
  INVX1 INVX1_1107 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n196) );
  INVX1 INVX1_1108 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n198) );
  INVX1 INVX1_1109 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n200), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n201) );
  INVX1 INVX1_111 ( .A(AES_CORE_DATAPATH__abc_16259_n3420), .Y(AES_CORE_DATAPATH__abc_16259_n3421) );
  INVX1 INVX1_1110 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n208), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n209) );
  INVX1 INVX1_1111 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n162), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n213) );
  INVX1 INVX1_1112 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n218) );
  INVX1 INVX1_1113 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n220) );
  INVX1 INVX1_1114 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n222), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n232) );
  INVX1 INVX1_1115 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n246), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n247) );
  INVX1 INVX1_1116 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n249), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n250) );
  INVX1 INVX1_1117 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n259) );
  INVX1 INVX1_1118 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n261) );
  INVX1 INVX1_1119 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n263), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n264) );
  INVX1 INVX1_112 ( .A(AES_CORE_DATAPATH_col_0__15_), .Y(AES_CORE_DATAPATH__abc_16259_n3433_1) );
  INVX1 INVX1_1120 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n265), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n266) );
  INVX1 INVX1_1121 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n267) );
  INVX1 INVX1_1122 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n269) );
  INVX1 INVX1_1123 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n271), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n272) );
  INVX1 INVX1_1124 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n273), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n275) );
  INVX1 INVX1_1125 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n284), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n285) );
  INVX1 INVX1_1126 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n282), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n289) );
  INVX1 INVX1_1127 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n292), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n293) );
  INVX1 INVX1_1128 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n277), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n295) );
  INVX1 INVX1_1129 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n303), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n304) );
  INVX1 INVX1_113 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_15_), .Y(AES_CORE_DATAPATH__abc_16259_n3435) );
  INVX1 INVX1_1130 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n306), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n307) );
  INVX1 INVX1_1131 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n310), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n311) );
  INVX1 INVX1_1132 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n297), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n313) );
  INVX1 INVX1_1133 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n315), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n318) );
  INVX1 INVX1_1134 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n321), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n322) );
  INVX1 INVX1_1135 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n323), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n324) );
  INVX1 INVX1_1136 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n327), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n328) );
  INVX1 INVX1_1137 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n330), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n331) );
  INVX1 INVX1_1138 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n333), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n335) );
  INVX1 INVX1_1139 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n337), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n338) );
  INVX1 INVX1_114 ( .A(AES_CORE_DATAPATH__abc_16259_n3442_1), .Y(AES_CORE_DATAPATH__abc_16259_n3443) );
  INVX1 INVX1_1140 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n344), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n345) );
  INVX1 INVX1_1141 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n347), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n348) );
  INVX1 INVX1_1142 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n352), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n353) );
  INVX1 INVX1_1143 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n356), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_1_2_) );
  INVX1 INVX1_1144 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n358), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n360) );
  INVX1 INVX1_1145 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n379), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n380) );
  INVX1 INVX1_1146 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n382), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n383) );
  INVX1 INVX1_1147 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_13_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n401) );
  INVX1 INVX1_1148 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n407), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n409) );
  INVX1 INVX1_1149 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n412), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n413) );
  INVX1 INVX1_115 ( .A(AES_CORE_DATAPATH__abc_16259_n3457), .Y(AES_CORE_DATAPATH__abc_16259_n3458) );
  INVX1 INVX1_1150 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n316), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n441) );
  INVX1 INVX1_1151 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n461), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_1_) );
  INVX1 INVX1_1152 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n469) );
  INVX1 INVX1_1153 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n470), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n471) );
  INVX1 INVX1_1154 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n472) );
  INVX1 INVX1_1155 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n478), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n479) );
  INVX1 INVX1_1156 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n484), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n485) );
  INVX1 INVX1_1157 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n486) );
  INVX1 INVX1_1158 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n493) );
  INVX1 INVX1_1159 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n497), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n498) );
  INVX1 INVX1_116 ( .A(AES_CORE_DATAPATH__abc_16259_n3460_1), .Y(AES_CORE_DATAPATH__abc_16259_n3461) );
  INVX1 INVX1_1160 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n501), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n502) );
  INVX1 INVX1_1161 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n504), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n505) );
  INVX1 INVX1_1162 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n481), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n507) );
  INVX1 INVX1_1163 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n475), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n510) );
  INVX1 INVX1_1164 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n512), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n513) );
  INVX1 INVX1_1165 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n514), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n515) );
  INVX1 INVX1_1166 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n524), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n525) );
  INVX1 INVX1_1167 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n529), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n542) );
  INVX1 INVX1_1168 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n550), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n551) );
  INVX1 INVX1_1169 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n552), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n553) );
  INVX1 INVX1_117 ( .A(AES_CORE_DATAPATH_col_0__16_), .Y(AES_CORE_DATAPATH__abc_16259_n3473_1) );
  INVX1 INVX1_1170 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n555), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n556) );
  INVX1 INVX1_1171 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n548), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n558) );
  INVX1 INVX1_1172 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n567), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n568) );
  INVX1 INVX1_1173 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n569), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n570) );
  INVX1 INVX1_1174 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n573), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n575) );
  INVX1 INVX1_1175 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n577), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n578) );
  INVX1 INVX1_1176 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_9_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n583) );
  INVX1 INVX1_1177 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n50) );
  INVX1 INVX1_1178 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n52) );
  INVX1 INVX1_1179 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n54_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n55) );
  INVX1 INVX1_118 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_16_), .Y(AES_CORE_DATAPATH__abc_16259_n3475_1) );
  INVX1 INVX1_1180 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n56) );
  INVX1 INVX1_1181 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n58) );
  INVX1 INVX1_1182 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n60), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n61) );
  INVX1 INVX1_1183 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n67) );
  INVX1 INVX1_1184 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n72) );
  INVX1 INVX1_1185 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n70), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n73) );
  INVX1 INVX1_1186 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n79) );
  INVX1 INVX1_1187 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n86_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n87) );
  INVX1 INVX1_1188 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n92), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n93) );
  INVX1 INVX1_1189 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n95), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n96) );
  INVX1 INVX1_119 ( .A(AES_CORE_DATAPATH__abc_16259_n3482), .Y(AES_CORE_DATAPATH__abc_16259_n3483) );
  INVX1 INVX1_1190 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n104_1) );
  INVX1 INVX1_1191 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n107), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n109) );
  INVX1 INVX1_1192 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n112), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n113) );
  INVX1 INVX1_1193 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n114), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_7_) );
  INVX1 INVX1_1194 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n116), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n117) );
  INVX1 INVX1_1195 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n121_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n122) );
  INVX1 INVX1_1196 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n126_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_0_) );
  INVX1 INVX1_1197 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n130), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n131) );
  INVX1 INVX1_1198 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n140), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_2_) );
  INVX1 INVX1_1199 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n102), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n142) );
  INVX1 INVX1_12 ( .A(start), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n131) );
  INVX1 INVX1_120 ( .A(AES_CORE_DATAPATH__abc_16259_n3497_1), .Y(AES_CORE_DATAPATH__abc_16259_n3498) );
  INVX1 INVX1_1200 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n149), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n150_1) );
  INVX1 INVX1_1201 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n157), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n158) );
  INVX1 INVX1_1202 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n159) );
  INVX1 INVX1_1203 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n161) );
  INVX1 INVX1_1204 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n167), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n168) );
  INVX1 INVX1_1205 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n173), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n174) );
  INVX1 INVX1_1206 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n164), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n175) );
  INVX1 INVX1_1207 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n176_1) );
  INVX1 INVX1_1208 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n180), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n181) );
  INVX1 INVX1_1209 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n156), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n186) );
  INVX1 INVX1_121 ( .A(AES_CORE_DATAPATH__abc_16259_n3500_1), .Y(AES_CORE_DATAPATH__abc_16259_n3501) );
  INVX1 INVX1_1210 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n163), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n187_1) );
  INVX1 INVX1_1211 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n196) );
  INVX1 INVX1_1212 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n198) );
  INVX1 INVX1_1213 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n200), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n201) );
  INVX1 INVX1_1214 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n208), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n209) );
  INVX1 INVX1_1215 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n162), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n213) );
  INVX1 INVX1_1216 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n218) );
  INVX1 INVX1_1217 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n220) );
  INVX1 INVX1_1218 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n222), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n232) );
  INVX1 INVX1_1219 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n246), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n247) );
  INVX1 INVX1_122 ( .A(AES_CORE_DATAPATH_col_0__17_), .Y(AES_CORE_DATAPATH__abc_16259_n3513) );
  INVX1 INVX1_1220 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n249), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n250) );
  INVX1 INVX1_1221 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n259) );
  INVX1 INVX1_1222 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n261) );
  INVX1 INVX1_1223 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n263), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n264) );
  INVX1 INVX1_1224 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n265), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n266) );
  INVX1 INVX1_1225 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n267) );
  INVX1 INVX1_1226 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n269) );
  INVX1 INVX1_1227 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n271), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n272) );
  INVX1 INVX1_1228 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n273), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n275) );
  INVX1 INVX1_1229 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n284), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n285) );
  INVX1 INVX1_123 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_17_), .Y(AES_CORE_DATAPATH__abc_16259_n3515) );
  INVX1 INVX1_1230 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n282), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n289) );
  INVX1 INVX1_1231 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n292), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n293) );
  INVX1 INVX1_1232 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n277), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n295) );
  INVX1 INVX1_1233 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n303), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n304) );
  INVX1 INVX1_1234 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n306), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n307) );
  INVX1 INVX1_1235 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n310), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n311) );
  INVX1 INVX1_1236 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n297), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n313) );
  INVX1 INVX1_1237 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n315), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n318) );
  INVX1 INVX1_1238 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n321), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n322) );
  INVX1 INVX1_1239 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n323), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n324) );
  INVX1 INVX1_124 ( .A(AES_CORE_DATAPATH__abc_16259_n3522), .Y(AES_CORE_DATAPATH__abc_16259_n3523) );
  INVX1 INVX1_1240 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n327), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n328) );
  INVX1 INVX1_1241 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n330), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n331) );
  INVX1 INVX1_1242 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n333), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n335) );
  INVX1 INVX1_1243 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n337), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n338) );
  INVX1 INVX1_1244 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n344), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n345) );
  INVX1 INVX1_1245 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n347), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n348) );
  INVX1 INVX1_1246 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n352), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n353) );
  INVX1 INVX1_1247 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n356), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_1_2_) );
  INVX1 INVX1_1248 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n358), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n360) );
  INVX1 INVX1_1249 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n379), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n380) );
  INVX1 INVX1_125 ( .A(AES_CORE_DATAPATH__abc_16259_n3537), .Y(AES_CORE_DATAPATH__abc_16259_n3538) );
  INVX1 INVX1_1250 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n382), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n383) );
  INVX1 INVX1_1251 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_21_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n401) );
  INVX1 INVX1_1252 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n407), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n409) );
  INVX1 INVX1_1253 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n412), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n413) );
  INVX1 INVX1_1254 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n316), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n441) );
  INVX1 INVX1_1255 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n461), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_1_) );
  INVX1 INVX1_1256 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n469) );
  INVX1 INVX1_1257 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n470), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n471) );
  INVX1 INVX1_1258 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n472) );
  INVX1 INVX1_1259 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n478), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n479) );
  INVX1 INVX1_126 ( .A(AES_CORE_DATAPATH__abc_16259_n3540), .Y(AES_CORE_DATAPATH__abc_16259_n3541) );
  INVX1 INVX1_1260 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n484), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n485) );
  INVX1 INVX1_1261 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n486) );
  INVX1 INVX1_1262 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n493) );
  INVX1 INVX1_1263 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n497), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n498) );
  INVX1 INVX1_1264 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n501), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n502) );
  INVX1 INVX1_1265 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n504), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n505) );
  INVX1 INVX1_1266 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n481), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n507) );
  INVX1 INVX1_1267 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n475), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n510) );
  INVX1 INVX1_1268 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n512), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n513) );
  INVX1 INVX1_1269 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n514), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n515) );
  INVX1 INVX1_127 ( .A(AES_CORE_DATAPATH_col_0__18_), .Y(AES_CORE_DATAPATH__abc_16259_n3553) );
  INVX1 INVX1_1270 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n524), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n525) );
  INVX1 INVX1_1271 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n529), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n542) );
  INVX1 INVX1_1272 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n550), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n551) );
  INVX1 INVX1_1273 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n552), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n553) );
  INVX1 INVX1_1274 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n555), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n556) );
  INVX1 INVX1_1275 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n548), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n558) );
  INVX1 INVX1_1276 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n567), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n568) );
  INVX1 INVX1_1277 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n569), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n570) );
  INVX1 INVX1_1278 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n573), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n575) );
  INVX1 INVX1_1279 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n577), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n578) );
  INVX1 INVX1_128 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_18_), .Y(AES_CORE_DATAPATH__abc_16259_n3555_1) );
  INVX1 INVX1_1280 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_17_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n583) );
  INVX1 INVX1_1281 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n50) );
  INVX1 INVX1_1282 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n52) );
  INVX1 INVX1_1283 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n54_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n55) );
  INVX1 INVX1_1284 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n56) );
  INVX1 INVX1_1285 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n58) );
  INVX1 INVX1_1286 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n60), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n61) );
  INVX1 INVX1_1287 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n67) );
  INVX1 INVX1_1288 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n72) );
  INVX1 INVX1_1289 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n70), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n73) );
  INVX1 INVX1_129 ( .A(AES_CORE_DATAPATH__abc_16259_n3562_1), .Y(AES_CORE_DATAPATH__abc_16259_n3563) );
  INVX1 INVX1_1290 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n79) );
  INVX1 INVX1_1291 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n86_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n87) );
  INVX1 INVX1_1292 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n92), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n93) );
  INVX1 INVX1_1293 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n95), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n96) );
  INVX1 INVX1_1294 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n104_1) );
  INVX1 INVX1_1295 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n107), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n109) );
  INVX1 INVX1_1296 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n112), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n113) );
  INVX1 INVX1_1297 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n114), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_7_) );
  INVX1 INVX1_1298 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n116), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n117) );
  INVX1 INVX1_1299 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n121_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n122) );
  INVX1 INVX1_13 ( .A(AES_CORE_CONTROL_UNIT_last_round_bF_buf4), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n142) );
  INVX1 INVX1_130 ( .A(AES_CORE_DATAPATH__abc_16259_n3577), .Y(AES_CORE_DATAPATH__abc_16259_n3578_1) );
  INVX1 INVX1_1300 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n126_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_0_) );
  INVX1 INVX1_1301 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n130), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n131) );
  INVX1 INVX1_1302 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n140), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_2_) );
  INVX1 INVX1_1303 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n102), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n142) );
  INVX1 INVX1_1304 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n149), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n150_1) );
  INVX1 INVX1_1305 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n157), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n158) );
  INVX1 INVX1_1306 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n159) );
  INVX1 INVX1_1307 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n161) );
  INVX1 INVX1_1308 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n167), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n168) );
  INVX1 INVX1_1309 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n173), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n174) );
  INVX1 INVX1_131 ( .A(AES_CORE_DATAPATH__abc_16259_n3580), .Y(AES_CORE_DATAPATH__abc_16259_n3581) );
  INVX1 INVX1_1310 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n164), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n175) );
  INVX1 INVX1_1311 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n176_1) );
  INVX1 INVX1_1312 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n180), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n181) );
  INVX1 INVX1_1313 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n156), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n186) );
  INVX1 INVX1_1314 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n163), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n187_1) );
  INVX1 INVX1_1315 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n196) );
  INVX1 INVX1_1316 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n198) );
  INVX1 INVX1_1317 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n200), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n201) );
  INVX1 INVX1_1318 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n208), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n209) );
  INVX1 INVX1_1319 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n162), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n213) );
  INVX1 INVX1_132 ( .A(AES_CORE_DATAPATH_col_0__19_), .Y(AES_CORE_DATAPATH__abc_16259_n3593_1) );
  INVX1 INVX1_1320 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n218) );
  INVX1 INVX1_1321 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n220) );
  INVX1 INVX1_1322 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n222), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n232) );
  INVX1 INVX1_1323 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n246), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n247) );
  INVX1 INVX1_1324 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n249), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n250) );
  INVX1 INVX1_1325 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n259) );
  INVX1 INVX1_1326 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n261) );
  INVX1 INVX1_1327 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n263), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n264) );
  INVX1 INVX1_1328 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n265), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n266) );
  INVX1 INVX1_1329 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n267) );
  INVX1 INVX1_133 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_19_), .Y(AES_CORE_DATAPATH__abc_16259_n3595) );
  INVX1 INVX1_1330 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n269) );
  INVX1 INVX1_1331 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n271), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n272) );
  INVX1 INVX1_1332 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n273), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n275) );
  INVX1 INVX1_1333 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n284), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n285) );
  INVX1 INVX1_1334 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n282), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n289) );
  INVX1 INVX1_1335 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n292), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n293) );
  INVX1 INVX1_1336 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n277), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n295) );
  INVX1 INVX1_1337 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n303), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n304) );
  INVX1 INVX1_1338 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n306), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n307) );
  INVX1 INVX1_1339 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n310), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n311) );
  INVX1 INVX1_134 ( .A(AES_CORE_DATAPATH__abc_16259_n3602), .Y(AES_CORE_DATAPATH__abc_16259_n3603) );
  INVX1 INVX1_1340 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n297), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n313) );
  INVX1 INVX1_1341 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n315), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n318) );
  INVX1 INVX1_1342 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n321), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n322) );
  INVX1 INVX1_1343 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n323), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n324) );
  INVX1 INVX1_1344 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n327), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n328) );
  INVX1 INVX1_1345 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n330), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n331) );
  INVX1 INVX1_1346 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n333), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n335) );
  INVX1 INVX1_1347 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n337), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n338) );
  INVX1 INVX1_1348 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n344), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n345) );
  INVX1 INVX1_1349 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n347), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n348) );
  INVX1 INVX1_135 ( .A(AES_CORE_DATAPATH__abc_16259_n3617), .Y(AES_CORE_DATAPATH__abc_16259_n3618_1) );
  INVX1 INVX1_1350 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n352), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n353) );
  INVX1 INVX1_1351 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n356), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_1_2_) );
  INVX1 INVX1_1352 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n358), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n360) );
  INVX1 INVX1_1353 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n379), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n380) );
  INVX1 INVX1_1354 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n382), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n383) );
  INVX1 INVX1_1355 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_29_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n401) );
  INVX1 INVX1_1356 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n407), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n409) );
  INVX1 INVX1_1357 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n412), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n413) );
  INVX1 INVX1_1358 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n316), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n441) );
  INVX1 INVX1_1359 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n461), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_1_) );
  INVX1 INVX1_136 ( .A(AES_CORE_DATAPATH__abc_16259_n3620_1), .Y(AES_CORE_DATAPATH__abc_16259_n3621) );
  INVX1 INVX1_1360 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n469) );
  INVX1 INVX1_1361 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n470), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n471) );
  INVX1 INVX1_1362 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n472) );
  INVX1 INVX1_1363 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n478), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n479) );
  INVX1 INVX1_1364 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n484), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n485) );
  INVX1 INVX1_1365 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n486) );
  INVX1 INVX1_1366 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n493) );
  INVX1 INVX1_1367 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n497), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n498) );
  INVX1 INVX1_1368 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n501), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n502) );
  INVX1 INVX1_1369 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n504), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n505) );
  INVX1 INVX1_137 ( .A(AES_CORE_DATAPATH_col_0__20_), .Y(AES_CORE_DATAPATH__abc_16259_n3633) );
  INVX1 INVX1_1370 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n481), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n507) );
  INVX1 INVX1_1371 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n475), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n510) );
  INVX1 INVX1_1372 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n512), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n513) );
  INVX1 INVX1_1373 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n514), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n515) );
  INVX1 INVX1_1374 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n524), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n525) );
  INVX1 INVX1_1375 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n529), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n542) );
  INVX1 INVX1_1376 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n550), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n551) );
  INVX1 INVX1_1377 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n552), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n553) );
  INVX1 INVX1_1378 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n555), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n556) );
  INVX1 INVX1_1379 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n548), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n558) );
  INVX1 INVX1_138 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_20_), .Y(AES_CORE_DATAPATH__abc_16259_n3635) );
  INVX1 INVX1_1380 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n567), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n568) );
  INVX1 INVX1_1381 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n569), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n570) );
  INVX1 INVX1_1382 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n573), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n575) );
  INVX1 INVX1_1383 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n577), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n578) );
  INVX1 INVX1_1384 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_25_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n583) );
  INVX1 INVX1_1385 ( .A(\data_type[0] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n69) );
  INVX1 INVX1_1386 ( .A(\data_type[1] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n73) );
  INVX1 INVX1_1387 ( .A(\data_type[0] ), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n69) );
  INVX1 INVX1_1388 ( .A(\data_type[1] ), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n73) );
  INVX1 INVX1_139 ( .A(AES_CORE_DATAPATH__abc_16259_n3642_1), .Y(AES_CORE_DATAPATH__abc_16259_n3643) );
  INVX1 INVX1_14 ( .A(AES_CORE_CONTROL_UNIT_state_0_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n163) );
  INVX1 INVX1_140 ( .A(AES_CORE_DATAPATH__abc_16259_n3657), .Y(AES_CORE_DATAPATH__abc_16259_n3658) );
  INVX1 INVX1_141 ( .A(AES_CORE_DATAPATH__abc_16259_n3660), .Y(AES_CORE_DATAPATH__abc_16259_n3661) );
  INVX1 INVX1_142 ( .A(AES_CORE_DATAPATH_col_0__21_), .Y(AES_CORE_DATAPATH__abc_16259_n3673_1) );
  INVX1 INVX1_143 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_21_), .Y(AES_CORE_DATAPATH__abc_16259_n3675) );
  INVX1 INVX1_144 ( .A(AES_CORE_DATAPATH__abc_16259_n3682), .Y(AES_CORE_DATAPATH__abc_16259_n3683) );
  INVX1 INVX1_145 ( .A(AES_CORE_DATAPATH__abc_16259_n3697_1), .Y(AES_CORE_DATAPATH__abc_16259_n3698) );
  INVX1 INVX1_146 ( .A(AES_CORE_DATAPATH__abc_16259_n3700), .Y(AES_CORE_DATAPATH__abc_16259_n3701) );
  INVX1 INVX1_147 ( .A(AES_CORE_DATAPATH_col_0__22_), .Y(AES_CORE_DATAPATH__abc_16259_n3713_1) );
  INVX1 INVX1_148 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_22_), .Y(AES_CORE_DATAPATH__abc_16259_n3715) );
  INVX1 INVX1_149 ( .A(AES_CORE_DATAPATH__abc_16259_n3722), .Y(AES_CORE_DATAPATH__abc_16259_n3723) );
  INVX1 INVX1_15 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n164), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n165) );
  INVX1 INVX1_150 ( .A(AES_CORE_DATAPATH__abc_16259_n3737_1), .Y(AES_CORE_DATAPATH__abc_16259_n3738) );
  INVX1 INVX1_151 ( .A(AES_CORE_DATAPATH__abc_16259_n3740), .Y(AES_CORE_DATAPATH__abc_16259_n3741) );
  INVX1 INVX1_152 ( .A(AES_CORE_DATAPATH_col_0__23_), .Y(AES_CORE_DATAPATH__abc_16259_n3753_1) );
  INVX1 INVX1_153 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_23_), .Y(AES_CORE_DATAPATH__abc_16259_n3755) );
  INVX1 INVX1_154 ( .A(AES_CORE_DATAPATH__abc_16259_n3762), .Y(AES_CORE_DATAPATH__abc_16259_n3763) );
  INVX1 INVX1_155 ( .A(AES_CORE_DATAPATH__abc_16259_n3777_1), .Y(AES_CORE_DATAPATH__abc_16259_n3778) );
  INVX1 INVX1_156 ( .A(AES_CORE_DATAPATH__abc_16259_n3780), .Y(AES_CORE_DATAPATH__abc_16259_n3781) );
  INVX1 INVX1_157 ( .A(AES_CORE_DATAPATH_col_0__24_), .Y(AES_CORE_DATAPATH__abc_16259_n3793_1) );
  INVX1 INVX1_158 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_24_), .Y(AES_CORE_DATAPATH__abc_16259_n3795) );
  INVX1 INVX1_159 ( .A(AES_CORE_DATAPATH__abc_16259_n3802), .Y(AES_CORE_DATAPATH__abc_16259_n3803) );
  INVX1 INVX1_16 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n169), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n170) );
  INVX1 INVX1_160 ( .A(AES_CORE_DATAPATH__abc_16259_n3817_1), .Y(AES_CORE_DATAPATH__abc_16259_n3818) );
  INVX1 INVX1_161 ( .A(AES_CORE_DATAPATH__abc_16259_n3820), .Y(AES_CORE_DATAPATH__abc_16259_n3821) );
  INVX1 INVX1_162 ( .A(AES_CORE_DATAPATH_col_0__25_), .Y(AES_CORE_DATAPATH__abc_16259_n3833_1) );
  INVX1 INVX1_163 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_25_), .Y(AES_CORE_DATAPATH__abc_16259_n3835) );
  INVX1 INVX1_164 ( .A(AES_CORE_DATAPATH__abc_16259_n3842), .Y(AES_CORE_DATAPATH__abc_16259_n3843) );
  INVX1 INVX1_165 ( .A(AES_CORE_DATAPATH__abc_16259_n3857_1), .Y(AES_CORE_DATAPATH__abc_16259_n3858) );
  INVX1 INVX1_166 ( .A(AES_CORE_DATAPATH__abc_16259_n3860), .Y(AES_CORE_DATAPATH__abc_16259_n3861) );
  INVX1 INVX1_167 ( .A(AES_CORE_DATAPATH_col_0__26_), .Y(AES_CORE_DATAPATH__abc_16259_n3873_1) );
  INVX1 INVX1_168 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_26_), .Y(AES_CORE_DATAPATH__abc_16259_n3875) );
  INVX1 INVX1_169 ( .A(AES_CORE_DATAPATH__abc_16259_n3882), .Y(AES_CORE_DATAPATH__abc_16259_n3883) );
  INVX1 INVX1_17 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n173), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n174) );
  INVX1 INVX1_170 ( .A(AES_CORE_DATAPATH__abc_16259_n3897_1), .Y(AES_CORE_DATAPATH__abc_16259_n3898) );
  INVX1 INVX1_171 ( .A(AES_CORE_DATAPATH__abc_16259_n3900), .Y(AES_CORE_DATAPATH__abc_16259_n3901) );
  INVX1 INVX1_172 ( .A(AES_CORE_DATAPATH_col_0__27_), .Y(AES_CORE_DATAPATH__abc_16259_n3913_1) );
  INVX1 INVX1_173 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_27_), .Y(AES_CORE_DATAPATH__abc_16259_n3915) );
  INVX1 INVX1_174 ( .A(AES_CORE_DATAPATH__abc_16259_n3922), .Y(AES_CORE_DATAPATH__abc_16259_n3923) );
  INVX1 INVX1_175 ( .A(AES_CORE_DATAPATH__abc_16259_n3937_1), .Y(AES_CORE_DATAPATH__abc_16259_n3938) );
  INVX1 INVX1_176 ( .A(AES_CORE_DATAPATH__abc_16259_n3940), .Y(AES_CORE_DATAPATH__abc_16259_n3941) );
  INVX1 INVX1_177 ( .A(AES_CORE_DATAPATH_col_0__28_), .Y(AES_CORE_DATAPATH__abc_16259_n3953_1) );
  INVX1 INVX1_178 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_28_), .Y(AES_CORE_DATAPATH__abc_16259_n3955) );
  INVX1 INVX1_179 ( .A(AES_CORE_DATAPATH__abc_16259_n3962), .Y(AES_CORE_DATAPATH__abc_16259_n3963) );
  INVX1 INVX1_18 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n178), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n179_1) );
  INVX1 INVX1_180 ( .A(AES_CORE_DATAPATH__abc_16259_n3977_1), .Y(AES_CORE_DATAPATH__abc_16259_n3978) );
  INVX1 INVX1_181 ( .A(AES_CORE_DATAPATH__abc_16259_n3980), .Y(AES_CORE_DATAPATH__abc_16259_n3981) );
  INVX1 INVX1_182 ( .A(AES_CORE_DATAPATH_col_0__29_), .Y(AES_CORE_DATAPATH__abc_16259_n3993_1) );
  INVX1 INVX1_183 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_29_), .Y(AES_CORE_DATAPATH__abc_16259_n3995) );
  INVX1 INVX1_184 ( .A(AES_CORE_DATAPATH__abc_16259_n4002), .Y(AES_CORE_DATAPATH__abc_16259_n4003) );
  INVX1 INVX1_185 ( .A(AES_CORE_DATAPATH__abc_16259_n4017_1), .Y(AES_CORE_DATAPATH__abc_16259_n4018) );
  INVX1 INVX1_186 ( .A(AES_CORE_DATAPATH__abc_16259_n4020), .Y(AES_CORE_DATAPATH__abc_16259_n4021) );
  INVX1 INVX1_187 ( .A(AES_CORE_DATAPATH_col_0__30_), .Y(AES_CORE_DATAPATH__abc_16259_n4033_1) );
  INVX1 INVX1_188 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_30_), .Y(AES_CORE_DATAPATH__abc_16259_n4035) );
  INVX1 INVX1_189 ( .A(AES_CORE_DATAPATH__abc_16259_n4042), .Y(AES_CORE_DATAPATH__abc_16259_n4043) );
  INVX1 INVX1_19 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n183_1), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n184_1) );
  INVX1 INVX1_190 ( .A(AES_CORE_DATAPATH__abc_16259_n4057_1), .Y(AES_CORE_DATAPATH__abc_16259_n4058) );
  INVX1 INVX1_191 ( .A(AES_CORE_DATAPATH__abc_16259_n4060), .Y(AES_CORE_DATAPATH__abc_16259_n4061) );
  INVX1 INVX1_192 ( .A(AES_CORE_DATAPATH_col_0__31_), .Y(AES_CORE_DATAPATH__abc_16259_n4073_1) );
  INVX1 INVX1_193 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_31_), .Y(AES_CORE_DATAPATH__abc_16259_n4075) );
  INVX1 INVX1_194 ( .A(AES_CORE_DATAPATH__abc_16259_n4082), .Y(AES_CORE_DATAPATH__abc_16259_n4083) );
  INVX1 INVX1_195 ( .A(AES_CORE_DATAPATH__abc_16259_n4097_1), .Y(AES_CORE_DATAPATH__abc_16259_n4098) );
  INVX1 INVX1_196 ( .A(AES_CORE_DATAPATH__abc_16259_n4100), .Y(AES_CORE_DATAPATH__abc_16259_n4101) );
  INVX1 INVX1_197 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_1_2_), .Y(AES_CORE_DATAPATH__abc_16259_n4210) );
  INVX1 INVX1_198 ( .A(_auto_iopadmap_cc_313_execute_26949_0_), .Y(AES_CORE_DATAPATH__abc_16259_n4212) );
  INVX1 INVX1_199 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_1_), .Y(AES_CORE_DATAPATH__abc_16259_n4218) );
  INVX1 INVX1_2 ( .A(\addr[0] ), .Y(_abc_15830_n12_1) );
  INVX1 INVX1_20 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n195), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n196) );
  INVX1 INVX1_200 ( .A(_auto_iopadmap_cc_313_execute_26949_1_), .Y(AES_CORE_DATAPATH__abc_16259_n4220) );
  INVX1 INVX1_201 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_2_), .Y(AES_CORE_DATAPATH__abc_16259_n4226) );
  INVX1 INVX1_202 ( .A(_auto_iopadmap_cc_313_execute_26949_2_), .Y(AES_CORE_DATAPATH__abc_16259_n4228) );
  INVX1 INVX1_203 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_3_), .Y(AES_CORE_DATAPATH__abc_16259_n4234) );
  INVX1 INVX1_204 ( .A(_auto_iopadmap_cc_313_execute_26949_3_), .Y(AES_CORE_DATAPATH__abc_16259_n4236) );
  INVX1 INVX1_205 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_4_), .Y(AES_CORE_DATAPATH__abc_16259_n4242) );
  INVX1 INVX1_206 ( .A(_auto_iopadmap_cc_313_execute_26949_4_), .Y(AES_CORE_DATAPATH__abc_16259_n4244) );
  INVX1 INVX1_207 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_5_), .Y(AES_CORE_DATAPATH__abc_16259_n4250) );
  INVX1 INVX1_208 ( .A(_auto_iopadmap_cc_313_execute_26949_5_), .Y(AES_CORE_DATAPATH__abc_16259_n4252) );
  INVX1 INVX1_209 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_6_), .Y(AES_CORE_DATAPATH__abc_16259_n4258) );
  INVX1 INVX1_21 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n216), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n217) );
  INVX1 INVX1_210 ( .A(_auto_iopadmap_cc_313_execute_26949_6_), .Y(AES_CORE_DATAPATH__abc_16259_n4260) );
  INVX1 INVX1_211 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_7_), .Y(AES_CORE_DATAPATH__abc_16259_n4266) );
  INVX1 INVX1_212 ( .A(_auto_iopadmap_cc_313_execute_26949_7_), .Y(AES_CORE_DATAPATH__abc_16259_n4268) );
  INVX1 INVX1_213 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_1_2_), .Y(AES_CORE_DATAPATH__abc_16259_n4274) );
  INVX1 INVX1_214 ( .A(_auto_iopadmap_cc_313_execute_26949_8_), .Y(AES_CORE_DATAPATH__abc_16259_n4276) );
  INVX1 INVX1_215 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_1_), .Y(AES_CORE_DATAPATH__abc_16259_n4282) );
  INVX1 INVX1_216 ( .A(_auto_iopadmap_cc_313_execute_26949_9_), .Y(AES_CORE_DATAPATH__abc_16259_n4284) );
  INVX1 INVX1_217 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_2_), .Y(AES_CORE_DATAPATH__abc_16259_n4290) );
  INVX1 INVX1_218 ( .A(_auto_iopadmap_cc_313_execute_26949_10_), .Y(AES_CORE_DATAPATH__abc_16259_n4292) );
  INVX1 INVX1_219 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_3_), .Y(AES_CORE_DATAPATH__abc_16259_n4298) );
  INVX1 INVX1_22 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n137), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n226) );
  INVX1 INVX1_220 ( .A(_auto_iopadmap_cc_313_execute_26949_11_), .Y(AES_CORE_DATAPATH__abc_16259_n4300) );
  INVX1 INVX1_221 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_4_), .Y(AES_CORE_DATAPATH__abc_16259_n4306) );
  INVX1 INVX1_222 ( .A(_auto_iopadmap_cc_313_execute_26949_12_), .Y(AES_CORE_DATAPATH__abc_16259_n4308) );
  INVX1 INVX1_223 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_5_), .Y(AES_CORE_DATAPATH__abc_16259_n4314) );
  INVX1 INVX1_224 ( .A(_auto_iopadmap_cc_313_execute_26949_13_), .Y(AES_CORE_DATAPATH__abc_16259_n4315) );
  INVX1 INVX1_225 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_6_), .Y(AES_CORE_DATAPATH__abc_16259_n4322) );
  INVX1 INVX1_226 ( .A(_auto_iopadmap_cc_313_execute_26949_14_), .Y(AES_CORE_DATAPATH__abc_16259_n4324) );
  INVX1 INVX1_227 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_7_), .Y(AES_CORE_DATAPATH__abc_16259_n4330) );
  INVX1 INVX1_228 ( .A(_auto_iopadmap_cc_313_execute_26949_15_), .Y(AES_CORE_DATAPATH__abc_16259_n4332) );
  INVX1 INVX1_229 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_1_2_), .Y(AES_CORE_DATAPATH__abc_16259_n4338) );
  INVX1 INVX1_23 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n140), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n227) );
  INVX1 INVX1_230 ( .A(_auto_iopadmap_cc_313_execute_26949_16_), .Y(AES_CORE_DATAPATH__abc_16259_n4340) );
  INVX1 INVX1_231 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_1_), .Y(AES_CORE_DATAPATH__abc_16259_n4346) );
  INVX1 INVX1_232 ( .A(_auto_iopadmap_cc_313_execute_26949_17_), .Y(AES_CORE_DATAPATH__abc_16259_n4348) );
  INVX1 INVX1_233 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_2_), .Y(AES_CORE_DATAPATH__abc_16259_n4354) );
  INVX1 INVX1_234 ( .A(_auto_iopadmap_cc_313_execute_26949_18_), .Y(AES_CORE_DATAPATH__abc_16259_n4356) );
  INVX1 INVX1_235 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_3_), .Y(AES_CORE_DATAPATH__abc_16259_n4362) );
  INVX1 INVX1_236 ( .A(_auto_iopadmap_cc_313_execute_26949_19_), .Y(AES_CORE_DATAPATH__abc_16259_n4364) );
  INVX1 INVX1_237 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_4_), .Y(AES_CORE_DATAPATH__abc_16259_n4370) );
  INVX1 INVX1_238 ( .A(_auto_iopadmap_cc_313_execute_26949_20_), .Y(AES_CORE_DATAPATH__abc_16259_n4372) );
  INVX1 INVX1_239 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_5_), .Y(AES_CORE_DATAPATH__abc_16259_n4378) );
  INVX1 INVX1_24 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n188), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n229) );
  INVX1 INVX1_240 ( .A(_auto_iopadmap_cc_313_execute_26949_21_), .Y(AES_CORE_DATAPATH__abc_16259_n4380) );
  INVX1 INVX1_241 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_6_), .Y(AES_CORE_DATAPATH__abc_16259_n4386) );
  INVX1 INVX1_242 ( .A(_auto_iopadmap_cc_313_execute_26949_22_), .Y(AES_CORE_DATAPATH__abc_16259_n4388) );
  INVX1 INVX1_243 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_7_), .Y(AES_CORE_DATAPATH__abc_16259_n4394) );
  INVX1 INVX1_244 ( .A(_auto_iopadmap_cc_313_execute_26949_23_), .Y(AES_CORE_DATAPATH__abc_16259_n4396) );
  INVX1 INVX1_245 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_1_2_), .Y(AES_CORE_DATAPATH__abc_16259_n4402) );
  INVX1 INVX1_246 ( .A(_auto_iopadmap_cc_313_execute_26949_24_), .Y(AES_CORE_DATAPATH__abc_16259_n4404) );
  INVX1 INVX1_247 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_1_), .Y(AES_CORE_DATAPATH__abc_16259_n4410) );
  INVX1 INVX1_248 ( .A(_auto_iopadmap_cc_313_execute_26949_25_), .Y(AES_CORE_DATAPATH__abc_16259_n4412) );
  INVX1 INVX1_249 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_2_), .Y(AES_CORE_DATAPATH__abc_16259_n4418) );
  INVX1 INVX1_25 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n206_1), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n230) );
  INVX1 INVX1_250 ( .A(_auto_iopadmap_cc_313_execute_26949_26_), .Y(AES_CORE_DATAPATH__abc_16259_n4419) );
  INVX1 INVX1_251 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_3_), .Y(AES_CORE_DATAPATH__abc_16259_n4426) );
  INVX1 INVX1_252 ( .A(_auto_iopadmap_cc_313_execute_26949_27_), .Y(AES_CORE_DATAPATH__abc_16259_n4428) );
  INVX1 INVX1_253 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_4_), .Y(AES_CORE_DATAPATH__abc_16259_n4434) );
  INVX1 INVX1_254 ( .A(_auto_iopadmap_cc_313_execute_26949_28_), .Y(AES_CORE_DATAPATH__abc_16259_n4436) );
  INVX1 INVX1_255 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_5_), .Y(AES_CORE_DATAPATH__abc_16259_n4442) );
  INVX1 INVX1_256 ( .A(_auto_iopadmap_cc_313_execute_26949_29_), .Y(AES_CORE_DATAPATH__abc_16259_n4444_1) );
  INVX1 INVX1_257 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_6_), .Y(AES_CORE_DATAPATH__abc_16259_n4450_1) );
  INVX1 INVX1_258 ( .A(_auto_iopadmap_cc_313_execute_26949_30_), .Y(AES_CORE_DATAPATH__abc_16259_n4452_1) );
  INVX1 INVX1_259 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_7_), .Y(AES_CORE_DATAPATH__abc_16259_n4458_1) );
  INVX1 INVX1_26 ( .A(AES_CORE_DATAPATH__abc_16259_n2462_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n2463_1) );
  INVX1 INVX1_260 ( .A(_auto_iopadmap_cc_313_execute_26949_31_), .Y(AES_CORE_DATAPATH__abc_16259_n4460_1) );
  INVX1 INVX1_261 ( .A(AES_CORE_DATAPATH__abc_16259_n4466_1), .Y(AES_CORE_DATAPATH__abc_16259_n4467_1) );
  INVX1 INVX1_262 ( .A(start), .Y(AES_CORE_DATAPATH__abc_16259_n4469_1) );
  INVX1 INVX1_263 ( .A(AES_CORE_DATAPATH__abc_16259_n4471_1), .Y(AES_CORE_DATAPATH__abc_16259_n4472_1) );
  INVX1 INVX1_264 ( .A(AES_CORE_DATAPATH__abc_16259_n4865_1), .Y(AES_CORE_DATAPATH__abc_16259_n4866_1) );
  INVX1 INVX1_265 ( .A(AES_CORE_DATAPATH__abc_16259_n4869_1), .Y(AES_CORE_DATAPATH__abc_16259_n4870_1) );
  INVX1 INVX1_266 ( .A(AES_CORE_DATAPATH__abc_16259_n5258_1), .Y(AES_CORE_DATAPATH__abc_16259_n5259_1) );
  INVX1 INVX1_267 ( .A(AES_CORE_DATAPATH__abc_16259_n5262_1), .Y(AES_CORE_DATAPATH__abc_16259_n5263_1) );
  INVX1 INVX1_268 ( .A(AES_CORE_DATAPATH__abc_16259_n5651), .Y(AES_CORE_DATAPATH__abc_16259_n5652) );
  INVX1 INVX1_269 ( .A(AES_CORE_DATAPATH__abc_16259_n5655), .Y(AES_CORE_DATAPATH__abc_16259_n5656) );
  INVX1 INVX1_27 ( .A(AES_CORE_DATAPATH_col_0__0_), .Y(AES_CORE_DATAPATH__abc_16259_n2770) );
  INVX1 INVX1_270 ( .A(AES_CORE_DATAPATH__abc_16259_n6048), .Y(AES_CORE_DATAPATH__abc_16259_n6049) );
  INVX1 INVX1_271 ( .A(AES_CORE_DATAPATH__abc_16259_n6052), .Y(AES_CORE_DATAPATH__abc_16259_n6055) );
  INVX1 INVX1_272 ( .A(AES_CORE_DATAPATH__abc_16259_n2801_1), .Y(AES_CORE_DATAPATH__abc_16259_n6078) );
  INVX1 INVX1_273 ( .A(AES_CORE_DATAPATH__abc_16259_n2865), .Y(AES_CORE_DATAPATH__abc_16259_n6079) );
  INVX1 INVX1_274 ( .A(AES_CORE_DATAPATH__abc_16259_n6061), .Y(AES_CORE_DATAPATH__abc_16259_n6084) );
  INVX1 INVX1_275 ( .A(AES_CORE_DATAPATH__abc_16259_n6076), .Y(AES_CORE_DATAPATH__abc_16259_n6086) );
  INVX1 INVX1_276 ( .A(AES_CORE_DATAPATH__abc_16259_n2902), .Y(AES_CORE_DATAPATH__abc_16259_n6132) );
  INVX1 INVX1_277 ( .A(AES_CORE_DATAPATH__abc_16259_n2908), .Y(AES_CORE_DATAPATH__abc_16259_n6135) );
  INVX1 INVX1_278 ( .A(AES_CORE_DATAPATH__abc_16259_n6117), .Y(AES_CORE_DATAPATH__abc_16259_n6138) );
  INVX1 INVX1_279 ( .A(AES_CORE_DATAPATH__abc_16259_n6130), .Y(AES_CORE_DATAPATH__abc_16259_n6140) );
  INVX1 INVX1_28 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_0_), .Y(AES_CORE_DATAPATH__abc_16259_n2776) );
  INVX1 INVX1_280 ( .A(AES_CORE_DATAPATH__abc_16259_n2942), .Y(AES_CORE_DATAPATH__abc_16259_n6181) );
  INVX1 INVX1_281 ( .A(AES_CORE_DATAPATH__abc_16259_n2948), .Y(AES_CORE_DATAPATH__abc_16259_n6184) );
  INVX1 INVX1_282 ( .A(AES_CORE_DATAPATH__abc_16259_n6166), .Y(AES_CORE_DATAPATH__abc_16259_n6187) );
  INVX1 INVX1_283 ( .A(AES_CORE_DATAPATH__abc_16259_n6179), .Y(AES_CORE_DATAPATH__abc_16259_n6189) );
  INVX1 INVX1_284 ( .A(AES_CORE_DATAPATH__abc_16259_n2982_1), .Y(AES_CORE_DATAPATH__abc_16259_n6230) );
  INVX1 INVX1_285 ( .A(AES_CORE_DATAPATH__abc_16259_n2988), .Y(AES_CORE_DATAPATH__abc_16259_n6233) );
  INVX1 INVX1_286 ( .A(AES_CORE_DATAPATH__abc_16259_n6215), .Y(AES_CORE_DATAPATH__abc_16259_n6236) );
  INVX1 INVX1_287 ( .A(AES_CORE_DATAPATH__abc_16259_n6228), .Y(AES_CORE_DATAPATH__abc_16259_n6238) );
  INVX1 INVX1_288 ( .A(AES_CORE_DATAPATH__abc_16259_n3022), .Y(AES_CORE_DATAPATH__abc_16259_n6279) );
  INVX1 INVX1_289 ( .A(AES_CORE_DATAPATH__abc_16259_n3028), .Y(AES_CORE_DATAPATH__abc_16259_n6282) );
  INVX1 INVX1_29 ( .A(AES_CORE_CONTROL_UNIT_sbox_sel_2_), .Y(AES_CORE_DATAPATH__abc_16259_n2777_1) );
  INVX1 INVX1_290 ( .A(AES_CORE_DATAPATH__abc_16259_n6264), .Y(AES_CORE_DATAPATH__abc_16259_n6285) );
  INVX1 INVX1_291 ( .A(AES_CORE_DATAPATH__abc_16259_n6277), .Y(AES_CORE_DATAPATH__abc_16259_n6287) );
  INVX1 INVX1_292 ( .A(AES_CORE_DATAPATH__abc_16259_n3062_1), .Y(AES_CORE_DATAPATH__abc_16259_n6328) );
  INVX1 INVX1_293 ( .A(AES_CORE_DATAPATH__abc_16259_n3068), .Y(AES_CORE_DATAPATH__abc_16259_n6331) );
  INVX1 INVX1_294 ( .A(AES_CORE_DATAPATH__abc_16259_n6313), .Y(AES_CORE_DATAPATH__abc_16259_n6334) );
  INVX1 INVX1_295 ( .A(AES_CORE_DATAPATH__abc_16259_n6326), .Y(AES_CORE_DATAPATH__abc_16259_n6336) );
  INVX1 INVX1_296 ( .A(AES_CORE_DATAPATH__abc_16259_n3102), .Y(AES_CORE_DATAPATH__abc_16259_n6377) );
  INVX1 INVX1_297 ( .A(AES_CORE_DATAPATH__abc_16259_n3108), .Y(AES_CORE_DATAPATH__abc_16259_n6380) );
  INVX1 INVX1_298 ( .A(AES_CORE_DATAPATH__abc_16259_n6362), .Y(AES_CORE_DATAPATH__abc_16259_n6383) );
  INVX1 INVX1_299 ( .A(AES_CORE_DATAPATH__abc_16259_n6375), .Y(AES_CORE_DATAPATH__abc_16259_n6385) );
  INVX1 INVX1_3 ( .A(\aes_mode[0] ), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n73) );
  INVX1 INVX1_30 ( .A(AES_CORE_DATAPATH__abc_16259_n2772_1), .Y(AES_CORE_DATAPATH__abc_16259_n2784) );
  INVX1 INVX1_300 ( .A(AES_CORE_DATAPATH__abc_16259_n3142), .Y(AES_CORE_DATAPATH__abc_16259_n6426) );
  INVX1 INVX1_301 ( .A(AES_CORE_DATAPATH__abc_16259_n3148_1), .Y(AES_CORE_DATAPATH__abc_16259_n6429) );
  INVX1 INVX1_302 ( .A(AES_CORE_DATAPATH__abc_16259_n6411), .Y(AES_CORE_DATAPATH__abc_16259_n6432) );
  INVX1 INVX1_303 ( .A(AES_CORE_DATAPATH__abc_16259_n6424), .Y(AES_CORE_DATAPATH__abc_16259_n6434) );
  INVX1 INVX1_304 ( .A(AES_CORE_DATAPATH__abc_16259_n3182), .Y(AES_CORE_DATAPATH__abc_16259_n6475) );
  INVX1 INVX1_305 ( .A(AES_CORE_DATAPATH__abc_16259_n3188), .Y(AES_CORE_DATAPATH__abc_16259_n6478) );
  INVX1 INVX1_306 ( .A(AES_CORE_DATAPATH__abc_16259_n6460), .Y(AES_CORE_DATAPATH__abc_16259_n6481) );
  INVX1 INVX1_307 ( .A(AES_CORE_DATAPATH__abc_16259_n6473), .Y(AES_CORE_DATAPATH__abc_16259_n6483) );
  INVX1 INVX1_308 ( .A(AES_CORE_DATAPATH__abc_16259_n3222), .Y(AES_CORE_DATAPATH__abc_16259_n6524) );
  INVX1 INVX1_309 ( .A(AES_CORE_DATAPATH__abc_16259_n3228_1), .Y(AES_CORE_DATAPATH__abc_16259_n6527) );
  INVX1 INVX1_31 ( .A(AES_CORE_DATAPATH__abc_16259_n2771_1), .Y(AES_CORE_DATAPATH__abc_16259_n2788) );
  INVX1 INVX1_310 ( .A(AES_CORE_DATAPATH__abc_16259_n6509), .Y(AES_CORE_DATAPATH__abc_16259_n6530) );
  INVX1 INVX1_311 ( .A(AES_CORE_DATAPATH__abc_16259_n6522), .Y(AES_CORE_DATAPATH__abc_16259_n6532) );
  INVX1 INVX1_312 ( .A(AES_CORE_DATAPATH__abc_16259_n3262), .Y(AES_CORE_DATAPATH__abc_16259_n6557) );
  INVX1 INVX1_313 ( .A(AES_CORE_DATAPATH__abc_16259_n3268_1), .Y(AES_CORE_DATAPATH__abc_16259_n6560) );
  INVX1 INVX1_314 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_10_), .Y(AES_CORE_DATAPATH__abc_16259_n6563) );
  INVX1 INVX1_315 ( .A(AES_CORE_DATAPATH__abc_16259_n6564), .Y(AES_CORE_DATAPATH__abc_16259_n6580) );
  INVX1 INVX1_316 ( .A(AES_CORE_DATAPATH__abc_16259_n6577), .Y(AES_CORE_DATAPATH__abc_16259_n6582) );
  INVX1 INVX1_317 ( .A(_auto_iopadmap_cc_313_execute_26916_10_), .Y(AES_CORE_DATAPATH__abc_16259_n6587) );
  INVX1 INVX1_318 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_42_), .Y(AES_CORE_DATAPATH__abc_16259_n6604) );
  INVX1 INVX1_319 ( .A(AES_CORE_DATAPATH__abc_16259_n6606), .Y(AES_CORE_DATAPATH__abc_16259_n6607) );
  INVX1 INVX1_32 ( .A(AES_CORE_DATAPATH__abc_16259_n2792), .Y(AES_CORE_DATAPATH__abc_16259_n2793_1) );
  INVX1 INVX1_320 ( .A(AES_CORE_DATAPATH__abc_16259_n6611), .Y(AES_CORE_DATAPATH__abc_16259_n6612) );
  INVX1 INVX1_321 ( .A(AES_CORE_DATAPATH__abc_16259_n3302), .Y(AES_CORE_DATAPATH__abc_16259_n6615) );
  INVX1 INVX1_322 ( .A(AES_CORE_DATAPATH__abc_16259_n3308), .Y(AES_CORE_DATAPATH__abc_16259_n6618) );
  INVX1 INVX1_323 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_11_), .Y(AES_CORE_DATAPATH__abc_16259_n6621) );
  INVX1 INVX1_324 ( .A(AES_CORE_DATAPATH__abc_16259_n6622), .Y(AES_CORE_DATAPATH__abc_16259_n6638) );
  INVX1 INVX1_325 ( .A(AES_CORE_DATAPATH__abc_16259_n6635), .Y(AES_CORE_DATAPATH__abc_16259_n6640) );
  INVX1 INVX1_326 ( .A(_auto_iopadmap_cc_313_execute_26916_11_), .Y(AES_CORE_DATAPATH__abc_16259_n6644) );
  INVX1 INVX1_327 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_43_), .Y(AES_CORE_DATAPATH__abc_16259_n6658) );
  INVX1 INVX1_328 ( .A(AES_CORE_DATAPATH__abc_16259_n6660), .Y(AES_CORE_DATAPATH__abc_16259_n6661) );
  INVX1 INVX1_329 ( .A(AES_CORE_DATAPATH__abc_16259_n6665), .Y(AES_CORE_DATAPATH__abc_16259_n6666) );
  INVX1 INVX1_33 ( .A(AES_CORE_DATAPATH__abc_16259_n2810_1), .Y(AES_CORE_DATAPATH__abc_16259_n2811) );
  INVX1 INVX1_330 ( .A(AES_CORE_DATAPATH__abc_16259_n3342), .Y(AES_CORE_DATAPATH__abc_16259_n6686) );
  INVX1 INVX1_331 ( .A(AES_CORE_DATAPATH__abc_16259_n3348), .Y(AES_CORE_DATAPATH__abc_16259_n6689) );
  INVX1 INVX1_332 ( .A(AES_CORE_DATAPATH__abc_16259_n6671), .Y(AES_CORE_DATAPATH__abc_16259_n6692) );
  INVX1 INVX1_333 ( .A(AES_CORE_DATAPATH__abc_16259_n6684), .Y(AES_CORE_DATAPATH__abc_16259_n6694) );
  INVX1 INVX1_334 ( .A(AES_CORE_DATAPATH__abc_16259_n3382), .Y(AES_CORE_DATAPATH__abc_16259_n6718) );
  INVX1 INVX1_335 ( .A(AES_CORE_DATAPATH__abc_16259_n3388_1), .Y(AES_CORE_DATAPATH__abc_16259_n6721) );
  INVX1 INVX1_336 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_13_), .Y(AES_CORE_DATAPATH__abc_16259_n6724) );
  INVX1 INVX1_337 ( .A(AES_CORE_DATAPATH__abc_16259_n6725), .Y(AES_CORE_DATAPATH__abc_16259_n6741) );
  INVX1 INVX1_338 ( .A(AES_CORE_DATAPATH__abc_16259_n6738), .Y(AES_CORE_DATAPATH__abc_16259_n6743) );
  INVX1 INVX1_339 ( .A(_auto_iopadmap_cc_313_execute_26916_13_), .Y(AES_CORE_DATAPATH__abc_16259_n6747) );
  INVX1 INVX1_34 ( .A(AES_CORE_DATAPATH__abc_16259_n2813), .Y(AES_CORE_DATAPATH__abc_16259_n2814) );
  INVX1 INVX1_340 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_45_), .Y(AES_CORE_DATAPATH__abc_16259_n6761) );
  INVX1 INVX1_341 ( .A(AES_CORE_DATAPATH__abc_16259_n6763), .Y(AES_CORE_DATAPATH__abc_16259_n6764) );
  INVX1 INVX1_342 ( .A(AES_CORE_DATAPATH__abc_16259_n6768), .Y(AES_CORE_DATAPATH__abc_16259_n6769) );
  INVX1 INVX1_343 ( .A(AES_CORE_DATAPATH__abc_16259_n3422), .Y(AES_CORE_DATAPATH__abc_16259_n6789) );
  INVX1 INVX1_344 ( .A(AES_CORE_DATAPATH__abc_16259_n3428), .Y(AES_CORE_DATAPATH__abc_16259_n6792) );
  INVX1 INVX1_345 ( .A(AES_CORE_DATAPATH__abc_16259_n6774), .Y(AES_CORE_DATAPATH__abc_16259_n6795) );
  INVX1 INVX1_346 ( .A(AES_CORE_DATAPATH__abc_16259_n6787), .Y(AES_CORE_DATAPATH__abc_16259_n6797) );
  INVX1 INVX1_347 ( .A(AES_CORE_DATAPATH__abc_16259_n3462_1), .Y(AES_CORE_DATAPATH__abc_16259_n6821) );
  INVX1 INVX1_348 ( .A(AES_CORE_DATAPATH__abc_16259_n3468_1), .Y(AES_CORE_DATAPATH__abc_16259_n6824) );
  INVX1 INVX1_349 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_15_), .Y(AES_CORE_DATAPATH__abc_16259_n6827) );
  INVX1 INVX1_35 ( .A(AES_CORE_DATAPATH_key_out_sel_pp1_0_), .Y(AES_CORE_DATAPATH__abc_16259_n2816) );
  INVX1 INVX1_350 ( .A(AES_CORE_DATAPATH__abc_16259_n6828), .Y(AES_CORE_DATAPATH__abc_16259_n6844) );
  INVX1 INVX1_351 ( .A(AES_CORE_DATAPATH__abc_16259_n6841), .Y(AES_CORE_DATAPATH__abc_16259_n6846) );
  INVX1 INVX1_352 ( .A(_auto_iopadmap_cc_313_execute_26916_15_), .Y(AES_CORE_DATAPATH__abc_16259_n6850) );
  INVX1 INVX1_353 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_47_), .Y(AES_CORE_DATAPATH__abc_16259_n6864) );
  INVX1 INVX1_354 ( .A(AES_CORE_DATAPATH__abc_16259_n6866), .Y(AES_CORE_DATAPATH__abc_16259_n6867) );
  INVX1 INVX1_355 ( .A(AES_CORE_DATAPATH__abc_16259_n6871), .Y(AES_CORE_DATAPATH__abc_16259_n6872) );
  INVX1 INVX1_356 ( .A(AES_CORE_DATAPATH__abc_16259_n3502_1), .Y(AES_CORE_DATAPATH__abc_16259_n6876) );
  INVX1 INVX1_357 ( .A(AES_CORE_DATAPATH__abc_16259_n3508), .Y(AES_CORE_DATAPATH__abc_16259_n6879) );
  INVX1 INVX1_358 ( .A(AES_CORE_DATAPATH__abc_16259_n6882), .Y(AES_CORE_DATAPATH__abc_16259_n6883) );
  INVX1 INVX1_359 ( .A(AES_CORE_DATAPATH__abc_16259_n6896), .Y(AES_CORE_DATAPATH__abc_16259_n6897) );
  INVX1 INVX1_36 ( .A(AES_CORE_DATAPATH_key_out_sel_pp2_0_), .Y(AES_CORE_DATAPATH__abc_16259_n2818) );
  INVX1 INVX1_360 ( .A(AES_CORE_DATAPATH__abc_16259_n3542), .Y(AES_CORE_DATAPATH__abc_16259_n6924) );
  INVX1 INVX1_361 ( .A(AES_CORE_DATAPATH__abc_16259_n3548), .Y(AES_CORE_DATAPATH__abc_16259_n6927) );
  INVX1 INVX1_362 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_17_), .Y(AES_CORE_DATAPATH__abc_16259_n6930) );
  INVX1 INVX1_363 ( .A(AES_CORE_DATAPATH__abc_16259_n6931), .Y(AES_CORE_DATAPATH__abc_16259_n6947) );
  INVX1 INVX1_364 ( .A(AES_CORE_DATAPATH__abc_16259_n6944), .Y(AES_CORE_DATAPATH__abc_16259_n6949) );
  INVX1 INVX1_365 ( .A(_auto_iopadmap_cc_313_execute_26916_17_), .Y(AES_CORE_DATAPATH__abc_16259_n6953) );
  INVX1 INVX1_366 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_17_), .Y(AES_CORE_DATAPATH__abc_16259_n6967) );
  INVX1 INVX1_367 ( .A(AES_CORE_DATAPATH__abc_16259_n6969), .Y(AES_CORE_DATAPATH__abc_16259_n6970) );
  INVX1 INVX1_368 ( .A(AES_CORE_DATAPATH__abc_16259_n6974), .Y(AES_CORE_DATAPATH__abc_16259_n6975) );
  INVX1 INVX1_369 ( .A(AES_CORE_DATAPATH__abc_16259_n3582), .Y(AES_CORE_DATAPATH__abc_16259_n6995) );
  INVX1 INVX1_37 ( .A(AES_CORE_DATAPATH__abc_16259_n2823), .Y(AES_CORE_DATAPATH__abc_16259_n2824_1) );
  INVX1 INVX1_370 ( .A(AES_CORE_DATAPATH__abc_16259_n3588), .Y(AES_CORE_DATAPATH__abc_16259_n6998) );
  INVX1 INVX1_371 ( .A(AES_CORE_DATAPATH__abc_16259_n6980), .Y(AES_CORE_DATAPATH__abc_16259_n7001) );
  INVX1 INVX1_372 ( .A(AES_CORE_DATAPATH__abc_16259_n6993), .Y(AES_CORE_DATAPATH__abc_16259_n7003) );
  INVX1 INVX1_373 ( .A(AES_CORE_DATAPATH__abc_16259_n3622_1), .Y(AES_CORE_DATAPATH__abc_16259_n7044) );
  INVX1 INVX1_374 ( .A(AES_CORE_DATAPATH__abc_16259_n3628), .Y(AES_CORE_DATAPATH__abc_16259_n7047) );
  INVX1 INVX1_375 ( .A(AES_CORE_DATAPATH__abc_16259_n7029), .Y(AES_CORE_DATAPATH__abc_16259_n7050) );
  INVX1 INVX1_376 ( .A(AES_CORE_DATAPATH__abc_16259_n7042), .Y(AES_CORE_DATAPATH__abc_16259_n7052) );
  INVX1 INVX1_377 ( .A(AES_CORE_DATAPATH__abc_16259_n3662), .Y(AES_CORE_DATAPATH__abc_16259_n7093) );
  INVX1 INVX1_378 ( .A(AES_CORE_DATAPATH__abc_16259_n3668), .Y(AES_CORE_DATAPATH__abc_16259_n7096) );
  INVX1 INVX1_379 ( .A(AES_CORE_DATAPATH__abc_16259_n7078), .Y(AES_CORE_DATAPATH__abc_16259_n7099) );
  INVX1 INVX1_38 ( .A(AES_CORE_DATAPATH__abc_16259_n2846), .Y(AES_CORE_DATAPATH__abc_16259_n2847) );
  INVX1 INVX1_380 ( .A(AES_CORE_DATAPATH__abc_16259_n7091), .Y(AES_CORE_DATAPATH__abc_16259_n7101) );
  INVX1 INVX1_381 ( .A(AES_CORE_DATAPATH__abc_16259_n3702_1), .Y(AES_CORE_DATAPATH__abc_16259_n7125) );
  INVX1 INVX1_382 ( .A(AES_CORE_DATAPATH__abc_16259_n3708), .Y(AES_CORE_DATAPATH__abc_16259_n7128) );
  INVX1 INVX1_383 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_21_), .Y(AES_CORE_DATAPATH__abc_16259_n7131) );
  INVX1 INVX1_384 ( .A(AES_CORE_DATAPATH__abc_16259_n7132), .Y(AES_CORE_DATAPATH__abc_16259_n7148) );
  INVX1 INVX1_385 ( .A(AES_CORE_DATAPATH__abc_16259_n7145), .Y(AES_CORE_DATAPATH__abc_16259_n7150) );
  INVX1 INVX1_386 ( .A(_auto_iopadmap_cc_313_execute_26916_21_), .Y(AES_CORE_DATAPATH__abc_16259_n7154) );
  INVX1 INVX1_387 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_21_), .Y(AES_CORE_DATAPATH__abc_16259_n7168) );
  INVX1 INVX1_388 ( .A(AES_CORE_DATAPATH__abc_16259_n7170), .Y(AES_CORE_DATAPATH__abc_16259_n7171) );
  INVX1 INVX1_389 ( .A(AES_CORE_DATAPATH__abc_16259_n7175), .Y(AES_CORE_DATAPATH__abc_16259_n7176) );
  INVX1 INVX1_39 ( .A(AES_CORE_DATAPATH__abc_16259_n2850), .Y(AES_CORE_DATAPATH__abc_16259_n2851_1) );
  INVX1 INVX1_390 ( .A(AES_CORE_DATAPATH__abc_16259_n3742_1), .Y(AES_CORE_DATAPATH__abc_16259_n7196) );
  INVX1 INVX1_391 ( .A(AES_CORE_DATAPATH__abc_16259_n3748), .Y(AES_CORE_DATAPATH__abc_16259_n7199) );
  INVX1 INVX1_392 ( .A(AES_CORE_DATAPATH__abc_16259_n7181), .Y(AES_CORE_DATAPATH__abc_16259_n7202) );
  INVX1 INVX1_393 ( .A(AES_CORE_DATAPATH__abc_16259_n7194), .Y(AES_CORE_DATAPATH__abc_16259_n7204) );
  INVX1 INVX1_394 ( .A(AES_CORE_DATAPATH__abc_16259_n3782_1), .Y(AES_CORE_DATAPATH__abc_16259_n7229) );
  INVX1 INVX1_395 ( .A(AES_CORE_DATAPATH__abc_16259_n3788), .Y(AES_CORE_DATAPATH__abc_16259_n7232) );
  INVX1 INVX1_396 ( .A(AES_CORE_DATAPATH__abc_16259_n7235), .Y(AES_CORE_DATAPATH__abc_16259_n7236) );
  INVX1 INVX1_397 ( .A(AES_CORE_DATAPATH__abc_16259_n7249), .Y(AES_CORE_DATAPATH__abc_16259_n7250) );
  INVX1 INVX1_398 ( .A(AES_CORE_DATAPATH__abc_16259_n3822_1), .Y(AES_CORE_DATAPATH__abc_16259_n7294) );
  INVX1 INVX1_399 ( .A(AES_CORE_DATAPATH__abc_16259_n3828), .Y(AES_CORE_DATAPATH__abc_16259_n7297) );
  INVX1 INVX1_4 ( .A(\op_mode[1] ), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n77) );
  INVX1 INVX1_40 ( .A(AES_CORE_DATAPATH__abc_16259_n2859_1), .Y(AES_CORE_DATAPATH__abc_16259_n2860) );
  INVX1 INVX1_400 ( .A(AES_CORE_DATAPATH__abc_16259_n7279), .Y(AES_CORE_DATAPATH__abc_16259_n7300) );
  INVX1 INVX1_401 ( .A(AES_CORE_DATAPATH__abc_16259_n7292), .Y(AES_CORE_DATAPATH__abc_16259_n7302) );
  INVX1 INVX1_402 ( .A(AES_CORE_DATAPATH__abc_16259_n3862_1), .Y(AES_CORE_DATAPATH__abc_16259_n7343) );
  INVX1 INVX1_403 ( .A(AES_CORE_DATAPATH__abc_16259_n3868), .Y(AES_CORE_DATAPATH__abc_16259_n7346) );
  INVX1 INVX1_404 ( .A(AES_CORE_DATAPATH__abc_16259_n7328), .Y(AES_CORE_DATAPATH__abc_16259_n7349) );
  INVX1 INVX1_405 ( .A(AES_CORE_DATAPATH__abc_16259_n7341), .Y(AES_CORE_DATAPATH__abc_16259_n7351) );
  INVX1 INVX1_406 ( .A(AES_CORE_DATAPATH__abc_16259_n3902_1), .Y(AES_CORE_DATAPATH__abc_16259_n7376) );
  INVX1 INVX1_407 ( .A(AES_CORE_DATAPATH__abc_16259_n3908), .Y(AES_CORE_DATAPATH__abc_16259_n7379) );
  INVX1 INVX1_408 ( .A(AES_CORE_DATAPATH__abc_16259_n7382), .Y(AES_CORE_DATAPATH__abc_16259_n7383) );
  INVX1 INVX1_409 ( .A(AES_CORE_DATAPATH__abc_16259_n7396), .Y(AES_CORE_DATAPATH__abc_16259_n7397) );
  INVX1 INVX1_41 ( .A(AES_CORE_DATAPATH__abc_16259_n2862_1), .Y(AES_CORE_DATAPATH__abc_16259_n2863) );
  INVX1 INVX1_410 ( .A(AES_CORE_DATAPATH__abc_16259_n3942_1), .Y(AES_CORE_DATAPATH__abc_16259_n7441) );
  INVX1 INVX1_411 ( .A(AES_CORE_DATAPATH__abc_16259_n3948), .Y(AES_CORE_DATAPATH__abc_16259_n7444) );
  INVX1 INVX1_412 ( .A(AES_CORE_DATAPATH__abc_16259_n7426), .Y(AES_CORE_DATAPATH__abc_16259_n7447) );
  INVX1 INVX1_413 ( .A(AES_CORE_DATAPATH__abc_16259_n7439), .Y(AES_CORE_DATAPATH__abc_16259_n7449) );
  INVX1 INVX1_414 ( .A(AES_CORE_DATAPATH__abc_16259_n3982_1), .Y(AES_CORE_DATAPATH__abc_16259_n7474) );
  INVX1 INVX1_415 ( .A(AES_CORE_DATAPATH__abc_16259_n3988), .Y(AES_CORE_DATAPATH__abc_16259_n7477) );
  INVX1 INVX1_416 ( .A(AES_CORE_DATAPATH__abc_16259_n7480), .Y(AES_CORE_DATAPATH__abc_16259_n7481) );
  INVX1 INVX1_417 ( .A(AES_CORE_DATAPATH__abc_16259_n7494), .Y(AES_CORE_DATAPATH__abc_16259_n7495) );
  INVX1 INVX1_418 ( .A(AES_CORE_DATAPATH__abc_16259_n4022_1), .Y(AES_CORE_DATAPATH__abc_16259_n7539) );
  INVX1 INVX1_419 ( .A(AES_CORE_DATAPATH__abc_16259_n4028), .Y(AES_CORE_DATAPATH__abc_16259_n7542) );
  INVX1 INVX1_42 ( .A(AES_CORE_DATAPATH_col_0__1_), .Y(AES_CORE_DATAPATH__abc_16259_n2872) );
  INVX1 INVX1_420 ( .A(AES_CORE_DATAPATH__abc_16259_n7524), .Y(AES_CORE_DATAPATH__abc_16259_n7545) );
  INVX1 INVX1_421 ( .A(AES_CORE_DATAPATH__abc_16259_n7537), .Y(AES_CORE_DATAPATH__abc_16259_n7547) );
  INVX1 INVX1_422 ( .A(AES_CORE_DATAPATH__abc_16259_n4062_1), .Y(AES_CORE_DATAPATH__abc_16259_n7588) );
  INVX1 INVX1_423 ( .A(AES_CORE_DATAPATH__abc_16259_n4068), .Y(AES_CORE_DATAPATH__abc_16259_n7591) );
  INVX1 INVX1_424 ( .A(AES_CORE_DATAPATH__abc_16259_n7573), .Y(AES_CORE_DATAPATH__abc_16259_n7594) );
  INVX1 INVX1_425 ( .A(AES_CORE_DATAPATH__abc_16259_n7586), .Y(AES_CORE_DATAPATH__abc_16259_n7596) );
  INVX1 INVX1_426 ( .A(AES_CORE_DATAPATH__abc_16259_n4102_1), .Y(AES_CORE_DATAPATH__abc_16259_n7637) );
  INVX1 INVX1_427 ( .A(AES_CORE_DATAPATH__abc_16259_n4108), .Y(AES_CORE_DATAPATH__abc_16259_n7640) );
  INVX1 INVX1_428 ( .A(AES_CORE_DATAPATH__abc_16259_n7622), .Y(AES_CORE_DATAPATH__abc_16259_n7643) );
  INVX1 INVX1_429 ( .A(AES_CORE_DATAPATH__abc_16259_n7635), .Y(AES_CORE_DATAPATH__abc_16259_n7645) );
  INVX1 INVX1_43 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_1_), .Y(AES_CORE_DATAPATH__abc_16259_n2874) );
  INVX1 INVX1_430 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_10_), .Y(AES_CORE_DATAPATH__abc_16259_n7751) );
  INVX1 INVX1_431 ( .A(AES_CORE_DATAPATH__abc_16259_n7753), .Y(AES_CORE_DATAPATH__abc_16259_n7754) );
  INVX1 INVX1_432 ( .A(AES_CORE_DATAPATH__abc_16259_n7758), .Y(AES_CORE_DATAPATH__abc_16259_n7759) );
  INVX1 INVX1_433 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_11_), .Y(AES_CORE_DATAPATH__abc_16259_n7761) );
  INVX1 INVX1_434 ( .A(AES_CORE_DATAPATH__abc_16259_n7763), .Y(AES_CORE_DATAPATH__abc_16259_n7764) );
  INVX1 INVX1_435 ( .A(AES_CORE_DATAPATH__abc_16259_n7768), .Y(AES_CORE_DATAPATH__abc_16259_n7769) );
  INVX1 INVX1_436 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_13_), .Y(AES_CORE_DATAPATH__abc_16259_n7780) );
  INVX1 INVX1_437 ( .A(AES_CORE_DATAPATH__abc_16259_n7782), .Y(AES_CORE_DATAPATH__abc_16259_n7783) );
  INVX1 INVX1_438 ( .A(AES_CORE_DATAPATH__abc_16259_n7787), .Y(AES_CORE_DATAPATH__abc_16259_n7788) );
  INVX1 INVX1_439 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_15_), .Y(AES_CORE_DATAPATH__abc_16259_n7799) );
  INVX1 INVX1_44 ( .A(AES_CORE_DATAPATH__abc_16259_n2881), .Y(AES_CORE_DATAPATH__abc_16259_n2882_1) );
  INVX1 INVX1_440 ( .A(AES_CORE_DATAPATH__abc_16259_n7801), .Y(AES_CORE_DATAPATH__abc_16259_n7802) );
  INVX1 INVX1_441 ( .A(AES_CORE_DATAPATH__abc_16259_n7806), .Y(AES_CORE_DATAPATH__abc_16259_n7807) );
  INVX1 INVX1_442 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_113_), .Y(AES_CORE_DATAPATH__abc_16259_n7818) );
  INVX1 INVX1_443 ( .A(AES_CORE_DATAPATH__abc_16259_n7820), .Y(AES_CORE_DATAPATH__abc_16259_n7821) );
  INVX1 INVX1_444 ( .A(AES_CORE_DATAPATH__abc_16259_n7825), .Y(AES_CORE_DATAPATH__abc_16259_n7826) );
  INVX1 INVX1_445 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_117_), .Y(AES_CORE_DATAPATH__abc_16259_n7853) );
  INVX1 INVX1_446 ( .A(AES_CORE_DATAPATH__abc_16259_n7855), .Y(AES_CORE_DATAPATH__abc_16259_n7856) );
  INVX1 INVX1_447 ( .A(AES_CORE_DATAPATH__abc_16259_n7860), .Y(AES_CORE_DATAPATH__abc_16259_n7861) );
  INVX1 INVX1_448 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_106_), .Y(AES_CORE_DATAPATH__abc_16259_n8025) );
  INVX1 INVX1_449 ( .A(AES_CORE_DATAPATH__abc_16259_n8027), .Y(AES_CORE_DATAPATH__abc_16259_n8028) );
  INVX1 INVX1_45 ( .A(AES_CORE_DATAPATH__abc_16259_n2897_1), .Y(AES_CORE_DATAPATH__abc_16259_n2898) );
  INVX1 INVX1_450 ( .A(AES_CORE_DATAPATH__abc_16259_n8032), .Y(AES_CORE_DATAPATH__abc_16259_n8033) );
  INVX1 INVX1_451 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_107_), .Y(AES_CORE_DATAPATH__abc_16259_n8037) );
  INVX1 INVX1_452 ( .A(AES_CORE_DATAPATH__abc_16259_n8039), .Y(AES_CORE_DATAPATH__abc_16259_n8040) );
  INVX1 INVX1_453 ( .A(AES_CORE_DATAPATH__abc_16259_n8044), .Y(AES_CORE_DATAPATH__abc_16259_n8045) );
  INVX1 INVX1_454 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_109_), .Y(AES_CORE_DATAPATH__abc_16259_n8055) );
  INVX1 INVX1_455 ( .A(AES_CORE_DATAPATH__abc_16259_n8057), .Y(AES_CORE_DATAPATH__abc_16259_n8058) );
  INVX1 INVX1_456 ( .A(AES_CORE_DATAPATH__abc_16259_n8062), .Y(AES_CORE_DATAPATH__abc_16259_n8063) );
  INVX1 INVX1_457 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_111_), .Y(AES_CORE_DATAPATH__abc_16259_n8074) );
  INVX1 INVX1_458 ( .A(AES_CORE_DATAPATH__abc_16259_n8076), .Y(AES_CORE_DATAPATH__abc_16259_n8077) );
  INVX1 INVX1_459 ( .A(AES_CORE_DATAPATH__abc_16259_n8081), .Y(AES_CORE_DATAPATH__abc_16259_n8082) );
  INVX1 INVX1_46 ( .A(AES_CORE_DATAPATH__abc_16259_n2900), .Y(AES_CORE_DATAPATH__abc_16259_n2901) );
  INVX1 INVX1_460 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_81_), .Y(AES_CORE_DATAPATH__abc_16259_n8093) );
  INVX1 INVX1_461 ( .A(AES_CORE_DATAPATH__abc_16259_n8095), .Y(AES_CORE_DATAPATH__abc_16259_n8096) );
  INVX1 INVX1_462 ( .A(AES_CORE_DATAPATH__abc_16259_n8100), .Y(AES_CORE_DATAPATH__abc_16259_n8101) );
  INVX1 INVX1_463 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_85_), .Y(AES_CORE_DATAPATH__abc_16259_n8128) );
  INVX1 INVX1_464 ( .A(AES_CORE_DATAPATH__abc_16259_n8130), .Y(AES_CORE_DATAPATH__abc_16259_n8131) );
  INVX1 INVX1_465 ( .A(AES_CORE_DATAPATH__abc_16259_n8135), .Y(AES_CORE_DATAPATH__abc_16259_n8136) );
  INVX1 INVX1_466 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_74_), .Y(AES_CORE_DATAPATH__abc_16259_n8300) );
  INVX1 INVX1_467 ( .A(AES_CORE_DATAPATH__abc_16259_n8302), .Y(AES_CORE_DATAPATH__abc_16259_n8303) );
  INVX1 INVX1_468 ( .A(AES_CORE_DATAPATH__abc_16259_n8307), .Y(AES_CORE_DATAPATH__abc_16259_n8308) );
  INVX1 INVX1_469 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_75_), .Y(AES_CORE_DATAPATH__abc_16259_n8311) );
  INVX1 INVX1_47 ( .A(AES_CORE_DATAPATH_col_0__2_), .Y(AES_CORE_DATAPATH__abc_16259_n2913) );
  INVX1 INVX1_470 ( .A(AES_CORE_DATAPATH__abc_16259_n8313), .Y(AES_CORE_DATAPATH__abc_16259_n8314) );
  INVX1 INVX1_471 ( .A(AES_CORE_DATAPATH__abc_16259_n8318), .Y(AES_CORE_DATAPATH__abc_16259_n8319) );
  INVX1 INVX1_472 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_77_), .Y(AES_CORE_DATAPATH__abc_16259_n8330) );
  INVX1 INVX1_473 ( .A(AES_CORE_DATAPATH__abc_16259_n8332), .Y(AES_CORE_DATAPATH__abc_16259_n8333) );
  INVX1 INVX1_474 ( .A(AES_CORE_DATAPATH__abc_16259_n8337), .Y(AES_CORE_DATAPATH__abc_16259_n8338) );
  INVX1 INVX1_475 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_79_), .Y(AES_CORE_DATAPATH__abc_16259_n8349) );
  INVX1 INVX1_476 ( .A(AES_CORE_DATAPATH__abc_16259_n8351), .Y(AES_CORE_DATAPATH__abc_16259_n8352) );
  INVX1 INVX1_477 ( .A(AES_CORE_DATAPATH__abc_16259_n8356), .Y(AES_CORE_DATAPATH__abc_16259_n8357) );
  INVX1 INVX1_478 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_49_), .Y(AES_CORE_DATAPATH__abc_16259_n8368) );
  INVX1 INVX1_479 ( .A(AES_CORE_DATAPATH__abc_16259_n8370), .Y(AES_CORE_DATAPATH__abc_16259_n8371) );
  INVX1 INVX1_48 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_2_), .Y(AES_CORE_DATAPATH__abc_16259_n2915) );
  INVX1 INVX1_480 ( .A(AES_CORE_DATAPATH__abc_16259_n8375), .Y(AES_CORE_DATAPATH__abc_16259_n8376) );
  INVX1 INVX1_481 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_53_), .Y(AES_CORE_DATAPATH__abc_16259_n8403) );
  INVX1 INVX1_482 ( .A(AES_CORE_DATAPATH__abc_16259_n8405), .Y(AES_CORE_DATAPATH__abc_16259_n8406) );
  INVX1 INVX1_483 ( .A(AES_CORE_DATAPATH__abc_16259_n8410), .Y(AES_CORE_DATAPATH__abc_16259_n8411) );
  INVX1 INVX1_484 ( .A(AES_CORE_DATAPATH__abc_16259_n8531), .Y(AES_CORE_DATAPATH__abc_16259_n8532) );
  INVX1 INVX1_485 ( .A(AES_CORE_DATAPATH__abc_16259_n8535), .Y(AES_CORE_DATAPATH__abc_16259_n8536) );
  INVX1 INVX1_486 ( .A(AES_CORE_DATAPATH__abc_16259_n8542), .Y(AES_CORE_DATAPATH__abc_16259_n8543) );
  INVX1 INVX1_487 ( .A(AES_CORE_DATAPATH__abc_16259_n8549), .Y(AES_CORE_DATAPATH__abc_16259_n8550) );
  INVX1 INVX1_488 ( .A(AES_CORE_DATAPATH__abc_16259_n8556), .Y(AES_CORE_DATAPATH__abc_16259_n8557) );
  INVX1 INVX1_489 ( .A(AES_CORE_DATAPATH__abc_16259_n8569), .Y(AES_CORE_DATAPATH__abc_16259_n8570) );
  INVX1 INVX1_49 ( .A(AES_CORE_DATAPATH__abc_16259_n2922_1), .Y(AES_CORE_DATAPATH__abc_16259_n2923) );
  INVX1 INVX1_490 ( .A(AES_CORE_DATAPATH__abc_16259_n8694), .Y(AES_CORE_DATAPATH__abc_16259_n8695) );
  INVX1 INVX1_491 ( .A(AES_CORE_DATAPATH__abc_16259_n8704), .Y(AES_CORE_DATAPATH__abc_16259_n8705) );
  INVX1 INVX1_492 ( .A(AES_CORE_DATAPATH__abc_16259_n8723), .Y(AES_CORE_DATAPATH__abc_16259_n8724) );
  INVX1 INVX1_493 ( .A(AES_CORE_DATAPATH__abc_16259_n8742), .Y(AES_CORE_DATAPATH__abc_16259_n8743) );
  INVX1 INVX1_494 ( .A(AES_CORE_DATAPATH__abc_16259_n8761), .Y(AES_CORE_DATAPATH__abc_16259_n8762) );
  INVX1 INVX1_495 ( .A(AES_CORE_DATAPATH__abc_16259_n8798), .Y(AES_CORE_DATAPATH__abc_16259_n8799) );
  INVX1 INVX1_496 ( .A(AES_CORE_DATAPATH__abc_16259_n8901), .Y(AES_CORE_DATAPATH__abc_16259_n8902) );
  INVX1 INVX1_497 ( .A(AES_CORE_DATAPATH__abc_16259_n8906), .Y(AES_CORE_DATAPATH__abc_16259_n8907) );
  INVX1 INVX1_498 ( .A(AES_CORE_DATAPATH__abc_16259_n8914), .Y(AES_CORE_DATAPATH__abc_16259_n8915) );
  INVX1 INVX1_499 ( .A(AES_CORE_DATAPATH__abc_16259_n8929), .Y(AES_CORE_DATAPATH__abc_16259_n8930) );
  INVX1 INVX1_5 ( .A(AES_CORE_CONTROL_UNIT_rd_count_2_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n81_1) );
  INVX1 INVX1_50 ( .A(AES_CORE_DATAPATH__abc_16259_n2937), .Y(AES_CORE_DATAPATH__abc_16259_n2938_1) );
  INVX1 INVX1_500 ( .A(AES_CORE_DATAPATH__abc_16259_n8941), .Y(AES_CORE_DATAPATH__abc_16259_n8942) );
  INVX1 INVX1_501 ( .A(AES_CORE_DATAPATH__abc_16259_n8951), .Y(AES_CORE_DATAPATH__abc_16259_n8952) );
  INVX1 INVX1_502 ( .A(AES_CORE_DATAPATH__abc_16259_n8961), .Y(AES_CORE_DATAPATH__abc_16259_n8962) );
  INVX1 INVX1_503 ( .A(AES_CORE_DATAPATH_iv_3__6_), .Y(AES_CORE_DATAPATH__abc_16259_n8971) );
  INVX1 INVX1_504 ( .A(AES_CORE_DATAPATH__abc_16259_n8980), .Y(AES_CORE_DATAPATH__abc_16259_n8981) );
  INVX1 INVX1_505 ( .A(AES_CORE_DATAPATH__abc_16259_n8990), .Y(AES_CORE_DATAPATH__abc_16259_n8991) );
  INVX1 INVX1_506 ( .A(AES_CORE_DATAPATH__abc_16259_n9003), .Y(AES_CORE_DATAPATH__abc_16259_n9004) );
  INVX1 INVX1_507 ( .A(AES_CORE_DATAPATH__abc_16259_n9014), .Y(AES_CORE_DATAPATH__abc_16259_n9015) );
  INVX1 INVX1_508 ( .A(AES_CORE_DATAPATH__abc_16259_n9027), .Y(AES_CORE_DATAPATH__abc_16259_n9028) );
  INVX1 INVX1_509 ( .A(AES_CORE_DATAPATH__abc_16259_n9037), .Y(AES_CORE_DATAPATH__abc_16259_n9038) );
  INVX1 INVX1_51 ( .A(AES_CORE_DATAPATH__abc_16259_n2940_1), .Y(AES_CORE_DATAPATH__abc_16259_n2941) );
  INVX1 INVX1_510 ( .A(AES_CORE_DATAPATH__abc_16259_n9049), .Y(AES_CORE_DATAPATH__abc_16259_n9050) );
  INVX1 INVX1_511 ( .A(AES_CORE_DATAPATH__abc_16259_n9061), .Y(AES_CORE_DATAPATH__abc_16259_n9062) );
  INVX1 INVX1_512 ( .A(AES_CORE_DATAPATH__abc_16259_n9073), .Y(AES_CORE_DATAPATH__abc_16259_n9074) );
  INVX1 INVX1_513 ( .A(AES_CORE_DATAPATH__abc_16259_n9085), .Y(AES_CORE_DATAPATH__abc_16259_n9086) );
  INVX1 INVX1_514 ( .A(AES_CORE_DATAPATH__abc_16259_n9097), .Y(AES_CORE_DATAPATH__abc_16259_n9098) );
  INVX1 INVX1_515 ( .A(AES_CORE_DATAPATH__abc_16259_n9111), .Y(AES_CORE_DATAPATH__abc_16259_n9112) );
  INVX1 INVX1_516 ( .A(AES_CORE_DATAPATH__abc_16259_n9122), .Y(AES_CORE_DATAPATH__abc_16259_n9123) );
  INVX1 INVX1_517 ( .A(AES_CORE_DATAPATH__abc_16259_n9137), .Y(AES_CORE_DATAPATH__abc_16259_n9138) );
  INVX1 INVX1_518 ( .A(AES_CORE_DATAPATH_iv_3__21_), .Y(AES_CORE_DATAPATH__abc_16259_n9149) );
  INVX1 INVX1_519 ( .A(AES_CORE_DATAPATH__abc_16259_n9164), .Y(AES_CORE_DATAPATH__abc_16259_n9165) );
  INVX1 INVX1_52 ( .A(AES_CORE_DATAPATH_col_0__3_), .Y(AES_CORE_DATAPATH__abc_16259_n2953_1) );
  INVX1 INVX1_520 ( .A(AES_CORE_DATAPATH__abc_16259_n9175), .Y(AES_CORE_DATAPATH__abc_16259_n9176) );
  INVX1 INVX1_521 ( .A(AES_CORE_DATAPATH__abc_16259_n9190), .Y(AES_CORE_DATAPATH__abc_16259_n9191) );
  INVX1 INVX1_522 ( .A(AES_CORE_DATAPATH_iv_3__25_), .Y(AES_CORE_DATAPATH__abc_16259_n9202) );
  INVX1 INVX1_523 ( .A(AES_CORE_DATAPATH__abc_16259_n9215), .Y(AES_CORE_DATAPATH__abc_16259_n9216) );
  INVX1 INVX1_524 ( .A(AES_CORE_DATAPATH__abc_16259_n9227), .Y(AES_CORE_DATAPATH__abc_16259_n9228) );
  INVX1 INVX1_525 ( .A(AES_CORE_DATAPATH__abc_16259_n9239), .Y(AES_CORE_DATAPATH__abc_16259_n9240) );
  INVX1 INVX1_526 ( .A(AES_CORE_DATAPATH__abc_16259_n9251), .Y(AES_CORE_DATAPATH__abc_16259_n9252) );
  INVX1 INVX1_527 ( .A(AES_CORE_DATAPATH__abc_16259_n9262), .Y(AES_CORE_DATAPATH__abc_16259_n9263) );
  INVX1 INVX1_528 ( .A(AES_CORE_DATAPATH_iv_3__31_), .Y(AES_CORE_DATAPATH__abc_16259_n9275) );
  INVX1 INVX1_529 ( .A(AES_CORE_DATAPATH__abc_16259_n9319), .Y(AES_CORE_DATAPATH__abc_16259_n9320) );
  INVX1 INVX1_53 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_3_), .Y(AES_CORE_DATAPATH__abc_16259_n2955_1) );
  INVX1 INVX1_530 ( .A(AES_CORE_DATAPATH__abc_16259_n9323), .Y(AES_CORE_DATAPATH__abc_16259_n9324) );
  INVX1 INVX1_531 ( .A(AES_CORE_DATAPATH__abc_16259_n9330), .Y(AES_CORE_DATAPATH__abc_16259_n9331) );
  INVX1 INVX1_532 ( .A(AES_CORE_DATAPATH__abc_16259_n9337), .Y(AES_CORE_DATAPATH__abc_16259_n9338) );
  INVX1 INVX1_533 ( .A(AES_CORE_DATAPATH__abc_16259_n9344), .Y(AES_CORE_DATAPATH__abc_16259_n9345) );
  INVX1 INVX1_534 ( .A(AES_CORE_DATAPATH__abc_16259_n9357), .Y(AES_CORE_DATAPATH__abc_16259_n9358) );
  INVX1 INVX1_535 ( .A(AES_CORE_DATAPATH__abc_16259_n9471), .Y(AES_CORE_DATAPATH__abc_16259_n9472) );
  INVX1 INVX1_536 ( .A(AES_CORE_DATAPATH__abc_16259_n9480), .Y(AES_CORE_DATAPATH__abc_16259_n9481) );
  INVX1 INVX1_537 ( .A(AES_CORE_DATAPATH__abc_16259_n9497), .Y(AES_CORE_DATAPATH__abc_16259_n9498) );
  INVX1 INVX1_538 ( .A(AES_CORE_DATAPATH__abc_16259_n9514), .Y(AES_CORE_DATAPATH__abc_16259_n9515) );
  INVX1 INVX1_539 ( .A(AES_CORE_DATAPATH__abc_16259_n9531), .Y(AES_CORE_DATAPATH__abc_16259_n9532) );
  INVX1 INVX1_54 ( .A(AES_CORE_DATAPATH__abc_16259_n2962), .Y(AES_CORE_DATAPATH__abc_16259_n2963) );
  INVX1 INVX1_540 ( .A(AES_CORE_DATAPATH__abc_16259_n9564), .Y(AES_CORE_DATAPATH__abc_16259_n9565) );
  INVX1 INVX1_541 ( .A(AES_CORE_DATAPATH__abc_16259_n9784), .Y(AES_CORE_DATAPATH__abc_16259_n9785) );
  INVX1 INVX1_542 ( .A(AES_CORE_DATAPATH__abc_16259_n9788), .Y(AES_CORE_DATAPATH__abc_16259_n9789) );
  INVX1 INVX1_543 ( .A(AES_CORE_DATAPATH__abc_16259_n9795), .Y(AES_CORE_DATAPATH__abc_16259_n9796) );
  INVX1 INVX1_544 ( .A(AES_CORE_DATAPATH__abc_16259_n9802), .Y(AES_CORE_DATAPATH__abc_16259_n9803) );
  INVX1 INVX1_545 ( .A(AES_CORE_DATAPATH__abc_16259_n9809), .Y(AES_CORE_DATAPATH__abc_16259_n9810) );
  INVX1 INVX1_546 ( .A(AES_CORE_DATAPATH__abc_16259_n9822), .Y(AES_CORE_DATAPATH__abc_16259_n9823) );
  INVX1 INVX1_547 ( .A(AES_CORE_DATAPATH__abc_16259_n9936), .Y(AES_CORE_DATAPATH__abc_16259_n9937) );
  INVX1 INVX1_548 ( .A(AES_CORE_DATAPATH__abc_16259_n9945), .Y(AES_CORE_DATAPATH__abc_16259_n9946) );
  INVX1 INVX1_549 ( .A(AES_CORE_DATAPATH__abc_16259_n9962), .Y(AES_CORE_DATAPATH__abc_16259_n9963) );
  INVX1 INVX1_55 ( .A(AES_CORE_DATAPATH__abc_16259_n2977), .Y(AES_CORE_DATAPATH__abc_16259_n2978_1) );
  INVX1 INVX1_550 ( .A(AES_CORE_DATAPATH__abc_16259_n9979), .Y(AES_CORE_DATAPATH__abc_16259_n9980) );
  INVX1 INVX1_551 ( .A(AES_CORE_DATAPATH__abc_16259_n9996), .Y(AES_CORE_DATAPATH__abc_16259_n9997) );
  INVX1 INVX1_552 ( .A(AES_CORE_DATAPATH__abc_16259_n10029), .Y(AES_CORE_DATAPATH__abc_16259_n10030) );
  INVX1 INVX1_553 ( .A(AES_CORE_DATAPATH__abc_16259_n10249), .Y(AES_CORE_DATAPATH__abc_16259_n10250) );
  INVX1 INVX1_554 ( .A(AES_CORE_DATAPATH__abc_16259_n10253), .Y(AES_CORE_DATAPATH__abc_16259_n10254) );
  INVX1 INVX1_555 ( .A(AES_CORE_DATAPATH__abc_16259_n10260), .Y(AES_CORE_DATAPATH__abc_16259_n10261) );
  INVX1 INVX1_556 ( .A(AES_CORE_DATAPATH__abc_16259_n10267), .Y(AES_CORE_DATAPATH__abc_16259_n10268) );
  INVX1 INVX1_557 ( .A(AES_CORE_DATAPATH__abc_16259_n10274), .Y(AES_CORE_DATAPATH__abc_16259_n10275) );
  INVX1 INVX1_558 ( .A(AES_CORE_DATAPATH__abc_16259_n10287), .Y(AES_CORE_DATAPATH__abc_16259_n10288) );
  INVX1 INVX1_559 ( .A(AES_CORE_DATAPATH__abc_16259_n10401), .Y(AES_CORE_DATAPATH__abc_16259_n10402) );
  INVX1 INVX1_56 ( .A(AES_CORE_DATAPATH__abc_16259_n2980_1), .Y(AES_CORE_DATAPATH__abc_16259_n2981) );
  INVX1 INVX1_560 ( .A(AES_CORE_DATAPATH__abc_16259_n10410), .Y(AES_CORE_DATAPATH__abc_16259_n10411) );
  INVX1 INVX1_561 ( .A(AES_CORE_DATAPATH__abc_16259_n10427), .Y(AES_CORE_DATAPATH__abc_16259_n10428) );
  INVX1 INVX1_562 ( .A(AES_CORE_DATAPATH__abc_16259_n10444), .Y(AES_CORE_DATAPATH__abc_16259_n10445) );
  INVX1 INVX1_563 ( .A(AES_CORE_DATAPATH__abc_16259_n10461), .Y(AES_CORE_DATAPATH__abc_16259_n10462) );
  INVX1 INVX1_564 ( .A(AES_CORE_DATAPATH__abc_16259_n10494), .Y(AES_CORE_DATAPATH__abc_16259_n10495) );
  INVX1 INVX1_565 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__0_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n327_1) );
  INVX1 INVX1_566 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__0_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n329_1) );
  INVX1 INVX1_567 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n331_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n332_1) );
  INVX1 INVX1_568 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n333_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n335_1) );
  INVX1 INVX1_569 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__1_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n338_1) );
  INVX1 INVX1_57 ( .A(AES_CORE_DATAPATH_col_0__4_), .Y(AES_CORE_DATAPATH__abc_16259_n2993) );
  INVX1 INVX1_570 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__1_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n340_1) );
  INVX1 INVX1_571 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n342_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n343_1) );
  INVX1 INVX1_572 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n344_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n346_1) );
  INVX1 INVX1_573 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__2_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n349_1) );
  INVX1 INVX1_574 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__2_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n351_1) );
  INVX1 INVX1_575 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n353_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n354_1) );
  INVX1 INVX1_576 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n355_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n357_1) );
  INVX1 INVX1_577 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__3_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n360_1) );
  INVX1 INVX1_578 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__3_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n362_1) );
  INVX1 INVX1_579 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n364_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n365_1) );
  INVX1 INVX1_58 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_4_), .Y(AES_CORE_DATAPATH__abc_16259_n2995) );
  INVX1 INVX1_580 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n366_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n368_1) );
  INVX1 INVX1_581 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__4_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n371_1) );
  INVX1 INVX1_582 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__4_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n373_1) );
  INVX1 INVX1_583 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n375_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n376_1) );
  INVX1 INVX1_584 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n377_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n379_1) );
  INVX1 INVX1_585 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__5_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n382_1) );
  INVX1 INVX1_586 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__5_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n384_1) );
  INVX1 INVX1_587 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n386_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n387_1) );
  INVX1 INVX1_588 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n388_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n390_1) );
  INVX1 INVX1_589 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__6_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n393_1) );
  INVX1 INVX1_59 ( .A(AES_CORE_DATAPATH__abc_16259_n3002), .Y(AES_CORE_DATAPATH__abc_16259_n3003_1) );
  INVX1 INVX1_590 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__6_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n395_1) );
  INVX1 INVX1_591 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n397_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n398_1) );
  INVX1 INVX1_592 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n399_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n401_1) );
  INVX1 INVX1_593 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__7_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n404_1) );
  INVX1 INVX1_594 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__7_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n406_1) );
  INVX1 INVX1_595 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n408_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n409_1) );
  INVX1 INVX1_596 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n410_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n412_1) );
  INVX1 INVX1_597 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__8_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n415_1) );
  INVX1 INVX1_598 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__8_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n417_1) );
  INVX1 INVX1_599 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n419_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n420_1) );
  INVX1 INVX1_6 ( .A(\aes_mode[1] ), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n88) );
  INVX1 INVX1_60 ( .A(AES_CORE_DATAPATH__abc_16259_n3017), .Y(AES_CORE_DATAPATH__abc_16259_n3018) );
  INVX1 INVX1_600 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n421_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n423_1) );
  INVX1 INVX1_601 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__9_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n426_1) );
  INVX1 INVX1_602 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__9_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n428_1) );
  INVX1 INVX1_603 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n430_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n431_1) );
  INVX1 INVX1_604 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n432_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n434_1) );
  INVX1 INVX1_605 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__10_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n437_1) );
  INVX1 INVX1_606 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__10_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n439_1) );
  INVX1 INVX1_607 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n441_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n442_1) );
  INVX1 INVX1_608 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n443_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n445_1) );
  INVX1 INVX1_609 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__11_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n448_1) );
  INVX1 INVX1_61 ( .A(AES_CORE_DATAPATH__abc_16259_n3020), .Y(AES_CORE_DATAPATH__abc_16259_n3021) );
  INVX1 INVX1_610 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__11_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n450_1) );
  INVX1 INVX1_611 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n452_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n453_1) );
  INVX1 INVX1_612 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n454_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n456_1) );
  INVX1 INVX1_613 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__12_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n459_1) );
  INVX1 INVX1_614 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__12_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n461_1) );
  INVX1 INVX1_615 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n463_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n464_1) );
  INVX1 INVX1_616 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n465_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n467_1) );
  INVX1 INVX1_617 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__13_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n470_1) );
  INVX1 INVX1_618 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__13_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n472_1) );
  INVX1 INVX1_619 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n474_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n475_1) );
  INVX1 INVX1_62 ( .A(AES_CORE_DATAPATH_col_0__5_), .Y(AES_CORE_DATAPATH__abc_16259_n3033_1) );
  INVX1 INVX1_620 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n476_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n478_1) );
  INVX1 INVX1_621 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__14_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n481_1) );
  INVX1 INVX1_622 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__14_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n483_1) );
  INVX1 INVX1_623 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n485_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n486_1) );
  INVX1 INVX1_624 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n487_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n489_1) );
  INVX1 INVX1_625 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__15_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n492_1) );
  INVX1 INVX1_626 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__15_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n494_1) );
  INVX1 INVX1_627 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n496_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n497_1) );
  INVX1 INVX1_628 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n498_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n500_1) );
  INVX1 INVX1_629 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__16_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n503) );
  INVX1 INVX1_63 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_5_), .Y(AES_CORE_DATAPATH__abc_16259_n3035) );
  INVX1 INVX1_630 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__16_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n505) );
  INVX1 INVX1_631 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n507), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n508) );
  INVX1 INVX1_632 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n509), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n511) );
  INVX1 INVX1_633 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__17_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n514) );
  INVX1 INVX1_634 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__17_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n516) );
  INVX1 INVX1_635 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n518), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n519) );
  INVX1 INVX1_636 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n520), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n522) );
  INVX1 INVX1_637 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__18_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n525) );
  INVX1 INVX1_638 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__18_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n527) );
  INVX1 INVX1_639 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n529), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n530) );
  INVX1 INVX1_64 ( .A(AES_CORE_DATAPATH__abc_16259_n3042_1), .Y(AES_CORE_DATAPATH__abc_16259_n3043) );
  INVX1 INVX1_640 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n531), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n533) );
  INVX1 INVX1_641 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__19_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n536) );
  INVX1 INVX1_642 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__19_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n538) );
  INVX1 INVX1_643 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n540), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n541) );
  INVX1 INVX1_644 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n542), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n544) );
  INVX1 INVX1_645 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__20_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n547) );
  INVX1 INVX1_646 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__20_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n549) );
  INVX1 INVX1_647 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n551), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n552) );
  INVX1 INVX1_648 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n553), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n555) );
  INVX1 INVX1_649 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__21_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n558) );
  INVX1 INVX1_65 ( .A(AES_CORE_DATAPATH__abc_16259_n3057), .Y(AES_CORE_DATAPATH__abc_16259_n3058) );
  INVX1 INVX1_650 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__21_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n560) );
  INVX1 INVX1_651 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n562), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n563) );
  INVX1 INVX1_652 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n564), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n566) );
  INVX1 INVX1_653 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__22_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n569) );
  INVX1 INVX1_654 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__22_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n571) );
  INVX1 INVX1_655 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n573), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n574) );
  INVX1 INVX1_656 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n575), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n577) );
  INVX1 INVX1_657 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__23_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n580) );
  INVX1 INVX1_658 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__23_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n582) );
  INVX1 INVX1_659 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n584), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n585) );
  INVX1 INVX1_66 ( .A(AES_CORE_DATAPATH__abc_16259_n3060), .Y(AES_CORE_DATAPATH__abc_16259_n3061_1) );
  INVX1 INVX1_660 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n586), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n588) );
  INVX1 INVX1_661 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n592), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n593) );
  INVX1 INVX1_662 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n594), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n595) );
  INVX1 INVX1_663 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_round_2_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n598) );
  INVX1 INVX1_664 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_round_1_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n599) );
  INVX1 INVX1_665 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n601), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n602) );
  INVX1 INVX1_666 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n608), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n609) );
  INVX1 INVX1_667 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n612), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n613) );
  INVX1 INVX1_668 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n618), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n619) );
  INVX1 INVX1_669 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n620), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n621) );
  INVX1 INVX1_67 ( .A(AES_CORE_DATAPATH_col_0__6_), .Y(AES_CORE_DATAPATH__abc_16259_n3073) );
  INVX1 INVX1_670 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_25_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n622) );
  INVX1 INVX1_671 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_round_0_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n623) );
  INVX1 INVX1_672 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n632), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n633) );
  INVX1 INVX1_673 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n637), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n638) );
  INVX1 INVX1_674 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n628), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n642) );
  INVX1 INVX1_675 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n634), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n643) );
  INVX1 INVX1_676 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n651), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n652) );
  INVX1 INVX1_677 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n653), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n654) );
  INVX1 INVX1_678 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_26_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n655) );
  INVX1 INVX1_679 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_round_3_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n656) );
  INVX1 INVX1_68 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_6_), .Y(AES_CORE_DATAPATH__abc_16259_n3075) );
  INVX1 INVX1_680 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n661), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n662) );
  INVX1 INVX1_681 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n670), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n671) );
  INVX1 INVX1_682 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n673), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n674) );
  INVX1 INVX1_683 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n604), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n679) );
  INVX1 INVX1_684 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n691), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n692) );
  INVX1 INVX1_685 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n693), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n694) );
  INVX1 INVX1_686 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n702), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n703) );
  INVX1 INVX1_687 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n706), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n708) );
  INVX1 INVX1_688 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n712), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n713) );
  INVX1 INVX1_689 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n714), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n715) );
  INVX1 INVX1_69 ( .A(AES_CORE_DATAPATH__abc_16259_n3082), .Y(AES_CORE_DATAPATH__abc_16259_n3083_1) );
  INVX1 INVX1_690 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_28_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n716) );
  INVX1 INVX1_691 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n720), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n721) );
  INVX1 INVX1_692 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n722), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n723) );
  INVX1 INVX1_693 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n725), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n728) );
  INVX1 INVX1_694 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n741), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n742) );
  INVX1 INVX1_695 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n743), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n744) );
  INVX1 INVX1_696 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_29_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n745) );
  INVX1 INVX1_697 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n719), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n746) );
  INVX1 INVX1_698 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n629), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n749) );
  INVX1 INVX1_699 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n753), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n754) );
  INVX1 INVX1_7 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n91), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n92) );
  INVX1 INVX1_70 ( .A(AES_CORE_DATAPATH__abc_16259_n3097), .Y(AES_CORE_DATAPATH__abc_16259_n3098_1) );
  INVX1 INVX1_700 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n751), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n761) );
  INVX1 INVX1_701 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n769), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n770) );
  INVX1 INVX1_702 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n771), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n772) );
  INVX1 INVX1_703 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_30_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n773) );
  INVX1 INVX1_704 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n666), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n774) );
  INVX1 INVX1_705 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n776), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n777) );
  INVX1 INVX1_706 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n778), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n779) );
  INVX1 INVX1_707 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n783), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n784) );
  INVX1 INVX1_708 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n801), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n802) );
  INVX1 INVX1_709 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n803), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n804) );
  INVX1 INVX1_71 ( .A(AES_CORE_DATAPATH__abc_16259_n3100_1), .Y(AES_CORE_DATAPATH__abc_16259_n3101) );
  INVX1 INVX1_710 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_31_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n805) );
  INVX1 INVX1_711 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n660), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n806) );
  INVX1 INVX1_712 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n808), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n809) );
  INVX1 INVX1_713 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n825), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n826) );
  INVX1 INVX1_714 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n832), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n833) );
  INVX1 INVX1_715 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n839), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n840) );
  INVX1 INVX1_716 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n846), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n847) );
  INVX1 INVX1_717 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n853), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n854) );
  INVX1 INVX1_718 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n860), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n861) );
  INVX1 INVX1_719 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n867), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n868) );
  INVX1 INVX1_72 ( .A(AES_CORE_DATAPATH_col_0__7_), .Y(AES_CORE_DATAPATH__abc_16259_n3113) );
  INVX1 INVX1_720 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n874), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n875) );
  INVX1 INVX1_721 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n881), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n882) );
  INVX1 INVX1_722 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n888), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n889) );
  INVX1 INVX1_723 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n895), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n896) );
  INVX1 INVX1_724 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n902), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n903) );
  INVX1 INVX1_725 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n909), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n910) );
  INVX1 INVX1_726 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n916), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n917) );
  INVX1 INVX1_727 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n923), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n924) );
  INVX1 INVX1_728 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n930), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n931) );
  INVX1 INVX1_729 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n937), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n938) );
  INVX1 INVX1_73 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_7_), .Y(AES_CORE_DATAPATH__abc_16259_n3115) );
  INVX1 INVX1_730 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n944), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n945) );
  INVX1 INVX1_731 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n951), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n952) );
  INVX1 INVX1_732 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n958), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n959) );
  INVX1 INVX1_733 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n965), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n966) );
  INVX1 INVX1_734 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n972), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n973) );
  INVX1 INVX1_735 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n979), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n980) );
  INVX1 INVX1_736 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n986), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n987) );
  INVX1 INVX1_737 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n993), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n994) );
  INVX1 INVX1_738 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1000), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1001) );
  INVX1 INVX1_739 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1007), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1008) );
  INVX1 INVX1_74 ( .A(AES_CORE_DATAPATH__abc_16259_n3122), .Y(AES_CORE_DATAPATH__abc_16259_n3123_1) );
  INVX1 INVX1_740 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1014), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1015) );
  INVX1 INVX1_741 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1021), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1022) );
  INVX1 INVX1_742 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1028), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1029) );
  INVX1 INVX1_743 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1035), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1036) );
  INVX1 INVX1_744 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1042), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1043) );
  INVX1 INVX1_745 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1049), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1050) );
  INVX1 INVX1_746 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1053), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1054) );
  INVX1 INVX1_747 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1057), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1058) );
  INVX1 INVX1_748 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1061), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1062) );
  INVX1 INVX1_749 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1065), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1066) );
  INVX1 INVX1_75 ( .A(AES_CORE_DATAPATH__abc_16259_n3137), .Y(AES_CORE_DATAPATH__abc_16259_n3138) );
  INVX1 INVX1_750 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1069), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1070) );
  INVX1 INVX1_751 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1073), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1074) );
  INVX1 INVX1_752 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1077), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1078) );
  INVX1 INVX1_753 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1081), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1082) );
  INVX1 INVX1_754 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1085), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1086) );
  INVX1 INVX1_755 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1089), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1090) );
  INVX1 INVX1_756 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1093), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1094) );
  INVX1 INVX1_757 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1097), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1098) );
  INVX1 INVX1_758 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1101), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1102) );
  INVX1 INVX1_759 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1105), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1106) );
  INVX1 INVX1_76 ( .A(AES_CORE_DATAPATH__abc_16259_n3140), .Y(AES_CORE_DATAPATH__abc_16259_n3141_1) );
  INVX1 INVX1_760 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1109), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1110) );
  INVX1 INVX1_761 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1113), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1114) );
  INVX1 INVX1_762 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1117), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1118) );
  INVX1 INVX1_763 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1121), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1122) );
  INVX1 INVX1_764 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1125), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1126) );
  INVX1 INVX1_765 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1129), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1130) );
  INVX1 INVX1_766 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1133), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1134) );
  INVX1 INVX1_767 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1137), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1138) );
  INVX1 INVX1_768 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1141), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1142) );
  INVX1 INVX1_769 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__24_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1144) );
  INVX1 INVX1_77 ( .A(AES_CORE_DATAPATH_col_0__8_), .Y(AES_CORE_DATAPATH__abc_16259_n3153) );
  INVX1 INVX1_770 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n611), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1145) );
  INVX1 INVX1_771 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__25_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1149) );
  INVX1 INVX1_772 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__26_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1154) );
  INVX1 INVX1_773 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__27_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1157) );
  INVX1 INVX1_774 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n705), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1158) );
  INVX1 INVX1_775 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__28_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1162) );
  INVX1 INVX1_776 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__29_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1167) );
  INVX1 INVX1_777 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__30_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1171) );
  INVX1 INVX1_778 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__31_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1175) );
  INVX1 INVX1_779 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1179), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1180) );
  INVX1 INVX1_78 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_8_), .Y(AES_CORE_DATAPATH__abc_16259_n3155) );
  INVX1 INVX1_780 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1183), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1184) );
  INVX1 INVX1_781 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1187), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1188) );
  INVX1 INVX1_782 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1191), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1192) );
  INVX1 INVX1_783 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1195), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1196) );
  INVX1 INVX1_784 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1199), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1200) );
  INVX1 INVX1_785 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1203), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1204) );
  INVX1 INVX1_786 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1207), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1208) );
  INVX1 INVX1_787 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1211), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1212) );
  INVX1 INVX1_788 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1215), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1216) );
  INVX1 INVX1_789 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1219), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1220) );
  INVX1 INVX1_79 ( .A(AES_CORE_DATAPATH__abc_16259_n3162), .Y(AES_CORE_DATAPATH__abc_16259_n3163) );
  INVX1 INVX1_790 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1223), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1224) );
  INVX1 INVX1_791 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1227), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1228) );
  INVX1 INVX1_792 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1231), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1232) );
  INVX1 INVX1_793 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1235), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1236) );
  INVX1 INVX1_794 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1239), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1240) );
  INVX1 INVX1_795 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1243), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1244) );
  INVX1 INVX1_796 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1247), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1248) );
  INVX1 INVX1_797 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1251), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1252) );
  INVX1 INVX1_798 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1255), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1256) );
  INVX1 INVX1_799 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1259), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1260) );
  INVX1 INVX1_8 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n90), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n96_1) );
  INVX1 INVX1_80 ( .A(AES_CORE_DATAPATH__abc_16259_n3177_1), .Y(AES_CORE_DATAPATH__abc_16259_n3178_1) );
  INVX1 INVX1_800 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1263), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1264) );
  INVX1 INVX1_801 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1267), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1268) );
  INVX1 INVX1_802 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1271), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1272) );
  INVX1 INVX1_803 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1275), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1276) );
  INVX1 INVX1_804 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1279), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1280) );
  INVX1 INVX1_805 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1283), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1284) );
  INVX1 INVX1_806 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1287), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1288) );
  INVX1 INVX1_807 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1291), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1292) );
  INVX1 INVX1_808 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1295), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1296) );
  INVX1 INVX1_809 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1299), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1300) );
  INVX1 INVX1_81 ( .A(AES_CORE_DATAPATH__abc_16259_n3180), .Y(AES_CORE_DATAPATH__abc_16259_n3181_1) );
  INVX1 INVX1_810 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1303), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1304) );
  INVX1 INVX1_811 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n97_1) );
  INVX1 INVX1_812 ( .A(AES_CORE_DATAPATH_MIX_COL_col_3__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n98) );
  INVX1 INVX1_813 ( .A(AES_CORE_DATAPATH_MIX_COL_col_3__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n102) );
  INVX1 INVX1_814 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n104) );
  INVX1 INVX1_815 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n109_1) );
  INVX1 INVX1_816 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n100), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n114) );
  INVX1 INVX1_817 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n111), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n116) );
  INVX1 INVX1_818 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n119_1) );
  INVX1 INVX1_819 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n120) );
  INVX1 INVX1_82 ( .A(AES_CORE_DATAPATH_col_0__9_), .Y(AES_CORE_DATAPATH__abc_16259_n3193) );
  INVX1 INVX1_820 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n121) );
  INVX1 INVX1_821 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n126), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n127_1) );
  INVX1 INVX1_822 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n130), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n131) );
  INVX1 INVX1_823 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n134_1) );
  INVX1 INVX1_824 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n138) );
  INVX1 INVX1_825 ( .A(AES_CORE_DATAPATH_MIX_COL_col_3__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n139) );
  INVX1 INVX1_826 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n123_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n146) );
  INVX1 INVX1_827 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n163), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n164) );
  INVX1 INVX1_828 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n166_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n167) );
  INVX1 INVX1_829 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n169), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n170) );
  INVX1 INVX1_83 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_9_), .Y(AES_CORE_DATAPATH__abc_16259_n3195) );
  INVX1 INVX1_830 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n173) );
  INVX1 INVX1_831 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n174_1) );
  INVX1 INVX1_832 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n179), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n180_1) );
  INVX1 INVX1_833 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n183_1), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_1_) );
  INVX1 INVX1_834 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n186), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n187_1) );
  INVX1 INVX1_835 ( .A(AES_CORE_DATAPATH_MIX_COL_col_3__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n196) );
  INVX1 INVX1_836 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n198_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n202) );
  INVX1 INVX1_837 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n222_1) );
  INVX1 INVX1_838 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n225_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n226) );
  INVX1 INVX1_839 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n228_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n229) );
  INVX1 INVX1_84 ( .A(AES_CORE_DATAPATH__abc_16259_n3202), .Y(AES_CORE_DATAPATH__abc_16259_n3203) );
  INVX1 INVX1_840 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n232) );
  INVX1 INVX1_841 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n234), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n235) );
  INVX1 INVX1_842 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n240), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n241) );
  INVX1 INVX1_843 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n248) );
  INVX1 INVX1_844 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n250), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n254) );
  INVX1 INVX1_845 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n263), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n264) );
  INVX1 INVX1_846 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n270), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n271) );
  INVX1 INVX1_847 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n273) );
  INVX1 INVX1_848 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n277) );
  INVX1 INVX1_849 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n280), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n281) );
  INVX1 INVX1_85 ( .A(AES_CORE_DATAPATH__abc_16259_n3217), .Y(AES_CORE_DATAPATH__abc_16259_n3218) );
  INVX1 INVX1_850 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n283), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n284) );
  INVX1 INVX1_851 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n287) );
  INVX1 INVX1_852 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n291) );
  INVX1 INVX1_853 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n289), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n292) );
  INVX1 INVX1_854 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n294), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n295) );
  INVX1 INVX1_855 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n298), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_3_) );
  INVX1 INVX1_856 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n316), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n317) );
  INVX1 INVX1_857 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n340) );
  INVX1 INVX1_858 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n343), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n344) );
  INVX1 INVX1_859 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n346), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n347) );
  INVX1 INVX1_86 ( .A(AES_CORE_DATAPATH__abc_16259_n3220), .Y(AES_CORE_DATAPATH__abc_16259_n3221) );
  INVX1 INVX1_860 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__4_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n348) );
  INVX1 INVX1_861 ( .A(AES_CORE_DATAPATH_MIX_COL_col_3__4_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n350) );
  INVX1 INVX1_862 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n352), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n353) );
  INVX1 INVX1_863 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__4_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n355) );
  INVX1 INVX1_864 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n357), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n358) );
  INVX1 INVX1_865 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n361), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_4_) );
  INVX1 INVX1_866 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n364) );
  INVX1 INVX1_867 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n366), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n368) );
  INVX1 INVX1_868 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n403), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n404) );
  INVX1 INVX1_869 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__4_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n405) );
  INVX1 INVX1_87 ( .A(AES_CORE_DATAPATH_col_0__10_), .Y(AES_CORE_DATAPATH__abc_16259_n3233) );
  INVX1 INVX1_870 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n408), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n409) );
  INVX1 INVX1_871 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n412), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_5_) );
  INVX1 INVX1_872 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n415), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n416) );
  INVX1 INVX1_873 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n417), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n418) );
  INVX1 INVX1_874 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n421), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n432) );
  INVX1 INVX1_875 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n447), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n448) );
  INVX1 INVX1_876 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n450), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n455) );
  INVX1 INVX1_877 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n453), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n456) );
  INVX1 INVX1_878 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n459) );
  INVX1 INVX1_879 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n465), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n466) );
  INVX1 INVX1_88 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_10_), .Y(AES_CORE_DATAPATH__abc_16259_n3235_1) );
  INVX1 INVX1_880 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n462), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n471) );
  INVX1 INVX1_881 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n469), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n472) );
  INVX1 INVX1_882 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n474), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n475) );
  INVX1 INVX1_883 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n481), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n482) );
  INVX1 INVX1_884 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n485), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n487) );
  INVX1 INVX1_885 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n490) );
  INVX1 INVX1_886 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n493), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n494) );
  INVX1 INVX1_887 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n497), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n499) );
  INVX1 INVX1_888 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n507), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n508) );
  INVX1 INVX1_889 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_8_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n513) );
  INVX1 INVX1_89 ( .A(AES_CORE_DATAPATH__abc_16259_n3242), .Y(AES_CORE_DATAPATH__abc_16259_n3243_1) );
  INVX1 INVX1_890 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n516), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n517) );
  INVX1 INVX1_891 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n523), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n524) );
  INVX1 INVX1_892 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n530), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n531) );
  INVX1 INVX1_893 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n532), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n533) );
  INVX1 INVX1_894 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n535), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_9_) );
  INVX1 INVX1_895 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n539), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n541) );
  INVX1 INVX1_896 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n549), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n550) );
  INVX1 INVX1_897 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n546), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n552) );
  INVX1 INVX1_898 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_10_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n555) );
  INVX1 INVX1_899 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n558), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n560) );
  INVX1 INVX1_9 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n76_1), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n103) );
  INVX1 INVX1_90 ( .A(AES_CORE_DATAPATH__abc_16259_n3257_1), .Y(AES_CORE_DATAPATH__abc_16259_n3258) );
  INVX1 INVX1_900 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n565), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n566) );
  INVX1 INVX1_901 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n569), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n570) );
  INVX1 INVX1_902 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n573), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n574) );
  INVX1 INVX1_903 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_11_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n582) );
  INVX1 INVX1_904 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n590), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n591) );
  INVX1 INVX1_905 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n594), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n595) );
  INVX1 INVX1_906 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n598), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n599) );
  INVX1 INVX1_907 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_12_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n607) );
  INVX1 INVX1_908 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n618), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n619) );
  INVX1 INVX1_909 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n615), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n621) );
  INVX1 INVX1_91 ( .A(AES_CORE_DATAPATH__abc_16259_n3260), .Y(AES_CORE_DATAPATH__abc_16259_n3261) );
  INVX1 INVX1_910 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_13_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n624) );
  INVX1 INVX1_911 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n636), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n637) );
  INVX1 INVX1_912 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n640), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n641) );
  INVX1 INVX1_913 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n644), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_14_) );
  INVX1 INVX1_914 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n648), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n650) );
  INVX1 INVX1_915 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n662), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n663) );
  INVX1 INVX1_916 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n655), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n665) );
  INVX1 INVX1_917 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n667), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_15_) );
  INVX1 INVX1_918 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n671), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n673) );
  INVX1 INVX1_919 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n681), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n682) );
  INVX1 INVX1_92 ( .A(AES_CORE_DATAPATH_col_0__11_), .Y(AES_CORE_DATAPATH__abc_16259_n3273) );
  INVX1 INVX1_920 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_16_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n687) );
  INVX1 INVX1_921 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n693), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n694) );
  INVX1 INVX1_922 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n697), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n698) );
  INVX1 INVX1_923 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n701), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n702) );
  INVX1 INVX1_924 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n705), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_17_) );
  INVX1 INVX1_925 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n712), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n717) );
  INVX1 INVX1_926 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n715), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n718) );
  INVX1 INVX1_927 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_18_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n721) );
  INVX1 INVX1_928 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n727), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n729) );
  INVX1 INVX1_929 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n735), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n736) );
  INVX1 INVX1_93 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_11_), .Y(AES_CORE_DATAPATH__abc_16259_n3275) );
  INVX1 INVX1_930 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_19_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n740) );
  INVX1 INVX1_931 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n746), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n747) );
  INVX1 INVX1_932 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n749), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n750) );
  INVX1 INVX1_933 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n753), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n754) );
  INVX1 INVX1_934 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n757), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_20_) );
  INVX1 INVX1_935 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n765), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n766) );
  INVX1 INVX1_936 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n768), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n770) );
  INVX1 INVX1_937 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n772), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_21_) );
  INVX1 INVX1_938 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n779), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n780) );
  INVX1 INVX1_939 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n783), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n784) );
  INVX1 INVX1_94 ( .A(AES_CORE_DATAPATH__abc_16259_n3282), .Y(AES_CORE_DATAPATH__abc_16259_n3283) );
  INVX1 INVX1_940 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_22_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n788) );
  INVX1 INVX1_941 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n797), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n798) );
  INVX1 INVX1_942 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n799), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n800) );
  INVX1 INVX1_943 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n802), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_23_) );
  INVX1 INVX1_944 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n809), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n810) );
  INVX1 INVX1_945 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_24_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n814) );
  INVX1 INVX1_946 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n821), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n822) );
  INVX1 INVX1_947 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n824), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n825) );
  INVX1 INVX1_948 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n829), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n830) );
  INVX1 INVX1_949 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n832), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_25_) );
  INVX1 INVX1_95 ( .A(AES_CORE_DATAPATH__abc_16259_n3297_1), .Y(AES_CORE_DATAPATH__abc_16259_n3298) );
  INVX1 INVX1_950 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n841), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n842) );
  INVX1 INVX1_951 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n843), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n844) );
  INVX1 INVX1_952 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n847), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_26_) );
  INVX1 INVX1_953 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n855), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n856) );
  INVX1 INVX1_954 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n858), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n859) );
  INVX1 INVX1_955 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n862), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n863) );
  INVX1 INVX1_956 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_27_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n868) );
  INVX1 INVX1_957 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n873), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n874) );
  INVX1 INVX1_958 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n878), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n879) );
  INVX1 INVX1_959 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n881), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n882) );
  INVX1 INVX1_96 ( .A(AES_CORE_DATAPATH__abc_16259_n3300), .Y(AES_CORE_DATAPATH__abc_16259_n3301_1) );
  INVX1 INVX1_960 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n885), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_28_) );
  INVX1 INVX1_961 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n892), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n893) );
  INVX1 INVX1_962 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n896), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n898) );
  INVX1 INVX1_963 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n900), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_29_) );
  INVX1 INVX1_964 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n907), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n909) );
  INVX1 INVX1_965 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n911), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n912) );
  INVX1 INVX1_966 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_30_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n916) );
  INVX1 INVX1_967 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n922), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n923) );
  INVX1 INVX1_968 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n926), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_31_) );
  INVX1 INVX1_969 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n50) );
  INVX1 INVX1_97 ( .A(AES_CORE_DATAPATH_col_0__12_), .Y(AES_CORE_DATAPATH__abc_16259_n3313) );
  INVX1 INVX1_970 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n52) );
  INVX1 INVX1_971 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n54_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n55) );
  INVX1 INVX1_972 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n56) );
  INVX1 INVX1_973 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n58) );
  INVX1 INVX1_974 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n60), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n61) );
  INVX1 INVX1_975 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n67) );
  INVX1 INVX1_976 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n72) );
  INVX1 INVX1_977 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n70), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n73) );
  INVX1 INVX1_978 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n79) );
  INVX1 INVX1_979 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n86_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n87) );
  INVX1 INVX1_98 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_12_), .Y(AES_CORE_DATAPATH__abc_16259_n3315_1) );
  INVX1 INVX1_980 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n92), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n93) );
  INVX1 INVX1_981 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n95), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n96) );
  INVX1 INVX1_982 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n104_1) );
  INVX1 INVX1_983 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n107), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n109) );
  INVX1 INVX1_984 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n112), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n113) );
  INVX1 INVX1_985 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n114), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_7_) );
  INVX1 INVX1_986 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n116), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n117) );
  INVX1 INVX1_987 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n121_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n122) );
  INVX1 INVX1_988 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n126_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_0_) );
  INVX1 INVX1_989 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n130), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n131) );
  INVX1 INVX1_99 ( .A(AES_CORE_DATAPATH__abc_16259_n3322_1), .Y(AES_CORE_DATAPATH__abc_16259_n3323_1) );
  INVX1 INVX1_990 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n140), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_2_) );
  INVX1 INVX1_991 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n102), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n142) );
  INVX1 INVX1_992 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n149), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n150_1) );
  INVX1 INVX1_993 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n157), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n158) );
  INVX1 INVX1_994 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n159) );
  INVX1 INVX1_995 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n161) );
  INVX1 INVX1_996 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n167), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n168) );
  INVX1 INVX1_997 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n173), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n174) );
  INVX1 INVX1_998 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n164), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n175) );
  INVX1 INVX1_999 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n176_1) );
  INVX2 INVX2_1 ( .A(disable_core), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n84_1) );
  INVX2 INVX2_10 ( .A(AES_CORE_DATAPATH__abc_16259_n3204), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_1_) );
  INVX2 INVX2_11 ( .A(AES_CORE_DATAPATH__abc_16259_n3244), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_2_) );
  INVX2 INVX2_12 ( .A(AES_CORE_DATAPATH__abc_16259_n3284), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_3_) );
  INVX2 INVX2_13 ( .A(AES_CORE_DATAPATH__abc_16259_n3364), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_5_) );
  INVX2 INVX2_14 ( .A(AES_CORE_DATAPATH__abc_16259_n3404_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_6_) );
  INVX2 INVX2_15 ( .A(AES_CORE_DATAPATH__abc_16259_n3444_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_7_) );
  INVX2 INVX2_16 ( .A(AES_CORE_DATAPATH__abc_16259_n3484), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_0_) );
  INVX2 INVX2_17 ( .A(AES_CORE_DATAPATH__abc_16259_n3524), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_1_) );
  INVX2 INVX2_18 ( .A(AES_CORE_DATAPATH__abc_16259_n3564_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_2_) );
  INVX2 INVX2_19 ( .A(AES_CORE_DATAPATH__abc_16259_n3604), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_3_) );
  INVX2 INVX2_2 ( .A(AES_CORE_DATAPATH__abc_16259_n2794), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_0_) );
  INVX2 INVX2_20 ( .A(AES_CORE_DATAPATH__abc_16259_n3684), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_5_) );
  INVX2 INVX2_21 ( .A(AES_CORE_DATAPATH__abc_16259_n3724), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_6_) );
  INVX2 INVX2_22 ( .A(AES_CORE_DATAPATH__abc_16259_n3764), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_7_) );
  INVX2 INVX2_23 ( .A(AES_CORE_DATAPATH__abc_16259_n3804), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_0_) );
  INVX2 INVX2_24 ( .A(AES_CORE_DATAPATH__abc_16259_n3844), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_1_) );
  INVX2 INVX2_25 ( .A(AES_CORE_DATAPATH__abc_16259_n3884), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_2_) );
  INVX2 INVX2_26 ( .A(AES_CORE_DATAPATH__abc_16259_n3924), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_3_) );
  INVX2 INVX2_27 ( .A(AES_CORE_DATAPATH__abc_16259_n4004), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_5_) );
  INVX2 INVX2_28 ( .A(AES_CORE_DATAPATH__abc_16259_n4044), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_6_) );
  INVX2 INVX2_29 ( .A(AES_CORE_DATAPATH__abc_16259_n4084), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_7_) );
  INVX2 INVX2_3 ( .A(AES_CORE_DATAPATH__abc_16259_n2883), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_1_) );
  INVX2 INVX2_30 ( .A(AES_CORE_CONTROL_UNIT_mode_cbc_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6091) );
  INVX2 INVX2_31 ( .A(AES_CORE_DATAPATH__abc_16259_n6056_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6556) );
  INVX2 INVX2_32 ( .A(AES_CORE_DATAPATH__abc_16259_n6092_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6586) );
  INVX2 INVX2_33 ( .A(AES_CORE_DATAPATH__abc_16259_n6101_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6595) );
  INVX2 INVX2_34 ( .A(AES_CORE_DATAPATH__abc_16259_n6053_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6600) );
  INVX2 INVX2_35 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out_bF_buf0), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n596) );
  INVX2 INVX2_36 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n106), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n107) );
  INVX2 INVX2_37 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n135) );
  INVX2 INVX2_38 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n160_1) );
  INVX2 INVX2_39 ( .A(AES_CORE_DATAPATH_MIX_COL_col_3__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n175) );
  INVX2 INVX2_4 ( .A(AES_CORE_DATAPATH__abc_16259_n2924_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_2_) );
  INVX2 INVX2_40 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n190) );
  INVX2 INVX2_41 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n195_1) );
  INVX2 INVX2_42 ( .A(AES_CORE_DATAPATH_MIX_COL_col_3__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n230) );
  INVX2 INVX2_43 ( .A(AES_CORE_DATAPATH_MIX_COL_col_3__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n285) );
  INVX2 INVX2_44 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n504), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n510) );
  INVX2 INVX2_45 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n658), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n659) );
  INVX2 INVX2_46 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n678), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n684) );
  INVX2 INVX2_47 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n66_1) );
  INVX2 INVX2_48 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n136), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_1_) );
  INVX2 INVX2_49 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n206), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n212) );
  INVX2 INVX2_5 ( .A(AES_CORE_DATAPATH__abc_16259_n2964), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_3_) );
  INVX2 INVX2_50 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n258), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n317) );
  INVX2 INVX2_51 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n490), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n491) );
  INVX2 INVX2_52 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n66_1) );
  INVX2 INVX2_53 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n136), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_1_) );
  INVX2 INVX2_54 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n206), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n212) );
  INVX2 INVX2_55 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n258), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n317) );
  INVX2 INVX2_56 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n490), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n491) );
  INVX2 INVX2_57 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n66_1) );
  INVX2 INVX2_58 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n136), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_1_) );
  INVX2 INVX2_59 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n206), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n212) );
  INVX2 INVX2_6 ( .A(AES_CORE_DATAPATH__abc_16259_n3044), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_5_) );
  INVX2 INVX2_60 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n258), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n317) );
  INVX2 INVX2_61 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n490), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n491) );
  INVX2 INVX2_62 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n66_1) );
  INVX2 INVX2_63 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n136), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_1_) );
  INVX2 INVX2_64 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n206), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n212) );
  INVX2 INVX2_65 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n258), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n317) );
  INVX2 INVX2_66 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n490), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n491) );
  INVX2 INVX2_7 ( .A(AES_CORE_DATAPATH__abc_16259_n3084), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_6_) );
  INVX2 INVX2_8 ( .A(AES_CORE_DATAPATH__abc_16259_n3124), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_7_) );
  INVX2 INVX2_9 ( .A(AES_CORE_DATAPATH__abc_16259_n3164), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_0_) );
  INVX4 INVX4_1 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n2457_1) );
  INVX4 INVX4_2 ( .A(AES_CORE_CONTROL_UNIT_bypass_key_en), .Y(AES_CORE_DATAPATH__abc_16259_n2806_1) );
  INVX4 INVX4_3 ( .A(AES_CORE_DATAPATH__abc_16259_n3004_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_4_) );
  INVX4 INVX4_4 ( .A(AES_CORE_DATAPATH__abc_16259_n3324), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_4_) );
  INVX4 INVX4_5 ( .A(AES_CORE_DATAPATH__abc_16259_n3644), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_4_) );
  INVX4 INVX4_6 ( .A(AES_CORE_DATAPATH__abc_16259_n3964), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_4_) );
  INVX8 INVX8_1 ( .A(AES_CORE_DATAPATH__abc_16259_n2483_1_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n2484) );
  INVX8 INVX8_10 ( .A(AES_CORE_DATAPATH__abc_16259_n4474_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n4475_1) );
  INVX8 INVX8_11 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf9), .Y(AES_CORE_DATAPATH__abc_16259_n4480_1) );
  INVX8 INVX8_12 ( .A(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf9), .Y(AES_CORE_DATAPATH__abc_16259_n4769) );
  INVX8 INVX8_13 ( .A(key_en_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n4867_1) );
  INVX8 INVX8_14 ( .A(AES_CORE_DATAPATH__abc_16259_n4872_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n4873_1) );
  INVX8 INVX8_15 ( .A(key_en_2_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5260_1) );
  INVX8 INVX8_16 ( .A(AES_CORE_DATAPATH__abc_16259_n5265_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5266_1) );
  INVX8 INVX8_17 ( .A(key_en_3_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5653) );
  INVX8 INVX8_18 ( .A(AES_CORE_DATAPATH__abc_16259_n5658_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5659) );
  INVX8 INVX8_19 ( .A(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6044) );
  INVX8 INVX8_2 ( .A(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n2485_1) );
  INVX8 INVX8_20 ( .A(AES_CORE_CONTROL_UNIT_last_round_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6057) );
  INVX8 INVX8_21 ( .A(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n6059) );
  INVX8 INVX8_22 ( .A(AES_CORE_DATAPATH__abc_16259_n6063_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6074) );
  INVX8 INVX8_23 ( .A(AES_CORE_DATAPATH__abc_16259_n6095_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6097) );
  INVX8 INVX8_24 ( .A(AES_CORE_DATAPATH__abc_16259_n6107_bF_buf9), .Y(AES_CORE_DATAPATH__abc_16259_n6603) );
  INVX8 INVX8_25 ( .A(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7669) );
  INVX8 INVX8_26 ( .A(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7944) );
  INVX8 INVX8_27 ( .A(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n8219) );
  INVX8 INVX8_28 ( .A(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n8500) );
  INVX8 INVX8_29 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf10), .Y(AES_CORE_DATAPATH__abc_16259_n8603) );
  INVX8 INVX8_3 ( .A(AES_CORE_DATAPATH_last_round_pp2_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n2798) );
  INVX8 INVX8_30 ( .A(AES_CORE_DATAPATH__abc_16259_n8898_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n8899) );
  INVX8 INVX8_31 ( .A(AES_CORE_CONTROL_UNIT_iv_cnt_en), .Y(AES_CORE_DATAPATH__abc_16259_n8918) );
  INVX8 INVX8_32 ( .A(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n9288) );
  INVX8 INVX8_33 ( .A(iv_en_2_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n9654) );
  INVX8 INVX8_34 ( .A(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n9753) );
  INVX8 INVX8_35 ( .A(iv_en_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n10119) );
  INVX8 INVX8_36 ( .A(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n10218) );
  INVX8 INVX8_37 ( .A(iv_en_0_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n10584) );
  INVX8 INVX8_38 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf7), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597) );
  INVX8 INVX8_4 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n2802) );
  INVX8 INVX8_5 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n2803) );
  INVX8 INVX8_6 ( .A(AES_CORE_DATAPATH__abc_16259_n2826_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n2841) );
  INVX8 INVX8_7 ( .A(AES_CORE_DATAPATH__abc_16259_n2852), .Y(AES_CORE_DATAPATH__abc_16259_n2853_1) );
  INVX8 INVX8_8 ( .A(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n2864_1) );
  INVX8 INVX8_9 ( .A(key_en_0_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n4468_1) );
  OR2X2 OR2X2_1 ( .A(AES_CORE_CONTROL_UNIT_state_7_), .B(AES_CORE_CONTROL_UNIT_state_11_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n75) );
  OR2X2 OR2X2_10 ( .A(AES_CORE_CONTROL_UNIT_rd_count_2_), .B(AES_CORE_CONTROL_UNIT_rd_count_3_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n110_1) );
  OR2X2 OR2X2_100 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf4), .B(AES_CORE_DATAPATH_iv_2__3_), .Y(AES_CORE_DATAPATH__abc_16259_n2513_1) );
  OR2X2 OR2X2_1000 ( .A(AES_CORE_DATAPATH__abc_16259_n4742), .B(AES_CORE_DATAPATH__abc_16259_n4743), .Y(AES_CORE_DATAPATH__abc_16259_n4744_1) );
  OR2X2 OR2X2_1001 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n4744_1), .Y(AES_CORE_DATAPATH__abc_16259_n4745) );
  OR2X2 OR2X2_1002 ( .A(AES_CORE_DATAPATH__abc_16259_n4747), .B(AES_CORE_DATAPATH__abc_16259_n4748), .Y(AES_CORE_DATAPATH__0key_0__31_0__29_) );
  OR2X2 OR2X2_1003 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_126_), .Y(AES_CORE_DATAPATH__abc_16259_n4750_1) );
  OR2X2 OR2X2_1004 ( .A(AES_CORE_DATAPATH__abc_16259_n4751), .B(AES_CORE_DATAPATH__abc_16259_n4752), .Y(AES_CORE_DATAPATH__abc_16259_n4753) );
  OR2X2 OR2X2_1005 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n4753), .Y(AES_CORE_DATAPATH__abc_16259_n4754) );
  OR2X2 OR2X2_1006 ( .A(AES_CORE_DATAPATH__abc_16259_n4756), .B(AES_CORE_DATAPATH__abc_16259_n4757_1), .Y(AES_CORE_DATAPATH__0key_0__31_0__30_) );
  OR2X2 OR2X2_1007 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_127_), .Y(AES_CORE_DATAPATH__abc_16259_n4759) );
  OR2X2 OR2X2_1008 ( .A(AES_CORE_DATAPATH__abc_16259_n4760), .B(AES_CORE_DATAPATH__abc_16259_n4761), .Y(AES_CORE_DATAPATH__abc_16259_n4762) );
  OR2X2 OR2X2_1009 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n4762), .Y(AES_CORE_DATAPATH__abc_16259_n4763_1) );
  OR2X2 OR2X2_101 ( .A(AES_CORE_DATAPATH__abc_16259_n2515), .B(AES_CORE_DATAPATH__abc_16259_n2516_1), .Y(_auto_iopadmap_cc_313_execute_26916_3_) );
  OR2X2 OR2X2_1010 ( .A(AES_CORE_DATAPATH__abc_16259_n4764), .B(AES_CORE_DATAPATH__abc_16259_n4474_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n4765) );
  OR2X2 OR2X2_1011 ( .A(AES_CORE_DATAPATH__abc_16259_n4475_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__31_), .Y(AES_CORE_DATAPATH__abc_16259_n4766) );
  OR2X2 OR2X2_1012 ( .A(AES_CORE_DATAPATH__abc_16259_n4770), .B(AES_CORE_DATAPATH__abc_16259_n4768), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__0_) );
  OR2X2 OR2X2_1013 ( .A(AES_CORE_DATAPATH__abc_16259_n4492_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf8), .Y(AES_CORE_DATAPATH__abc_16259_n4772_1) );
  OR2X2 OR2X2_1014 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf9), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__1_), .Y(AES_CORE_DATAPATH__abc_16259_n4773) );
  OR2X2 OR2X2_1015 ( .A(AES_CORE_DATAPATH__abc_16259_n4501_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n4775) );
  OR2X2 OR2X2_1016 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf8), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__2_), .Y(AES_CORE_DATAPATH__abc_16259_n4776) );
  OR2X2 OR2X2_1017 ( .A(AES_CORE_DATAPATH__abc_16259_n4510_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n4778_1) );
  OR2X2 OR2X2_1018 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf7), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__3_), .Y(AES_CORE_DATAPATH__abc_16259_n4779) );
  OR2X2 OR2X2_1019 ( .A(AES_CORE_DATAPATH__abc_16259_n4519_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n4781) );
  OR2X2 OR2X2_102 ( .A(AES_CORE_DATAPATH__abc_16259_n2519_1), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n2520) );
  OR2X2 OR2X2_1020 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf6), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__4_), .Y(AES_CORE_DATAPATH__abc_16259_n4782) );
  OR2X2 OR2X2_1021 ( .A(AES_CORE_DATAPATH__abc_16259_n4528_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n4784) );
  OR2X2 OR2X2_1022 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf5), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__5_), .Y(AES_CORE_DATAPATH__abc_16259_n4785_1) );
  OR2X2 OR2X2_1023 ( .A(AES_CORE_DATAPATH__abc_16259_n4537_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n4787) );
  OR2X2 OR2X2_1024 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__6_), .Y(AES_CORE_DATAPATH__abc_16259_n4788) );
  OR2X2 OR2X2_1025 ( .A(AES_CORE_DATAPATH__abc_16259_n4546_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n4790) );
  OR2X2 OR2X2_1026 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__7_), .Y(AES_CORE_DATAPATH__abc_16259_n4791_1) );
  OR2X2 OR2X2_1027 ( .A(AES_CORE_DATAPATH__abc_16259_n4555_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n4793) );
  OR2X2 OR2X2_1028 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__8_), .Y(AES_CORE_DATAPATH__abc_16259_n4794) );
  OR2X2 OR2X2_1029 ( .A(AES_CORE_DATAPATH__abc_16259_n4564_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n4796) );
  OR2X2 OR2X2_103 ( .A(AES_CORE_DATAPATH__abc_16259_n2518_1), .B(AES_CORE_DATAPATH__abc_16259_n2520), .Y(AES_CORE_DATAPATH__abc_16259_n2521_1) );
  OR2X2 OR2X2_1030 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__9_), .Y(AES_CORE_DATAPATH__abc_16259_n4797) );
  OR2X2 OR2X2_1031 ( .A(AES_CORE_DATAPATH__abc_16259_n4573_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf10), .Y(AES_CORE_DATAPATH__abc_16259_n4799_1) );
  OR2X2 OR2X2_1032 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__10_), .Y(AES_CORE_DATAPATH__abc_16259_n4800) );
  OR2X2 OR2X2_1033 ( .A(AES_CORE_DATAPATH__abc_16259_n4582_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf9), .Y(AES_CORE_DATAPATH__abc_16259_n4802) );
  OR2X2 OR2X2_1034 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf10), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__11_), .Y(AES_CORE_DATAPATH__abc_16259_n4803) );
  OR2X2 OR2X2_1035 ( .A(AES_CORE_DATAPATH__abc_16259_n4591_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf8), .Y(AES_CORE_DATAPATH__abc_16259_n4805_1) );
  OR2X2 OR2X2_1036 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf9), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__12_), .Y(AES_CORE_DATAPATH__abc_16259_n4806) );
  OR2X2 OR2X2_1037 ( .A(AES_CORE_DATAPATH__abc_16259_n4600_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n4808) );
  OR2X2 OR2X2_1038 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf8), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__13_), .Y(AES_CORE_DATAPATH__abc_16259_n4809) );
  OR2X2 OR2X2_1039 ( .A(AES_CORE_DATAPATH__abc_16259_n4609), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n4811) );
  OR2X2 OR2X2_104 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf3), .B(AES_CORE_DATAPATH_iv_2__4_), .Y(AES_CORE_DATAPATH__abc_16259_n2522) );
  OR2X2 OR2X2_1040 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf7), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__14_), .Y(AES_CORE_DATAPATH__abc_16259_n4812_1) );
  OR2X2 OR2X2_1041 ( .A(AES_CORE_DATAPATH__abc_16259_n4618), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n4814) );
  OR2X2 OR2X2_1042 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf6), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__15_), .Y(AES_CORE_DATAPATH__abc_16259_n4815) );
  OR2X2 OR2X2_1043 ( .A(AES_CORE_DATAPATH__abc_16259_n4627), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n4817) );
  OR2X2 OR2X2_1044 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf5), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__16_), .Y(AES_CORE_DATAPATH__abc_16259_n4818_1) );
  OR2X2 OR2X2_1045 ( .A(AES_CORE_DATAPATH__abc_16259_n4636), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n4820_1) );
  OR2X2 OR2X2_1046 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__17_), .Y(AES_CORE_DATAPATH__abc_16259_n4821_1) );
  OR2X2 OR2X2_1047 ( .A(AES_CORE_DATAPATH__abc_16259_n4645), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n4823_1) );
  OR2X2 OR2X2_1048 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__18_), .Y(AES_CORE_DATAPATH__abc_16259_n4824_1) );
  OR2X2 OR2X2_1049 ( .A(AES_CORE_DATAPATH__abc_16259_n4654_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n4826_1) );
  OR2X2 OR2X2_105 ( .A(AES_CORE_DATAPATH__abc_16259_n2524_1), .B(AES_CORE_DATAPATH__abc_16259_n2525), .Y(_auto_iopadmap_cc_313_execute_26916_4_) );
  OR2X2 OR2X2_1050 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__19_), .Y(AES_CORE_DATAPATH__abc_16259_n4827_1) );
  OR2X2 OR2X2_1051 ( .A(AES_CORE_DATAPATH__abc_16259_n4663), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n4829_1) );
  OR2X2 OR2X2_1052 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__20_), .Y(AES_CORE_DATAPATH__abc_16259_n4830_1) );
  OR2X2 OR2X2_1053 ( .A(AES_CORE_DATAPATH__abc_16259_n4672), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf10), .Y(AES_CORE_DATAPATH__abc_16259_n4832_1) );
  OR2X2 OR2X2_1054 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__21_), .Y(AES_CORE_DATAPATH__abc_16259_n4833_1) );
  OR2X2 OR2X2_1055 ( .A(AES_CORE_DATAPATH__abc_16259_n4681_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf9), .Y(AES_CORE_DATAPATH__abc_16259_n4835_1) );
  OR2X2 OR2X2_1056 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf10), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__22_), .Y(AES_CORE_DATAPATH__abc_16259_n4836_1) );
  OR2X2 OR2X2_1057 ( .A(AES_CORE_DATAPATH__abc_16259_n4690), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf8), .Y(AES_CORE_DATAPATH__abc_16259_n4838_1) );
  OR2X2 OR2X2_1058 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf9), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__23_), .Y(AES_CORE_DATAPATH__abc_16259_n4839_1) );
  OR2X2 OR2X2_1059 ( .A(AES_CORE_DATAPATH__abc_16259_n4699), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n4841_1) );
  OR2X2 OR2X2_106 ( .A(AES_CORE_DATAPATH__abc_16259_n2528_1), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n2529_1) );
  OR2X2 OR2X2_1060 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf8), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__24_), .Y(AES_CORE_DATAPATH__abc_16259_n4842_1) );
  OR2X2 OR2X2_1061 ( .A(AES_CORE_DATAPATH__abc_16259_n4708_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n4844_1) );
  OR2X2 OR2X2_1062 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf7), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__25_), .Y(AES_CORE_DATAPATH__abc_16259_n4845_1) );
  OR2X2 OR2X2_1063 ( .A(AES_CORE_DATAPATH__abc_16259_n4717_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n4847_1) );
  OR2X2 OR2X2_1064 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf6), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__26_), .Y(AES_CORE_DATAPATH__abc_16259_n4848_1) );
  OR2X2 OR2X2_1065 ( .A(AES_CORE_DATAPATH__abc_16259_n4726), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n4850_1) );
  OR2X2 OR2X2_1066 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf5), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__27_), .Y(AES_CORE_DATAPATH__abc_16259_n4851_1) );
  OR2X2 OR2X2_1067 ( .A(AES_CORE_DATAPATH__abc_16259_n4735), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n4853_1) );
  OR2X2 OR2X2_1068 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__28_), .Y(AES_CORE_DATAPATH__abc_16259_n4854_1) );
  OR2X2 OR2X2_1069 ( .A(AES_CORE_DATAPATH__abc_16259_n4744_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n4856_1) );
  OR2X2 OR2X2_107 ( .A(AES_CORE_DATAPATH__abc_16259_n2527), .B(AES_CORE_DATAPATH__abc_16259_n2529_1), .Y(AES_CORE_DATAPATH__abc_16259_n2530) );
  OR2X2 OR2X2_1070 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__29_), .Y(AES_CORE_DATAPATH__abc_16259_n4857_1) );
  OR2X2 OR2X2_1071 ( .A(AES_CORE_DATAPATH__abc_16259_n4753), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n4859_1) );
  OR2X2 OR2X2_1072 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__30_), .Y(AES_CORE_DATAPATH__abc_16259_n4860_1) );
  OR2X2 OR2X2_1073 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__31_), .Y(AES_CORE_DATAPATH__abc_16259_n4862_1) );
  OR2X2 OR2X2_1074 ( .A(AES_CORE_DATAPATH__abc_16259_n4762), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n4863_1) );
  OR2X2 OR2X2_1075 ( .A(AES_CORE_DATAPATH__abc_16259_n4876_1), .B(AES_CORE_DATAPATH__abc_16259_n4875_1), .Y(AES_CORE_DATAPATH__abc_16259_n4877_1) );
  OR2X2 OR2X2_1076 ( .A(AES_CORE_DATAPATH__abc_16259_n4878_1), .B(AES_CORE_DATAPATH__abc_16259_n4874_1), .Y(AES_CORE_DATAPATH__abc_16259_n4879_1) );
  OR2X2 OR2X2_1077 ( .A(AES_CORE_DATAPATH__abc_16259_n4880_1), .B(AES_CORE_DATAPATH__abc_16259_n4881_1), .Y(AES_CORE_DATAPATH__0key_1__31_0__0_) );
  OR2X2 OR2X2_1078 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf10), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_65_), .Y(AES_CORE_DATAPATH__abc_16259_n4883_1) );
  OR2X2 OR2X2_1079 ( .A(AES_CORE_DATAPATH__abc_16259_n4884), .B(AES_CORE_DATAPATH__abc_16259_n4885), .Y(AES_CORE_DATAPATH__abc_16259_n4886_1) );
  OR2X2 OR2X2_108 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf2), .B(AES_CORE_DATAPATH_iv_2__5_), .Y(AES_CORE_DATAPATH__abc_16259_n2531_1) );
  OR2X2 OR2X2_1080 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf9), .B(AES_CORE_DATAPATH__abc_16259_n4886_1), .Y(AES_CORE_DATAPATH__abc_16259_n4887) );
  OR2X2 OR2X2_1081 ( .A(AES_CORE_DATAPATH__abc_16259_n4889_1), .B(AES_CORE_DATAPATH__abc_16259_n4890), .Y(AES_CORE_DATAPATH__0key_1__31_0__1_) );
  OR2X2 OR2X2_1082 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf9), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_66_), .Y(AES_CORE_DATAPATH__abc_16259_n4892_1) );
  OR2X2 OR2X2_1083 ( .A(AES_CORE_DATAPATH__abc_16259_n4893), .B(AES_CORE_DATAPATH__abc_16259_n4894), .Y(AES_CORE_DATAPATH__abc_16259_n4895_1) );
  OR2X2 OR2X2_1084 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf8), .B(AES_CORE_DATAPATH__abc_16259_n4895_1), .Y(AES_CORE_DATAPATH__abc_16259_n4896) );
  OR2X2 OR2X2_1085 ( .A(AES_CORE_DATAPATH__abc_16259_n4897), .B(AES_CORE_DATAPATH__abc_16259_n4872_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n4898_1) );
  OR2X2 OR2X2_1086 ( .A(AES_CORE_DATAPATH__abc_16259_n4873_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__2_), .Y(AES_CORE_DATAPATH__abc_16259_n4899) );
  OR2X2 OR2X2_1087 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf8), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_67_), .Y(AES_CORE_DATAPATH__abc_16259_n4901_1) );
  OR2X2 OR2X2_1088 ( .A(AES_CORE_DATAPATH__abc_16259_n4902), .B(AES_CORE_DATAPATH__abc_16259_n4903), .Y(AES_CORE_DATAPATH__abc_16259_n4904_1) );
  OR2X2 OR2X2_1089 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf7), .B(AES_CORE_DATAPATH__abc_16259_n4904_1), .Y(AES_CORE_DATAPATH__abc_16259_n4905) );
  OR2X2 OR2X2_109 ( .A(AES_CORE_DATAPATH__abc_16259_n2533_1), .B(AES_CORE_DATAPATH__abc_16259_n2534_1), .Y(_auto_iopadmap_cc_313_execute_26916_5_) );
  OR2X2 OR2X2_1090 ( .A(AES_CORE_DATAPATH__abc_16259_n4907_1), .B(AES_CORE_DATAPATH__abc_16259_n4908), .Y(AES_CORE_DATAPATH__0key_1__31_0__3_) );
  OR2X2 OR2X2_1091 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf7), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_68_), .Y(AES_CORE_DATAPATH__abc_16259_n4910_1) );
  OR2X2 OR2X2_1092 ( .A(AES_CORE_DATAPATH__abc_16259_n4911), .B(AES_CORE_DATAPATH__abc_16259_n4912), .Y(AES_CORE_DATAPATH__abc_16259_n4913_1) );
  OR2X2 OR2X2_1093 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf6), .B(AES_CORE_DATAPATH__abc_16259_n4913_1), .Y(AES_CORE_DATAPATH__abc_16259_n4914) );
  OR2X2 OR2X2_1094 ( .A(AES_CORE_DATAPATH__abc_16259_n4916_1), .B(AES_CORE_DATAPATH__abc_16259_n4917), .Y(AES_CORE_DATAPATH__0key_1__31_0__4_) );
  OR2X2 OR2X2_1095 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf6), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_69_), .Y(AES_CORE_DATAPATH__abc_16259_n4919_1) );
  OR2X2 OR2X2_1096 ( .A(AES_CORE_DATAPATH__abc_16259_n4920), .B(AES_CORE_DATAPATH__abc_16259_n4921), .Y(AES_CORE_DATAPATH__abc_16259_n4922_1) );
  OR2X2 OR2X2_1097 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf5), .B(AES_CORE_DATAPATH__abc_16259_n4922_1), .Y(AES_CORE_DATAPATH__abc_16259_n4923) );
  OR2X2 OR2X2_1098 ( .A(AES_CORE_DATAPATH__abc_16259_n4924), .B(AES_CORE_DATAPATH__abc_16259_n4872_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n4925_1) );
  OR2X2 OR2X2_1099 ( .A(AES_CORE_DATAPATH__abc_16259_n4873_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__5_), .Y(AES_CORE_DATAPATH__abc_16259_n4926) );
  OR2X2 OR2X2_11 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n109_1), .B(AES_CORE_CONTROL_UNIT__abc_15841_n110_1), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n111) );
  OR2X2 OR2X2_110 ( .A(AES_CORE_DATAPATH__abc_16259_n2537), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n2538_1) );
  OR2X2 OR2X2_1100 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf5), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_70_), .Y(AES_CORE_DATAPATH__abc_16259_n4928_1) );
  OR2X2 OR2X2_1101 ( .A(AES_CORE_DATAPATH__abc_16259_n4929), .B(AES_CORE_DATAPATH__abc_16259_n4930), .Y(AES_CORE_DATAPATH__abc_16259_n4931_1) );
  OR2X2 OR2X2_1102 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n4931_1), .Y(AES_CORE_DATAPATH__abc_16259_n4932) );
  OR2X2 OR2X2_1103 ( .A(AES_CORE_DATAPATH__abc_16259_n4933), .B(AES_CORE_DATAPATH__abc_16259_n4872_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n4934_1) );
  OR2X2 OR2X2_1104 ( .A(AES_CORE_DATAPATH__abc_16259_n4873_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__6_), .Y(AES_CORE_DATAPATH__abc_16259_n4935) );
  OR2X2 OR2X2_1105 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_71_), .Y(AES_CORE_DATAPATH__abc_16259_n4937_1) );
  OR2X2 OR2X2_1106 ( .A(AES_CORE_DATAPATH__abc_16259_n4938), .B(AES_CORE_DATAPATH__abc_16259_n4939), .Y(AES_CORE_DATAPATH__abc_16259_n4940_1) );
  OR2X2 OR2X2_1107 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n4940_1), .Y(AES_CORE_DATAPATH__abc_16259_n4941) );
  OR2X2 OR2X2_1108 ( .A(AES_CORE_DATAPATH__abc_16259_n4943_1), .B(AES_CORE_DATAPATH__abc_16259_n4944), .Y(AES_CORE_DATAPATH__0key_1__31_0__7_) );
  OR2X2 OR2X2_1109 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_72_), .Y(AES_CORE_DATAPATH__abc_16259_n4946_1) );
  OR2X2 OR2X2_111 ( .A(AES_CORE_DATAPATH__abc_16259_n2536_1), .B(AES_CORE_DATAPATH__abc_16259_n2538_1), .Y(AES_CORE_DATAPATH__abc_16259_n2539_1) );
  OR2X2 OR2X2_1110 ( .A(AES_CORE_DATAPATH__abc_16259_n4947), .B(AES_CORE_DATAPATH__abc_16259_n4948), .Y(AES_CORE_DATAPATH__abc_16259_n4949_1) );
  OR2X2 OR2X2_1111 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n4949_1), .Y(AES_CORE_DATAPATH__abc_16259_n4950) );
  OR2X2 OR2X2_1112 ( .A(AES_CORE_DATAPATH__abc_16259_n4952_1), .B(AES_CORE_DATAPATH__abc_16259_n4953), .Y(AES_CORE_DATAPATH__0key_1__31_0__8_) );
  OR2X2 OR2X2_1113 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_73_), .Y(AES_CORE_DATAPATH__abc_16259_n4955_1) );
  OR2X2 OR2X2_1114 ( .A(AES_CORE_DATAPATH__abc_16259_n4956), .B(AES_CORE_DATAPATH__abc_16259_n4957), .Y(AES_CORE_DATAPATH__abc_16259_n4958_1) );
  OR2X2 OR2X2_1115 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n4958_1), .Y(AES_CORE_DATAPATH__abc_16259_n4959) );
  OR2X2 OR2X2_1116 ( .A(AES_CORE_DATAPATH__abc_16259_n4961_1), .B(AES_CORE_DATAPATH__abc_16259_n4962), .Y(AES_CORE_DATAPATH__0key_1__31_0__9_) );
  OR2X2 OR2X2_1117 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_74_), .Y(AES_CORE_DATAPATH__abc_16259_n4964_1) );
  OR2X2 OR2X2_1118 ( .A(AES_CORE_DATAPATH__abc_16259_n4965), .B(AES_CORE_DATAPATH__abc_16259_n4966), .Y(AES_CORE_DATAPATH__abc_16259_n4967_1) );
  OR2X2 OR2X2_1119 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n4967_1), .Y(AES_CORE_DATAPATH__abc_16259_n4968) );
  OR2X2 OR2X2_112 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf1), .B(AES_CORE_DATAPATH_iv_2__6_), .Y(AES_CORE_DATAPATH__abc_16259_n2540) );
  OR2X2 OR2X2_1120 ( .A(AES_CORE_DATAPATH__abc_16259_n4969), .B(AES_CORE_DATAPATH__abc_16259_n4872_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n4970_1) );
  OR2X2 OR2X2_1121 ( .A(AES_CORE_DATAPATH__abc_16259_n4873_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__10_), .Y(AES_CORE_DATAPATH__abc_16259_n4971) );
  OR2X2 OR2X2_1122 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_75_), .Y(AES_CORE_DATAPATH__abc_16259_n4973_1) );
  OR2X2 OR2X2_1123 ( .A(AES_CORE_DATAPATH__abc_16259_n4974), .B(AES_CORE_DATAPATH__abc_16259_n4975), .Y(AES_CORE_DATAPATH__abc_16259_n4976_1) );
  OR2X2 OR2X2_1124 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf10), .B(AES_CORE_DATAPATH__abc_16259_n4976_1), .Y(AES_CORE_DATAPATH__abc_16259_n4977) );
  OR2X2 OR2X2_1125 ( .A(AES_CORE_DATAPATH__abc_16259_n4979_1), .B(AES_CORE_DATAPATH__abc_16259_n4980_1), .Y(AES_CORE_DATAPATH__0key_1__31_0__11_) );
  OR2X2 OR2X2_1126 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf10), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_76_), .Y(AES_CORE_DATAPATH__abc_16259_n4982_1) );
  OR2X2 OR2X2_1127 ( .A(AES_CORE_DATAPATH__abc_16259_n4983_1), .B(AES_CORE_DATAPATH__abc_16259_n4984_1), .Y(AES_CORE_DATAPATH__abc_16259_n4985_1) );
  OR2X2 OR2X2_1128 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf9), .B(AES_CORE_DATAPATH__abc_16259_n4985_1), .Y(AES_CORE_DATAPATH__abc_16259_n4986_1) );
  OR2X2 OR2X2_1129 ( .A(AES_CORE_DATAPATH__abc_16259_n4988_1), .B(AES_CORE_DATAPATH__abc_16259_n4989_1), .Y(AES_CORE_DATAPATH__0key_1__31_0__12_) );
  OR2X2 OR2X2_113 ( .A(AES_CORE_DATAPATH__abc_16259_n2542), .B(AES_CORE_DATAPATH__abc_16259_n2543_1), .Y(_auto_iopadmap_cc_313_execute_26916_6_) );
  OR2X2 OR2X2_1130 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf9), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_77_), .Y(AES_CORE_DATAPATH__abc_16259_n4991_1) );
  OR2X2 OR2X2_1131 ( .A(AES_CORE_DATAPATH__abc_16259_n4992_1), .B(AES_CORE_DATAPATH__abc_16259_n4993_1), .Y(AES_CORE_DATAPATH__abc_16259_n4994_1) );
  OR2X2 OR2X2_1132 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf8), .B(AES_CORE_DATAPATH__abc_16259_n4994_1), .Y(AES_CORE_DATAPATH__abc_16259_n4995_1) );
  OR2X2 OR2X2_1133 ( .A(AES_CORE_DATAPATH__abc_16259_n4996_1), .B(AES_CORE_DATAPATH__abc_16259_n4872_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n4997_1) );
  OR2X2 OR2X2_1134 ( .A(AES_CORE_DATAPATH__abc_16259_n4873_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__13_), .Y(AES_CORE_DATAPATH__abc_16259_n4998_1) );
  OR2X2 OR2X2_1135 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf8), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_78_), .Y(AES_CORE_DATAPATH__abc_16259_n5000_1) );
  OR2X2 OR2X2_1136 ( .A(AES_CORE_DATAPATH__abc_16259_n5001_1), .B(AES_CORE_DATAPATH__abc_16259_n5002_1), .Y(AES_CORE_DATAPATH__abc_16259_n5003_1) );
  OR2X2 OR2X2_1137 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf7), .B(AES_CORE_DATAPATH__abc_16259_n5003_1), .Y(AES_CORE_DATAPATH__abc_16259_n5004_1) );
  OR2X2 OR2X2_1138 ( .A(AES_CORE_DATAPATH__abc_16259_n5006_1), .B(AES_CORE_DATAPATH__abc_16259_n5007_1), .Y(AES_CORE_DATAPATH__0key_1__31_0__14_) );
  OR2X2 OR2X2_1139 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf7), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_79_), .Y(AES_CORE_DATAPATH__abc_16259_n5009_1) );
  OR2X2 OR2X2_114 ( .A(AES_CORE_DATAPATH__abc_16259_n2546_1), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n2547) );
  OR2X2 OR2X2_1140 ( .A(AES_CORE_DATAPATH__abc_16259_n5010_1), .B(AES_CORE_DATAPATH__abc_16259_n5011_1), .Y(AES_CORE_DATAPATH__abc_16259_n5012_1) );
  OR2X2 OR2X2_1141 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf6), .B(AES_CORE_DATAPATH__abc_16259_n5012_1), .Y(AES_CORE_DATAPATH__abc_16259_n5013) );
  OR2X2 OR2X2_1142 ( .A(AES_CORE_DATAPATH__abc_16259_n5015_1), .B(AES_CORE_DATAPATH__abc_16259_n5016_1), .Y(AES_CORE_DATAPATH__0key_1__31_0__15_) );
  OR2X2 OR2X2_1143 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf6), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_80_), .Y(AES_CORE_DATAPATH__abc_16259_n5018_1) );
  OR2X2 OR2X2_1144 ( .A(AES_CORE_DATAPATH__abc_16259_n5019_1), .B(AES_CORE_DATAPATH__abc_16259_n5020_1), .Y(AES_CORE_DATAPATH__abc_16259_n5021_1) );
  OR2X2 OR2X2_1145 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf5), .B(AES_CORE_DATAPATH__abc_16259_n5021_1), .Y(AES_CORE_DATAPATH__abc_16259_n5022_1) );
  OR2X2 OR2X2_1146 ( .A(AES_CORE_DATAPATH__abc_16259_n5024_1), .B(AES_CORE_DATAPATH__abc_16259_n5025_1), .Y(AES_CORE_DATAPATH__0key_1__31_0__16_) );
  OR2X2 OR2X2_1147 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf5), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_81_), .Y(AES_CORE_DATAPATH__abc_16259_n5027_1) );
  OR2X2 OR2X2_1148 ( .A(AES_CORE_DATAPATH__abc_16259_n5028_1), .B(AES_CORE_DATAPATH__abc_16259_n5029_1), .Y(AES_CORE_DATAPATH__abc_16259_n5030_1) );
  OR2X2 OR2X2_1149 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n5030_1), .Y(AES_CORE_DATAPATH__abc_16259_n5031_1) );
  OR2X2 OR2X2_115 ( .A(AES_CORE_DATAPATH__abc_16259_n2545), .B(AES_CORE_DATAPATH__abc_16259_n2547), .Y(AES_CORE_DATAPATH__abc_16259_n2548_1) );
  OR2X2 OR2X2_1150 ( .A(AES_CORE_DATAPATH__abc_16259_n5032_1), .B(AES_CORE_DATAPATH__abc_16259_n4872_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n5033_1) );
  OR2X2 OR2X2_1151 ( .A(AES_CORE_DATAPATH__abc_16259_n4873_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__17_), .Y(AES_CORE_DATAPATH__abc_16259_n5034_1) );
  OR2X2 OR2X2_1152 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_82_), .Y(AES_CORE_DATAPATH__abc_16259_n5036_1) );
  OR2X2 OR2X2_1153 ( .A(AES_CORE_DATAPATH__abc_16259_n5037_1), .B(AES_CORE_DATAPATH__abc_16259_n5038_1), .Y(AES_CORE_DATAPATH__abc_16259_n5039_1) );
  OR2X2 OR2X2_1154 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n5039_1), .Y(AES_CORE_DATAPATH__abc_16259_n5040_1) );
  OR2X2 OR2X2_1155 ( .A(AES_CORE_DATAPATH__abc_16259_n5042_1), .B(AES_CORE_DATAPATH__abc_16259_n5043_1), .Y(AES_CORE_DATAPATH__0key_1__31_0__18_) );
  OR2X2 OR2X2_1156 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_83_), .Y(AES_CORE_DATAPATH__abc_16259_n5045_1) );
  OR2X2 OR2X2_1157 ( .A(AES_CORE_DATAPATH__abc_16259_n5046_1), .B(AES_CORE_DATAPATH__abc_16259_n5047_1), .Y(AES_CORE_DATAPATH__abc_16259_n5048_1) );
  OR2X2 OR2X2_1158 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n5048_1), .Y(AES_CORE_DATAPATH__abc_16259_n5049_1) );
  OR2X2 OR2X2_1159 ( .A(AES_CORE_DATAPATH__abc_16259_n5050_1), .B(AES_CORE_DATAPATH__abc_16259_n4872_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5051_1) );
  OR2X2 OR2X2_116 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf0), .B(AES_CORE_DATAPATH_iv_2__7_), .Y(AES_CORE_DATAPATH__abc_16259_n2549_1) );
  OR2X2 OR2X2_1160 ( .A(AES_CORE_DATAPATH__abc_16259_n4873_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__19_), .Y(AES_CORE_DATAPATH__abc_16259_n5052_1) );
  OR2X2 OR2X2_1161 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_84_), .Y(AES_CORE_DATAPATH__abc_16259_n5054_1) );
  OR2X2 OR2X2_1162 ( .A(AES_CORE_DATAPATH__abc_16259_n5055_1), .B(AES_CORE_DATAPATH__abc_16259_n5056_1), .Y(AES_CORE_DATAPATH__abc_16259_n5057_1) );
  OR2X2 OR2X2_1163 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n5057_1), .Y(AES_CORE_DATAPATH__abc_16259_n5058_1) );
  OR2X2 OR2X2_1164 ( .A(AES_CORE_DATAPATH__abc_16259_n5060_1), .B(AES_CORE_DATAPATH__abc_16259_n5061_1), .Y(AES_CORE_DATAPATH__0key_1__31_0__20_) );
  OR2X2 OR2X2_1165 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_85_), .Y(AES_CORE_DATAPATH__abc_16259_n5063_1) );
  OR2X2 OR2X2_1166 ( .A(AES_CORE_DATAPATH__abc_16259_n5064_1), .B(AES_CORE_DATAPATH__abc_16259_n5065_1), .Y(AES_CORE_DATAPATH__abc_16259_n5066_1) );
  OR2X2 OR2X2_1167 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n5066_1), .Y(AES_CORE_DATAPATH__abc_16259_n5067_1) );
  OR2X2 OR2X2_1168 ( .A(AES_CORE_DATAPATH__abc_16259_n5068_1), .B(AES_CORE_DATAPATH__abc_16259_n4872_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n5069_1) );
  OR2X2 OR2X2_1169 ( .A(AES_CORE_DATAPATH__abc_16259_n4873_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__21_), .Y(AES_CORE_DATAPATH__abc_16259_n5070_1) );
  OR2X2 OR2X2_117 ( .A(AES_CORE_DATAPATH__abc_16259_n2551_1), .B(AES_CORE_DATAPATH__abc_16259_n2552), .Y(_auto_iopadmap_cc_313_execute_26916_7_) );
  OR2X2 OR2X2_1170 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_86_), .Y(AES_CORE_DATAPATH__abc_16259_n5072_1) );
  OR2X2 OR2X2_1171 ( .A(AES_CORE_DATAPATH__abc_16259_n5073_1), .B(AES_CORE_DATAPATH__abc_16259_n5074_1), .Y(AES_CORE_DATAPATH__abc_16259_n5075_1) );
  OR2X2 OR2X2_1172 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf10), .B(AES_CORE_DATAPATH__abc_16259_n5075_1), .Y(AES_CORE_DATAPATH__abc_16259_n5076_1) );
  OR2X2 OR2X2_1173 ( .A(AES_CORE_DATAPATH__abc_16259_n5077_1), .B(AES_CORE_DATAPATH__abc_16259_n4872_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n5078) );
  OR2X2 OR2X2_1174 ( .A(AES_CORE_DATAPATH__abc_16259_n4873_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__22_), .Y(AES_CORE_DATAPATH__abc_16259_n5079) );
  OR2X2 OR2X2_1175 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf10), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_87_), .Y(AES_CORE_DATAPATH__abc_16259_n5081) );
  OR2X2 OR2X2_1176 ( .A(AES_CORE_DATAPATH__abc_16259_n5082), .B(AES_CORE_DATAPATH__abc_16259_n5083_1), .Y(AES_CORE_DATAPATH__abc_16259_n5084) );
  OR2X2 OR2X2_1177 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf9), .B(AES_CORE_DATAPATH__abc_16259_n5084), .Y(AES_CORE_DATAPATH__abc_16259_n5085) );
  OR2X2 OR2X2_1178 ( .A(AES_CORE_DATAPATH__abc_16259_n5087), .B(AES_CORE_DATAPATH__abc_16259_n5088), .Y(AES_CORE_DATAPATH__0key_1__31_0__23_) );
  OR2X2 OR2X2_1179 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf9), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_88_), .Y(AES_CORE_DATAPATH__abc_16259_n5090) );
  OR2X2 OR2X2_118 ( .A(AES_CORE_DATAPATH__abc_16259_n2555), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n2556_1) );
  OR2X2 OR2X2_1180 ( .A(AES_CORE_DATAPATH__abc_16259_n5091), .B(AES_CORE_DATAPATH__abc_16259_n5092_1), .Y(AES_CORE_DATAPATH__abc_16259_n5093) );
  OR2X2 OR2X2_1181 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf8), .B(AES_CORE_DATAPATH__abc_16259_n5093), .Y(AES_CORE_DATAPATH__abc_16259_n5094) );
  OR2X2 OR2X2_1182 ( .A(AES_CORE_DATAPATH__abc_16259_n5095_1), .B(AES_CORE_DATAPATH__abc_16259_n4872_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5096) );
  OR2X2 OR2X2_1183 ( .A(AES_CORE_DATAPATH__abc_16259_n4873_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__24_), .Y(AES_CORE_DATAPATH__abc_16259_n5097) );
  OR2X2 OR2X2_1184 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf8), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_89_), .Y(AES_CORE_DATAPATH__abc_16259_n5099) );
  OR2X2 OR2X2_1185 ( .A(AES_CORE_DATAPATH__abc_16259_n5100), .B(AES_CORE_DATAPATH__abc_16259_n5101_1), .Y(AES_CORE_DATAPATH__abc_16259_n5102) );
  OR2X2 OR2X2_1186 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf7), .B(AES_CORE_DATAPATH__abc_16259_n5102), .Y(AES_CORE_DATAPATH__abc_16259_n5103) );
  OR2X2 OR2X2_1187 ( .A(AES_CORE_DATAPATH__abc_16259_n5105), .B(AES_CORE_DATAPATH__abc_16259_n5106), .Y(AES_CORE_DATAPATH__0key_1__31_0__25_) );
  OR2X2 OR2X2_1188 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf7), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_90_), .Y(AES_CORE_DATAPATH__abc_16259_n5108) );
  OR2X2 OR2X2_1189 ( .A(AES_CORE_DATAPATH__abc_16259_n5109), .B(AES_CORE_DATAPATH__abc_16259_n5110_1), .Y(AES_CORE_DATAPATH__abc_16259_n5111) );
  OR2X2 OR2X2_119 ( .A(AES_CORE_DATAPATH__abc_16259_n2554_1), .B(AES_CORE_DATAPATH__abc_16259_n2556_1), .Y(AES_CORE_DATAPATH__abc_16259_n2557) );
  OR2X2 OR2X2_1190 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf6), .B(AES_CORE_DATAPATH__abc_16259_n5111), .Y(AES_CORE_DATAPATH__abc_16259_n5112) );
  OR2X2 OR2X2_1191 ( .A(AES_CORE_DATAPATH__abc_16259_n5113_1), .B(AES_CORE_DATAPATH__abc_16259_n4872_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n5114) );
  OR2X2 OR2X2_1192 ( .A(AES_CORE_DATAPATH__abc_16259_n4873_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__26_), .Y(AES_CORE_DATAPATH__abc_16259_n5115) );
  OR2X2 OR2X2_1193 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf6), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_91_), .Y(AES_CORE_DATAPATH__abc_16259_n5117) );
  OR2X2 OR2X2_1194 ( .A(AES_CORE_DATAPATH__abc_16259_n5118), .B(AES_CORE_DATAPATH__abc_16259_n5119_1), .Y(AES_CORE_DATAPATH__abc_16259_n5120) );
  OR2X2 OR2X2_1195 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf5), .B(AES_CORE_DATAPATH__abc_16259_n5120), .Y(AES_CORE_DATAPATH__abc_16259_n5121) );
  OR2X2 OR2X2_1196 ( .A(AES_CORE_DATAPATH__abc_16259_n5123), .B(AES_CORE_DATAPATH__abc_16259_n5124), .Y(AES_CORE_DATAPATH__0key_1__31_0__27_) );
  OR2X2 OR2X2_1197 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf5), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_92_), .Y(AES_CORE_DATAPATH__abc_16259_n5126) );
  OR2X2 OR2X2_1198 ( .A(AES_CORE_DATAPATH__abc_16259_n5127), .B(AES_CORE_DATAPATH__abc_16259_n5128_1), .Y(AES_CORE_DATAPATH__abc_16259_n5129) );
  OR2X2 OR2X2_1199 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n5129), .Y(AES_CORE_DATAPATH__abc_16259_n5130) );
  OR2X2 OR2X2_12 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n113), .B(AES_CORE_CONTROL_UNIT_state_15_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n114_1) );
  OR2X2 OR2X2_120 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf7), .B(AES_CORE_DATAPATH_iv_2__8_), .Y(AES_CORE_DATAPATH__abc_16259_n2558_1) );
  OR2X2 OR2X2_1200 ( .A(AES_CORE_DATAPATH__abc_16259_n5131_1), .B(AES_CORE_DATAPATH__abc_16259_n4872_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n5132) );
  OR2X2 OR2X2_1201 ( .A(AES_CORE_DATAPATH__abc_16259_n4873_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__28_), .Y(AES_CORE_DATAPATH__abc_16259_n5133) );
  OR2X2 OR2X2_1202 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_93_), .Y(AES_CORE_DATAPATH__abc_16259_n5135) );
  OR2X2 OR2X2_1203 ( .A(AES_CORE_DATAPATH__abc_16259_n5136), .B(AES_CORE_DATAPATH__abc_16259_n5137_1), .Y(AES_CORE_DATAPATH__abc_16259_n5138) );
  OR2X2 OR2X2_1204 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n5138), .Y(AES_CORE_DATAPATH__abc_16259_n5139) );
  OR2X2 OR2X2_1205 ( .A(AES_CORE_DATAPATH__abc_16259_n5140_1), .B(AES_CORE_DATAPATH__abc_16259_n4872_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5141) );
  OR2X2 OR2X2_1206 ( .A(AES_CORE_DATAPATH__abc_16259_n4873_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__29_), .Y(AES_CORE_DATAPATH__abc_16259_n5142) );
  OR2X2 OR2X2_1207 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_94_), .Y(AES_CORE_DATAPATH__abc_16259_n5144) );
  OR2X2 OR2X2_1208 ( .A(AES_CORE_DATAPATH__abc_16259_n5145), .B(AES_CORE_DATAPATH__abc_16259_n5146_1), .Y(AES_CORE_DATAPATH__abc_16259_n5147) );
  OR2X2 OR2X2_1209 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n5147), .Y(AES_CORE_DATAPATH__abc_16259_n5148) );
  OR2X2 OR2X2_121 ( .A(AES_CORE_DATAPATH__abc_16259_n2560), .B(AES_CORE_DATAPATH__abc_16259_n2561_1), .Y(_auto_iopadmap_cc_313_execute_26916_8_) );
  OR2X2 OR2X2_1210 ( .A(AES_CORE_DATAPATH__abc_16259_n5149_1), .B(AES_CORE_DATAPATH__abc_16259_n4872_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n5150) );
  OR2X2 OR2X2_1211 ( .A(AES_CORE_DATAPATH__abc_16259_n4873_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__30_), .Y(AES_CORE_DATAPATH__abc_16259_n5151) );
  OR2X2 OR2X2_1212 ( .A(AES_CORE_DATAPATH__abc_16259_n5153), .B(AES_CORE_DATAPATH__abc_16259_n5154), .Y(AES_CORE_DATAPATH__abc_16259_n5155_1) );
  OR2X2 OR2X2_1213 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n5155_1), .Y(AES_CORE_DATAPATH__abc_16259_n5156) );
  OR2X2 OR2X2_1214 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_95_), .Y(AES_CORE_DATAPATH__abc_16259_n5157) );
  OR2X2 OR2X2_1215 ( .A(AES_CORE_DATAPATH__abc_16259_n5159), .B(AES_CORE_DATAPATH__abc_16259_n5160), .Y(AES_CORE_DATAPATH__0key_1__31_0__31_) );
  OR2X2 OR2X2_1216 ( .A(AES_CORE_DATAPATH__abc_16259_n5163), .B(AES_CORE_DATAPATH__abc_16259_n5162), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__0_) );
  OR2X2 OR2X2_1217 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf10), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__1_), .Y(AES_CORE_DATAPATH__abc_16259_n5165) );
  OR2X2 OR2X2_1218 ( .A(AES_CORE_DATAPATH__abc_16259_n4886_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf9), .Y(AES_CORE_DATAPATH__abc_16259_n5166) );
  OR2X2 OR2X2_1219 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf9), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__2_), .Y(AES_CORE_DATAPATH__abc_16259_n5168) );
  OR2X2 OR2X2_122 ( .A(AES_CORE_DATAPATH__abc_16259_n2564_1), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n2565) );
  OR2X2 OR2X2_1220 ( .A(AES_CORE_DATAPATH__abc_16259_n4895_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf8), .Y(AES_CORE_DATAPATH__abc_16259_n5169) );
  OR2X2 OR2X2_1221 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf8), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__3_), .Y(AES_CORE_DATAPATH__abc_16259_n5171) );
  OR2X2 OR2X2_1222 ( .A(AES_CORE_DATAPATH__abc_16259_n4904_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n5172) );
  OR2X2 OR2X2_1223 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf7), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__4_), .Y(AES_CORE_DATAPATH__abc_16259_n5174_1) );
  OR2X2 OR2X2_1224 ( .A(AES_CORE_DATAPATH__abc_16259_n4913_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n5175_1) );
  OR2X2 OR2X2_1225 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf6), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__5_), .Y(AES_CORE_DATAPATH__abc_16259_n5177_1) );
  OR2X2 OR2X2_1226 ( .A(AES_CORE_DATAPATH__abc_16259_n4922_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n5178_1) );
  OR2X2 OR2X2_1227 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf5), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__6_), .Y(AES_CORE_DATAPATH__abc_16259_n5180_1) );
  OR2X2 OR2X2_1228 ( .A(AES_CORE_DATAPATH__abc_16259_n4931_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5181_1) );
  OR2X2 OR2X2_1229 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__7_), .Y(AES_CORE_DATAPATH__abc_16259_n5183_1) );
  OR2X2 OR2X2_123 ( .A(AES_CORE_DATAPATH__abc_16259_n2563_1), .B(AES_CORE_DATAPATH__abc_16259_n2565), .Y(AES_CORE_DATAPATH__abc_16259_n2566_1) );
  OR2X2 OR2X2_1230 ( .A(AES_CORE_DATAPATH__abc_16259_n4940_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n5184_1) );
  OR2X2 OR2X2_1231 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__8_), .Y(AES_CORE_DATAPATH__abc_16259_n5186_1) );
  OR2X2 OR2X2_1232 ( .A(AES_CORE_DATAPATH__abc_16259_n4949_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n5187_1) );
  OR2X2 OR2X2_1233 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__9_), .Y(AES_CORE_DATAPATH__abc_16259_n5189_1) );
  OR2X2 OR2X2_1234 ( .A(AES_CORE_DATAPATH__abc_16259_n4958_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n5190_1) );
  OR2X2 OR2X2_1235 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__10_), .Y(AES_CORE_DATAPATH__abc_16259_n5192_1) );
  OR2X2 OR2X2_1236 ( .A(AES_CORE_DATAPATH__abc_16259_n4967_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n5193_1) );
  OR2X2 OR2X2_1237 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__11_), .Y(AES_CORE_DATAPATH__abc_16259_n5195_1) );
  OR2X2 OR2X2_1238 ( .A(AES_CORE_DATAPATH__abc_16259_n4976_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf10), .Y(AES_CORE_DATAPATH__abc_16259_n5196_1) );
  OR2X2 OR2X2_1239 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf10), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__12_), .Y(AES_CORE_DATAPATH__abc_16259_n5198_1) );
  OR2X2 OR2X2_124 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf6), .B(AES_CORE_DATAPATH_iv_2__9_), .Y(AES_CORE_DATAPATH__abc_16259_n2567) );
  OR2X2 OR2X2_1240 ( .A(AES_CORE_DATAPATH__abc_16259_n4985_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf9), .Y(AES_CORE_DATAPATH__abc_16259_n5199_1) );
  OR2X2 OR2X2_1241 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf9), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__13_), .Y(AES_CORE_DATAPATH__abc_16259_n5201_1) );
  OR2X2 OR2X2_1242 ( .A(AES_CORE_DATAPATH__abc_16259_n4994_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf8), .Y(AES_CORE_DATAPATH__abc_16259_n5202_1) );
  OR2X2 OR2X2_1243 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf8), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__14_), .Y(AES_CORE_DATAPATH__abc_16259_n5204_1) );
  OR2X2 OR2X2_1244 ( .A(AES_CORE_DATAPATH__abc_16259_n5003_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n5205_1) );
  OR2X2 OR2X2_1245 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf7), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__15_), .Y(AES_CORE_DATAPATH__abc_16259_n5207) );
  OR2X2 OR2X2_1246 ( .A(AES_CORE_DATAPATH__abc_16259_n5012_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n5208_1) );
  OR2X2 OR2X2_1247 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf6), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__16_), .Y(AES_CORE_DATAPATH__abc_16259_n5210_1) );
  OR2X2 OR2X2_1248 ( .A(AES_CORE_DATAPATH__abc_16259_n5021_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n5211_1) );
  OR2X2 OR2X2_1249 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf5), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__17_), .Y(AES_CORE_DATAPATH__abc_16259_n5213_1) );
  OR2X2 OR2X2_125 ( .A(AES_CORE_DATAPATH__abc_16259_n2569_1), .B(AES_CORE_DATAPATH__abc_16259_n2570), .Y(_auto_iopadmap_cc_313_execute_26916_9_) );
  OR2X2 OR2X2_1250 ( .A(AES_CORE_DATAPATH__abc_16259_n5030_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5214_1) );
  OR2X2 OR2X2_1251 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__18_), .Y(AES_CORE_DATAPATH__abc_16259_n5216_1) );
  OR2X2 OR2X2_1252 ( .A(AES_CORE_DATAPATH__abc_16259_n5039_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n5217_1) );
  OR2X2 OR2X2_1253 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__19_), .Y(AES_CORE_DATAPATH__abc_16259_n5219_1) );
  OR2X2 OR2X2_1254 ( .A(AES_CORE_DATAPATH__abc_16259_n5048_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n5220_1) );
  OR2X2 OR2X2_1255 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__20_), .Y(AES_CORE_DATAPATH__abc_16259_n5222_1) );
  OR2X2 OR2X2_1256 ( .A(AES_CORE_DATAPATH__abc_16259_n5057_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n5223_1) );
  OR2X2 OR2X2_1257 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__21_), .Y(AES_CORE_DATAPATH__abc_16259_n5225_1) );
  OR2X2 OR2X2_1258 ( .A(AES_CORE_DATAPATH__abc_16259_n5066_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n5226_1) );
  OR2X2 OR2X2_1259 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__22_), .Y(AES_CORE_DATAPATH__abc_16259_n5228_1) );
  OR2X2 OR2X2_126 ( .A(AES_CORE_DATAPATH__abc_16259_n2573_1), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n2574_1) );
  OR2X2 OR2X2_1260 ( .A(AES_CORE_DATAPATH__abc_16259_n5075_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf10), .Y(AES_CORE_DATAPATH__abc_16259_n5229_1) );
  OR2X2 OR2X2_1261 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf10), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__23_), .Y(AES_CORE_DATAPATH__abc_16259_n5231_1) );
  OR2X2 OR2X2_1262 ( .A(AES_CORE_DATAPATH__abc_16259_n5084), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf9), .Y(AES_CORE_DATAPATH__abc_16259_n5232_1) );
  OR2X2 OR2X2_1263 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf9), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__24_), .Y(AES_CORE_DATAPATH__abc_16259_n5234_1) );
  OR2X2 OR2X2_1264 ( .A(AES_CORE_DATAPATH__abc_16259_n5093), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf8), .Y(AES_CORE_DATAPATH__abc_16259_n5235_1) );
  OR2X2 OR2X2_1265 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf8), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__25_), .Y(AES_CORE_DATAPATH__abc_16259_n5237_1) );
  OR2X2 OR2X2_1266 ( .A(AES_CORE_DATAPATH__abc_16259_n5102), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n5238_1) );
  OR2X2 OR2X2_1267 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf7), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__26_), .Y(AES_CORE_DATAPATH__abc_16259_n5240_1) );
  OR2X2 OR2X2_1268 ( .A(AES_CORE_DATAPATH__abc_16259_n5111), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n5241_1) );
  OR2X2 OR2X2_1269 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf6), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__27_), .Y(AES_CORE_DATAPATH__abc_16259_n5243_1) );
  OR2X2 OR2X2_127 ( .A(AES_CORE_DATAPATH__abc_16259_n2572), .B(AES_CORE_DATAPATH__abc_16259_n2574_1), .Y(AES_CORE_DATAPATH__abc_16259_n2575) );
  OR2X2 OR2X2_1270 ( .A(AES_CORE_DATAPATH__abc_16259_n5120), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n5244_1) );
  OR2X2 OR2X2_1271 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf5), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__28_), .Y(AES_CORE_DATAPATH__abc_16259_n5246_1) );
  OR2X2 OR2X2_1272 ( .A(AES_CORE_DATAPATH__abc_16259_n5129), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5247_1) );
  OR2X2 OR2X2_1273 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__29_), .Y(AES_CORE_DATAPATH__abc_16259_n5249_1) );
  OR2X2 OR2X2_1274 ( .A(AES_CORE_DATAPATH__abc_16259_n5138), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n5250_1) );
  OR2X2 OR2X2_1275 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__30_), .Y(AES_CORE_DATAPATH__abc_16259_n5252_1) );
  OR2X2 OR2X2_1276 ( .A(AES_CORE_DATAPATH__abc_16259_n5147), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n5253_1) );
  OR2X2 OR2X2_1277 ( .A(AES_CORE_DATAPATH__abc_16259_n5155_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n5255_1) );
  OR2X2 OR2X2_1278 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__31_), .Y(AES_CORE_DATAPATH__abc_16259_n5256_1) );
  OR2X2 OR2X2_1279 ( .A(AES_CORE_DATAPATH__abc_16259_n5269_1), .B(AES_CORE_DATAPATH__abc_16259_n5268_1), .Y(AES_CORE_DATAPATH__abc_16259_n5270_1) );
  OR2X2 OR2X2_128 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf5), .B(AES_CORE_DATAPATH_iv_2__10_), .Y(AES_CORE_DATAPATH__abc_16259_n2576_1) );
  OR2X2 OR2X2_1280 ( .A(AES_CORE_DATAPATH__abc_16259_n5271_1), .B(AES_CORE_DATAPATH__abc_16259_n5267_1), .Y(AES_CORE_DATAPATH__abc_16259_n5272) );
  OR2X2 OR2X2_1281 ( .A(AES_CORE_DATAPATH__abc_16259_n5273), .B(AES_CORE_DATAPATH__abc_16259_n5274_1), .Y(AES_CORE_DATAPATH__0key_2__31_0__0_) );
  OR2X2 OR2X2_1282 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_33_), .Y(AES_CORE_DATAPATH__abc_16259_n5276) );
  OR2X2 OR2X2_1283 ( .A(AES_CORE_DATAPATH__abc_16259_n5277_1), .B(AES_CORE_DATAPATH__abc_16259_n5278), .Y(AES_CORE_DATAPATH__abc_16259_n5279) );
  OR2X2 OR2X2_1284 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf10), .B(AES_CORE_DATAPATH__abc_16259_n5279), .Y(AES_CORE_DATAPATH__abc_16259_n5280_1) );
  OR2X2 OR2X2_1285 ( .A(AES_CORE_DATAPATH__abc_16259_n5282), .B(AES_CORE_DATAPATH__abc_16259_n5283_1), .Y(AES_CORE_DATAPATH__0key_2__31_0__1_) );
  OR2X2 OR2X2_1286 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf10), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_34_), .Y(AES_CORE_DATAPATH__abc_16259_n5285) );
  OR2X2 OR2X2_1287 ( .A(AES_CORE_DATAPATH__abc_16259_n5286_1), .B(AES_CORE_DATAPATH__abc_16259_n5287), .Y(AES_CORE_DATAPATH__abc_16259_n5288) );
  OR2X2 OR2X2_1288 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf9), .B(AES_CORE_DATAPATH__abc_16259_n5288), .Y(AES_CORE_DATAPATH__abc_16259_n5289_1) );
  OR2X2 OR2X2_1289 ( .A(AES_CORE_DATAPATH__abc_16259_n5291), .B(AES_CORE_DATAPATH__abc_16259_n5292_1), .Y(AES_CORE_DATAPATH__0key_2__31_0__2_) );
  OR2X2 OR2X2_129 ( .A(AES_CORE_DATAPATH__abc_16259_n2578_1), .B(AES_CORE_DATAPATH__abc_16259_n2579_1), .Y(_auto_iopadmap_cc_313_execute_26916_10_) );
  OR2X2 OR2X2_1290 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf9), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_35_), .Y(AES_CORE_DATAPATH__abc_16259_n5294) );
  OR2X2 OR2X2_1291 ( .A(AES_CORE_DATAPATH__abc_16259_n5295_1), .B(AES_CORE_DATAPATH__abc_16259_n5296), .Y(AES_CORE_DATAPATH__abc_16259_n5297) );
  OR2X2 OR2X2_1292 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf8), .B(AES_CORE_DATAPATH__abc_16259_n5297), .Y(AES_CORE_DATAPATH__abc_16259_n5298_1) );
  OR2X2 OR2X2_1293 ( .A(AES_CORE_DATAPATH__abc_16259_n5300), .B(AES_CORE_DATAPATH__abc_16259_n5301_1), .Y(AES_CORE_DATAPATH__0key_2__31_0__3_) );
  OR2X2 OR2X2_1294 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf8), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_36_), .Y(AES_CORE_DATAPATH__abc_16259_n5303) );
  OR2X2 OR2X2_1295 ( .A(AES_CORE_DATAPATH__abc_16259_n5304_1), .B(AES_CORE_DATAPATH__abc_16259_n5305), .Y(AES_CORE_DATAPATH__abc_16259_n5306) );
  OR2X2 OR2X2_1296 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf7), .B(AES_CORE_DATAPATH__abc_16259_n5306), .Y(AES_CORE_DATAPATH__abc_16259_n5307_1) );
  OR2X2 OR2X2_1297 ( .A(AES_CORE_DATAPATH__abc_16259_n5309), .B(AES_CORE_DATAPATH__abc_16259_n5310_1), .Y(AES_CORE_DATAPATH__0key_2__31_0__4_) );
  OR2X2 OR2X2_1298 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf7), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_37_), .Y(AES_CORE_DATAPATH__abc_16259_n5312) );
  OR2X2 OR2X2_1299 ( .A(AES_CORE_DATAPATH__abc_16259_n5313_1), .B(AES_CORE_DATAPATH__abc_16259_n5314), .Y(AES_CORE_DATAPATH__abc_16259_n5315) );
  OR2X2 OR2X2_13 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n115), .B(AES_CORE_CONTROL_UNIT__abc_15841_n108), .Y(AES_CORE_CONTROL_UNIT__abc_10818_n12) );
  OR2X2 OR2X2_130 ( .A(AES_CORE_DATAPATH__abc_16259_n2582), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n2583_1) );
  OR2X2 OR2X2_1300 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf6), .B(AES_CORE_DATAPATH__abc_16259_n5315), .Y(AES_CORE_DATAPATH__abc_16259_n5316_1) );
  OR2X2 OR2X2_1301 ( .A(AES_CORE_DATAPATH__abc_16259_n5318), .B(AES_CORE_DATAPATH__abc_16259_n5319_1), .Y(AES_CORE_DATAPATH__0key_2__31_0__5_) );
  OR2X2 OR2X2_1302 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf6), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_38_), .Y(AES_CORE_DATAPATH__abc_16259_n5321) );
  OR2X2 OR2X2_1303 ( .A(AES_CORE_DATAPATH__abc_16259_n5322_1), .B(AES_CORE_DATAPATH__abc_16259_n5323), .Y(AES_CORE_DATAPATH__abc_16259_n5324) );
  OR2X2 OR2X2_1304 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf5), .B(AES_CORE_DATAPATH__abc_16259_n5324), .Y(AES_CORE_DATAPATH__abc_16259_n5325_1) );
  OR2X2 OR2X2_1305 ( .A(AES_CORE_DATAPATH__abc_16259_n5327), .B(AES_CORE_DATAPATH__abc_16259_n5328_1), .Y(AES_CORE_DATAPATH__0key_2__31_0__6_) );
  OR2X2 OR2X2_1306 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf5), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_39_), .Y(AES_CORE_DATAPATH__abc_16259_n5330) );
  OR2X2 OR2X2_1307 ( .A(AES_CORE_DATAPATH__abc_16259_n5331_1), .B(AES_CORE_DATAPATH__abc_16259_n5332), .Y(AES_CORE_DATAPATH__abc_16259_n5333) );
  OR2X2 OR2X2_1308 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n5333), .Y(AES_CORE_DATAPATH__abc_16259_n5334_1) );
  OR2X2 OR2X2_1309 ( .A(AES_CORE_DATAPATH__abc_16259_n5336), .B(AES_CORE_DATAPATH__abc_16259_n5337_1), .Y(AES_CORE_DATAPATH__0key_2__31_0__7_) );
  OR2X2 OR2X2_131 ( .A(AES_CORE_DATAPATH__abc_16259_n2581_1), .B(AES_CORE_DATAPATH__abc_16259_n2583_1), .Y(AES_CORE_DATAPATH__abc_16259_n2584_1) );
  OR2X2 OR2X2_1310 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_40_), .Y(AES_CORE_DATAPATH__abc_16259_n5339) );
  OR2X2 OR2X2_1311 ( .A(AES_CORE_DATAPATH__abc_16259_n5340_1), .B(AES_CORE_DATAPATH__abc_16259_n5341), .Y(AES_CORE_DATAPATH__abc_16259_n5342) );
  OR2X2 OR2X2_1312 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n5342), .Y(AES_CORE_DATAPATH__abc_16259_n5343_1) );
  OR2X2 OR2X2_1313 ( .A(AES_CORE_DATAPATH__abc_16259_n5345), .B(AES_CORE_DATAPATH__abc_16259_n5346_1), .Y(AES_CORE_DATAPATH__0key_2__31_0__8_) );
  OR2X2 OR2X2_1314 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_41_), .Y(AES_CORE_DATAPATH__abc_16259_n5348) );
  OR2X2 OR2X2_1315 ( .A(AES_CORE_DATAPATH__abc_16259_n5349_1), .B(AES_CORE_DATAPATH__abc_16259_n5350), .Y(AES_CORE_DATAPATH__abc_16259_n5351) );
  OR2X2 OR2X2_1316 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n5351), .Y(AES_CORE_DATAPATH__abc_16259_n5352_1) );
  OR2X2 OR2X2_1317 ( .A(AES_CORE_DATAPATH__abc_16259_n5354), .B(AES_CORE_DATAPATH__abc_16259_n5355_1), .Y(AES_CORE_DATAPATH__0key_2__31_0__9_) );
  OR2X2 OR2X2_1318 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_42_), .Y(AES_CORE_DATAPATH__abc_16259_n5357) );
  OR2X2 OR2X2_1319 ( .A(AES_CORE_DATAPATH__abc_16259_n5358_1), .B(AES_CORE_DATAPATH__abc_16259_n5359), .Y(AES_CORE_DATAPATH__abc_16259_n5360) );
  OR2X2 OR2X2_132 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf4), .B(AES_CORE_DATAPATH_iv_2__11_), .Y(AES_CORE_DATAPATH__abc_16259_n2585) );
  OR2X2 OR2X2_1320 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n5360), .Y(AES_CORE_DATAPATH__abc_16259_n5361_1) );
  OR2X2 OR2X2_1321 ( .A(AES_CORE_DATAPATH__abc_16259_n5363), .B(AES_CORE_DATAPATH__abc_16259_n5364_1), .Y(AES_CORE_DATAPATH__0key_2__31_0__10_) );
  OR2X2 OR2X2_1322 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_43_), .Y(AES_CORE_DATAPATH__abc_16259_n5366) );
  OR2X2 OR2X2_1323 ( .A(AES_CORE_DATAPATH__abc_16259_n5367_1), .B(AES_CORE_DATAPATH__abc_16259_n5368_1), .Y(AES_CORE_DATAPATH__abc_16259_n5369_1) );
  OR2X2 OR2X2_1324 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n5369_1), .Y(AES_CORE_DATAPATH__abc_16259_n5370_1) );
  OR2X2 OR2X2_1325 ( .A(AES_CORE_DATAPATH__abc_16259_n5372_1), .B(AES_CORE_DATAPATH__abc_16259_n5373_1), .Y(AES_CORE_DATAPATH__0key_2__31_0__11_) );
  OR2X2 OR2X2_1326 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_44_), .Y(AES_CORE_DATAPATH__abc_16259_n5375_1) );
  OR2X2 OR2X2_1327 ( .A(AES_CORE_DATAPATH__abc_16259_n5376_1), .B(AES_CORE_DATAPATH__abc_16259_n5377_1), .Y(AES_CORE_DATAPATH__abc_16259_n5378_1) );
  OR2X2 OR2X2_1328 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf10), .B(AES_CORE_DATAPATH__abc_16259_n5378_1), .Y(AES_CORE_DATAPATH__abc_16259_n5379_1) );
  OR2X2 OR2X2_1329 ( .A(AES_CORE_DATAPATH__abc_16259_n5381_1), .B(AES_CORE_DATAPATH__abc_16259_n5382_1), .Y(AES_CORE_DATAPATH__0key_2__31_0__12_) );
  OR2X2 OR2X2_133 ( .A(AES_CORE_DATAPATH__abc_16259_n2587), .B(AES_CORE_DATAPATH__abc_16259_n2588_1), .Y(_auto_iopadmap_cc_313_execute_26916_11_) );
  OR2X2 OR2X2_1330 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf10), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_45_), .Y(AES_CORE_DATAPATH__abc_16259_n5384_1) );
  OR2X2 OR2X2_1331 ( .A(AES_CORE_DATAPATH__abc_16259_n5385_1), .B(AES_CORE_DATAPATH__abc_16259_n5386_1), .Y(AES_CORE_DATAPATH__abc_16259_n5387_1) );
  OR2X2 OR2X2_1332 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf9), .B(AES_CORE_DATAPATH__abc_16259_n5387_1), .Y(AES_CORE_DATAPATH__abc_16259_n5388_1) );
  OR2X2 OR2X2_1333 ( .A(AES_CORE_DATAPATH__abc_16259_n5390_1), .B(AES_CORE_DATAPATH__abc_16259_n5391_1), .Y(AES_CORE_DATAPATH__0key_2__31_0__13_) );
  OR2X2 OR2X2_1334 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf9), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_46_), .Y(AES_CORE_DATAPATH__abc_16259_n5393_1) );
  OR2X2 OR2X2_1335 ( .A(AES_CORE_DATAPATH__abc_16259_n5394_1), .B(AES_CORE_DATAPATH__abc_16259_n5395_1), .Y(AES_CORE_DATAPATH__abc_16259_n5396_1) );
  OR2X2 OR2X2_1336 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf8), .B(AES_CORE_DATAPATH__abc_16259_n5396_1), .Y(AES_CORE_DATAPATH__abc_16259_n5397_1) );
  OR2X2 OR2X2_1337 ( .A(AES_CORE_DATAPATH__abc_16259_n5399_1), .B(AES_CORE_DATAPATH__abc_16259_n5400_1), .Y(AES_CORE_DATAPATH__0key_2__31_0__14_) );
  OR2X2 OR2X2_1338 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf8), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_47_), .Y(AES_CORE_DATAPATH__abc_16259_n5402_1) );
  OR2X2 OR2X2_1339 ( .A(AES_CORE_DATAPATH__abc_16259_n5403_1), .B(AES_CORE_DATAPATH__abc_16259_n5404_1), .Y(AES_CORE_DATAPATH__abc_16259_n5405_1) );
  OR2X2 OR2X2_134 ( .A(AES_CORE_DATAPATH__abc_16259_n2591_1), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n2592) );
  OR2X2 OR2X2_1340 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf7), .B(AES_CORE_DATAPATH__abc_16259_n5405_1), .Y(AES_CORE_DATAPATH__abc_16259_n5406_1) );
  OR2X2 OR2X2_1341 ( .A(AES_CORE_DATAPATH__abc_16259_n5408_1), .B(AES_CORE_DATAPATH__abc_16259_n5409_1), .Y(AES_CORE_DATAPATH__0key_2__31_0__15_) );
  OR2X2 OR2X2_1342 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf7), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_48_), .Y(AES_CORE_DATAPATH__abc_16259_n5411_1) );
  OR2X2 OR2X2_1343 ( .A(AES_CORE_DATAPATH__abc_16259_n5412_1), .B(AES_CORE_DATAPATH__abc_16259_n5413_1), .Y(AES_CORE_DATAPATH__abc_16259_n5414_1) );
  OR2X2 OR2X2_1344 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf6), .B(AES_CORE_DATAPATH__abc_16259_n5414_1), .Y(AES_CORE_DATAPATH__abc_16259_n5415_1) );
  OR2X2 OR2X2_1345 ( .A(AES_CORE_DATAPATH__abc_16259_n5417_1), .B(AES_CORE_DATAPATH__abc_16259_n5418_1), .Y(AES_CORE_DATAPATH__0key_2__31_0__16_) );
  OR2X2 OR2X2_1346 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf6), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_49_), .Y(AES_CORE_DATAPATH__abc_16259_n5420_1) );
  OR2X2 OR2X2_1347 ( .A(AES_CORE_DATAPATH__abc_16259_n5421_1), .B(AES_CORE_DATAPATH__abc_16259_n5422_1), .Y(AES_CORE_DATAPATH__abc_16259_n5423_1) );
  OR2X2 OR2X2_1348 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf5), .B(AES_CORE_DATAPATH__abc_16259_n5423_1), .Y(AES_CORE_DATAPATH__abc_16259_n5424_1) );
  OR2X2 OR2X2_1349 ( .A(AES_CORE_DATAPATH__abc_16259_n5426_1), .B(AES_CORE_DATAPATH__abc_16259_n5427_1), .Y(AES_CORE_DATAPATH__0key_2__31_0__17_) );
  OR2X2 OR2X2_135 ( .A(AES_CORE_DATAPATH__abc_16259_n2590), .B(AES_CORE_DATAPATH__abc_16259_n2592), .Y(AES_CORE_DATAPATH__abc_16259_n2593_1) );
  OR2X2 OR2X2_1350 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf5), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_50_), .Y(AES_CORE_DATAPATH__abc_16259_n5429_1) );
  OR2X2 OR2X2_1351 ( .A(AES_CORE_DATAPATH__abc_16259_n5430_1), .B(AES_CORE_DATAPATH__abc_16259_n5431_1), .Y(AES_CORE_DATAPATH__abc_16259_n5432_1) );
  OR2X2 OR2X2_1352 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n5432_1), .Y(AES_CORE_DATAPATH__abc_16259_n5433_1) );
  OR2X2 OR2X2_1353 ( .A(AES_CORE_DATAPATH__abc_16259_n5435_1), .B(AES_CORE_DATAPATH__abc_16259_n5436_1), .Y(AES_CORE_DATAPATH__0key_2__31_0__18_) );
  OR2X2 OR2X2_1354 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_51_), .Y(AES_CORE_DATAPATH__abc_16259_n5438_1) );
  OR2X2 OR2X2_1355 ( .A(AES_CORE_DATAPATH__abc_16259_n5439_1), .B(AES_CORE_DATAPATH__abc_16259_n5440_1), .Y(AES_CORE_DATAPATH__abc_16259_n5441_1) );
  OR2X2 OR2X2_1356 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n5441_1), .Y(AES_CORE_DATAPATH__abc_16259_n5442_1) );
  OR2X2 OR2X2_1357 ( .A(AES_CORE_DATAPATH__abc_16259_n5444_1), .B(AES_CORE_DATAPATH__abc_16259_n5445_1), .Y(AES_CORE_DATAPATH__0key_2__31_0__19_) );
  OR2X2 OR2X2_1358 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_52_), .Y(AES_CORE_DATAPATH__abc_16259_n5447_1) );
  OR2X2 OR2X2_1359 ( .A(AES_CORE_DATAPATH__abc_16259_n5448_1), .B(AES_CORE_DATAPATH__abc_16259_n5449_1), .Y(AES_CORE_DATAPATH__abc_16259_n5450_1) );
  OR2X2 OR2X2_136 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf3), .B(AES_CORE_DATAPATH_iv_2__12_), .Y(AES_CORE_DATAPATH__abc_16259_n2594_1) );
  OR2X2 OR2X2_1360 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n5450_1), .Y(AES_CORE_DATAPATH__abc_16259_n5451_1) );
  OR2X2 OR2X2_1361 ( .A(AES_CORE_DATAPATH__abc_16259_n5453), .B(AES_CORE_DATAPATH__abc_16259_n5454), .Y(AES_CORE_DATAPATH__0key_2__31_0__20_) );
  OR2X2 OR2X2_1362 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_53_), .Y(AES_CORE_DATAPATH__abc_16259_n5456) );
  OR2X2 OR2X2_1363 ( .A(AES_CORE_DATAPATH__abc_16259_n5457), .B(AES_CORE_DATAPATH__abc_16259_n5458), .Y(AES_CORE_DATAPATH__abc_16259_n5459) );
  OR2X2 OR2X2_1364 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n5459), .Y(AES_CORE_DATAPATH__abc_16259_n5460) );
  OR2X2 OR2X2_1365 ( .A(AES_CORE_DATAPATH__abc_16259_n5462), .B(AES_CORE_DATAPATH__abc_16259_n5463), .Y(AES_CORE_DATAPATH__0key_2__31_0__21_) );
  OR2X2 OR2X2_1366 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_54_), .Y(AES_CORE_DATAPATH__abc_16259_n5465) );
  OR2X2 OR2X2_1367 ( .A(AES_CORE_DATAPATH__abc_16259_n5466), .B(AES_CORE_DATAPATH__abc_16259_n5467), .Y(AES_CORE_DATAPATH__abc_16259_n5468) );
  OR2X2 OR2X2_1368 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n5468), .Y(AES_CORE_DATAPATH__abc_16259_n5469) );
  OR2X2 OR2X2_1369 ( .A(AES_CORE_DATAPATH__abc_16259_n5471), .B(AES_CORE_DATAPATH__abc_16259_n5472), .Y(AES_CORE_DATAPATH__0key_2__31_0__22_) );
  OR2X2 OR2X2_137 ( .A(AES_CORE_DATAPATH__abc_16259_n2596_1), .B(AES_CORE_DATAPATH__abc_16259_n2597), .Y(_auto_iopadmap_cc_313_execute_26916_12_) );
  OR2X2 OR2X2_1370 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_55_), .Y(AES_CORE_DATAPATH__abc_16259_n5474) );
  OR2X2 OR2X2_1371 ( .A(AES_CORE_DATAPATH__abc_16259_n5475), .B(AES_CORE_DATAPATH__abc_16259_n5476), .Y(AES_CORE_DATAPATH__abc_16259_n5477) );
  OR2X2 OR2X2_1372 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf10), .B(AES_CORE_DATAPATH__abc_16259_n5477), .Y(AES_CORE_DATAPATH__abc_16259_n5478) );
  OR2X2 OR2X2_1373 ( .A(AES_CORE_DATAPATH__abc_16259_n5480), .B(AES_CORE_DATAPATH__abc_16259_n5481), .Y(AES_CORE_DATAPATH__0key_2__31_0__23_) );
  OR2X2 OR2X2_1374 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf10), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_56_), .Y(AES_CORE_DATAPATH__abc_16259_n5483) );
  OR2X2 OR2X2_1375 ( .A(AES_CORE_DATAPATH__abc_16259_n5484), .B(AES_CORE_DATAPATH__abc_16259_n5485), .Y(AES_CORE_DATAPATH__abc_16259_n5486) );
  OR2X2 OR2X2_1376 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf9), .B(AES_CORE_DATAPATH__abc_16259_n5486), .Y(AES_CORE_DATAPATH__abc_16259_n5487) );
  OR2X2 OR2X2_1377 ( .A(AES_CORE_DATAPATH__abc_16259_n5489), .B(AES_CORE_DATAPATH__abc_16259_n5490), .Y(AES_CORE_DATAPATH__0key_2__31_0__24_) );
  OR2X2 OR2X2_1378 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf9), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_57_), .Y(AES_CORE_DATAPATH__abc_16259_n5492) );
  OR2X2 OR2X2_1379 ( .A(AES_CORE_DATAPATH__abc_16259_n5493), .B(AES_CORE_DATAPATH__abc_16259_n5494), .Y(AES_CORE_DATAPATH__abc_16259_n5495) );
  OR2X2 OR2X2_138 ( .A(AES_CORE_DATAPATH__abc_16259_n2600), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n2601_1) );
  OR2X2 OR2X2_1380 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf8), .B(AES_CORE_DATAPATH__abc_16259_n5495), .Y(AES_CORE_DATAPATH__abc_16259_n5496) );
  OR2X2 OR2X2_1381 ( .A(AES_CORE_DATAPATH__abc_16259_n5498), .B(AES_CORE_DATAPATH__abc_16259_n5499), .Y(AES_CORE_DATAPATH__0key_2__31_0__25_) );
  OR2X2 OR2X2_1382 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf8), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_58_), .Y(AES_CORE_DATAPATH__abc_16259_n5501) );
  OR2X2 OR2X2_1383 ( .A(AES_CORE_DATAPATH__abc_16259_n5502), .B(AES_CORE_DATAPATH__abc_16259_n5503), .Y(AES_CORE_DATAPATH__abc_16259_n5504) );
  OR2X2 OR2X2_1384 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf7), .B(AES_CORE_DATAPATH__abc_16259_n5504), .Y(AES_CORE_DATAPATH__abc_16259_n5505) );
  OR2X2 OR2X2_1385 ( .A(AES_CORE_DATAPATH__abc_16259_n5507), .B(AES_CORE_DATAPATH__abc_16259_n5508), .Y(AES_CORE_DATAPATH__0key_2__31_0__26_) );
  OR2X2 OR2X2_1386 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf7), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_59_), .Y(AES_CORE_DATAPATH__abc_16259_n5510) );
  OR2X2 OR2X2_1387 ( .A(AES_CORE_DATAPATH__abc_16259_n5511), .B(AES_CORE_DATAPATH__abc_16259_n5512), .Y(AES_CORE_DATAPATH__abc_16259_n5513) );
  OR2X2 OR2X2_1388 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf6), .B(AES_CORE_DATAPATH__abc_16259_n5513), .Y(AES_CORE_DATAPATH__abc_16259_n5514) );
  OR2X2 OR2X2_1389 ( .A(AES_CORE_DATAPATH__abc_16259_n5516), .B(AES_CORE_DATAPATH__abc_16259_n5517), .Y(AES_CORE_DATAPATH__0key_2__31_0__27_) );
  OR2X2 OR2X2_139 ( .A(AES_CORE_DATAPATH__abc_16259_n2599_1), .B(AES_CORE_DATAPATH__abc_16259_n2601_1), .Y(AES_CORE_DATAPATH__abc_16259_n2602) );
  OR2X2 OR2X2_1390 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf6), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_60_), .Y(AES_CORE_DATAPATH__abc_16259_n5519) );
  OR2X2 OR2X2_1391 ( .A(AES_CORE_DATAPATH__abc_16259_n5520), .B(AES_CORE_DATAPATH__abc_16259_n5521), .Y(AES_CORE_DATAPATH__abc_16259_n5522) );
  OR2X2 OR2X2_1392 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf5), .B(AES_CORE_DATAPATH__abc_16259_n5522), .Y(AES_CORE_DATAPATH__abc_16259_n5523) );
  OR2X2 OR2X2_1393 ( .A(AES_CORE_DATAPATH__abc_16259_n5525), .B(AES_CORE_DATAPATH__abc_16259_n5526), .Y(AES_CORE_DATAPATH__0key_2__31_0__28_) );
  OR2X2 OR2X2_1394 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf5), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_61_), .Y(AES_CORE_DATAPATH__abc_16259_n5528) );
  OR2X2 OR2X2_1395 ( .A(AES_CORE_DATAPATH__abc_16259_n5529), .B(AES_CORE_DATAPATH__abc_16259_n5530), .Y(AES_CORE_DATAPATH__abc_16259_n5531) );
  OR2X2 OR2X2_1396 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n5531), .Y(AES_CORE_DATAPATH__abc_16259_n5532) );
  OR2X2 OR2X2_1397 ( .A(AES_CORE_DATAPATH__abc_16259_n5534), .B(AES_CORE_DATAPATH__abc_16259_n5535), .Y(AES_CORE_DATAPATH__0key_2__31_0__29_) );
  OR2X2 OR2X2_1398 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_62_), .Y(AES_CORE_DATAPATH__abc_16259_n5537) );
  OR2X2 OR2X2_1399 ( .A(AES_CORE_DATAPATH__abc_16259_n5538), .B(AES_CORE_DATAPATH__abc_16259_n5539), .Y(AES_CORE_DATAPATH__abc_16259_n5540) );
  OR2X2 OR2X2_14 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n117_1), .B(AES_CORE_CONTROL_UNIT__abc_15841_n118), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n119) );
  OR2X2 OR2X2_140 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf2), .B(AES_CORE_DATAPATH_iv_2__13_), .Y(AES_CORE_DATAPATH__abc_16259_n2603_1) );
  OR2X2 OR2X2_1400 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n5540), .Y(AES_CORE_DATAPATH__abc_16259_n5541) );
  OR2X2 OR2X2_1401 ( .A(AES_CORE_DATAPATH__abc_16259_n5543), .B(AES_CORE_DATAPATH__abc_16259_n5544), .Y(AES_CORE_DATAPATH__0key_2__31_0__30_) );
  OR2X2 OR2X2_1402 ( .A(AES_CORE_DATAPATH__abc_16259_n5546), .B(AES_CORE_DATAPATH__abc_16259_n5547), .Y(AES_CORE_DATAPATH__abc_16259_n5548) );
  OR2X2 OR2X2_1403 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n5548), .Y(AES_CORE_DATAPATH__abc_16259_n5549) );
  OR2X2 OR2X2_1404 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_63_), .Y(AES_CORE_DATAPATH__abc_16259_n5550) );
  OR2X2 OR2X2_1405 ( .A(AES_CORE_DATAPATH__abc_16259_n5552), .B(AES_CORE_DATAPATH__abc_16259_n5553), .Y(AES_CORE_DATAPATH__0key_2__31_0__31_) );
  OR2X2 OR2X2_1406 ( .A(AES_CORE_DATAPATH__abc_16259_n5556), .B(AES_CORE_DATAPATH__abc_16259_n5555), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__0_) );
  OR2X2 OR2X2_1407 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__1_), .Y(AES_CORE_DATAPATH__abc_16259_n5558) );
  OR2X2 OR2X2_1408 ( .A(AES_CORE_DATAPATH__abc_16259_n5279), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf10), .Y(AES_CORE_DATAPATH__abc_16259_n5559) );
  OR2X2 OR2X2_1409 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf10), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__2_), .Y(AES_CORE_DATAPATH__abc_16259_n5561) );
  OR2X2 OR2X2_141 ( .A(AES_CORE_DATAPATH__abc_16259_n2605), .B(AES_CORE_DATAPATH__abc_16259_n2606_1), .Y(_auto_iopadmap_cc_313_execute_26916_13_) );
  OR2X2 OR2X2_1410 ( .A(AES_CORE_DATAPATH__abc_16259_n5288), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf9), .Y(AES_CORE_DATAPATH__abc_16259_n5562) );
  OR2X2 OR2X2_1411 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf9), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__3_), .Y(AES_CORE_DATAPATH__abc_16259_n5564) );
  OR2X2 OR2X2_1412 ( .A(AES_CORE_DATAPATH__abc_16259_n5297), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf8), .Y(AES_CORE_DATAPATH__abc_16259_n5565) );
  OR2X2 OR2X2_1413 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf8), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__4_), .Y(AES_CORE_DATAPATH__abc_16259_n5567) );
  OR2X2 OR2X2_1414 ( .A(AES_CORE_DATAPATH__abc_16259_n5306), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n5568) );
  OR2X2 OR2X2_1415 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf7), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__5_), .Y(AES_CORE_DATAPATH__abc_16259_n5570) );
  OR2X2 OR2X2_1416 ( .A(AES_CORE_DATAPATH__abc_16259_n5315), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n5571) );
  OR2X2 OR2X2_1417 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf6), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__6_), .Y(AES_CORE_DATAPATH__abc_16259_n5573) );
  OR2X2 OR2X2_1418 ( .A(AES_CORE_DATAPATH__abc_16259_n5324), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n5574) );
  OR2X2 OR2X2_1419 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf5), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__7_), .Y(AES_CORE_DATAPATH__abc_16259_n5576) );
  OR2X2 OR2X2_142 ( .A(AES_CORE_DATAPATH__abc_16259_n2609_1), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n2610) );
  OR2X2 OR2X2_1420 ( .A(AES_CORE_DATAPATH__abc_16259_n5333), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5577) );
  OR2X2 OR2X2_1421 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__8_), .Y(AES_CORE_DATAPATH__abc_16259_n5579) );
  OR2X2 OR2X2_1422 ( .A(AES_CORE_DATAPATH__abc_16259_n5342), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n5580) );
  OR2X2 OR2X2_1423 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__9_), .Y(AES_CORE_DATAPATH__abc_16259_n5582) );
  OR2X2 OR2X2_1424 ( .A(AES_CORE_DATAPATH__abc_16259_n5351), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n5583) );
  OR2X2 OR2X2_1425 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__10_), .Y(AES_CORE_DATAPATH__abc_16259_n5585) );
  OR2X2 OR2X2_1426 ( .A(AES_CORE_DATAPATH__abc_16259_n5360), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n5586) );
  OR2X2 OR2X2_1427 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__11_), .Y(AES_CORE_DATAPATH__abc_16259_n5588) );
  OR2X2 OR2X2_1428 ( .A(AES_CORE_DATAPATH__abc_16259_n5369_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n5589) );
  OR2X2 OR2X2_1429 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__12_), .Y(AES_CORE_DATAPATH__abc_16259_n5591) );
  OR2X2 OR2X2_143 ( .A(AES_CORE_DATAPATH__abc_16259_n2608_1), .B(AES_CORE_DATAPATH__abc_16259_n2610), .Y(AES_CORE_DATAPATH__abc_16259_n2611_1) );
  OR2X2 OR2X2_1430 ( .A(AES_CORE_DATAPATH__abc_16259_n5378_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf10), .Y(AES_CORE_DATAPATH__abc_16259_n5592) );
  OR2X2 OR2X2_1431 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf10), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__13_), .Y(AES_CORE_DATAPATH__abc_16259_n5594) );
  OR2X2 OR2X2_1432 ( .A(AES_CORE_DATAPATH__abc_16259_n5387_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf9), .Y(AES_CORE_DATAPATH__abc_16259_n5595) );
  OR2X2 OR2X2_1433 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf9), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__14_), .Y(AES_CORE_DATAPATH__abc_16259_n5597) );
  OR2X2 OR2X2_1434 ( .A(AES_CORE_DATAPATH__abc_16259_n5396_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf8), .Y(AES_CORE_DATAPATH__abc_16259_n5598) );
  OR2X2 OR2X2_1435 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf8), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__15_), .Y(AES_CORE_DATAPATH__abc_16259_n5600) );
  OR2X2 OR2X2_1436 ( .A(AES_CORE_DATAPATH__abc_16259_n5405_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n5601) );
  OR2X2 OR2X2_1437 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf7), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__16_), .Y(AES_CORE_DATAPATH__abc_16259_n5603) );
  OR2X2 OR2X2_1438 ( .A(AES_CORE_DATAPATH__abc_16259_n5414_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n5604) );
  OR2X2 OR2X2_1439 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf6), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__17_), .Y(AES_CORE_DATAPATH__abc_16259_n5606) );
  OR2X2 OR2X2_144 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf1), .B(AES_CORE_DATAPATH_iv_2__14_), .Y(AES_CORE_DATAPATH__abc_16259_n2612) );
  OR2X2 OR2X2_1440 ( .A(AES_CORE_DATAPATH__abc_16259_n5423_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n5607) );
  OR2X2 OR2X2_1441 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf5), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__18_), .Y(AES_CORE_DATAPATH__abc_16259_n5609) );
  OR2X2 OR2X2_1442 ( .A(AES_CORE_DATAPATH__abc_16259_n5432_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5610) );
  OR2X2 OR2X2_1443 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__19_), .Y(AES_CORE_DATAPATH__abc_16259_n5612) );
  OR2X2 OR2X2_1444 ( .A(AES_CORE_DATAPATH__abc_16259_n5441_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n5613) );
  OR2X2 OR2X2_1445 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__20_), .Y(AES_CORE_DATAPATH__abc_16259_n5615) );
  OR2X2 OR2X2_1446 ( .A(AES_CORE_DATAPATH__abc_16259_n5450_1), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n5616) );
  OR2X2 OR2X2_1447 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__21_), .Y(AES_CORE_DATAPATH__abc_16259_n5618) );
  OR2X2 OR2X2_1448 ( .A(AES_CORE_DATAPATH__abc_16259_n5459), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n5619) );
  OR2X2 OR2X2_1449 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__22_), .Y(AES_CORE_DATAPATH__abc_16259_n5621) );
  OR2X2 OR2X2_145 ( .A(AES_CORE_DATAPATH__abc_16259_n2614_1), .B(AES_CORE_DATAPATH__abc_16259_n2615), .Y(_auto_iopadmap_cc_313_execute_26916_14_) );
  OR2X2 OR2X2_1450 ( .A(AES_CORE_DATAPATH__abc_16259_n5468), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n5622) );
  OR2X2 OR2X2_1451 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__23_), .Y(AES_CORE_DATAPATH__abc_16259_n5624) );
  OR2X2 OR2X2_1452 ( .A(AES_CORE_DATAPATH__abc_16259_n5477), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf10), .Y(AES_CORE_DATAPATH__abc_16259_n5625) );
  OR2X2 OR2X2_1453 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf10), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__24_), .Y(AES_CORE_DATAPATH__abc_16259_n5627) );
  OR2X2 OR2X2_1454 ( .A(AES_CORE_DATAPATH__abc_16259_n5486), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf9), .Y(AES_CORE_DATAPATH__abc_16259_n5628) );
  OR2X2 OR2X2_1455 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf9), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__25_), .Y(AES_CORE_DATAPATH__abc_16259_n5630) );
  OR2X2 OR2X2_1456 ( .A(AES_CORE_DATAPATH__abc_16259_n5495), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf8), .Y(AES_CORE_DATAPATH__abc_16259_n5631) );
  OR2X2 OR2X2_1457 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf8), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__26_), .Y(AES_CORE_DATAPATH__abc_16259_n5633) );
  OR2X2 OR2X2_1458 ( .A(AES_CORE_DATAPATH__abc_16259_n5504), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n5634) );
  OR2X2 OR2X2_1459 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf7), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__27_), .Y(AES_CORE_DATAPATH__abc_16259_n5636) );
  OR2X2 OR2X2_146 ( .A(AES_CORE_DATAPATH__abc_16259_n2618_1), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n2619_1) );
  OR2X2 OR2X2_1460 ( .A(AES_CORE_DATAPATH__abc_16259_n5513), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n5637) );
  OR2X2 OR2X2_1461 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf6), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__28_), .Y(AES_CORE_DATAPATH__abc_16259_n5639) );
  OR2X2 OR2X2_1462 ( .A(AES_CORE_DATAPATH__abc_16259_n5522), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n5640) );
  OR2X2 OR2X2_1463 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf5), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__29_), .Y(AES_CORE_DATAPATH__abc_16259_n5642) );
  OR2X2 OR2X2_1464 ( .A(AES_CORE_DATAPATH__abc_16259_n5531), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5643) );
  OR2X2 OR2X2_1465 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__30_), .Y(AES_CORE_DATAPATH__abc_16259_n5645) );
  OR2X2 OR2X2_1466 ( .A(AES_CORE_DATAPATH__abc_16259_n5540), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n5646) );
  OR2X2 OR2X2_1467 ( .A(AES_CORE_DATAPATH__abc_16259_n5548), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n5648) );
  OR2X2 OR2X2_1468 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__31_), .Y(AES_CORE_DATAPATH__abc_16259_n5649) );
  OR2X2 OR2X2_1469 ( .A(AES_CORE_DATAPATH__abc_16259_n5662), .B(AES_CORE_DATAPATH__abc_16259_n5661), .Y(AES_CORE_DATAPATH__abc_16259_n5663) );
  OR2X2 OR2X2_147 ( .A(AES_CORE_DATAPATH__abc_16259_n2617), .B(AES_CORE_DATAPATH__abc_16259_n2619_1), .Y(AES_CORE_DATAPATH__abc_16259_n2620) );
  OR2X2 OR2X2_1470 ( .A(AES_CORE_DATAPATH__abc_16259_n5664), .B(AES_CORE_DATAPATH__abc_16259_n5660), .Y(AES_CORE_DATAPATH__abc_16259_n5665) );
  OR2X2 OR2X2_1471 ( .A(AES_CORE_DATAPATH__abc_16259_n5666), .B(AES_CORE_DATAPATH__abc_16259_n5667), .Y(AES_CORE_DATAPATH__0key_3__31_0__0_) );
  OR2X2 OR2X2_1472 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_1_), .Y(AES_CORE_DATAPATH__abc_16259_n5669) );
  OR2X2 OR2X2_1473 ( .A(AES_CORE_DATAPATH__abc_16259_n5670), .B(AES_CORE_DATAPATH__abc_16259_n5671), .Y(AES_CORE_DATAPATH__abc_16259_n5672) );
  OR2X2 OR2X2_1474 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n5672), .Y(AES_CORE_DATAPATH__abc_16259_n5673) );
  OR2X2 OR2X2_1475 ( .A(AES_CORE_DATAPATH__abc_16259_n5675), .B(AES_CORE_DATAPATH__abc_16259_n5676), .Y(AES_CORE_DATAPATH__0key_3__31_0__1_) );
  OR2X2 OR2X2_1476 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_2_), .Y(AES_CORE_DATAPATH__abc_16259_n5678) );
  OR2X2 OR2X2_1477 ( .A(AES_CORE_DATAPATH__abc_16259_n5679), .B(AES_CORE_DATAPATH__abc_16259_n5680), .Y(AES_CORE_DATAPATH__abc_16259_n5681) );
  OR2X2 OR2X2_1478 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf10), .B(AES_CORE_DATAPATH__abc_16259_n5681), .Y(AES_CORE_DATAPATH__abc_16259_n5682) );
  OR2X2 OR2X2_1479 ( .A(AES_CORE_DATAPATH__abc_16259_n5684), .B(AES_CORE_DATAPATH__abc_16259_n5685), .Y(AES_CORE_DATAPATH__0key_3__31_0__2_) );
  OR2X2 OR2X2_148 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf0), .B(AES_CORE_DATAPATH_iv_2__15_), .Y(AES_CORE_DATAPATH__abc_16259_n2621_1) );
  OR2X2 OR2X2_1480 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf10), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_3_), .Y(AES_CORE_DATAPATH__abc_16259_n5687) );
  OR2X2 OR2X2_1481 ( .A(AES_CORE_DATAPATH__abc_16259_n5688), .B(AES_CORE_DATAPATH__abc_16259_n5689), .Y(AES_CORE_DATAPATH__abc_16259_n5690) );
  OR2X2 OR2X2_1482 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf9), .B(AES_CORE_DATAPATH__abc_16259_n5690), .Y(AES_CORE_DATAPATH__abc_16259_n5691) );
  OR2X2 OR2X2_1483 ( .A(AES_CORE_DATAPATH__abc_16259_n5693), .B(AES_CORE_DATAPATH__abc_16259_n5694), .Y(AES_CORE_DATAPATH__0key_3__31_0__3_) );
  OR2X2 OR2X2_1484 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf9), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_4_), .Y(AES_CORE_DATAPATH__abc_16259_n5696) );
  OR2X2 OR2X2_1485 ( .A(AES_CORE_DATAPATH__abc_16259_n5697), .B(AES_CORE_DATAPATH__abc_16259_n5698), .Y(AES_CORE_DATAPATH__abc_16259_n5699) );
  OR2X2 OR2X2_1486 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf8), .B(AES_CORE_DATAPATH__abc_16259_n5699), .Y(AES_CORE_DATAPATH__abc_16259_n5700) );
  OR2X2 OR2X2_1487 ( .A(AES_CORE_DATAPATH__abc_16259_n5702), .B(AES_CORE_DATAPATH__abc_16259_n5703), .Y(AES_CORE_DATAPATH__0key_3__31_0__4_) );
  OR2X2 OR2X2_1488 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf8), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_5_), .Y(AES_CORE_DATAPATH__abc_16259_n5705) );
  OR2X2 OR2X2_1489 ( .A(AES_CORE_DATAPATH__abc_16259_n5706), .B(AES_CORE_DATAPATH__abc_16259_n5707), .Y(AES_CORE_DATAPATH__abc_16259_n5708) );
  OR2X2 OR2X2_149 ( .A(AES_CORE_DATAPATH__abc_16259_n2623_1), .B(AES_CORE_DATAPATH__abc_16259_n2624_1), .Y(_auto_iopadmap_cc_313_execute_26916_15_) );
  OR2X2 OR2X2_1490 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf7), .B(AES_CORE_DATAPATH__abc_16259_n5708), .Y(AES_CORE_DATAPATH__abc_16259_n5709) );
  OR2X2 OR2X2_1491 ( .A(AES_CORE_DATAPATH__abc_16259_n5711), .B(AES_CORE_DATAPATH__abc_16259_n5712), .Y(AES_CORE_DATAPATH__0key_3__31_0__5_) );
  OR2X2 OR2X2_1492 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf7), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_6_), .Y(AES_CORE_DATAPATH__abc_16259_n5714) );
  OR2X2 OR2X2_1493 ( .A(AES_CORE_DATAPATH__abc_16259_n5715), .B(AES_CORE_DATAPATH__abc_16259_n5716), .Y(AES_CORE_DATAPATH__abc_16259_n5717) );
  OR2X2 OR2X2_1494 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf6), .B(AES_CORE_DATAPATH__abc_16259_n5717), .Y(AES_CORE_DATAPATH__abc_16259_n5718) );
  OR2X2 OR2X2_1495 ( .A(AES_CORE_DATAPATH__abc_16259_n5719), .B(AES_CORE_DATAPATH__abc_16259_n5658_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n5720) );
  OR2X2 OR2X2_1496 ( .A(AES_CORE_DATAPATH__abc_16259_n5659_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__6_), .Y(AES_CORE_DATAPATH__abc_16259_n5721) );
  OR2X2 OR2X2_1497 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf6), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_7_), .Y(AES_CORE_DATAPATH__abc_16259_n5723) );
  OR2X2 OR2X2_1498 ( .A(AES_CORE_DATAPATH__abc_16259_n5724), .B(AES_CORE_DATAPATH__abc_16259_n5725), .Y(AES_CORE_DATAPATH__abc_16259_n5726) );
  OR2X2 OR2X2_1499 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf5), .B(AES_CORE_DATAPATH__abc_16259_n5726), .Y(AES_CORE_DATAPATH__abc_16259_n5727) );
  OR2X2 OR2X2_15 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n122), .B(AES_CORE_CONTROL_UNIT__abc_15841_n121), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n123) );
  OR2X2 OR2X2_150 ( .A(AES_CORE_DATAPATH__abc_16259_n2627), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n2628_1) );
  OR2X2 OR2X2_1500 ( .A(AES_CORE_DATAPATH__abc_16259_n5729), .B(AES_CORE_DATAPATH__abc_16259_n5730), .Y(AES_CORE_DATAPATH__0key_3__31_0__7_) );
  OR2X2 OR2X2_1501 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf5), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_8_), .Y(AES_CORE_DATAPATH__abc_16259_n5732) );
  OR2X2 OR2X2_1502 ( .A(AES_CORE_DATAPATH__abc_16259_n5733), .B(AES_CORE_DATAPATH__abc_16259_n5734), .Y(AES_CORE_DATAPATH__abc_16259_n5735) );
  OR2X2 OR2X2_1503 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n5735), .Y(AES_CORE_DATAPATH__abc_16259_n5736) );
  OR2X2 OR2X2_1504 ( .A(AES_CORE_DATAPATH__abc_16259_n5737), .B(AES_CORE_DATAPATH__abc_16259_n5658_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n5738) );
  OR2X2 OR2X2_1505 ( .A(AES_CORE_DATAPATH__abc_16259_n5659_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__8_), .Y(AES_CORE_DATAPATH__abc_16259_n5739) );
  OR2X2 OR2X2_1506 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_9_), .Y(AES_CORE_DATAPATH__abc_16259_n5741) );
  OR2X2 OR2X2_1507 ( .A(AES_CORE_DATAPATH__abc_16259_n5742), .B(AES_CORE_DATAPATH__abc_16259_n5743), .Y(AES_CORE_DATAPATH__abc_16259_n5744) );
  OR2X2 OR2X2_1508 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n5744), .Y(AES_CORE_DATAPATH__abc_16259_n5745) );
  OR2X2 OR2X2_1509 ( .A(AES_CORE_DATAPATH__abc_16259_n5747), .B(AES_CORE_DATAPATH__abc_16259_n5748), .Y(AES_CORE_DATAPATH__0key_3__31_0__9_) );
  OR2X2 OR2X2_151 ( .A(AES_CORE_DATAPATH__abc_16259_n2626_1), .B(AES_CORE_DATAPATH__abc_16259_n2628_1), .Y(AES_CORE_DATAPATH__abc_16259_n2629_1) );
  OR2X2 OR2X2_1510 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_10_), .Y(AES_CORE_DATAPATH__abc_16259_n5750) );
  OR2X2 OR2X2_1511 ( .A(AES_CORE_DATAPATH__abc_16259_n5751), .B(AES_CORE_DATAPATH__abc_16259_n5752), .Y(AES_CORE_DATAPATH__abc_16259_n5753) );
  OR2X2 OR2X2_1512 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n5753), .Y(AES_CORE_DATAPATH__abc_16259_n5754) );
  OR2X2 OR2X2_1513 ( .A(AES_CORE_DATAPATH__abc_16259_n5756), .B(AES_CORE_DATAPATH__abc_16259_n5757), .Y(AES_CORE_DATAPATH__0key_3__31_0__10_) );
  OR2X2 OR2X2_1514 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_11_), .Y(AES_CORE_DATAPATH__abc_16259_n5759) );
  OR2X2 OR2X2_1515 ( .A(AES_CORE_DATAPATH__abc_16259_n5760), .B(AES_CORE_DATAPATH__abc_16259_n5761), .Y(AES_CORE_DATAPATH__abc_16259_n5762) );
  OR2X2 OR2X2_1516 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n5762), .Y(AES_CORE_DATAPATH__abc_16259_n5763) );
  OR2X2 OR2X2_1517 ( .A(AES_CORE_DATAPATH__abc_16259_n5765), .B(AES_CORE_DATAPATH__abc_16259_n5766), .Y(AES_CORE_DATAPATH__0key_3__31_0__11_) );
  OR2X2 OR2X2_1518 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_12_), .Y(AES_CORE_DATAPATH__abc_16259_n5768) );
  OR2X2 OR2X2_1519 ( .A(AES_CORE_DATAPATH__abc_16259_n5769), .B(AES_CORE_DATAPATH__abc_16259_n5770), .Y(AES_CORE_DATAPATH__abc_16259_n5771) );
  OR2X2 OR2X2_152 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf7), .B(AES_CORE_DATAPATH_iv_2__16_), .Y(AES_CORE_DATAPATH__abc_16259_n2630) );
  OR2X2 OR2X2_1520 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n5771), .Y(AES_CORE_DATAPATH__abc_16259_n5772) );
  OR2X2 OR2X2_1521 ( .A(AES_CORE_DATAPATH__abc_16259_n5773), .B(AES_CORE_DATAPATH__abc_16259_n5658_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n5774) );
  OR2X2 OR2X2_1522 ( .A(AES_CORE_DATAPATH__abc_16259_n5659_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__12_), .Y(AES_CORE_DATAPATH__abc_16259_n5775) );
  OR2X2 OR2X2_1523 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_13_), .Y(AES_CORE_DATAPATH__abc_16259_n5777) );
  OR2X2 OR2X2_1524 ( .A(AES_CORE_DATAPATH__abc_16259_n5778), .B(AES_CORE_DATAPATH__abc_16259_n5779), .Y(AES_CORE_DATAPATH__abc_16259_n5780) );
  OR2X2 OR2X2_1525 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf10), .B(AES_CORE_DATAPATH__abc_16259_n5780), .Y(AES_CORE_DATAPATH__abc_16259_n5781) );
  OR2X2 OR2X2_1526 ( .A(AES_CORE_DATAPATH__abc_16259_n5783), .B(AES_CORE_DATAPATH__abc_16259_n5784), .Y(AES_CORE_DATAPATH__0key_3__31_0__13_) );
  OR2X2 OR2X2_1527 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf10), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_14_), .Y(AES_CORE_DATAPATH__abc_16259_n5786) );
  OR2X2 OR2X2_1528 ( .A(AES_CORE_DATAPATH__abc_16259_n5787), .B(AES_CORE_DATAPATH__abc_16259_n5788), .Y(AES_CORE_DATAPATH__abc_16259_n5789) );
  OR2X2 OR2X2_1529 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf9), .B(AES_CORE_DATAPATH__abc_16259_n5789), .Y(AES_CORE_DATAPATH__abc_16259_n5790) );
  OR2X2 OR2X2_153 ( .A(AES_CORE_DATAPATH__abc_16259_n2632), .B(AES_CORE_DATAPATH__abc_16259_n2633_1), .Y(_auto_iopadmap_cc_313_execute_26916_16_) );
  OR2X2 OR2X2_1530 ( .A(AES_CORE_DATAPATH__abc_16259_n5791), .B(AES_CORE_DATAPATH__abc_16259_n5658_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5792) );
  OR2X2 OR2X2_1531 ( .A(AES_CORE_DATAPATH__abc_16259_n5659_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__14_), .Y(AES_CORE_DATAPATH__abc_16259_n5793) );
  OR2X2 OR2X2_1532 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf9), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_15_), .Y(AES_CORE_DATAPATH__abc_16259_n5795) );
  OR2X2 OR2X2_1533 ( .A(AES_CORE_DATAPATH__abc_16259_n5796), .B(AES_CORE_DATAPATH__abc_16259_n5797), .Y(AES_CORE_DATAPATH__abc_16259_n5798) );
  OR2X2 OR2X2_1534 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf8), .B(AES_CORE_DATAPATH__abc_16259_n5798), .Y(AES_CORE_DATAPATH__abc_16259_n5799) );
  OR2X2 OR2X2_1535 ( .A(AES_CORE_DATAPATH__abc_16259_n5801), .B(AES_CORE_DATAPATH__abc_16259_n5802), .Y(AES_CORE_DATAPATH__0key_3__31_0__15_) );
  OR2X2 OR2X2_1536 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf8), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_16_), .Y(AES_CORE_DATAPATH__abc_16259_n5804) );
  OR2X2 OR2X2_1537 ( .A(AES_CORE_DATAPATH__abc_16259_n5805), .B(AES_CORE_DATAPATH__abc_16259_n5806), .Y(AES_CORE_DATAPATH__abc_16259_n5807) );
  OR2X2 OR2X2_1538 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf7), .B(AES_CORE_DATAPATH__abc_16259_n5807), .Y(AES_CORE_DATAPATH__abc_16259_n5808) );
  OR2X2 OR2X2_1539 ( .A(AES_CORE_DATAPATH__abc_16259_n5809), .B(AES_CORE_DATAPATH__abc_16259_n5658_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n5810) );
  OR2X2 OR2X2_154 ( .A(AES_CORE_DATAPATH__abc_16259_n2636_1), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n2637) );
  OR2X2 OR2X2_1540 ( .A(AES_CORE_DATAPATH__abc_16259_n5659_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__16_), .Y(AES_CORE_DATAPATH__abc_16259_n5811) );
  OR2X2 OR2X2_1541 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf7), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_17_), .Y(AES_CORE_DATAPATH__abc_16259_n5813) );
  OR2X2 OR2X2_1542 ( .A(AES_CORE_DATAPATH__abc_16259_n5814), .B(AES_CORE_DATAPATH__abc_16259_n5815), .Y(AES_CORE_DATAPATH__abc_16259_n5816) );
  OR2X2 OR2X2_1543 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf6), .B(AES_CORE_DATAPATH__abc_16259_n5816), .Y(AES_CORE_DATAPATH__abc_16259_n5817) );
  OR2X2 OR2X2_1544 ( .A(AES_CORE_DATAPATH__abc_16259_n5819), .B(AES_CORE_DATAPATH__abc_16259_n5820), .Y(AES_CORE_DATAPATH__0key_3__31_0__17_) );
  OR2X2 OR2X2_1545 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf6), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_18_), .Y(AES_CORE_DATAPATH__abc_16259_n5822) );
  OR2X2 OR2X2_1546 ( .A(AES_CORE_DATAPATH__abc_16259_n5823), .B(AES_CORE_DATAPATH__abc_16259_n5824), .Y(AES_CORE_DATAPATH__abc_16259_n5825) );
  OR2X2 OR2X2_1547 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf5), .B(AES_CORE_DATAPATH__abc_16259_n5825), .Y(AES_CORE_DATAPATH__abc_16259_n5826) );
  OR2X2 OR2X2_1548 ( .A(AES_CORE_DATAPATH__abc_16259_n5828), .B(AES_CORE_DATAPATH__abc_16259_n5829), .Y(AES_CORE_DATAPATH__0key_3__31_0__18_) );
  OR2X2 OR2X2_1549 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf5), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_19_), .Y(AES_CORE_DATAPATH__abc_16259_n5831) );
  OR2X2 OR2X2_155 ( .A(AES_CORE_DATAPATH__abc_16259_n2635), .B(AES_CORE_DATAPATH__abc_16259_n2637), .Y(AES_CORE_DATAPATH__abc_16259_n2638_1) );
  OR2X2 OR2X2_1550 ( .A(AES_CORE_DATAPATH__abc_16259_n5832), .B(AES_CORE_DATAPATH__abc_16259_n5833), .Y(AES_CORE_DATAPATH__abc_16259_n5834) );
  OR2X2 OR2X2_1551 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n5834), .Y(AES_CORE_DATAPATH__abc_16259_n5835) );
  OR2X2 OR2X2_1552 ( .A(AES_CORE_DATAPATH__abc_16259_n5837), .B(AES_CORE_DATAPATH__abc_16259_n5838), .Y(AES_CORE_DATAPATH__0key_3__31_0__19_) );
  OR2X2 OR2X2_1553 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_20_), .Y(AES_CORE_DATAPATH__abc_16259_n5840) );
  OR2X2 OR2X2_1554 ( .A(AES_CORE_DATAPATH__abc_16259_n5841), .B(AES_CORE_DATAPATH__abc_16259_n5842), .Y(AES_CORE_DATAPATH__abc_16259_n5843) );
  OR2X2 OR2X2_1555 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n5843), .Y(AES_CORE_DATAPATH__abc_16259_n5844) );
  OR2X2 OR2X2_1556 ( .A(AES_CORE_DATAPATH__abc_16259_n5846), .B(AES_CORE_DATAPATH__abc_16259_n5847), .Y(AES_CORE_DATAPATH__0key_3__31_0__20_) );
  OR2X2 OR2X2_1557 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_21_), .Y(AES_CORE_DATAPATH__abc_16259_n5849) );
  OR2X2 OR2X2_1558 ( .A(AES_CORE_DATAPATH__abc_16259_n5850), .B(AES_CORE_DATAPATH__abc_16259_n5851), .Y(AES_CORE_DATAPATH__abc_16259_n5852) );
  OR2X2 OR2X2_1559 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n5852), .Y(AES_CORE_DATAPATH__abc_16259_n5853) );
  OR2X2 OR2X2_156 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf6), .B(AES_CORE_DATAPATH_iv_2__17_), .Y(AES_CORE_DATAPATH__abc_16259_n2639_1) );
  OR2X2 OR2X2_1560 ( .A(AES_CORE_DATAPATH__abc_16259_n5854), .B(AES_CORE_DATAPATH__abc_16259_n5658_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n5855) );
  OR2X2 OR2X2_1561 ( .A(AES_CORE_DATAPATH__abc_16259_n5659_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__21_), .Y(AES_CORE_DATAPATH__abc_16259_n5856) );
  OR2X2 OR2X2_1562 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_22_), .Y(AES_CORE_DATAPATH__abc_16259_n5858) );
  OR2X2 OR2X2_1563 ( .A(AES_CORE_DATAPATH__abc_16259_n5859), .B(AES_CORE_DATAPATH__abc_16259_n5860), .Y(AES_CORE_DATAPATH__abc_16259_n5861) );
  OR2X2 OR2X2_1564 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n5861), .Y(AES_CORE_DATAPATH__abc_16259_n5862) );
  OR2X2 OR2X2_1565 ( .A(AES_CORE_DATAPATH__abc_16259_n5864), .B(AES_CORE_DATAPATH__abc_16259_n5865), .Y(AES_CORE_DATAPATH__0key_3__31_0__22_) );
  OR2X2 OR2X2_1566 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_23_), .Y(AES_CORE_DATAPATH__abc_16259_n5867) );
  OR2X2 OR2X2_1567 ( .A(AES_CORE_DATAPATH__abc_16259_n5868), .B(AES_CORE_DATAPATH__abc_16259_n5869), .Y(AES_CORE_DATAPATH__abc_16259_n5870) );
  OR2X2 OR2X2_1568 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n5870), .Y(AES_CORE_DATAPATH__abc_16259_n5871) );
  OR2X2 OR2X2_1569 ( .A(AES_CORE_DATAPATH__abc_16259_n5872), .B(AES_CORE_DATAPATH__abc_16259_n5658_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n5873) );
  OR2X2 OR2X2_157 ( .A(AES_CORE_DATAPATH__abc_16259_n2641_1), .B(AES_CORE_DATAPATH__abc_16259_n2642), .Y(_auto_iopadmap_cc_313_execute_26916_17_) );
  OR2X2 OR2X2_1570 ( .A(AES_CORE_DATAPATH__abc_16259_n5659_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__23_), .Y(AES_CORE_DATAPATH__abc_16259_n5874) );
  OR2X2 OR2X2_1571 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_24_), .Y(AES_CORE_DATAPATH__abc_16259_n5876) );
  OR2X2 OR2X2_1572 ( .A(AES_CORE_DATAPATH__abc_16259_n5877), .B(AES_CORE_DATAPATH__abc_16259_n5878), .Y(AES_CORE_DATAPATH__abc_16259_n5879) );
  OR2X2 OR2X2_1573 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf10), .B(AES_CORE_DATAPATH__abc_16259_n5879), .Y(AES_CORE_DATAPATH__abc_16259_n5880) );
  OR2X2 OR2X2_1574 ( .A(AES_CORE_DATAPATH__abc_16259_n5882), .B(AES_CORE_DATAPATH__abc_16259_n5883), .Y(AES_CORE_DATAPATH__0key_3__31_0__24_) );
  OR2X2 OR2X2_1575 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf10), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_25_), .Y(AES_CORE_DATAPATH__abc_16259_n5885) );
  OR2X2 OR2X2_1576 ( .A(AES_CORE_DATAPATH__abc_16259_n5886), .B(AES_CORE_DATAPATH__abc_16259_n5887), .Y(AES_CORE_DATAPATH__abc_16259_n5888) );
  OR2X2 OR2X2_1577 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf9), .B(AES_CORE_DATAPATH__abc_16259_n5888), .Y(AES_CORE_DATAPATH__abc_16259_n5889) );
  OR2X2 OR2X2_1578 ( .A(AES_CORE_DATAPATH__abc_16259_n5890), .B(AES_CORE_DATAPATH__abc_16259_n5658_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n5891) );
  OR2X2 OR2X2_1579 ( .A(AES_CORE_DATAPATH__abc_16259_n5659_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__25_), .Y(AES_CORE_DATAPATH__abc_16259_n5892) );
  OR2X2 OR2X2_158 ( .A(AES_CORE_DATAPATH__abc_16259_n2645), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n2646_1) );
  OR2X2 OR2X2_1580 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf9), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_26_), .Y(AES_CORE_DATAPATH__abc_16259_n5894) );
  OR2X2 OR2X2_1581 ( .A(AES_CORE_DATAPATH__abc_16259_n5895), .B(AES_CORE_DATAPATH__abc_16259_n5896), .Y(AES_CORE_DATAPATH__abc_16259_n5897) );
  OR2X2 OR2X2_1582 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf8), .B(AES_CORE_DATAPATH__abc_16259_n5897), .Y(AES_CORE_DATAPATH__abc_16259_n5898) );
  OR2X2 OR2X2_1583 ( .A(AES_CORE_DATAPATH__abc_16259_n5900), .B(AES_CORE_DATAPATH__abc_16259_n5901), .Y(AES_CORE_DATAPATH__0key_3__31_0__26_) );
  OR2X2 OR2X2_1584 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf8), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_27_), .Y(AES_CORE_DATAPATH__abc_16259_n5903) );
  OR2X2 OR2X2_1585 ( .A(AES_CORE_DATAPATH__abc_16259_n5904), .B(AES_CORE_DATAPATH__abc_16259_n5905), .Y(AES_CORE_DATAPATH__abc_16259_n5906) );
  OR2X2 OR2X2_1586 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf7), .B(AES_CORE_DATAPATH__abc_16259_n5906), .Y(AES_CORE_DATAPATH__abc_16259_n5907) );
  OR2X2 OR2X2_1587 ( .A(AES_CORE_DATAPATH__abc_16259_n5909), .B(AES_CORE_DATAPATH__abc_16259_n5910), .Y(AES_CORE_DATAPATH__0key_3__31_0__27_) );
  OR2X2 OR2X2_1588 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf7), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_28_), .Y(AES_CORE_DATAPATH__abc_16259_n5912) );
  OR2X2 OR2X2_1589 ( .A(AES_CORE_DATAPATH__abc_16259_n5913), .B(AES_CORE_DATAPATH__abc_16259_n5914), .Y(AES_CORE_DATAPATH__abc_16259_n5915) );
  OR2X2 OR2X2_159 ( .A(AES_CORE_DATAPATH__abc_16259_n2644_1), .B(AES_CORE_DATAPATH__abc_16259_n2646_1), .Y(AES_CORE_DATAPATH__abc_16259_n2647) );
  OR2X2 OR2X2_1590 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf6), .B(AES_CORE_DATAPATH__abc_16259_n5915), .Y(AES_CORE_DATAPATH__abc_16259_n5916) );
  OR2X2 OR2X2_1591 ( .A(AES_CORE_DATAPATH__abc_16259_n5918), .B(AES_CORE_DATAPATH__abc_16259_n5919), .Y(AES_CORE_DATAPATH__0key_3__31_0__28_) );
  OR2X2 OR2X2_1592 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf6), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_29_), .Y(AES_CORE_DATAPATH__abc_16259_n5921) );
  OR2X2 OR2X2_1593 ( .A(AES_CORE_DATAPATH__abc_16259_n5922), .B(AES_CORE_DATAPATH__abc_16259_n5923), .Y(AES_CORE_DATAPATH__abc_16259_n5924) );
  OR2X2 OR2X2_1594 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf5), .B(AES_CORE_DATAPATH__abc_16259_n5924), .Y(AES_CORE_DATAPATH__abc_16259_n5925) );
  OR2X2 OR2X2_1595 ( .A(AES_CORE_DATAPATH__abc_16259_n5927), .B(AES_CORE_DATAPATH__abc_16259_n5928), .Y(AES_CORE_DATAPATH__0key_3__31_0__29_) );
  OR2X2 OR2X2_1596 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf5), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_30_), .Y(AES_CORE_DATAPATH__abc_16259_n5930) );
  OR2X2 OR2X2_1597 ( .A(AES_CORE_DATAPATH__abc_16259_n5931), .B(AES_CORE_DATAPATH__abc_16259_n5932), .Y(AES_CORE_DATAPATH__abc_16259_n5933) );
  OR2X2 OR2X2_1598 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n5933), .Y(AES_CORE_DATAPATH__abc_16259_n5934) );
  OR2X2 OR2X2_1599 ( .A(AES_CORE_DATAPATH__abc_16259_n5936), .B(AES_CORE_DATAPATH__abc_16259_n5937), .Y(AES_CORE_DATAPATH__0key_3__31_0__30_) );
  OR2X2 OR2X2_16 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n124_1), .B(AES_CORE_CONTROL_UNIT__abc_15841_n123), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n125) );
  OR2X2 OR2X2_160 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf5), .B(AES_CORE_DATAPATH_iv_2__18_), .Y(AES_CORE_DATAPATH__abc_16259_n2648_1) );
  OR2X2 OR2X2_1600 ( .A(AES_CORE_DATAPATH__abc_16259_n5939), .B(AES_CORE_DATAPATH__abc_16259_n5940), .Y(AES_CORE_DATAPATH__abc_16259_n5941) );
  OR2X2 OR2X2_1601 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n5941), .Y(AES_CORE_DATAPATH__abc_16259_n5942) );
  OR2X2 OR2X2_1602 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_31_), .Y(AES_CORE_DATAPATH__abc_16259_n5943) );
  OR2X2 OR2X2_1603 ( .A(AES_CORE_DATAPATH__abc_16259_n5945), .B(AES_CORE_DATAPATH__abc_16259_n5946), .Y(AES_CORE_DATAPATH__0key_3__31_0__31_) );
  OR2X2 OR2X2_1604 ( .A(AES_CORE_DATAPATH__abc_16259_n5949), .B(AES_CORE_DATAPATH__abc_16259_n5948), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__0_) );
  OR2X2 OR2X2_1605 ( .A(AES_CORE_DATAPATH__abc_16259_n5672), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n5951) );
  OR2X2 OR2X2_1606 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__1_), .Y(AES_CORE_DATAPATH__abc_16259_n5952) );
  OR2X2 OR2X2_1607 ( .A(AES_CORE_DATAPATH__abc_16259_n5681), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf10), .Y(AES_CORE_DATAPATH__abc_16259_n5954) );
  OR2X2 OR2X2_1608 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__2_), .Y(AES_CORE_DATAPATH__abc_16259_n5955) );
  OR2X2 OR2X2_1609 ( .A(AES_CORE_DATAPATH__abc_16259_n5690), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf9), .Y(AES_CORE_DATAPATH__abc_16259_n5957) );
  OR2X2 OR2X2_161 ( .A(AES_CORE_DATAPATH__abc_16259_n2650), .B(AES_CORE_DATAPATH__abc_16259_n2651_1), .Y(_auto_iopadmap_cc_313_execute_26916_18_) );
  OR2X2 OR2X2_1610 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf10), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__3_), .Y(AES_CORE_DATAPATH__abc_16259_n5958) );
  OR2X2 OR2X2_1611 ( .A(AES_CORE_DATAPATH__abc_16259_n5699), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf8), .Y(AES_CORE_DATAPATH__abc_16259_n5960) );
  OR2X2 OR2X2_1612 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf9), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__4_), .Y(AES_CORE_DATAPATH__abc_16259_n5961) );
  OR2X2 OR2X2_1613 ( .A(AES_CORE_DATAPATH__abc_16259_n5708), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n5963) );
  OR2X2 OR2X2_1614 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf8), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__5_), .Y(AES_CORE_DATAPATH__abc_16259_n5964) );
  OR2X2 OR2X2_1615 ( .A(AES_CORE_DATAPATH__abc_16259_n5717), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n5966) );
  OR2X2 OR2X2_1616 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf7), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__6_), .Y(AES_CORE_DATAPATH__abc_16259_n5967) );
  OR2X2 OR2X2_1617 ( .A(AES_CORE_DATAPATH__abc_16259_n5726), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n5969) );
  OR2X2 OR2X2_1618 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf6), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__7_), .Y(AES_CORE_DATAPATH__abc_16259_n5970) );
  OR2X2 OR2X2_1619 ( .A(AES_CORE_DATAPATH__abc_16259_n5735), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n5972) );
  OR2X2 OR2X2_162 ( .A(AES_CORE_DATAPATH__abc_16259_n2654_1), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n2655) );
  OR2X2 OR2X2_1620 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf5), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__8_), .Y(AES_CORE_DATAPATH__abc_16259_n5973) );
  OR2X2 OR2X2_1621 ( .A(AES_CORE_DATAPATH__abc_16259_n5744), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n5975) );
  OR2X2 OR2X2_1622 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__9_), .Y(AES_CORE_DATAPATH__abc_16259_n5976) );
  OR2X2 OR2X2_1623 ( .A(AES_CORE_DATAPATH__abc_16259_n5753), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n5978) );
  OR2X2 OR2X2_1624 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__10_), .Y(AES_CORE_DATAPATH__abc_16259_n5979) );
  OR2X2 OR2X2_1625 ( .A(AES_CORE_DATAPATH__abc_16259_n5762), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n5981) );
  OR2X2 OR2X2_1626 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__11_), .Y(AES_CORE_DATAPATH__abc_16259_n5982) );
  OR2X2 OR2X2_1627 ( .A(AES_CORE_DATAPATH__abc_16259_n5771), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n5984) );
  OR2X2 OR2X2_1628 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__12_), .Y(AES_CORE_DATAPATH__abc_16259_n5985) );
  OR2X2 OR2X2_1629 ( .A(AES_CORE_DATAPATH__abc_16259_n5780), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf10), .Y(AES_CORE_DATAPATH__abc_16259_n5987) );
  OR2X2 OR2X2_163 ( .A(AES_CORE_DATAPATH__abc_16259_n2653_1), .B(AES_CORE_DATAPATH__abc_16259_n2655), .Y(AES_CORE_DATAPATH__abc_16259_n2656_1) );
  OR2X2 OR2X2_1630 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__13_), .Y(AES_CORE_DATAPATH__abc_16259_n5988) );
  OR2X2 OR2X2_1631 ( .A(AES_CORE_DATAPATH__abc_16259_n5789), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf9), .Y(AES_CORE_DATAPATH__abc_16259_n5990) );
  OR2X2 OR2X2_1632 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf10), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__14_), .Y(AES_CORE_DATAPATH__abc_16259_n5991) );
  OR2X2 OR2X2_1633 ( .A(AES_CORE_DATAPATH__abc_16259_n5798), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf8), .Y(AES_CORE_DATAPATH__abc_16259_n5993) );
  OR2X2 OR2X2_1634 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf9), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__15_), .Y(AES_CORE_DATAPATH__abc_16259_n5994) );
  OR2X2 OR2X2_1635 ( .A(AES_CORE_DATAPATH__abc_16259_n5807), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n5996) );
  OR2X2 OR2X2_1636 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf8), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__16_), .Y(AES_CORE_DATAPATH__abc_16259_n5997) );
  OR2X2 OR2X2_1637 ( .A(AES_CORE_DATAPATH__abc_16259_n5816), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n5999) );
  OR2X2 OR2X2_1638 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf7), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__17_), .Y(AES_CORE_DATAPATH__abc_16259_n6000) );
  OR2X2 OR2X2_1639 ( .A(AES_CORE_DATAPATH__abc_16259_n5825), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n6002) );
  OR2X2 OR2X2_164 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf4), .B(AES_CORE_DATAPATH_iv_2__19_), .Y(AES_CORE_DATAPATH__abc_16259_n2657) );
  OR2X2 OR2X2_1640 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf6), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__18_), .Y(AES_CORE_DATAPATH__abc_16259_n6003) );
  OR2X2 OR2X2_1641 ( .A(AES_CORE_DATAPATH__abc_16259_n5834), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6005) );
  OR2X2 OR2X2_1642 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf5), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__19_), .Y(AES_CORE_DATAPATH__abc_16259_n6006) );
  OR2X2 OR2X2_1643 ( .A(AES_CORE_DATAPATH__abc_16259_n5843), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6008) );
  OR2X2 OR2X2_1644 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__20_), .Y(AES_CORE_DATAPATH__abc_16259_n6009) );
  OR2X2 OR2X2_1645 ( .A(AES_CORE_DATAPATH__abc_16259_n5852), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6011) );
  OR2X2 OR2X2_1646 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__21_), .Y(AES_CORE_DATAPATH__abc_16259_n6012) );
  OR2X2 OR2X2_1647 ( .A(AES_CORE_DATAPATH__abc_16259_n5861), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6014) );
  OR2X2 OR2X2_1648 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__22_), .Y(AES_CORE_DATAPATH__abc_16259_n6015) );
  OR2X2 OR2X2_1649 ( .A(AES_CORE_DATAPATH__abc_16259_n5870), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n6017) );
  OR2X2 OR2X2_165 ( .A(AES_CORE_DATAPATH__abc_16259_n2659), .B(AES_CORE_DATAPATH__abc_16259_n2660), .Y(_auto_iopadmap_cc_313_execute_26916_19_) );
  OR2X2 OR2X2_1650 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__23_), .Y(AES_CORE_DATAPATH__abc_16259_n6018) );
  OR2X2 OR2X2_1651 ( .A(AES_CORE_DATAPATH__abc_16259_n5879), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf10), .Y(AES_CORE_DATAPATH__abc_16259_n6020) );
  OR2X2 OR2X2_1652 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__24_), .Y(AES_CORE_DATAPATH__abc_16259_n6021) );
  OR2X2 OR2X2_1653 ( .A(AES_CORE_DATAPATH__abc_16259_n5888), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf9), .Y(AES_CORE_DATAPATH__abc_16259_n6023) );
  OR2X2 OR2X2_1654 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf10), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__25_), .Y(AES_CORE_DATAPATH__abc_16259_n6024) );
  OR2X2 OR2X2_1655 ( .A(AES_CORE_DATAPATH__abc_16259_n5897), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf8), .Y(AES_CORE_DATAPATH__abc_16259_n6026) );
  OR2X2 OR2X2_1656 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf9), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__26_), .Y(AES_CORE_DATAPATH__abc_16259_n6027) );
  OR2X2 OR2X2_1657 ( .A(AES_CORE_DATAPATH__abc_16259_n5906), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n6029) );
  OR2X2 OR2X2_1658 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf8), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__27_), .Y(AES_CORE_DATAPATH__abc_16259_n6030) );
  OR2X2 OR2X2_1659 ( .A(AES_CORE_DATAPATH__abc_16259_n5915), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n6032) );
  OR2X2 OR2X2_166 ( .A(AES_CORE_DATAPATH__abc_16259_n2663_1), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n2664) );
  OR2X2 OR2X2_1660 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf7), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__28_), .Y(AES_CORE_DATAPATH__abc_16259_n6033) );
  OR2X2 OR2X2_1661 ( .A(AES_CORE_DATAPATH__abc_16259_n5924), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n6035) );
  OR2X2 OR2X2_1662 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf6), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__29_), .Y(AES_CORE_DATAPATH__abc_16259_n6036) );
  OR2X2 OR2X2_1663 ( .A(AES_CORE_DATAPATH__abc_16259_n5933), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6038) );
  OR2X2 OR2X2_1664 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf5), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__30_), .Y(AES_CORE_DATAPATH__abc_16259_n6039) );
  OR2X2 OR2X2_1665 ( .A(AES_CORE_DATAPATH__abc_16259_n4769_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__31_), .Y(AES_CORE_DATAPATH__abc_16259_n6041) );
  OR2X2 OR2X2_1666 ( .A(AES_CORE_DATAPATH__abc_16259_n5941), .B(AES_CORE_CONTROL_UNIT_key_derivation_en_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6042) );
  OR2X2 OR2X2_1667 ( .A(AES_CORE_DATAPATH__abc_16259_n6046), .B(AES_CORE_DATAPATH__abc_16259_n6047), .Y(AES_CORE_DATAPATH__abc_16259_n6048) );
  OR2X2 OR2X2_1668 ( .A(AES_CORE_DATAPATH__abc_16259_n6050), .B(AES_CORE_DATAPATH__abc_16259_n6051), .Y(AES_CORE_DATAPATH__abc_16259_n6052) );
  OR2X2 OR2X2_1669 ( .A(AES_CORE_DATAPATH__abc_16259_n6060), .B(AES_CORE_DATAPATH__abc_16259_n6061), .Y(AES_CORE_DATAPATH__abc_16259_n6062) );
  OR2X2 OR2X2_167 ( .A(AES_CORE_DATAPATH__abc_16259_n2662), .B(AES_CORE_DATAPATH__abc_16259_n2664), .Y(AES_CORE_DATAPATH__abc_16259_n2665_1) );
  OR2X2 OR2X2_1670 ( .A(AES_CORE_DATAPATH__abc_16259_n6066), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n6067) );
  OR2X2 OR2X2_1671 ( .A(AES_CORE_DATAPATH__abc_16259_n6065), .B(AES_CORE_DATAPATH__abc_16259_n6067), .Y(AES_CORE_DATAPATH__abc_16259_n6068) );
  OR2X2 OR2X2_1672 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf7), .B(AES_CORE_DATAPATH_bkp_2__0_), .Y(AES_CORE_DATAPATH__abc_16259_n6069) );
  OR2X2 OR2X2_1673 ( .A(AES_CORE_DATAPATH__abc_16259_n6071), .B(AES_CORE_DATAPATH__abc_16259_n6064), .Y(AES_CORE_DATAPATH__abc_16259_n6072) );
  OR2X2 OR2X2_1674 ( .A(AES_CORE_DATAPATH__abc_16259_n6072), .B(AES_CORE_DATAPATH__abc_16259_n6063_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6073) );
  OR2X2 OR2X2_1675 ( .A(_auto_iopadmap_cc_313_execute_26916_0_), .B(AES_CORE_DATAPATH__abc_16259_n6074_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6075) );
  OR2X2 OR2X2_1676 ( .A(AES_CORE_DATAPATH__abc_16259_n6062), .B(AES_CORE_DATAPATH__abc_16259_n6076), .Y(AES_CORE_DATAPATH__abc_16259_n6077) );
  OR2X2 OR2X2_1677 ( .A(AES_CORE_DATAPATH__abc_16259_n6081), .B(AES_CORE_DATAPATH__abc_16259_n6078), .Y(AES_CORE_DATAPATH__abc_16259_n6082) );
  OR2X2 OR2X2_1678 ( .A(AES_CORE_DATAPATH__abc_16259_n6082), .B(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6083) );
  OR2X2 OR2X2_1679 ( .A(AES_CORE_DATAPATH__abc_16259_n6085), .B(AES_CORE_DATAPATH__abc_16259_n6086), .Y(AES_CORE_DATAPATH__abc_16259_n6087) );
  OR2X2 OR2X2_168 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf3), .B(AES_CORE_DATAPATH_iv_2__20_), .Y(AES_CORE_DATAPATH__abc_16259_n2666) );
  OR2X2 OR2X2_1680 ( .A(AES_CORE_DATAPATH__abc_16259_n6088), .B(AES_CORE_DATAPATH__abc_16259_n6057_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6089) );
  OR2X2 OR2X2_1681 ( .A(_auto_iopadmap_cc_313_execute_26916_0_), .B(AES_CORE_CONTROL_UNIT_last_round_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6090) );
  OR2X2 OR2X2_1682 ( .A(AES_CORE_DATAPATH__abc_16259_n6088), .B(AES_CORE_DATAPATH__abc_16259_n6095_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6096) );
  OR2X2 OR2X2_1683 ( .A(AES_CORE_DATAPATH__abc_16259_n6097_bF_buf4), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_0_), .Y(AES_CORE_DATAPATH__abc_16259_n6098) );
  OR2X2 OR2X2_1684 ( .A(AES_CORE_DATAPATH__abc_16259_n6100), .B(AES_CORE_DATAPATH__abc_16259_n6102), .Y(AES_CORE_DATAPATH__abc_16259_n6103) );
  OR2X2 OR2X2_1685 ( .A(AES_CORE_DATAPATH__abc_16259_n6103), .B(AES_CORE_DATAPATH__abc_16259_n6094), .Y(AES_CORE_DATAPATH__abc_16259_n6104) );
  OR2X2 OR2X2_1686 ( .A(AES_CORE_DATAPATH__abc_16259_n6105), .B(AES_CORE_DATAPATH__abc_16259_n6054), .Y(AES_CORE_DATAPATH__abc_16259_n6106) );
  OR2X2 OR2X2_1687 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf11), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_0_), .Y(AES_CORE_DATAPATH__abc_16259_n6108) );
  OR2X2 OR2X2_1688 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf14), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_64_), .Y(AES_CORE_DATAPATH__abc_16259_n6109) );
  OR2X2 OR2X2_1689 ( .A(AES_CORE_DATAPATH__abc_16259_n6106), .B(AES_CORE_DATAPATH__abc_16259_n6111), .Y(AES_CORE_DATAPATH__abc_16259_n6112) );
  OR2X2 OR2X2_169 ( .A(AES_CORE_DATAPATH__abc_16259_n2668), .B(AES_CORE_DATAPATH__abc_16259_n2669_1), .Y(_auto_iopadmap_cc_313_execute_26916_20_) );
  OR2X2 OR2X2_1690 ( .A(AES_CORE_DATAPATH__abc_16259_n6113), .B(AES_CORE_DATAPATH__abc_16259_n6045), .Y(AES_CORE_DATAPATH__0col_0__31_0__0_) );
  OR2X2 OR2X2_1691 ( .A(AES_CORE_DATAPATH__abc_16259_n2909_1), .B(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6116) );
  OR2X2 OR2X2_1692 ( .A(AES_CORE_DATAPATH__abc_16259_n6059_bF_buf4), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_1_), .Y(AES_CORE_DATAPATH__abc_16259_n6117) );
  OR2X2 OR2X2_1693 ( .A(AES_CORE_DATAPATH__abc_16259_n6120), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n6121) );
  OR2X2 OR2X2_1694 ( .A(AES_CORE_DATAPATH__abc_16259_n6119), .B(AES_CORE_DATAPATH__abc_16259_n6121), .Y(AES_CORE_DATAPATH__abc_16259_n6122) );
  OR2X2 OR2X2_1695 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf6), .B(AES_CORE_DATAPATH_bkp_2__1_), .Y(AES_CORE_DATAPATH__abc_16259_n6123) );
  OR2X2 OR2X2_1696 ( .A(AES_CORE_DATAPATH__abc_16259_n6125), .B(AES_CORE_DATAPATH__abc_16259_n6126), .Y(AES_CORE_DATAPATH__abc_16259_n6127) );
  OR2X2 OR2X2_1697 ( .A(AES_CORE_DATAPATH__abc_16259_n6127), .B(AES_CORE_DATAPATH__abc_16259_n6063_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6128) );
  OR2X2 OR2X2_1698 ( .A(_auto_iopadmap_cc_313_execute_26916_1_), .B(AES_CORE_DATAPATH__abc_16259_n6074_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6129) );
  OR2X2 OR2X2_1699 ( .A(AES_CORE_DATAPATH__abc_16259_n6118), .B(AES_CORE_DATAPATH__abc_16259_n6130), .Y(AES_CORE_DATAPATH__abc_16259_n6131) );
  OR2X2 OR2X2_17 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n128), .B(AES_CORE_CONTROL_UNIT__abc_15841_n127), .Y(AES_CORE_CONTROL_UNIT__abc_10818_n41) );
  OR2X2 OR2X2_170 ( .A(AES_CORE_DATAPATH__abc_16259_n2672), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n2673_1) );
  OR2X2 OR2X2_1700 ( .A(AES_CORE_DATAPATH__abc_16259_n6134), .B(AES_CORE_DATAPATH__abc_16259_n6135), .Y(AES_CORE_DATAPATH__abc_16259_n6136) );
  OR2X2 OR2X2_1701 ( .A(AES_CORE_DATAPATH__abc_16259_n6137), .B(AES_CORE_DATAPATH__abc_16259_n6138), .Y(AES_CORE_DATAPATH__abc_16259_n6139) );
  OR2X2 OR2X2_1702 ( .A(AES_CORE_DATAPATH__abc_16259_n6139), .B(AES_CORE_DATAPATH__abc_16259_n6140), .Y(AES_CORE_DATAPATH__abc_16259_n6141) );
  OR2X2 OR2X2_1703 ( .A(AES_CORE_DATAPATH__abc_16259_n6142), .B(AES_CORE_DATAPATH__abc_16259_n6057_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6143) );
  OR2X2 OR2X2_1704 ( .A(_auto_iopadmap_cc_313_execute_26916_1_), .B(AES_CORE_CONTROL_UNIT_last_round_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6144) );
  OR2X2 OR2X2_1705 ( .A(AES_CORE_DATAPATH__abc_16259_n6142), .B(AES_CORE_DATAPATH__abc_16259_n6095_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6147) );
  OR2X2 OR2X2_1706 ( .A(AES_CORE_DATAPATH__abc_16259_n6097_bF_buf3), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_1_), .Y(AES_CORE_DATAPATH__abc_16259_n6148) );
  OR2X2 OR2X2_1707 ( .A(AES_CORE_DATAPATH__abc_16259_n6150), .B(AES_CORE_DATAPATH__abc_16259_n6151), .Y(AES_CORE_DATAPATH__abc_16259_n6152) );
  OR2X2 OR2X2_1708 ( .A(AES_CORE_DATAPATH__abc_16259_n6152), .B(AES_CORE_DATAPATH__abc_16259_n6146), .Y(AES_CORE_DATAPATH__abc_16259_n6153) );
  OR2X2 OR2X2_1709 ( .A(AES_CORE_DATAPATH__abc_16259_n6154), .B(AES_CORE_DATAPATH__abc_16259_n6155), .Y(AES_CORE_DATAPATH__abc_16259_n6156) );
  OR2X2 OR2X2_171 ( .A(AES_CORE_DATAPATH__abc_16259_n2671_1), .B(AES_CORE_DATAPATH__abc_16259_n2673_1), .Y(AES_CORE_DATAPATH__abc_16259_n2674) );
  OR2X2 OR2X2_1710 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf10), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_1_), .Y(AES_CORE_DATAPATH__abc_16259_n6157) );
  OR2X2 OR2X2_1711 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf13), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_65_), .Y(AES_CORE_DATAPATH__abc_16259_n6158) );
  OR2X2 OR2X2_1712 ( .A(AES_CORE_DATAPATH__abc_16259_n6156), .B(AES_CORE_DATAPATH__abc_16259_n6160), .Y(AES_CORE_DATAPATH__abc_16259_n6161) );
  OR2X2 OR2X2_1713 ( .A(AES_CORE_DATAPATH__abc_16259_n6162), .B(AES_CORE_DATAPATH__abc_16259_n6115), .Y(AES_CORE_DATAPATH__0col_0__31_0__1_) );
  OR2X2 OR2X2_1714 ( .A(AES_CORE_DATAPATH__abc_16259_n6165), .B(AES_CORE_DATAPATH__abc_16259_n6166), .Y(AES_CORE_DATAPATH__abc_16259_n6167) );
  OR2X2 OR2X2_1715 ( .A(AES_CORE_DATAPATH__abc_16259_n6169), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6170) );
  OR2X2 OR2X2_1716 ( .A(AES_CORE_DATAPATH__abc_16259_n6168), .B(AES_CORE_DATAPATH__abc_16259_n6170), .Y(AES_CORE_DATAPATH__abc_16259_n6171) );
  OR2X2 OR2X2_1717 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf5), .B(AES_CORE_DATAPATH_bkp_2__2_), .Y(AES_CORE_DATAPATH__abc_16259_n6172) );
  OR2X2 OR2X2_1718 ( .A(AES_CORE_DATAPATH__abc_16259_n6174), .B(AES_CORE_DATAPATH__abc_16259_n6175), .Y(AES_CORE_DATAPATH__abc_16259_n6176) );
  OR2X2 OR2X2_1719 ( .A(AES_CORE_DATAPATH__abc_16259_n6176), .B(AES_CORE_DATAPATH__abc_16259_n6063_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6177) );
  OR2X2 OR2X2_172 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf2), .B(AES_CORE_DATAPATH_iv_2__21_), .Y(AES_CORE_DATAPATH__abc_16259_n2675_1) );
  OR2X2 OR2X2_1720 ( .A(_auto_iopadmap_cc_313_execute_26916_2_), .B(AES_CORE_DATAPATH__abc_16259_n6074_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6178) );
  OR2X2 OR2X2_1721 ( .A(AES_CORE_DATAPATH__abc_16259_n6167), .B(AES_CORE_DATAPATH__abc_16259_n6179), .Y(AES_CORE_DATAPATH__abc_16259_n6180) );
  OR2X2 OR2X2_1722 ( .A(AES_CORE_DATAPATH__abc_16259_n6183), .B(AES_CORE_DATAPATH__abc_16259_n6184), .Y(AES_CORE_DATAPATH__abc_16259_n6185) );
  OR2X2 OR2X2_1723 ( .A(AES_CORE_DATAPATH__abc_16259_n6185), .B(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6186) );
  OR2X2 OR2X2_1724 ( .A(AES_CORE_DATAPATH__abc_16259_n6188), .B(AES_CORE_DATAPATH__abc_16259_n6189), .Y(AES_CORE_DATAPATH__abc_16259_n6190) );
  OR2X2 OR2X2_1725 ( .A(AES_CORE_DATAPATH__abc_16259_n6191), .B(AES_CORE_DATAPATH__abc_16259_n6057_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6192) );
  OR2X2 OR2X2_1726 ( .A(_auto_iopadmap_cc_313_execute_26916_2_), .B(AES_CORE_CONTROL_UNIT_last_round_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n6193) );
  OR2X2 OR2X2_1727 ( .A(AES_CORE_DATAPATH__abc_16259_n6191), .B(AES_CORE_DATAPATH__abc_16259_n6095_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6196) );
  OR2X2 OR2X2_1728 ( .A(AES_CORE_DATAPATH__abc_16259_n6097_bF_buf2), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_2_), .Y(AES_CORE_DATAPATH__abc_16259_n6197) );
  OR2X2 OR2X2_1729 ( .A(AES_CORE_DATAPATH__abc_16259_n6199), .B(AES_CORE_DATAPATH__abc_16259_n6200), .Y(AES_CORE_DATAPATH__abc_16259_n6201) );
  OR2X2 OR2X2_173 ( .A(AES_CORE_DATAPATH__abc_16259_n2677_1), .B(AES_CORE_DATAPATH__abc_16259_n2678), .Y(_auto_iopadmap_cc_313_execute_26916_21_) );
  OR2X2 OR2X2_1730 ( .A(AES_CORE_DATAPATH__abc_16259_n6201), .B(AES_CORE_DATAPATH__abc_16259_n6195), .Y(AES_CORE_DATAPATH__abc_16259_n6202) );
  OR2X2 OR2X2_1731 ( .A(AES_CORE_DATAPATH__abc_16259_n6203), .B(AES_CORE_DATAPATH__abc_16259_n6204), .Y(AES_CORE_DATAPATH__abc_16259_n6205) );
  OR2X2 OR2X2_1732 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf9), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_2_), .Y(AES_CORE_DATAPATH__abc_16259_n6206) );
  OR2X2 OR2X2_1733 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf12), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_66_), .Y(AES_CORE_DATAPATH__abc_16259_n6207) );
  OR2X2 OR2X2_1734 ( .A(AES_CORE_DATAPATH__abc_16259_n6205), .B(AES_CORE_DATAPATH__abc_16259_n6209), .Y(AES_CORE_DATAPATH__abc_16259_n6210) );
  OR2X2 OR2X2_1735 ( .A(AES_CORE_DATAPATH__abc_16259_n6211), .B(AES_CORE_DATAPATH__abc_16259_n6164), .Y(AES_CORE_DATAPATH__0col_0__31_0__2_) );
  OR2X2 OR2X2_1736 ( .A(AES_CORE_DATAPATH__abc_16259_n6214), .B(AES_CORE_DATAPATH__abc_16259_n6215), .Y(AES_CORE_DATAPATH__abc_16259_n6216) );
  OR2X2 OR2X2_1737 ( .A(AES_CORE_DATAPATH__abc_16259_n6218), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6219) );
  OR2X2 OR2X2_1738 ( .A(AES_CORE_DATAPATH__abc_16259_n6217), .B(AES_CORE_DATAPATH__abc_16259_n6219), .Y(AES_CORE_DATAPATH__abc_16259_n6220) );
  OR2X2 OR2X2_1739 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf4), .B(AES_CORE_DATAPATH_bkp_2__3_), .Y(AES_CORE_DATAPATH__abc_16259_n6221) );
  OR2X2 OR2X2_174 ( .A(AES_CORE_DATAPATH__abc_16259_n2681_1), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n2682) );
  OR2X2 OR2X2_1740 ( .A(AES_CORE_DATAPATH__abc_16259_n6223), .B(AES_CORE_DATAPATH__abc_16259_n6224), .Y(AES_CORE_DATAPATH__abc_16259_n6225) );
  OR2X2 OR2X2_1741 ( .A(AES_CORE_DATAPATH__abc_16259_n6225), .B(AES_CORE_DATAPATH__abc_16259_n6063_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n6226) );
  OR2X2 OR2X2_1742 ( .A(_auto_iopadmap_cc_313_execute_26916_3_), .B(AES_CORE_DATAPATH__abc_16259_n6074_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6227) );
  OR2X2 OR2X2_1743 ( .A(AES_CORE_DATAPATH__abc_16259_n6216), .B(AES_CORE_DATAPATH__abc_16259_n6228), .Y(AES_CORE_DATAPATH__abc_16259_n6229) );
  OR2X2 OR2X2_1744 ( .A(AES_CORE_DATAPATH__abc_16259_n6232), .B(AES_CORE_DATAPATH__abc_16259_n6233), .Y(AES_CORE_DATAPATH__abc_16259_n6234) );
  OR2X2 OR2X2_1745 ( .A(AES_CORE_DATAPATH__abc_16259_n6234), .B(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n6235) );
  OR2X2 OR2X2_1746 ( .A(AES_CORE_DATAPATH__abc_16259_n6237), .B(AES_CORE_DATAPATH__abc_16259_n6238), .Y(AES_CORE_DATAPATH__abc_16259_n6239) );
  OR2X2 OR2X2_1747 ( .A(AES_CORE_DATAPATH__abc_16259_n6240), .B(AES_CORE_DATAPATH__abc_16259_n6057_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n6241) );
  OR2X2 OR2X2_1748 ( .A(_auto_iopadmap_cc_313_execute_26916_3_), .B(AES_CORE_CONTROL_UNIT_last_round_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n6242) );
  OR2X2 OR2X2_1749 ( .A(AES_CORE_DATAPATH__abc_16259_n6240), .B(AES_CORE_DATAPATH__abc_16259_n6095_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n6245) );
  OR2X2 OR2X2_175 ( .A(AES_CORE_DATAPATH__abc_16259_n2680), .B(AES_CORE_DATAPATH__abc_16259_n2682), .Y(AES_CORE_DATAPATH__abc_16259_n2683_1) );
  OR2X2 OR2X2_1750 ( .A(AES_CORE_DATAPATH__abc_16259_n6097_bF_buf1), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_3_), .Y(AES_CORE_DATAPATH__abc_16259_n6246) );
  OR2X2 OR2X2_1751 ( .A(AES_CORE_DATAPATH__abc_16259_n6248), .B(AES_CORE_DATAPATH__abc_16259_n6249), .Y(AES_CORE_DATAPATH__abc_16259_n6250) );
  OR2X2 OR2X2_1752 ( .A(AES_CORE_DATAPATH__abc_16259_n6250), .B(AES_CORE_DATAPATH__abc_16259_n6244), .Y(AES_CORE_DATAPATH__abc_16259_n6251) );
  OR2X2 OR2X2_1753 ( .A(AES_CORE_DATAPATH__abc_16259_n6252), .B(AES_CORE_DATAPATH__abc_16259_n6253), .Y(AES_CORE_DATAPATH__abc_16259_n6254) );
  OR2X2 OR2X2_1754 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf8), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_3_), .Y(AES_CORE_DATAPATH__abc_16259_n6255) );
  OR2X2 OR2X2_1755 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf11), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_67_), .Y(AES_CORE_DATAPATH__abc_16259_n6256) );
  OR2X2 OR2X2_1756 ( .A(AES_CORE_DATAPATH__abc_16259_n6254), .B(AES_CORE_DATAPATH__abc_16259_n6258), .Y(AES_CORE_DATAPATH__abc_16259_n6259) );
  OR2X2 OR2X2_1757 ( .A(AES_CORE_DATAPATH__abc_16259_n6260), .B(AES_CORE_DATAPATH__abc_16259_n6213), .Y(AES_CORE_DATAPATH__0col_0__31_0__3_) );
  OR2X2 OR2X2_1758 ( .A(AES_CORE_DATAPATH__abc_16259_n6263), .B(AES_CORE_DATAPATH__abc_16259_n6264), .Y(AES_CORE_DATAPATH__abc_16259_n6265) );
  OR2X2 OR2X2_1759 ( .A(AES_CORE_DATAPATH__abc_16259_n6267), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6268) );
  OR2X2 OR2X2_176 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf1), .B(AES_CORE_DATAPATH_iv_2__22_), .Y(AES_CORE_DATAPATH__abc_16259_n2684) );
  OR2X2 OR2X2_1760 ( .A(AES_CORE_DATAPATH__abc_16259_n6266), .B(AES_CORE_DATAPATH__abc_16259_n6268), .Y(AES_CORE_DATAPATH__abc_16259_n6269) );
  OR2X2 OR2X2_1761 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf3), .B(AES_CORE_DATAPATH_bkp_2__4_), .Y(AES_CORE_DATAPATH__abc_16259_n6270) );
  OR2X2 OR2X2_1762 ( .A(AES_CORE_DATAPATH__abc_16259_n6272), .B(AES_CORE_DATAPATH__abc_16259_n6273), .Y(AES_CORE_DATAPATH__abc_16259_n6274) );
  OR2X2 OR2X2_1763 ( .A(AES_CORE_DATAPATH__abc_16259_n6274), .B(AES_CORE_DATAPATH__abc_16259_n6063_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6275) );
  OR2X2 OR2X2_1764 ( .A(_auto_iopadmap_cc_313_execute_26916_4_), .B(AES_CORE_DATAPATH__abc_16259_n6074_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n6276) );
  OR2X2 OR2X2_1765 ( .A(AES_CORE_DATAPATH__abc_16259_n6265), .B(AES_CORE_DATAPATH__abc_16259_n6277), .Y(AES_CORE_DATAPATH__abc_16259_n6278) );
  OR2X2 OR2X2_1766 ( .A(AES_CORE_DATAPATH__abc_16259_n6281), .B(AES_CORE_DATAPATH__abc_16259_n6282), .Y(AES_CORE_DATAPATH__abc_16259_n6283) );
  OR2X2 OR2X2_1767 ( .A(AES_CORE_DATAPATH__abc_16259_n6283), .B(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6284) );
  OR2X2 OR2X2_1768 ( .A(AES_CORE_DATAPATH__abc_16259_n6286), .B(AES_CORE_DATAPATH__abc_16259_n6287), .Y(AES_CORE_DATAPATH__abc_16259_n6288) );
  OR2X2 OR2X2_1769 ( .A(AES_CORE_DATAPATH__abc_16259_n6289), .B(AES_CORE_DATAPATH__abc_16259_n6057_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6290) );
  OR2X2 OR2X2_177 ( .A(AES_CORE_DATAPATH__abc_16259_n2686), .B(AES_CORE_DATAPATH__abc_16259_n2687_1), .Y(_auto_iopadmap_cc_313_execute_26916_22_) );
  OR2X2 OR2X2_1770 ( .A(_auto_iopadmap_cc_313_execute_26916_4_), .B(AES_CORE_CONTROL_UNIT_last_round_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6291) );
  OR2X2 OR2X2_1771 ( .A(AES_CORE_DATAPATH__abc_16259_n6289), .B(AES_CORE_DATAPATH__abc_16259_n6095_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6294) );
  OR2X2 OR2X2_1772 ( .A(AES_CORE_DATAPATH__abc_16259_n6097_bF_buf0), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_4_), .Y(AES_CORE_DATAPATH__abc_16259_n6295) );
  OR2X2 OR2X2_1773 ( .A(AES_CORE_DATAPATH__abc_16259_n6297), .B(AES_CORE_DATAPATH__abc_16259_n6298), .Y(AES_CORE_DATAPATH__abc_16259_n6299) );
  OR2X2 OR2X2_1774 ( .A(AES_CORE_DATAPATH__abc_16259_n6299), .B(AES_CORE_DATAPATH__abc_16259_n6293), .Y(AES_CORE_DATAPATH__abc_16259_n6300) );
  OR2X2 OR2X2_1775 ( .A(AES_CORE_DATAPATH__abc_16259_n6301), .B(AES_CORE_DATAPATH__abc_16259_n6302), .Y(AES_CORE_DATAPATH__abc_16259_n6303) );
  OR2X2 OR2X2_1776 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf7), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_4_), .Y(AES_CORE_DATAPATH__abc_16259_n6304) );
  OR2X2 OR2X2_1777 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf10), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_68_), .Y(AES_CORE_DATAPATH__abc_16259_n6305) );
  OR2X2 OR2X2_1778 ( .A(AES_CORE_DATAPATH__abc_16259_n6303), .B(AES_CORE_DATAPATH__abc_16259_n6307), .Y(AES_CORE_DATAPATH__abc_16259_n6308) );
  OR2X2 OR2X2_1779 ( .A(AES_CORE_DATAPATH__abc_16259_n6309), .B(AES_CORE_DATAPATH__abc_16259_n6262), .Y(AES_CORE_DATAPATH__0col_0__31_0__4_) );
  OR2X2 OR2X2_178 ( .A(AES_CORE_DATAPATH__abc_16259_n2690), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n2691_1) );
  OR2X2 OR2X2_1780 ( .A(AES_CORE_DATAPATH__abc_16259_n6312), .B(AES_CORE_DATAPATH__abc_16259_n6313), .Y(AES_CORE_DATAPATH__abc_16259_n6314) );
  OR2X2 OR2X2_1781 ( .A(AES_CORE_DATAPATH__abc_16259_n6316), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6317) );
  OR2X2 OR2X2_1782 ( .A(AES_CORE_DATAPATH__abc_16259_n6315), .B(AES_CORE_DATAPATH__abc_16259_n6317), .Y(AES_CORE_DATAPATH__abc_16259_n6318) );
  OR2X2 OR2X2_1783 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf2), .B(AES_CORE_DATAPATH_bkp_2__5_), .Y(AES_CORE_DATAPATH__abc_16259_n6319) );
  OR2X2 OR2X2_1784 ( .A(AES_CORE_DATAPATH__abc_16259_n6321), .B(AES_CORE_DATAPATH__abc_16259_n6322), .Y(AES_CORE_DATAPATH__abc_16259_n6323) );
  OR2X2 OR2X2_1785 ( .A(AES_CORE_DATAPATH__abc_16259_n6323), .B(AES_CORE_DATAPATH__abc_16259_n6063_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6324) );
  OR2X2 OR2X2_1786 ( .A(_auto_iopadmap_cc_313_execute_26916_5_), .B(AES_CORE_DATAPATH__abc_16259_n6074_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6325) );
  OR2X2 OR2X2_1787 ( .A(AES_CORE_DATAPATH__abc_16259_n6314), .B(AES_CORE_DATAPATH__abc_16259_n6326), .Y(AES_CORE_DATAPATH__abc_16259_n6327) );
  OR2X2 OR2X2_1788 ( .A(AES_CORE_DATAPATH__abc_16259_n6330), .B(AES_CORE_DATAPATH__abc_16259_n6331), .Y(AES_CORE_DATAPATH__abc_16259_n6332) );
  OR2X2 OR2X2_1789 ( .A(AES_CORE_DATAPATH__abc_16259_n6332), .B(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6333) );
  OR2X2 OR2X2_179 ( .A(AES_CORE_DATAPATH__abc_16259_n2689_1), .B(AES_CORE_DATAPATH__abc_16259_n2691_1), .Y(AES_CORE_DATAPATH__abc_16259_n2692) );
  OR2X2 OR2X2_1790 ( .A(AES_CORE_DATAPATH__abc_16259_n6335), .B(AES_CORE_DATAPATH__abc_16259_n6336), .Y(AES_CORE_DATAPATH__abc_16259_n6337) );
  OR2X2 OR2X2_1791 ( .A(AES_CORE_DATAPATH__abc_16259_n6338), .B(AES_CORE_DATAPATH__abc_16259_n6057_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6339) );
  OR2X2 OR2X2_1792 ( .A(_auto_iopadmap_cc_313_execute_26916_5_), .B(AES_CORE_CONTROL_UNIT_last_round_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6340) );
  OR2X2 OR2X2_1793 ( .A(AES_CORE_DATAPATH__abc_16259_n6338), .B(AES_CORE_DATAPATH__abc_16259_n6095_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6343) );
  OR2X2 OR2X2_1794 ( .A(AES_CORE_DATAPATH__abc_16259_n6097_bF_buf4), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_5_), .Y(AES_CORE_DATAPATH__abc_16259_n6344) );
  OR2X2 OR2X2_1795 ( .A(AES_CORE_DATAPATH__abc_16259_n6346), .B(AES_CORE_DATAPATH__abc_16259_n6347), .Y(AES_CORE_DATAPATH__abc_16259_n6348) );
  OR2X2 OR2X2_1796 ( .A(AES_CORE_DATAPATH__abc_16259_n6348), .B(AES_CORE_DATAPATH__abc_16259_n6342), .Y(AES_CORE_DATAPATH__abc_16259_n6349) );
  OR2X2 OR2X2_1797 ( .A(AES_CORE_DATAPATH__abc_16259_n6350), .B(AES_CORE_DATAPATH__abc_16259_n6351), .Y(AES_CORE_DATAPATH__abc_16259_n6352) );
  OR2X2 OR2X2_1798 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf6), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_5_), .Y(AES_CORE_DATAPATH__abc_16259_n6353) );
  OR2X2 OR2X2_1799 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf9), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_69_), .Y(AES_CORE_DATAPATH__abc_16259_n6354) );
  OR2X2 OR2X2_18 ( .A(disable_core), .B(_auto_iopadmap_cc_313_execute_26914), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n130_1) );
  OR2X2 OR2X2_180 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf0), .B(AES_CORE_DATAPATH_iv_2__23_), .Y(AES_CORE_DATAPATH__abc_16259_n2693_1) );
  OR2X2 OR2X2_1800 ( .A(AES_CORE_DATAPATH__abc_16259_n6352), .B(AES_CORE_DATAPATH__abc_16259_n6356), .Y(AES_CORE_DATAPATH__abc_16259_n6357) );
  OR2X2 OR2X2_1801 ( .A(AES_CORE_DATAPATH__abc_16259_n6358), .B(AES_CORE_DATAPATH__abc_16259_n6311), .Y(AES_CORE_DATAPATH__0col_0__31_0__5_) );
  OR2X2 OR2X2_1802 ( .A(AES_CORE_DATAPATH__abc_16259_n6361), .B(AES_CORE_DATAPATH__abc_16259_n6362), .Y(AES_CORE_DATAPATH__abc_16259_n6363) );
  OR2X2 OR2X2_1803 ( .A(AES_CORE_DATAPATH__abc_16259_n6365), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n6366) );
  OR2X2 OR2X2_1804 ( .A(AES_CORE_DATAPATH__abc_16259_n6364), .B(AES_CORE_DATAPATH__abc_16259_n6366), .Y(AES_CORE_DATAPATH__abc_16259_n6367) );
  OR2X2 OR2X2_1805 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf1), .B(AES_CORE_DATAPATH_bkp_2__6_), .Y(AES_CORE_DATAPATH__abc_16259_n6368) );
  OR2X2 OR2X2_1806 ( .A(AES_CORE_DATAPATH__abc_16259_n6370), .B(AES_CORE_DATAPATH__abc_16259_n6371), .Y(AES_CORE_DATAPATH__abc_16259_n6372) );
  OR2X2 OR2X2_1807 ( .A(AES_CORE_DATAPATH__abc_16259_n6372), .B(AES_CORE_DATAPATH__abc_16259_n6063_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6373) );
  OR2X2 OR2X2_1808 ( .A(_auto_iopadmap_cc_313_execute_26916_6_), .B(AES_CORE_DATAPATH__abc_16259_n6074_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6374) );
  OR2X2 OR2X2_1809 ( .A(AES_CORE_DATAPATH__abc_16259_n6363), .B(AES_CORE_DATAPATH__abc_16259_n6375), .Y(AES_CORE_DATAPATH__abc_16259_n6376) );
  OR2X2 OR2X2_181 ( .A(AES_CORE_DATAPATH__abc_16259_n2695_1), .B(AES_CORE_DATAPATH__abc_16259_n2696), .Y(_auto_iopadmap_cc_313_execute_26916_23_) );
  OR2X2 OR2X2_1810 ( .A(AES_CORE_DATAPATH__abc_16259_n6379), .B(AES_CORE_DATAPATH__abc_16259_n6380), .Y(AES_CORE_DATAPATH__abc_16259_n6381) );
  OR2X2 OR2X2_1811 ( .A(AES_CORE_DATAPATH__abc_16259_n6381), .B(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n6382) );
  OR2X2 OR2X2_1812 ( .A(AES_CORE_DATAPATH__abc_16259_n6384), .B(AES_CORE_DATAPATH__abc_16259_n6385), .Y(AES_CORE_DATAPATH__abc_16259_n6386) );
  OR2X2 OR2X2_1813 ( .A(AES_CORE_DATAPATH__abc_16259_n6387), .B(AES_CORE_DATAPATH__abc_16259_n6057_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6388) );
  OR2X2 OR2X2_1814 ( .A(_auto_iopadmap_cc_313_execute_26916_6_), .B(AES_CORE_CONTROL_UNIT_last_round_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6389) );
  OR2X2 OR2X2_1815 ( .A(AES_CORE_DATAPATH__abc_16259_n6387), .B(AES_CORE_DATAPATH__abc_16259_n6095_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6392) );
  OR2X2 OR2X2_1816 ( .A(AES_CORE_DATAPATH__abc_16259_n6097_bF_buf3), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_6_), .Y(AES_CORE_DATAPATH__abc_16259_n6393) );
  OR2X2 OR2X2_1817 ( .A(AES_CORE_DATAPATH__abc_16259_n6395), .B(AES_CORE_DATAPATH__abc_16259_n6396), .Y(AES_CORE_DATAPATH__abc_16259_n6397) );
  OR2X2 OR2X2_1818 ( .A(AES_CORE_DATAPATH__abc_16259_n6397), .B(AES_CORE_DATAPATH__abc_16259_n6391), .Y(AES_CORE_DATAPATH__abc_16259_n6398) );
  OR2X2 OR2X2_1819 ( .A(AES_CORE_DATAPATH__abc_16259_n6399), .B(AES_CORE_DATAPATH__abc_16259_n6400), .Y(AES_CORE_DATAPATH__abc_16259_n6401) );
  OR2X2 OR2X2_182 ( .A(AES_CORE_DATAPATH__abc_16259_n2699_1), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n2700) );
  OR2X2 OR2X2_1820 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf5), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_6_), .Y(AES_CORE_DATAPATH__abc_16259_n6402) );
  OR2X2 OR2X2_1821 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf8), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_70_), .Y(AES_CORE_DATAPATH__abc_16259_n6403) );
  OR2X2 OR2X2_1822 ( .A(AES_CORE_DATAPATH__abc_16259_n6401), .B(AES_CORE_DATAPATH__abc_16259_n6405), .Y(AES_CORE_DATAPATH__abc_16259_n6406) );
  OR2X2 OR2X2_1823 ( .A(AES_CORE_DATAPATH__abc_16259_n6407), .B(AES_CORE_DATAPATH__abc_16259_n6360), .Y(AES_CORE_DATAPATH__0col_0__31_0__6_) );
  OR2X2 OR2X2_1824 ( .A(AES_CORE_DATAPATH__abc_16259_n6410), .B(AES_CORE_DATAPATH__abc_16259_n6411), .Y(AES_CORE_DATAPATH__abc_16259_n6412) );
  OR2X2 OR2X2_1825 ( .A(AES_CORE_DATAPATH__abc_16259_n6414), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n6415) );
  OR2X2 OR2X2_1826 ( .A(AES_CORE_DATAPATH__abc_16259_n6413), .B(AES_CORE_DATAPATH__abc_16259_n6415), .Y(AES_CORE_DATAPATH__abc_16259_n6416) );
  OR2X2 OR2X2_1827 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf0), .B(AES_CORE_DATAPATH_bkp_2__7_), .Y(AES_CORE_DATAPATH__abc_16259_n6417) );
  OR2X2 OR2X2_1828 ( .A(AES_CORE_DATAPATH__abc_16259_n6419), .B(AES_CORE_DATAPATH__abc_16259_n6420), .Y(AES_CORE_DATAPATH__abc_16259_n6421) );
  OR2X2 OR2X2_1829 ( .A(AES_CORE_DATAPATH__abc_16259_n6421), .B(AES_CORE_DATAPATH__abc_16259_n6063_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6422) );
  OR2X2 OR2X2_183 ( .A(AES_CORE_DATAPATH__abc_16259_n2698), .B(AES_CORE_DATAPATH__abc_16259_n2700), .Y(AES_CORE_DATAPATH__abc_16259_n2701_1) );
  OR2X2 OR2X2_1830 ( .A(_auto_iopadmap_cc_313_execute_26916_7_), .B(AES_CORE_DATAPATH__abc_16259_n6074_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6423) );
  OR2X2 OR2X2_1831 ( .A(AES_CORE_DATAPATH__abc_16259_n6412), .B(AES_CORE_DATAPATH__abc_16259_n6424), .Y(AES_CORE_DATAPATH__abc_16259_n6425) );
  OR2X2 OR2X2_1832 ( .A(AES_CORE_DATAPATH__abc_16259_n6428), .B(AES_CORE_DATAPATH__abc_16259_n6429), .Y(AES_CORE_DATAPATH__abc_16259_n6430) );
  OR2X2 OR2X2_1833 ( .A(AES_CORE_DATAPATH__abc_16259_n6430), .B(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n6431) );
  OR2X2 OR2X2_1834 ( .A(AES_CORE_DATAPATH__abc_16259_n6433), .B(AES_CORE_DATAPATH__abc_16259_n6434), .Y(AES_CORE_DATAPATH__abc_16259_n6435) );
  OR2X2 OR2X2_1835 ( .A(AES_CORE_DATAPATH__abc_16259_n6436), .B(AES_CORE_DATAPATH__abc_16259_n6057_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6437) );
  OR2X2 OR2X2_1836 ( .A(_auto_iopadmap_cc_313_execute_26916_7_), .B(AES_CORE_CONTROL_UNIT_last_round_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6438) );
  OR2X2 OR2X2_1837 ( .A(AES_CORE_DATAPATH__abc_16259_n6436), .B(AES_CORE_DATAPATH__abc_16259_n6095_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6441) );
  OR2X2 OR2X2_1838 ( .A(AES_CORE_DATAPATH__abc_16259_n6097_bF_buf2), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_7_), .Y(AES_CORE_DATAPATH__abc_16259_n6442) );
  OR2X2 OR2X2_1839 ( .A(AES_CORE_DATAPATH__abc_16259_n6444), .B(AES_CORE_DATAPATH__abc_16259_n6445), .Y(AES_CORE_DATAPATH__abc_16259_n6446) );
  OR2X2 OR2X2_184 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf7), .B(AES_CORE_DATAPATH_iv_2__24_), .Y(AES_CORE_DATAPATH__abc_16259_n2702) );
  OR2X2 OR2X2_1840 ( .A(AES_CORE_DATAPATH__abc_16259_n6446), .B(AES_CORE_DATAPATH__abc_16259_n6440), .Y(AES_CORE_DATAPATH__abc_16259_n6447) );
  OR2X2 OR2X2_1841 ( .A(AES_CORE_DATAPATH__abc_16259_n6448), .B(AES_CORE_DATAPATH__abc_16259_n6449), .Y(AES_CORE_DATAPATH__abc_16259_n6450) );
  OR2X2 OR2X2_1842 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf4), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_7_), .Y(AES_CORE_DATAPATH__abc_16259_n6451) );
  OR2X2 OR2X2_1843 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf7), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_71_), .Y(AES_CORE_DATAPATH__abc_16259_n6452) );
  OR2X2 OR2X2_1844 ( .A(AES_CORE_DATAPATH__abc_16259_n6450), .B(AES_CORE_DATAPATH__abc_16259_n6454), .Y(AES_CORE_DATAPATH__abc_16259_n6455) );
  OR2X2 OR2X2_1845 ( .A(AES_CORE_DATAPATH__abc_16259_n6456), .B(AES_CORE_DATAPATH__abc_16259_n6409), .Y(AES_CORE_DATAPATH__0col_0__31_0__7_) );
  OR2X2 OR2X2_1846 ( .A(AES_CORE_DATAPATH__abc_16259_n6459), .B(AES_CORE_DATAPATH__abc_16259_n6460), .Y(AES_CORE_DATAPATH__abc_16259_n6461) );
  OR2X2 OR2X2_1847 ( .A(AES_CORE_DATAPATH__abc_16259_n6463), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n6464) );
  OR2X2 OR2X2_1848 ( .A(AES_CORE_DATAPATH__abc_16259_n6462), .B(AES_CORE_DATAPATH__abc_16259_n6464), .Y(AES_CORE_DATAPATH__abc_16259_n6465) );
  OR2X2 OR2X2_1849 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf7), .B(AES_CORE_DATAPATH_bkp_2__8_), .Y(AES_CORE_DATAPATH__abc_16259_n6466) );
  OR2X2 OR2X2_185 ( .A(AES_CORE_DATAPATH__abc_16259_n2704), .B(AES_CORE_DATAPATH__abc_16259_n2705_1), .Y(_auto_iopadmap_cc_313_execute_26916_24_) );
  OR2X2 OR2X2_1850 ( .A(AES_CORE_DATAPATH__abc_16259_n6468), .B(AES_CORE_DATAPATH__abc_16259_n6469), .Y(AES_CORE_DATAPATH__abc_16259_n6470) );
  OR2X2 OR2X2_1851 ( .A(AES_CORE_DATAPATH__abc_16259_n6470), .B(AES_CORE_DATAPATH__abc_16259_n6063_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n6471) );
  OR2X2 OR2X2_1852 ( .A(_auto_iopadmap_cc_313_execute_26916_8_), .B(AES_CORE_DATAPATH__abc_16259_n6074_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6472) );
  OR2X2 OR2X2_1853 ( .A(AES_CORE_DATAPATH__abc_16259_n6461), .B(AES_CORE_DATAPATH__abc_16259_n6473), .Y(AES_CORE_DATAPATH__abc_16259_n6474) );
  OR2X2 OR2X2_1854 ( .A(AES_CORE_DATAPATH__abc_16259_n6477), .B(AES_CORE_DATAPATH__abc_16259_n6478), .Y(AES_CORE_DATAPATH__abc_16259_n6479) );
  OR2X2 OR2X2_1855 ( .A(AES_CORE_DATAPATH__abc_16259_n6479), .B(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6480) );
  OR2X2 OR2X2_1856 ( .A(AES_CORE_DATAPATH__abc_16259_n6482), .B(AES_CORE_DATAPATH__abc_16259_n6483), .Y(AES_CORE_DATAPATH__abc_16259_n6484) );
  OR2X2 OR2X2_1857 ( .A(AES_CORE_DATAPATH__abc_16259_n6485), .B(AES_CORE_DATAPATH__abc_16259_n6057_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n6486) );
  OR2X2 OR2X2_1858 ( .A(_auto_iopadmap_cc_313_execute_26916_8_), .B(AES_CORE_CONTROL_UNIT_last_round_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n6487) );
  OR2X2 OR2X2_1859 ( .A(AES_CORE_DATAPATH__abc_16259_n6485), .B(AES_CORE_DATAPATH__abc_16259_n6095_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n6490) );
  OR2X2 OR2X2_186 ( .A(AES_CORE_DATAPATH__abc_16259_n2708), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n2709_1) );
  OR2X2 OR2X2_1860 ( .A(AES_CORE_DATAPATH__abc_16259_n6097_bF_buf1), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_8_), .Y(AES_CORE_DATAPATH__abc_16259_n6491) );
  OR2X2 OR2X2_1861 ( .A(AES_CORE_DATAPATH__abc_16259_n6493), .B(AES_CORE_DATAPATH__abc_16259_n6494), .Y(AES_CORE_DATAPATH__abc_16259_n6495) );
  OR2X2 OR2X2_1862 ( .A(AES_CORE_DATAPATH__abc_16259_n6495), .B(AES_CORE_DATAPATH__abc_16259_n6489), .Y(AES_CORE_DATAPATH__abc_16259_n6496) );
  OR2X2 OR2X2_1863 ( .A(AES_CORE_DATAPATH__abc_16259_n6497), .B(AES_CORE_DATAPATH__abc_16259_n6498), .Y(AES_CORE_DATAPATH__abc_16259_n6499) );
  OR2X2 OR2X2_1864 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf3), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_40_), .Y(AES_CORE_DATAPATH__abc_16259_n6500) );
  OR2X2 OR2X2_1865 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf6), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_40_), .Y(AES_CORE_DATAPATH__abc_16259_n6501) );
  OR2X2 OR2X2_1866 ( .A(AES_CORE_DATAPATH__abc_16259_n6499), .B(AES_CORE_DATAPATH__abc_16259_n6503), .Y(AES_CORE_DATAPATH__abc_16259_n6504) );
  OR2X2 OR2X2_1867 ( .A(AES_CORE_DATAPATH__abc_16259_n6505), .B(AES_CORE_DATAPATH__abc_16259_n6458), .Y(AES_CORE_DATAPATH__0col_0__31_0__8_) );
  OR2X2 OR2X2_1868 ( .A(AES_CORE_DATAPATH__abc_16259_n6508), .B(AES_CORE_DATAPATH__abc_16259_n6509), .Y(AES_CORE_DATAPATH__abc_16259_n6510) );
  OR2X2 OR2X2_1869 ( .A(AES_CORE_DATAPATH__abc_16259_n6512), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n6513) );
  OR2X2 OR2X2_187 ( .A(AES_CORE_DATAPATH__abc_16259_n2707_1), .B(AES_CORE_DATAPATH__abc_16259_n2709_1), .Y(AES_CORE_DATAPATH__abc_16259_n2710) );
  OR2X2 OR2X2_1870 ( .A(AES_CORE_DATAPATH__abc_16259_n6511), .B(AES_CORE_DATAPATH__abc_16259_n6513), .Y(AES_CORE_DATAPATH__abc_16259_n6514) );
  OR2X2 OR2X2_1871 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf6), .B(AES_CORE_DATAPATH_bkp_2__9_), .Y(AES_CORE_DATAPATH__abc_16259_n6515) );
  OR2X2 OR2X2_1872 ( .A(AES_CORE_DATAPATH__abc_16259_n6517), .B(AES_CORE_DATAPATH__abc_16259_n6518), .Y(AES_CORE_DATAPATH__abc_16259_n6519) );
  OR2X2 OR2X2_1873 ( .A(AES_CORE_DATAPATH__abc_16259_n6519), .B(AES_CORE_DATAPATH__abc_16259_n6063_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6520) );
  OR2X2 OR2X2_1874 ( .A(_auto_iopadmap_cc_313_execute_26916_9_), .B(AES_CORE_DATAPATH__abc_16259_n6074_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n6521) );
  OR2X2 OR2X2_1875 ( .A(AES_CORE_DATAPATH__abc_16259_n6510), .B(AES_CORE_DATAPATH__abc_16259_n6522), .Y(AES_CORE_DATAPATH__abc_16259_n6523) );
  OR2X2 OR2X2_1876 ( .A(AES_CORE_DATAPATH__abc_16259_n6526), .B(AES_CORE_DATAPATH__abc_16259_n6527), .Y(AES_CORE_DATAPATH__abc_16259_n6528) );
  OR2X2 OR2X2_1877 ( .A(AES_CORE_DATAPATH__abc_16259_n6528), .B(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6529) );
  OR2X2 OR2X2_1878 ( .A(AES_CORE_DATAPATH__abc_16259_n6531), .B(AES_CORE_DATAPATH__abc_16259_n6532), .Y(AES_CORE_DATAPATH__abc_16259_n6533) );
  OR2X2 OR2X2_1879 ( .A(AES_CORE_DATAPATH__abc_16259_n6534), .B(AES_CORE_DATAPATH__abc_16259_n6057_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6535) );
  OR2X2 OR2X2_188 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf6), .B(AES_CORE_DATAPATH_iv_2__25_), .Y(AES_CORE_DATAPATH__abc_16259_n2711_1) );
  OR2X2 OR2X2_1880 ( .A(_auto_iopadmap_cc_313_execute_26916_9_), .B(AES_CORE_CONTROL_UNIT_last_round_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n6536) );
  OR2X2 OR2X2_1881 ( .A(AES_CORE_DATAPATH__abc_16259_n6534), .B(AES_CORE_DATAPATH__abc_16259_n6095_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6539) );
  OR2X2 OR2X2_1882 ( .A(AES_CORE_DATAPATH__abc_16259_n6097_bF_buf0), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_9_), .Y(AES_CORE_DATAPATH__abc_16259_n6540) );
  OR2X2 OR2X2_1883 ( .A(AES_CORE_DATAPATH__abc_16259_n6542), .B(AES_CORE_DATAPATH__abc_16259_n6543), .Y(AES_CORE_DATAPATH__abc_16259_n6544) );
  OR2X2 OR2X2_1884 ( .A(AES_CORE_DATAPATH__abc_16259_n6544), .B(AES_CORE_DATAPATH__abc_16259_n6538), .Y(AES_CORE_DATAPATH__abc_16259_n6545) );
  OR2X2 OR2X2_1885 ( .A(AES_CORE_DATAPATH__abc_16259_n6546), .B(AES_CORE_DATAPATH__abc_16259_n6547), .Y(AES_CORE_DATAPATH__abc_16259_n6548) );
  OR2X2 OR2X2_1886 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf2), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_41_), .Y(AES_CORE_DATAPATH__abc_16259_n6549) );
  OR2X2 OR2X2_1887 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf5), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_41_), .Y(AES_CORE_DATAPATH__abc_16259_n6550) );
  OR2X2 OR2X2_1888 ( .A(AES_CORE_DATAPATH__abc_16259_n6548), .B(AES_CORE_DATAPATH__abc_16259_n6552), .Y(AES_CORE_DATAPATH__abc_16259_n6553) );
  OR2X2 OR2X2_1889 ( .A(AES_CORE_DATAPATH__abc_16259_n6554), .B(AES_CORE_DATAPATH__abc_16259_n6507), .Y(AES_CORE_DATAPATH__0col_0__31_0__9_) );
  OR2X2 OR2X2_189 ( .A(AES_CORE_DATAPATH__abc_16259_n2713_1), .B(AES_CORE_DATAPATH__abc_16259_n2714), .Y(_auto_iopadmap_cc_313_execute_26916_25_) );
  OR2X2 OR2X2_1890 ( .A(AES_CORE_DATAPATH__abc_16259_n6559), .B(AES_CORE_DATAPATH__abc_16259_n6560), .Y(AES_CORE_DATAPATH__abc_16259_n6561) );
  OR2X2 OR2X2_1891 ( .A(AES_CORE_DATAPATH__abc_16259_n6562), .B(AES_CORE_DATAPATH__abc_16259_n6564), .Y(AES_CORE_DATAPATH__abc_16259_n6565) );
  OR2X2 OR2X2_1892 ( .A(AES_CORE_DATAPATH__abc_16259_n6567), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6568) );
  OR2X2 OR2X2_1893 ( .A(AES_CORE_DATAPATH__abc_16259_n6566), .B(AES_CORE_DATAPATH__abc_16259_n6568), .Y(AES_CORE_DATAPATH__abc_16259_n6569) );
  OR2X2 OR2X2_1894 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf5), .B(AES_CORE_DATAPATH_bkp_2__10_), .Y(AES_CORE_DATAPATH__abc_16259_n6570) );
  OR2X2 OR2X2_1895 ( .A(AES_CORE_DATAPATH__abc_16259_n6572), .B(AES_CORE_DATAPATH__abc_16259_n6573), .Y(AES_CORE_DATAPATH__abc_16259_n6574) );
  OR2X2 OR2X2_1896 ( .A(AES_CORE_DATAPATH__abc_16259_n6574), .B(AES_CORE_DATAPATH__abc_16259_n6063_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6575) );
  OR2X2 OR2X2_1897 ( .A(_auto_iopadmap_cc_313_execute_26916_10_), .B(AES_CORE_DATAPATH__abc_16259_n6074_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6576) );
  OR2X2 OR2X2_1898 ( .A(AES_CORE_DATAPATH__abc_16259_n6565), .B(AES_CORE_DATAPATH__abc_16259_n6577), .Y(AES_CORE_DATAPATH__abc_16259_n6578) );
  OR2X2 OR2X2_1899 ( .A(AES_CORE_DATAPATH__abc_16259_n3269), .B(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n6579) );
  OR2X2 OR2X2_19 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n132), .B(AES_CORE_CONTROL_UNIT__abc_15841_n130_1), .Y(AES_CORE_CONTROL_UNIT__abc_10818_n59) );
  OR2X2 OR2X2_190 ( .A(AES_CORE_DATAPATH__abc_16259_n2717_1), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n2718) );
  OR2X2 OR2X2_1900 ( .A(AES_CORE_DATAPATH__abc_16259_n6581), .B(AES_CORE_DATAPATH__abc_16259_n6582), .Y(AES_CORE_DATAPATH__abc_16259_n6583) );
  OR2X2 OR2X2_1901 ( .A(AES_CORE_DATAPATH__abc_16259_n6588), .B(AES_CORE_DATAPATH__abc_16259_n6586), .Y(AES_CORE_DATAPATH__abc_16259_n6589) );
  OR2X2 OR2X2_1902 ( .A(AES_CORE_DATAPATH__abc_16259_n6585), .B(AES_CORE_DATAPATH__abc_16259_n6589), .Y(AES_CORE_DATAPATH__abc_16259_n6590) );
  OR2X2 OR2X2_1903 ( .A(AES_CORE_DATAPATH__abc_16259_n6592), .B(AES_CORE_DATAPATH__abc_16259_n6091), .Y(AES_CORE_DATAPATH__abc_16259_n6593) );
  OR2X2 OR2X2_1904 ( .A(AES_CORE_DATAPATH__abc_16259_n6591), .B(AES_CORE_DATAPATH__abc_16259_n6593), .Y(AES_CORE_DATAPATH__abc_16259_n6594) );
  OR2X2 OR2X2_1905 ( .A(AES_CORE_DATAPATH__abc_16259_n6595), .B(AES_CORE_DATAPATH__abc_16259_n6563), .Y(AES_CORE_DATAPATH__abc_16259_n6596) );
  OR2X2 OR2X2_1906 ( .A(AES_CORE_DATAPATH__abc_16259_n6598), .B(AES_CORE_DATAPATH__abc_16259_n6556), .Y(AES_CORE_DATAPATH__abc_16259_n6599) );
  OR2X2 OR2X2_1907 ( .A(AES_CORE_DATAPATH__abc_16259_n6561), .B(AES_CORE_DATAPATH__abc_16259_n6600), .Y(AES_CORE_DATAPATH__abc_16259_n6601) );
  OR2X2 OR2X2_1908 ( .A(AES_CORE_DATAPATH__abc_16259_n6604), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6605) );
  OR2X2 OR2X2_1909 ( .A(AES_CORE_DATAPATH__abc_16259_n6603_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n6608), .Y(AES_CORE_DATAPATH__abc_16259_n6609) );
  OR2X2 OR2X2_191 ( .A(AES_CORE_DATAPATH__abc_16259_n2716), .B(AES_CORE_DATAPATH__abc_16259_n2718), .Y(AES_CORE_DATAPATH__abc_16259_n2719_1) );
  OR2X2 OR2X2_1910 ( .A(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf4), .B(AES_CORE_DATAPATH_col_0__10_), .Y(AES_CORE_DATAPATH__abc_16259_n6613) );
  OR2X2 OR2X2_1911 ( .A(AES_CORE_DATAPATH__abc_16259_n6617), .B(AES_CORE_DATAPATH__abc_16259_n6618), .Y(AES_CORE_DATAPATH__abc_16259_n6619) );
  OR2X2 OR2X2_1912 ( .A(AES_CORE_DATAPATH__abc_16259_n6620), .B(AES_CORE_DATAPATH__abc_16259_n6622), .Y(AES_CORE_DATAPATH__abc_16259_n6623) );
  OR2X2 OR2X2_1913 ( .A(AES_CORE_DATAPATH__abc_16259_n6625), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6626) );
  OR2X2 OR2X2_1914 ( .A(AES_CORE_DATAPATH__abc_16259_n6624), .B(AES_CORE_DATAPATH__abc_16259_n6626), .Y(AES_CORE_DATAPATH__abc_16259_n6627) );
  OR2X2 OR2X2_1915 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf4), .B(AES_CORE_DATAPATH_bkp_2__11_), .Y(AES_CORE_DATAPATH__abc_16259_n6628) );
  OR2X2 OR2X2_1916 ( .A(AES_CORE_DATAPATH__abc_16259_n6630), .B(AES_CORE_DATAPATH__abc_16259_n6631), .Y(AES_CORE_DATAPATH__abc_16259_n6632) );
  OR2X2 OR2X2_1917 ( .A(AES_CORE_DATAPATH__abc_16259_n6632), .B(AES_CORE_DATAPATH__abc_16259_n6063_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6633) );
  OR2X2 OR2X2_1918 ( .A(_auto_iopadmap_cc_313_execute_26916_11_), .B(AES_CORE_DATAPATH__abc_16259_n6074_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6634) );
  OR2X2 OR2X2_1919 ( .A(AES_CORE_DATAPATH__abc_16259_n6623), .B(AES_CORE_DATAPATH__abc_16259_n6635), .Y(AES_CORE_DATAPATH__abc_16259_n6636) );
  OR2X2 OR2X2_192 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf5), .B(AES_CORE_DATAPATH_iv_2__26_), .Y(AES_CORE_DATAPATH__abc_16259_n2720) );
  OR2X2 OR2X2_1920 ( .A(AES_CORE_DATAPATH__abc_16259_n3309), .B(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6637) );
  OR2X2 OR2X2_1921 ( .A(AES_CORE_DATAPATH__abc_16259_n6639), .B(AES_CORE_DATAPATH__abc_16259_n6640), .Y(AES_CORE_DATAPATH__abc_16259_n6641) );
  OR2X2 OR2X2_1922 ( .A(AES_CORE_DATAPATH__abc_16259_n6645), .B(AES_CORE_DATAPATH__abc_16259_n6586), .Y(AES_CORE_DATAPATH__abc_16259_n6646) );
  OR2X2 OR2X2_1923 ( .A(AES_CORE_DATAPATH__abc_16259_n6643), .B(AES_CORE_DATAPATH__abc_16259_n6646), .Y(AES_CORE_DATAPATH__abc_16259_n6647) );
  OR2X2 OR2X2_1924 ( .A(AES_CORE_DATAPATH__abc_16259_n6649), .B(AES_CORE_DATAPATH__abc_16259_n6091), .Y(AES_CORE_DATAPATH__abc_16259_n6650) );
  OR2X2 OR2X2_1925 ( .A(AES_CORE_DATAPATH__abc_16259_n6648), .B(AES_CORE_DATAPATH__abc_16259_n6650), .Y(AES_CORE_DATAPATH__abc_16259_n6651) );
  OR2X2 OR2X2_1926 ( .A(AES_CORE_DATAPATH__abc_16259_n6595), .B(AES_CORE_DATAPATH__abc_16259_n6621), .Y(AES_CORE_DATAPATH__abc_16259_n6652) );
  OR2X2 OR2X2_1927 ( .A(AES_CORE_DATAPATH__abc_16259_n6654), .B(AES_CORE_DATAPATH__abc_16259_n6556), .Y(AES_CORE_DATAPATH__abc_16259_n6655) );
  OR2X2 OR2X2_1928 ( .A(AES_CORE_DATAPATH__abc_16259_n6619), .B(AES_CORE_DATAPATH__abc_16259_n6600), .Y(AES_CORE_DATAPATH__abc_16259_n6656) );
  OR2X2 OR2X2_1929 ( .A(AES_CORE_DATAPATH__abc_16259_n6658), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6659) );
  OR2X2 OR2X2_193 ( .A(AES_CORE_DATAPATH__abc_16259_n2722), .B(AES_CORE_DATAPATH__abc_16259_n2723_1), .Y(_auto_iopadmap_cc_313_execute_26916_26_) );
  OR2X2 OR2X2_1930 ( .A(AES_CORE_DATAPATH__abc_16259_n6603_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n6662), .Y(AES_CORE_DATAPATH__abc_16259_n6663) );
  OR2X2 OR2X2_1931 ( .A(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf2), .B(AES_CORE_DATAPATH_col_0__11_), .Y(AES_CORE_DATAPATH__abc_16259_n6667) );
  OR2X2 OR2X2_1932 ( .A(AES_CORE_DATAPATH__abc_16259_n6670), .B(AES_CORE_DATAPATH__abc_16259_n6671), .Y(AES_CORE_DATAPATH__abc_16259_n6672) );
  OR2X2 OR2X2_1933 ( .A(AES_CORE_DATAPATH__abc_16259_n6674), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6675) );
  OR2X2 OR2X2_1934 ( .A(AES_CORE_DATAPATH__abc_16259_n6673), .B(AES_CORE_DATAPATH__abc_16259_n6675), .Y(AES_CORE_DATAPATH__abc_16259_n6676) );
  OR2X2 OR2X2_1935 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf3), .B(AES_CORE_DATAPATH_bkp_2__12_), .Y(AES_CORE_DATAPATH__abc_16259_n6677) );
  OR2X2 OR2X2_1936 ( .A(AES_CORE_DATAPATH__abc_16259_n6679), .B(AES_CORE_DATAPATH__abc_16259_n6680), .Y(AES_CORE_DATAPATH__abc_16259_n6681) );
  OR2X2 OR2X2_1937 ( .A(AES_CORE_DATAPATH__abc_16259_n6681), .B(AES_CORE_DATAPATH__abc_16259_n6063_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6682) );
  OR2X2 OR2X2_1938 ( .A(_auto_iopadmap_cc_313_execute_26916_12_), .B(AES_CORE_DATAPATH__abc_16259_n6074_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6683) );
  OR2X2 OR2X2_1939 ( .A(AES_CORE_DATAPATH__abc_16259_n6672), .B(AES_CORE_DATAPATH__abc_16259_n6684), .Y(AES_CORE_DATAPATH__abc_16259_n6685) );
  OR2X2 OR2X2_194 ( .A(AES_CORE_DATAPATH__abc_16259_n2726), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n2727_1) );
  OR2X2 OR2X2_1940 ( .A(AES_CORE_DATAPATH__abc_16259_n6688), .B(AES_CORE_DATAPATH__abc_16259_n6689), .Y(AES_CORE_DATAPATH__abc_16259_n6690) );
  OR2X2 OR2X2_1941 ( .A(AES_CORE_DATAPATH__abc_16259_n6690), .B(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6691) );
  OR2X2 OR2X2_1942 ( .A(AES_CORE_DATAPATH__abc_16259_n6693), .B(AES_CORE_DATAPATH__abc_16259_n6694), .Y(AES_CORE_DATAPATH__abc_16259_n6695) );
  OR2X2 OR2X2_1943 ( .A(AES_CORE_DATAPATH__abc_16259_n6696), .B(AES_CORE_DATAPATH__abc_16259_n6057_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6697) );
  OR2X2 OR2X2_1944 ( .A(_auto_iopadmap_cc_313_execute_26916_12_), .B(AES_CORE_CONTROL_UNIT_last_round_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6698) );
  OR2X2 OR2X2_1945 ( .A(AES_CORE_DATAPATH__abc_16259_n6696), .B(AES_CORE_DATAPATH__abc_16259_n6095_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6701) );
  OR2X2 OR2X2_1946 ( .A(AES_CORE_DATAPATH__abc_16259_n6097_bF_buf2), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_12_), .Y(AES_CORE_DATAPATH__abc_16259_n6702) );
  OR2X2 OR2X2_1947 ( .A(AES_CORE_DATAPATH__abc_16259_n6704), .B(AES_CORE_DATAPATH__abc_16259_n6705), .Y(AES_CORE_DATAPATH__abc_16259_n6706) );
  OR2X2 OR2X2_1948 ( .A(AES_CORE_DATAPATH__abc_16259_n6706), .B(AES_CORE_DATAPATH__abc_16259_n6700), .Y(AES_CORE_DATAPATH__abc_16259_n6707) );
  OR2X2 OR2X2_1949 ( .A(AES_CORE_DATAPATH__abc_16259_n6708), .B(AES_CORE_DATAPATH__abc_16259_n6709), .Y(AES_CORE_DATAPATH__abc_16259_n6710) );
  OR2X2 OR2X2_195 ( .A(AES_CORE_DATAPATH__abc_16259_n2725), .B(AES_CORE_DATAPATH__abc_16259_n2727_1), .Y(AES_CORE_DATAPATH__abc_16259_n2728) );
  OR2X2 OR2X2_1950 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf1), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_44_), .Y(AES_CORE_DATAPATH__abc_16259_n6711) );
  OR2X2 OR2X2_1951 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf0), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_44_), .Y(AES_CORE_DATAPATH__abc_16259_n6712) );
  OR2X2 OR2X2_1952 ( .A(AES_CORE_DATAPATH__abc_16259_n6710), .B(AES_CORE_DATAPATH__abc_16259_n6714), .Y(AES_CORE_DATAPATH__abc_16259_n6715) );
  OR2X2 OR2X2_1953 ( .A(AES_CORE_DATAPATH__abc_16259_n6716), .B(AES_CORE_DATAPATH__abc_16259_n6669), .Y(AES_CORE_DATAPATH__0col_0__31_0__12_) );
  OR2X2 OR2X2_1954 ( .A(AES_CORE_DATAPATH__abc_16259_n6720), .B(AES_CORE_DATAPATH__abc_16259_n6721), .Y(AES_CORE_DATAPATH__abc_16259_n6722) );
  OR2X2 OR2X2_1955 ( .A(AES_CORE_DATAPATH__abc_16259_n6723), .B(AES_CORE_DATAPATH__abc_16259_n6725), .Y(AES_CORE_DATAPATH__abc_16259_n6726) );
  OR2X2 OR2X2_1956 ( .A(AES_CORE_DATAPATH__abc_16259_n6728), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6729) );
  OR2X2 OR2X2_1957 ( .A(AES_CORE_DATAPATH__abc_16259_n6727), .B(AES_CORE_DATAPATH__abc_16259_n6729), .Y(AES_CORE_DATAPATH__abc_16259_n6730) );
  OR2X2 OR2X2_1958 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf2), .B(AES_CORE_DATAPATH_bkp_2__13_), .Y(AES_CORE_DATAPATH__abc_16259_n6731) );
  OR2X2 OR2X2_1959 ( .A(AES_CORE_DATAPATH__abc_16259_n6733), .B(AES_CORE_DATAPATH__abc_16259_n6734), .Y(AES_CORE_DATAPATH__abc_16259_n6735) );
  OR2X2 OR2X2_196 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf4), .B(AES_CORE_DATAPATH_iv_2__27_), .Y(AES_CORE_DATAPATH__abc_16259_n2729) );
  OR2X2 OR2X2_1960 ( .A(AES_CORE_DATAPATH__abc_16259_n6735), .B(AES_CORE_DATAPATH__abc_16259_n6063_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n6736) );
  OR2X2 OR2X2_1961 ( .A(_auto_iopadmap_cc_313_execute_26916_13_), .B(AES_CORE_DATAPATH__abc_16259_n6074_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6737) );
  OR2X2 OR2X2_1962 ( .A(AES_CORE_DATAPATH__abc_16259_n6726), .B(AES_CORE_DATAPATH__abc_16259_n6738), .Y(AES_CORE_DATAPATH__abc_16259_n6739) );
  OR2X2 OR2X2_1963 ( .A(AES_CORE_DATAPATH__abc_16259_n3389), .B(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n6740) );
  OR2X2 OR2X2_1964 ( .A(AES_CORE_DATAPATH__abc_16259_n6742), .B(AES_CORE_DATAPATH__abc_16259_n6743), .Y(AES_CORE_DATAPATH__abc_16259_n6744) );
  OR2X2 OR2X2_1965 ( .A(AES_CORE_DATAPATH__abc_16259_n6748), .B(AES_CORE_DATAPATH__abc_16259_n6586), .Y(AES_CORE_DATAPATH__abc_16259_n6749) );
  OR2X2 OR2X2_1966 ( .A(AES_CORE_DATAPATH__abc_16259_n6746), .B(AES_CORE_DATAPATH__abc_16259_n6749), .Y(AES_CORE_DATAPATH__abc_16259_n6750) );
  OR2X2 OR2X2_1967 ( .A(AES_CORE_DATAPATH__abc_16259_n6752), .B(AES_CORE_DATAPATH__abc_16259_n6091), .Y(AES_CORE_DATAPATH__abc_16259_n6753) );
  OR2X2 OR2X2_1968 ( .A(AES_CORE_DATAPATH__abc_16259_n6751), .B(AES_CORE_DATAPATH__abc_16259_n6753), .Y(AES_CORE_DATAPATH__abc_16259_n6754) );
  OR2X2 OR2X2_1969 ( .A(AES_CORE_DATAPATH__abc_16259_n6595), .B(AES_CORE_DATAPATH__abc_16259_n6724), .Y(AES_CORE_DATAPATH__abc_16259_n6755) );
  OR2X2 OR2X2_197 ( .A(AES_CORE_DATAPATH__abc_16259_n2731_1), .B(AES_CORE_DATAPATH__abc_16259_n2732), .Y(_auto_iopadmap_cc_313_execute_26916_27_) );
  OR2X2 OR2X2_1970 ( .A(AES_CORE_DATAPATH__abc_16259_n6757), .B(AES_CORE_DATAPATH__abc_16259_n6556), .Y(AES_CORE_DATAPATH__abc_16259_n6758) );
  OR2X2 OR2X2_1971 ( .A(AES_CORE_DATAPATH__abc_16259_n6722), .B(AES_CORE_DATAPATH__abc_16259_n6600), .Y(AES_CORE_DATAPATH__abc_16259_n6759) );
  OR2X2 OR2X2_1972 ( .A(AES_CORE_DATAPATH__abc_16259_n6761), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf14), .Y(AES_CORE_DATAPATH__abc_16259_n6762) );
  OR2X2 OR2X2_1973 ( .A(AES_CORE_DATAPATH__abc_16259_n6603_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n6765), .Y(AES_CORE_DATAPATH__abc_16259_n6766) );
  OR2X2 OR2X2_1974 ( .A(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf5), .B(AES_CORE_DATAPATH_col_0__13_), .Y(AES_CORE_DATAPATH__abc_16259_n6770) );
  OR2X2 OR2X2_1975 ( .A(AES_CORE_DATAPATH__abc_16259_n6773), .B(AES_CORE_DATAPATH__abc_16259_n6774), .Y(AES_CORE_DATAPATH__abc_16259_n6775) );
  OR2X2 OR2X2_1976 ( .A(AES_CORE_DATAPATH__abc_16259_n6777), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n6778) );
  OR2X2 OR2X2_1977 ( .A(AES_CORE_DATAPATH__abc_16259_n6776), .B(AES_CORE_DATAPATH__abc_16259_n6778), .Y(AES_CORE_DATAPATH__abc_16259_n6779) );
  OR2X2 OR2X2_1978 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf1), .B(AES_CORE_DATAPATH_bkp_2__14_), .Y(AES_CORE_DATAPATH__abc_16259_n6780) );
  OR2X2 OR2X2_1979 ( .A(AES_CORE_DATAPATH__abc_16259_n6782), .B(AES_CORE_DATAPATH__abc_16259_n6783), .Y(AES_CORE_DATAPATH__abc_16259_n6784) );
  OR2X2 OR2X2_198 ( .A(AES_CORE_DATAPATH__abc_16259_n2735_1), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n2736) );
  OR2X2 OR2X2_1980 ( .A(AES_CORE_DATAPATH__abc_16259_n6784), .B(AES_CORE_DATAPATH__abc_16259_n6063_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6785) );
  OR2X2 OR2X2_1981 ( .A(_auto_iopadmap_cc_313_execute_26916_14_), .B(AES_CORE_DATAPATH__abc_16259_n6074_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n6786) );
  OR2X2 OR2X2_1982 ( .A(AES_CORE_DATAPATH__abc_16259_n6775), .B(AES_CORE_DATAPATH__abc_16259_n6787), .Y(AES_CORE_DATAPATH__abc_16259_n6788) );
  OR2X2 OR2X2_1983 ( .A(AES_CORE_DATAPATH__abc_16259_n6791), .B(AES_CORE_DATAPATH__abc_16259_n6792), .Y(AES_CORE_DATAPATH__abc_16259_n6793) );
  OR2X2 OR2X2_1984 ( .A(AES_CORE_DATAPATH__abc_16259_n6793), .B(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n6794) );
  OR2X2 OR2X2_1985 ( .A(AES_CORE_DATAPATH__abc_16259_n6796), .B(AES_CORE_DATAPATH__abc_16259_n6797), .Y(AES_CORE_DATAPATH__abc_16259_n6798) );
  OR2X2 OR2X2_1986 ( .A(AES_CORE_DATAPATH__abc_16259_n6799), .B(AES_CORE_DATAPATH__abc_16259_n6057_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6800) );
  OR2X2 OR2X2_1987 ( .A(_auto_iopadmap_cc_313_execute_26916_14_), .B(AES_CORE_CONTROL_UNIT_last_round_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n6801) );
  OR2X2 OR2X2_1988 ( .A(AES_CORE_DATAPATH__abc_16259_n6799), .B(AES_CORE_DATAPATH__abc_16259_n6095_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6804) );
  OR2X2 OR2X2_1989 ( .A(AES_CORE_DATAPATH__abc_16259_n6097_bF_buf0), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_14_), .Y(AES_CORE_DATAPATH__abc_16259_n6805) );
  OR2X2 OR2X2_199 ( .A(AES_CORE_DATAPATH__abc_16259_n2734), .B(AES_CORE_DATAPATH__abc_16259_n2736), .Y(AES_CORE_DATAPATH__abc_16259_n2737_1) );
  OR2X2 OR2X2_1990 ( .A(AES_CORE_DATAPATH__abc_16259_n6807), .B(AES_CORE_DATAPATH__abc_16259_n6808), .Y(AES_CORE_DATAPATH__abc_16259_n6809) );
  OR2X2 OR2X2_1991 ( .A(AES_CORE_DATAPATH__abc_16259_n6809), .B(AES_CORE_DATAPATH__abc_16259_n6803), .Y(AES_CORE_DATAPATH__abc_16259_n6810) );
  OR2X2 OR2X2_1992 ( .A(AES_CORE_DATAPATH__abc_16259_n6811), .B(AES_CORE_DATAPATH__abc_16259_n6812), .Y(AES_CORE_DATAPATH__abc_16259_n6813) );
  OR2X2 OR2X2_1993 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf0), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_46_), .Y(AES_CORE_DATAPATH__abc_16259_n6814) );
  OR2X2 OR2X2_1994 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf12), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_46_), .Y(AES_CORE_DATAPATH__abc_16259_n6815) );
  OR2X2 OR2X2_1995 ( .A(AES_CORE_DATAPATH__abc_16259_n6813), .B(AES_CORE_DATAPATH__abc_16259_n6817), .Y(AES_CORE_DATAPATH__abc_16259_n6818) );
  OR2X2 OR2X2_1996 ( .A(AES_CORE_DATAPATH__abc_16259_n6819), .B(AES_CORE_DATAPATH__abc_16259_n6772), .Y(AES_CORE_DATAPATH__0col_0__31_0__14_) );
  OR2X2 OR2X2_1997 ( .A(AES_CORE_DATAPATH__abc_16259_n6823), .B(AES_CORE_DATAPATH__abc_16259_n6824), .Y(AES_CORE_DATAPATH__abc_16259_n6825) );
  OR2X2 OR2X2_1998 ( .A(AES_CORE_DATAPATH__abc_16259_n6826), .B(AES_CORE_DATAPATH__abc_16259_n6828), .Y(AES_CORE_DATAPATH__abc_16259_n6829) );
  OR2X2 OR2X2_1999 ( .A(AES_CORE_DATAPATH__abc_16259_n6831), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n6832) );
  OR2X2 OR2X2_2 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n75), .B(AES_CORE_CONTROL_UNIT_state_3_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n76_1) );
  OR2X2 OR2X2_20 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n134), .B(AES_CORE_CONTROL_UNIT__abc_15841_n135), .Y(AES_CORE_CONTROL_UNIT__abc_10818_n79) );
  OR2X2 OR2X2_200 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf3), .B(AES_CORE_DATAPATH_iv_2__28_), .Y(AES_CORE_DATAPATH__abc_16259_n2738) );
  OR2X2 OR2X2_2000 ( .A(AES_CORE_DATAPATH__abc_16259_n6830), .B(AES_CORE_DATAPATH__abc_16259_n6832), .Y(AES_CORE_DATAPATH__abc_16259_n6833) );
  OR2X2 OR2X2_2001 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf0), .B(AES_CORE_DATAPATH_bkp_2__15_), .Y(AES_CORE_DATAPATH__abc_16259_n6834) );
  OR2X2 OR2X2_2002 ( .A(AES_CORE_DATAPATH__abc_16259_n6836), .B(AES_CORE_DATAPATH__abc_16259_n6837), .Y(AES_CORE_DATAPATH__abc_16259_n6838) );
  OR2X2 OR2X2_2003 ( .A(AES_CORE_DATAPATH__abc_16259_n6838), .B(AES_CORE_DATAPATH__abc_16259_n6063_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6839) );
  OR2X2 OR2X2_2004 ( .A(_auto_iopadmap_cc_313_execute_26916_15_), .B(AES_CORE_DATAPATH__abc_16259_n6074_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6840) );
  OR2X2 OR2X2_2005 ( .A(AES_CORE_DATAPATH__abc_16259_n6829), .B(AES_CORE_DATAPATH__abc_16259_n6841), .Y(AES_CORE_DATAPATH__abc_16259_n6842) );
  OR2X2 OR2X2_2006 ( .A(AES_CORE_DATAPATH__abc_16259_n3469), .B(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6843) );
  OR2X2 OR2X2_2007 ( .A(AES_CORE_DATAPATH__abc_16259_n6845), .B(AES_CORE_DATAPATH__abc_16259_n6846), .Y(AES_CORE_DATAPATH__abc_16259_n6847) );
  OR2X2 OR2X2_2008 ( .A(AES_CORE_DATAPATH__abc_16259_n6851), .B(AES_CORE_DATAPATH__abc_16259_n6586), .Y(AES_CORE_DATAPATH__abc_16259_n6852) );
  OR2X2 OR2X2_2009 ( .A(AES_CORE_DATAPATH__abc_16259_n6849), .B(AES_CORE_DATAPATH__abc_16259_n6852), .Y(AES_CORE_DATAPATH__abc_16259_n6853) );
  OR2X2 OR2X2_201 ( .A(AES_CORE_DATAPATH__abc_16259_n2740), .B(AES_CORE_DATAPATH__abc_16259_n2741), .Y(_auto_iopadmap_cc_313_execute_26916_28_) );
  OR2X2 OR2X2_2010 ( .A(AES_CORE_DATAPATH__abc_16259_n6855), .B(AES_CORE_DATAPATH__abc_16259_n6091), .Y(AES_CORE_DATAPATH__abc_16259_n6856) );
  OR2X2 OR2X2_2011 ( .A(AES_CORE_DATAPATH__abc_16259_n6854), .B(AES_CORE_DATAPATH__abc_16259_n6856), .Y(AES_CORE_DATAPATH__abc_16259_n6857) );
  OR2X2 OR2X2_2012 ( .A(AES_CORE_DATAPATH__abc_16259_n6595), .B(AES_CORE_DATAPATH__abc_16259_n6827), .Y(AES_CORE_DATAPATH__abc_16259_n6858) );
  OR2X2 OR2X2_2013 ( .A(AES_CORE_DATAPATH__abc_16259_n6860), .B(AES_CORE_DATAPATH__abc_16259_n6556), .Y(AES_CORE_DATAPATH__abc_16259_n6861) );
  OR2X2 OR2X2_2014 ( .A(AES_CORE_DATAPATH__abc_16259_n6825), .B(AES_CORE_DATAPATH__abc_16259_n6600), .Y(AES_CORE_DATAPATH__abc_16259_n6862) );
  OR2X2 OR2X2_2015 ( .A(AES_CORE_DATAPATH__abc_16259_n6864), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf11), .Y(AES_CORE_DATAPATH__abc_16259_n6865) );
  OR2X2 OR2X2_2016 ( .A(AES_CORE_DATAPATH__abc_16259_n6603_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n6868), .Y(AES_CORE_DATAPATH__abc_16259_n6869) );
  OR2X2 OR2X2_2017 ( .A(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf2), .B(AES_CORE_DATAPATH_col_0__15_), .Y(AES_CORE_DATAPATH__abc_16259_n6873) );
  OR2X2 OR2X2_2018 ( .A(AES_CORE_DATAPATH__abc_16259_n6878), .B(AES_CORE_DATAPATH__abc_16259_n6879), .Y(AES_CORE_DATAPATH__abc_16259_n6880) );
  OR2X2 OR2X2_2019 ( .A(AES_CORE_DATAPATH__abc_16259_n6059_bF_buf5), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_16_), .Y(AES_CORE_DATAPATH__abc_16259_n6882) );
  OR2X2 OR2X2_202 ( .A(AES_CORE_DATAPATH__abc_16259_n2744), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n2745) );
  OR2X2 OR2X2_2020 ( .A(AES_CORE_DATAPATH__abc_16259_n6881), .B(AES_CORE_DATAPATH__abc_16259_n6883), .Y(AES_CORE_DATAPATH__abc_16259_n6884) );
  OR2X2 OR2X2_2021 ( .A(AES_CORE_DATAPATH__abc_16259_n6886), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n6887) );
  OR2X2 OR2X2_2022 ( .A(AES_CORE_DATAPATH__abc_16259_n6885), .B(AES_CORE_DATAPATH__abc_16259_n6887), .Y(AES_CORE_DATAPATH__abc_16259_n6888) );
  OR2X2 OR2X2_2023 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf7), .B(AES_CORE_DATAPATH_bkp_2__16_), .Y(AES_CORE_DATAPATH__abc_16259_n6889) );
  OR2X2 OR2X2_2024 ( .A(AES_CORE_DATAPATH__abc_16259_n6891), .B(AES_CORE_DATAPATH__abc_16259_n6892), .Y(AES_CORE_DATAPATH__abc_16259_n6893) );
  OR2X2 OR2X2_2025 ( .A(AES_CORE_DATAPATH__abc_16259_n6893), .B(AES_CORE_DATAPATH__abc_16259_n6063_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6894) );
  OR2X2 OR2X2_2026 ( .A(_auto_iopadmap_cc_313_execute_26916_16_), .B(AES_CORE_DATAPATH__abc_16259_n6074_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n6895) );
  OR2X2 OR2X2_2027 ( .A(AES_CORE_DATAPATH__abc_16259_n6884), .B(AES_CORE_DATAPATH__abc_16259_n6897), .Y(AES_CORE_DATAPATH__abc_16259_n6898) );
  OR2X2 OR2X2_2028 ( .A(AES_CORE_DATAPATH__abc_16259_n3509), .B(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6899) );
  OR2X2 OR2X2_2029 ( .A(AES_CORE_DATAPATH__abc_16259_n6900), .B(AES_CORE_DATAPATH__abc_16259_n6896), .Y(AES_CORE_DATAPATH__abc_16259_n6901) );
  OR2X2 OR2X2_203 ( .A(AES_CORE_DATAPATH__abc_16259_n2743), .B(AES_CORE_DATAPATH__abc_16259_n2745), .Y(AES_CORE_DATAPATH__abc_16259_n2746_1) );
  OR2X2 OR2X2_2030 ( .A(AES_CORE_DATAPATH__abc_16259_n6902), .B(AES_CORE_DATAPATH__abc_16259_n6057_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6903) );
  OR2X2 OR2X2_2031 ( .A(_auto_iopadmap_cc_313_execute_26916_16_), .B(AES_CORE_CONTROL_UNIT_last_round_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6904) );
  OR2X2 OR2X2_2032 ( .A(AES_CORE_DATAPATH__abc_16259_n6902), .B(AES_CORE_DATAPATH__abc_16259_n6095_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6907) );
  OR2X2 OR2X2_2033 ( .A(AES_CORE_DATAPATH__abc_16259_n6097_bF_buf3), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_16_), .Y(AES_CORE_DATAPATH__abc_16259_n6908) );
  OR2X2 OR2X2_2034 ( .A(AES_CORE_DATAPATH__abc_16259_n6910), .B(AES_CORE_DATAPATH__abc_16259_n6911), .Y(AES_CORE_DATAPATH__abc_16259_n6912) );
  OR2X2 OR2X2_2035 ( .A(AES_CORE_DATAPATH__abc_16259_n6912), .B(AES_CORE_DATAPATH__abc_16259_n6906), .Y(AES_CORE_DATAPATH__abc_16259_n6913) );
  OR2X2 OR2X2_2036 ( .A(AES_CORE_DATAPATH__abc_16259_n6914), .B(AES_CORE_DATAPATH__abc_16259_n6915), .Y(AES_CORE_DATAPATH__abc_16259_n6916) );
  OR2X2 OR2X2_2037 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf12), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_80_), .Y(AES_CORE_DATAPATH__abc_16259_n6917) );
  OR2X2 OR2X2_2038 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf9), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_16_), .Y(AES_CORE_DATAPATH__abc_16259_n6918) );
  OR2X2 OR2X2_2039 ( .A(AES_CORE_DATAPATH__abc_16259_n6916), .B(AES_CORE_DATAPATH__abc_16259_n6920), .Y(AES_CORE_DATAPATH__abc_16259_n6921) );
  OR2X2 OR2X2_204 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf2), .B(AES_CORE_DATAPATH_iv_2__29_), .Y(AES_CORE_DATAPATH__abc_16259_n2747) );
  OR2X2 OR2X2_2040 ( .A(AES_CORE_DATAPATH__abc_16259_n6922), .B(AES_CORE_DATAPATH__abc_16259_n6875), .Y(AES_CORE_DATAPATH__0col_0__31_0__16_) );
  OR2X2 OR2X2_2041 ( .A(AES_CORE_DATAPATH__abc_16259_n6926), .B(AES_CORE_DATAPATH__abc_16259_n6927), .Y(AES_CORE_DATAPATH__abc_16259_n6928) );
  OR2X2 OR2X2_2042 ( .A(AES_CORE_DATAPATH__abc_16259_n6929), .B(AES_CORE_DATAPATH__abc_16259_n6931), .Y(AES_CORE_DATAPATH__abc_16259_n6932) );
  OR2X2 OR2X2_2043 ( .A(AES_CORE_DATAPATH__abc_16259_n6934), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n6935) );
  OR2X2 OR2X2_2044 ( .A(AES_CORE_DATAPATH__abc_16259_n6933), .B(AES_CORE_DATAPATH__abc_16259_n6935), .Y(AES_CORE_DATAPATH__abc_16259_n6936) );
  OR2X2 OR2X2_2045 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf6), .B(AES_CORE_DATAPATH_bkp_2__17_), .Y(AES_CORE_DATAPATH__abc_16259_n6937) );
  OR2X2 OR2X2_2046 ( .A(AES_CORE_DATAPATH__abc_16259_n6939), .B(AES_CORE_DATAPATH__abc_16259_n6940), .Y(AES_CORE_DATAPATH__abc_16259_n6941) );
  OR2X2 OR2X2_2047 ( .A(AES_CORE_DATAPATH__abc_16259_n6941), .B(AES_CORE_DATAPATH__abc_16259_n6063_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6942) );
  OR2X2 OR2X2_2048 ( .A(_auto_iopadmap_cc_313_execute_26916_17_), .B(AES_CORE_DATAPATH__abc_16259_n6074_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n6943) );
  OR2X2 OR2X2_2049 ( .A(AES_CORE_DATAPATH__abc_16259_n6932), .B(AES_CORE_DATAPATH__abc_16259_n6944), .Y(AES_CORE_DATAPATH__abc_16259_n6945) );
  OR2X2 OR2X2_205 ( .A(AES_CORE_DATAPATH__abc_16259_n2749), .B(AES_CORE_DATAPATH__abc_16259_n2750), .Y(_auto_iopadmap_cc_313_execute_26916_29_) );
  OR2X2 OR2X2_2050 ( .A(AES_CORE_DATAPATH__abc_16259_n3549_1), .B(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n6946) );
  OR2X2 OR2X2_2051 ( .A(AES_CORE_DATAPATH__abc_16259_n6948), .B(AES_CORE_DATAPATH__abc_16259_n6949), .Y(AES_CORE_DATAPATH__abc_16259_n6950) );
  OR2X2 OR2X2_2052 ( .A(AES_CORE_DATAPATH__abc_16259_n6954), .B(AES_CORE_DATAPATH__abc_16259_n6586), .Y(AES_CORE_DATAPATH__abc_16259_n6955) );
  OR2X2 OR2X2_2053 ( .A(AES_CORE_DATAPATH__abc_16259_n6952), .B(AES_CORE_DATAPATH__abc_16259_n6955), .Y(AES_CORE_DATAPATH__abc_16259_n6956) );
  OR2X2 OR2X2_2054 ( .A(AES_CORE_DATAPATH__abc_16259_n6958), .B(AES_CORE_DATAPATH__abc_16259_n6091), .Y(AES_CORE_DATAPATH__abc_16259_n6959) );
  OR2X2 OR2X2_2055 ( .A(AES_CORE_DATAPATH__abc_16259_n6957), .B(AES_CORE_DATAPATH__abc_16259_n6959), .Y(AES_CORE_DATAPATH__abc_16259_n6960) );
  OR2X2 OR2X2_2056 ( .A(AES_CORE_DATAPATH__abc_16259_n6595), .B(AES_CORE_DATAPATH__abc_16259_n6930), .Y(AES_CORE_DATAPATH__abc_16259_n6961) );
  OR2X2 OR2X2_2057 ( .A(AES_CORE_DATAPATH__abc_16259_n6963), .B(AES_CORE_DATAPATH__abc_16259_n6556), .Y(AES_CORE_DATAPATH__abc_16259_n6964) );
  OR2X2 OR2X2_2058 ( .A(AES_CORE_DATAPATH__abc_16259_n6928), .B(AES_CORE_DATAPATH__abc_16259_n6600), .Y(AES_CORE_DATAPATH__abc_16259_n6965) );
  OR2X2 OR2X2_2059 ( .A(AES_CORE_DATAPATH__abc_16259_n6967), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf8), .Y(AES_CORE_DATAPATH__abc_16259_n6968) );
  OR2X2 OR2X2_206 ( .A(AES_CORE_DATAPATH__abc_16259_n2753_1), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n2754) );
  OR2X2 OR2X2_2060 ( .A(AES_CORE_DATAPATH__abc_16259_n6603_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n6971), .Y(AES_CORE_DATAPATH__abc_16259_n6972) );
  OR2X2 OR2X2_2061 ( .A(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf5), .B(AES_CORE_DATAPATH_col_0__17_), .Y(AES_CORE_DATAPATH__abc_16259_n6976) );
  OR2X2 OR2X2_2062 ( .A(AES_CORE_DATAPATH__abc_16259_n6979), .B(AES_CORE_DATAPATH__abc_16259_n6980), .Y(AES_CORE_DATAPATH__abc_16259_n6981) );
  OR2X2 OR2X2_2063 ( .A(AES_CORE_DATAPATH__abc_16259_n6983), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n6984) );
  OR2X2 OR2X2_2064 ( .A(AES_CORE_DATAPATH__abc_16259_n6982), .B(AES_CORE_DATAPATH__abc_16259_n6984), .Y(AES_CORE_DATAPATH__abc_16259_n6985) );
  OR2X2 OR2X2_2065 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf5), .B(AES_CORE_DATAPATH_bkp_2__18_), .Y(AES_CORE_DATAPATH__abc_16259_n6986) );
  OR2X2 OR2X2_2066 ( .A(AES_CORE_DATAPATH__abc_16259_n6988), .B(AES_CORE_DATAPATH__abc_16259_n6989), .Y(AES_CORE_DATAPATH__abc_16259_n6990) );
  OR2X2 OR2X2_2067 ( .A(AES_CORE_DATAPATH__abc_16259_n6990), .B(AES_CORE_DATAPATH__abc_16259_n6063_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n6991) );
  OR2X2 OR2X2_2068 ( .A(_auto_iopadmap_cc_313_execute_26916_18_), .B(AES_CORE_DATAPATH__abc_16259_n6074_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n6992) );
  OR2X2 OR2X2_2069 ( .A(AES_CORE_DATAPATH__abc_16259_n6981), .B(AES_CORE_DATAPATH__abc_16259_n6993), .Y(AES_CORE_DATAPATH__abc_16259_n6994) );
  OR2X2 OR2X2_207 ( .A(AES_CORE_DATAPATH__abc_16259_n2752_1), .B(AES_CORE_DATAPATH__abc_16259_n2754), .Y(AES_CORE_DATAPATH__abc_16259_n2755_1) );
  OR2X2 OR2X2_2070 ( .A(AES_CORE_DATAPATH__abc_16259_n6997), .B(AES_CORE_DATAPATH__abc_16259_n6998), .Y(AES_CORE_DATAPATH__abc_16259_n6999) );
  OR2X2 OR2X2_2071 ( .A(AES_CORE_DATAPATH__abc_16259_n6999), .B(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n7000) );
  OR2X2 OR2X2_2072 ( .A(AES_CORE_DATAPATH__abc_16259_n7002), .B(AES_CORE_DATAPATH__abc_16259_n7003), .Y(AES_CORE_DATAPATH__abc_16259_n7004) );
  OR2X2 OR2X2_2073 ( .A(AES_CORE_DATAPATH__abc_16259_n7005), .B(AES_CORE_DATAPATH__abc_16259_n6057_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n7006) );
  OR2X2 OR2X2_2074 ( .A(_auto_iopadmap_cc_313_execute_26916_18_), .B(AES_CORE_CONTROL_UNIT_last_round_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n7007) );
  OR2X2 OR2X2_2075 ( .A(AES_CORE_DATAPATH__abc_16259_n7005), .B(AES_CORE_DATAPATH__abc_16259_n6095_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n7010) );
  OR2X2 OR2X2_2076 ( .A(AES_CORE_DATAPATH__abc_16259_n6097_bF_buf1), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_18_), .Y(AES_CORE_DATAPATH__abc_16259_n7011) );
  OR2X2 OR2X2_2077 ( .A(AES_CORE_DATAPATH__abc_16259_n7013), .B(AES_CORE_DATAPATH__abc_16259_n7014), .Y(AES_CORE_DATAPATH__abc_16259_n7015) );
  OR2X2 OR2X2_2078 ( .A(AES_CORE_DATAPATH__abc_16259_n7015), .B(AES_CORE_DATAPATH__abc_16259_n7009), .Y(AES_CORE_DATAPATH__abc_16259_n7016) );
  OR2X2 OR2X2_2079 ( .A(AES_CORE_DATAPATH__abc_16259_n7017), .B(AES_CORE_DATAPATH__abc_16259_n7018), .Y(AES_CORE_DATAPATH__abc_16259_n7019) );
  OR2X2 OR2X2_208 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf1), .B(AES_CORE_DATAPATH_iv_2__30_), .Y(AES_CORE_DATAPATH__abc_16259_n2756_1) );
  OR2X2 OR2X2_2080 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf11), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_82_), .Y(AES_CORE_DATAPATH__abc_16259_n7020) );
  OR2X2 OR2X2_2081 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf6), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_18_), .Y(AES_CORE_DATAPATH__abc_16259_n7021) );
  OR2X2 OR2X2_2082 ( .A(AES_CORE_DATAPATH__abc_16259_n7019), .B(AES_CORE_DATAPATH__abc_16259_n7023), .Y(AES_CORE_DATAPATH__abc_16259_n7024) );
  OR2X2 OR2X2_2083 ( .A(AES_CORE_DATAPATH__abc_16259_n7025), .B(AES_CORE_DATAPATH__abc_16259_n6978), .Y(AES_CORE_DATAPATH__0col_0__31_0__18_) );
  OR2X2 OR2X2_2084 ( .A(AES_CORE_DATAPATH__abc_16259_n7028), .B(AES_CORE_DATAPATH__abc_16259_n7029), .Y(AES_CORE_DATAPATH__abc_16259_n7030) );
  OR2X2 OR2X2_2085 ( .A(AES_CORE_DATAPATH__abc_16259_n7032), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7033) );
  OR2X2 OR2X2_2086 ( .A(AES_CORE_DATAPATH__abc_16259_n7031), .B(AES_CORE_DATAPATH__abc_16259_n7033), .Y(AES_CORE_DATAPATH__abc_16259_n7034) );
  OR2X2 OR2X2_2087 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf4), .B(AES_CORE_DATAPATH_bkp_2__19_), .Y(AES_CORE_DATAPATH__abc_16259_n7035) );
  OR2X2 OR2X2_2088 ( .A(AES_CORE_DATAPATH__abc_16259_n7037), .B(AES_CORE_DATAPATH__abc_16259_n7038), .Y(AES_CORE_DATAPATH__abc_16259_n7039) );
  OR2X2 OR2X2_2089 ( .A(AES_CORE_DATAPATH__abc_16259_n7039), .B(AES_CORE_DATAPATH__abc_16259_n6063_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7040) );
  OR2X2 OR2X2_209 ( .A(AES_CORE_DATAPATH__abc_16259_n2758), .B(AES_CORE_DATAPATH__abc_16259_n2759), .Y(_auto_iopadmap_cc_313_execute_26916_30_) );
  OR2X2 OR2X2_2090 ( .A(_auto_iopadmap_cc_313_execute_26916_19_), .B(AES_CORE_DATAPATH__abc_16259_n6074_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n7041) );
  OR2X2 OR2X2_2091 ( .A(AES_CORE_DATAPATH__abc_16259_n7030), .B(AES_CORE_DATAPATH__abc_16259_n7042), .Y(AES_CORE_DATAPATH__abc_16259_n7043) );
  OR2X2 OR2X2_2092 ( .A(AES_CORE_DATAPATH__abc_16259_n7046), .B(AES_CORE_DATAPATH__abc_16259_n7047), .Y(AES_CORE_DATAPATH__abc_16259_n7048) );
  OR2X2 OR2X2_2093 ( .A(AES_CORE_DATAPATH__abc_16259_n7048), .B(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7049) );
  OR2X2 OR2X2_2094 ( .A(AES_CORE_DATAPATH__abc_16259_n7051), .B(AES_CORE_DATAPATH__abc_16259_n7052), .Y(AES_CORE_DATAPATH__abc_16259_n7053) );
  OR2X2 OR2X2_2095 ( .A(AES_CORE_DATAPATH__abc_16259_n7054), .B(AES_CORE_DATAPATH__abc_16259_n6057_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7055) );
  OR2X2 OR2X2_2096 ( .A(_auto_iopadmap_cc_313_execute_26916_19_), .B(AES_CORE_CONTROL_UNIT_last_round_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n7056) );
  OR2X2 OR2X2_2097 ( .A(AES_CORE_DATAPATH__abc_16259_n7054), .B(AES_CORE_DATAPATH__abc_16259_n6095_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7059) );
  OR2X2 OR2X2_2098 ( .A(AES_CORE_DATAPATH__abc_16259_n6097_bF_buf0), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_19_), .Y(AES_CORE_DATAPATH__abc_16259_n7060) );
  OR2X2 OR2X2_2099 ( .A(AES_CORE_DATAPATH__abc_16259_n7062), .B(AES_CORE_DATAPATH__abc_16259_n7063), .Y(AES_CORE_DATAPATH__abc_16259_n7064) );
  OR2X2 OR2X2_21 ( .A(AES_CORE_CONTROL_UNIT_state_12_), .B(AES_CORE_CONTROL_UNIT_state_4_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n137) );
  OR2X2 OR2X2_210 ( .A(AES_CORE_DATAPATH__abc_16259_n2762_1), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n2763) );
  OR2X2 OR2X2_2100 ( .A(AES_CORE_DATAPATH__abc_16259_n7064), .B(AES_CORE_DATAPATH__abc_16259_n7058), .Y(AES_CORE_DATAPATH__abc_16259_n7065) );
  OR2X2 OR2X2_2101 ( .A(AES_CORE_DATAPATH__abc_16259_n7066), .B(AES_CORE_DATAPATH__abc_16259_n7067), .Y(AES_CORE_DATAPATH__abc_16259_n7068) );
  OR2X2 OR2X2_2102 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf10), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_83_), .Y(AES_CORE_DATAPATH__abc_16259_n7069) );
  OR2X2 OR2X2_2103 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf5), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_19_), .Y(AES_CORE_DATAPATH__abc_16259_n7070) );
  OR2X2 OR2X2_2104 ( .A(AES_CORE_DATAPATH__abc_16259_n7068), .B(AES_CORE_DATAPATH__abc_16259_n7072), .Y(AES_CORE_DATAPATH__abc_16259_n7073) );
  OR2X2 OR2X2_2105 ( .A(AES_CORE_DATAPATH__abc_16259_n7074), .B(AES_CORE_DATAPATH__abc_16259_n7027), .Y(AES_CORE_DATAPATH__0col_0__31_0__19_) );
  OR2X2 OR2X2_2106 ( .A(AES_CORE_DATAPATH__abc_16259_n3669), .B(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n7077) );
  OR2X2 OR2X2_2107 ( .A(AES_CORE_DATAPATH__abc_16259_n6059_bF_buf1), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_20_), .Y(AES_CORE_DATAPATH__abc_16259_n7078) );
  OR2X2 OR2X2_2108 ( .A(AES_CORE_DATAPATH__abc_16259_n7081), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n7082) );
  OR2X2 OR2X2_2109 ( .A(AES_CORE_DATAPATH__abc_16259_n7080), .B(AES_CORE_DATAPATH__abc_16259_n7082), .Y(AES_CORE_DATAPATH__abc_16259_n7083) );
  OR2X2 OR2X2_211 ( .A(AES_CORE_DATAPATH__abc_16259_n2761), .B(AES_CORE_DATAPATH__abc_16259_n2763), .Y(AES_CORE_DATAPATH__abc_16259_n2764_1) );
  OR2X2 OR2X2_2110 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf3), .B(AES_CORE_DATAPATH_bkp_2__20_), .Y(AES_CORE_DATAPATH__abc_16259_n7084) );
  OR2X2 OR2X2_2111 ( .A(AES_CORE_DATAPATH__abc_16259_n7086), .B(AES_CORE_DATAPATH__abc_16259_n7087), .Y(AES_CORE_DATAPATH__abc_16259_n7088) );
  OR2X2 OR2X2_2112 ( .A(AES_CORE_DATAPATH__abc_16259_n7088), .B(AES_CORE_DATAPATH__abc_16259_n6063_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7089) );
  OR2X2 OR2X2_2113 ( .A(_auto_iopadmap_cc_313_execute_26916_20_), .B(AES_CORE_DATAPATH__abc_16259_n6074_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7090) );
  OR2X2 OR2X2_2114 ( .A(AES_CORE_DATAPATH__abc_16259_n7079), .B(AES_CORE_DATAPATH__abc_16259_n7091), .Y(AES_CORE_DATAPATH__abc_16259_n7092) );
  OR2X2 OR2X2_2115 ( .A(AES_CORE_DATAPATH__abc_16259_n7095), .B(AES_CORE_DATAPATH__abc_16259_n7096), .Y(AES_CORE_DATAPATH__abc_16259_n7097) );
  OR2X2 OR2X2_2116 ( .A(AES_CORE_DATAPATH__abc_16259_n7098), .B(AES_CORE_DATAPATH__abc_16259_n7099), .Y(AES_CORE_DATAPATH__abc_16259_n7100) );
  OR2X2 OR2X2_2117 ( .A(AES_CORE_DATAPATH__abc_16259_n7100), .B(AES_CORE_DATAPATH__abc_16259_n7101), .Y(AES_CORE_DATAPATH__abc_16259_n7102) );
  OR2X2 OR2X2_2118 ( .A(AES_CORE_DATAPATH__abc_16259_n7103), .B(AES_CORE_DATAPATH__abc_16259_n6057_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7104) );
  OR2X2 OR2X2_2119 ( .A(_auto_iopadmap_cc_313_execute_26916_20_), .B(AES_CORE_CONTROL_UNIT_last_round_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n7105) );
  OR2X2 OR2X2_212 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf0), .B(AES_CORE_DATAPATH_iv_2__31_), .Y(AES_CORE_DATAPATH__abc_16259_n2765) );
  OR2X2 OR2X2_2120 ( .A(AES_CORE_DATAPATH__abc_16259_n7103), .B(AES_CORE_DATAPATH__abc_16259_n6095_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7108) );
  OR2X2 OR2X2_2121 ( .A(AES_CORE_DATAPATH__abc_16259_n6097_bF_buf4), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_20_), .Y(AES_CORE_DATAPATH__abc_16259_n7109) );
  OR2X2 OR2X2_2122 ( .A(AES_CORE_DATAPATH__abc_16259_n7111), .B(AES_CORE_DATAPATH__abc_16259_n7112), .Y(AES_CORE_DATAPATH__abc_16259_n7113) );
  OR2X2 OR2X2_2123 ( .A(AES_CORE_DATAPATH__abc_16259_n7113), .B(AES_CORE_DATAPATH__abc_16259_n7107), .Y(AES_CORE_DATAPATH__abc_16259_n7114) );
  OR2X2 OR2X2_2124 ( .A(AES_CORE_DATAPATH__abc_16259_n7115), .B(AES_CORE_DATAPATH__abc_16259_n7116), .Y(AES_CORE_DATAPATH__abc_16259_n7117) );
  OR2X2 OR2X2_2125 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf9), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_84_), .Y(AES_CORE_DATAPATH__abc_16259_n7118) );
  OR2X2 OR2X2_2126 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf4), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_20_), .Y(AES_CORE_DATAPATH__abc_16259_n7119) );
  OR2X2 OR2X2_2127 ( .A(AES_CORE_DATAPATH__abc_16259_n7117), .B(AES_CORE_DATAPATH__abc_16259_n7121), .Y(AES_CORE_DATAPATH__abc_16259_n7122) );
  OR2X2 OR2X2_2128 ( .A(AES_CORE_DATAPATH__abc_16259_n7123), .B(AES_CORE_DATAPATH__abc_16259_n7076), .Y(AES_CORE_DATAPATH__0col_0__31_0__20_) );
  OR2X2 OR2X2_2129 ( .A(AES_CORE_DATAPATH__abc_16259_n7127), .B(AES_CORE_DATAPATH__abc_16259_n7128), .Y(AES_CORE_DATAPATH__abc_16259_n7129) );
  OR2X2 OR2X2_213 ( .A(AES_CORE_DATAPATH__abc_16259_n2767), .B(AES_CORE_DATAPATH__abc_16259_n2768), .Y(_auto_iopadmap_cc_313_execute_26916_31_) );
  OR2X2 OR2X2_2130 ( .A(AES_CORE_DATAPATH__abc_16259_n7130), .B(AES_CORE_DATAPATH__abc_16259_n7132), .Y(AES_CORE_DATAPATH__abc_16259_n7133) );
  OR2X2 OR2X2_2131 ( .A(AES_CORE_DATAPATH__abc_16259_n7135), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n7136) );
  OR2X2 OR2X2_2132 ( .A(AES_CORE_DATAPATH__abc_16259_n7134), .B(AES_CORE_DATAPATH__abc_16259_n7136), .Y(AES_CORE_DATAPATH__abc_16259_n7137) );
  OR2X2 OR2X2_2133 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf2), .B(AES_CORE_DATAPATH_bkp_2__21_), .Y(AES_CORE_DATAPATH__abc_16259_n7138) );
  OR2X2 OR2X2_2134 ( .A(AES_CORE_DATAPATH__abc_16259_n7140), .B(AES_CORE_DATAPATH__abc_16259_n7141), .Y(AES_CORE_DATAPATH__abc_16259_n7142) );
  OR2X2 OR2X2_2135 ( .A(AES_CORE_DATAPATH__abc_16259_n7142), .B(AES_CORE_DATAPATH__abc_16259_n6063_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n7143) );
  OR2X2 OR2X2_2136 ( .A(_auto_iopadmap_cc_313_execute_26916_21_), .B(AES_CORE_DATAPATH__abc_16259_n6074_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7144) );
  OR2X2 OR2X2_2137 ( .A(AES_CORE_DATAPATH__abc_16259_n7133), .B(AES_CORE_DATAPATH__abc_16259_n7145), .Y(AES_CORE_DATAPATH__abc_16259_n7146) );
  OR2X2 OR2X2_2138 ( .A(AES_CORE_DATAPATH__abc_16259_n3709), .B(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n7147) );
  OR2X2 OR2X2_2139 ( .A(AES_CORE_DATAPATH__abc_16259_n7149), .B(AES_CORE_DATAPATH__abc_16259_n7150), .Y(AES_CORE_DATAPATH__abc_16259_n7151) );
  OR2X2 OR2X2_214 ( .A(AES_CORE_DATAPATH_col_sel_host_0_), .B(AES_CORE_CONTROL_UNIT_sbox_sel_0_), .Y(AES_CORE_DATAPATH__abc_16259_n2771_1) );
  OR2X2 OR2X2_2140 ( .A(AES_CORE_DATAPATH__abc_16259_n7155), .B(AES_CORE_DATAPATH__abc_16259_n6586), .Y(AES_CORE_DATAPATH__abc_16259_n7156) );
  OR2X2 OR2X2_2141 ( .A(AES_CORE_DATAPATH__abc_16259_n7153), .B(AES_CORE_DATAPATH__abc_16259_n7156), .Y(AES_CORE_DATAPATH__abc_16259_n7157) );
  OR2X2 OR2X2_2142 ( .A(AES_CORE_DATAPATH__abc_16259_n7159), .B(AES_CORE_DATAPATH__abc_16259_n6091), .Y(AES_CORE_DATAPATH__abc_16259_n7160) );
  OR2X2 OR2X2_2143 ( .A(AES_CORE_DATAPATH__abc_16259_n7158), .B(AES_CORE_DATAPATH__abc_16259_n7160), .Y(AES_CORE_DATAPATH__abc_16259_n7161) );
  OR2X2 OR2X2_2144 ( .A(AES_CORE_DATAPATH__abc_16259_n6595), .B(AES_CORE_DATAPATH__abc_16259_n7131), .Y(AES_CORE_DATAPATH__abc_16259_n7162) );
  OR2X2 OR2X2_2145 ( .A(AES_CORE_DATAPATH__abc_16259_n7164), .B(AES_CORE_DATAPATH__abc_16259_n6556), .Y(AES_CORE_DATAPATH__abc_16259_n7165) );
  OR2X2 OR2X2_2146 ( .A(AES_CORE_DATAPATH__abc_16259_n7129), .B(AES_CORE_DATAPATH__abc_16259_n6600), .Y(AES_CORE_DATAPATH__abc_16259_n7166) );
  OR2X2 OR2X2_2147 ( .A(AES_CORE_DATAPATH__abc_16259_n7168), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7169) );
  OR2X2 OR2X2_2148 ( .A(AES_CORE_DATAPATH__abc_16259_n6603_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n7172), .Y(AES_CORE_DATAPATH__abc_16259_n7173) );
  OR2X2 OR2X2_2149 ( .A(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf0), .B(AES_CORE_DATAPATH_col_0__21_), .Y(AES_CORE_DATAPATH__abc_16259_n7177) );
  OR2X2 OR2X2_215 ( .A(AES_CORE_DATAPATH_col_sel_host_1_), .B(AES_CORE_CONTROL_UNIT_sbox_sel_1_), .Y(AES_CORE_DATAPATH__abc_16259_n2772_1) );
  OR2X2 OR2X2_2150 ( .A(AES_CORE_DATAPATH__abc_16259_n7180), .B(AES_CORE_DATAPATH__abc_16259_n7181), .Y(AES_CORE_DATAPATH__abc_16259_n7182) );
  OR2X2 OR2X2_2151 ( .A(AES_CORE_DATAPATH__abc_16259_n7184), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n7185) );
  OR2X2 OR2X2_2152 ( .A(AES_CORE_DATAPATH__abc_16259_n7183), .B(AES_CORE_DATAPATH__abc_16259_n7185), .Y(AES_CORE_DATAPATH__abc_16259_n7186) );
  OR2X2 OR2X2_2153 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf1), .B(AES_CORE_DATAPATH_bkp_2__22_), .Y(AES_CORE_DATAPATH__abc_16259_n7187) );
  OR2X2 OR2X2_2154 ( .A(AES_CORE_DATAPATH__abc_16259_n7189), .B(AES_CORE_DATAPATH__abc_16259_n7190), .Y(AES_CORE_DATAPATH__abc_16259_n7191) );
  OR2X2 OR2X2_2155 ( .A(AES_CORE_DATAPATH__abc_16259_n7191), .B(AES_CORE_DATAPATH__abc_16259_n6063_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n7192) );
  OR2X2 OR2X2_2156 ( .A(_auto_iopadmap_cc_313_execute_26916_22_), .B(AES_CORE_DATAPATH__abc_16259_n6074_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n7193) );
  OR2X2 OR2X2_2157 ( .A(AES_CORE_DATAPATH__abc_16259_n7182), .B(AES_CORE_DATAPATH__abc_16259_n7194), .Y(AES_CORE_DATAPATH__abc_16259_n7195) );
  OR2X2 OR2X2_2158 ( .A(AES_CORE_DATAPATH__abc_16259_n7198), .B(AES_CORE_DATAPATH__abc_16259_n7199), .Y(AES_CORE_DATAPATH__abc_16259_n7200) );
  OR2X2 OR2X2_2159 ( .A(AES_CORE_DATAPATH__abc_16259_n7200), .B(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n7201) );
  OR2X2 OR2X2_216 ( .A(AES_CORE_DATAPATH__abc_16259_n2771_1), .B(AES_CORE_DATAPATH__abc_16259_n2772_1), .Y(AES_CORE_DATAPATH__abc_16259_n2773) );
  OR2X2 OR2X2_2160 ( .A(AES_CORE_DATAPATH__abc_16259_n7203), .B(AES_CORE_DATAPATH__abc_16259_n7204), .Y(AES_CORE_DATAPATH__abc_16259_n7205) );
  OR2X2 OR2X2_2161 ( .A(AES_CORE_DATAPATH__abc_16259_n7206), .B(AES_CORE_DATAPATH__abc_16259_n6057_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n7207) );
  OR2X2 OR2X2_2162 ( .A(_auto_iopadmap_cc_313_execute_26916_22_), .B(AES_CORE_CONTROL_UNIT_last_round_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7208) );
  OR2X2 OR2X2_2163 ( .A(AES_CORE_DATAPATH__abc_16259_n7206), .B(AES_CORE_DATAPATH__abc_16259_n6095_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n7211) );
  OR2X2 OR2X2_2164 ( .A(AES_CORE_DATAPATH__abc_16259_n6097_bF_buf2), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_22_), .Y(AES_CORE_DATAPATH__abc_16259_n7212) );
  OR2X2 OR2X2_2165 ( .A(AES_CORE_DATAPATH__abc_16259_n7214), .B(AES_CORE_DATAPATH__abc_16259_n7215), .Y(AES_CORE_DATAPATH__abc_16259_n7216) );
  OR2X2 OR2X2_2166 ( .A(AES_CORE_DATAPATH__abc_16259_n7216), .B(AES_CORE_DATAPATH__abc_16259_n7210), .Y(AES_CORE_DATAPATH__abc_16259_n7217) );
  OR2X2 OR2X2_2167 ( .A(AES_CORE_DATAPATH__abc_16259_n7218), .B(AES_CORE_DATAPATH__abc_16259_n7219), .Y(AES_CORE_DATAPATH__abc_16259_n7220) );
  OR2X2 OR2X2_2168 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf8), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_86_), .Y(AES_CORE_DATAPATH__abc_16259_n7221) );
  OR2X2 OR2X2_2169 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf1), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_22_), .Y(AES_CORE_DATAPATH__abc_16259_n7222) );
  OR2X2 OR2X2_217 ( .A(AES_CORE_DATAPATH__abc_16259_n2773), .B(AES_CORE_CONTROL_UNIT_sbox_sel_2_), .Y(AES_CORE_DATAPATH__abc_16259_n2774) );
  OR2X2 OR2X2_2170 ( .A(AES_CORE_DATAPATH__abc_16259_n7220), .B(AES_CORE_DATAPATH__abc_16259_n7224), .Y(AES_CORE_DATAPATH__abc_16259_n7225) );
  OR2X2 OR2X2_2171 ( .A(AES_CORE_DATAPATH__abc_16259_n7226), .B(AES_CORE_DATAPATH__abc_16259_n7179), .Y(AES_CORE_DATAPATH__0col_0__31_0__22_) );
  OR2X2 OR2X2_2172 ( .A(AES_CORE_DATAPATH__abc_16259_n7231), .B(AES_CORE_DATAPATH__abc_16259_n7232), .Y(AES_CORE_DATAPATH__abc_16259_n7233) );
  OR2X2 OR2X2_2173 ( .A(AES_CORE_DATAPATH__abc_16259_n6059_bF_buf2), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_23_), .Y(AES_CORE_DATAPATH__abc_16259_n7235) );
  OR2X2 OR2X2_2174 ( .A(AES_CORE_DATAPATH__abc_16259_n7234), .B(AES_CORE_DATAPATH__abc_16259_n7236), .Y(AES_CORE_DATAPATH__abc_16259_n7237) );
  OR2X2 OR2X2_2175 ( .A(AES_CORE_DATAPATH__abc_16259_n7239), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n7240) );
  OR2X2 OR2X2_2176 ( .A(AES_CORE_DATAPATH__abc_16259_n7238), .B(AES_CORE_DATAPATH__abc_16259_n7240), .Y(AES_CORE_DATAPATH__abc_16259_n7241) );
  OR2X2 OR2X2_2177 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf0), .B(AES_CORE_DATAPATH_bkp_2__23_), .Y(AES_CORE_DATAPATH__abc_16259_n7242) );
  OR2X2 OR2X2_2178 ( .A(AES_CORE_DATAPATH__abc_16259_n7244), .B(AES_CORE_DATAPATH__abc_16259_n7245), .Y(AES_CORE_DATAPATH__abc_16259_n7246) );
  OR2X2 OR2X2_2179 ( .A(AES_CORE_DATAPATH__abc_16259_n7246), .B(AES_CORE_DATAPATH__abc_16259_n6063_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n7247) );
  OR2X2 OR2X2_218 ( .A(AES_CORE_DATAPATH__abc_16259_n2774_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n2770), .Y(AES_CORE_DATAPATH__abc_16259_n2775_1) );
  OR2X2 OR2X2_2180 ( .A(_auto_iopadmap_cc_313_execute_26916_23_), .B(AES_CORE_DATAPATH__abc_16259_n6074_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n7248) );
  OR2X2 OR2X2_2181 ( .A(AES_CORE_DATAPATH__abc_16259_n7237), .B(AES_CORE_DATAPATH__abc_16259_n7250), .Y(AES_CORE_DATAPATH__abc_16259_n7251) );
  OR2X2 OR2X2_2182 ( .A(AES_CORE_DATAPATH__abc_16259_n3789), .B(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7252) );
  OR2X2 OR2X2_2183 ( .A(AES_CORE_DATAPATH__abc_16259_n7253), .B(AES_CORE_DATAPATH__abc_16259_n7249), .Y(AES_CORE_DATAPATH__abc_16259_n7254) );
  OR2X2 OR2X2_2184 ( .A(AES_CORE_DATAPATH__abc_16259_n7255), .B(AES_CORE_DATAPATH__abc_16259_n6057_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n7256) );
  OR2X2 OR2X2_2185 ( .A(_auto_iopadmap_cc_313_execute_26916_23_), .B(AES_CORE_CONTROL_UNIT_last_round_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7257) );
  OR2X2 OR2X2_2186 ( .A(AES_CORE_DATAPATH__abc_16259_n7255), .B(AES_CORE_DATAPATH__abc_16259_n6095_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n7260) );
  OR2X2 OR2X2_2187 ( .A(AES_CORE_DATAPATH__abc_16259_n6097_bF_buf1), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_23_), .Y(AES_CORE_DATAPATH__abc_16259_n7261) );
  OR2X2 OR2X2_2188 ( .A(AES_CORE_DATAPATH__abc_16259_n7263), .B(AES_CORE_DATAPATH__abc_16259_n7264), .Y(AES_CORE_DATAPATH__abc_16259_n7265) );
  OR2X2 OR2X2_2189 ( .A(AES_CORE_DATAPATH__abc_16259_n7265), .B(AES_CORE_DATAPATH__abc_16259_n7259), .Y(AES_CORE_DATAPATH__abc_16259_n7266) );
  OR2X2 OR2X2_219 ( .A(AES_CORE_DATAPATH__abc_16259_n2773), .B(AES_CORE_DATAPATH__abc_16259_n2777_1), .Y(AES_CORE_DATAPATH__abc_16259_n2778) );
  OR2X2 OR2X2_2190 ( .A(AES_CORE_DATAPATH__abc_16259_n7267), .B(AES_CORE_DATAPATH__abc_16259_n7268), .Y(AES_CORE_DATAPATH__abc_16259_n7269) );
  OR2X2 OR2X2_2191 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf7), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_87_), .Y(AES_CORE_DATAPATH__abc_16259_n7270) );
  OR2X2 OR2X2_2192 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf0), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_23_), .Y(AES_CORE_DATAPATH__abc_16259_n7271) );
  OR2X2 OR2X2_2193 ( .A(AES_CORE_DATAPATH__abc_16259_n7269), .B(AES_CORE_DATAPATH__abc_16259_n7273), .Y(AES_CORE_DATAPATH__abc_16259_n7274) );
  OR2X2 OR2X2_2194 ( .A(AES_CORE_DATAPATH__abc_16259_n7275), .B(AES_CORE_DATAPATH__abc_16259_n7228), .Y(AES_CORE_DATAPATH__0col_0__31_0__23_) );
  OR2X2 OR2X2_2195 ( .A(AES_CORE_DATAPATH__abc_16259_n7278), .B(AES_CORE_DATAPATH__abc_16259_n7279), .Y(AES_CORE_DATAPATH__abc_16259_n7280) );
  OR2X2 OR2X2_2196 ( .A(AES_CORE_DATAPATH__abc_16259_n7282), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n7283) );
  OR2X2 OR2X2_2197 ( .A(AES_CORE_DATAPATH__abc_16259_n7281), .B(AES_CORE_DATAPATH__abc_16259_n7283), .Y(AES_CORE_DATAPATH__abc_16259_n7284) );
  OR2X2 OR2X2_2198 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf7), .B(AES_CORE_DATAPATH_bkp_2__24_), .Y(AES_CORE_DATAPATH__abc_16259_n7285) );
  OR2X2 OR2X2_2199 ( .A(AES_CORE_DATAPATH__abc_16259_n7287), .B(AES_CORE_DATAPATH__abc_16259_n7288), .Y(AES_CORE_DATAPATH__abc_16259_n7289) );
  OR2X2 OR2X2_22 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n137), .B(AES_CORE_CONTROL_UNIT_state_2_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n138) );
  OR2X2 OR2X2_220 ( .A(AES_CORE_DATAPATH__abc_16259_n2778_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n2776), .Y(AES_CORE_DATAPATH__abc_16259_n2779_1) );
  OR2X2 OR2X2_2200 ( .A(AES_CORE_DATAPATH__abc_16259_n7289), .B(AES_CORE_DATAPATH__abc_16259_n6063_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7290) );
  OR2X2 OR2X2_2201 ( .A(_auto_iopadmap_cc_313_execute_26916_24_), .B(AES_CORE_DATAPATH__abc_16259_n6074_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n7291) );
  OR2X2 OR2X2_2202 ( .A(AES_CORE_DATAPATH__abc_16259_n7280), .B(AES_CORE_DATAPATH__abc_16259_n7292), .Y(AES_CORE_DATAPATH__abc_16259_n7293) );
  OR2X2 OR2X2_2203 ( .A(AES_CORE_DATAPATH__abc_16259_n7296), .B(AES_CORE_DATAPATH__abc_16259_n7297), .Y(AES_CORE_DATAPATH__abc_16259_n7298) );
  OR2X2 OR2X2_2204 ( .A(AES_CORE_DATAPATH__abc_16259_n7298), .B(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n7299) );
  OR2X2 OR2X2_2205 ( .A(AES_CORE_DATAPATH__abc_16259_n7301), .B(AES_CORE_DATAPATH__abc_16259_n7302), .Y(AES_CORE_DATAPATH__abc_16259_n7303) );
  OR2X2 OR2X2_2206 ( .A(AES_CORE_DATAPATH__abc_16259_n7304), .B(AES_CORE_DATAPATH__abc_16259_n6057_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7305) );
  OR2X2 OR2X2_2207 ( .A(_auto_iopadmap_cc_313_execute_26916_24_), .B(AES_CORE_CONTROL_UNIT_last_round_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n7306) );
  OR2X2 OR2X2_2208 ( .A(AES_CORE_DATAPATH__abc_16259_n7304), .B(AES_CORE_DATAPATH__abc_16259_n6095_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7309) );
  OR2X2 OR2X2_2209 ( .A(AES_CORE_DATAPATH__abc_16259_n6097_bF_buf0), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_24_), .Y(AES_CORE_DATAPATH__abc_16259_n7310) );
  OR2X2 OR2X2_221 ( .A(AES_CORE_DATAPATH__abc_16259_n2787), .B(AES_CORE_DATAPATH__abc_16259_n2790), .Y(AES_CORE_DATAPATH__abc_16259_n2791) );
  OR2X2 OR2X2_2210 ( .A(AES_CORE_DATAPATH__abc_16259_n7312), .B(AES_CORE_DATAPATH__abc_16259_n7313), .Y(AES_CORE_DATAPATH__abc_16259_n7314) );
  OR2X2 OR2X2_2211 ( .A(AES_CORE_DATAPATH__abc_16259_n7314), .B(AES_CORE_DATAPATH__abc_16259_n7308), .Y(AES_CORE_DATAPATH__abc_16259_n7315) );
  OR2X2 OR2X2_2212 ( .A(AES_CORE_DATAPATH__abc_16259_n7316), .B(AES_CORE_DATAPATH__abc_16259_n7317), .Y(AES_CORE_DATAPATH__abc_16259_n7318) );
  OR2X2 OR2X2_2213 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf6), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_120_), .Y(AES_CORE_DATAPATH__abc_16259_n7319) );
  OR2X2 OR2X2_2214 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf14), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_120_), .Y(AES_CORE_DATAPATH__abc_16259_n7320) );
  OR2X2 OR2X2_2215 ( .A(AES_CORE_DATAPATH__abc_16259_n7318), .B(AES_CORE_DATAPATH__abc_16259_n7322), .Y(AES_CORE_DATAPATH__abc_16259_n7323) );
  OR2X2 OR2X2_2216 ( .A(AES_CORE_DATAPATH__abc_16259_n7324), .B(AES_CORE_DATAPATH__abc_16259_n7277), .Y(AES_CORE_DATAPATH__0col_0__31_0__24_) );
  OR2X2 OR2X2_2217 ( .A(AES_CORE_DATAPATH__abc_16259_n7327), .B(AES_CORE_DATAPATH__abc_16259_n7328), .Y(AES_CORE_DATAPATH__abc_16259_n7329) );
  OR2X2 OR2X2_2218 ( .A(AES_CORE_DATAPATH__abc_16259_n7331), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n7332) );
  OR2X2 OR2X2_2219 ( .A(AES_CORE_DATAPATH__abc_16259_n7330), .B(AES_CORE_DATAPATH__abc_16259_n7332), .Y(AES_CORE_DATAPATH__abc_16259_n7333) );
  OR2X2 OR2X2_222 ( .A(AES_CORE_DATAPATH__abc_16259_n2791), .B(AES_CORE_DATAPATH__abc_16259_n2783), .Y(AES_CORE_DATAPATH__abc_16259_n2792) );
  OR2X2 OR2X2_2220 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf6), .B(AES_CORE_DATAPATH_bkp_2__25_), .Y(AES_CORE_DATAPATH__abc_16259_n7334) );
  OR2X2 OR2X2_2221 ( .A(AES_CORE_DATAPATH__abc_16259_n7336), .B(AES_CORE_DATAPATH__abc_16259_n7337), .Y(AES_CORE_DATAPATH__abc_16259_n7338) );
  OR2X2 OR2X2_2222 ( .A(AES_CORE_DATAPATH__abc_16259_n7338), .B(AES_CORE_DATAPATH__abc_16259_n6063_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7339) );
  OR2X2 OR2X2_2223 ( .A(_auto_iopadmap_cc_313_execute_26916_25_), .B(AES_CORE_DATAPATH__abc_16259_n6074_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7340) );
  OR2X2 OR2X2_2224 ( .A(AES_CORE_DATAPATH__abc_16259_n7329), .B(AES_CORE_DATAPATH__abc_16259_n7341), .Y(AES_CORE_DATAPATH__abc_16259_n7342) );
  OR2X2 OR2X2_2225 ( .A(AES_CORE_DATAPATH__abc_16259_n7345), .B(AES_CORE_DATAPATH__abc_16259_n7346), .Y(AES_CORE_DATAPATH__abc_16259_n7347) );
  OR2X2 OR2X2_2226 ( .A(AES_CORE_DATAPATH__abc_16259_n7347), .B(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n7348) );
  OR2X2 OR2X2_2227 ( .A(AES_CORE_DATAPATH__abc_16259_n7350), .B(AES_CORE_DATAPATH__abc_16259_n7351), .Y(AES_CORE_DATAPATH__abc_16259_n7352) );
  OR2X2 OR2X2_2228 ( .A(AES_CORE_DATAPATH__abc_16259_n7353), .B(AES_CORE_DATAPATH__abc_16259_n6057_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7354) );
  OR2X2 OR2X2_2229 ( .A(_auto_iopadmap_cc_313_execute_26916_25_), .B(AES_CORE_CONTROL_UNIT_last_round_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n7355) );
  OR2X2 OR2X2_223 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk_bF_buf1), .B(AES_CORE_DATAPATH_rk_out_sel_pp2), .Y(AES_CORE_DATAPATH__abc_16259_n2796) );
  OR2X2 OR2X2_2230 ( .A(AES_CORE_DATAPATH__abc_16259_n7353), .B(AES_CORE_DATAPATH__abc_16259_n6095_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7358) );
  OR2X2 OR2X2_2231 ( .A(AES_CORE_DATAPATH__abc_16259_n6097_bF_buf4), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_25_), .Y(AES_CORE_DATAPATH__abc_16259_n7359) );
  OR2X2 OR2X2_2232 ( .A(AES_CORE_DATAPATH__abc_16259_n7361), .B(AES_CORE_DATAPATH__abc_16259_n7362), .Y(AES_CORE_DATAPATH__abc_16259_n7363) );
  OR2X2 OR2X2_2233 ( .A(AES_CORE_DATAPATH__abc_16259_n7363), .B(AES_CORE_DATAPATH__abc_16259_n7357), .Y(AES_CORE_DATAPATH__abc_16259_n7364) );
  OR2X2 OR2X2_2234 ( .A(AES_CORE_DATAPATH__abc_16259_n7365), .B(AES_CORE_DATAPATH__abc_16259_n7366), .Y(AES_CORE_DATAPATH__abc_16259_n7367) );
  OR2X2 OR2X2_2235 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf5), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_121_), .Y(AES_CORE_DATAPATH__abc_16259_n7368) );
  OR2X2 OR2X2_2236 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf13), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_121_), .Y(AES_CORE_DATAPATH__abc_16259_n7369) );
  OR2X2 OR2X2_2237 ( .A(AES_CORE_DATAPATH__abc_16259_n7367), .B(AES_CORE_DATAPATH__abc_16259_n7371), .Y(AES_CORE_DATAPATH__abc_16259_n7372) );
  OR2X2 OR2X2_2238 ( .A(AES_CORE_DATAPATH__abc_16259_n7373), .B(AES_CORE_DATAPATH__abc_16259_n7326), .Y(AES_CORE_DATAPATH__0col_0__31_0__25_) );
  OR2X2 OR2X2_2239 ( .A(AES_CORE_DATAPATH__abc_16259_n7378), .B(AES_CORE_DATAPATH__abc_16259_n7379), .Y(AES_CORE_DATAPATH__abc_16259_n7380) );
  OR2X2 OR2X2_224 ( .A(AES_CORE_DATAPATH__abc_16259_n2799), .B(AES_CORE_DATAPATH__abc_16259_n2797), .Y(AES_CORE_DATAPATH__abc_16259_n2800_1) );
  OR2X2 OR2X2_2240 ( .A(AES_CORE_DATAPATH__abc_16259_n6059_bF_buf4), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_26_), .Y(AES_CORE_DATAPATH__abc_16259_n7382) );
  OR2X2 OR2X2_2241 ( .A(AES_CORE_DATAPATH__abc_16259_n7381), .B(AES_CORE_DATAPATH__abc_16259_n7383), .Y(AES_CORE_DATAPATH__abc_16259_n7384) );
  OR2X2 OR2X2_2242 ( .A(AES_CORE_DATAPATH__abc_16259_n7386), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7387) );
  OR2X2 OR2X2_2243 ( .A(AES_CORE_DATAPATH__abc_16259_n7385), .B(AES_CORE_DATAPATH__abc_16259_n7387), .Y(AES_CORE_DATAPATH__abc_16259_n7388) );
  OR2X2 OR2X2_2244 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf5), .B(AES_CORE_DATAPATH_bkp_2__26_), .Y(AES_CORE_DATAPATH__abc_16259_n7389) );
  OR2X2 OR2X2_2245 ( .A(AES_CORE_DATAPATH__abc_16259_n7391), .B(AES_CORE_DATAPATH__abc_16259_n7392), .Y(AES_CORE_DATAPATH__abc_16259_n7393) );
  OR2X2 OR2X2_2246 ( .A(AES_CORE_DATAPATH__abc_16259_n7393), .B(AES_CORE_DATAPATH__abc_16259_n6063_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n7394) );
  OR2X2 OR2X2_2247 ( .A(_auto_iopadmap_cc_313_execute_26916_26_), .B(AES_CORE_DATAPATH__abc_16259_n6074_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7395) );
  OR2X2 OR2X2_2248 ( .A(AES_CORE_DATAPATH__abc_16259_n7384), .B(AES_CORE_DATAPATH__abc_16259_n7397), .Y(AES_CORE_DATAPATH__abc_16259_n7398) );
  OR2X2 OR2X2_2249 ( .A(AES_CORE_DATAPATH__abc_16259_n3909), .B(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n7399) );
  OR2X2 OR2X2_225 ( .A(AES_CORE_DATAPATH__abc_16259_n2800_1), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n2801_1) );
  OR2X2 OR2X2_2250 ( .A(AES_CORE_DATAPATH__abc_16259_n7400), .B(AES_CORE_DATAPATH__abc_16259_n7396), .Y(AES_CORE_DATAPATH__abc_16259_n7401) );
  OR2X2 OR2X2_2251 ( .A(AES_CORE_DATAPATH__abc_16259_n7402), .B(AES_CORE_DATAPATH__abc_16259_n6057_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n7403) );
  OR2X2 OR2X2_2252 ( .A(_auto_iopadmap_cc_313_execute_26916_26_), .B(AES_CORE_CONTROL_UNIT_last_round_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n7404) );
  OR2X2 OR2X2_2253 ( .A(AES_CORE_DATAPATH__abc_16259_n7402), .B(AES_CORE_DATAPATH__abc_16259_n6095_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n7407) );
  OR2X2 OR2X2_2254 ( .A(AES_CORE_DATAPATH__abc_16259_n6097_bF_buf3), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_26_), .Y(AES_CORE_DATAPATH__abc_16259_n7408) );
  OR2X2 OR2X2_2255 ( .A(AES_CORE_DATAPATH__abc_16259_n7410), .B(AES_CORE_DATAPATH__abc_16259_n7411), .Y(AES_CORE_DATAPATH__abc_16259_n7412) );
  OR2X2 OR2X2_2256 ( .A(AES_CORE_DATAPATH__abc_16259_n7412), .B(AES_CORE_DATAPATH__abc_16259_n7406), .Y(AES_CORE_DATAPATH__abc_16259_n7413) );
  OR2X2 OR2X2_2257 ( .A(AES_CORE_DATAPATH__abc_16259_n7414), .B(AES_CORE_DATAPATH__abc_16259_n7415), .Y(AES_CORE_DATAPATH__abc_16259_n7416) );
  OR2X2 OR2X2_2258 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf4), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_122_), .Y(AES_CORE_DATAPATH__abc_16259_n7417) );
  OR2X2 OR2X2_2259 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf12), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_122_), .Y(AES_CORE_DATAPATH__abc_16259_n7418) );
  OR2X2 OR2X2_226 ( .A(AES_CORE_DATAPATH__abc_16259_n2804_1_bF_buf4), .B(AES_CORE_DATAPATH_key_out_sel_pp2_1_), .Y(AES_CORE_DATAPATH__abc_16259_n2805) );
  OR2X2 OR2X2_2260 ( .A(AES_CORE_DATAPATH__abc_16259_n7416), .B(AES_CORE_DATAPATH__abc_16259_n7420), .Y(AES_CORE_DATAPATH__abc_16259_n7421) );
  OR2X2 OR2X2_2261 ( .A(AES_CORE_DATAPATH__abc_16259_n7422), .B(AES_CORE_DATAPATH__abc_16259_n7375), .Y(AES_CORE_DATAPATH__0col_0__31_0__26_) );
  OR2X2 OR2X2_2262 ( .A(AES_CORE_DATAPATH__abc_16259_n7425), .B(AES_CORE_DATAPATH__abc_16259_n7426), .Y(AES_CORE_DATAPATH__abc_16259_n7427) );
  OR2X2 OR2X2_2263 ( .A(AES_CORE_DATAPATH__abc_16259_n7429), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7430) );
  OR2X2 OR2X2_2264 ( .A(AES_CORE_DATAPATH__abc_16259_n7428), .B(AES_CORE_DATAPATH__abc_16259_n7430), .Y(AES_CORE_DATAPATH__abc_16259_n7431) );
  OR2X2 OR2X2_2265 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf4), .B(AES_CORE_DATAPATH_bkp_2__27_), .Y(AES_CORE_DATAPATH__abc_16259_n7432) );
  OR2X2 OR2X2_2266 ( .A(AES_CORE_DATAPATH__abc_16259_n7434), .B(AES_CORE_DATAPATH__abc_16259_n7435), .Y(AES_CORE_DATAPATH__abc_16259_n7436) );
  OR2X2 OR2X2_2267 ( .A(AES_CORE_DATAPATH__abc_16259_n7436), .B(AES_CORE_DATAPATH__abc_16259_n6063_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n7437) );
  OR2X2 OR2X2_2268 ( .A(_auto_iopadmap_cc_313_execute_26916_27_), .B(AES_CORE_DATAPATH__abc_16259_n6074_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n7438) );
  OR2X2 OR2X2_2269 ( .A(AES_CORE_DATAPATH__abc_16259_n7427), .B(AES_CORE_DATAPATH__abc_16259_n7439), .Y(AES_CORE_DATAPATH__abc_16259_n7440) );
  OR2X2 OR2X2_227 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf5), .B(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n2807) );
  OR2X2 OR2X2_2270 ( .A(AES_CORE_DATAPATH__abc_16259_n7443), .B(AES_CORE_DATAPATH__abc_16259_n7444), .Y(AES_CORE_DATAPATH__abc_16259_n7445) );
  OR2X2 OR2X2_2271 ( .A(AES_CORE_DATAPATH__abc_16259_n7445), .B(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7446) );
  OR2X2 OR2X2_2272 ( .A(AES_CORE_DATAPATH__abc_16259_n7448), .B(AES_CORE_DATAPATH__abc_16259_n7449), .Y(AES_CORE_DATAPATH__abc_16259_n7450) );
  OR2X2 OR2X2_2273 ( .A(AES_CORE_DATAPATH__abc_16259_n7451), .B(AES_CORE_DATAPATH__abc_16259_n6057_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n7452) );
  OR2X2 OR2X2_2274 ( .A(_auto_iopadmap_cc_313_execute_26916_27_), .B(AES_CORE_CONTROL_UNIT_last_round_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n7453) );
  OR2X2 OR2X2_2275 ( .A(AES_CORE_DATAPATH__abc_16259_n7451), .B(AES_CORE_DATAPATH__abc_16259_n6095_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n7456) );
  OR2X2 OR2X2_2276 ( .A(AES_CORE_DATAPATH__abc_16259_n6097_bF_buf2), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_27_), .Y(AES_CORE_DATAPATH__abc_16259_n7457) );
  OR2X2 OR2X2_2277 ( .A(AES_CORE_DATAPATH__abc_16259_n7459), .B(AES_CORE_DATAPATH__abc_16259_n7460), .Y(AES_CORE_DATAPATH__abc_16259_n7461) );
  OR2X2 OR2X2_2278 ( .A(AES_CORE_DATAPATH__abc_16259_n7461), .B(AES_CORE_DATAPATH__abc_16259_n7455), .Y(AES_CORE_DATAPATH__abc_16259_n7462) );
  OR2X2 OR2X2_2279 ( .A(AES_CORE_DATAPATH__abc_16259_n7463), .B(AES_CORE_DATAPATH__abc_16259_n7464), .Y(AES_CORE_DATAPATH__abc_16259_n7465) );
  OR2X2 OR2X2_228 ( .A(AES_CORE_DATAPATH__abc_16259_n2807_bF_buf5), .B(AES_CORE_DATAPATH_key_out_sel_pp1_1_), .Y(AES_CORE_DATAPATH__abc_16259_n2808_1) );
  OR2X2 OR2X2_2280 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf3), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_123_), .Y(AES_CORE_DATAPATH__abc_16259_n7466) );
  OR2X2 OR2X2_2281 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf11), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_123_), .Y(AES_CORE_DATAPATH__abc_16259_n7467) );
  OR2X2 OR2X2_2282 ( .A(AES_CORE_DATAPATH__abc_16259_n7465), .B(AES_CORE_DATAPATH__abc_16259_n7469), .Y(AES_CORE_DATAPATH__abc_16259_n7470) );
  OR2X2 OR2X2_2283 ( .A(AES_CORE_DATAPATH__abc_16259_n7471), .B(AES_CORE_DATAPATH__abc_16259_n7424), .Y(AES_CORE_DATAPATH__0col_0__31_0__27_) );
  OR2X2 OR2X2_2284 ( .A(AES_CORE_DATAPATH__abc_16259_n7476), .B(AES_CORE_DATAPATH__abc_16259_n7477), .Y(AES_CORE_DATAPATH__abc_16259_n7478) );
  OR2X2 OR2X2_2285 ( .A(AES_CORE_DATAPATH__abc_16259_n6059_bF_buf1), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_28_), .Y(AES_CORE_DATAPATH__abc_16259_n7480) );
  OR2X2 OR2X2_2286 ( .A(AES_CORE_DATAPATH__abc_16259_n7479), .B(AES_CORE_DATAPATH__abc_16259_n7481), .Y(AES_CORE_DATAPATH__abc_16259_n7482) );
  OR2X2 OR2X2_2287 ( .A(AES_CORE_DATAPATH__abc_16259_n7484), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n7485) );
  OR2X2 OR2X2_2288 ( .A(AES_CORE_DATAPATH__abc_16259_n7483), .B(AES_CORE_DATAPATH__abc_16259_n7485), .Y(AES_CORE_DATAPATH__abc_16259_n7486) );
  OR2X2 OR2X2_2289 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf3), .B(AES_CORE_DATAPATH_bkp_2__28_), .Y(AES_CORE_DATAPATH__abc_16259_n7487) );
  OR2X2 OR2X2_229 ( .A(AES_CORE_DATAPATH__abc_16259_n2812), .B(\key_sel_rd[1] ), .Y(AES_CORE_DATAPATH__abc_16259_n2813) );
  OR2X2 OR2X2_2290 ( .A(AES_CORE_DATAPATH__abc_16259_n7489), .B(AES_CORE_DATAPATH__abc_16259_n7490), .Y(AES_CORE_DATAPATH__abc_16259_n7491) );
  OR2X2 OR2X2_2291 ( .A(AES_CORE_DATAPATH__abc_16259_n7491), .B(AES_CORE_DATAPATH__abc_16259_n6063_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n7492) );
  OR2X2 OR2X2_2292 ( .A(_auto_iopadmap_cc_313_execute_26916_28_), .B(AES_CORE_DATAPATH__abc_16259_n6074_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n7493) );
  OR2X2 OR2X2_2293 ( .A(AES_CORE_DATAPATH__abc_16259_n7482), .B(AES_CORE_DATAPATH__abc_16259_n7495), .Y(AES_CORE_DATAPATH__abc_16259_n7496) );
  OR2X2 OR2X2_2294 ( .A(AES_CORE_DATAPATH__abc_16259_n3989), .B(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7497) );
  OR2X2 OR2X2_2295 ( .A(AES_CORE_DATAPATH__abc_16259_n7498), .B(AES_CORE_DATAPATH__abc_16259_n7494), .Y(AES_CORE_DATAPATH__abc_16259_n7499) );
  OR2X2 OR2X2_2296 ( .A(AES_CORE_DATAPATH__abc_16259_n7500), .B(AES_CORE_DATAPATH__abc_16259_n6057_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n7501) );
  OR2X2 OR2X2_2297 ( .A(_auto_iopadmap_cc_313_execute_26916_28_), .B(AES_CORE_CONTROL_UNIT_last_round_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7502) );
  OR2X2 OR2X2_2298 ( .A(AES_CORE_DATAPATH__abc_16259_n7500), .B(AES_CORE_DATAPATH__abc_16259_n6095_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n7505) );
  OR2X2 OR2X2_2299 ( .A(AES_CORE_DATAPATH__abc_16259_n6097_bF_buf1), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_28_), .Y(AES_CORE_DATAPATH__abc_16259_n7506) );
  OR2X2 OR2X2_23 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n138), .B(AES_CORE_CONTROL_UNIT_state_8_), .Y(AES_CORE_CONTROL_UNIT_bypass_rk) );
  OR2X2 OR2X2_230 ( .A(AES_CORE_DATAPATH__abc_16259_n2807_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n2816), .Y(AES_CORE_DATAPATH__abc_16259_n2817) );
  OR2X2 OR2X2_2300 ( .A(AES_CORE_DATAPATH__abc_16259_n7508), .B(AES_CORE_DATAPATH__abc_16259_n7509), .Y(AES_CORE_DATAPATH__abc_16259_n7510) );
  OR2X2 OR2X2_2301 ( .A(AES_CORE_DATAPATH__abc_16259_n7510), .B(AES_CORE_DATAPATH__abc_16259_n7504), .Y(AES_CORE_DATAPATH__abc_16259_n7511) );
  OR2X2 OR2X2_2302 ( .A(AES_CORE_DATAPATH__abc_16259_n7512), .B(AES_CORE_DATAPATH__abc_16259_n7513), .Y(AES_CORE_DATAPATH__abc_16259_n7514) );
  OR2X2 OR2X2_2303 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf2), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_124_), .Y(AES_CORE_DATAPATH__abc_16259_n7515) );
  OR2X2 OR2X2_2304 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf10), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_124_), .Y(AES_CORE_DATAPATH__abc_16259_n7516) );
  OR2X2 OR2X2_2305 ( .A(AES_CORE_DATAPATH__abc_16259_n7514), .B(AES_CORE_DATAPATH__abc_16259_n7518), .Y(AES_CORE_DATAPATH__abc_16259_n7519) );
  OR2X2 OR2X2_2306 ( .A(AES_CORE_DATAPATH__abc_16259_n7520), .B(AES_CORE_DATAPATH__abc_16259_n7473), .Y(AES_CORE_DATAPATH__0col_0__31_0__28_) );
  OR2X2 OR2X2_2307 ( .A(AES_CORE_DATAPATH__abc_16259_n7523), .B(AES_CORE_DATAPATH__abc_16259_n7524), .Y(AES_CORE_DATAPATH__abc_16259_n7525) );
  OR2X2 OR2X2_2308 ( .A(AES_CORE_DATAPATH__abc_16259_n7527), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n7528) );
  OR2X2 OR2X2_2309 ( .A(AES_CORE_DATAPATH__abc_16259_n7526), .B(AES_CORE_DATAPATH__abc_16259_n7528), .Y(AES_CORE_DATAPATH__abc_16259_n7529) );
  OR2X2 OR2X2_231 ( .A(AES_CORE_DATAPATH__abc_16259_n2804_1_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n2818), .Y(AES_CORE_DATAPATH__abc_16259_n2819) );
  OR2X2 OR2X2_2310 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf2), .B(AES_CORE_DATAPATH_bkp_2__29_), .Y(AES_CORE_DATAPATH__abc_16259_n7530) );
  OR2X2 OR2X2_2311 ( .A(AES_CORE_DATAPATH__abc_16259_n7532), .B(AES_CORE_DATAPATH__abc_16259_n7533), .Y(AES_CORE_DATAPATH__abc_16259_n7534) );
  OR2X2 OR2X2_2312 ( .A(AES_CORE_DATAPATH__abc_16259_n7534), .B(AES_CORE_DATAPATH__abc_16259_n6063_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7535) );
  OR2X2 OR2X2_2313 ( .A(_auto_iopadmap_cc_313_execute_26916_29_), .B(AES_CORE_DATAPATH__abc_16259_n6074_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n7536) );
  OR2X2 OR2X2_2314 ( .A(AES_CORE_DATAPATH__abc_16259_n7525), .B(AES_CORE_DATAPATH__abc_16259_n7537), .Y(AES_CORE_DATAPATH__abc_16259_n7538) );
  OR2X2 OR2X2_2315 ( .A(AES_CORE_DATAPATH__abc_16259_n7541), .B(AES_CORE_DATAPATH__abc_16259_n7542), .Y(AES_CORE_DATAPATH__abc_16259_n7543) );
  OR2X2 OR2X2_2316 ( .A(AES_CORE_DATAPATH__abc_16259_n7543), .B(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n7544) );
  OR2X2 OR2X2_2317 ( .A(AES_CORE_DATAPATH__abc_16259_n7546), .B(AES_CORE_DATAPATH__abc_16259_n7547), .Y(AES_CORE_DATAPATH__abc_16259_n7548) );
  OR2X2 OR2X2_2318 ( .A(AES_CORE_DATAPATH__abc_16259_n7549), .B(AES_CORE_DATAPATH__abc_16259_n6057_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7550) );
  OR2X2 OR2X2_2319 ( .A(_auto_iopadmap_cc_313_execute_26916_29_), .B(AES_CORE_CONTROL_UNIT_last_round_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7551) );
  OR2X2 OR2X2_232 ( .A(AES_CORE_DATAPATH__abc_16259_n2820), .B(AES_CORE_CONTROL_UNIT_bypass_key_en), .Y(AES_CORE_DATAPATH__abc_16259_n2821) );
  OR2X2 OR2X2_2320 ( .A(AES_CORE_DATAPATH__abc_16259_n7549), .B(AES_CORE_DATAPATH__abc_16259_n6095_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7554) );
  OR2X2 OR2X2_2321 ( .A(AES_CORE_DATAPATH__abc_16259_n6097_bF_buf0), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_29_), .Y(AES_CORE_DATAPATH__abc_16259_n7555) );
  OR2X2 OR2X2_2322 ( .A(AES_CORE_DATAPATH__abc_16259_n7557), .B(AES_CORE_DATAPATH__abc_16259_n7558), .Y(AES_CORE_DATAPATH__abc_16259_n7559) );
  OR2X2 OR2X2_2323 ( .A(AES_CORE_DATAPATH__abc_16259_n7559), .B(AES_CORE_DATAPATH__abc_16259_n7553), .Y(AES_CORE_DATAPATH__abc_16259_n7560) );
  OR2X2 OR2X2_2324 ( .A(AES_CORE_DATAPATH__abc_16259_n7561), .B(AES_CORE_DATAPATH__abc_16259_n7562), .Y(AES_CORE_DATAPATH__abc_16259_n7563) );
  OR2X2 OR2X2_2325 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf1), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_125_), .Y(AES_CORE_DATAPATH__abc_16259_n7564) );
  OR2X2 OR2X2_2326 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf9), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_125_), .Y(AES_CORE_DATAPATH__abc_16259_n7565) );
  OR2X2 OR2X2_2327 ( .A(AES_CORE_DATAPATH__abc_16259_n7563), .B(AES_CORE_DATAPATH__abc_16259_n7567), .Y(AES_CORE_DATAPATH__abc_16259_n7568) );
  OR2X2 OR2X2_2328 ( .A(AES_CORE_DATAPATH__abc_16259_n7569), .B(AES_CORE_DATAPATH__abc_16259_n7522), .Y(AES_CORE_DATAPATH__0col_0__31_0__29_) );
  OR2X2 OR2X2_2329 ( .A(AES_CORE_DATAPATH__abc_16259_n7572), .B(AES_CORE_DATAPATH__abc_16259_n7573), .Y(AES_CORE_DATAPATH__abc_16259_n7574) );
  OR2X2 OR2X2_233 ( .A(AES_CORE_DATAPATH__abc_16259_n2822_1), .B(\key_sel_rd[0] ), .Y(AES_CORE_DATAPATH__abc_16259_n2823) );
  OR2X2 OR2X2_2330 ( .A(AES_CORE_DATAPATH__abc_16259_n7576), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n7577) );
  OR2X2 OR2X2_2331 ( .A(AES_CORE_DATAPATH__abc_16259_n7575), .B(AES_CORE_DATAPATH__abc_16259_n7577), .Y(AES_CORE_DATAPATH__abc_16259_n7578) );
  OR2X2 OR2X2_2332 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf1), .B(AES_CORE_DATAPATH_bkp_2__30_), .Y(AES_CORE_DATAPATH__abc_16259_n7579) );
  OR2X2 OR2X2_2333 ( .A(AES_CORE_DATAPATH__abc_16259_n7581), .B(AES_CORE_DATAPATH__abc_16259_n7582), .Y(AES_CORE_DATAPATH__abc_16259_n7583) );
  OR2X2 OR2X2_2334 ( .A(AES_CORE_DATAPATH__abc_16259_n7583), .B(AES_CORE_DATAPATH__abc_16259_n6063_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7584) );
  OR2X2 OR2X2_2335 ( .A(_auto_iopadmap_cc_313_execute_26916_30_), .B(AES_CORE_DATAPATH__abc_16259_n6074_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7585) );
  OR2X2 OR2X2_2336 ( .A(AES_CORE_DATAPATH__abc_16259_n7574), .B(AES_CORE_DATAPATH__abc_16259_n7586), .Y(AES_CORE_DATAPATH__abc_16259_n7587) );
  OR2X2 OR2X2_2337 ( .A(AES_CORE_DATAPATH__abc_16259_n7590), .B(AES_CORE_DATAPATH__abc_16259_n7591), .Y(AES_CORE_DATAPATH__abc_16259_n7592) );
  OR2X2 OR2X2_2338 ( .A(AES_CORE_DATAPATH__abc_16259_n7592), .B(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n7593) );
  OR2X2 OR2X2_2339 ( .A(AES_CORE_DATAPATH__abc_16259_n7595), .B(AES_CORE_DATAPATH__abc_16259_n7596), .Y(AES_CORE_DATAPATH__abc_16259_n7597) );
  OR2X2 OR2X2_234 ( .A(AES_CORE_DATAPATH__abc_16259_n2826_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n2827), .Y(AES_CORE_DATAPATH__abc_16259_n2828) );
  OR2X2 OR2X2_2340 ( .A(AES_CORE_DATAPATH__abc_16259_n7598), .B(AES_CORE_DATAPATH__abc_16259_n6057_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7599) );
  OR2X2 OR2X2_2341 ( .A(_auto_iopadmap_cc_313_execute_26916_30_), .B(AES_CORE_CONTROL_UNIT_last_round_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n7600) );
  OR2X2 OR2X2_2342 ( .A(AES_CORE_DATAPATH__abc_16259_n7598), .B(AES_CORE_DATAPATH__abc_16259_n6095_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7603) );
  OR2X2 OR2X2_2343 ( .A(AES_CORE_DATAPATH__abc_16259_n6097_bF_buf4), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_30_), .Y(AES_CORE_DATAPATH__abc_16259_n7604) );
  OR2X2 OR2X2_2344 ( .A(AES_CORE_DATAPATH__abc_16259_n7606), .B(AES_CORE_DATAPATH__abc_16259_n7607), .Y(AES_CORE_DATAPATH__abc_16259_n7608) );
  OR2X2 OR2X2_2345 ( .A(AES_CORE_DATAPATH__abc_16259_n7608), .B(AES_CORE_DATAPATH__abc_16259_n7602), .Y(AES_CORE_DATAPATH__abc_16259_n7609) );
  OR2X2 OR2X2_2346 ( .A(AES_CORE_DATAPATH__abc_16259_n7610), .B(AES_CORE_DATAPATH__abc_16259_n7611), .Y(AES_CORE_DATAPATH__abc_16259_n7612) );
  OR2X2 OR2X2_2347 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf0), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_126_), .Y(AES_CORE_DATAPATH__abc_16259_n7613) );
  OR2X2 OR2X2_2348 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf8), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_126_), .Y(AES_CORE_DATAPATH__abc_16259_n7614) );
  OR2X2 OR2X2_2349 ( .A(AES_CORE_DATAPATH__abc_16259_n7612), .B(AES_CORE_DATAPATH__abc_16259_n7616), .Y(AES_CORE_DATAPATH__abc_16259_n7617) );
  OR2X2 OR2X2_235 ( .A(AES_CORE_DATAPATH__abc_16259_n2810_1), .B(AES_CORE_DATAPATH__abc_16259_n2813), .Y(AES_CORE_DATAPATH__abc_16259_n2829_1) );
  OR2X2 OR2X2_2350 ( .A(AES_CORE_DATAPATH__abc_16259_n7618), .B(AES_CORE_DATAPATH__abc_16259_n7571), .Y(AES_CORE_DATAPATH__0col_0__31_0__30_) );
  OR2X2 OR2X2_2351 ( .A(AES_CORE_DATAPATH__abc_16259_n7621), .B(AES_CORE_DATAPATH__abc_16259_n7622), .Y(AES_CORE_DATAPATH__abc_16259_n7623) );
  OR2X2 OR2X2_2352 ( .A(AES_CORE_DATAPATH__abc_16259_n7625), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n7626) );
  OR2X2 OR2X2_2353 ( .A(AES_CORE_DATAPATH__abc_16259_n7624), .B(AES_CORE_DATAPATH__abc_16259_n7626), .Y(AES_CORE_DATAPATH__abc_16259_n7627) );
  OR2X2 OR2X2_2354 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf0), .B(AES_CORE_DATAPATH_bkp_2__31_), .Y(AES_CORE_DATAPATH__abc_16259_n7628) );
  OR2X2 OR2X2_2355 ( .A(AES_CORE_DATAPATH__abc_16259_n7630), .B(AES_CORE_DATAPATH__abc_16259_n7631), .Y(AES_CORE_DATAPATH__abc_16259_n7632) );
  OR2X2 OR2X2_2356 ( .A(AES_CORE_DATAPATH__abc_16259_n7632), .B(AES_CORE_DATAPATH__abc_16259_n6063_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n7633) );
  OR2X2 OR2X2_2357 ( .A(_auto_iopadmap_cc_313_execute_26916_31_), .B(AES_CORE_DATAPATH__abc_16259_n6074_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7634) );
  OR2X2 OR2X2_2358 ( .A(AES_CORE_DATAPATH__abc_16259_n7623), .B(AES_CORE_DATAPATH__abc_16259_n7635), .Y(AES_CORE_DATAPATH__abc_16259_n7636) );
  OR2X2 OR2X2_2359 ( .A(AES_CORE_DATAPATH__abc_16259_n7639), .B(AES_CORE_DATAPATH__abc_16259_n7640), .Y(AES_CORE_DATAPATH__abc_16259_n7641) );
  OR2X2 OR2X2_236 ( .A(AES_CORE_DATAPATH__abc_16259_n2832), .B(AES_CORE_DATAPATH__abc_16259_n2833_1), .Y(AES_CORE_DATAPATH__abc_16259_n2834) );
  OR2X2 OR2X2_2360 ( .A(AES_CORE_DATAPATH__abc_16259_n7641), .B(AES_CORE_DATAPATH__abc_16259_n6058_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n7642) );
  OR2X2 OR2X2_2361 ( .A(AES_CORE_DATAPATH__abc_16259_n7644), .B(AES_CORE_DATAPATH__abc_16259_n7645), .Y(AES_CORE_DATAPATH__abc_16259_n7646) );
  OR2X2 OR2X2_2362 ( .A(AES_CORE_DATAPATH__abc_16259_n7647), .B(AES_CORE_DATAPATH__abc_16259_n6057_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n7648) );
  OR2X2 OR2X2_2363 ( .A(_auto_iopadmap_cc_313_execute_26916_31_), .B(AES_CORE_CONTROL_UNIT_last_round_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n7649) );
  OR2X2 OR2X2_2364 ( .A(AES_CORE_DATAPATH__abc_16259_n7647), .B(AES_CORE_DATAPATH__abc_16259_n6095_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n7652) );
  OR2X2 OR2X2_2365 ( .A(AES_CORE_DATAPATH__abc_16259_n6097_bF_buf3), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_31_), .Y(AES_CORE_DATAPATH__abc_16259_n7653) );
  OR2X2 OR2X2_2366 ( .A(AES_CORE_DATAPATH__abc_16259_n7655), .B(AES_CORE_DATAPATH__abc_16259_n7656), .Y(AES_CORE_DATAPATH__abc_16259_n7657) );
  OR2X2 OR2X2_2367 ( .A(AES_CORE_DATAPATH__abc_16259_n7657), .B(AES_CORE_DATAPATH__abc_16259_n7651), .Y(AES_CORE_DATAPATH__abc_16259_n7658) );
  OR2X2 OR2X2_2368 ( .A(AES_CORE_DATAPATH__abc_16259_n7659), .B(AES_CORE_DATAPATH__abc_16259_n7660), .Y(AES_CORE_DATAPATH__abc_16259_n7661) );
  OR2X2 OR2X2_2369 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf12), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_127_), .Y(AES_CORE_DATAPATH__abc_16259_n7662) );
  OR2X2 OR2X2_237 ( .A(AES_CORE_DATAPATH__abc_16259_n2835_1), .B(AES_CORE_DATAPATH__abc_16259_n2823), .Y(AES_CORE_DATAPATH__abc_16259_n2836) );
  OR2X2 OR2X2_2370 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf7), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_127_), .Y(AES_CORE_DATAPATH__abc_16259_n7663) );
  OR2X2 OR2X2_2371 ( .A(AES_CORE_DATAPATH__abc_16259_n7661), .B(AES_CORE_DATAPATH__abc_16259_n7665), .Y(AES_CORE_DATAPATH__abc_16259_n7666) );
  OR2X2 OR2X2_2372 ( .A(AES_CORE_DATAPATH__abc_16259_n7667), .B(AES_CORE_DATAPATH__abc_16259_n7620), .Y(AES_CORE_DATAPATH__0col_0__31_0__31_) );
  OR2X2 OR2X2_2373 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf11), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_96_), .Y(AES_CORE_DATAPATH__abc_16259_n7671) );
  OR2X2 OR2X2_2374 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf6), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_32_), .Y(AES_CORE_DATAPATH__abc_16259_n7672) );
  OR2X2 OR2X2_2375 ( .A(AES_CORE_DATAPATH__abc_16259_n6106), .B(AES_CORE_DATAPATH__abc_16259_n7674), .Y(AES_CORE_DATAPATH__abc_16259_n7675) );
  OR2X2 OR2X2_2376 ( .A(AES_CORE_DATAPATH__abc_16259_n7676), .B(AES_CORE_DATAPATH__abc_16259_n7670), .Y(AES_CORE_DATAPATH__0col_1__31_0__0_) );
  OR2X2 OR2X2_2377 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf10), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_97_), .Y(AES_CORE_DATAPATH__abc_16259_n7679) );
  OR2X2 OR2X2_2378 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf5), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_33_), .Y(AES_CORE_DATAPATH__abc_16259_n7680) );
  OR2X2 OR2X2_2379 ( .A(AES_CORE_DATAPATH__abc_16259_n6156), .B(AES_CORE_DATAPATH__abc_16259_n7682), .Y(AES_CORE_DATAPATH__abc_16259_n7683) );
  OR2X2 OR2X2_238 ( .A(AES_CORE_DATAPATH__abc_16259_n2831), .B(AES_CORE_DATAPATH__abc_16259_n2838), .Y(AES_CORE_DATAPATH__abc_16259_n2839_1) );
  OR2X2 OR2X2_2380 ( .A(AES_CORE_DATAPATH__abc_16259_n7684), .B(AES_CORE_DATAPATH__abc_16259_n7678), .Y(AES_CORE_DATAPATH__0col_1__31_0__1_) );
  OR2X2 OR2X2_2381 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf9), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_98_), .Y(AES_CORE_DATAPATH__abc_16259_n7687) );
  OR2X2 OR2X2_2382 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf4), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_34_), .Y(AES_CORE_DATAPATH__abc_16259_n7688) );
  OR2X2 OR2X2_2383 ( .A(AES_CORE_DATAPATH__abc_16259_n6205), .B(AES_CORE_DATAPATH__abc_16259_n7690), .Y(AES_CORE_DATAPATH__abc_16259_n7691) );
  OR2X2 OR2X2_2384 ( .A(AES_CORE_DATAPATH__abc_16259_n7692), .B(AES_CORE_DATAPATH__abc_16259_n7686), .Y(AES_CORE_DATAPATH__0col_1__31_0__2_) );
  OR2X2 OR2X2_2385 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf8), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_99_), .Y(AES_CORE_DATAPATH__abc_16259_n7695) );
  OR2X2 OR2X2_2386 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf3), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_35_), .Y(AES_CORE_DATAPATH__abc_16259_n7696) );
  OR2X2 OR2X2_2387 ( .A(AES_CORE_DATAPATH__abc_16259_n6254), .B(AES_CORE_DATAPATH__abc_16259_n7698), .Y(AES_CORE_DATAPATH__abc_16259_n7699) );
  OR2X2 OR2X2_2388 ( .A(AES_CORE_DATAPATH__abc_16259_n7700), .B(AES_CORE_DATAPATH__abc_16259_n7694), .Y(AES_CORE_DATAPATH__0col_1__31_0__3_) );
  OR2X2 OR2X2_2389 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf7), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_100_), .Y(AES_CORE_DATAPATH__abc_16259_n7703) );
  OR2X2 OR2X2_239 ( .A(AES_CORE_DATAPATH__abc_16259_n2839_1), .B(AES_CORE_DATAPATH__abc_16259_n2828), .Y(AES_CORE_DATAPATH__abc_16259_n2840) );
  OR2X2 OR2X2_2390 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf2), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_36_), .Y(AES_CORE_DATAPATH__abc_16259_n7704) );
  OR2X2 OR2X2_2391 ( .A(AES_CORE_DATAPATH__abc_16259_n6303), .B(AES_CORE_DATAPATH__abc_16259_n7706), .Y(AES_CORE_DATAPATH__abc_16259_n7707) );
  OR2X2 OR2X2_2392 ( .A(AES_CORE_DATAPATH__abc_16259_n7708), .B(AES_CORE_DATAPATH__abc_16259_n7702), .Y(AES_CORE_DATAPATH__0col_1__31_0__4_) );
  OR2X2 OR2X2_2393 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf6), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_101_), .Y(AES_CORE_DATAPATH__abc_16259_n7711) );
  OR2X2 OR2X2_2394 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf1), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_37_), .Y(AES_CORE_DATAPATH__abc_16259_n7712) );
  OR2X2 OR2X2_2395 ( .A(AES_CORE_DATAPATH__abc_16259_n6352), .B(AES_CORE_DATAPATH__abc_16259_n7714), .Y(AES_CORE_DATAPATH__abc_16259_n7715) );
  OR2X2 OR2X2_2396 ( .A(AES_CORE_DATAPATH__abc_16259_n7716), .B(AES_CORE_DATAPATH__abc_16259_n7710), .Y(AES_CORE_DATAPATH__0col_1__31_0__5_) );
  OR2X2 OR2X2_2397 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf5), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_102_), .Y(AES_CORE_DATAPATH__abc_16259_n7719) );
  OR2X2 OR2X2_2398 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf0), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_38_), .Y(AES_CORE_DATAPATH__abc_16259_n7720) );
  OR2X2 OR2X2_2399 ( .A(AES_CORE_DATAPATH__abc_16259_n6401), .B(AES_CORE_DATAPATH__abc_16259_n7722), .Y(AES_CORE_DATAPATH__abc_16259_n7723) );
  OR2X2 OR2X2_24 ( .A(AES_CORE_CONTROL_UNIT_state_8_), .B(AES_CORE_CONTROL_UNIT_state_6_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n140) );
  OR2X2 OR2X2_240 ( .A(AES_CORE_DATAPATH__abc_16259_n2841_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__0_), .Y(AES_CORE_DATAPATH__abc_16259_n2842) );
  OR2X2 OR2X2_2400 ( .A(AES_CORE_DATAPATH__abc_16259_n7724), .B(AES_CORE_DATAPATH__abc_16259_n7718), .Y(AES_CORE_DATAPATH__0col_1__31_0__6_) );
  OR2X2 OR2X2_2401 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf4), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_103_), .Y(AES_CORE_DATAPATH__abc_16259_n7727) );
  OR2X2 OR2X2_2402 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf14), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_39_), .Y(AES_CORE_DATAPATH__abc_16259_n7728) );
  OR2X2 OR2X2_2403 ( .A(AES_CORE_DATAPATH__abc_16259_n6450), .B(AES_CORE_DATAPATH__abc_16259_n7730), .Y(AES_CORE_DATAPATH__abc_16259_n7731) );
  OR2X2 OR2X2_2404 ( .A(AES_CORE_DATAPATH__abc_16259_n7732), .B(AES_CORE_DATAPATH__abc_16259_n7726), .Y(AES_CORE_DATAPATH__0col_1__31_0__7_) );
  OR2X2 OR2X2_2405 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf3), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_8_), .Y(AES_CORE_DATAPATH__abc_16259_n7735) );
  OR2X2 OR2X2_2406 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf13), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_8_), .Y(AES_CORE_DATAPATH__abc_16259_n7736) );
  OR2X2 OR2X2_2407 ( .A(AES_CORE_DATAPATH__abc_16259_n6499), .B(AES_CORE_DATAPATH__abc_16259_n7738), .Y(AES_CORE_DATAPATH__abc_16259_n7739) );
  OR2X2 OR2X2_2408 ( .A(AES_CORE_DATAPATH__abc_16259_n7740), .B(AES_CORE_DATAPATH__abc_16259_n7734), .Y(AES_CORE_DATAPATH__0col_1__31_0__8_) );
  OR2X2 OR2X2_2409 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf2), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_9_), .Y(AES_CORE_DATAPATH__abc_16259_n7743) );
  OR2X2 OR2X2_241 ( .A(AES_CORE_DATAPATH__abc_16259_n2844), .B(AES_CORE_DATAPATH__abc_16259_n2845), .Y(AES_CORE_DATAPATH__abc_16259_n2846) );
  OR2X2 OR2X2_2410 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf12), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_9_), .Y(AES_CORE_DATAPATH__abc_16259_n7744) );
  OR2X2 OR2X2_2411 ( .A(AES_CORE_DATAPATH__abc_16259_n6548), .B(AES_CORE_DATAPATH__abc_16259_n7746), .Y(AES_CORE_DATAPATH__abc_16259_n7747) );
  OR2X2 OR2X2_2412 ( .A(AES_CORE_DATAPATH__abc_16259_n7748), .B(AES_CORE_DATAPATH__abc_16259_n7742), .Y(AES_CORE_DATAPATH__0col_1__31_0__9_) );
  OR2X2 OR2X2_2413 ( .A(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf5), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_74_), .Y(AES_CORE_DATAPATH__abc_16259_n7750) );
  OR2X2 OR2X2_2414 ( .A(AES_CORE_DATAPATH__abc_16259_n7751), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf11), .Y(AES_CORE_DATAPATH__abc_16259_n7752) );
  OR2X2 OR2X2_2415 ( .A(AES_CORE_DATAPATH__abc_16259_n6603_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n7755), .Y(AES_CORE_DATAPATH__abc_16259_n7756) );
  OR2X2 OR2X2_2416 ( .A(AES_CORE_DATAPATH__abc_16259_n7761), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf9), .Y(AES_CORE_DATAPATH__abc_16259_n7762) );
  OR2X2 OR2X2_2417 ( .A(AES_CORE_DATAPATH__abc_16259_n6603_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n7765), .Y(AES_CORE_DATAPATH__abc_16259_n7766) );
  OR2X2 OR2X2_2418 ( .A(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf2), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_75_), .Y(AES_CORE_DATAPATH__abc_16259_n7770) );
  OR2X2 OR2X2_2419 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf1), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_12_), .Y(AES_CORE_DATAPATH__abc_16259_n7773) );
  OR2X2 OR2X2_242 ( .A(AES_CORE_DATAPATH__abc_16259_n2848), .B(AES_CORE_DATAPATH__abc_16259_n2849), .Y(AES_CORE_DATAPATH__abc_16259_n2850) );
  OR2X2 OR2X2_2420 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf7), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_12_), .Y(AES_CORE_DATAPATH__abc_16259_n7774) );
  OR2X2 OR2X2_2421 ( .A(AES_CORE_DATAPATH__abc_16259_n6710), .B(AES_CORE_DATAPATH__abc_16259_n7776), .Y(AES_CORE_DATAPATH__abc_16259_n7777) );
  OR2X2 OR2X2_2422 ( .A(AES_CORE_DATAPATH__abc_16259_n7778), .B(AES_CORE_DATAPATH__abc_16259_n7772), .Y(AES_CORE_DATAPATH__0col_1__31_0__12_) );
  OR2X2 OR2X2_2423 ( .A(AES_CORE_DATAPATH__abc_16259_n7780), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n7781) );
  OR2X2 OR2X2_2424 ( .A(AES_CORE_DATAPATH__abc_16259_n6603_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n7784), .Y(AES_CORE_DATAPATH__abc_16259_n7785) );
  OR2X2 OR2X2_2425 ( .A(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf5), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_77_), .Y(AES_CORE_DATAPATH__abc_16259_n7789) );
  OR2X2 OR2X2_2426 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf0), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_14_), .Y(AES_CORE_DATAPATH__abc_16259_n7792) );
  OR2X2 OR2X2_2427 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf4), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_14_), .Y(AES_CORE_DATAPATH__abc_16259_n7793) );
  OR2X2 OR2X2_2428 ( .A(AES_CORE_DATAPATH__abc_16259_n6813), .B(AES_CORE_DATAPATH__abc_16259_n7795), .Y(AES_CORE_DATAPATH__abc_16259_n7796) );
  OR2X2 OR2X2_2429 ( .A(AES_CORE_DATAPATH__abc_16259_n7797), .B(AES_CORE_DATAPATH__abc_16259_n7791), .Y(AES_CORE_DATAPATH__0col_1__31_0__14_) );
  OR2X2 OR2X2_243 ( .A(AES_CORE_DATAPATH__abc_16259_n2794), .B(AES_CORE_DATAPATH__abc_16259_n2853_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n2854) );
  OR2X2 OR2X2_2430 ( .A(AES_CORE_DATAPATH__abc_16259_n7799), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n7800) );
  OR2X2 OR2X2_2431 ( .A(AES_CORE_DATAPATH__abc_16259_n6603_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n7803), .Y(AES_CORE_DATAPATH__abc_16259_n7804) );
  OR2X2 OR2X2_2432 ( .A(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf2), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_79_), .Y(AES_CORE_DATAPATH__abc_16259_n7808) );
  OR2X2 OR2X2_2433 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf12), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_48_), .Y(AES_CORE_DATAPATH__abc_16259_n7811) );
  OR2X2 OR2X2_2434 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf1), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_112_), .Y(AES_CORE_DATAPATH__abc_16259_n7812) );
  OR2X2 OR2X2_2435 ( .A(AES_CORE_DATAPATH__abc_16259_n6916), .B(AES_CORE_DATAPATH__abc_16259_n7814), .Y(AES_CORE_DATAPATH__abc_16259_n7815) );
  OR2X2 OR2X2_2436 ( .A(AES_CORE_DATAPATH__abc_16259_n7816), .B(AES_CORE_DATAPATH__abc_16259_n7810), .Y(AES_CORE_DATAPATH__0col_1__31_0__16_) );
  OR2X2 OR2X2_2437 ( .A(AES_CORE_DATAPATH__abc_16259_n7818), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n7819) );
  OR2X2 OR2X2_2438 ( .A(AES_CORE_DATAPATH__abc_16259_n6603_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n7822), .Y(AES_CORE_DATAPATH__abc_16259_n7823) );
  OR2X2 OR2X2_2439 ( .A(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf5), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_81_), .Y(AES_CORE_DATAPATH__abc_16259_n7827) );
  OR2X2 OR2X2_244 ( .A(AES_CORE_DATAPATH__abc_16259_n2856), .B(AES_CORE_DATAPATH__abc_16259_n2858_1), .Y(AES_CORE_DATAPATH__abc_16259_n2859_1) );
  OR2X2 OR2X2_2440 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf11), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_50_), .Y(AES_CORE_DATAPATH__abc_16259_n7830) );
  OR2X2 OR2X2_2441 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf13), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_114_), .Y(AES_CORE_DATAPATH__abc_16259_n7831) );
  OR2X2 OR2X2_2442 ( .A(AES_CORE_DATAPATH__abc_16259_n7019), .B(AES_CORE_DATAPATH__abc_16259_n7833), .Y(AES_CORE_DATAPATH__abc_16259_n7834) );
  OR2X2 OR2X2_2443 ( .A(AES_CORE_DATAPATH__abc_16259_n7835), .B(AES_CORE_DATAPATH__abc_16259_n7829), .Y(AES_CORE_DATAPATH__0col_1__31_0__18_) );
  OR2X2 OR2X2_2444 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf10), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_51_), .Y(AES_CORE_DATAPATH__abc_16259_n7838) );
  OR2X2 OR2X2_2445 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf12), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_115_), .Y(AES_CORE_DATAPATH__abc_16259_n7839) );
  OR2X2 OR2X2_2446 ( .A(AES_CORE_DATAPATH__abc_16259_n7068), .B(AES_CORE_DATAPATH__abc_16259_n7841), .Y(AES_CORE_DATAPATH__abc_16259_n7842) );
  OR2X2 OR2X2_2447 ( .A(AES_CORE_DATAPATH__abc_16259_n7843), .B(AES_CORE_DATAPATH__abc_16259_n7837), .Y(AES_CORE_DATAPATH__0col_1__31_0__19_) );
  OR2X2 OR2X2_2448 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf9), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_52_), .Y(AES_CORE_DATAPATH__abc_16259_n7846) );
  OR2X2 OR2X2_2449 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf11), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_116_), .Y(AES_CORE_DATAPATH__abc_16259_n7847) );
  OR2X2 OR2X2_245 ( .A(_auto_iopadmap_cc_313_execute_26949_0_), .B(AES_CORE_DATAPATH__abc_16259_n2861), .Y(AES_CORE_DATAPATH__abc_16259_n2862_1) );
  OR2X2 OR2X2_2450 ( .A(AES_CORE_DATAPATH__abc_16259_n7117), .B(AES_CORE_DATAPATH__abc_16259_n7849), .Y(AES_CORE_DATAPATH__abc_16259_n7850) );
  OR2X2 OR2X2_2451 ( .A(AES_CORE_DATAPATH__abc_16259_n7851), .B(AES_CORE_DATAPATH__abc_16259_n7845), .Y(AES_CORE_DATAPATH__0col_1__31_0__20_) );
  OR2X2 OR2X2_2452 ( .A(AES_CORE_DATAPATH__abc_16259_n7853), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf10), .Y(AES_CORE_DATAPATH__abc_16259_n7854) );
  OR2X2 OR2X2_2453 ( .A(AES_CORE_DATAPATH__abc_16259_n6603_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n7857), .Y(AES_CORE_DATAPATH__abc_16259_n7858) );
  OR2X2 OR2X2_2454 ( .A(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf0), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_85_), .Y(AES_CORE_DATAPATH__abc_16259_n7862) );
  OR2X2 OR2X2_2455 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf8), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_54_), .Y(AES_CORE_DATAPATH__abc_16259_n7865) );
  OR2X2 OR2X2_2456 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf8), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_118_), .Y(AES_CORE_DATAPATH__abc_16259_n7866) );
  OR2X2 OR2X2_2457 ( .A(AES_CORE_DATAPATH__abc_16259_n7220), .B(AES_CORE_DATAPATH__abc_16259_n7868), .Y(AES_CORE_DATAPATH__abc_16259_n7869) );
  OR2X2 OR2X2_2458 ( .A(AES_CORE_DATAPATH__abc_16259_n7870), .B(AES_CORE_DATAPATH__abc_16259_n7864), .Y(AES_CORE_DATAPATH__0col_1__31_0__22_) );
  OR2X2 OR2X2_2459 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf7), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_55_), .Y(AES_CORE_DATAPATH__abc_16259_n7873) );
  OR2X2 OR2X2_246 ( .A(AES_CORE_DATAPATH__abc_16259_n2865), .B(AES_CORE_DATAPATH__abc_16259_n2864_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n2866_1) );
  OR2X2 OR2X2_2460 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf7), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_119_), .Y(AES_CORE_DATAPATH__abc_16259_n7874) );
  OR2X2 OR2X2_2461 ( .A(AES_CORE_DATAPATH__abc_16259_n7269), .B(AES_CORE_DATAPATH__abc_16259_n7876), .Y(AES_CORE_DATAPATH__abc_16259_n7877) );
  OR2X2 OR2X2_2462 ( .A(AES_CORE_DATAPATH__abc_16259_n7878), .B(AES_CORE_DATAPATH__abc_16259_n7872), .Y(AES_CORE_DATAPATH__0col_1__31_0__23_) );
  OR2X2 OR2X2_2463 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf6), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_88_), .Y(AES_CORE_DATAPATH__abc_16259_n7881) );
  OR2X2 OR2X2_2464 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf6), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_88_), .Y(AES_CORE_DATAPATH__abc_16259_n7882) );
  OR2X2 OR2X2_2465 ( .A(AES_CORE_DATAPATH__abc_16259_n7318), .B(AES_CORE_DATAPATH__abc_16259_n7884), .Y(AES_CORE_DATAPATH__abc_16259_n7885) );
  OR2X2 OR2X2_2466 ( .A(AES_CORE_DATAPATH__abc_16259_n7886), .B(AES_CORE_DATAPATH__abc_16259_n7880), .Y(AES_CORE_DATAPATH__0col_1__31_0__24_) );
  OR2X2 OR2X2_2467 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf5), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_89_), .Y(AES_CORE_DATAPATH__abc_16259_n7889) );
  OR2X2 OR2X2_2468 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf5), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_89_), .Y(AES_CORE_DATAPATH__abc_16259_n7890) );
  OR2X2 OR2X2_2469 ( .A(AES_CORE_DATAPATH__abc_16259_n7367), .B(AES_CORE_DATAPATH__abc_16259_n7892), .Y(AES_CORE_DATAPATH__abc_16259_n7893) );
  OR2X2 OR2X2_247 ( .A(AES_CORE_DATAPATH__abc_16259_n2866_1), .B(AES_CORE_DATAPATH__abc_16259_n2863), .Y(AES_CORE_DATAPATH__abc_16259_n2867) );
  OR2X2 OR2X2_2470 ( .A(AES_CORE_DATAPATH__abc_16259_n7894), .B(AES_CORE_DATAPATH__abc_16259_n7888), .Y(AES_CORE_DATAPATH__0col_1__31_0__25_) );
  OR2X2 OR2X2_2471 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf4), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_90_), .Y(AES_CORE_DATAPATH__abc_16259_n7897) );
  OR2X2 OR2X2_2472 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf4), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_90_), .Y(AES_CORE_DATAPATH__abc_16259_n7898) );
  OR2X2 OR2X2_2473 ( .A(AES_CORE_DATAPATH__abc_16259_n7416), .B(AES_CORE_DATAPATH__abc_16259_n7900), .Y(AES_CORE_DATAPATH__abc_16259_n7901) );
  OR2X2 OR2X2_2474 ( .A(AES_CORE_DATAPATH__abc_16259_n7902), .B(AES_CORE_DATAPATH__abc_16259_n7896), .Y(AES_CORE_DATAPATH__0col_1__31_0__26_) );
  OR2X2 OR2X2_2475 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf3), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_91_), .Y(AES_CORE_DATAPATH__abc_16259_n7905) );
  OR2X2 OR2X2_2476 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf3), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_91_), .Y(AES_CORE_DATAPATH__abc_16259_n7906) );
  OR2X2 OR2X2_2477 ( .A(AES_CORE_DATAPATH__abc_16259_n7465), .B(AES_CORE_DATAPATH__abc_16259_n7908), .Y(AES_CORE_DATAPATH__abc_16259_n7909) );
  OR2X2 OR2X2_2478 ( .A(AES_CORE_DATAPATH__abc_16259_n7910), .B(AES_CORE_DATAPATH__abc_16259_n7904), .Y(AES_CORE_DATAPATH__0col_1__31_0__27_) );
  OR2X2 OR2X2_2479 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf2), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_92_), .Y(AES_CORE_DATAPATH__abc_16259_n7913) );
  OR2X2 OR2X2_248 ( .A(AES_CORE_DATAPATH__abc_16259_n2869), .B(AES_CORE_DATAPATH__abc_16259_n2870), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_0_) );
  OR2X2 OR2X2_2480 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf2), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_92_), .Y(AES_CORE_DATAPATH__abc_16259_n7914) );
  OR2X2 OR2X2_2481 ( .A(AES_CORE_DATAPATH__abc_16259_n7514), .B(AES_CORE_DATAPATH__abc_16259_n7916), .Y(AES_CORE_DATAPATH__abc_16259_n7917) );
  OR2X2 OR2X2_2482 ( .A(AES_CORE_DATAPATH__abc_16259_n7918), .B(AES_CORE_DATAPATH__abc_16259_n7912), .Y(AES_CORE_DATAPATH__0col_1__31_0__28_) );
  OR2X2 OR2X2_2483 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf1), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_93_), .Y(AES_CORE_DATAPATH__abc_16259_n7921) );
  OR2X2 OR2X2_2484 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf1), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_93_), .Y(AES_CORE_DATAPATH__abc_16259_n7922) );
  OR2X2 OR2X2_2485 ( .A(AES_CORE_DATAPATH__abc_16259_n7563), .B(AES_CORE_DATAPATH__abc_16259_n7924), .Y(AES_CORE_DATAPATH__abc_16259_n7925) );
  OR2X2 OR2X2_2486 ( .A(AES_CORE_DATAPATH__abc_16259_n7926), .B(AES_CORE_DATAPATH__abc_16259_n7920), .Y(AES_CORE_DATAPATH__0col_1__31_0__29_) );
  OR2X2 OR2X2_2487 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf0), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_94_), .Y(AES_CORE_DATAPATH__abc_16259_n7929) );
  OR2X2 OR2X2_2488 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf0), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_94_), .Y(AES_CORE_DATAPATH__abc_16259_n7930) );
  OR2X2 OR2X2_2489 ( .A(AES_CORE_DATAPATH__abc_16259_n7612), .B(AES_CORE_DATAPATH__abc_16259_n7932), .Y(AES_CORE_DATAPATH__abc_16259_n7933) );
  OR2X2 OR2X2_249 ( .A(AES_CORE_DATAPATH__abc_16259_n2774_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n2872), .Y(AES_CORE_DATAPATH__abc_16259_n2873) );
  OR2X2 OR2X2_2490 ( .A(AES_CORE_DATAPATH__abc_16259_n7934), .B(AES_CORE_DATAPATH__abc_16259_n7928), .Y(AES_CORE_DATAPATH__0col_1__31_0__30_) );
  OR2X2 OR2X2_2491 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf12), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_95_), .Y(AES_CORE_DATAPATH__abc_16259_n7937) );
  OR2X2 OR2X2_2492 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf14), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_95_), .Y(AES_CORE_DATAPATH__abc_16259_n7938) );
  OR2X2 OR2X2_2493 ( .A(AES_CORE_DATAPATH__abc_16259_n7661), .B(AES_CORE_DATAPATH__abc_16259_n7940), .Y(AES_CORE_DATAPATH__abc_16259_n7941) );
  OR2X2 OR2X2_2494 ( .A(AES_CORE_DATAPATH__abc_16259_n7942), .B(AES_CORE_DATAPATH__abc_16259_n7936), .Y(AES_CORE_DATAPATH__0col_1__31_0__31_) );
  OR2X2 OR2X2_2495 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf11), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_64_), .Y(AES_CORE_DATAPATH__abc_16259_n7946) );
  OR2X2 OR2X2_2496 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf13), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_0_), .Y(AES_CORE_DATAPATH__abc_16259_n7947) );
  OR2X2 OR2X2_2497 ( .A(AES_CORE_DATAPATH__abc_16259_n6106), .B(AES_CORE_DATAPATH__abc_16259_n7949), .Y(AES_CORE_DATAPATH__abc_16259_n7950) );
  OR2X2 OR2X2_2498 ( .A(AES_CORE_DATAPATH__abc_16259_n7951), .B(AES_CORE_DATAPATH__abc_16259_n7945), .Y(AES_CORE_DATAPATH__0col_2__31_0__0_) );
  OR2X2 OR2X2_2499 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf10), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_65_), .Y(AES_CORE_DATAPATH__abc_16259_n7954) );
  OR2X2 OR2X2_25 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n143), .B(AES_CORE_CONTROL_UNIT_state_2_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n144) );
  OR2X2 OR2X2_250 ( .A(AES_CORE_DATAPATH__abc_16259_n2778_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n2874), .Y(AES_CORE_DATAPATH__abc_16259_n2875) );
  OR2X2 OR2X2_2500 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf12), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_1_), .Y(AES_CORE_DATAPATH__abc_16259_n7955) );
  OR2X2 OR2X2_2501 ( .A(AES_CORE_DATAPATH__abc_16259_n6156), .B(AES_CORE_DATAPATH__abc_16259_n7957), .Y(AES_CORE_DATAPATH__abc_16259_n7958) );
  OR2X2 OR2X2_2502 ( .A(AES_CORE_DATAPATH__abc_16259_n7959), .B(AES_CORE_DATAPATH__abc_16259_n7953), .Y(AES_CORE_DATAPATH__0col_2__31_0__1_) );
  OR2X2 OR2X2_2503 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf9), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_66_), .Y(AES_CORE_DATAPATH__abc_16259_n7962) );
  OR2X2 OR2X2_2504 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf11), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_2_), .Y(AES_CORE_DATAPATH__abc_16259_n7963) );
  OR2X2 OR2X2_2505 ( .A(AES_CORE_DATAPATH__abc_16259_n6205), .B(AES_CORE_DATAPATH__abc_16259_n7965), .Y(AES_CORE_DATAPATH__abc_16259_n7966) );
  OR2X2 OR2X2_2506 ( .A(AES_CORE_DATAPATH__abc_16259_n7967), .B(AES_CORE_DATAPATH__abc_16259_n7961), .Y(AES_CORE_DATAPATH__0col_2__31_0__2_) );
  OR2X2 OR2X2_2507 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf8), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_67_), .Y(AES_CORE_DATAPATH__abc_16259_n7970) );
  OR2X2 OR2X2_2508 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf10), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_3_), .Y(AES_CORE_DATAPATH__abc_16259_n7971) );
  OR2X2 OR2X2_2509 ( .A(AES_CORE_DATAPATH__abc_16259_n6254), .B(AES_CORE_DATAPATH__abc_16259_n7973), .Y(AES_CORE_DATAPATH__abc_16259_n7974) );
  OR2X2 OR2X2_251 ( .A(AES_CORE_DATAPATH__abc_16259_n2878), .B(AES_CORE_DATAPATH__abc_16259_n2879), .Y(AES_CORE_DATAPATH__abc_16259_n2880_1) );
  OR2X2 OR2X2_2510 ( .A(AES_CORE_DATAPATH__abc_16259_n7975), .B(AES_CORE_DATAPATH__abc_16259_n7969), .Y(AES_CORE_DATAPATH__0col_2__31_0__3_) );
  OR2X2 OR2X2_2511 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf7), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_68_), .Y(AES_CORE_DATAPATH__abc_16259_n7978) );
  OR2X2 OR2X2_2512 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf9), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_4_), .Y(AES_CORE_DATAPATH__abc_16259_n7979) );
  OR2X2 OR2X2_2513 ( .A(AES_CORE_DATAPATH__abc_16259_n6303), .B(AES_CORE_DATAPATH__abc_16259_n7981), .Y(AES_CORE_DATAPATH__abc_16259_n7982) );
  OR2X2 OR2X2_2514 ( .A(AES_CORE_DATAPATH__abc_16259_n7983), .B(AES_CORE_DATAPATH__abc_16259_n7977), .Y(AES_CORE_DATAPATH__0col_2__31_0__4_) );
  OR2X2 OR2X2_2515 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf6), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_69_), .Y(AES_CORE_DATAPATH__abc_16259_n7986) );
  OR2X2 OR2X2_2516 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf8), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_5_), .Y(AES_CORE_DATAPATH__abc_16259_n7987) );
  OR2X2 OR2X2_2517 ( .A(AES_CORE_DATAPATH__abc_16259_n6352), .B(AES_CORE_DATAPATH__abc_16259_n7989), .Y(AES_CORE_DATAPATH__abc_16259_n7990) );
  OR2X2 OR2X2_2518 ( .A(AES_CORE_DATAPATH__abc_16259_n7991), .B(AES_CORE_DATAPATH__abc_16259_n7985), .Y(AES_CORE_DATAPATH__0col_2__31_0__5_) );
  OR2X2 OR2X2_2519 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf5), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_70_), .Y(AES_CORE_DATAPATH__abc_16259_n7994) );
  OR2X2 OR2X2_252 ( .A(AES_CORE_DATAPATH__abc_16259_n2880_1), .B(AES_CORE_DATAPATH__abc_16259_n2877), .Y(AES_CORE_DATAPATH__abc_16259_n2881) );
  OR2X2 OR2X2_2520 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf7), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_6_), .Y(AES_CORE_DATAPATH__abc_16259_n7995) );
  OR2X2 OR2X2_2521 ( .A(AES_CORE_DATAPATH__abc_16259_n6401), .B(AES_CORE_DATAPATH__abc_16259_n7997), .Y(AES_CORE_DATAPATH__abc_16259_n7998) );
  OR2X2 OR2X2_2522 ( .A(AES_CORE_DATAPATH__abc_16259_n7999), .B(AES_CORE_DATAPATH__abc_16259_n7993), .Y(AES_CORE_DATAPATH__0col_2__31_0__6_) );
  OR2X2 OR2X2_2523 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf4), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_71_), .Y(AES_CORE_DATAPATH__abc_16259_n8002) );
  OR2X2 OR2X2_2524 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf6), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_7_), .Y(AES_CORE_DATAPATH__abc_16259_n8003) );
  OR2X2 OR2X2_2525 ( .A(AES_CORE_DATAPATH__abc_16259_n6450), .B(AES_CORE_DATAPATH__abc_16259_n8005), .Y(AES_CORE_DATAPATH__abc_16259_n8006) );
  OR2X2 OR2X2_2526 ( .A(AES_CORE_DATAPATH__abc_16259_n8007), .B(AES_CORE_DATAPATH__abc_16259_n8001), .Y(AES_CORE_DATAPATH__0col_2__31_0__7_) );
  OR2X2 OR2X2_2527 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf3), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_104_), .Y(AES_CORE_DATAPATH__abc_16259_n8010) );
  OR2X2 OR2X2_2528 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf5), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_104_), .Y(AES_CORE_DATAPATH__abc_16259_n8011) );
  OR2X2 OR2X2_2529 ( .A(AES_CORE_DATAPATH__abc_16259_n6499), .B(AES_CORE_DATAPATH__abc_16259_n8013), .Y(AES_CORE_DATAPATH__abc_16259_n8014) );
  OR2X2 OR2X2_253 ( .A(AES_CORE_DATAPATH__abc_16259_n2885), .B(AES_CORE_DATAPATH__abc_16259_n2826_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n2886) );
  OR2X2 OR2X2_2530 ( .A(AES_CORE_DATAPATH__abc_16259_n8015), .B(AES_CORE_DATAPATH__abc_16259_n8009), .Y(AES_CORE_DATAPATH__0col_2__31_0__8_) );
  OR2X2 OR2X2_2531 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf2), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_105_), .Y(AES_CORE_DATAPATH__abc_16259_n8018) );
  OR2X2 OR2X2_2532 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf4), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_105_), .Y(AES_CORE_DATAPATH__abc_16259_n8019) );
  OR2X2 OR2X2_2533 ( .A(AES_CORE_DATAPATH__abc_16259_n6548), .B(AES_CORE_DATAPATH__abc_16259_n8021), .Y(AES_CORE_DATAPATH__abc_16259_n8022) );
  OR2X2 OR2X2_2534 ( .A(AES_CORE_DATAPATH__abc_16259_n8023), .B(AES_CORE_DATAPATH__abc_16259_n8017), .Y(AES_CORE_DATAPATH__0col_2__31_0__9_) );
  OR2X2 OR2X2_2535 ( .A(AES_CORE_DATAPATH__abc_16259_n8025), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n8026) );
  OR2X2 OR2X2_2536 ( .A(AES_CORE_DATAPATH__abc_16259_n6603_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n8029), .Y(AES_CORE_DATAPATH__abc_16259_n8030) );
  OR2X2 OR2X2_2537 ( .A(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf4), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_42_), .Y(AES_CORE_DATAPATH__abc_16259_n8034) );
  OR2X2 OR2X2_2538 ( .A(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf3), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_43_), .Y(AES_CORE_DATAPATH__abc_16259_n8036) );
  OR2X2 OR2X2_2539 ( .A(AES_CORE_DATAPATH__abc_16259_n8037), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n8038) );
  OR2X2 OR2X2_254 ( .A(AES_CORE_DATAPATH__abc_16259_n2888_1), .B(AES_CORE_DATAPATH__abc_16259_n2889), .Y(AES_CORE_DATAPATH__abc_16259_n2890) );
  OR2X2 OR2X2_2540 ( .A(AES_CORE_DATAPATH__abc_16259_n6603_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n8041), .Y(AES_CORE_DATAPATH__abc_16259_n8042) );
  OR2X2 OR2X2_2541 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf1), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_108_), .Y(AES_CORE_DATAPATH__abc_16259_n8048) );
  OR2X2 OR2X2_2542 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf14), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_108_), .Y(AES_CORE_DATAPATH__abc_16259_n8049) );
  OR2X2 OR2X2_2543 ( .A(AES_CORE_DATAPATH__abc_16259_n6710), .B(AES_CORE_DATAPATH__abc_16259_n8051), .Y(AES_CORE_DATAPATH__abc_16259_n8052) );
  OR2X2 OR2X2_2544 ( .A(AES_CORE_DATAPATH__abc_16259_n8053), .B(AES_CORE_DATAPATH__abc_16259_n8047), .Y(AES_CORE_DATAPATH__0col_2__31_0__12_) );
  OR2X2 OR2X2_2545 ( .A(AES_CORE_DATAPATH__abc_16259_n8055), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf13), .Y(AES_CORE_DATAPATH__abc_16259_n8056) );
  OR2X2 OR2X2_2546 ( .A(AES_CORE_DATAPATH__abc_16259_n6603_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n8059), .Y(AES_CORE_DATAPATH__abc_16259_n8060) );
  OR2X2 OR2X2_2547 ( .A(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf5), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_45_), .Y(AES_CORE_DATAPATH__abc_16259_n8064) );
  OR2X2 OR2X2_2548 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf0), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_110_), .Y(AES_CORE_DATAPATH__abc_16259_n8067) );
  OR2X2 OR2X2_2549 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf11), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_110_), .Y(AES_CORE_DATAPATH__abc_16259_n8068) );
  OR2X2 OR2X2_255 ( .A(AES_CORE_DATAPATH__abc_16259_n2890), .B(AES_CORE_DATAPATH__abc_16259_n2886), .Y(AES_CORE_DATAPATH__abc_16259_n2891_1) );
  OR2X2 OR2X2_2550 ( .A(AES_CORE_DATAPATH__abc_16259_n6813), .B(AES_CORE_DATAPATH__abc_16259_n8070), .Y(AES_CORE_DATAPATH__abc_16259_n8071) );
  OR2X2 OR2X2_2551 ( .A(AES_CORE_DATAPATH__abc_16259_n8072), .B(AES_CORE_DATAPATH__abc_16259_n8066), .Y(AES_CORE_DATAPATH__0col_2__31_0__14_) );
  OR2X2 OR2X2_2552 ( .A(AES_CORE_DATAPATH__abc_16259_n8074), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf10), .Y(AES_CORE_DATAPATH__abc_16259_n8075) );
  OR2X2 OR2X2_2553 ( .A(AES_CORE_DATAPATH__abc_16259_n6603_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n8078), .Y(AES_CORE_DATAPATH__abc_16259_n8079) );
  OR2X2 OR2X2_2554 ( .A(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf2), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_47_), .Y(AES_CORE_DATAPATH__abc_16259_n8083) );
  OR2X2 OR2X2_2555 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf12), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_16_), .Y(AES_CORE_DATAPATH__abc_16259_n8086) );
  OR2X2 OR2X2_2556 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf8), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_80_), .Y(AES_CORE_DATAPATH__abc_16259_n8087) );
  OR2X2 OR2X2_2557 ( .A(AES_CORE_DATAPATH__abc_16259_n6916), .B(AES_CORE_DATAPATH__abc_16259_n8089), .Y(AES_CORE_DATAPATH__abc_16259_n8090) );
  OR2X2 OR2X2_2558 ( .A(AES_CORE_DATAPATH__abc_16259_n8091), .B(AES_CORE_DATAPATH__abc_16259_n8085), .Y(AES_CORE_DATAPATH__0col_2__31_0__16_) );
  OR2X2 OR2X2_2559 ( .A(AES_CORE_DATAPATH__abc_16259_n8093), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n8094) );
  OR2X2 OR2X2_256 ( .A(AES_CORE_DATAPATH__abc_16259_n2841_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__1_), .Y(AES_CORE_DATAPATH__abc_16259_n2892) );
  OR2X2 OR2X2_2560 ( .A(AES_CORE_DATAPATH__abc_16259_n6603_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n8097), .Y(AES_CORE_DATAPATH__abc_16259_n8098) );
  OR2X2 OR2X2_2561 ( .A(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf5), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_49_), .Y(AES_CORE_DATAPATH__abc_16259_n8102) );
  OR2X2 OR2X2_2562 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf11), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_18_), .Y(AES_CORE_DATAPATH__abc_16259_n8105) );
  OR2X2 OR2X2_2563 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf5), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_82_), .Y(AES_CORE_DATAPATH__abc_16259_n8106) );
  OR2X2 OR2X2_2564 ( .A(AES_CORE_DATAPATH__abc_16259_n7019), .B(AES_CORE_DATAPATH__abc_16259_n8108), .Y(AES_CORE_DATAPATH__abc_16259_n8109) );
  OR2X2 OR2X2_2565 ( .A(AES_CORE_DATAPATH__abc_16259_n8110), .B(AES_CORE_DATAPATH__abc_16259_n8104), .Y(AES_CORE_DATAPATH__0col_2__31_0__18_) );
  OR2X2 OR2X2_2566 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf10), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_19_), .Y(AES_CORE_DATAPATH__abc_16259_n8113) );
  OR2X2 OR2X2_2567 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf4), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_83_), .Y(AES_CORE_DATAPATH__abc_16259_n8114) );
  OR2X2 OR2X2_2568 ( .A(AES_CORE_DATAPATH__abc_16259_n7068), .B(AES_CORE_DATAPATH__abc_16259_n8116), .Y(AES_CORE_DATAPATH__abc_16259_n8117) );
  OR2X2 OR2X2_2569 ( .A(AES_CORE_DATAPATH__abc_16259_n8118), .B(AES_CORE_DATAPATH__abc_16259_n8112), .Y(AES_CORE_DATAPATH__0col_2__31_0__19_) );
  OR2X2 OR2X2_257 ( .A(AES_CORE_DATAPATH__abc_16259_n2883), .B(AES_CORE_DATAPATH__abc_16259_n2853_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n2894) );
  OR2X2 OR2X2_2570 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf9), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_20_), .Y(AES_CORE_DATAPATH__abc_16259_n8121) );
  OR2X2 OR2X2_2571 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf3), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_84_), .Y(AES_CORE_DATAPATH__abc_16259_n8122) );
  OR2X2 OR2X2_2572 ( .A(AES_CORE_DATAPATH__abc_16259_n7117), .B(AES_CORE_DATAPATH__abc_16259_n8124), .Y(AES_CORE_DATAPATH__abc_16259_n8125) );
  OR2X2 OR2X2_2573 ( .A(AES_CORE_DATAPATH__abc_16259_n8126), .B(AES_CORE_DATAPATH__abc_16259_n8120), .Y(AES_CORE_DATAPATH__0col_2__31_0__20_) );
  OR2X2 OR2X2_2574 ( .A(AES_CORE_DATAPATH__abc_16259_n8128), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n8129) );
  OR2X2 OR2X2_2575 ( .A(AES_CORE_DATAPATH__abc_16259_n6603_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n8132), .Y(AES_CORE_DATAPATH__abc_16259_n8133) );
  OR2X2 OR2X2_2576 ( .A(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf0), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_53_), .Y(AES_CORE_DATAPATH__abc_16259_n8137) );
  OR2X2 OR2X2_2577 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf8), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_22_), .Y(AES_CORE_DATAPATH__abc_16259_n8140) );
  OR2X2 OR2X2_2578 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf0), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_86_), .Y(AES_CORE_DATAPATH__abc_16259_n8141) );
  OR2X2 OR2X2_2579 ( .A(AES_CORE_DATAPATH__abc_16259_n7220), .B(AES_CORE_DATAPATH__abc_16259_n8143), .Y(AES_CORE_DATAPATH__abc_16259_n8144) );
  OR2X2 OR2X2_258 ( .A(AES_CORE_DATAPATH__abc_16259_n2895_1), .B(AES_CORE_DATAPATH__abc_16259_n2896), .Y(AES_CORE_DATAPATH__abc_16259_n2897_1) );
  OR2X2 OR2X2_2580 ( .A(AES_CORE_DATAPATH__abc_16259_n8145), .B(AES_CORE_DATAPATH__abc_16259_n8139), .Y(AES_CORE_DATAPATH__0col_2__31_0__22_) );
  OR2X2 OR2X2_2581 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf7), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_23_), .Y(AES_CORE_DATAPATH__abc_16259_n8148) );
  OR2X2 OR2X2_2582 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf14), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_87_), .Y(AES_CORE_DATAPATH__abc_16259_n8149) );
  OR2X2 OR2X2_2583 ( .A(AES_CORE_DATAPATH__abc_16259_n7269), .B(AES_CORE_DATAPATH__abc_16259_n8151), .Y(AES_CORE_DATAPATH__abc_16259_n8152) );
  OR2X2 OR2X2_2584 ( .A(AES_CORE_DATAPATH__abc_16259_n8153), .B(AES_CORE_DATAPATH__abc_16259_n8147), .Y(AES_CORE_DATAPATH__0col_2__31_0__23_) );
  OR2X2 OR2X2_2585 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf6), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_56_), .Y(AES_CORE_DATAPATH__abc_16259_n8156) );
  OR2X2 OR2X2_2586 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf13), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_56_), .Y(AES_CORE_DATAPATH__abc_16259_n8157) );
  OR2X2 OR2X2_2587 ( .A(AES_CORE_DATAPATH__abc_16259_n7318), .B(AES_CORE_DATAPATH__abc_16259_n8159), .Y(AES_CORE_DATAPATH__abc_16259_n8160) );
  OR2X2 OR2X2_2588 ( .A(AES_CORE_DATAPATH__abc_16259_n8161), .B(AES_CORE_DATAPATH__abc_16259_n8155), .Y(AES_CORE_DATAPATH__0col_2__31_0__24_) );
  OR2X2 OR2X2_2589 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf5), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_57_), .Y(AES_CORE_DATAPATH__abc_16259_n8164) );
  OR2X2 OR2X2_259 ( .A(_auto_iopadmap_cc_313_execute_26949_1_), .B(AES_CORE_DATAPATH__abc_16259_n2899), .Y(AES_CORE_DATAPATH__abc_16259_n2900) );
  OR2X2 OR2X2_2590 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf12), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_57_), .Y(AES_CORE_DATAPATH__abc_16259_n8165) );
  OR2X2 OR2X2_2591 ( .A(AES_CORE_DATAPATH__abc_16259_n7367), .B(AES_CORE_DATAPATH__abc_16259_n8167), .Y(AES_CORE_DATAPATH__abc_16259_n8168) );
  OR2X2 OR2X2_2592 ( .A(AES_CORE_DATAPATH__abc_16259_n8169), .B(AES_CORE_DATAPATH__abc_16259_n8163), .Y(AES_CORE_DATAPATH__0col_2__31_0__25_) );
  OR2X2 OR2X2_2593 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf4), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_58_), .Y(AES_CORE_DATAPATH__abc_16259_n8172) );
  OR2X2 OR2X2_2594 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf11), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_58_), .Y(AES_CORE_DATAPATH__abc_16259_n8173) );
  OR2X2 OR2X2_2595 ( .A(AES_CORE_DATAPATH__abc_16259_n7416), .B(AES_CORE_DATAPATH__abc_16259_n8175), .Y(AES_CORE_DATAPATH__abc_16259_n8176) );
  OR2X2 OR2X2_2596 ( .A(AES_CORE_DATAPATH__abc_16259_n8177), .B(AES_CORE_DATAPATH__abc_16259_n8171), .Y(AES_CORE_DATAPATH__0col_2__31_0__26_) );
  OR2X2 OR2X2_2597 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf3), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_59_), .Y(AES_CORE_DATAPATH__abc_16259_n8180) );
  OR2X2 OR2X2_2598 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf10), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_59_), .Y(AES_CORE_DATAPATH__abc_16259_n8181) );
  OR2X2 OR2X2_2599 ( .A(AES_CORE_DATAPATH__abc_16259_n7465), .B(AES_CORE_DATAPATH__abc_16259_n8183), .Y(AES_CORE_DATAPATH__abc_16259_n8184) );
  OR2X2 OR2X2_26 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n145), .B(AES_CORE_CONTROL_UNIT__abc_15841_n141_1), .Y(AES_CORE_CONTROL_UNIT__abc_10818_n97) );
  OR2X2 OR2X2_260 ( .A(AES_CORE_DATAPATH__abc_16259_n2902), .B(AES_CORE_DATAPATH__abc_16259_n2864_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n2903) );
  OR2X2 OR2X2_2600 ( .A(AES_CORE_DATAPATH__abc_16259_n8185), .B(AES_CORE_DATAPATH__abc_16259_n8179), .Y(AES_CORE_DATAPATH__0col_2__31_0__27_) );
  OR2X2 OR2X2_2601 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf2), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_60_), .Y(AES_CORE_DATAPATH__abc_16259_n8188) );
  OR2X2 OR2X2_2602 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf9), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_60_), .Y(AES_CORE_DATAPATH__abc_16259_n8189) );
  OR2X2 OR2X2_2603 ( .A(AES_CORE_DATAPATH__abc_16259_n7514), .B(AES_CORE_DATAPATH__abc_16259_n8191), .Y(AES_CORE_DATAPATH__abc_16259_n8192) );
  OR2X2 OR2X2_2604 ( .A(AES_CORE_DATAPATH__abc_16259_n8193), .B(AES_CORE_DATAPATH__abc_16259_n8187), .Y(AES_CORE_DATAPATH__0col_2__31_0__28_) );
  OR2X2 OR2X2_2605 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf1), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_61_), .Y(AES_CORE_DATAPATH__abc_16259_n8196) );
  OR2X2 OR2X2_2606 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf8), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_61_), .Y(AES_CORE_DATAPATH__abc_16259_n8197) );
  OR2X2 OR2X2_2607 ( .A(AES_CORE_DATAPATH__abc_16259_n7563), .B(AES_CORE_DATAPATH__abc_16259_n8199), .Y(AES_CORE_DATAPATH__abc_16259_n8200) );
  OR2X2 OR2X2_2608 ( .A(AES_CORE_DATAPATH__abc_16259_n8201), .B(AES_CORE_DATAPATH__abc_16259_n8195), .Y(AES_CORE_DATAPATH__0col_2__31_0__29_) );
  OR2X2 OR2X2_2609 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf0), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_62_), .Y(AES_CORE_DATAPATH__abc_16259_n8204) );
  OR2X2 OR2X2_261 ( .A(AES_CORE_DATAPATH__abc_16259_n2903), .B(AES_CORE_DATAPATH__abc_16259_n2901), .Y(AES_CORE_DATAPATH__abc_16259_n2904) );
  OR2X2 OR2X2_2610 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf7), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_62_), .Y(AES_CORE_DATAPATH__abc_16259_n8205) );
  OR2X2 OR2X2_2611 ( .A(AES_CORE_DATAPATH__abc_16259_n7612), .B(AES_CORE_DATAPATH__abc_16259_n8207), .Y(AES_CORE_DATAPATH__abc_16259_n8208) );
  OR2X2 OR2X2_2612 ( .A(AES_CORE_DATAPATH__abc_16259_n8209), .B(AES_CORE_DATAPATH__abc_16259_n8203), .Y(AES_CORE_DATAPATH__0col_2__31_0__30_) );
  OR2X2 OR2X2_2613 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf12), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_63_), .Y(AES_CORE_DATAPATH__abc_16259_n8212) );
  OR2X2 OR2X2_2614 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf6), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_63_), .Y(AES_CORE_DATAPATH__abc_16259_n8213) );
  OR2X2 OR2X2_2615 ( .A(AES_CORE_DATAPATH__abc_16259_n7661), .B(AES_CORE_DATAPATH__abc_16259_n8215), .Y(AES_CORE_DATAPATH__abc_16259_n8216) );
  OR2X2 OR2X2_2616 ( .A(AES_CORE_DATAPATH__abc_16259_n8217), .B(AES_CORE_DATAPATH__abc_16259_n8211), .Y(AES_CORE_DATAPATH__0col_2__31_0__31_) );
  OR2X2 OR2X2_2617 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf11), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_32_), .Y(AES_CORE_DATAPATH__abc_16259_n8221) );
  OR2X2 OR2X2_2618 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf5), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_96_), .Y(AES_CORE_DATAPATH__abc_16259_n8222) );
  OR2X2 OR2X2_2619 ( .A(AES_CORE_DATAPATH__abc_16259_n6106), .B(AES_CORE_DATAPATH__abc_16259_n8224), .Y(AES_CORE_DATAPATH__abc_16259_n8225) );
  OR2X2 OR2X2_262 ( .A(AES_CORE_DATAPATH__abc_16259_n2906), .B(AES_CORE_DATAPATH__abc_16259_n2905), .Y(AES_CORE_DATAPATH__abc_16259_n2907) );
  OR2X2 OR2X2_2620 ( .A(AES_CORE_DATAPATH__abc_16259_n8226), .B(AES_CORE_DATAPATH__abc_16259_n8220), .Y(AES_CORE_DATAPATH__0col_3__31_0__0_) );
  OR2X2 OR2X2_2621 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf10), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_33_), .Y(AES_CORE_DATAPATH__abc_16259_n8229) );
  OR2X2 OR2X2_2622 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf4), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_97_), .Y(AES_CORE_DATAPATH__abc_16259_n8230) );
  OR2X2 OR2X2_2623 ( .A(AES_CORE_DATAPATH__abc_16259_n6156), .B(AES_CORE_DATAPATH__abc_16259_n8232), .Y(AES_CORE_DATAPATH__abc_16259_n8233) );
  OR2X2 OR2X2_2624 ( .A(AES_CORE_DATAPATH__abc_16259_n8234), .B(AES_CORE_DATAPATH__abc_16259_n8228), .Y(AES_CORE_DATAPATH__0col_3__31_0__1_) );
  OR2X2 OR2X2_2625 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf9), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_34_), .Y(AES_CORE_DATAPATH__abc_16259_n8237) );
  OR2X2 OR2X2_2626 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf3), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_98_), .Y(AES_CORE_DATAPATH__abc_16259_n8238) );
  OR2X2 OR2X2_2627 ( .A(AES_CORE_DATAPATH__abc_16259_n6205), .B(AES_CORE_DATAPATH__abc_16259_n8240), .Y(AES_CORE_DATAPATH__abc_16259_n8241) );
  OR2X2 OR2X2_2628 ( .A(AES_CORE_DATAPATH__abc_16259_n8242), .B(AES_CORE_DATAPATH__abc_16259_n8236), .Y(AES_CORE_DATAPATH__0col_3__31_0__2_) );
  OR2X2 OR2X2_2629 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf8), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_35_), .Y(AES_CORE_DATAPATH__abc_16259_n8245) );
  OR2X2 OR2X2_263 ( .A(AES_CORE_DATAPATH__abc_16259_n2907), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n2908) );
  OR2X2 OR2X2_2630 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf2), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_99_), .Y(AES_CORE_DATAPATH__abc_16259_n8246) );
  OR2X2 OR2X2_2631 ( .A(AES_CORE_DATAPATH__abc_16259_n6254), .B(AES_CORE_DATAPATH__abc_16259_n8248), .Y(AES_CORE_DATAPATH__abc_16259_n8249) );
  OR2X2 OR2X2_2632 ( .A(AES_CORE_DATAPATH__abc_16259_n8250), .B(AES_CORE_DATAPATH__abc_16259_n8244), .Y(AES_CORE_DATAPATH__0col_3__31_0__3_) );
  OR2X2 OR2X2_2633 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf7), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_36_), .Y(AES_CORE_DATAPATH__abc_16259_n8253) );
  OR2X2 OR2X2_2634 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf1), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_100_), .Y(AES_CORE_DATAPATH__abc_16259_n8254) );
  OR2X2 OR2X2_2635 ( .A(AES_CORE_DATAPATH__abc_16259_n6303), .B(AES_CORE_DATAPATH__abc_16259_n8256), .Y(AES_CORE_DATAPATH__abc_16259_n8257) );
  OR2X2 OR2X2_2636 ( .A(AES_CORE_DATAPATH__abc_16259_n8258), .B(AES_CORE_DATAPATH__abc_16259_n8252), .Y(AES_CORE_DATAPATH__0col_3__31_0__4_) );
  OR2X2 OR2X2_2637 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf6), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_37_), .Y(AES_CORE_DATAPATH__abc_16259_n8261) );
  OR2X2 OR2X2_2638 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf0), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_101_), .Y(AES_CORE_DATAPATH__abc_16259_n8262) );
  OR2X2 OR2X2_2639 ( .A(AES_CORE_DATAPATH__abc_16259_n6352), .B(AES_CORE_DATAPATH__abc_16259_n8264), .Y(AES_CORE_DATAPATH__abc_16259_n8265) );
  OR2X2 OR2X2_264 ( .A(AES_CORE_DATAPATH__abc_16259_n2910), .B(AES_CORE_DATAPATH__abc_16259_n2911_1), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_1_) );
  OR2X2 OR2X2_2640 ( .A(AES_CORE_DATAPATH__abc_16259_n8266), .B(AES_CORE_DATAPATH__abc_16259_n8260), .Y(AES_CORE_DATAPATH__0col_3__31_0__5_) );
  OR2X2 OR2X2_2641 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf5), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_38_), .Y(AES_CORE_DATAPATH__abc_16259_n8269) );
  OR2X2 OR2X2_2642 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf14), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_102_), .Y(AES_CORE_DATAPATH__abc_16259_n8270) );
  OR2X2 OR2X2_2643 ( .A(AES_CORE_DATAPATH__abc_16259_n6401), .B(AES_CORE_DATAPATH__abc_16259_n8272), .Y(AES_CORE_DATAPATH__abc_16259_n8273) );
  OR2X2 OR2X2_2644 ( .A(AES_CORE_DATAPATH__abc_16259_n8274), .B(AES_CORE_DATAPATH__abc_16259_n8268), .Y(AES_CORE_DATAPATH__0col_3__31_0__6_) );
  OR2X2 OR2X2_2645 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf4), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_39_), .Y(AES_CORE_DATAPATH__abc_16259_n8277) );
  OR2X2 OR2X2_2646 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf13), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_103_), .Y(AES_CORE_DATAPATH__abc_16259_n8278) );
  OR2X2 OR2X2_2647 ( .A(AES_CORE_DATAPATH__abc_16259_n6450), .B(AES_CORE_DATAPATH__abc_16259_n8280), .Y(AES_CORE_DATAPATH__abc_16259_n8281) );
  OR2X2 OR2X2_2648 ( .A(AES_CORE_DATAPATH__abc_16259_n8282), .B(AES_CORE_DATAPATH__abc_16259_n8276), .Y(AES_CORE_DATAPATH__0col_3__31_0__7_) );
  OR2X2 OR2X2_2649 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf3), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_72_), .Y(AES_CORE_DATAPATH__abc_16259_n8285) );
  OR2X2 OR2X2_265 ( .A(AES_CORE_DATAPATH__abc_16259_n2774_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n2913), .Y(AES_CORE_DATAPATH__abc_16259_n2914) );
  OR2X2 OR2X2_2650 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf12), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_72_), .Y(AES_CORE_DATAPATH__abc_16259_n8286) );
  OR2X2 OR2X2_2651 ( .A(AES_CORE_DATAPATH__abc_16259_n6499), .B(AES_CORE_DATAPATH__abc_16259_n8288), .Y(AES_CORE_DATAPATH__abc_16259_n8289) );
  OR2X2 OR2X2_2652 ( .A(AES_CORE_DATAPATH__abc_16259_n8290), .B(AES_CORE_DATAPATH__abc_16259_n8284), .Y(AES_CORE_DATAPATH__0col_3__31_0__8_) );
  OR2X2 OR2X2_2653 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf2), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_73_), .Y(AES_CORE_DATAPATH__abc_16259_n8293) );
  OR2X2 OR2X2_2654 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf11), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_73_), .Y(AES_CORE_DATAPATH__abc_16259_n8294) );
  OR2X2 OR2X2_2655 ( .A(AES_CORE_DATAPATH__abc_16259_n6548), .B(AES_CORE_DATAPATH__abc_16259_n8296), .Y(AES_CORE_DATAPATH__abc_16259_n8297) );
  OR2X2 OR2X2_2656 ( .A(AES_CORE_DATAPATH__abc_16259_n8298), .B(AES_CORE_DATAPATH__abc_16259_n8292), .Y(AES_CORE_DATAPATH__0col_3__31_0__9_) );
  OR2X2 OR2X2_2657 ( .A(AES_CORE_DATAPATH__abc_16259_n8300), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf10), .Y(AES_CORE_DATAPATH__abc_16259_n8301) );
  OR2X2 OR2X2_2658 ( .A(AES_CORE_DATAPATH__abc_16259_n6603_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n8304), .Y(AES_CORE_DATAPATH__abc_16259_n8305) );
  OR2X2 OR2X2_2659 ( .A(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf4), .B(AES_CORE_DATAPATH_col_3__10_), .Y(AES_CORE_DATAPATH__abc_16259_n8309) );
  OR2X2 OR2X2_266 ( .A(AES_CORE_DATAPATH__abc_16259_n2778_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n2915), .Y(AES_CORE_DATAPATH__abc_16259_n2916_1) );
  OR2X2 OR2X2_2660 ( .A(AES_CORE_DATAPATH__abc_16259_n8311), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf8), .Y(AES_CORE_DATAPATH__abc_16259_n8312) );
  OR2X2 OR2X2_2661 ( .A(AES_CORE_DATAPATH__abc_16259_n6603_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n8315), .Y(AES_CORE_DATAPATH__abc_16259_n8316) );
  OR2X2 OR2X2_2662 ( .A(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf2), .B(AES_CORE_DATAPATH_col_3__11_), .Y(AES_CORE_DATAPATH__abc_16259_n8320) );
  OR2X2 OR2X2_2663 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf1), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_76_), .Y(AES_CORE_DATAPATH__abc_16259_n8323) );
  OR2X2 OR2X2_2664 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf6), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_76_), .Y(AES_CORE_DATAPATH__abc_16259_n8324) );
  OR2X2 OR2X2_2665 ( .A(AES_CORE_DATAPATH__abc_16259_n6710), .B(AES_CORE_DATAPATH__abc_16259_n8326), .Y(AES_CORE_DATAPATH__abc_16259_n8327) );
  OR2X2 OR2X2_2666 ( .A(AES_CORE_DATAPATH__abc_16259_n8328), .B(AES_CORE_DATAPATH__abc_16259_n8322), .Y(AES_CORE_DATAPATH__0col_3__31_0__12_) );
  OR2X2 OR2X2_2667 ( .A(AES_CORE_DATAPATH__abc_16259_n8330), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n8331) );
  OR2X2 OR2X2_2668 ( .A(AES_CORE_DATAPATH__abc_16259_n6603_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n8334), .Y(AES_CORE_DATAPATH__abc_16259_n8335) );
  OR2X2 OR2X2_2669 ( .A(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf5), .B(AES_CORE_DATAPATH_col_3__13_), .Y(AES_CORE_DATAPATH__abc_16259_n8339) );
  OR2X2 OR2X2_267 ( .A(AES_CORE_DATAPATH__abc_16259_n2919), .B(AES_CORE_DATAPATH__abc_16259_n2920_1), .Y(AES_CORE_DATAPATH__abc_16259_n2921) );
  OR2X2 OR2X2_2670 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf0), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_78_), .Y(AES_CORE_DATAPATH__abc_16259_n8342) );
  OR2X2 OR2X2_2671 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf3), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_78_), .Y(AES_CORE_DATAPATH__abc_16259_n8343) );
  OR2X2 OR2X2_2672 ( .A(AES_CORE_DATAPATH__abc_16259_n6813), .B(AES_CORE_DATAPATH__abc_16259_n8345), .Y(AES_CORE_DATAPATH__abc_16259_n8346) );
  OR2X2 OR2X2_2673 ( .A(AES_CORE_DATAPATH__abc_16259_n8347), .B(AES_CORE_DATAPATH__abc_16259_n8341), .Y(AES_CORE_DATAPATH__0col_3__31_0__14_) );
  OR2X2 OR2X2_2674 ( .A(AES_CORE_DATAPATH__abc_16259_n8349), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n8350) );
  OR2X2 OR2X2_2675 ( .A(AES_CORE_DATAPATH__abc_16259_n6603_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n8353), .Y(AES_CORE_DATAPATH__abc_16259_n8354) );
  OR2X2 OR2X2_2676 ( .A(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf2), .B(AES_CORE_DATAPATH_col_3__15_), .Y(AES_CORE_DATAPATH__abc_16259_n8358) );
  OR2X2 OR2X2_2677 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf12), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_112_), .Y(AES_CORE_DATAPATH__abc_16259_n8361) );
  OR2X2 OR2X2_2678 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf0), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_48_), .Y(AES_CORE_DATAPATH__abc_16259_n8362) );
  OR2X2 OR2X2_2679 ( .A(AES_CORE_DATAPATH__abc_16259_n6916), .B(AES_CORE_DATAPATH__abc_16259_n8364), .Y(AES_CORE_DATAPATH__abc_16259_n8365) );
  OR2X2 OR2X2_268 ( .A(AES_CORE_DATAPATH__abc_16259_n2921), .B(AES_CORE_DATAPATH__abc_16259_n2918), .Y(AES_CORE_DATAPATH__abc_16259_n2922_1) );
  OR2X2 OR2X2_2680 ( .A(AES_CORE_DATAPATH__abc_16259_n8366), .B(AES_CORE_DATAPATH__abc_16259_n8360), .Y(AES_CORE_DATAPATH__0col_3__31_0__16_) );
  OR2X2 OR2X2_2681 ( .A(AES_CORE_DATAPATH__abc_16259_n8368), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf14), .Y(AES_CORE_DATAPATH__abc_16259_n8369) );
  OR2X2 OR2X2_2682 ( .A(AES_CORE_DATAPATH__abc_16259_n6603_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n8372), .Y(AES_CORE_DATAPATH__abc_16259_n8373) );
  OR2X2 OR2X2_2683 ( .A(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf5), .B(AES_CORE_DATAPATH_col_3__17_), .Y(AES_CORE_DATAPATH__abc_16259_n8377) );
  OR2X2 OR2X2_2684 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf11), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_114_), .Y(AES_CORE_DATAPATH__abc_16259_n8380) );
  OR2X2 OR2X2_2685 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf12), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_50_), .Y(AES_CORE_DATAPATH__abc_16259_n8381) );
  OR2X2 OR2X2_2686 ( .A(AES_CORE_DATAPATH__abc_16259_n7019), .B(AES_CORE_DATAPATH__abc_16259_n8383), .Y(AES_CORE_DATAPATH__abc_16259_n8384) );
  OR2X2 OR2X2_2687 ( .A(AES_CORE_DATAPATH__abc_16259_n8385), .B(AES_CORE_DATAPATH__abc_16259_n8379), .Y(AES_CORE_DATAPATH__0col_3__31_0__18_) );
  OR2X2 OR2X2_2688 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf10), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_115_), .Y(AES_CORE_DATAPATH__abc_16259_n8388) );
  OR2X2 OR2X2_2689 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf11), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_51_), .Y(AES_CORE_DATAPATH__abc_16259_n8389) );
  OR2X2 OR2X2_269 ( .A(AES_CORE_DATAPATH__abc_16259_n2926_1), .B(AES_CORE_DATAPATH__abc_16259_n2826_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n2927) );
  OR2X2 OR2X2_2690 ( .A(AES_CORE_DATAPATH__abc_16259_n7068), .B(AES_CORE_DATAPATH__abc_16259_n8391), .Y(AES_CORE_DATAPATH__abc_16259_n8392) );
  OR2X2 OR2X2_2691 ( .A(AES_CORE_DATAPATH__abc_16259_n8393), .B(AES_CORE_DATAPATH__abc_16259_n8387), .Y(AES_CORE_DATAPATH__0col_3__31_0__19_) );
  OR2X2 OR2X2_2692 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf9), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_116_), .Y(AES_CORE_DATAPATH__abc_16259_n8396) );
  OR2X2 OR2X2_2693 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf10), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_52_), .Y(AES_CORE_DATAPATH__abc_16259_n8397) );
  OR2X2 OR2X2_2694 ( .A(AES_CORE_DATAPATH__abc_16259_n7117), .B(AES_CORE_DATAPATH__abc_16259_n8399), .Y(AES_CORE_DATAPATH__abc_16259_n8400) );
  OR2X2 OR2X2_2695 ( .A(AES_CORE_DATAPATH__abc_16259_n8401), .B(AES_CORE_DATAPATH__abc_16259_n8395), .Y(AES_CORE_DATAPATH__0col_3__31_0__20_) );
  OR2X2 OR2X2_2696 ( .A(AES_CORE_DATAPATH__abc_16259_n8403), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf9), .Y(AES_CORE_DATAPATH__abc_16259_n8404) );
  OR2X2 OR2X2_2697 ( .A(AES_CORE_DATAPATH__abc_16259_n6603_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n8407), .Y(AES_CORE_DATAPATH__abc_16259_n8408) );
  OR2X2 OR2X2_2698 ( .A(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf0), .B(AES_CORE_DATAPATH_col_3__21_), .Y(AES_CORE_DATAPATH__abc_16259_n8412) );
  OR2X2 OR2X2_2699 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf8), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_118_), .Y(AES_CORE_DATAPATH__abc_16259_n8415) );
  OR2X2 OR2X2_27 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk_bF_buf3), .B(AES_CORE_CONTROL_UNIT__abc_15841_n76_1), .Y(AES_CORE_CONTROL_UNIT_bypass_key_en) );
  OR2X2 OR2X2_270 ( .A(AES_CORE_DATAPATH__abc_16259_n2928), .B(AES_CORE_DATAPATH__abc_16259_n2929), .Y(AES_CORE_DATAPATH__abc_16259_n2930) );
  OR2X2 OR2X2_2700 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf7), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_54_), .Y(AES_CORE_DATAPATH__abc_16259_n8416) );
  OR2X2 OR2X2_2701 ( .A(AES_CORE_DATAPATH__abc_16259_n7220), .B(AES_CORE_DATAPATH__abc_16259_n8418), .Y(AES_CORE_DATAPATH__abc_16259_n8419) );
  OR2X2 OR2X2_2702 ( .A(AES_CORE_DATAPATH__abc_16259_n8420), .B(AES_CORE_DATAPATH__abc_16259_n8414), .Y(AES_CORE_DATAPATH__0col_3__31_0__22_) );
  OR2X2 OR2X2_2703 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf7), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_119_), .Y(AES_CORE_DATAPATH__abc_16259_n8423) );
  OR2X2 OR2X2_2704 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf6), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_55_), .Y(AES_CORE_DATAPATH__abc_16259_n8424) );
  OR2X2 OR2X2_2705 ( .A(AES_CORE_DATAPATH__abc_16259_n7269), .B(AES_CORE_DATAPATH__abc_16259_n8426), .Y(AES_CORE_DATAPATH__abc_16259_n8427) );
  OR2X2 OR2X2_2706 ( .A(AES_CORE_DATAPATH__abc_16259_n8428), .B(AES_CORE_DATAPATH__abc_16259_n8422), .Y(AES_CORE_DATAPATH__0col_3__31_0__23_) );
  OR2X2 OR2X2_2707 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf6), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_24_), .Y(AES_CORE_DATAPATH__abc_16259_n8431) );
  OR2X2 OR2X2_2708 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf5), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_24_), .Y(AES_CORE_DATAPATH__abc_16259_n8432) );
  OR2X2 OR2X2_2709 ( .A(AES_CORE_DATAPATH__abc_16259_n7318), .B(AES_CORE_DATAPATH__abc_16259_n8434), .Y(AES_CORE_DATAPATH__abc_16259_n8435) );
  OR2X2 OR2X2_271 ( .A(AES_CORE_DATAPATH__abc_16259_n2930), .B(AES_CORE_DATAPATH__abc_16259_n2927), .Y(AES_CORE_DATAPATH__abc_16259_n2931) );
  OR2X2 OR2X2_2710 ( .A(AES_CORE_DATAPATH__abc_16259_n8436), .B(AES_CORE_DATAPATH__abc_16259_n8430), .Y(AES_CORE_DATAPATH__0col_3__31_0__24_) );
  OR2X2 OR2X2_2711 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf5), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_25_), .Y(AES_CORE_DATAPATH__abc_16259_n8439) );
  OR2X2 OR2X2_2712 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf4), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_25_), .Y(AES_CORE_DATAPATH__abc_16259_n8440) );
  OR2X2 OR2X2_2713 ( .A(AES_CORE_DATAPATH__abc_16259_n7367), .B(AES_CORE_DATAPATH__abc_16259_n8442), .Y(AES_CORE_DATAPATH__abc_16259_n8443) );
  OR2X2 OR2X2_2714 ( .A(AES_CORE_DATAPATH__abc_16259_n8444), .B(AES_CORE_DATAPATH__abc_16259_n8438), .Y(AES_CORE_DATAPATH__0col_3__31_0__25_) );
  OR2X2 OR2X2_2715 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf4), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_26_), .Y(AES_CORE_DATAPATH__abc_16259_n8447) );
  OR2X2 OR2X2_2716 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf3), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_26_), .Y(AES_CORE_DATAPATH__abc_16259_n8448) );
  OR2X2 OR2X2_2717 ( .A(AES_CORE_DATAPATH__abc_16259_n7416), .B(AES_CORE_DATAPATH__abc_16259_n8450), .Y(AES_CORE_DATAPATH__abc_16259_n8451) );
  OR2X2 OR2X2_2718 ( .A(AES_CORE_DATAPATH__abc_16259_n8452), .B(AES_CORE_DATAPATH__abc_16259_n8446), .Y(AES_CORE_DATAPATH__0col_3__31_0__26_) );
  OR2X2 OR2X2_2719 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf3), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_27_), .Y(AES_CORE_DATAPATH__abc_16259_n8455) );
  OR2X2 OR2X2_272 ( .A(AES_CORE_DATAPATH__abc_16259_n2841_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__2_), .Y(AES_CORE_DATAPATH__abc_16259_n2932) );
  OR2X2 OR2X2_2720 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf2), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_27_), .Y(AES_CORE_DATAPATH__abc_16259_n8456) );
  OR2X2 OR2X2_2721 ( .A(AES_CORE_DATAPATH__abc_16259_n7465), .B(AES_CORE_DATAPATH__abc_16259_n8458), .Y(AES_CORE_DATAPATH__abc_16259_n8459) );
  OR2X2 OR2X2_2722 ( .A(AES_CORE_DATAPATH__abc_16259_n8460), .B(AES_CORE_DATAPATH__abc_16259_n8454), .Y(AES_CORE_DATAPATH__0col_3__31_0__27_) );
  OR2X2 OR2X2_2723 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf2), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_28_), .Y(AES_CORE_DATAPATH__abc_16259_n8463) );
  OR2X2 OR2X2_2724 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf1), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_28_), .Y(AES_CORE_DATAPATH__abc_16259_n8464) );
  OR2X2 OR2X2_2725 ( .A(AES_CORE_DATAPATH__abc_16259_n7514), .B(AES_CORE_DATAPATH__abc_16259_n8466), .Y(AES_CORE_DATAPATH__abc_16259_n8467) );
  OR2X2 OR2X2_2726 ( .A(AES_CORE_DATAPATH__abc_16259_n8468), .B(AES_CORE_DATAPATH__abc_16259_n8462), .Y(AES_CORE_DATAPATH__0col_3__31_0__28_) );
  OR2X2 OR2X2_2727 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf1), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_29_), .Y(AES_CORE_DATAPATH__abc_16259_n8471) );
  OR2X2 OR2X2_2728 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf0), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_29_), .Y(AES_CORE_DATAPATH__abc_16259_n8472) );
  OR2X2 OR2X2_2729 ( .A(AES_CORE_DATAPATH__abc_16259_n7563), .B(AES_CORE_DATAPATH__abc_16259_n8474), .Y(AES_CORE_DATAPATH__abc_16259_n8475) );
  OR2X2 OR2X2_273 ( .A(AES_CORE_DATAPATH__abc_16259_n2924_1), .B(AES_CORE_DATAPATH__abc_16259_n2853_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n2934) );
  OR2X2 OR2X2_2730 ( .A(AES_CORE_DATAPATH__abc_16259_n8476), .B(AES_CORE_DATAPATH__abc_16259_n8470), .Y(AES_CORE_DATAPATH__0col_3__31_0__29_) );
  OR2X2 OR2X2_2731 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf0), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_30_), .Y(AES_CORE_DATAPATH__abc_16259_n8479) );
  OR2X2 OR2X2_2732 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf14), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_30_), .Y(AES_CORE_DATAPATH__abc_16259_n8480) );
  OR2X2 OR2X2_2733 ( .A(AES_CORE_DATAPATH__abc_16259_n7612), .B(AES_CORE_DATAPATH__abc_16259_n8482), .Y(AES_CORE_DATAPATH__abc_16259_n8483) );
  OR2X2 OR2X2_2734 ( .A(AES_CORE_DATAPATH__abc_16259_n8484), .B(AES_CORE_DATAPATH__abc_16259_n8478), .Y(AES_CORE_DATAPATH__0col_3__31_0__30_) );
  OR2X2 OR2X2_2735 ( .A(AES_CORE_DATAPATH__abc_16259_n2802_bF_buf12), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_31_), .Y(AES_CORE_DATAPATH__abc_16259_n8487) );
  OR2X2 OR2X2_2736 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf13), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_31_), .Y(AES_CORE_DATAPATH__abc_16259_n8488) );
  OR2X2 OR2X2_2737 ( .A(AES_CORE_DATAPATH__abc_16259_n7661), .B(AES_CORE_DATAPATH__abc_16259_n8490), .Y(AES_CORE_DATAPATH__abc_16259_n8491) );
  OR2X2 OR2X2_2738 ( .A(AES_CORE_DATAPATH__abc_16259_n8492), .B(AES_CORE_DATAPATH__abc_16259_n8486), .Y(AES_CORE_DATAPATH__0col_3__31_0__31_) );
  OR2X2 OR2X2_2739 ( .A(AES_CORE_DATAPATH__abc_16259_n8495), .B(AES_CORE_DATAPATH__abc_16259_n8498), .Y(AES_CORE_DATAPATH__abc_16259_n8499) );
  OR2X2 OR2X2_274 ( .A(AES_CORE_DATAPATH__abc_16259_n2935), .B(AES_CORE_DATAPATH__abc_16259_n2936), .Y(AES_CORE_DATAPATH__abc_16259_n2937) );
  OR2X2 OR2X2_2740 ( .A(AES_CORE_DATAPATH__abc_16259_n8502), .B(AES_CORE_DATAPATH__abc_16259_n8501), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__0_) );
  OR2X2 OR2X2_2741 ( .A(AES_CORE_DATAPATH__abc_16259_n8505), .B(AES_CORE_DATAPATH__abc_16259_n8504), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__1_) );
  OR2X2 OR2X2_2742 ( .A(AES_CORE_DATAPATH__abc_16259_n8508), .B(AES_CORE_DATAPATH__abc_16259_n8507), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__2_) );
  OR2X2 OR2X2_2743 ( .A(AES_CORE_DATAPATH__abc_16259_n8511), .B(AES_CORE_DATAPATH__abc_16259_n8510), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__3_) );
  OR2X2 OR2X2_2744 ( .A(AES_CORE_DATAPATH__abc_16259_n8514), .B(AES_CORE_DATAPATH__abc_16259_n8513), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__4_) );
  OR2X2 OR2X2_2745 ( .A(AES_CORE_DATAPATH__abc_16259_n8517), .B(AES_CORE_DATAPATH__abc_16259_n8516), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__5_) );
  OR2X2 OR2X2_2746 ( .A(AES_CORE_DATAPATH__abc_16259_n8520), .B(AES_CORE_DATAPATH__abc_16259_n8519), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__6_) );
  OR2X2 OR2X2_2747 ( .A(AES_CORE_DATAPATH__abc_16259_n8523), .B(AES_CORE_DATAPATH__abc_16259_n8522), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__7_) );
  OR2X2 OR2X2_2748 ( .A(AES_CORE_DATAPATH__abc_16259_n8526), .B(AES_CORE_DATAPATH__abc_16259_n8525), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__8_) );
  OR2X2 OR2X2_2749 ( .A(AES_CORE_DATAPATH__abc_16259_n8529), .B(AES_CORE_DATAPATH__abc_16259_n8528), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__9_) );
  OR2X2 OR2X2_275 ( .A(_auto_iopadmap_cc_313_execute_26949_2_), .B(AES_CORE_DATAPATH__abc_16259_n2939), .Y(AES_CORE_DATAPATH__abc_16259_n2940_1) );
  OR2X2 OR2X2_2750 ( .A(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1_3__10_), .Y(AES_CORE_DATAPATH__abc_16259_n8533) );
  OR2X2 OR2X2_2751 ( .A(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf1), .B(AES_CORE_DATAPATH_bkp_1_3__11_), .Y(AES_CORE_DATAPATH__abc_16259_n8537) );
  OR2X2 OR2X2_2752 ( .A(AES_CORE_DATAPATH__abc_16259_n8540), .B(AES_CORE_DATAPATH__abc_16259_n8539), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__12_) );
  OR2X2 OR2X2_2753 ( .A(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf6), .B(AES_CORE_DATAPATH_bkp_1_3__13_), .Y(AES_CORE_DATAPATH__abc_16259_n8544) );
  OR2X2 OR2X2_2754 ( .A(AES_CORE_DATAPATH__abc_16259_n8547), .B(AES_CORE_DATAPATH__abc_16259_n8546), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__14_) );
  OR2X2 OR2X2_2755 ( .A(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1_3__15_), .Y(AES_CORE_DATAPATH__abc_16259_n8551) );
  OR2X2 OR2X2_2756 ( .A(AES_CORE_DATAPATH__abc_16259_n8554), .B(AES_CORE_DATAPATH__abc_16259_n8553), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__16_) );
  OR2X2 OR2X2_2757 ( .A(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf0), .B(AES_CORE_DATAPATH_bkp_1_3__17_), .Y(AES_CORE_DATAPATH__abc_16259_n8558) );
  OR2X2 OR2X2_2758 ( .A(AES_CORE_DATAPATH__abc_16259_n8561), .B(AES_CORE_DATAPATH__abc_16259_n8560), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__18_) );
  OR2X2 OR2X2_2759 ( .A(AES_CORE_DATAPATH__abc_16259_n8564), .B(AES_CORE_DATAPATH__abc_16259_n8563), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__19_) );
  OR2X2 OR2X2_276 ( .A(AES_CORE_DATAPATH__abc_16259_n2942), .B(AES_CORE_DATAPATH__abc_16259_n2864_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n2943) );
  OR2X2 OR2X2_2760 ( .A(AES_CORE_DATAPATH__abc_16259_n8567), .B(AES_CORE_DATAPATH__abc_16259_n8566), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__20_) );
  OR2X2 OR2X2_2761 ( .A(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1_3__21_), .Y(AES_CORE_DATAPATH__abc_16259_n8571) );
  OR2X2 OR2X2_2762 ( .A(AES_CORE_DATAPATH__abc_16259_n8574), .B(AES_CORE_DATAPATH__abc_16259_n8573), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__22_) );
  OR2X2 OR2X2_2763 ( .A(AES_CORE_DATAPATH__abc_16259_n8577), .B(AES_CORE_DATAPATH__abc_16259_n8576), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__23_) );
  OR2X2 OR2X2_2764 ( .A(AES_CORE_DATAPATH__abc_16259_n8580), .B(AES_CORE_DATAPATH__abc_16259_n8579), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__24_) );
  OR2X2 OR2X2_2765 ( .A(AES_CORE_DATAPATH__abc_16259_n8583), .B(AES_CORE_DATAPATH__abc_16259_n8582), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__25_) );
  OR2X2 OR2X2_2766 ( .A(AES_CORE_DATAPATH__abc_16259_n8586), .B(AES_CORE_DATAPATH__abc_16259_n8585), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__26_) );
  OR2X2 OR2X2_2767 ( .A(AES_CORE_DATAPATH__abc_16259_n8589), .B(AES_CORE_DATAPATH__abc_16259_n8588), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__27_) );
  OR2X2 OR2X2_2768 ( .A(AES_CORE_DATAPATH__abc_16259_n8592), .B(AES_CORE_DATAPATH__abc_16259_n8591), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__28_) );
  OR2X2 OR2X2_2769 ( .A(AES_CORE_DATAPATH__abc_16259_n8595), .B(AES_CORE_DATAPATH__abc_16259_n8594), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__29_) );
  OR2X2 OR2X2_277 ( .A(AES_CORE_DATAPATH__abc_16259_n2943), .B(AES_CORE_DATAPATH__abc_16259_n2941), .Y(AES_CORE_DATAPATH__abc_16259_n2944) );
  OR2X2 OR2X2_2770 ( .A(AES_CORE_DATAPATH__abc_16259_n8598), .B(AES_CORE_DATAPATH__abc_16259_n8597), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__30_) );
  OR2X2 OR2X2_2771 ( .A(AES_CORE_DATAPATH__abc_16259_n8601), .B(AES_CORE_DATAPATH__abc_16259_n8600), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__31_) );
  OR2X2 OR2X2_2772 ( .A(AES_CORE_DATAPATH__abc_16259_n6112), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf9), .Y(AES_CORE_DATAPATH__abc_16259_n8604) );
  OR2X2 OR2X2_2773 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf9), .B(AES_CORE_DATAPATH_bkp_1_3__0_), .Y(AES_CORE_DATAPATH__abc_16259_n8605) );
  OR2X2 OR2X2_2774 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n8608), .Y(AES_CORE_DATAPATH__abc_16259_n8609) );
  OR2X2 OR2X2_2775 ( .A(AES_CORE_DATAPATH__abc_16259_n8607), .B(AES_CORE_DATAPATH__abc_16259_n8609), .Y(AES_CORE_DATAPATH__abc_16259_n8610) );
  OR2X2 OR2X2_2776 ( .A(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf0), .B(AES_CORE_DATAPATH_bkp_3__0_), .Y(AES_CORE_DATAPATH__abc_16259_n8611) );
  OR2X2 OR2X2_2777 ( .A(AES_CORE_DATAPATH__abc_16259_n6161), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf8), .Y(AES_CORE_DATAPATH__abc_16259_n8613) );
  OR2X2 OR2X2_2778 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf8), .B(AES_CORE_DATAPATH_bkp_1_3__1_), .Y(AES_CORE_DATAPATH__abc_16259_n8614) );
  OR2X2 OR2X2_2779 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n8617), .Y(AES_CORE_DATAPATH__abc_16259_n8618) );
  OR2X2 OR2X2_278 ( .A(AES_CORE_DATAPATH__abc_16259_n2946_1), .B(AES_CORE_DATAPATH__abc_16259_n2945_1), .Y(AES_CORE_DATAPATH__abc_16259_n2947) );
  OR2X2 OR2X2_2780 ( .A(AES_CORE_DATAPATH__abc_16259_n8616), .B(AES_CORE_DATAPATH__abc_16259_n8618), .Y(AES_CORE_DATAPATH__abc_16259_n8619) );
  OR2X2 OR2X2_2781 ( .A(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf7), .B(AES_CORE_DATAPATH_bkp_3__1_), .Y(AES_CORE_DATAPATH__abc_16259_n8620) );
  OR2X2 OR2X2_2782 ( .A(AES_CORE_DATAPATH__abc_16259_n6210), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n8622) );
  OR2X2 OR2X2_2783 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf7), .B(AES_CORE_DATAPATH_bkp_1_3__2_), .Y(AES_CORE_DATAPATH__abc_16259_n8623) );
  OR2X2 OR2X2_2784 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf6), .B(AES_CORE_DATAPATH__abc_16259_n8626), .Y(AES_CORE_DATAPATH__abc_16259_n8627) );
  OR2X2 OR2X2_2785 ( .A(AES_CORE_DATAPATH__abc_16259_n8625), .B(AES_CORE_DATAPATH__abc_16259_n8627), .Y(AES_CORE_DATAPATH__abc_16259_n8628) );
  OR2X2 OR2X2_2786 ( .A(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf6), .B(AES_CORE_DATAPATH_bkp_3__2_), .Y(AES_CORE_DATAPATH__abc_16259_n8629) );
  OR2X2 OR2X2_2787 ( .A(AES_CORE_DATAPATH__abc_16259_n6259), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n8631) );
  OR2X2 OR2X2_2788 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf6), .B(AES_CORE_DATAPATH_bkp_1_3__3_), .Y(AES_CORE_DATAPATH__abc_16259_n8632) );
  OR2X2 OR2X2_2789 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf5), .B(AES_CORE_DATAPATH__abc_16259_n8635), .Y(AES_CORE_DATAPATH__abc_16259_n8636) );
  OR2X2 OR2X2_279 ( .A(AES_CORE_DATAPATH__abc_16259_n2947), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n2948) );
  OR2X2 OR2X2_2790 ( .A(AES_CORE_DATAPATH__abc_16259_n8634), .B(AES_CORE_DATAPATH__abc_16259_n8636), .Y(AES_CORE_DATAPATH__abc_16259_n8637) );
  OR2X2 OR2X2_2791 ( .A(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf5), .B(AES_CORE_DATAPATH_bkp_3__3_), .Y(AES_CORE_DATAPATH__abc_16259_n8638) );
  OR2X2 OR2X2_2792 ( .A(AES_CORE_DATAPATH__abc_16259_n6308), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n8640) );
  OR2X2 OR2X2_2793 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf5), .B(AES_CORE_DATAPATH_bkp_1_3__4_), .Y(AES_CORE_DATAPATH__abc_16259_n8641) );
  OR2X2 OR2X2_2794 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n8644), .Y(AES_CORE_DATAPATH__abc_16259_n8645) );
  OR2X2 OR2X2_2795 ( .A(AES_CORE_DATAPATH__abc_16259_n8643), .B(AES_CORE_DATAPATH__abc_16259_n8645), .Y(AES_CORE_DATAPATH__abc_16259_n8646) );
  OR2X2 OR2X2_2796 ( .A(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf4), .B(AES_CORE_DATAPATH_bkp_3__4_), .Y(AES_CORE_DATAPATH__abc_16259_n8647) );
  OR2X2 OR2X2_2797 ( .A(AES_CORE_DATAPATH__abc_16259_n6357), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n8649) );
  OR2X2 OR2X2_2798 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf4), .B(AES_CORE_DATAPATH_bkp_1_3__5_), .Y(AES_CORE_DATAPATH__abc_16259_n8650) );
  OR2X2 OR2X2_2799 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n8653), .Y(AES_CORE_DATAPATH__abc_16259_n8654) );
  OR2X2 OR2X2_28 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n148), .B(AES_CORE_CONTROL_UNIT__abc_15841_n149), .Y(AES_CORE_CONTROL_UNIT__abc_10818_n109) );
  OR2X2 OR2X2_280 ( .A(AES_CORE_DATAPATH__abc_16259_n2950), .B(AES_CORE_DATAPATH__abc_16259_n2951_1), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_2_) );
  OR2X2 OR2X2_2800 ( .A(AES_CORE_DATAPATH__abc_16259_n8652), .B(AES_CORE_DATAPATH__abc_16259_n8654), .Y(AES_CORE_DATAPATH__abc_16259_n8655) );
  OR2X2 OR2X2_2801 ( .A(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf3), .B(AES_CORE_DATAPATH_bkp_3__5_), .Y(AES_CORE_DATAPATH__abc_16259_n8656) );
  OR2X2 OR2X2_2802 ( .A(AES_CORE_DATAPATH__abc_16259_n6406), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n8658) );
  OR2X2 OR2X2_2803 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1_3__6_), .Y(AES_CORE_DATAPATH__abc_16259_n8659) );
  OR2X2 OR2X2_2804 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n8662), .Y(AES_CORE_DATAPATH__abc_16259_n8663) );
  OR2X2 OR2X2_2805 ( .A(AES_CORE_DATAPATH__abc_16259_n8661), .B(AES_CORE_DATAPATH__abc_16259_n8663), .Y(AES_CORE_DATAPATH__abc_16259_n8664) );
  OR2X2 OR2X2_2806 ( .A(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf2), .B(AES_CORE_DATAPATH_bkp_3__6_), .Y(AES_CORE_DATAPATH__abc_16259_n8665) );
  OR2X2 OR2X2_2807 ( .A(AES_CORE_DATAPATH__abc_16259_n6455), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n8667) );
  OR2X2 OR2X2_2808 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf2), .B(AES_CORE_DATAPATH_bkp_1_3__7_), .Y(AES_CORE_DATAPATH__abc_16259_n8668) );
  OR2X2 OR2X2_2809 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n8671), .Y(AES_CORE_DATAPATH__abc_16259_n8672) );
  OR2X2 OR2X2_281 ( .A(AES_CORE_DATAPATH__abc_16259_n2774_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n2953_1), .Y(AES_CORE_DATAPATH__abc_16259_n2954) );
  OR2X2 OR2X2_2810 ( .A(AES_CORE_DATAPATH__abc_16259_n8670), .B(AES_CORE_DATAPATH__abc_16259_n8672), .Y(AES_CORE_DATAPATH__abc_16259_n8673) );
  OR2X2 OR2X2_2811 ( .A(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf1), .B(AES_CORE_DATAPATH_bkp_3__7_), .Y(AES_CORE_DATAPATH__abc_16259_n8674) );
  OR2X2 OR2X2_2812 ( .A(AES_CORE_DATAPATH__abc_16259_n6504), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n8676) );
  OR2X2 OR2X2_2813 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf1), .B(AES_CORE_DATAPATH_bkp_1_3__8_), .Y(AES_CORE_DATAPATH__abc_16259_n8677) );
  OR2X2 OR2X2_2814 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n8680), .Y(AES_CORE_DATAPATH__abc_16259_n8681) );
  OR2X2 OR2X2_2815 ( .A(AES_CORE_DATAPATH__abc_16259_n8679), .B(AES_CORE_DATAPATH__abc_16259_n8681), .Y(AES_CORE_DATAPATH__abc_16259_n8682) );
  OR2X2 OR2X2_2816 ( .A(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf0), .B(AES_CORE_DATAPATH_bkp_3__8_), .Y(AES_CORE_DATAPATH__abc_16259_n8683) );
  OR2X2 OR2X2_2817 ( .A(AES_CORE_DATAPATH__abc_16259_n6553), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n8685) );
  OR2X2 OR2X2_2818 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf0), .B(AES_CORE_DATAPATH_bkp_1_3__9_), .Y(AES_CORE_DATAPATH__abc_16259_n8686) );
  OR2X2 OR2X2_2819 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf6), .B(AES_CORE_DATAPATH__abc_16259_n8689), .Y(AES_CORE_DATAPATH__abc_16259_n8690) );
  OR2X2 OR2X2_282 ( .A(AES_CORE_DATAPATH__abc_16259_n2778_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n2955_1), .Y(AES_CORE_DATAPATH__abc_16259_n2956) );
  OR2X2 OR2X2_2820 ( .A(AES_CORE_DATAPATH__abc_16259_n8688), .B(AES_CORE_DATAPATH__abc_16259_n8690), .Y(AES_CORE_DATAPATH__abc_16259_n8691) );
  OR2X2 OR2X2_2821 ( .A(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf7), .B(AES_CORE_DATAPATH_bkp_3__9_), .Y(AES_CORE_DATAPATH__abc_16259_n8692) );
  OR2X2 OR2X2_2822 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf10), .B(AES_CORE_DATAPATH_bkp_1_3__10_), .Y(AES_CORE_DATAPATH__abc_16259_n8696) );
  OR2X2 OR2X2_2823 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf5), .B(AES_CORE_DATAPATH__abc_16259_n8699), .Y(AES_CORE_DATAPATH__abc_16259_n8700) );
  OR2X2 OR2X2_2824 ( .A(AES_CORE_DATAPATH__abc_16259_n8698), .B(AES_CORE_DATAPATH__abc_16259_n8700), .Y(AES_CORE_DATAPATH__abc_16259_n8701) );
  OR2X2 OR2X2_2825 ( .A(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf6), .B(AES_CORE_DATAPATH_bkp_3__10_), .Y(AES_CORE_DATAPATH__abc_16259_n8702) );
  OR2X2 OR2X2_2826 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf8), .B(AES_CORE_DATAPATH_bkp_1_3__11_), .Y(AES_CORE_DATAPATH__abc_16259_n8706) );
  OR2X2 OR2X2_2827 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n8709), .Y(AES_CORE_DATAPATH__abc_16259_n8710) );
  OR2X2 OR2X2_2828 ( .A(AES_CORE_DATAPATH__abc_16259_n8708), .B(AES_CORE_DATAPATH__abc_16259_n8710), .Y(AES_CORE_DATAPATH__abc_16259_n8711) );
  OR2X2 OR2X2_2829 ( .A(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf5), .B(AES_CORE_DATAPATH_bkp_3__11_), .Y(AES_CORE_DATAPATH__abc_16259_n8712) );
  OR2X2 OR2X2_283 ( .A(AES_CORE_DATAPATH__abc_16259_n2959), .B(AES_CORE_DATAPATH__abc_16259_n2960), .Y(AES_CORE_DATAPATH__abc_16259_n2961) );
  OR2X2 OR2X2_2830 ( .A(AES_CORE_DATAPATH__abc_16259_n6715), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf9), .Y(AES_CORE_DATAPATH__abc_16259_n8714) );
  OR2X2 OR2X2_2831 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf7), .B(AES_CORE_DATAPATH_bkp_1_3__12_), .Y(AES_CORE_DATAPATH__abc_16259_n8715) );
  OR2X2 OR2X2_2832 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n8718), .Y(AES_CORE_DATAPATH__abc_16259_n8719) );
  OR2X2 OR2X2_2833 ( .A(AES_CORE_DATAPATH__abc_16259_n8717), .B(AES_CORE_DATAPATH__abc_16259_n8719), .Y(AES_CORE_DATAPATH__abc_16259_n8720) );
  OR2X2 OR2X2_2834 ( .A(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf4), .B(AES_CORE_DATAPATH_bkp_3__12_), .Y(AES_CORE_DATAPATH__abc_16259_n8721) );
  OR2X2 OR2X2_2835 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf5), .B(AES_CORE_DATAPATH_bkp_1_3__13_), .Y(AES_CORE_DATAPATH__abc_16259_n8725) );
  OR2X2 OR2X2_2836 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n8728), .Y(AES_CORE_DATAPATH__abc_16259_n8729) );
  OR2X2 OR2X2_2837 ( .A(AES_CORE_DATAPATH__abc_16259_n8727), .B(AES_CORE_DATAPATH__abc_16259_n8729), .Y(AES_CORE_DATAPATH__abc_16259_n8730) );
  OR2X2 OR2X2_2838 ( .A(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf3), .B(AES_CORE_DATAPATH_bkp_3__13_), .Y(AES_CORE_DATAPATH__abc_16259_n8731) );
  OR2X2 OR2X2_2839 ( .A(AES_CORE_DATAPATH__abc_16259_n6818), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf8), .Y(AES_CORE_DATAPATH__abc_16259_n8733) );
  OR2X2 OR2X2_284 ( .A(AES_CORE_DATAPATH__abc_16259_n2961), .B(AES_CORE_DATAPATH__abc_16259_n2958), .Y(AES_CORE_DATAPATH__abc_16259_n2962) );
  OR2X2 OR2X2_2840 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf4), .B(AES_CORE_DATAPATH_bkp_1_3__14_), .Y(AES_CORE_DATAPATH__abc_16259_n8734) );
  OR2X2 OR2X2_2841 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n8737), .Y(AES_CORE_DATAPATH__abc_16259_n8738) );
  OR2X2 OR2X2_2842 ( .A(AES_CORE_DATAPATH__abc_16259_n8736), .B(AES_CORE_DATAPATH__abc_16259_n8738), .Y(AES_CORE_DATAPATH__abc_16259_n8739) );
  OR2X2 OR2X2_2843 ( .A(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf2), .B(AES_CORE_DATAPATH_bkp_3__14_), .Y(AES_CORE_DATAPATH__abc_16259_n8740) );
  OR2X2 OR2X2_2844 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf2), .B(AES_CORE_DATAPATH_bkp_1_3__15_), .Y(AES_CORE_DATAPATH__abc_16259_n8744) );
  OR2X2 OR2X2_2845 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n8747), .Y(AES_CORE_DATAPATH__abc_16259_n8748) );
  OR2X2 OR2X2_2846 ( .A(AES_CORE_DATAPATH__abc_16259_n8746), .B(AES_CORE_DATAPATH__abc_16259_n8748), .Y(AES_CORE_DATAPATH__abc_16259_n8749) );
  OR2X2 OR2X2_2847 ( .A(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf1), .B(AES_CORE_DATAPATH_bkp_3__15_), .Y(AES_CORE_DATAPATH__abc_16259_n8750) );
  OR2X2 OR2X2_2848 ( .A(AES_CORE_DATAPATH__abc_16259_n6921), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n8752) );
  OR2X2 OR2X2_2849 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf1), .B(AES_CORE_DATAPATH_bkp_1_3__16_), .Y(AES_CORE_DATAPATH__abc_16259_n8753) );
  OR2X2 OR2X2_285 ( .A(AES_CORE_DATAPATH__abc_16259_n2966), .B(AES_CORE_DATAPATH__abc_16259_n2826_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n2967_1) );
  OR2X2 OR2X2_2850 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf6), .B(AES_CORE_DATAPATH__abc_16259_n8756), .Y(AES_CORE_DATAPATH__abc_16259_n8757) );
  OR2X2 OR2X2_2851 ( .A(AES_CORE_DATAPATH__abc_16259_n8755), .B(AES_CORE_DATAPATH__abc_16259_n8757), .Y(AES_CORE_DATAPATH__abc_16259_n8758) );
  OR2X2 OR2X2_2852 ( .A(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf0), .B(AES_CORE_DATAPATH_bkp_3__16_), .Y(AES_CORE_DATAPATH__abc_16259_n8759) );
  OR2X2 OR2X2_2853 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf11), .B(AES_CORE_DATAPATH_bkp_1_3__17_), .Y(AES_CORE_DATAPATH__abc_16259_n8763) );
  OR2X2 OR2X2_2854 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf5), .B(AES_CORE_DATAPATH__abc_16259_n8766), .Y(AES_CORE_DATAPATH__abc_16259_n8767) );
  OR2X2 OR2X2_2855 ( .A(AES_CORE_DATAPATH__abc_16259_n8765), .B(AES_CORE_DATAPATH__abc_16259_n8767), .Y(AES_CORE_DATAPATH__abc_16259_n8768) );
  OR2X2 OR2X2_2856 ( .A(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf7), .B(AES_CORE_DATAPATH_bkp_3__17_), .Y(AES_CORE_DATAPATH__abc_16259_n8769) );
  OR2X2 OR2X2_2857 ( .A(AES_CORE_DATAPATH__abc_16259_n7024), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n8771) );
  OR2X2 OR2X2_2858 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf10), .B(AES_CORE_DATAPATH_bkp_1_3__18_), .Y(AES_CORE_DATAPATH__abc_16259_n8772) );
  OR2X2 OR2X2_2859 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n8775), .Y(AES_CORE_DATAPATH__abc_16259_n8776) );
  OR2X2 OR2X2_286 ( .A(AES_CORE_DATAPATH__abc_16259_n2968), .B(AES_CORE_DATAPATH__abc_16259_n2969_1), .Y(AES_CORE_DATAPATH__abc_16259_n2970) );
  OR2X2 OR2X2_2860 ( .A(AES_CORE_DATAPATH__abc_16259_n8774), .B(AES_CORE_DATAPATH__abc_16259_n8776), .Y(AES_CORE_DATAPATH__abc_16259_n8777) );
  OR2X2 OR2X2_2861 ( .A(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf6), .B(AES_CORE_DATAPATH_bkp_3__18_), .Y(AES_CORE_DATAPATH__abc_16259_n8778) );
  OR2X2 OR2X2_2862 ( .A(AES_CORE_DATAPATH__abc_16259_n7073), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n8780) );
  OR2X2 OR2X2_2863 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf9), .B(AES_CORE_DATAPATH_bkp_1_3__19_), .Y(AES_CORE_DATAPATH__abc_16259_n8781) );
  OR2X2 OR2X2_2864 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n8784), .Y(AES_CORE_DATAPATH__abc_16259_n8785) );
  OR2X2 OR2X2_2865 ( .A(AES_CORE_DATAPATH__abc_16259_n8783), .B(AES_CORE_DATAPATH__abc_16259_n8785), .Y(AES_CORE_DATAPATH__abc_16259_n8786) );
  OR2X2 OR2X2_2866 ( .A(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf5), .B(AES_CORE_DATAPATH_bkp_3__19_), .Y(AES_CORE_DATAPATH__abc_16259_n8787) );
  OR2X2 OR2X2_2867 ( .A(AES_CORE_DATAPATH__abc_16259_n7122), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n8789) );
  OR2X2 OR2X2_2868 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf8), .B(AES_CORE_DATAPATH_bkp_1_3__20_), .Y(AES_CORE_DATAPATH__abc_16259_n8790) );
  OR2X2 OR2X2_2869 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n8793), .Y(AES_CORE_DATAPATH__abc_16259_n8794) );
  OR2X2 OR2X2_287 ( .A(AES_CORE_DATAPATH__abc_16259_n2970), .B(AES_CORE_DATAPATH__abc_16259_n2967_1), .Y(AES_CORE_DATAPATH__abc_16259_n2971) );
  OR2X2 OR2X2_2870 ( .A(AES_CORE_DATAPATH__abc_16259_n8792), .B(AES_CORE_DATAPATH__abc_16259_n8794), .Y(AES_CORE_DATAPATH__abc_16259_n8795) );
  OR2X2 OR2X2_2871 ( .A(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf4), .B(AES_CORE_DATAPATH_bkp_3__20_), .Y(AES_CORE_DATAPATH__abc_16259_n8796) );
  OR2X2 OR2X2_2872 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf6), .B(AES_CORE_DATAPATH_bkp_1_3__21_), .Y(AES_CORE_DATAPATH__abc_16259_n8800) );
  OR2X2 OR2X2_2873 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n8803), .Y(AES_CORE_DATAPATH__abc_16259_n8804) );
  OR2X2 OR2X2_2874 ( .A(AES_CORE_DATAPATH__abc_16259_n8802), .B(AES_CORE_DATAPATH__abc_16259_n8804), .Y(AES_CORE_DATAPATH__abc_16259_n8805) );
  OR2X2 OR2X2_2875 ( .A(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf3), .B(AES_CORE_DATAPATH_bkp_3__21_), .Y(AES_CORE_DATAPATH__abc_16259_n8806) );
  OR2X2 OR2X2_2876 ( .A(AES_CORE_DATAPATH__abc_16259_n7225), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n8808) );
  OR2X2 OR2X2_2877 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf5), .B(AES_CORE_DATAPATH_bkp_1_3__22_), .Y(AES_CORE_DATAPATH__abc_16259_n8809) );
  OR2X2 OR2X2_2878 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n8812), .Y(AES_CORE_DATAPATH__abc_16259_n8813) );
  OR2X2 OR2X2_2879 ( .A(AES_CORE_DATAPATH__abc_16259_n8811), .B(AES_CORE_DATAPATH__abc_16259_n8813), .Y(AES_CORE_DATAPATH__abc_16259_n8814) );
  OR2X2 OR2X2_288 ( .A(AES_CORE_DATAPATH__abc_16259_n2841_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__3_), .Y(AES_CORE_DATAPATH__abc_16259_n2972) );
  OR2X2 OR2X2_2880 ( .A(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf2), .B(AES_CORE_DATAPATH_bkp_3__22_), .Y(AES_CORE_DATAPATH__abc_16259_n8815) );
  OR2X2 OR2X2_2881 ( .A(AES_CORE_DATAPATH__abc_16259_n7274), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n8817) );
  OR2X2 OR2X2_2882 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf4), .B(AES_CORE_DATAPATH_bkp_1_3__23_), .Y(AES_CORE_DATAPATH__abc_16259_n8818) );
  OR2X2 OR2X2_2883 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf6), .B(AES_CORE_DATAPATH__abc_16259_n8821), .Y(AES_CORE_DATAPATH__abc_16259_n8822) );
  OR2X2 OR2X2_2884 ( .A(AES_CORE_DATAPATH__abc_16259_n8820), .B(AES_CORE_DATAPATH__abc_16259_n8822), .Y(AES_CORE_DATAPATH__abc_16259_n8823) );
  OR2X2 OR2X2_2885 ( .A(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf1), .B(AES_CORE_DATAPATH_bkp_3__23_), .Y(AES_CORE_DATAPATH__abc_16259_n8824) );
  OR2X2 OR2X2_2886 ( .A(AES_CORE_DATAPATH__abc_16259_n7323), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n8826) );
  OR2X2 OR2X2_2887 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1_3__24_), .Y(AES_CORE_DATAPATH__abc_16259_n8827) );
  OR2X2 OR2X2_2888 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf5), .B(AES_CORE_DATAPATH__abc_16259_n8830), .Y(AES_CORE_DATAPATH__abc_16259_n8831) );
  OR2X2 OR2X2_2889 ( .A(AES_CORE_DATAPATH__abc_16259_n8829), .B(AES_CORE_DATAPATH__abc_16259_n8831), .Y(AES_CORE_DATAPATH__abc_16259_n8832) );
  OR2X2 OR2X2_289 ( .A(AES_CORE_DATAPATH__abc_16259_n2964), .B(AES_CORE_DATAPATH__abc_16259_n2853_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n2974_1) );
  OR2X2 OR2X2_2890 ( .A(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf0), .B(AES_CORE_DATAPATH_bkp_3__24_), .Y(AES_CORE_DATAPATH__abc_16259_n8833) );
  OR2X2 OR2X2_2891 ( .A(AES_CORE_DATAPATH__abc_16259_n7372), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n8835) );
  OR2X2 OR2X2_2892 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf2), .B(AES_CORE_DATAPATH_bkp_1_3__25_), .Y(AES_CORE_DATAPATH__abc_16259_n8836) );
  OR2X2 OR2X2_2893 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n8839), .Y(AES_CORE_DATAPATH__abc_16259_n8840) );
  OR2X2 OR2X2_2894 ( .A(AES_CORE_DATAPATH__abc_16259_n8838), .B(AES_CORE_DATAPATH__abc_16259_n8840), .Y(AES_CORE_DATAPATH__abc_16259_n8841) );
  OR2X2 OR2X2_2895 ( .A(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf7), .B(AES_CORE_DATAPATH_bkp_3__25_), .Y(AES_CORE_DATAPATH__abc_16259_n8842) );
  OR2X2 OR2X2_2896 ( .A(AES_CORE_DATAPATH__abc_16259_n7421), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf9), .Y(AES_CORE_DATAPATH__abc_16259_n8844) );
  OR2X2 OR2X2_2897 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf1), .B(AES_CORE_DATAPATH_bkp_1_3__26_), .Y(AES_CORE_DATAPATH__abc_16259_n8845) );
  OR2X2 OR2X2_2898 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n8848), .Y(AES_CORE_DATAPATH__abc_16259_n8849) );
  OR2X2 OR2X2_2899 ( .A(AES_CORE_DATAPATH__abc_16259_n8847), .B(AES_CORE_DATAPATH__abc_16259_n8849), .Y(AES_CORE_DATAPATH__abc_16259_n8850) );
  OR2X2 OR2X2_29 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n151), .B(AES_CORE_CONTROL_UNIT__abc_15841_n152), .Y(AES_CORE_CONTROL_UNIT__abc_10818_n112) );
  OR2X2 OR2X2_290 ( .A(AES_CORE_DATAPATH__abc_16259_n2975_1), .B(AES_CORE_DATAPATH__abc_16259_n2976), .Y(AES_CORE_DATAPATH__abc_16259_n2977) );
  OR2X2 OR2X2_2900 ( .A(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf6), .B(AES_CORE_DATAPATH_bkp_3__26_), .Y(AES_CORE_DATAPATH__abc_16259_n8851) );
  OR2X2 OR2X2_2901 ( .A(AES_CORE_DATAPATH__abc_16259_n7470), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf8), .Y(AES_CORE_DATAPATH__abc_16259_n8853) );
  OR2X2 OR2X2_2902 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf0), .B(AES_CORE_DATAPATH_bkp_1_3__27_), .Y(AES_CORE_DATAPATH__abc_16259_n8854) );
  OR2X2 OR2X2_2903 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n8857), .Y(AES_CORE_DATAPATH__abc_16259_n8858) );
  OR2X2 OR2X2_2904 ( .A(AES_CORE_DATAPATH__abc_16259_n8856), .B(AES_CORE_DATAPATH__abc_16259_n8858), .Y(AES_CORE_DATAPATH__abc_16259_n8859) );
  OR2X2 OR2X2_2905 ( .A(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf5), .B(AES_CORE_DATAPATH_bkp_3__27_), .Y(AES_CORE_DATAPATH__abc_16259_n8860) );
  OR2X2 OR2X2_2906 ( .A(AES_CORE_DATAPATH__abc_16259_n7519), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n8862) );
  OR2X2 OR2X2_2907 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf11), .B(AES_CORE_DATAPATH_bkp_1_3__28_), .Y(AES_CORE_DATAPATH__abc_16259_n8863) );
  OR2X2 OR2X2_2908 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n8866), .Y(AES_CORE_DATAPATH__abc_16259_n8867) );
  OR2X2 OR2X2_2909 ( .A(AES_CORE_DATAPATH__abc_16259_n8865), .B(AES_CORE_DATAPATH__abc_16259_n8867), .Y(AES_CORE_DATAPATH__abc_16259_n8868) );
  OR2X2 OR2X2_291 ( .A(_auto_iopadmap_cc_313_execute_26949_3_), .B(AES_CORE_DATAPATH__abc_16259_n2979), .Y(AES_CORE_DATAPATH__abc_16259_n2980_1) );
  OR2X2 OR2X2_2910 ( .A(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf4), .B(AES_CORE_DATAPATH_bkp_3__28_), .Y(AES_CORE_DATAPATH__abc_16259_n8869) );
  OR2X2 OR2X2_2911 ( .A(AES_CORE_DATAPATH__abc_16259_n7568), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n8871) );
  OR2X2 OR2X2_2912 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf10), .B(AES_CORE_DATAPATH_bkp_1_3__29_), .Y(AES_CORE_DATAPATH__abc_16259_n8872) );
  OR2X2 OR2X2_2913 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n8875), .Y(AES_CORE_DATAPATH__abc_16259_n8876) );
  OR2X2 OR2X2_2914 ( .A(AES_CORE_DATAPATH__abc_16259_n8874), .B(AES_CORE_DATAPATH__abc_16259_n8876), .Y(AES_CORE_DATAPATH__abc_16259_n8877) );
  OR2X2 OR2X2_2915 ( .A(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf3), .B(AES_CORE_DATAPATH_bkp_3__29_), .Y(AES_CORE_DATAPATH__abc_16259_n8878) );
  OR2X2 OR2X2_2916 ( .A(AES_CORE_DATAPATH__abc_16259_n7617), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n8880) );
  OR2X2 OR2X2_2917 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf9), .B(AES_CORE_DATAPATH_bkp_1_3__30_), .Y(AES_CORE_DATAPATH__abc_16259_n8881) );
  OR2X2 OR2X2_2918 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf6), .B(AES_CORE_DATAPATH__abc_16259_n8884), .Y(AES_CORE_DATAPATH__abc_16259_n8885) );
  OR2X2 OR2X2_2919 ( .A(AES_CORE_DATAPATH__abc_16259_n8883), .B(AES_CORE_DATAPATH__abc_16259_n8885), .Y(AES_CORE_DATAPATH__abc_16259_n8886) );
  OR2X2 OR2X2_292 ( .A(AES_CORE_DATAPATH__abc_16259_n2982_1), .B(AES_CORE_DATAPATH__abc_16259_n2864_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n2983) );
  OR2X2 OR2X2_2920 ( .A(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf2), .B(AES_CORE_DATAPATH_bkp_3__30_), .Y(AES_CORE_DATAPATH__abc_16259_n8887) );
  OR2X2 OR2X2_2921 ( .A(AES_CORE_DATAPATH__abc_16259_n7666), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n8889) );
  OR2X2 OR2X2_2922 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf8), .B(AES_CORE_DATAPATH_bkp_1_3__31_), .Y(AES_CORE_DATAPATH__abc_16259_n8890) );
  OR2X2 OR2X2_2923 ( .A(AES_CORE_DATAPATH__abc_16259_n8500_bF_buf5), .B(AES_CORE_DATAPATH__abc_16259_n8893), .Y(AES_CORE_DATAPATH__abc_16259_n8894) );
  OR2X2 OR2X2_2924 ( .A(AES_CORE_DATAPATH__abc_16259_n8892), .B(AES_CORE_DATAPATH__abc_16259_n8894), .Y(AES_CORE_DATAPATH__abc_16259_n8895) );
  OR2X2 OR2X2_2925 ( .A(AES_CORE_DATAPATH__abc_16259_n8499_bF_buf1), .B(AES_CORE_DATAPATH_bkp_3__31_), .Y(AES_CORE_DATAPATH__abc_16259_n8896) );
  OR2X2 OR2X2_2926 ( .A(AES_CORE_CONTROL_UNIT_iv_cnt_en), .B(\iv_en[3] ), .Y(AES_CORE_DATAPATH__abc_16259_n8898) );
  OR2X2 OR2X2_2927 ( .A(AES_CORE_DATAPATH__abc_16259_n8899_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n8900_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n8901) );
  OR2X2 OR2X2_2928 ( .A(AES_CORE_DATAPATH__abc_16259_n8902), .B(AES_CORE_DATAPATH_iv_3__0_), .Y(AES_CORE_DATAPATH__abc_16259_n8903) );
  OR2X2 OR2X2_2929 ( .A(\bus_in[0] ), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .Y(AES_CORE_DATAPATH__abc_16259_n8904) );
  OR2X2 OR2X2_293 ( .A(AES_CORE_DATAPATH__abc_16259_n2983), .B(AES_CORE_DATAPATH__abc_16259_n2981), .Y(AES_CORE_DATAPATH__abc_16259_n2984_1) );
  OR2X2 OR2X2_2930 ( .A(AES_CORE_DATAPATH__abc_16259_n8908), .B(AES_CORE_DATAPATH__abc_16259_n8899_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n8909) );
  OR2X2 OR2X2_2931 ( .A(\bus_in[1] ), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .Y(AES_CORE_DATAPATH__abc_16259_n8911) );
  OR2X2 OR2X2_2932 ( .A(AES_CORE_DATAPATH__abc_16259_n8916), .B(AES_CORE_DATAPATH__abc_16259_n8899_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n8917) );
  OR2X2 OR2X2_2933 ( .A(AES_CORE_DATAPATH__abc_16259_n8919), .B(AES_CORE_DATAPATH__abc_16259_n8918_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n8920) );
  OR2X2 OR2X2_2934 ( .A(AES_CORE_DATAPATH__abc_16259_n8921), .B(AES_CORE_DATAPATH_iv_3__1_), .Y(AES_CORE_DATAPATH__abc_16259_n8922) );
  OR2X2 OR2X2_2935 ( .A(AES_CORE_DATAPATH__abc_16259_n8913), .B(AES_CORE_DATAPATH__abc_16259_n8918_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n8924) );
  OR2X2 OR2X2_2936 ( .A(AES_CORE_DATAPATH__abc_16259_n8925), .B(AES_CORE_DATAPATH_iv_3__2_), .Y(AES_CORE_DATAPATH__abc_16259_n8926) );
  OR2X2 OR2X2_2937 ( .A(\bus_in[2] ), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .Y(AES_CORE_DATAPATH__abc_16259_n8927) );
  OR2X2 OR2X2_2938 ( .A(AES_CORE_DATAPATH__abc_16259_n8931), .B(AES_CORE_DATAPATH__abc_16259_n8899_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n8932) );
  OR2X2 OR2X2_2939 ( .A(AES_CORE_DATAPATH__abc_16259_n8928), .B(AES_CORE_DATAPATH__abc_16259_n8918_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n8934) );
  OR2X2 OR2X2_294 ( .A(AES_CORE_DATAPATH__abc_16259_n2986), .B(AES_CORE_DATAPATH__abc_16259_n2985), .Y(AES_CORE_DATAPATH__abc_16259_n2987) );
  OR2X2 OR2X2_2940 ( .A(AES_CORE_DATAPATH__abc_16259_n8935), .B(AES_CORE_DATAPATH_iv_3__3_), .Y(AES_CORE_DATAPATH__abc_16259_n8936) );
  OR2X2 OR2X2_2941 ( .A(\bus_in[3] ), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .Y(AES_CORE_DATAPATH__abc_16259_n8937) );
  OR2X2 OR2X2_2942 ( .A(AES_CORE_DATAPATH__abc_16259_n8943), .B(AES_CORE_DATAPATH__abc_16259_n8899_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n8944) );
  OR2X2 OR2X2_2943 ( .A(AES_CORE_DATAPATH__abc_16259_n8940), .B(AES_CORE_DATAPATH__abc_16259_n8918_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n8946) );
  OR2X2 OR2X2_2944 ( .A(AES_CORE_DATAPATH__abc_16259_n8947), .B(AES_CORE_DATAPATH_iv_3__4_), .Y(AES_CORE_DATAPATH__abc_16259_n8948) );
  OR2X2 OR2X2_2945 ( .A(\bus_in[4] ), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .Y(AES_CORE_DATAPATH__abc_16259_n8949) );
  OR2X2 OR2X2_2946 ( .A(AES_CORE_DATAPATH__abc_16259_n8953), .B(AES_CORE_DATAPATH__abc_16259_n8899_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n8954) );
  OR2X2 OR2X2_2947 ( .A(AES_CORE_DATAPATH__abc_16259_n8950), .B(AES_CORE_DATAPATH__abc_16259_n8956), .Y(AES_CORE_DATAPATH__abc_16259_n8957) );
  OR2X2 OR2X2_2948 ( .A(AES_CORE_DATAPATH__abc_16259_n8958), .B(AES_CORE_DATAPATH_iv_3__5_), .Y(AES_CORE_DATAPATH__abc_16259_n8959) );
  OR2X2 OR2X2_2949 ( .A(AES_CORE_DATAPATH__abc_16259_n8899_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n8956), .Y(AES_CORE_DATAPATH__abc_16259_n8964) );
  OR2X2 OR2X2_295 ( .A(AES_CORE_DATAPATH__abc_16259_n2987), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n2988) );
  OR2X2 OR2X2_2950 ( .A(AES_CORE_DATAPATH__abc_16259_n8963), .B(AES_CORE_DATAPATH__abc_16259_n8964), .Y(AES_CORE_DATAPATH__abc_16259_n8965) );
  OR2X2 OR2X2_2951 ( .A(\bus_in[6] ), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .Y(AES_CORE_DATAPATH__abc_16259_n8968) );
  OR2X2 OR2X2_2952 ( .A(AES_CORE_DATAPATH__abc_16259_n8970), .B(AES_CORE_DATAPATH__abc_16259_n8972), .Y(AES_CORE_DATAPATH__abc_16259_n8973) );
  OR2X2 OR2X2_2953 ( .A(AES_CORE_DATAPATH__abc_16259_n8973), .B(AES_CORE_DATAPATH__abc_16259_n8918_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n8974) );
  OR2X2 OR2X2_2954 ( .A(AES_CORE_DATAPATH__abc_16259_n8975), .B(AES_CORE_DATAPATH__abc_16259_n8967), .Y(AES_CORE_DATAPATH__0iv_3__31_0__6_) );
  OR2X2 OR2X2_2955 ( .A(AES_CORE_DATAPATH__abc_16259_n8983), .B(AES_CORE_DATAPATH__abc_16259_n8977), .Y(AES_CORE_DATAPATH__abc_16259_n8984) );
  OR2X2 OR2X2_2956 ( .A(AES_CORE_DATAPATH__abc_16259_n8982), .B(AES_CORE_DATAPATH__abc_16259_n8901), .Y(AES_CORE_DATAPATH__abc_16259_n8986) );
  OR2X2 OR2X2_2957 ( .A(AES_CORE_DATAPATH__abc_16259_n8985), .B(AES_CORE_DATAPATH__abc_16259_n8987), .Y(AES_CORE_DATAPATH__0iv_3__31_0__7_) );
  OR2X2 OR2X2_2958 ( .A(AES_CORE_DATAPATH__abc_16259_n8993), .B(AES_CORE_DATAPATH__abc_16259_n8989), .Y(AES_CORE_DATAPATH__abc_16259_n8994) );
  OR2X2 OR2X2_2959 ( .A(AES_CORE_DATAPATH__abc_16259_n8992), .B(AES_CORE_DATAPATH__abc_16259_n8901), .Y(AES_CORE_DATAPATH__abc_16259_n8996) );
  OR2X2 OR2X2_296 ( .A(AES_CORE_DATAPATH__abc_16259_n2990), .B(AES_CORE_DATAPATH__abc_16259_n2991), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_3_) );
  OR2X2 OR2X2_2960 ( .A(AES_CORE_DATAPATH__abc_16259_n8995), .B(AES_CORE_DATAPATH__abc_16259_n8997), .Y(AES_CORE_DATAPATH__0iv_3__31_0__8_) );
  OR2X2 OR2X2_2961 ( .A(AES_CORE_DATAPATH__abc_16259_n8898_bF_buf0), .B(AES_CORE_DATAPATH_iv_3__9_), .Y(AES_CORE_DATAPATH__abc_16259_n8999) );
  OR2X2 OR2X2_2962 ( .A(AES_CORE_DATAPATH__abc_16259_n8990), .B(AES_CORE_DATAPATH_iv_3__9_), .Y(AES_CORE_DATAPATH__abc_16259_n9000) );
  OR2X2 OR2X2_2963 ( .A(AES_CORE_DATAPATH__abc_16259_n9005), .B(AES_CORE_DATAPATH__abc_16259_n9001), .Y(AES_CORE_DATAPATH__abc_16259_n9006) );
  OR2X2 OR2X2_2964 ( .A(AES_CORE_DATAPATH__abc_16259_n8899_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n9008), .Y(AES_CORE_DATAPATH__abc_16259_n9009) );
  OR2X2 OR2X2_2965 ( .A(AES_CORE_DATAPATH__abc_16259_n9007), .B(AES_CORE_DATAPATH__abc_16259_n9009), .Y(AES_CORE_DATAPATH__abc_16259_n9010) );
  OR2X2 OR2X2_2966 ( .A(AES_CORE_DATAPATH__abc_16259_n8898_bF_buf4), .B(AES_CORE_DATAPATH_iv_3__10_), .Y(AES_CORE_DATAPATH__abc_16259_n9012) );
  OR2X2 OR2X2_2967 ( .A(AES_CORE_DATAPATH__abc_16259_n9003), .B(AES_CORE_DATAPATH_iv_3__10_), .Y(AES_CORE_DATAPATH__abc_16259_n9013) );
  OR2X2 OR2X2_2968 ( .A(AES_CORE_DATAPATH__abc_16259_n9018), .B(AES_CORE_DATAPATH__abc_16259_n9019), .Y(AES_CORE_DATAPATH__abc_16259_n9020) );
  OR2X2 OR2X2_2969 ( .A(AES_CORE_DATAPATH__abc_16259_n9020), .B(AES_CORE_DATAPATH__abc_16259_n8899_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n9021) );
  OR2X2 OR2X2_297 ( .A(AES_CORE_DATAPATH__abc_16259_n2774_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n2993), .Y(AES_CORE_DATAPATH__abc_16259_n2994) );
  OR2X2 OR2X2_2970 ( .A(AES_CORE_DATAPATH__abc_16259_n9017), .B(AES_CORE_DATAPATH__abc_16259_n9021), .Y(AES_CORE_DATAPATH__abc_16259_n9022) );
  OR2X2 OR2X2_2971 ( .A(AES_CORE_DATAPATH__abc_16259_n8898_bF_buf3), .B(AES_CORE_DATAPATH_iv_3__11_), .Y(AES_CORE_DATAPATH__abc_16259_n9024) );
  OR2X2 OR2X2_2972 ( .A(AES_CORE_DATAPATH__abc_16259_n9014), .B(AES_CORE_DATAPATH_iv_3__11_), .Y(AES_CORE_DATAPATH__abc_16259_n9025) );
  OR2X2 OR2X2_2973 ( .A(AES_CORE_DATAPATH__abc_16259_n9029), .B(AES_CORE_DATAPATH__abc_16259_n9026), .Y(AES_CORE_DATAPATH__abc_16259_n9030) );
  OR2X2 OR2X2_2974 ( .A(AES_CORE_DATAPATH__abc_16259_n8899_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n9032), .Y(AES_CORE_DATAPATH__abc_16259_n9033) );
  OR2X2 OR2X2_2975 ( .A(AES_CORE_DATAPATH__abc_16259_n9031), .B(AES_CORE_DATAPATH__abc_16259_n9033), .Y(AES_CORE_DATAPATH__abc_16259_n9034) );
  OR2X2 OR2X2_2976 ( .A(AES_CORE_DATAPATH__abc_16259_n8898_bF_buf2), .B(AES_CORE_DATAPATH_iv_3__12_), .Y(AES_CORE_DATAPATH__abc_16259_n9036) );
  OR2X2 OR2X2_2977 ( .A(AES_CORE_DATAPATH__abc_16259_n9027), .B(AES_CORE_DATAPATH_iv_3__12_), .Y(AES_CORE_DATAPATH__abc_16259_n9039) );
  OR2X2 OR2X2_2978 ( .A(AES_CORE_DATAPATH__abc_16259_n8899_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n9043), .Y(AES_CORE_DATAPATH__abc_16259_n9044) );
  OR2X2 OR2X2_2979 ( .A(AES_CORE_DATAPATH__abc_16259_n9044), .B(AES_CORE_DATAPATH__abc_16259_n9042), .Y(AES_CORE_DATAPATH__abc_16259_n9045) );
  OR2X2 OR2X2_298 ( .A(AES_CORE_DATAPATH__abc_16259_n2778_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n2995), .Y(AES_CORE_DATAPATH__abc_16259_n2996_1) );
  OR2X2 OR2X2_2980 ( .A(AES_CORE_DATAPATH__abc_16259_n9041), .B(AES_CORE_DATAPATH__abc_16259_n9045), .Y(AES_CORE_DATAPATH__abc_16259_n9046) );
  OR2X2 OR2X2_2981 ( .A(AES_CORE_DATAPATH__abc_16259_n8898_bF_buf1), .B(AES_CORE_DATAPATH_iv_3__13_), .Y(AES_CORE_DATAPATH__abc_16259_n9048) );
  OR2X2 OR2X2_2982 ( .A(AES_CORE_DATAPATH__abc_16259_n9037), .B(AES_CORE_DATAPATH_iv_3__13_), .Y(AES_CORE_DATAPATH__abc_16259_n9051) );
  OR2X2 OR2X2_2983 ( .A(AES_CORE_DATAPATH__abc_16259_n8899_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n9055), .Y(AES_CORE_DATAPATH__abc_16259_n9056) );
  OR2X2 OR2X2_2984 ( .A(AES_CORE_DATAPATH__abc_16259_n9056), .B(AES_CORE_DATAPATH__abc_16259_n9054), .Y(AES_CORE_DATAPATH__abc_16259_n9057) );
  OR2X2 OR2X2_2985 ( .A(AES_CORE_DATAPATH__abc_16259_n9053), .B(AES_CORE_DATAPATH__abc_16259_n9057), .Y(AES_CORE_DATAPATH__abc_16259_n9058) );
  OR2X2 OR2X2_2986 ( .A(AES_CORE_DATAPATH__abc_16259_n8898_bF_buf0), .B(AES_CORE_DATAPATH_iv_3__14_), .Y(AES_CORE_DATAPATH__abc_16259_n9060) );
  OR2X2 OR2X2_2987 ( .A(AES_CORE_DATAPATH__abc_16259_n9049), .B(AES_CORE_DATAPATH_iv_3__14_), .Y(AES_CORE_DATAPATH__abc_16259_n9063) );
  OR2X2 OR2X2_2988 ( .A(AES_CORE_DATAPATH__abc_16259_n8899_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n9067), .Y(AES_CORE_DATAPATH__abc_16259_n9068) );
  OR2X2 OR2X2_2989 ( .A(AES_CORE_DATAPATH__abc_16259_n9068), .B(AES_CORE_DATAPATH__abc_16259_n9066), .Y(AES_CORE_DATAPATH__abc_16259_n9069) );
  OR2X2 OR2X2_299 ( .A(AES_CORE_DATAPATH__abc_16259_n2999), .B(AES_CORE_DATAPATH__abc_16259_n3000), .Y(AES_CORE_DATAPATH__abc_16259_n3001) );
  OR2X2 OR2X2_2990 ( .A(AES_CORE_DATAPATH__abc_16259_n9065), .B(AES_CORE_DATAPATH__abc_16259_n9069), .Y(AES_CORE_DATAPATH__abc_16259_n9070) );
  OR2X2 OR2X2_2991 ( .A(AES_CORE_DATAPATH__abc_16259_n8898_bF_buf4), .B(AES_CORE_DATAPATH_iv_3__15_), .Y(AES_CORE_DATAPATH__abc_16259_n9072) );
  OR2X2 OR2X2_2992 ( .A(AES_CORE_DATAPATH__abc_16259_n9061), .B(AES_CORE_DATAPATH_iv_3__15_), .Y(AES_CORE_DATAPATH__abc_16259_n9075) );
  OR2X2 OR2X2_2993 ( .A(AES_CORE_DATAPATH__abc_16259_n8899_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n9079), .Y(AES_CORE_DATAPATH__abc_16259_n9080) );
  OR2X2 OR2X2_2994 ( .A(AES_CORE_DATAPATH__abc_16259_n9080), .B(AES_CORE_DATAPATH__abc_16259_n9078), .Y(AES_CORE_DATAPATH__abc_16259_n9081) );
  OR2X2 OR2X2_2995 ( .A(AES_CORE_DATAPATH__abc_16259_n9077), .B(AES_CORE_DATAPATH__abc_16259_n9081), .Y(AES_CORE_DATAPATH__abc_16259_n9082) );
  OR2X2 OR2X2_2996 ( .A(AES_CORE_DATAPATH__abc_16259_n8898_bF_buf3), .B(AES_CORE_DATAPATH_iv_3__16_), .Y(AES_CORE_DATAPATH__abc_16259_n9084) );
  OR2X2 OR2X2_2997 ( .A(AES_CORE_DATAPATH__abc_16259_n9073), .B(AES_CORE_DATAPATH_iv_3__16_), .Y(AES_CORE_DATAPATH__abc_16259_n9087) );
  OR2X2 OR2X2_2998 ( .A(AES_CORE_DATAPATH__abc_16259_n8899_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n9091), .Y(AES_CORE_DATAPATH__abc_16259_n9092) );
  OR2X2 OR2X2_2999 ( .A(AES_CORE_DATAPATH__abc_16259_n9092), .B(AES_CORE_DATAPATH__abc_16259_n9090), .Y(AES_CORE_DATAPATH__abc_16259_n9093) );
  OR2X2 OR2X2_3 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr_bF_buf5), .B(AES_CORE_CONTROL_UNIT__abc_15841_n77), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n78) );
  OR2X2 OR2X2_30 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n155_1), .B(AES_CORE_CONTROL_UNIT__abc_15841_n156), .Y(AES_CORE_CONTROL_UNIT__abc_10818_n118) );
  OR2X2 OR2X2_300 ( .A(AES_CORE_DATAPATH__abc_16259_n3001), .B(AES_CORE_DATAPATH__abc_16259_n2998_1), .Y(AES_CORE_DATAPATH__abc_16259_n3002) );
  OR2X2 OR2X2_3000 ( .A(AES_CORE_DATAPATH__abc_16259_n9089), .B(AES_CORE_DATAPATH__abc_16259_n9093), .Y(AES_CORE_DATAPATH__abc_16259_n9094) );
  OR2X2 OR2X2_3001 ( .A(AES_CORE_DATAPATH__abc_16259_n8898_bF_buf2), .B(AES_CORE_DATAPATH_iv_3__17_), .Y(AES_CORE_DATAPATH__abc_16259_n9096) );
  OR2X2 OR2X2_3002 ( .A(AES_CORE_DATAPATH__abc_16259_n9085), .B(AES_CORE_DATAPATH_iv_3__17_), .Y(AES_CORE_DATAPATH__abc_16259_n9099) );
  OR2X2 OR2X2_3003 ( .A(AES_CORE_DATAPATH__abc_16259_n8899_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n9103), .Y(AES_CORE_DATAPATH__abc_16259_n9104) );
  OR2X2 OR2X2_3004 ( .A(AES_CORE_DATAPATH__abc_16259_n9104), .B(AES_CORE_DATAPATH__abc_16259_n9102), .Y(AES_CORE_DATAPATH__abc_16259_n9105) );
  OR2X2 OR2X2_3005 ( .A(AES_CORE_DATAPATH__abc_16259_n9101), .B(AES_CORE_DATAPATH__abc_16259_n9105), .Y(AES_CORE_DATAPATH__abc_16259_n9106) );
  OR2X2 OR2X2_3006 ( .A(AES_CORE_DATAPATH__abc_16259_n8898_bF_buf1), .B(AES_CORE_DATAPATH_iv_3__18_), .Y(AES_CORE_DATAPATH__abc_16259_n9108) );
  OR2X2 OR2X2_3007 ( .A(AES_CORE_DATAPATH__abc_16259_n9097), .B(AES_CORE_DATAPATH_iv_3__18_), .Y(AES_CORE_DATAPATH__abc_16259_n9109) );
  OR2X2 OR2X2_3008 ( .A(AES_CORE_DATAPATH__abc_16259_n8899_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n9116), .Y(AES_CORE_DATAPATH__abc_16259_n9117) );
  OR2X2 OR2X2_3009 ( .A(AES_CORE_DATAPATH__abc_16259_n9117), .B(AES_CORE_DATAPATH__abc_16259_n9115), .Y(AES_CORE_DATAPATH__abc_16259_n9118) );
  OR2X2 OR2X2_301 ( .A(AES_CORE_DATAPATH__abc_16259_n3006), .B(AES_CORE_DATAPATH__abc_16259_n2826_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n3007_1) );
  OR2X2 OR2X2_3010 ( .A(AES_CORE_DATAPATH__abc_16259_n9114), .B(AES_CORE_DATAPATH__abc_16259_n9118), .Y(AES_CORE_DATAPATH__abc_16259_n9119) );
  OR2X2 OR2X2_3011 ( .A(AES_CORE_DATAPATH__abc_16259_n8898_bF_buf0), .B(AES_CORE_DATAPATH_iv_3__19_), .Y(AES_CORE_DATAPATH__abc_16259_n9121) );
  OR2X2 OR2X2_3012 ( .A(AES_CORE_DATAPATH__abc_16259_n9111), .B(AES_CORE_DATAPATH_iv_3__19_), .Y(AES_CORE_DATAPATH__abc_16259_n9124) );
  OR2X2 OR2X2_3013 ( .A(AES_CORE_DATAPATH__abc_16259_n8899_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n9128), .Y(AES_CORE_DATAPATH__abc_16259_n9129) );
  OR2X2 OR2X2_3014 ( .A(AES_CORE_DATAPATH__abc_16259_n9129), .B(AES_CORE_DATAPATH__abc_16259_n9127), .Y(AES_CORE_DATAPATH__abc_16259_n9130) );
  OR2X2 OR2X2_3015 ( .A(AES_CORE_DATAPATH__abc_16259_n9126), .B(AES_CORE_DATAPATH__abc_16259_n9130), .Y(AES_CORE_DATAPATH__abc_16259_n9131) );
  OR2X2 OR2X2_3016 ( .A(AES_CORE_DATAPATH__abc_16259_n8898_bF_buf4), .B(AES_CORE_DATAPATH_iv_3__20_), .Y(AES_CORE_DATAPATH__abc_16259_n9133) );
  OR2X2 OR2X2_3017 ( .A(AES_CORE_DATAPATH__abc_16259_n9135), .B(AES_CORE_DATAPATH_iv_3__20_), .Y(AES_CORE_DATAPATH__abc_16259_n9136) );
  OR2X2 OR2X2_3018 ( .A(AES_CORE_DATAPATH__abc_16259_n8899_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n9142), .Y(AES_CORE_DATAPATH__abc_16259_n9143) );
  OR2X2 OR2X2_3019 ( .A(AES_CORE_DATAPATH__abc_16259_n9143), .B(AES_CORE_DATAPATH__abc_16259_n9141), .Y(AES_CORE_DATAPATH__abc_16259_n9144) );
  OR2X2 OR2X2_302 ( .A(AES_CORE_DATAPATH__abc_16259_n3008), .B(AES_CORE_DATAPATH__abc_16259_n3009_1), .Y(AES_CORE_DATAPATH__abc_16259_n3010) );
  OR2X2 OR2X2_3020 ( .A(AES_CORE_DATAPATH__abc_16259_n9140), .B(AES_CORE_DATAPATH__abc_16259_n9144), .Y(AES_CORE_DATAPATH__abc_16259_n9145) );
  OR2X2 OR2X2_3021 ( .A(AES_CORE_DATAPATH__abc_16259_n8898_bF_buf3), .B(AES_CORE_DATAPATH_iv_3__21_), .Y(AES_CORE_DATAPATH__abc_16259_n9147) );
  OR2X2 OR2X2_3022 ( .A(AES_CORE_DATAPATH__abc_16259_n9148), .B(AES_CORE_DATAPATH__abc_16259_n9150), .Y(AES_CORE_DATAPATH__abc_16259_n9151) );
  OR2X2 OR2X2_3023 ( .A(AES_CORE_DATAPATH__abc_16259_n8899_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n9154), .Y(AES_CORE_DATAPATH__abc_16259_n9155) );
  OR2X2 OR2X2_3024 ( .A(AES_CORE_DATAPATH__abc_16259_n9155), .B(AES_CORE_DATAPATH__abc_16259_n9153), .Y(AES_CORE_DATAPATH__abc_16259_n9156) );
  OR2X2 OR2X2_3025 ( .A(AES_CORE_DATAPATH__abc_16259_n9152), .B(AES_CORE_DATAPATH__abc_16259_n9156), .Y(AES_CORE_DATAPATH__abc_16259_n9157) );
  OR2X2 OR2X2_3026 ( .A(AES_CORE_DATAPATH__abc_16259_n8898_bF_buf2), .B(AES_CORE_DATAPATH_iv_3__22_), .Y(AES_CORE_DATAPATH__abc_16259_n9159) );
  OR2X2 OR2X2_3027 ( .A(AES_CORE_DATAPATH__abc_16259_n9160), .B(AES_CORE_DATAPATH_iv_3__22_), .Y(AES_CORE_DATAPATH__abc_16259_n9161) );
  OR2X2 OR2X2_3028 ( .A(AES_CORE_DATAPATH__abc_16259_n8899_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n9169), .Y(AES_CORE_DATAPATH__abc_16259_n9170) );
  OR2X2 OR2X2_3029 ( .A(AES_CORE_DATAPATH__abc_16259_n9170), .B(AES_CORE_DATAPATH__abc_16259_n9168), .Y(AES_CORE_DATAPATH__abc_16259_n9171) );
  OR2X2 OR2X2_303 ( .A(AES_CORE_DATAPATH__abc_16259_n3010), .B(AES_CORE_DATAPATH__abc_16259_n3007_1), .Y(AES_CORE_DATAPATH__abc_16259_n3011_1) );
  OR2X2 OR2X2_3030 ( .A(AES_CORE_DATAPATH__abc_16259_n9167), .B(AES_CORE_DATAPATH__abc_16259_n9171), .Y(AES_CORE_DATAPATH__abc_16259_n9172) );
  OR2X2 OR2X2_3031 ( .A(AES_CORE_DATAPATH__abc_16259_n8898_bF_buf1), .B(AES_CORE_DATAPATH_iv_3__23_), .Y(AES_CORE_DATAPATH__abc_16259_n9174) );
  OR2X2 OR2X2_3032 ( .A(AES_CORE_DATAPATH__abc_16259_n9164), .B(AES_CORE_DATAPATH_iv_3__23_), .Y(AES_CORE_DATAPATH__abc_16259_n9177) );
  OR2X2 OR2X2_3033 ( .A(AES_CORE_DATAPATH__abc_16259_n8899_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n9181), .Y(AES_CORE_DATAPATH__abc_16259_n9182) );
  OR2X2 OR2X2_3034 ( .A(AES_CORE_DATAPATH__abc_16259_n9182), .B(AES_CORE_DATAPATH__abc_16259_n9180), .Y(AES_CORE_DATAPATH__abc_16259_n9183) );
  OR2X2 OR2X2_3035 ( .A(AES_CORE_DATAPATH__abc_16259_n9179), .B(AES_CORE_DATAPATH__abc_16259_n9183), .Y(AES_CORE_DATAPATH__abc_16259_n9184) );
  OR2X2 OR2X2_3036 ( .A(AES_CORE_DATAPATH__abc_16259_n8898_bF_buf0), .B(AES_CORE_DATAPATH_iv_3__24_), .Y(AES_CORE_DATAPATH__abc_16259_n9186) );
  OR2X2 OR2X2_3037 ( .A(AES_CORE_DATAPATH__abc_16259_n9188), .B(AES_CORE_DATAPATH_iv_3__24_), .Y(AES_CORE_DATAPATH__abc_16259_n9189) );
  OR2X2 OR2X2_3038 ( .A(AES_CORE_DATAPATH__abc_16259_n8899_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n9195), .Y(AES_CORE_DATAPATH__abc_16259_n9196) );
  OR2X2 OR2X2_3039 ( .A(AES_CORE_DATAPATH__abc_16259_n9196), .B(AES_CORE_DATAPATH__abc_16259_n9194), .Y(AES_CORE_DATAPATH__abc_16259_n9197) );
  OR2X2 OR2X2_304 ( .A(AES_CORE_DATAPATH__abc_16259_n2841_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__4_), .Y(AES_CORE_DATAPATH__abc_16259_n3012) );
  OR2X2 OR2X2_3040 ( .A(AES_CORE_DATAPATH__abc_16259_n9193), .B(AES_CORE_DATAPATH__abc_16259_n9197), .Y(AES_CORE_DATAPATH__abc_16259_n9198) );
  OR2X2 OR2X2_3041 ( .A(AES_CORE_DATAPATH__abc_16259_n8898_bF_buf4), .B(AES_CORE_DATAPATH_iv_3__25_), .Y(AES_CORE_DATAPATH__abc_16259_n9200) );
  OR2X2 OR2X2_3042 ( .A(AES_CORE_DATAPATH__abc_16259_n9201), .B(AES_CORE_DATAPATH__abc_16259_n9203), .Y(AES_CORE_DATAPATH__abc_16259_n9204) );
  OR2X2 OR2X2_3043 ( .A(AES_CORE_DATAPATH__abc_16259_n8899_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n9207), .Y(AES_CORE_DATAPATH__abc_16259_n9208) );
  OR2X2 OR2X2_3044 ( .A(AES_CORE_DATAPATH__abc_16259_n9208), .B(AES_CORE_DATAPATH__abc_16259_n9206), .Y(AES_CORE_DATAPATH__abc_16259_n9209) );
  OR2X2 OR2X2_3045 ( .A(AES_CORE_DATAPATH__abc_16259_n9205), .B(AES_CORE_DATAPATH__abc_16259_n9209), .Y(AES_CORE_DATAPATH__abc_16259_n9210) );
  OR2X2 OR2X2_3046 ( .A(AES_CORE_DATAPATH__abc_16259_n8898_bF_buf3), .B(AES_CORE_DATAPATH_iv_3__26_), .Y(AES_CORE_DATAPATH__abc_16259_n9212) );
  OR2X2 OR2X2_3047 ( .A(AES_CORE_DATAPATH__abc_16259_n9213), .B(AES_CORE_DATAPATH_iv_3__26_), .Y(AES_CORE_DATAPATH__abc_16259_n9214) );
  OR2X2 OR2X2_3048 ( .A(AES_CORE_DATAPATH__abc_16259_n8899_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n9220), .Y(AES_CORE_DATAPATH__abc_16259_n9221) );
  OR2X2 OR2X2_3049 ( .A(AES_CORE_DATAPATH__abc_16259_n9221), .B(AES_CORE_DATAPATH__abc_16259_n9219), .Y(AES_CORE_DATAPATH__abc_16259_n9222) );
  OR2X2 OR2X2_305 ( .A(AES_CORE_DATAPATH__abc_16259_n3004_1), .B(AES_CORE_DATAPATH__abc_16259_n2853_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n3014) );
  OR2X2 OR2X2_3050 ( .A(AES_CORE_DATAPATH__abc_16259_n9218), .B(AES_CORE_DATAPATH__abc_16259_n9222), .Y(AES_CORE_DATAPATH__abc_16259_n9223) );
  OR2X2 OR2X2_3051 ( .A(AES_CORE_DATAPATH__abc_16259_n8898_bF_buf2), .B(AES_CORE_DATAPATH_iv_3__27_), .Y(AES_CORE_DATAPATH__abc_16259_n9225) );
  OR2X2 OR2X2_3052 ( .A(AES_CORE_DATAPATH__abc_16259_n9215), .B(AES_CORE_DATAPATH_iv_3__27_), .Y(AES_CORE_DATAPATH__abc_16259_n9226) );
  OR2X2 OR2X2_3053 ( .A(AES_CORE_DATAPATH__abc_16259_n8899_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n9232), .Y(AES_CORE_DATAPATH__abc_16259_n9233) );
  OR2X2 OR2X2_3054 ( .A(AES_CORE_DATAPATH__abc_16259_n9233), .B(AES_CORE_DATAPATH__abc_16259_n9231), .Y(AES_CORE_DATAPATH__abc_16259_n9234) );
  OR2X2 OR2X2_3055 ( .A(AES_CORE_DATAPATH__abc_16259_n9230), .B(AES_CORE_DATAPATH__abc_16259_n9234), .Y(AES_CORE_DATAPATH__abc_16259_n9235) );
  OR2X2 OR2X2_3056 ( .A(AES_CORE_DATAPATH__abc_16259_n8898_bF_buf1), .B(AES_CORE_DATAPATH_iv_3__28_), .Y(AES_CORE_DATAPATH__abc_16259_n9237) );
  OR2X2 OR2X2_3057 ( .A(AES_CORE_DATAPATH__abc_16259_n9227), .B(AES_CORE_DATAPATH_iv_3__28_), .Y(AES_CORE_DATAPATH__abc_16259_n9238) );
  OR2X2 OR2X2_3058 ( .A(AES_CORE_DATAPATH__abc_16259_n8899_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n9244), .Y(AES_CORE_DATAPATH__abc_16259_n9245) );
  OR2X2 OR2X2_3059 ( .A(AES_CORE_DATAPATH__abc_16259_n9245), .B(AES_CORE_DATAPATH__abc_16259_n9243), .Y(AES_CORE_DATAPATH__abc_16259_n9246) );
  OR2X2 OR2X2_306 ( .A(AES_CORE_DATAPATH__abc_16259_n3015), .B(AES_CORE_DATAPATH__abc_16259_n3016), .Y(AES_CORE_DATAPATH__abc_16259_n3017) );
  OR2X2 OR2X2_3060 ( .A(AES_CORE_DATAPATH__abc_16259_n9242), .B(AES_CORE_DATAPATH__abc_16259_n9246), .Y(AES_CORE_DATAPATH__abc_16259_n9247) );
  OR2X2 OR2X2_3061 ( .A(AES_CORE_DATAPATH__abc_16259_n8898_bF_buf0), .B(AES_CORE_DATAPATH_iv_3__29_), .Y(AES_CORE_DATAPATH__abc_16259_n9249) );
  OR2X2 OR2X2_3062 ( .A(AES_CORE_DATAPATH__abc_16259_n9239), .B(AES_CORE_DATAPATH_iv_3__29_), .Y(AES_CORE_DATAPATH__abc_16259_n9250) );
  OR2X2 OR2X2_3063 ( .A(AES_CORE_DATAPATH__abc_16259_n8899_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n9256), .Y(AES_CORE_DATAPATH__abc_16259_n9257) );
  OR2X2 OR2X2_3064 ( .A(AES_CORE_DATAPATH__abc_16259_n9257), .B(AES_CORE_DATAPATH__abc_16259_n9255), .Y(AES_CORE_DATAPATH__abc_16259_n9258) );
  OR2X2 OR2X2_3065 ( .A(AES_CORE_DATAPATH__abc_16259_n9254), .B(AES_CORE_DATAPATH__abc_16259_n9258), .Y(AES_CORE_DATAPATH__abc_16259_n9259) );
  OR2X2 OR2X2_3066 ( .A(AES_CORE_DATAPATH__abc_16259_n8898_bF_buf4), .B(AES_CORE_DATAPATH_iv_3__30_), .Y(AES_CORE_DATAPATH__abc_16259_n9261) );
  OR2X2 OR2X2_3067 ( .A(AES_CORE_DATAPATH__abc_16259_n9251), .B(AES_CORE_DATAPATH_iv_3__30_), .Y(AES_CORE_DATAPATH__abc_16259_n9264) );
  OR2X2 OR2X2_3068 ( .A(AES_CORE_DATAPATH__abc_16259_n8899_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n9268), .Y(AES_CORE_DATAPATH__abc_16259_n9269) );
  OR2X2 OR2X2_3069 ( .A(AES_CORE_DATAPATH__abc_16259_n9269), .B(AES_CORE_DATAPATH__abc_16259_n9267), .Y(AES_CORE_DATAPATH__abc_16259_n9270) );
  OR2X2 OR2X2_307 ( .A(_auto_iopadmap_cc_313_execute_26949_4_), .B(AES_CORE_DATAPATH__abc_16259_n3019), .Y(AES_CORE_DATAPATH__abc_16259_n3020) );
  OR2X2 OR2X2_3070 ( .A(AES_CORE_DATAPATH__abc_16259_n9266), .B(AES_CORE_DATAPATH__abc_16259_n9270), .Y(AES_CORE_DATAPATH__abc_16259_n9271) );
  OR2X2 OR2X2_3071 ( .A(AES_CORE_DATAPATH__abc_16259_n8898_bF_buf3), .B(AES_CORE_DATAPATH_iv_3__31_), .Y(AES_CORE_DATAPATH__abc_16259_n9273) );
  OR2X2 OR2X2_3072 ( .A(AES_CORE_DATAPATH__abc_16259_n9274), .B(AES_CORE_DATAPATH__abc_16259_n9276), .Y(AES_CORE_DATAPATH__abc_16259_n9277) );
  OR2X2 OR2X2_3073 ( .A(AES_CORE_DATAPATH__abc_16259_n8899_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n9280), .Y(AES_CORE_DATAPATH__abc_16259_n9281) );
  OR2X2 OR2X2_3074 ( .A(AES_CORE_DATAPATH__abc_16259_n9281), .B(AES_CORE_DATAPATH__abc_16259_n9279), .Y(AES_CORE_DATAPATH__abc_16259_n9282) );
  OR2X2 OR2X2_3075 ( .A(AES_CORE_DATAPATH__abc_16259_n9278), .B(AES_CORE_DATAPATH__abc_16259_n9282), .Y(AES_CORE_DATAPATH__abc_16259_n9283) );
  OR2X2 OR2X2_3076 ( .A(AES_CORE_DATAPATH__abc_16259_n9285), .B(AES_CORE_DATAPATH__abc_16259_n9286), .Y(AES_CORE_DATAPATH__abc_16259_n9287) );
  OR2X2 OR2X2_3077 ( .A(AES_CORE_DATAPATH__abc_16259_n9290), .B(AES_CORE_DATAPATH__abc_16259_n9289), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__0_) );
  OR2X2 OR2X2_3078 ( .A(AES_CORE_DATAPATH__abc_16259_n9293), .B(AES_CORE_DATAPATH__abc_16259_n9292), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__1_) );
  OR2X2 OR2X2_3079 ( .A(AES_CORE_DATAPATH__abc_16259_n9296), .B(AES_CORE_DATAPATH__abc_16259_n9295), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__2_) );
  OR2X2 OR2X2_308 ( .A(AES_CORE_DATAPATH__abc_16259_n3022), .B(AES_CORE_DATAPATH__abc_16259_n2864_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n3023) );
  OR2X2 OR2X2_3080 ( .A(AES_CORE_DATAPATH__abc_16259_n9299), .B(AES_CORE_DATAPATH__abc_16259_n9298), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__3_) );
  OR2X2 OR2X2_3081 ( .A(AES_CORE_DATAPATH__abc_16259_n9302), .B(AES_CORE_DATAPATH__abc_16259_n9301), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__4_) );
  OR2X2 OR2X2_3082 ( .A(AES_CORE_DATAPATH__abc_16259_n9305), .B(AES_CORE_DATAPATH__abc_16259_n9304), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__5_) );
  OR2X2 OR2X2_3083 ( .A(AES_CORE_DATAPATH__abc_16259_n9308), .B(AES_CORE_DATAPATH__abc_16259_n9307), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__6_) );
  OR2X2 OR2X2_3084 ( .A(AES_CORE_DATAPATH__abc_16259_n9311), .B(AES_CORE_DATAPATH__abc_16259_n9310), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__7_) );
  OR2X2 OR2X2_3085 ( .A(AES_CORE_DATAPATH__abc_16259_n9314), .B(AES_CORE_DATAPATH__abc_16259_n9313), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__8_) );
  OR2X2 OR2X2_3086 ( .A(AES_CORE_DATAPATH__abc_16259_n9317), .B(AES_CORE_DATAPATH__abc_16259_n9316), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__9_) );
  OR2X2 OR2X2_3087 ( .A(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1_2__10_), .Y(AES_CORE_DATAPATH__abc_16259_n9321) );
  OR2X2 OR2X2_3088 ( .A(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf1), .B(AES_CORE_DATAPATH_bkp_1_2__11_), .Y(AES_CORE_DATAPATH__abc_16259_n9325) );
  OR2X2 OR2X2_3089 ( .A(AES_CORE_DATAPATH__abc_16259_n9328), .B(AES_CORE_DATAPATH__abc_16259_n9327), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__12_) );
  OR2X2 OR2X2_309 ( .A(AES_CORE_DATAPATH__abc_16259_n3023), .B(AES_CORE_DATAPATH__abc_16259_n3021), .Y(AES_CORE_DATAPATH__abc_16259_n3024) );
  OR2X2 OR2X2_3090 ( .A(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf6), .B(AES_CORE_DATAPATH_bkp_1_2__13_), .Y(AES_CORE_DATAPATH__abc_16259_n9332) );
  OR2X2 OR2X2_3091 ( .A(AES_CORE_DATAPATH__abc_16259_n9335), .B(AES_CORE_DATAPATH__abc_16259_n9334), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__14_) );
  OR2X2 OR2X2_3092 ( .A(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1_2__15_), .Y(AES_CORE_DATAPATH__abc_16259_n9339) );
  OR2X2 OR2X2_3093 ( .A(AES_CORE_DATAPATH__abc_16259_n9342), .B(AES_CORE_DATAPATH__abc_16259_n9341), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__16_) );
  OR2X2 OR2X2_3094 ( .A(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf0), .B(AES_CORE_DATAPATH_bkp_1_2__17_), .Y(AES_CORE_DATAPATH__abc_16259_n9346) );
  OR2X2 OR2X2_3095 ( .A(AES_CORE_DATAPATH__abc_16259_n9349), .B(AES_CORE_DATAPATH__abc_16259_n9348), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__18_) );
  OR2X2 OR2X2_3096 ( .A(AES_CORE_DATAPATH__abc_16259_n9352), .B(AES_CORE_DATAPATH__abc_16259_n9351), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__19_) );
  OR2X2 OR2X2_3097 ( .A(AES_CORE_DATAPATH__abc_16259_n9355), .B(AES_CORE_DATAPATH__abc_16259_n9354), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__20_) );
  OR2X2 OR2X2_3098 ( .A(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1_2__21_), .Y(AES_CORE_DATAPATH__abc_16259_n9359) );
  OR2X2 OR2X2_3099 ( .A(AES_CORE_DATAPATH__abc_16259_n9362), .B(AES_CORE_DATAPATH__abc_16259_n9361), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__22_) );
  OR2X2 OR2X2_31 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n158), .B(AES_CORE_CONTROL_UNIT__abc_15841_n159), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n160) );
  OR2X2 OR2X2_310 ( .A(AES_CORE_DATAPATH__abc_16259_n3026), .B(AES_CORE_DATAPATH__abc_16259_n3025_1), .Y(AES_CORE_DATAPATH__abc_16259_n3027_1) );
  OR2X2 OR2X2_3100 ( .A(AES_CORE_DATAPATH__abc_16259_n9365), .B(AES_CORE_DATAPATH__abc_16259_n9364), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__23_) );
  OR2X2 OR2X2_3101 ( .A(AES_CORE_DATAPATH__abc_16259_n9368), .B(AES_CORE_DATAPATH__abc_16259_n9367), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__24_) );
  OR2X2 OR2X2_3102 ( .A(AES_CORE_DATAPATH__abc_16259_n9371), .B(AES_CORE_DATAPATH__abc_16259_n9370), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__25_) );
  OR2X2 OR2X2_3103 ( .A(AES_CORE_DATAPATH__abc_16259_n9374), .B(AES_CORE_DATAPATH__abc_16259_n9373), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__26_) );
  OR2X2 OR2X2_3104 ( .A(AES_CORE_DATAPATH__abc_16259_n9377), .B(AES_CORE_DATAPATH__abc_16259_n9376), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__27_) );
  OR2X2 OR2X2_3105 ( .A(AES_CORE_DATAPATH__abc_16259_n9380), .B(AES_CORE_DATAPATH__abc_16259_n9379), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__28_) );
  OR2X2 OR2X2_3106 ( .A(AES_CORE_DATAPATH__abc_16259_n9383), .B(AES_CORE_DATAPATH__abc_16259_n9382), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__29_) );
  OR2X2 OR2X2_3107 ( .A(AES_CORE_DATAPATH__abc_16259_n9386), .B(AES_CORE_DATAPATH__abc_16259_n9385), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__30_) );
  OR2X2 OR2X2_3108 ( .A(AES_CORE_DATAPATH__abc_16259_n9389), .B(AES_CORE_DATAPATH__abc_16259_n9388), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__31_) );
  OR2X2 OR2X2_3109 ( .A(AES_CORE_DATAPATH__abc_16259_n7675), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n9391) );
  OR2X2 OR2X2_311 ( .A(AES_CORE_DATAPATH__abc_16259_n3027_1), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n3028) );
  OR2X2 OR2X2_3110 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf7), .B(AES_CORE_DATAPATH_bkp_1_2__0_), .Y(AES_CORE_DATAPATH__abc_16259_n9392) );
  OR2X2 OR2X2_3111 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n8608), .Y(AES_CORE_DATAPATH__abc_16259_n9395) );
  OR2X2 OR2X2_3112 ( .A(AES_CORE_DATAPATH__abc_16259_n9394), .B(AES_CORE_DATAPATH__abc_16259_n9395), .Y(AES_CORE_DATAPATH__abc_16259_n9396) );
  OR2X2 OR2X2_3113 ( .A(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf0), .B(AES_CORE_DATAPATH_bkp_2__0_), .Y(AES_CORE_DATAPATH__abc_16259_n9397) );
  OR2X2 OR2X2_3114 ( .A(AES_CORE_DATAPATH__abc_16259_n7683), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n9399) );
  OR2X2 OR2X2_3115 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf6), .B(AES_CORE_DATAPATH_bkp_1_2__1_), .Y(AES_CORE_DATAPATH__abc_16259_n9400) );
  OR2X2 OR2X2_3116 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n8617), .Y(AES_CORE_DATAPATH__abc_16259_n9403) );
  OR2X2 OR2X2_3117 ( .A(AES_CORE_DATAPATH__abc_16259_n9402), .B(AES_CORE_DATAPATH__abc_16259_n9403), .Y(AES_CORE_DATAPATH__abc_16259_n9404) );
  OR2X2 OR2X2_3118 ( .A(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf7), .B(AES_CORE_DATAPATH_bkp_2__1_), .Y(AES_CORE_DATAPATH__abc_16259_n9405) );
  OR2X2 OR2X2_3119 ( .A(AES_CORE_DATAPATH__abc_16259_n7691), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n9407) );
  OR2X2 OR2X2_312 ( .A(AES_CORE_DATAPATH__abc_16259_n3030), .B(AES_CORE_DATAPATH__abc_16259_n3031), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_4_) );
  OR2X2 OR2X2_3120 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf5), .B(AES_CORE_DATAPATH_bkp_1_2__2_), .Y(AES_CORE_DATAPATH__abc_16259_n9408) );
  OR2X2 OR2X2_3121 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf6), .B(AES_CORE_DATAPATH__abc_16259_n8626), .Y(AES_CORE_DATAPATH__abc_16259_n9411) );
  OR2X2 OR2X2_3122 ( .A(AES_CORE_DATAPATH__abc_16259_n9410), .B(AES_CORE_DATAPATH__abc_16259_n9411), .Y(AES_CORE_DATAPATH__abc_16259_n9412) );
  OR2X2 OR2X2_3123 ( .A(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf6), .B(AES_CORE_DATAPATH_bkp_2__2_), .Y(AES_CORE_DATAPATH__abc_16259_n9413) );
  OR2X2 OR2X2_3124 ( .A(AES_CORE_DATAPATH__abc_16259_n7699), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n9415) );
  OR2X2 OR2X2_3125 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf4), .B(AES_CORE_DATAPATH_bkp_1_2__3_), .Y(AES_CORE_DATAPATH__abc_16259_n9416) );
  OR2X2 OR2X2_3126 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf5), .B(AES_CORE_DATAPATH__abc_16259_n8635), .Y(AES_CORE_DATAPATH__abc_16259_n9419) );
  OR2X2 OR2X2_3127 ( .A(AES_CORE_DATAPATH__abc_16259_n9418), .B(AES_CORE_DATAPATH__abc_16259_n9419), .Y(AES_CORE_DATAPATH__abc_16259_n9420) );
  OR2X2 OR2X2_3128 ( .A(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf5), .B(AES_CORE_DATAPATH_bkp_2__3_), .Y(AES_CORE_DATAPATH__abc_16259_n9421) );
  OR2X2 OR2X2_3129 ( .A(AES_CORE_DATAPATH__abc_16259_n7707), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf9), .Y(AES_CORE_DATAPATH__abc_16259_n9423) );
  OR2X2 OR2X2_313 ( .A(AES_CORE_DATAPATH__abc_16259_n2774_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n3033_1), .Y(AES_CORE_DATAPATH__abc_16259_n3034) );
  OR2X2 OR2X2_3130 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1_2__4_), .Y(AES_CORE_DATAPATH__abc_16259_n9424) );
  OR2X2 OR2X2_3131 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n8644), .Y(AES_CORE_DATAPATH__abc_16259_n9427) );
  OR2X2 OR2X2_3132 ( .A(AES_CORE_DATAPATH__abc_16259_n9426), .B(AES_CORE_DATAPATH__abc_16259_n9427), .Y(AES_CORE_DATAPATH__abc_16259_n9428) );
  OR2X2 OR2X2_3133 ( .A(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf4), .B(AES_CORE_DATAPATH_bkp_2__4_), .Y(AES_CORE_DATAPATH__abc_16259_n9429) );
  OR2X2 OR2X2_3134 ( .A(AES_CORE_DATAPATH__abc_16259_n7715), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf8), .Y(AES_CORE_DATAPATH__abc_16259_n9431) );
  OR2X2 OR2X2_3135 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf2), .B(AES_CORE_DATAPATH_bkp_1_2__5_), .Y(AES_CORE_DATAPATH__abc_16259_n9432) );
  OR2X2 OR2X2_3136 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n8653), .Y(AES_CORE_DATAPATH__abc_16259_n9435) );
  OR2X2 OR2X2_3137 ( .A(AES_CORE_DATAPATH__abc_16259_n9434), .B(AES_CORE_DATAPATH__abc_16259_n9435), .Y(AES_CORE_DATAPATH__abc_16259_n9436) );
  OR2X2 OR2X2_3138 ( .A(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf3), .B(AES_CORE_DATAPATH_bkp_2__5_), .Y(AES_CORE_DATAPATH__abc_16259_n9437) );
  OR2X2 OR2X2_3139 ( .A(AES_CORE_DATAPATH__abc_16259_n7723), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n9439) );
  OR2X2 OR2X2_314 ( .A(AES_CORE_DATAPATH__abc_16259_n2778_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n3035), .Y(AES_CORE_DATAPATH__abc_16259_n3036_1) );
  OR2X2 OR2X2_3140 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf1), .B(AES_CORE_DATAPATH_bkp_1_2__6_), .Y(AES_CORE_DATAPATH__abc_16259_n9440) );
  OR2X2 OR2X2_3141 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n8662), .Y(AES_CORE_DATAPATH__abc_16259_n9443) );
  OR2X2 OR2X2_3142 ( .A(AES_CORE_DATAPATH__abc_16259_n9442), .B(AES_CORE_DATAPATH__abc_16259_n9443), .Y(AES_CORE_DATAPATH__abc_16259_n9444) );
  OR2X2 OR2X2_3143 ( .A(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf2), .B(AES_CORE_DATAPATH_bkp_2__6_), .Y(AES_CORE_DATAPATH__abc_16259_n9445) );
  OR2X2 OR2X2_3144 ( .A(AES_CORE_DATAPATH__abc_16259_n7731), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n9447) );
  OR2X2 OR2X2_3145 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf0), .B(AES_CORE_DATAPATH_bkp_1_2__7_), .Y(AES_CORE_DATAPATH__abc_16259_n9448) );
  OR2X2 OR2X2_3146 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n8671), .Y(AES_CORE_DATAPATH__abc_16259_n9451) );
  OR2X2 OR2X2_3147 ( .A(AES_CORE_DATAPATH__abc_16259_n9450), .B(AES_CORE_DATAPATH__abc_16259_n9451), .Y(AES_CORE_DATAPATH__abc_16259_n9452) );
  OR2X2 OR2X2_3148 ( .A(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf1), .B(AES_CORE_DATAPATH_bkp_2__7_), .Y(AES_CORE_DATAPATH__abc_16259_n9453) );
  OR2X2 OR2X2_3149 ( .A(AES_CORE_DATAPATH__abc_16259_n7739), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n9455) );
  OR2X2 OR2X2_315 ( .A(AES_CORE_DATAPATH__abc_16259_n3039), .B(AES_CORE_DATAPATH__abc_16259_n3040_1), .Y(AES_CORE_DATAPATH__abc_16259_n3041) );
  OR2X2 OR2X2_3150 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf11), .B(AES_CORE_DATAPATH_bkp_1_2__8_), .Y(AES_CORE_DATAPATH__abc_16259_n9456) );
  OR2X2 OR2X2_3151 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n8680), .Y(AES_CORE_DATAPATH__abc_16259_n9459) );
  OR2X2 OR2X2_3152 ( .A(AES_CORE_DATAPATH__abc_16259_n9458), .B(AES_CORE_DATAPATH__abc_16259_n9459), .Y(AES_CORE_DATAPATH__abc_16259_n9460) );
  OR2X2 OR2X2_3153 ( .A(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf0), .B(AES_CORE_DATAPATH_bkp_2__8_), .Y(AES_CORE_DATAPATH__abc_16259_n9461) );
  OR2X2 OR2X2_3154 ( .A(AES_CORE_DATAPATH__abc_16259_n7747), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n9463) );
  OR2X2 OR2X2_3155 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf10), .B(AES_CORE_DATAPATH_bkp_1_2__9_), .Y(AES_CORE_DATAPATH__abc_16259_n9464) );
  OR2X2 OR2X2_3156 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf6), .B(AES_CORE_DATAPATH__abc_16259_n8689), .Y(AES_CORE_DATAPATH__abc_16259_n9467) );
  OR2X2 OR2X2_3157 ( .A(AES_CORE_DATAPATH__abc_16259_n9466), .B(AES_CORE_DATAPATH__abc_16259_n9467), .Y(AES_CORE_DATAPATH__abc_16259_n9468) );
  OR2X2 OR2X2_3158 ( .A(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf7), .B(AES_CORE_DATAPATH_bkp_2__9_), .Y(AES_CORE_DATAPATH__abc_16259_n9469) );
  OR2X2 OR2X2_3159 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf8), .B(AES_CORE_DATAPATH_bkp_1_2__10_), .Y(AES_CORE_DATAPATH__abc_16259_n9473) );
  OR2X2 OR2X2_316 ( .A(AES_CORE_DATAPATH__abc_16259_n3041), .B(AES_CORE_DATAPATH__abc_16259_n3038_1), .Y(AES_CORE_DATAPATH__abc_16259_n3042_1) );
  OR2X2 OR2X2_3160 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf5), .B(AES_CORE_DATAPATH__abc_16259_n8699), .Y(AES_CORE_DATAPATH__abc_16259_n9476) );
  OR2X2 OR2X2_3161 ( .A(AES_CORE_DATAPATH__abc_16259_n9475), .B(AES_CORE_DATAPATH__abc_16259_n9476), .Y(AES_CORE_DATAPATH__abc_16259_n9477) );
  OR2X2 OR2X2_3162 ( .A(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf6), .B(AES_CORE_DATAPATH_bkp_2__10_), .Y(AES_CORE_DATAPATH__abc_16259_n9478) );
  OR2X2 OR2X2_3163 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf6), .B(AES_CORE_DATAPATH_bkp_1_2__11_), .Y(AES_CORE_DATAPATH__abc_16259_n9482) );
  OR2X2 OR2X2_3164 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n8709), .Y(AES_CORE_DATAPATH__abc_16259_n9485) );
  OR2X2 OR2X2_3165 ( .A(AES_CORE_DATAPATH__abc_16259_n9484), .B(AES_CORE_DATAPATH__abc_16259_n9485), .Y(AES_CORE_DATAPATH__abc_16259_n9486) );
  OR2X2 OR2X2_3166 ( .A(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf5), .B(AES_CORE_DATAPATH_bkp_2__11_), .Y(AES_CORE_DATAPATH__abc_16259_n9487) );
  OR2X2 OR2X2_3167 ( .A(AES_CORE_DATAPATH__abc_16259_n7777), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n9489) );
  OR2X2 OR2X2_3168 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf5), .B(AES_CORE_DATAPATH_bkp_1_2__12_), .Y(AES_CORE_DATAPATH__abc_16259_n9490) );
  OR2X2 OR2X2_3169 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n8718), .Y(AES_CORE_DATAPATH__abc_16259_n9493) );
  OR2X2 OR2X2_317 ( .A(AES_CORE_DATAPATH__abc_16259_n3046), .B(AES_CORE_DATAPATH__abc_16259_n2826_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n3047) );
  OR2X2 OR2X2_3170 ( .A(AES_CORE_DATAPATH__abc_16259_n9492), .B(AES_CORE_DATAPATH__abc_16259_n9493), .Y(AES_CORE_DATAPATH__abc_16259_n9494) );
  OR2X2 OR2X2_3171 ( .A(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf4), .B(AES_CORE_DATAPATH_bkp_2__12_), .Y(AES_CORE_DATAPATH__abc_16259_n9495) );
  OR2X2 OR2X2_3172 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1_2__13_), .Y(AES_CORE_DATAPATH__abc_16259_n9499) );
  OR2X2 OR2X2_3173 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n8728), .Y(AES_CORE_DATAPATH__abc_16259_n9502) );
  OR2X2 OR2X2_3174 ( .A(AES_CORE_DATAPATH__abc_16259_n9501), .B(AES_CORE_DATAPATH__abc_16259_n9502), .Y(AES_CORE_DATAPATH__abc_16259_n9503) );
  OR2X2 OR2X2_3175 ( .A(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf3), .B(AES_CORE_DATAPATH_bkp_2__13_), .Y(AES_CORE_DATAPATH__abc_16259_n9504) );
  OR2X2 OR2X2_3176 ( .A(AES_CORE_DATAPATH__abc_16259_n7796), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n9506) );
  OR2X2 OR2X2_3177 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf2), .B(AES_CORE_DATAPATH_bkp_1_2__14_), .Y(AES_CORE_DATAPATH__abc_16259_n9507) );
  OR2X2 OR2X2_3178 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n8737), .Y(AES_CORE_DATAPATH__abc_16259_n9510) );
  OR2X2 OR2X2_3179 ( .A(AES_CORE_DATAPATH__abc_16259_n9509), .B(AES_CORE_DATAPATH__abc_16259_n9510), .Y(AES_CORE_DATAPATH__abc_16259_n9511) );
  OR2X2 OR2X2_318 ( .A(AES_CORE_DATAPATH__abc_16259_n3048), .B(AES_CORE_DATAPATH__abc_16259_n3049), .Y(AES_CORE_DATAPATH__abc_16259_n3050) );
  OR2X2 OR2X2_3180 ( .A(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf2), .B(AES_CORE_DATAPATH_bkp_2__14_), .Y(AES_CORE_DATAPATH__abc_16259_n9512) );
  OR2X2 OR2X2_3181 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf0), .B(AES_CORE_DATAPATH_bkp_1_2__15_), .Y(AES_CORE_DATAPATH__abc_16259_n9516) );
  OR2X2 OR2X2_3182 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n8747), .Y(AES_CORE_DATAPATH__abc_16259_n9519) );
  OR2X2 OR2X2_3183 ( .A(AES_CORE_DATAPATH__abc_16259_n9518), .B(AES_CORE_DATAPATH__abc_16259_n9519), .Y(AES_CORE_DATAPATH__abc_16259_n9520) );
  OR2X2 OR2X2_3184 ( .A(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf1), .B(AES_CORE_DATAPATH_bkp_2__15_), .Y(AES_CORE_DATAPATH__abc_16259_n9521) );
  OR2X2 OR2X2_3185 ( .A(AES_CORE_DATAPATH__abc_16259_n7815), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n9523) );
  OR2X2 OR2X2_3186 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf11), .B(AES_CORE_DATAPATH_bkp_1_2__16_), .Y(AES_CORE_DATAPATH__abc_16259_n9524) );
  OR2X2 OR2X2_3187 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf6), .B(AES_CORE_DATAPATH__abc_16259_n8756), .Y(AES_CORE_DATAPATH__abc_16259_n9527) );
  OR2X2 OR2X2_3188 ( .A(AES_CORE_DATAPATH__abc_16259_n9526), .B(AES_CORE_DATAPATH__abc_16259_n9527), .Y(AES_CORE_DATAPATH__abc_16259_n9528) );
  OR2X2 OR2X2_3189 ( .A(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf0), .B(AES_CORE_DATAPATH_bkp_2__16_), .Y(AES_CORE_DATAPATH__abc_16259_n9529) );
  OR2X2 OR2X2_319 ( .A(AES_CORE_DATAPATH__abc_16259_n3050), .B(AES_CORE_DATAPATH__abc_16259_n3047), .Y(AES_CORE_DATAPATH__abc_16259_n3051) );
  OR2X2 OR2X2_3190 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf9), .B(AES_CORE_DATAPATH_bkp_1_2__17_), .Y(AES_CORE_DATAPATH__abc_16259_n9533) );
  OR2X2 OR2X2_3191 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf5), .B(AES_CORE_DATAPATH__abc_16259_n8766), .Y(AES_CORE_DATAPATH__abc_16259_n9536) );
  OR2X2 OR2X2_3192 ( .A(AES_CORE_DATAPATH__abc_16259_n9535), .B(AES_CORE_DATAPATH__abc_16259_n9536), .Y(AES_CORE_DATAPATH__abc_16259_n9537) );
  OR2X2 OR2X2_3193 ( .A(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf7), .B(AES_CORE_DATAPATH_bkp_2__17_), .Y(AES_CORE_DATAPATH__abc_16259_n9538) );
  OR2X2 OR2X2_3194 ( .A(AES_CORE_DATAPATH__abc_16259_n7834), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n9540) );
  OR2X2 OR2X2_3195 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf8), .B(AES_CORE_DATAPATH_bkp_1_2__18_), .Y(AES_CORE_DATAPATH__abc_16259_n9541) );
  OR2X2 OR2X2_3196 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n8775), .Y(AES_CORE_DATAPATH__abc_16259_n9544) );
  OR2X2 OR2X2_3197 ( .A(AES_CORE_DATAPATH__abc_16259_n9543), .B(AES_CORE_DATAPATH__abc_16259_n9544), .Y(AES_CORE_DATAPATH__abc_16259_n9545) );
  OR2X2 OR2X2_3198 ( .A(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf6), .B(AES_CORE_DATAPATH_bkp_2__18_), .Y(AES_CORE_DATAPATH__abc_16259_n9546) );
  OR2X2 OR2X2_3199 ( .A(AES_CORE_DATAPATH__abc_16259_n7842), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf9), .Y(AES_CORE_DATAPATH__abc_16259_n9548) );
  OR2X2 OR2X2_32 ( .A(AES_CORE_CONTROL_UNIT_state_13_), .B(AES_CORE_CONTROL_UNIT_key_gen), .Y(AES_CORE_CONTROL_UNIT_sbox_sel_2_) );
  OR2X2 OR2X2_320 ( .A(AES_CORE_DATAPATH__abc_16259_n2841_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__5_), .Y(AES_CORE_DATAPATH__abc_16259_n3052) );
  OR2X2 OR2X2_3200 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf7), .B(AES_CORE_DATAPATH_bkp_1_2__19_), .Y(AES_CORE_DATAPATH__abc_16259_n9549) );
  OR2X2 OR2X2_3201 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n8784), .Y(AES_CORE_DATAPATH__abc_16259_n9552) );
  OR2X2 OR2X2_3202 ( .A(AES_CORE_DATAPATH__abc_16259_n9551), .B(AES_CORE_DATAPATH__abc_16259_n9552), .Y(AES_CORE_DATAPATH__abc_16259_n9553) );
  OR2X2 OR2X2_3203 ( .A(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf5), .B(AES_CORE_DATAPATH_bkp_2__19_), .Y(AES_CORE_DATAPATH__abc_16259_n9554) );
  OR2X2 OR2X2_3204 ( .A(AES_CORE_DATAPATH__abc_16259_n7850), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf8), .Y(AES_CORE_DATAPATH__abc_16259_n9556) );
  OR2X2 OR2X2_3205 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf6), .B(AES_CORE_DATAPATH_bkp_1_2__20_), .Y(AES_CORE_DATAPATH__abc_16259_n9557) );
  OR2X2 OR2X2_3206 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n8793), .Y(AES_CORE_DATAPATH__abc_16259_n9560) );
  OR2X2 OR2X2_3207 ( .A(AES_CORE_DATAPATH__abc_16259_n9559), .B(AES_CORE_DATAPATH__abc_16259_n9560), .Y(AES_CORE_DATAPATH__abc_16259_n9561) );
  OR2X2 OR2X2_3208 ( .A(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf4), .B(AES_CORE_DATAPATH_bkp_2__20_), .Y(AES_CORE_DATAPATH__abc_16259_n9562) );
  OR2X2 OR2X2_3209 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf4), .B(AES_CORE_DATAPATH_bkp_1_2__21_), .Y(AES_CORE_DATAPATH__abc_16259_n9566) );
  OR2X2 OR2X2_321 ( .A(AES_CORE_DATAPATH__abc_16259_n3044), .B(AES_CORE_DATAPATH__abc_16259_n2853_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n3054_1) );
  OR2X2 OR2X2_3210 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n8803), .Y(AES_CORE_DATAPATH__abc_16259_n9569) );
  OR2X2 OR2X2_3211 ( .A(AES_CORE_DATAPATH__abc_16259_n9568), .B(AES_CORE_DATAPATH__abc_16259_n9569), .Y(AES_CORE_DATAPATH__abc_16259_n9570) );
  OR2X2 OR2X2_3212 ( .A(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf3), .B(AES_CORE_DATAPATH_bkp_2__21_), .Y(AES_CORE_DATAPATH__abc_16259_n9571) );
  OR2X2 OR2X2_3213 ( .A(AES_CORE_DATAPATH__abc_16259_n7869), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n9573) );
  OR2X2 OR2X2_3214 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1_2__22_), .Y(AES_CORE_DATAPATH__abc_16259_n9574) );
  OR2X2 OR2X2_3215 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n8812), .Y(AES_CORE_DATAPATH__abc_16259_n9577) );
  OR2X2 OR2X2_3216 ( .A(AES_CORE_DATAPATH__abc_16259_n9576), .B(AES_CORE_DATAPATH__abc_16259_n9577), .Y(AES_CORE_DATAPATH__abc_16259_n9578) );
  OR2X2 OR2X2_3217 ( .A(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf2), .B(AES_CORE_DATAPATH_bkp_2__22_), .Y(AES_CORE_DATAPATH__abc_16259_n9579) );
  OR2X2 OR2X2_3218 ( .A(AES_CORE_DATAPATH__abc_16259_n7877), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n9581) );
  OR2X2 OR2X2_3219 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf2), .B(AES_CORE_DATAPATH_bkp_1_2__23_), .Y(AES_CORE_DATAPATH__abc_16259_n9582) );
  OR2X2 OR2X2_322 ( .A(AES_CORE_DATAPATH__abc_16259_n3055), .B(AES_CORE_DATAPATH__abc_16259_n3056_1), .Y(AES_CORE_DATAPATH__abc_16259_n3057) );
  OR2X2 OR2X2_3220 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf6), .B(AES_CORE_DATAPATH__abc_16259_n8821), .Y(AES_CORE_DATAPATH__abc_16259_n9585) );
  OR2X2 OR2X2_3221 ( .A(AES_CORE_DATAPATH__abc_16259_n9584), .B(AES_CORE_DATAPATH__abc_16259_n9585), .Y(AES_CORE_DATAPATH__abc_16259_n9586) );
  OR2X2 OR2X2_3222 ( .A(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf1), .B(AES_CORE_DATAPATH_bkp_2__23_), .Y(AES_CORE_DATAPATH__abc_16259_n9587) );
  OR2X2 OR2X2_3223 ( .A(AES_CORE_DATAPATH__abc_16259_n7885), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n9589) );
  OR2X2 OR2X2_3224 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf1), .B(AES_CORE_DATAPATH_bkp_1_2__24_), .Y(AES_CORE_DATAPATH__abc_16259_n9590) );
  OR2X2 OR2X2_3225 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf5), .B(AES_CORE_DATAPATH__abc_16259_n8830), .Y(AES_CORE_DATAPATH__abc_16259_n9593) );
  OR2X2 OR2X2_3226 ( .A(AES_CORE_DATAPATH__abc_16259_n9592), .B(AES_CORE_DATAPATH__abc_16259_n9593), .Y(AES_CORE_DATAPATH__abc_16259_n9594) );
  OR2X2 OR2X2_3227 ( .A(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf0), .B(AES_CORE_DATAPATH_bkp_2__24_), .Y(AES_CORE_DATAPATH__abc_16259_n9595) );
  OR2X2 OR2X2_3228 ( .A(AES_CORE_DATAPATH__abc_16259_n7893), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n9597) );
  OR2X2 OR2X2_3229 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf0), .B(AES_CORE_DATAPATH_bkp_1_2__25_), .Y(AES_CORE_DATAPATH__abc_16259_n9598) );
  OR2X2 OR2X2_323 ( .A(_auto_iopadmap_cc_313_execute_26949_5_), .B(AES_CORE_DATAPATH__abc_16259_n3059), .Y(AES_CORE_DATAPATH__abc_16259_n3060) );
  OR2X2 OR2X2_3230 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n8839), .Y(AES_CORE_DATAPATH__abc_16259_n9601) );
  OR2X2 OR2X2_3231 ( .A(AES_CORE_DATAPATH__abc_16259_n9600), .B(AES_CORE_DATAPATH__abc_16259_n9601), .Y(AES_CORE_DATAPATH__abc_16259_n9602) );
  OR2X2 OR2X2_3232 ( .A(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf7), .B(AES_CORE_DATAPATH_bkp_2__25_), .Y(AES_CORE_DATAPATH__abc_16259_n9603) );
  OR2X2 OR2X2_3233 ( .A(AES_CORE_DATAPATH__abc_16259_n7901), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n9605) );
  OR2X2 OR2X2_3234 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf11), .B(AES_CORE_DATAPATH_bkp_1_2__26_), .Y(AES_CORE_DATAPATH__abc_16259_n9606) );
  OR2X2 OR2X2_3235 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n8848), .Y(AES_CORE_DATAPATH__abc_16259_n9609) );
  OR2X2 OR2X2_3236 ( .A(AES_CORE_DATAPATH__abc_16259_n9608), .B(AES_CORE_DATAPATH__abc_16259_n9609), .Y(AES_CORE_DATAPATH__abc_16259_n9610) );
  OR2X2 OR2X2_3237 ( .A(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf6), .B(AES_CORE_DATAPATH_bkp_2__26_), .Y(AES_CORE_DATAPATH__abc_16259_n9611) );
  OR2X2 OR2X2_3238 ( .A(AES_CORE_DATAPATH__abc_16259_n7909), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n9613) );
  OR2X2 OR2X2_3239 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf10), .B(AES_CORE_DATAPATH_bkp_1_2__27_), .Y(AES_CORE_DATAPATH__abc_16259_n9614) );
  OR2X2 OR2X2_324 ( .A(AES_CORE_DATAPATH__abc_16259_n3062_1), .B(AES_CORE_DATAPATH__abc_16259_n2864_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n3063) );
  OR2X2 OR2X2_3240 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n8857), .Y(AES_CORE_DATAPATH__abc_16259_n9617) );
  OR2X2 OR2X2_3241 ( .A(AES_CORE_DATAPATH__abc_16259_n9616), .B(AES_CORE_DATAPATH__abc_16259_n9617), .Y(AES_CORE_DATAPATH__abc_16259_n9618) );
  OR2X2 OR2X2_3242 ( .A(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf5), .B(AES_CORE_DATAPATH_bkp_2__27_), .Y(AES_CORE_DATAPATH__abc_16259_n9619) );
  OR2X2 OR2X2_3243 ( .A(AES_CORE_DATAPATH__abc_16259_n7917), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n9621) );
  OR2X2 OR2X2_3244 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf9), .B(AES_CORE_DATAPATH_bkp_1_2__28_), .Y(AES_CORE_DATAPATH__abc_16259_n9622) );
  OR2X2 OR2X2_3245 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n8866), .Y(AES_CORE_DATAPATH__abc_16259_n9625) );
  OR2X2 OR2X2_3246 ( .A(AES_CORE_DATAPATH__abc_16259_n9624), .B(AES_CORE_DATAPATH__abc_16259_n9625), .Y(AES_CORE_DATAPATH__abc_16259_n9626) );
  OR2X2 OR2X2_3247 ( .A(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf4), .B(AES_CORE_DATAPATH_bkp_2__28_), .Y(AES_CORE_DATAPATH__abc_16259_n9627) );
  OR2X2 OR2X2_3248 ( .A(AES_CORE_DATAPATH__abc_16259_n7925), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n9629) );
  OR2X2 OR2X2_3249 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf8), .B(AES_CORE_DATAPATH_bkp_1_2__29_), .Y(AES_CORE_DATAPATH__abc_16259_n9630) );
  OR2X2 OR2X2_325 ( .A(AES_CORE_DATAPATH__abc_16259_n3063), .B(AES_CORE_DATAPATH__abc_16259_n3061_1), .Y(AES_CORE_DATAPATH__abc_16259_n3064) );
  OR2X2 OR2X2_3250 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n8875), .Y(AES_CORE_DATAPATH__abc_16259_n9633) );
  OR2X2 OR2X2_3251 ( .A(AES_CORE_DATAPATH__abc_16259_n9632), .B(AES_CORE_DATAPATH__abc_16259_n9633), .Y(AES_CORE_DATAPATH__abc_16259_n9634) );
  OR2X2 OR2X2_3252 ( .A(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf3), .B(AES_CORE_DATAPATH_bkp_2__29_), .Y(AES_CORE_DATAPATH__abc_16259_n9635) );
  OR2X2 OR2X2_3253 ( .A(AES_CORE_DATAPATH__abc_16259_n7933), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf9), .Y(AES_CORE_DATAPATH__abc_16259_n9637) );
  OR2X2 OR2X2_3254 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf7), .B(AES_CORE_DATAPATH_bkp_1_2__30_), .Y(AES_CORE_DATAPATH__abc_16259_n9638) );
  OR2X2 OR2X2_3255 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf6), .B(AES_CORE_DATAPATH__abc_16259_n8884), .Y(AES_CORE_DATAPATH__abc_16259_n9641) );
  OR2X2 OR2X2_3256 ( .A(AES_CORE_DATAPATH__abc_16259_n9640), .B(AES_CORE_DATAPATH__abc_16259_n9641), .Y(AES_CORE_DATAPATH__abc_16259_n9642) );
  OR2X2 OR2X2_3257 ( .A(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf2), .B(AES_CORE_DATAPATH_bkp_2__30_), .Y(AES_CORE_DATAPATH__abc_16259_n9643) );
  OR2X2 OR2X2_3258 ( .A(AES_CORE_DATAPATH__abc_16259_n7941), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf8), .Y(AES_CORE_DATAPATH__abc_16259_n9645) );
  OR2X2 OR2X2_3259 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf6), .B(AES_CORE_DATAPATH_bkp_1_2__31_), .Y(AES_CORE_DATAPATH__abc_16259_n9646) );
  OR2X2 OR2X2_326 ( .A(AES_CORE_DATAPATH__abc_16259_n3066), .B(AES_CORE_DATAPATH__abc_16259_n3065_1), .Y(AES_CORE_DATAPATH__abc_16259_n3067_1) );
  OR2X2 OR2X2_3260 ( .A(AES_CORE_DATAPATH__abc_16259_n9288_bF_buf5), .B(AES_CORE_DATAPATH__abc_16259_n8893), .Y(AES_CORE_DATAPATH__abc_16259_n9649) );
  OR2X2 OR2X2_3261 ( .A(AES_CORE_DATAPATH__abc_16259_n9648), .B(AES_CORE_DATAPATH__abc_16259_n9649), .Y(AES_CORE_DATAPATH__abc_16259_n9650) );
  OR2X2 OR2X2_3262 ( .A(AES_CORE_DATAPATH__abc_16259_n9287_bF_buf1), .B(AES_CORE_DATAPATH_bkp_2__31_), .Y(AES_CORE_DATAPATH__abc_16259_n9651) );
  OR2X2 OR2X2_3263 ( .A(AES_CORE_DATAPATH_iv_2__0_), .B(iv_en_2_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n9653) );
  OR2X2 OR2X2_3264 ( .A(AES_CORE_DATAPATH__abc_16259_n9654_bF_buf4), .B(\bus_in[0] ), .Y(AES_CORE_DATAPATH__abc_16259_n9655) );
  OR2X2 OR2X2_3265 ( .A(AES_CORE_DATAPATH_iv_2__1_), .B(iv_en_2_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n9657) );
  OR2X2 OR2X2_3266 ( .A(AES_CORE_DATAPATH__abc_16259_n9654_bF_buf3), .B(\bus_in[1] ), .Y(AES_CORE_DATAPATH__abc_16259_n9658) );
  OR2X2 OR2X2_3267 ( .A(AES_CORE_DATAPATH_iv_2__2_), .B(iv_en_2_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n9660) );
  OR2X2 OR2X2_3268 ( .A(AES_CORE_DATAPATH__abc_16259_n9654_bF_buf2), .B(\bus_in[2] ), .Y(AES_CORE_DATAPATH__abc_16259_n9661) );
  OR2X2 OR2X2_3269 ( .A(AES_CORE_DATAPATH_iv_2__3_), .B(iv_en_2_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n9663) );
  OR2X2 OR2X2_327 ( .A(AES_CORE_DATAPATH__abc_16259_n3067_1), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n3068) );
  OR2X2 OR2X2_3270 ( .A(AES_CORE_DATAPATH__abc_16259_n9654_bF_buf1), .B(\bus_in[3] ), .Y(AES_CORE_DATAPATH__abc_16259_n9664) );
  OR2X2 OR2X2_3271 ( .A(AES_CORE_DATAPATH_iv_2__4_), .B(iv_en_2_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n9666) );
  OR2X2 OR2X2_3272 ( .A(AES_CORE_DATAPATH__abc_16259_n9654_bF_buf0), .B(\bus_in[4] ), .Y(AES_CORE_DATAPATH__abc_16259_n9667) );
  OR2X2 OR2X2_3273 ( .A(AES_CORE_DATAPATH_iv_2__5_), .B(iv_en_2_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n9669) );
  OR2X2 OR2X2_3274 ( .A(AES_CORE_DATAPATH__abc_16259_n9654_bF_buf4), .B(\bus_in[5] ), .Y(AES_CORE_DATAPATH__abc_16259_n9670) );
  OR2X2 OR2X2_3275 ( .A(AES_CORE_DATAPATH_iv_2__6_), .B(iv_en_2_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n9672) );
  OR2X2 OR2X2_3276 ( .A(AES_CORE_DATAPATH__abc_16259_n9654_bF_buf3), .B(\bus_in[6] ), .Y(AES_CORE_DATAPATH__abc_16259_n9673) );
  OR2X2 OR2X2_3277 ( .A(AES_CORE_DATAPATH_iv_2__7_), .B(iv_en_2_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n9675) );
  OR2X2 OR2X2_3278 ( .A(AES_CORE_DATAPATH__abc_16259_n9654_bF_buf2), .B(\bus_in[7] ), .Y(AES_CORE_DATAPATH__abc_16259_n9676) );
  OR2X2 OR2X2_3279 ( .A(AES_CORE_DATAPATH_iv_2__8_), .B(iv_en_2_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n9678) );
  OR2X2 OR2X2_328 ( .A(AES_CORE_DATAPATH__abc_16259_n3070), .B(AES_CORE_DATAPATH__abc_16259_n3071_1), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_5_) );
  OR2X2 OR2X2_3280 ( .A(AES_CORE_DATAPATH__abc_16259_n9654_bF_buf1), .B(\bus_in[8] ), .Y(AES_CORE_DATAPATH__abc_16259_n9679) );
  OR2X2 OR2X2_3281 ( .A(AES_CORE_DATAPATH_iv_2__9_), .B(iv_en_2_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n9681) );
  OR2X2 OR2X2_3282 ( .A(AES_CORE_DATAPATH__abc_16259_n9654_bF_buf0), .B(\bus_in[9] ), .Y(AES_CORE_DATAPATH__abc_16259_n9682) );
  OR2X2 OR2X2_3283 ( .A(AES_CORE_DATAPATH_iv_2__10_), .B(iv_en_2_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n9684) );
  OR2X2 OR2X2_3284 ( .A(AES_CORE_DATAPATH__abc_16259_n9654_bF_buf4), .B(\bus_in[10] ), .Y(AES_CORE_DATAPATH__abc_16259_n9685) );
  OR2X2 OR2X2_3285 ( .A(AES_CORE_DATAPATH_iv_2__11_), .B(iv_en_2_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n9687) );
  OR2X2 OR2X2_3286 ( .A(AES_CORE_DATAPATH__abc_16259_n9654_bF_buf3), .B(\bus_in[11] ), .Y(AES_CORE_DATAPATH__abc_16259_n9688) );
  OR2X2 OR2X2_3287 ( .A(AES_CORE_DATAPATH_iv_2__12_), .B(iv_en_2_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n9690) );
  OR2X2 OR2X2_3288 ( .A(AES_CORE_DATAPATH__abc_16259_n9654_bF_buf2), .B(\bus_in[12] ), .Y(AES_CORE_DATAPATH__abc_16259_n9691) );
  OR2X2 OR2X2_3289 ( .A(AES_CORE_DATAPATH_iv_2__13_), .B(iv_en_2_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n9693) );
  OR2X2 OR2X2_329 ( .A(AES_CORE_DATAPATH__abc_16259_n2774_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n3073), .Y(AES_CORE_DATAPATH__abc_16259_n3074) );
  OR2X2 OR2X2_3290 ( .A(AES_CORE_DATAPATH__abc_16259_n9654_bF_buf1), .B(\bus_in[13] ), .Y(AES_CORE_DATAPATH__abc_16259_n9694) );
  OR2X2 OR2X2_3291 ( .A(AES_CORE_DATAPATH_iv_2__14_), .B(iv_en_2_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n9696) );
  OR2X2 OR2X2_3292 ( .A(AES_CORE_DATAPATH__abc_16259_n9654_bF_buf0), .B(\bus_in[14] ), .Y(AES_CORE_DATAPATH__abc_16259_n9697) );
  OR2X2 OR2X2_3293 ( .A(AES_CORE_DATAPATH_iv_2__15_), .B(iv_en_2_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n9699) );
  OR2X2 OR2X2_3294 ( .A(AES_CORE_DATAPATH__abc_16259_n9654_bF_buf4), .B(\bus_in[15] ), .Y(AES_CORE_DATAPATH__abc_16259_n9700) );
  OR2X2 OR2X2_3295 ( .A(AES_CORE_DATAPATH_iv_2__16_), .B(iv_en_2_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n9702) );
  OR2X2 OR2X2_3296 ( .A(AES_CORE_DATAPATH__abc_16259_n9654_bF_buf3), .B(\bus_in[16] ), .Y(AES_CORE_DATAPATH__abc_16259_n9703) );
  OR2X2 OR2X2_3297 ( .A(AES_CORE_DATAPATH_iv_2__17_), .B(iv_en_2_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n9705) );
  OR2X2 OR2X2_3298 ( .A(AES_CORE_DATAPATH__abc_16259_n9654_bF_buf2), .B(\bus_in[17] ), .Y(AES_CORE_DATAPATH__abc_16259_n9706) );
  OR2X2 OR2X2_3299 ( .A(AES_CORE_DATAPATH_iv_2__18_), .B(iv_en_2_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n9708) );
  OR2X2 OR2X2_33 ( .A(AES_CORE_CONTROL_UNIT_sbox_sel_2_), .B(AES_CORE_CONTROL_UNIT_rd_count_0_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n168) );
  OR2X2 OR2X2_330 ( .A(AES_CORE_DATAPATH__abc_16259_n2778_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n3075), .Y(AES_CORE_DATAPATH__abc_16259_n3076) );
  OR2X2 OR2X2_3300 ( .A(AES_CORE_DATAPATH__abc_16259_n9654_bF_buf1), .B(\bus_in[18] ), .Y(AES_CORE_DATAPATH__abc_16259_n9709) );
  OR2X2 OR2X2_3301 ( .A(AES_CORE_DATAPATH_iv_2__19_), .B(iv_en_2_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n9711) );
  OR2X2 OR2X2_3302 ( .A(AES_CORE_DATAPATH__abc_16259_n9654_bF_buf0), .B(\bus_in[19] ), .Y(AES_CORE_DATAPATH__abc_16259_n9712) );
  OR2X2 OR2X2_3303 ( .A(AES_CORE_DATAPATH_iv_2__20_), .B(iv_en_2_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n9714) );
  OR2X2 OR2X2_3304 ( .A(AES_CORE_DATAPATH__abc_16259_n9654_bF_buf4), .B(\bus_in[20] ), .Y(AES_CORE_DATAPATH__abc_16259_n9715) );
  OR2X2 OR2X2_3305 ( .A(AES_CORE_DATAPATH_iv_2__21_), .B(iv_en_2_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n9717) );
  OR2X2 OR2X2_3306 ( .A(AES_CORE_DATAPATH__abc_16259_n9654_bF_buf3), .B(\bus_in[21] ), .Y(AES_CORE_DATAPATH__abc_16259_n9718) );
  OR2X2 OR2X2_3307 ( .A(AES_CORE_DATAPATH_iv_2__22_), .B(iv_en_2_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n9720) );
  OR2X2 OR2X2_3308 ( .A(AES_CORE_DATAPATH__abc_16259_n9654_bF_buf2), .B(\bus_in[22] ), .Y(AES_CORE_DATAPATH__abc_16259_n9721) );
  OR2X2 OR2X2_3309 ( .A(AES_CORE_DATAPATH_iv_2__23_), .B(iv_en_2_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n9723) );
  OR2X2 OR2X2_331 ( .A(AES_CORE_DATAPATH__abc_16259_n3079), .B(AES_CORE_DATAPATH__abc_16259_n3080), .Y(AES_CORE_DATAPATH__abc_16259_n3081) );
  OR2X2 OR2X2_3310 ( .A(AES_CORE_DATAPATH__abc_16259_n9654_bF_buf1), .B(\bus_in[23] ), .Y(AES_CORE_DATAPATH__abc_16259_n9724) );
  OR2X2 OR2X2_3311 ( .A(AES_CORE_DATAPATH_iv_2__24_), .B(iv_en_2_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n9726) );
  OR2X2 OR2X2_3312 ( .A(AES_CORE_DATAPATH__abc_16259_n9654_bF_buf0), .B(\bus_in[24] ), .Y(AES_CORE_DATAPATH__abc_16259_n9727) );
  OR2X2 OR2X2_3313 ( .A(AES_CORE_DATAPATH_iv_2__25_), .B(iv_en_2_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n9729) );
  OR2X2 OR2X2_3314 ( .A(AES_CORE_DATAPATH__abc_16259_n9654_bF_buf4), .B(\bus_in[25] ), .Y(AES_CORE_DATAPATH__abc_16259_n9730) );
  OR2X2 OR2X2_3315 ( .A(AES_CORE_DATAPATH_iv_2__26_), .B(iv_en_2_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n9732) );
  OR2X2 OR2X2_3316 ( .A(AES_CORE_DATAPATH__abc_16259_n9654_bF_buf3), .B(\bus_in[26] ), .Y(AES_CORE_DATAPATH__abc_16259_n9733) );
  OR2X2 OR2X2_3317 ( .A(AES_CORE_DATAPATH_iv_2__27_), .B(iv_en_2_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n9735) );
  OR2X2 OR2X2_3318 ( .A(AES_CORE_DATAPATH__abc_16259_n9654_bF_buf2), .B(\bus_in[27] ), .Y(AES_CORE_DATAPATH__abc_16259_n9736) );
  OR2X2 OR2X2_3319 ( .A(AES_CORE_DATAPATH_iv_2__28_), .B(iv_en_2_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n9738) );
  OR2X2 OR2X2_332 ( .A(AES_CORE_DATAPATH__abc_16259_n3081), .B(AES_CORE_DATAPATH__abc_16259_n3078), .Y(AES_CORE_DATAPATH__abc_16259_n3082) );
  OR2X2 OR2X2_3320 ( .A(AES_CORE_DATAPATH__abc_16259_n9654_bF_buf1), .B(\bus_in[28] ), .Y(AES_CORE_DATAPATH__abc_16259_n9739) );
  OR2X2 OR2X2_3321 ( .A(AES_CORE_DATAPATH_iv_2__29_), .B(iv_en_2_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n9741) );
  OR2X2 OR2X2_3322 ( .A(AES_CORE_DATAPATH__abc_16259_n9654_bF_buf0), .B(\bus_in[29] ), .Y(AES_CORE_DATAPATH__abc_16259_n9742) );
  OR2X2 OR2X2_3323 ( .A(AES_CORE_DATAPATH_iv_2__30_), .B(iv_en_2_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n9744) );
  OR2X2 OR2X2_3324 ( .A(AES_CORE_DATAPATH__abc_16259_n9654_bF_buf4), .B(\bus_in[30] ), .Y(AES_CORE_DATAPATH__abc_16259_n9745) );
  OR2X2 OR2X2_3325 ( .A(AES_CORE_DATAPATH_iv_2__31_), .B(iv_en_2_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n9747) );
  OR2X2 OR2X2_3326 ( .A(AES_CORE_DATAPATH__abc_16259_n9654_bF_buf3), .B(\bus_in[31] ), .Y(AES_CORE_DATAPATH__abc_16259_n9748) );
  OR2X2 OR2X2_3327 ( .A(AES_CORE_DATAPATH__abc_16259_n9750), .B(AES_CORE_DATAPATH__abc_16259_n9751), .Y(AES_CORE_DATAPATH__abc_16259_n9752) );
  OR2X2 OR2X2_3328 ( .A(AES_CORE_DATAPATH__abc_16259_n9755), .B(AES_CORE_DATAPATH__abc_16259_n9754), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__0_) );
  OR2X2 OR2X2_3329 ( .A(AES_CORE_DATAPATH__abc_16259_n9758), .B(AES_CORE_DATAPATH__abc_16259_n9757), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__1_) );
  OR2X2 OR2X2_333 ( .A(AES_CORE_DATAPATH__abc_16259_n3086), .B(AES_CORE_DATAPATH__abc_16259_n2826_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n3087) );
  OR2X2 OR2X2_3330 ( .A(AES_CORE_DATAPATH__abc_16259_n9761), .B(AES_CORE_DATAPATH__abc_16259_n9760), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__2_) );
  OR2X2 OR2X2_3331 ( .A(AES_CORE_DATAPATH__abc_16259_n9764), .B(AES_CORE_DATAPATH__abc_16259_n9763), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__3_) );
  OR2X2 OR2X2_3332 ( .A(AES_CORE_DATAPATH__abc_16259_n9767), .B(AES_CORE_DATAPATH__abc_16259_n9766), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__4_) );
  OR2X2 OR2X2_3333 ( .A(AES_CORE_DATAPATH__abc_16259_n9770), .B(AES_CORE_DATAPATH__abc_16259_n9769), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__5_) );
  OR2X2 OR2X2_3334 ( .A(AES_CORE_DATAPATH__abc_16259_n9773), .B(AES_CORE_DATAPATH__abc_16259_n9772), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__6_) );
  OR2X2 OR2X2_3335 ( .A(AES_CORE_DATAPATH__abc_16259_n9776), .B(AES_CORE_DATAPATH__abc_16259_n9775), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__7_) );
  OR2X2 OR2X2_3336 ( .A(AES_CORE_DATAPATH__abc_16259_n9779), .B(AES_CORE_DATAPATH__abc_16259_n9778), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__8_) );
  OR2X2 OR2X2_3337 ( .A(AES_CORE_DATAPATH__abc_16259_n9782), .B(AES_CORE_DATAPATH__abc_16259_n9781), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__9_) );
  OR2X2 OR2X2_3338 ( .A(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1_1__10_), .Y(AES_CORE_DATAPATH__abc_16259_n9786) );
  OR2X2 OR2X2_3339 ( .A(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf1), .B(AES_CORE_DATAPATH_bkp_1_1__11_), .Y(AES_CORE_DATAPATH__abc_16259_n9790) );
  OR2X2 OR2X2_334 ( .A(AES_CORE_DATAPATH__abc_16259_n3088), .B(AES_CORE_DATAPATH__abc_16259_n3089), .Y(AES_CORE_DATAPATH__abc_16259_n3090_1) );
  OR2X2 OR2X2_3340 ( .A(AES_CORE_DATAPATH__abc_16259_n9793), .B(AES_CORE_DATAPATH__abc_16259_n9792), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__12_) );
  OR2X2 OR2X2_3341 ( .A(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf6), .B(AES_CORE_DATAPATH_bkp_1_1__13_), .Y(AES_CORE_DATAPATH__abc_16259_n9797) );
  OR2X2 OR2X2_3342 ( .A(AES_CORE_DATAPATH__abc_16259_n9800), .B(AES_CORE_DATAPATH__abc_16259_n9799), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__14_) );
  OR2X2 OR2X2_3343 ( .A(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1_1__15_), .Y(AES_CORE_DATAPATH__abc_16259_n9804) );
  OR2X2 OR2X2_3344 ( .A(AES_CORE_DATAPATH__abc_16259_n9807), .B(AES_CORE_DATAPATH__abc_16259_n9806), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__16_) );
  OR2X2 OR2X2_3345 ( .A(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf0), .B(AES_CORE_DATAPATH_bkp_1_1__17_), .Y(AES_CORE_DATAPATH__abc_16259_n9811) );
  OR2X2 OR2X2_3346 ( .A(AES_CORE_DATAPATH__abc_16259_n9814), .B(AES_CORE_DATAPATH__abc_16259_n9813), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__18_) );
  OR2X2 OR2X2_3347 ( .A(AES_CORE_DATAPATH__abc_16259_n9817), .B(AES_CORE_DATAPATH__abc_16259_n9816), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__19_) );
  OR2X2 OR2X2_3348 ( .A(AES_CORE_DATAPATH__abc_16259_n9820), .B(AES_CORE_DATAPATH__abc_16259_n9819), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__20_) );
  OR2X2 OR2X2_3349 ( .A(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1_1__21_), .Y(AES_CORE_DATAPATH__abc_16259_n9824) );
  OR2X2 OR2X2_335 ( .A(AES_CORE_DATAPATH__abc_16259_n3090_1), .B(AES_CORE_DATAPATH__abc_16259_n3087), .Y(AES_CORE_DATAPATH__abc_16259_n3091_1) );
  OR2X2 OR2X2_3350 ( .A(AES_CORE_DATAPATH__abc_16259_n9827), .B(AES_CORE_DATAPATH__abc_16259_n9826), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__22_) );
  OR2X2 OR2X2_3351 ( .A(AES_CORE_DATAPATH__abc_16259_n9830), .B(AES_CORE_DATAPATH__abc_16259_n9829), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__23_) );
  OR2X2 OR2X2_3352 ( .A(AES_CORE_DATAPATH__abc_16259_n9833), .B(AES_CORE_DATAPATH__abc_16259_n9832), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__24_) );
  OR2X2 OR2X2_3353 ( .A(AES_CORE_DATAPATH__abc_16259_n9836), .B(AES_CORE_DATAPATH__abc_16259_n9835), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__25_) );
  OR2X2 OR2X2_3354 ( .A(AES_CORE_DATAPATH__abc_16259_n9839), .B(AES_CORE_DATAPATH__abc_16259_n9838), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__26_) );
  OR2X2 OR2X2_3355 ( .A(AES_CORE_DATAPATH__abc_16259_n9842), .B(AES_CORE_DATAPATH__abc_16259_n9841), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__27_) );
  OR2X2 OR2X2_3356 ( .A(AES_CORE_DATAPATH__abc_16259_n9845), .B(AES_CORE_DATAPATH__abc_16259_n9844), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__28_) );
  OR2X2 OR2X2_3357 ( .A(AES_CORE_DATAPATH__abc_16259_n9848), .B(AES_CORE_DATAPATH__abc_16259_n9847), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__29_) );
  OR2X2 OR2X2_3358 ( .A(AES_CORE_DATAPATH__abc_16259_n9851), .B(AES_CORE_DATAPATH__abc_16259_n9850), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__30_) );
  OR2X2 OR2X2_3359 ( .A(AES_CORE_DATAPATH__abc_16259_n9854), .B(AES_CORE_DATAPATH__abc_16259_n9853), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__31_) );
  OR2X2 OR2X2_336 ( .A(AES_CORE_DATAPATH__abc_16259_n2841_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__6_), .Y(AES_CORE_DATAPATH__abc_16259_n3092) );
  OR2X2 OR2X2_3360 ( .A(AES_CORE_DATAPATH__abc_16259_n7950), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n9856) );
  OR2X2 OR2X2_3361 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf5), .B(AES_CORE_DATAPATH_bkp_1_1__0_), .Y(AES_CORE_DATAPATH__abc_16259_n9857) );
  OR2X2 OR2X2_3362 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n8608), .Y(AES_CORE_DATAPATH__abc_16259_n9860) );
  OR2X2 OR2X2_3363 ( .A(AES_CORE_DATAPATH__abc_16259_n9859), .B(AES_CORE_DATAPATH__abc_16259_n9860), .Y(AES_CORE_DATAPATH__abc_16259_n9861) );
  OR2X2 OR2X2_3364 ( .A(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf0), .B(AES_CORE_DATAPATH_bkp_1__0_), .Y(AES_CORE_DATAPATH__abc_16259_n9862) );
  OR2X2 OR2X2_3365 ( .A(AES_CORE_DATAPATH__abc_16259_n7958), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n9864) );
  OR2X2 OR2X2_3366 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf4), .B(AES_CORE_DATAPATH_bkp_1_1__1_), .Y(AES_CORE_DATAPATH__abc_16259_n9865) );
  OR2X2 OR2X2_3367 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n8617), .Y(AES_CORE_DATAPATH__abc_16259_n9868) );
  OR2X2 OR2X2_3368 ( .A(AES_CORE_DATAPATH__abc_16259_n9867), .B(AES_CORE_DATAPATH__abc_16259_n9868), .Y(AES_CORE_DATAPATH__abc_16259_n9869) );
  OR2X2 OR2X2_3369 ( .A(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf7), .B(AES_CORE_DATAPATH_bkp_1__1_), .Y(AES_CORE_DATAPATH__abc_16259_n9870) );
  OR2X2 OR2X2_337 ( .A(AES_CORE_DATAPATH__abc_16259_n3084), .B(AES_CORE_DATAPATH__abc_16259_n2853_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n3094_1) );
  OR2X2 OR2X2_3370 ( .A(AES_CORE_DATAPATH__abc_16259_n7966), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n9872) );
  OR2X2 OR2X2_3371 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1_1__2_), .Y(AES_CORE_DATAPATH__abc_16259_n9873) );
  OR2X2 OR2X2_3372 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf6), .B(AES_CORE_DATAPATH__abc_16259_n8626), .Y(AES_CORE_DATAPATH__abc_16259_n9876) );
  OR2X2 OR2X2_3373 ( .A(AES_CORE_DATAPATH__abc_16259_n9875), .B(AES_CORE_DATAPATH__abc_16259_n9876), .Y(AES_CORE_DATAPATH__abc_16259_n9877) );
  OR2X2 OR2X2_3374 ( .A(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf6), .B(AES_CORE_DATAPATH_bkp_1__2_), .Y(AES_CORE_DATAPATH__abc_16259_n9878) );
  OR2X2 OR2X2_3375 ( .A(AES_CORE_DATAPATH__abc_16259_n7974), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n9880) );
  OR2X2 OR2X2_3376 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf2), .B(AES_CORE_DATAPATH_bkp_1_1__3_), .Y(AES_CORE_DATAPATH__abc_16259_n9881) );
  OR2X2 OR2X2_3377 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf5), .B(AES_CORE_DATAPATH__abc_16259_n8635), .Y(AES_CORE_DATAPATH__abc_16259_n9884) );
  OR2X2 OR2X2_3378 ( .A(AES_CORE_DATAPATH__abc_16259_n9883), .B(AES_CORE_DATAPATH__abc_16259_n9884), .Y(AES_CORE_DATAPATH__abc_16259_n9885) );
  OR2X2 OR2X2_3379 ( .A(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf5), .B(AES_CORE_DATAPATH_bkp_1__3_), .Y(AES_CORE_DATAPATH__abc_16259_n9886) );
  OR2X2 OR2X2_338 ( .A(AES_CORE_DATAPATH__abc_16259_n3095), .B(AES_CORE_DATAPATH__abc_16259_n3096_1), .Y(AES_CORE_DATAPATH__abc_16259_n3097) );
  OR2X2 OR2X2_3380 ( .A(AES_CORE_DATAPATH__abc_16259_n7982), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n9888) );
  OR2X2 OR2X2_3381 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf1), .B(AES_CORE_DATAPATH_bkp_1_1__4_), .Y(AES_CORE_DATAPATH__abc_16259_n9889) );
  OR2X2 OR2X2_3382 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n8644), .Y(AES_CORE_DATAPATH__abc_16259_n9892) );
  OR2X2 OR2X2_3383 ( .A(AES_CORE_DATAPATH__abc_16259_n9891), .B(AES_CORE_DATAPATH__abc_16259_n9892), .Y(AES_CORE_DATAPATH__abc_16259_n9893) );
  OR2X2 OR2X2_3384 ( .A(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf4), .B(AES_CORE_DATAPATH_bkp_1__4_), .Y(AES_CORE_DATAPATH__abc_16259_n9894) );
  OR2X2 OR2X2_3385 ( .A(AES_CORE_DATAPATH__abc_16259_n7990), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n9896) );
  OR2X2 OR2X2_3386 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf0), .B(AES_CORE_DATAPATH_bkp_1_1__5_), .Y(AES_CORE_DATAPATH__abc_16259_n9897) );
  OR2X2 OR2X2_3387 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n8653), .Y(AES_CORE_DATAPATH__abc_16259_n9900) );
  OR2X2 OR2X2_3388 ( .A(AES_CORE_DATAPATH__abc_16259_n9899), .B(AES_CORE_DATAPATH__abc_16259_n9900), .Y(AES_CORE_DATAPATH__abc_16259_n9901) );
  OR2X2 OR2X2_3389 ( .A(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1__5_), .Y(AES_CORE_DATAPATH__abc_16259_n9902) );
  OR2X2 OR2X2_339 ( .A(_auto_iopadmap_cc_313_execute_26949_6_), .B(AES_CORE_DATAPATH__abc_16259_n3099), .Y(AES_CORE_DATAPATH__abc_16259_n3100_1) );
  OR2X2 OR2X2_3390 ( .A(AES_CORE_DATAPATH__abc_16259_n7998), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n9904) );
  OR2X2 OR2X2_3391 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf11), .B(AES_CORE_DATAPATH_bkp_1_1__6_), .Y(AES_CORE_DATAPATH__abc_16259_n9905) );
  OR2X2 OR2X2_3392 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n8662), .Y(AES_CORE_DATAPATH__abc_16259_n9908) );
  OR2X2 OR2X2_3393 ( .A(AES_CORE_DATAPATH__abc_16259_n9907), .B(AES_CORE_DATAPATH__abc_16259_n9908), .Y(AES_CORE_DATAPATH__abc_16259_n9909) );
  OR2X2 OR2X2_3394 ( .A(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf2), .B(AES_CORE_DATAPATH_bkp_1__6_), .Y(AES_CORE_DATAPATH__abc_16259_n9910) );
  OR2X2 OR2X2_3395 ( .A(AES_CORE_DATAPATH__abc_16259_n8006), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n9912) );
  OR2X2 OR2X2_3396 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf10), .B(AES_CORE_DATAPATH_bkp_1_1__7_), .Y(AES_CORE_DATAPATH__abc_16259_n9913) );
  OR2X2 OR2X2_3397 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n8671), .Y(AES_CORE_DATAPATH__abc_16259_n9916) );
  OR2X2 OR2X2_3398 ( .A(AES_CORE_DATAPATH__abc_16259_n9915), .B(AES_CORE_DATAPATH__abc_16259_n9916), .Y(AES_CORE_DATAPATH__abc_16259_n9917) );
  OR2X2 OR2X2_3399 ( .A(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf1), .B(AES_CORE_DATAPATH_bkp_1__7_), .Y(AES_CORE_DATAPATH__abc_16259_n9918) );
  OR2X2 OR2X2_34 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n169), .B(AES_CORE_CONTROL_UNIT_rd_count_1_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n175_1) );
  OR2X2 OR2X2_340 ( .A(AES_CORE_DATAPATH__abc_16259_n3102), .B(AES_CORE_DATAPATH__abc_16259_n2864_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n3103) );
  OR2X2 OR2X2_3400 ( .A(AES_CORE_DATAPATH__abc_16259_n8014), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf9), .Y(AES_CORE_DATAPATH__abc_16259_n9920) );
  OR2X2 OR2X2_3401 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf9), .B(AES_CORE_DATAPATH_bkp_1_1__8_), .Y(AES_CORE_DATAPATH__abc_16259_n9921) );
  OR2X2 OR2X2_3402 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n8680), .Y(AES_CORE_DATAPATH__abc_16259_n9924) );
  OR2X2 OR2X2_3403 ( .A(AES_CORE_DATAPATH__abc_16259_n9923), .B(AES_CORE_DATAPATH__abc_16259_n9924), .Y(AES_CORE_DATAPATH__abc_16259_n9925) );
  OR2X2 OR2X2_3404 ( .A(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf0), .B(AES_CORE_DATAPATH_bkp_1__8_), .Y(AES_CORE_DATAPATH__abc_16259_n9926) );
  OR2X2 OR2X2_3405 ( .A(AES_CORE_DATAPATH__abc_16259_n8022), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf8), .Y(AES_CORE_DATAPATH__abc_16259_n9928) );
  OR2X2 OR2X2_3406 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf8), .B(AES_CORE_DATAPATH_bkp_1_1__9_), .Y(AES_CORE_DATAPATH__abc_16259_n9929) );
  OR2X2 OR2X2_3407 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf6), .B(AES_CORE_DATAPATH__abc_16259_n8689), .Y(AES_CORE_DATAPATH__abc_16259_n9932) );
  OR2X2 OR2X2_3408 ( .A(AES_CORE_DATAPATH__abc_16259_n9931), .B(AES_CORE_DATAPATH__abc_16259_n9932), .Y(AES_CORE_DATAPATH__abc_16259_n9933) );
  OR2X2 OR2X2_3409 ( .A(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf7), .B(AES_CORE_DATAPATH_bkp_1__9_), .Y(AES_CORE_DATAPATH__abc_16259_n9934) );
  OR2X2 OR2X2_341 ( .A(AES_CORE_DATAPATH__abc_16259_n3103), .B(AES_CORE_DATAPATH__abc_16259_n3101), .Y(AES_CORE_DATAPATH__abc_16259_n3104) );
  OR2X2 OR2X2_3410 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf6), .B(AES_CORE_DATAPATH_bkp_1_1__10_), .Y(AES_CORE_DATAPATH__abc_16259_n9938) );
  OR2X2 OR2X2_3411 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf5), .B(AES_CORE_DATAPATH__abc_16259_n8699), .Y(AES_CORE_DATAPATH__abc_16259_n9941) );
  OR2X2 OR2X2_3412 ( .A(AES_CORE_DATAPATH__abc_16259_n9940), .B(AES_CORE_DATAPATH__abc_16259_n9941), .Y(AES_CORE_DATAPATH__abc_16259_n9942) );
  OR2X2 OR2X2_3413 ( .A(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf6), .B(AES_CORE_DATAPATH_bkp_1__10_), .Y(AES_CORE_DATAPATH__abc_16259_n9943) );
  OR2X2 OR2X2_3414 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf4), .B(AES_CORE_DATAPATH_bkp_1_1__11_), .Y(AES_CORE_DATAPATH__abc_16259_n9947) );
  OR2X2 OR2X2_3415 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n8709), .Y(AES_CORE_DATAPATH__abc_16259_n9950) );
  OR2X2 OR2X2_3416 ( .A(AES_CORE_DATAPATH__abc_16259_n9949), .B(AES_CORE_DATAPATH__abc_16259_n9950), .Y(AES_CORE_DATAPATH__abc_16259_n9951) );
  OR2X2 OR2X2_3417 ( .A(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf5), .B(AES_CORE_DATAPATH_bkp_1__11_), .Y(AES_CORE_DATAPATH__abc_16259_n9952) );
  OR2X2 OR2X2_3418 ( .A(AES_CORE_DATAPATH__abc_16259_n8052), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n9954) );
  OR2X2 OR2X2_3419 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1_1__12_), .Y(AES_CORE_DATAPATH__abc_16259_n9955) );
  OR2X2 OR2X2_342 ( .A(AES_CORE_DATAPATH__abc_16259_n3106), .B(AES_CORE_DATAPATH__abc_16259_n3105), .Y(AES_CORE_DATAPATH__abc_16259_n3107) );
  OR2X2 OR2X2_3420 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n8718), .Y(AES_CORE_DATAPATH__abc_16259_n9958) );
  OR2X2 OR2X2_3421 ( .A(AES_CORE_DATAPATH__abc_16259_n9957), .B(AES_CORE_DATAPATH__abc_16259_n9958), .Y(AES_CORE_DATAPATH__abc_16259_n9959) );
  OR2X2 OR2X2_3422 ( .A(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf4), .B(AES_CORE_DATAPATH_bkp_1__12_), .Y(AES_CORE_DATAPATH__abc_16259_n9960) );
  OR2X2 OR2X2_3423 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf1), .B(AES_CORE_DATAPATH_bkp_1_1__13_), .Y(AES_CORE_DATAPATH__abc_16259_n9964) );
  OR2X2 OR2X2_3424 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n8728), .Y(AES_CORE_DATAPATH__abc_16259_n9967) );
  OR2X2 OR2X2_3425 ( .A(AES_CORE_DATAPATH__abc_16259_n9966), .B(AES_CORE_DATAPATH__abc_16259_n9967), .Y(AES_CORE_DATAPATH__abc_16259_n9968) );
  OR2X2 OR2X2_3426 ( .A(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1__13_), .Y(AES_CORE_DATAPATH__abc_16259_n9969) );
  OR2X2 OR2X2_3427 ( .A(AES_CORE_DATAPATH__abc_16259_n8071), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n9971) );
  OR2X2 OR2X2_3428 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf0), .B(AES_CORE_DATAPATH_bkp_1_1__14_), .Y(AES_CORE_DATAPATH__abc_16259_n9972) );
  OR2X2 OR2X2_3429 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n8737), .Y(AES_CORE_DATAPATH__abc_16259_n9975) );
  OR2X2 OR2X2_343 ( .A(AES_CORE_DATAPATH__abc_16259_n3107), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n3108) );
  OR2X2 OR2X2_3430 ( .A(AES_CORE_DATAPATH__abc_16259_n9974), .B(AES_CORE_DATAPATH__abc_16259_n9975), .Y(AES_CORE_DATAPATH__abc_16259_n9976) );
  OR2X2 OR2X2_3431 ( .A(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf2), .B(AES_CORE_DATAPATH_bkp_1__14_), .Y(AES_CORE_DATAPATH__abc_16259_n9977) );
  OR2X2 OR2X2_3432 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf10), .B(AES_CORE_DATAPATH_bkp_1_1__15_), .Y(AES_CORE_DATAPATH__abc_16259_n9981) );
  OR2X2 OR2X2_3433 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n8747), .Y(AES_CORE_DATAPATH__abc_16259_n9984) );
  OR2X2 OR2X2_3434 ( .A(AES_CORE_DATAPATH__abc_16259_n9983), .B(AES_CORE_DATAPATH__abc_16259_n9984), .Y(AES_CORE_DATAPATH__abc_16259_n9985) );
  OR2X2 OR2X2_3435 ( .A(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf1), .B(AES_CORE_DATAPATH_bkp_1__15_), .Y(AES_CORE_DATAPATH__abc_16259_n9986) );
  OR2X2 OR2X2_3436 ( .A(AES_CORE_DATAPATH__abc_16259_n8090), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n9988) );
  OR2X2 OR2X2_3437 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf9), .B(AES_CORE_DATAPATH_bkp_1_1__16_), .Y(AES_CORE_DATAPATH__abc_16259_n9989) );
  OR2X2 OR2X2_3438 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf6), .B(AES_CORE_DATAPATH__abc_16259_n8756), .Y(AES_CORE_DATAPATH__abc_16259_n9992) );
  OR2X2 OR2X2_3439 ( .A(AES_CORE_DATAPATH__abc_16259_n9991), .B(AES_CORE_DATAPATH__abc_16259_n9992), .Y(AES_CORE_DATAPATH__abc_16259_n9993) );
  OR2X2 OR2X2_344 ( .A(AES_CORE_DATAPATH__abc_16259_n3110), .B(AES_CORE_DATAPATH__abc_16259_n3111), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_6_) );
  OR2X2 OR2X2_3440 ( .A(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf0), .B(AES_CORE_DATAPATH_bkp_1__16_), .Y(AES_CORE_DATAPATH__abc_16259_n9994) );
  OR2X2 OR2X2_3441 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf7), .B(AES_CORE_DATAPATH_bkp_1_1__17_), .Y(AES_CORE_DATAPATH__abc_16259_n9998) );
  OR2X2 OR2X2_3442 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf5), .B(AES_CORE_DATAPATH__abc_16259_n8766), .Y(AES_CORE_DATAPATH__abc_16259_n10001) );
  OR2X2 OR2X2_3443 ( .A(AES_CORE_DATAPATH__abc_16259_n10000), .B(AES_CORE_DATAPATH__abc_16259_n10001), .Y(AES_CORE_DATAPATH__abc_16259_n10002) );
  OR2X2 OR2X2_3444 ( .A(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf7), .B(AES_CORE_DATAPATH_bkp_1__17_), .Y(AES_CORE_DATAPATH__abc_16259_n10003) );
  OR2X2 OR2X2_3445 ( .A(AES_CORE_DATAPATH__abc_16259_n8109), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n10005) );
  OR2X2 OR2X2_3446 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf6), .B(AES_CORE_DATAPATH_bkp_1_1__18_), .Y(AES_CORE_DATAPATH__abc_16259_n10006) );
  OR2X2 OR2X2_3447 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n8775), .Y(AES_CORE_DATAPATH__abc_16259_n10009) );
  OR2X2 OR2X2_3448 ( .A(AES_CORE_DATAPATH__abc_16259_n10008), .B(AES_CORE_DATAPATH__abc_16259_n10009), .Y(AES_CORE_DATAPATH__abc_16259_n10010) );
  OR2X2 OR2X2_3449 ( .A(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf6), .B(AES_CORE_DATAPATH_bkp_1__18_), .Y(AES_CORE_DATAPATH__abc_16259_n10011) );
  OR2X2 OR2X2_345 ( .A(AES_CORE_DATAPATH__abc_16259_n2774_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n3113), .Y(AES_CORE_DATAPATH__abc_16259_n3114_1) );
  OR2X2 OR2X2_3450 ( .A(AES_CORE_DATAPATH__abc_16259_n8117), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n10013) );
  OR2X2 OR2X2_3451 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf5), .B(AES_CORE_DATAPATH_bkp_1_1__19_), .Y(AES_CORE_DATAPATH__abc_16259_n10014) );
  OR2X2 OR2X2_3452 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n8784), .Y(AES_CORE_DATAPATH__abc_16259_n10017) );
  OR2X2 OR2X2_3453 ( .A(AES_CORE_DATAPATH__abc_16259_n10016), .B(AES_CORE_DATAPATH__abc_16259_n10017), .Y(AES_CORE_DATAPATH__abc_16259_n10018) );
  OR2X2 OR2X2_3454 ( .A(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf5), .B(AES_CORE_DATAPATH_bkp_1__19_), .Y(AES_CORE_DATAPATH__abc_16259_n10019) );
  OR2X2 OR2X2_3455 ( .A(AES_CORE_DATAPATH__abc_16259_n8125), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n10021) );
  OR2X2 OR2X2_3456 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf4), .B(AES_CORE_DATAPATH_bkp_1_1__20_), .Y(AES_CORE_DATAPATH__abc_16259_n10022) );
  OR2X2 OR2X2_3457 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n8793), .Y(AES_CORE_DATAPATH__abc_16259_n10025) );
  OR2X2 OR2X2_3458 ( .A(AES_CORE_DATAPATH__abc_16259_n10024), .B(AES_CORE_DATAPATH__abc_16259_n10025), .Y(AES_CORE_DATAPATH__abc_16259_n10026) );
  OR2X2 OR2X2_3459 ( .A(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf4), .B(AES_CORE_DATAPATH_bkp_1__20_), .Y(AES_CORE_DATAPATH__abc_16259_n10027) );
  OR2X2 OR2X2_346 ( .A(AES_CORE_DATAPATH__abc_16259_n2778_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n3115), .Y(AES_CORE_DATAPATH__abc_16259_n3116) );
  OR2X2 OR2X2_3460 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf2), .B(AES_CORE_DATAPATH_bkp_1_1__21_), .Y(AES_CORE_DATAPATH__abc_16259_n10031) );
  OR2X2 OR2X2_3461 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n8803), .Y(AES_CORE_DATAPATH__abc_16259_n10034) );
  OR2X2 OR2X2_3462 ( .A(AES_CORE_DATAPATH__abc_16259_n10033), .B(AES_CORE_DATAPATH__abc_16259_n10034), .Y(AES_CORE_DATAPATH__abc_16259_n10035) );
  OR2X2 OR2X2_3463 ( .A(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1__21_), .Y(AES_CORE_DATAPATH__abc_16259_n10036) );
  OR2X2 OR2X2_3464 ( .A(AES_CORE_DATAPATH__abc_16259_n8144), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n10038) );
  OR2X2 OR2X2_3465 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf1), .B(AES_CORE_DATAPATH_bkp_1_1__22_), .Y(AES_CORE_DATAPATH__abc_16259_n10039) );
  OR2X2 OR2X2_3466 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n8812), .Y(AES_CORE_DATAPATH__abc_16259_n10042) );
  OR2X2 OR2X2_3467 ( .A(AES_CORE_DATAPATH__abc_16259_n10041), .B(AES_CORE_DATAPATH__abc_16259_n10042), .Y(AES_CORE_DATAPATH__abc_16259_n10043) );
  OR2X2 OR2X2_3468 ( .A(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf2), .B(AES_CORE_DATAPATH_bkp_1__22_), .Y(AES_CORE_DATAPATH__abc_16259_n10044) );
  OR2X2 OR2X2_3469 ( .A(AES_CORE_DATAPATH__abc_16259_n8152), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n10046) );
  OR2X2 OR2X2_347 ( .A(AES_CORE_DATAPATH__abc_16259_n3119_1), .B(AES_CORE_DATAPATH__abc_16259_n3120_1), .Y(AES_CORE_DATAPATH__abc_16259_n3121) );
  OR2X2 OR2X2_3470 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf0), .B(AES_CORE_DATAPATH_bkp_1_1__23_), .Y(AES_CORE_DATAPATH__abc_16259_n10047) );
  OR2X2 OR2X2_3471 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf6), .B(AES_CORE_DATAPATH__abc_16259_n8821), .Y(AES_CORE_DATAPATH__abc_16259_n10050) );
  OR2X2 OR2X2_3472 ( .A(AES_CORE_DATAPATH__abc_16259_n10049), .B(AES_CORE_DATAPATH__abc_16259_n10050), .Y(AES_CORE_DATAPATH__abc_16259_n10051) );
  OR2X2 OR2X2_3473 ( .A(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf1), .B(AES_CORE_DATAPATH_bkp_1__23_), .Y(AES_CORE_DATAPATH__abc_16259_n10052) );
  OR2X2 OR2X2_3474 ( .A(AES_CORE_DATAPATH__abc_16259_n8160), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf9), .Y(AES_CORE_DATAPATH__abc_16259_n10054) );
  OR2X2 OR2X2_3475 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf11), .B(AES_CORE_DATAPATH_bkp_1_1__24_), .Y(AES_CORE_DATAPATH__abc_16259_n10055) );
  OR2X2 OR2X2_3476 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf5), .B(AES_CORE_DATAPATH__abc_16259_n8830), .Y(AES_CORE_DATAPATH__abc_16259_n10058) );
  OR2X2 OR2X2_3477 ( .A(AES_CORE_DATAPATH__abc_16259_n10057), .B(AES_CORE_DATAPATH__abc_16259_n10058), .Y(AES_CORE_DATAPATH__abc_16259_n10059) );
  OR2X2 OR2X2_3478 ( .A(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf0), .B(AES_CORE_DATAPATH_bkp_1__24_), .Y(AES_CORE_DATAPATH__abc_16259_n10060) );
  OR2X2 OR2X2_3479 ( .A(AES_CORE_DATAPATH__abc_16259_n8168), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf8), .Y(AES_CORE_DATAPATH__abc_16259_n10062) );
  OR2X2 OR2X2_348 ( .A(AES_CORE_DATAPATH__abc_16259_n3121), .B(AES_CORE_DATAPATH__abc_16259_n3118), .Y(AES_CORE_DATAPATH__abc_16259_n3122) );
  OR2X2 OR2X2_3480 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf10), .B(AES_CORE_DATAPATH_bkp_1_1__25_), .Y(AES_CORE_DATAPATH__abc_16259_n10063) );
  OR2X2 OR2X2_3481 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n8839), .Y(AES_CORE_DATAPATH__abc_16259_n10066) );
  OR2X2 OR2X2_3482 ( .A(AES_CORE_DATAPATH__abc_16259_n10065), .B(AES_CORE_DATAPATH__abc_16259_n10066), .Y(AES_CORE_DATAPATH__abc_16259_n10067) );
  OR2X2 OR2X2_3483 ( .A(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf7), .B(AES_CORE_DATAPATH_bkp_1__25_), .Y(AES_CORE_DATAPATH__abc_16259_n10068) );
  OR2X2 OR2X2_3484 ( .A(AES_CORE_DATAPATH__abc_16259_n8176), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n10070) );
  OR2X2 OR2X2_3485 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf9), .B(AES_CORE_DATAPATH_bkp_1_1__26_), .Y(AES_CORE_DATAPATH__abc_16259_n10071) );
  OR2X2 OR2X2_3486 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n8848), .Y(AES_CORE_DATAPATH__abc_16259_n10074) );
  OR2X2 OR2X2_3487 ( .A(AES_CORE_DATAPATH__abc_16259_n10073), .B(AES_CORE_DATAPATH__abc_16259_n10074), .Y(AES_CORE_DATAPATH__abc_16259_n10075) );
  OR2X2 OR2X2_3488 ( .A(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf6), .B(AES_CORE_DATAPATH_bkp_1__26_), .Y(AES_CORE_DATAPATH__abc_16259_n10076) );
  OR2X2 OR2X2_3489 ( .A(AES_CORE_DATAPATH__abc_16259_n8184), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n10078) );
  OR2X2 OR2X2_349 ( .A(AES_CORE_DATAPATH__abc_16259_n3126), .B(AES_CORE_DATAPATH__abc_16259_n2826_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n3127_1) );
  OR2X2 OR2X2_3490 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf8), .B(AES_CORE_DATAPATH_bkp_1_1__27_), .Y(AES_CORE_DATAPATH__abc_16259_n10079) );
  OR2X2 OR2X2_3491 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n8857), .Y(AES_CORE_DATAPATH__abc_16259_n10082) );
  OR2X2 OR2X2_3492 ( .A(AES_CORE_DATAPATH__abc_16259_n10081), .B(AES_CORE_DATAPATH__abc_16259_n10082), .Y(AES_CORE_DATAPATH__abc_16259_n10083) );
  OR2X2 OR2X2_3493 ( .A(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf5), .B(AES_CORE_DATAPATH_bkp_1__27_), .Y(AES_CORE_DATAPATH__abc_16259_n10084) );
  OR2X2 OR2X2_3494 ( .A(AES_CORE_DATAPATH__abc_16259_n8192), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n10086) );
  OR2X2 OR2X2_3495 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf7), .B(AES_CORE_DATAPATH_bkp_1_1__28_), .Y(AES_CORE_DATAPATH__abc_16259_n10087) );
  OR2X2 OR2X2_3496 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n8866), .Y(AES_CORE_DATAPATH__abc_16259_n10090) );
  OR2X2 OR2X2_3497 ( .A(AES_CORE_DATAPATH__abc_16259_n10089), .B(AES_CORE_DATAPATH__abc_16259_n10090), .Y(AES_CORE_DATAPATH__abc_16259_n10091) );
  OR2X2 OR2X2_3498 ( .A(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf4), .B(AES_CORE_DATAPATH_bkp_1__28_), .Y(AES_CORE_DATAPATH__abc_16259_n10092) );
  OR2X2 OR2X2_3499 ( .A(AES_CORE_DATAPATH__abc_16259_n8200), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n10094) );
  OR2X2 OR2X2_35 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n173), .B(AES_CORE_CONTROL_UNIT_rd_count_2_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n180) );
  OR2X2 OR2X2_350 ( .A(AES_CORE_DATAPATH__abc_16259_n3128), .B(AES_CORE_DATAPATH__abc_16259_n3129_1), .Y(AES_CORE_DATAPATH__abc_16259_n3130) );
  OR2X2 OR2X2_3500 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf6), .B(AES_CORE_DATAPATH_bkp_1_1__29_), .Y(AES_CORE_DATAPATH__abc_16259_n10095) );
  OR2X2 OR2X2_3501 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n8875), .Y(AES_CORE_DATAPATH__abc_16259_n10098) );
  OR2X2 OR2X2_3502 ( .A(AES_CORE_DATAPATH__abc_16259_n10097), .B(AES_CORE_DATAPATH__abc_16259_n10098), .Y(AES_CORE_DATAPATH__abc_16259_n10099) );
  OR2X2 OR2X2_3503 ( .A(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1__29_), .Y(AES_CORE_DATAPATH__abc_16259_n10100) );
  OR2X2 OR2X2_3504 ( .A(AES_CORE_DATAPATH__abc_16259_n8208), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n10102) );
  OR2X2 OR2X2_3505 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf5), .B(AES_CORE_DATAPATH_bkp_1_1__30_), .Y(AES_CORE_DATAPATH__abc_16259_n10103) );
  OR2X2 OR2X2_3506 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf6), .B(AES_CORE_DATAPATH__abc_16259_n8884), .Y(AES_CORE_DATAPATH__abc_16259_n10106) );
  OR2X2 OR2X2_3507 ( .A(AES_CORE_DATAPATH__abc_16259_n10105), .B(AES_CORE_DATAPATH__abc_16259_n10106), .Y(AES_CORE_DATAPATH__abc_16259_n10107) );
  OR2X2 OR2X2_3508 ( .A(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf2), .B(AES_CORE_DATAPATH_bkp_1__30_), .Y(AES_CORE_DATAPATH__abc_16259_n10108) );
  OR2X2 OR2X2_3509 ( .A(AES_CORE_DATAPATH__abc_16259_n8216), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n10110) );
  OR2X2 OR2X2_351 ( .A(AES_CORE_DATAPATH__abc_16259_n3130), .B(AES_CORE_DATAPATH__abc_16259_n3127_1), .Y(AES_CORE_DATAPATH__abc_16259_n3131) );
  OR2X2 OR2X2_3510 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf4), .B(AES_CORE_DATAPATH_bkp_1_1__31_), .Y(AES_CORE_DATAPATH__abc_16259_n10111) );
  OR2X2 OR2X2_3511 ( .A(AES_CORE_DATAPATH__abc_16259_n9753_bF_buf5), .B(AES_CORE_DATAPATH__abc_16259_n8893), .Y(AES_CORE_DATAPATH__abc_16259_n10114) );
  OR2X2 OR2X2_3512 ( .A(AES_CORE_DATAPATH__abc_16259_n10113), .B(AES_CORE_DATAPATH__abc_16259_n10114), .Y(AES_CORE_DATAPATH__abc_16259_n10115) );
  OR2X2 OR2X2_3513 ( .A(AES_CORE_DATAPATH__abc_16259_n9752_bF_buf1), .B(AES_CORE_DATAPATH_bkp_1__31_), .Y(AES_CORE_DATAPATH__abc_16259_n10116) );
  OR2X2 OR2X2_3514 ( .A(AES_CORE_DATAPATH_iv_1__0_), .B(iv_en_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n10118) );
  OR2X2 OR2X2_3515 ( .A(AES_CORE_DATAPATH__abc_16259_n10119_bF_buf4), .B(\bus_in[0] ), .Y(AES_CORE_DATAPATH__abc_16259_n10120) );
  OR2X2 OR2X2_3516 ( .A(AES_CORE_DATAPATH_iv_1__1_), .B(iv_en_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n10122) );
  OR2X2 OR2X2_3517 ( .A(AES_CORE_DATAPATH__abc_16259_n10119_bF_buf3), .B(\bus_in[1] ), .Y(AES_CORE_DATAPATH__abc_16259_n10123) );
  OR2X2 OR2X2_3518 ( .A(AES_CORE_DATAPATH_iv_1__2_), .B(iv_en_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n10125) );
  OR2X2 OR2X2_3519 ( .A(AES_CORE_DATAPATH__abc_16259_n10119_bF_buf2), .B(\bus_in[2] ), .Y(AES_CORE_DATAPATH__abc_16259_n10126) );
  OR2X2 OR2X2_352 ( .A(AES_CORE_DATAPATH__abc_16259_n2841_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__7_), .Y(AES_CORE_DATAPATH__abc_16259_n3132) );
  OR2X2 OR2X2_3520 ( .A(AES_CORE_DATAPATH_iv_1__3_), .B(iv_en_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n10128) );
  OR2X2 OR2X2_3521 ( .A(AES_CORE_DATAPATH__abc_16259_n10119_bF_buf1), .B(\bus_in[3] ), .Y(AES_CORE_DATAPATH__abc_16259_n10129) );
  OR2X2 OR2X2_3522 ( .A(AES_CORE_DATAPATH_iv_1__4_), .B(iv_en_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n10131) );
  OR2X2 OR2X2_3523 ( .A(AES_CORE_DATAPATH__abc_16259_n10119_bF_buf0), .B(\bus_in[4] ), .Y(AES_CORE_DATAPATH__abc_16259_n10132) );
  OR2X2 OR2X2_3524 ( .A(AES_CORE_DATAPATH_iv_1__5_), .B(iv_en_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n10134) );
  OR2X2 OR2X2_3525 ( .A(AES_CORE_DATAPATH__abc_16259_n10119_bF_buf4), .B(\bus_in[5] ), .Y(AES_CORE_DATAPATH__abc_16259_n10135) );
  OR2X2 OR2X2_3526 ( .A(AES_CORE_DATAPATH_iv_1__6_), .B(iv_en_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n10137) );
  OR2X2 OR2X2_3527 ( .A(AES_CORE_DATAPATH__abc_16259_n10119_bF_buf3), .B(\bus_in[6] ), .Y(AES_CORE_DATAPATH__abc_16259_n10138) );
  OR2X2 OR2X2_3528 ( .A(AES_CORE_DATAPATH_iv_1__7_), .B(iv_en_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n10140) );
  OR2X2 OR2X2_3529 ( .A(AES_CORE_DATAPATH__abc_16259_n10119_bF_buf2), .B(\bus_in[7] ), .Y(AES_CORE_DATAPATH__abc_16259_n10141) );
  OR2X2 OR2X2_353 ( .A(AES_CORE_DATAPATH__abc_16259_n3124), .B(AES_CORE_DATAPATH__abc_16259_n2853_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n3134) );
  OR2X2 OR2X2_3530 ( .A(AES_CORE_DATAPATH_iv_1__8_), .B(iv_en_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n10143) );
  OR2X2 OR2X2_3531 ( .A(AES_CORE_DATAPATH__abc_16259_n10119_bF_buf1), .B(\bus_in[8] ), .Y(AES_CORE_DATAPATH__abc_16259_n10144) );
  OR2X2 OR2X2_3532 ( .A(AES_CORE_DATAPATH_iv_1__9_), .B(iv_en_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n10146) );
  OR2X2 OR2X2_3533 ( .A(AES_CORE_DATAPATH__abc_16259_n10119_bF_buf0), .B(\bus_in[9] ), .Y(AES_CORE_DATAPATH__abc_16259_n10147) );
  OR2X2 OR2X2_3534 ( .A(AES_CORE_DATAPATH_iv_1__10_), .B(iv_en_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n10149) );
  OR2X2 OR2X2_3535 ( .A(AES_CORE_DATAPATH__abc_16259_n10119_bF_buf4), .B(\bus_in[10] ), .Y(AES_CORE_DATAPATH__abc_16259_n10150) );
  OR2X2 OR2X2_3536 ( .A(AES_CORE_DATAPATH_iv_1__11_), .B(iv_en_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n10152) );
  OR2X2 OR2X2_3537 ( .A(AES_CORE_DATAPATH__abc_16259_n10119_bF_buf3), .B(\bus_in[11] ), .Y(AES_CORE_DATAPATH__abc_16259_n10153) );
  OR2X2 OR2X2_3538 ( .A(AES_CORE_DATAPATH_iv_1__12_), .B(iv_en_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n10155) );
  OR2X2 OR2X2_3539 ( .A(AES_CORE_DATAPATH__abc_16259_n10119_bF_buf2), .B(\bus_in[12] ), .Y(AES_CORE_DATAPATH__abc_16259_n10156) );
  OR2X2 OR2X2_354 ( .A(AES_CORE_DATAPATH__abc_16259_n3135), .B(AES_CORE_DATAPATH__abc_16259_n3136), .Y(AES_CORE_DATAPATH__abc_16259_n3137) );
  OR2X2 OR2X2_3540 ( .A(AES_CORE_DATAPATH_iv_1__13_), .B(iv_en_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n10158) );
  OR2X2 OR2X2_3541 ( .A(AES_CORE_DATAPATH__abc_16259_n10119_bF_buf1), .B(\bus_in[13] ), .Y(AES_CORE_DATAPATH__abc_16259_n10159) );
  OR2X2 OR2X2_3542 ( .A(AES_CORE_DATAPATH_iv_1__14_), .B(iv_en_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n10161) );
  OR2X2 OR2X2_3543 ( .A(AES_CORE_DATAPATH__abc_16259_n10119_bF_buf0), .B(\bus_in[14] ), .Y(AES_CORE_DATAPATH__abc_16259_n10162) );
  OR2X2 OR2X2_3544 ( .A(AES_CORE_DATAPATH_iv_1__15_), .B(iv_en_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n10164) );
  OR2X2 OR2X2_3545 ( .A(AES_CORE_DATAPATH__abc_16259_n10119_bF_buf4), .B(\bus_in[15] ), .Y(AES_CORE_DATAPATH__abc_16259_n10165) );
  OR2X2 OR2X2_3546 ( .A(AES_CORE_DATAPATH_iv_1__16_), .B(iv_en_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n10167) );
  OR2X2 OR2X2_3547 ( .A(AES_CORE_DATAPATH__abc_16259_n10119_bF_buf3), .B(\bus_in[16] ), .Y(AES_CORE_DATAPATH__abc_16259_n10168) );
  OR2X2 OR2X2_3548 ( .A(AES_CORE_DATAPATH_iv_1__17_), .B(iv_en_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n10170) );
  OR2X2 OR2X2_3549 ( .A(AES_CORE_DATAPATH__abc_16259_n10119_bF_buf2), .B(\bus_in[17] ), .Y(AES_CORE_DATAPATH__abc_16259_n10171) );
  OR2X2 OR2X2_355 ( .A(_auto_iopadmap_cc_313_execute_26949_7_), .B(AES_CORE_DATAPATH__abc_16259_n3139), .Y(AES_CORE_DATAPATH__abc_16259_n3140) );
  OR2X2 OR2X2_3550 ( .A(AES_CORE_DATAPATH_iv_1__18_), .B(iv_en_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n10173) );
  OR2X2 OR2X2_3551 ( .A(AES_CORE_DATAPATH__abc_16259_n10119_bF_buf1), .B(\bus_in[18] ), .Y(AES_CORE_DATAPATH__abc_16259_n10174) );
  OR2X2 OR2X2_3552 ( .A(AES_CORE_DATAPATH_iv_1__19_), .B(iv_en_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n10176) );
  OR2X2 OR2X2_3553 ( .A(AES_CORE_DATAPATH__abc_16259_n10119_bF_buf0), .B(\bus_in[19] ), .Y(AES_CORE_DATAPATH__abc_16259_n10177) );
  OR2X2 OR2X2_3554 ( .A(AES_CORE_DATAPATH_iv_1__20_), .B(iv_en_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n10179) );
  OR2X2 OR2X2_3555 ( .A(AES_CORE_DATAPATH__abc_16259_n10119_bF_buf4), .B(\bus_in[20] ), .Y(AES_CORE_DATAPATH__abc_16259_n10180) );
  OR2X2 OR2X2_3556 ( .A(AES_CORE_DATAPATH_iv_1__21_), .B(iv_en_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n10182) );
  OR2X2 OR2X2_3557 ( .A(AES_CORE_DATAPATH__abc_16259_n10119_bF_buf3), .B(\bus_in[21] ), .Y(AES_CORE_DATAPATH__abc_16259_n10183) );
  OR2X2 OR2X2_3558 ( .A(AES_CORE_DATAPATH_iv_1__22_), .B(iv_en_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n10185) );
  OR2X2 OR2X2_3559 ( .A(AES_CORE_DATAPATH__abc_16259_n10119_bF_buf2), .B(\bus_in[22] ), .Y(AES_CORE_DATAPATH__abc_16259_n10186) );
  OR2X2 OR2X2_356 ( .A(AES_CORE_DATAPATH__abc_16259_n3142), .B(AES_CORE_DATAPATH__abc_16259_n2864_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n3143_1) );
  OR2X2 OR2X2_3560 ( .A(AES_CORE_DATAPATH_iv_1__23_), .B(iv_en_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n10188) );
  OR2X2 OR2X2_3561 ( .A(AES_CORE_DATAPATH__abc_16259_n10119_bF_buf1), .B(\bus_in[23] ), .Y(AES_CORE_DATAPATH__abc_16259_n10189) );
  OR2X2 OR2X2_3562 ( .A(AES_CORE_DATAPATH_iv_1__24_), .B(iv_en_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n10191) );
  OR2X2 OR2X2_3563 ( .A(AES_CORE_DATAPATH__abc_16259_n10119_bF_buf0), .B(\bus_in[24] ), .Y(AES_CORE_DATAPATH__abc_16259_n10192) );
  OR2X2 OR2X2_3564 ( .A(AES_CORE_DATAPATH_iv_1__25_), .B(iv_en_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n10194) );
  OR2X2 OR2X2_3565 ( .A(AES_CORE_DATAPATH__abc_16259_n10119_bF_buf4), .B(\bus_in[25] ), .Y(AES_CORE_DATAPATH__abc_16259_n10195) );
  OR2X2 OR2X2_3566 ( .A(AES_CORE_DATAPATH_iv_1__26_), .B(iv_en_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n10197) );
  OR2X2 OR2X2_3567 ( .A(AES_CORE_DATAPATH__abc_16259_n10119_bF_buf3), .B(\bus_in[26] ), .Y(AES_CORE_DATAPATH__abc_16259_n10198) );
  OR2X2 OR2X2_3568 ( .A(AES_CORE_DATAPATH_iv_1__27_), .B(iv_en_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n10200) );
  OR2X2 OR2X2_3569 ( .A(AES_CORE_DATAPATH__abc_16259_n10119_bF_buf2), .B(\bus_in[27] ), .Y(AES_CORE_DATAPATH__abc_16259_n10201) );
  OR2X2 OR2X2_357 ( .A(AES_CORE_DATAPATH__abc_16259_n3143_1), .B(AES_CORE_DATAPATH__abc_16259_n3141_1), .Y(AES_CORE_DATAPATH__abc_16259_n3144) );
  OR2X2 OR2X2_3570 ( .A(AES_CORE_DATAPATH_iv_1__28_), .B(iv_en_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n10203) );
  OR2X2 OR2X2_3571 ( .A(AES_CORE_DATAPATH__abc_16259_n10119_bF_buf1), .B(\bus_in[28] ), .Y(AES_CORE_DATAPATH__abc_16259_n10204) );
  OR2X2 OR2X2_3572 ( .A(AES_CORE_DATAPATH_iv_1__29_), .B(iv_en_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n10206) );
  OR2X2 OR2X2_3573 ( .A(AES_CORE_DATAPATH__abc_16259_n10119_bF_buf0), .B(\bus_in[29] ), .Y(AES_CORE_DATAPATH__abc_16259_n10207) );
  OR2X2 OR2X2_3574 ( .A(AES_CORE_DATAPATH_iv_1__30_), .B(iv_en_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n10209) );
  OR2X2 OR2X2_3575 ( .A(AES_CORE_DATAPATH__abc_16259_n10119_bF_buf4), .B(\bus_in[30] ), .Y(AES_CORE_DATAPATH__abc_16259_n10210) );
  OR2X2 OR2X2_3576 ( .A(AES_CORE_DATAPATH_iv_1__31_), .B(iv_en_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n10212) );
  OR2X2 OR2X2_3577 ( .A(AES_CORE_DATAPATH__abc_16259_n10119_bF_buf3), .B(\bus_in[31] ), .Y(AES_CORE_DATAPATH__abc_16259_n10213) );
  OR2X2 OR2X2_3578 ( .A(AES_CORE_DATAPATH__abc_16259_n10215), .B(AES_CORE_DATAPATH__abc_16259_n10216), .Y(AES_CORE_DATAPATH__abc_16259_n10217) );
  OR2X2 OR2X2_3579 ( .A(AES_CORE_DATAPATH__abc_16259_n10220), .B(AES_CORE_DATAPATH__abc_16259_n10219), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__0_) );
  OR2X2 OR2X2_358 ( .A(AES_CORE_DATAPATH__abc_16259_n3146), .B(AES_CORE_DATAPATH__abc_16259_n3145), .Y(AES_CORE_DATAPATH__abc_16259_n3147) );
  OR2X2 OR2X2_3580 ( .A(AES_CORE_DATAPATH__abc_16259_n10223), .B(AES_CORE_DATAPATH__abc_16259_n10222), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__1_) );
  OR2X2 OR2X2_3581 ( .A(AES_CORE_DATAPATH__abc_16259_n10226), .B(AES_CORE_DATAPATH__abc_16259_n10225), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__2_) );
  OR2X2 OR2X2_3582 ( .A(AES_CORE_DATAPATH__abc_16259_n10229), .B(AES_CORE_DATAPATH__abc_16259_n10228), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__3_) );
  OR2X2 OR2X2_3583 ( .A(AES_CORE_DATAPATH__abc_16259_n10232), .B(AES_CORE_DATAPATH__abc_16259_n10231), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__4_) );
  OR2X2 OR2X2_3584 ( .A(AES_CORE_DATAPATH__abc_16259_n10235), .B(AES_CORE_DATAPATH__abc_16259_n10234), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__5_) );
  OR2X2 OR2X2_3585 ( .A(AES_CORE_DATAPATH__abc_16259_n10238), .B(AES_CORE_DATAPATH__abc_16259_n10237), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__6_) );
  OR2X2 OR2X2_3586 ( .A(AES_CORE_DATAPATH__abc_16259_n10241), .B(AES_CORE_DATAPATH__abc_16259_n10240), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__7_) );
  OR2X2 OR2X2_3587 ( .A(AES_CORE_DATAPATH__abc_16259_n10244), .B(AES_CORE_DATAPATH__abc_16259_n10243), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__8_) );
  OR2X2 OR2X2_3588 ( .A(AES_CORE_DATAPATH__abc_16259_n10247), .B(AES_CORE_DATAPATH__abc_16259_n10246), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__9_) );
  OR2X2 OR2X2_3589 ( .A(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1_0__10_), .Y(AES_CORE_DATAPATH__abc_16259_n10251) );
  OR2X2 OR2X2_359 ( .A(AES_CORE_DATAPATH__abc_16259_n3147), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n3148_1) );
  OR2X2 OR2X2_3590 ( .A(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf1), .B(AES_CORE_DATAPATH_bkp_1_0__11_), .Y(AES_CORE_DATAPATH__abc_16259_n10255) );
  OR2X2 OR2X2_3591 ( .A(AES_CORE_DATAPATH__abc_16259_n10258), .B(AES_CORE_DATAPATH__abc_16259_n10257), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__12_) );
  OR2X2 OR2X2_3592 ( .A(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf6), .B(AES_CORE_DATAPATH_bkp_1_0__13_), .Y(AES_CORE_DATAPATH__abc_16259_n10262) );
  OR2X2 OR2X2_3593 ( .A(AES_CORE_DATAPATH__abc_16259_n10265), .B(AES_CORE_DATAPATH__abc_16259_n10264), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__14_) );
  OR2X2 OR2X2_3594 ( .A(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1_0__15_), .Y(AES_CORE_DATAPATH__abc_16259_n10269) );
  OR2X2 OR2X2_3595 ( .A(AES_CORE_DATAPATH__abc_16259_n10272), .B(AES_CORE_DATAPATH__abc_16259_n10271), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__16_) );
  OR2X2 OR2X2_3596 ( .A(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf0), .B(AES_CORE_DATAPATH_bkp_1_0__17_), .Y(AES_CORE_DATAPATH__abc_16259_n10276) );
  OR2X2 OR2X2_3597 ( .A(AES_CORE_DATAPATH__abc_16259_n10279), .B(AES_CORE_DATAPATH__abc_16259_n10278), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__18_) );
  OR2X2 OR2X2_3598 ( .A(AES_CORE_DATAPATH__abc_16259_n10282), .B(AES_CORE_DATAPATH__abc_16259_n10281), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__19_) );
  OR2X2 OR2X2_3599 ( .A(AES_CORE_DATAPATH__abc_16259_n10285), .B(AES_CORE_DATAPATH__abc_16259_n10284), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__20_) );
  OR2X2 OR2X2_36 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n178), .B(AES_CORE_CONTROL_UNIT_rd_count_3_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n185) );
  OR2X2 OR2X2_360 ( .A(AES_CORE_DATAPATH__abc_16259_n3150), .B(AES_CORE_DATAPATH__abc_16259_n3151), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_7_) );
  OR2X2 OR2X2_3600 ( .A(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1_0__21_), .Y(AES_CORE_DATAPATH__abc_16259_n10289) );
  OR2X2 OR2X2_3601 ( .A(AES_CORE_DATAPATH__abc_16259_n10292), .B(AES_CORE_DATAPATH__abc_16259_n10291), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__22_) );
  OR2X2 OR2X2_3602 ( .A(AES_CORE_DATAPATH__abc_16259_n10295), .B(AES_CORE_DATAPATH__abc_16259_n10294), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__23_) );
  OR2X2 OR2X2_3603 ( .A(AES_CORE_DATAPATH__abc_16259_n10298), .B(AES_CORE_DATAPATH__abc_16259_n10297), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__24_) );
  OR2X2 OR2X2_3604 ( .A(AES_CORE_DATAPATH__abc_16259_n10301), .B(AES_CORE_DATAPATH__abc_16259_n10300), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__25_) );
  OR2X2 OR2X2_3605 ( .A(AES_CORE_DATAPATH__abc_16259_n10304), .B(AES_CORE_DATAPATH__abc_16259_n10303), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__26_) );
  OR2X2 OR2X2_3606 ( .A(AES_CORE_DATAPATH__abc_16259_n10307), .B(AES_CORE_DATAPATH__abc_16259_n10306), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__27_) );
  OR2X2 OR2X2_3607 ( .A(AES_CORE_DATAPATH__abc_16259_n10310), .B(AES_CORE_DATAPATH__abc_16259_n10309), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__28_) );
  OR2X2 OR2X2_3608 ( .A(AES_CORE_DATAPATH__abc_16259_n10313), .B(AES_CORE_DATAPATH__abc_16259_n10312), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__29_) );
  OR2X2 OR2X2_3609 ( .A(AES_CORE_DATAPATH__abc_16259_n10316), .B(AES_CORE_DATAPATH__abc_16259_n10315), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__30_) );
  OR2X2 OR2X2_361 ( .A(AES_CORE_DATAPATH__abc_16259_n2774_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n3153), .Y(AES_CORE_DATAPATH__abc_16259_n3154_1) );
  OR2X2 OR2X2_3610 ( .A(AES_CORE_DATAPATH__abc_16259_n10319), .B(AES_CORE_DATAPATH__abc_16259_n10318), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__31_) );
  OR2X2 OR2X2_3611 ( .A(AES_CORE_DATAPATH__abc_16259_n8225), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n10321) );
  OR2X2 OR2X2_3612 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1_0__0_), .Y(AES_CORE_DATAPATH__abc_16259_n10322) );
  OR2X2 OR2X2_3613 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n8608), .Y(AES_CORE_DATAPATH__abc_16259_n10325) );
  OR2X2 OR2X2_3614 ( .A(AES_CORE_DATAPATH__abc_16259_n10324), .B(AES_CORE_DATAPATH__abc_16259_n10325), .Y(AES_CORE_DATAPATH__abc_16259_n10326) );
  OR2X2 OR2X2_3615 ( .A(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf0), .B(AES_CORE_DATAPATH_bkp_0__0_), .Y(AES_CORE_DATAPATH__abc_16259_n10327) );
  OR2X2 OR2X2_3616 ( .A(AES_CORE_DATAPATH__abc_16259_n8233), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n10329) );
  OR2X2 OR2X2_3617 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf2), .B(AES_CORE_DATAPATH_bkp_1_0__1_), .Y(AES_CORE_DATAPATH__abc_16259_n10330) );
  OR2X2 OR2X2_3618 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n8617), .Y(AES_CORE_DATAPATH__abc_16259_n10333) );
  OR2X2 OR2X2_3619 ( .A(AES_CORE_DATAPATH__abc_16259_n10332), .B(AES_CORE_DATAPATH__abc_16259_n10333), .Y(AES_CORE_DATAPATH__abc_16259_n10334) );
  OR2X2 OR2X2_362 ( .A(AES_CORE_DATAPATH__abc_16259_n2778_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n3155), .Y(AES_CORE_DATAPATH__abc_16259_n3156_1) );
  OR2X2 OR2X2_3620 ( .A(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf7), .B(AES_CORE_DATAPATH_bkp_0__1_), .Y(AES_CORE_DATAPATH__abc_16259_n10335) );
  OR2X2 OR2X2_3621 ( .A(AES_CORE_DATAPATH__abc_16259_n8241), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf9), .Y(AES_CORE_DATAPATH__abc_16259_n10337) );
  OR2X2 OR2X2_3622 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf1), .B(AES_CORE_DATAPATH_bkp_1_0__2_), .Y(AES_CORE_DATAPATH__abc_16259_n10338) );
  OR2X2 OR2X2_3623 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf6), .B(AES_CORE_DATAPATH__abc_16259_n8626), .Y(AES_CORE_DATAPATH__abc_16259_n10341) );
  OR2X2 OR2X2_3624 ( .A(AES_CORE_DATAPATH__abc_16259_n10340), .B(AES_CORE_DATAPATH__abc_16259_n10341), .Y(AES_CORE_DATAPATH__abc_16259_n10342) );
  OR2X2 OR2X2_3625 ( .A(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf6), .B(AES_CORE_DATAPATH_bkp_0__2_), .Y(AES_CORE_DATAPATH__abc_16259_n10343) );
  OR2X2 OR2X2_3626 ( .A(AES_CORE_DATAPATH__abc_16259_n8249), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf8), .Y(AES_CORE_DATAPATH__abc_16259_n10345) );
  OR2X2 OR2X2_3627 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf0), .B(AES_CORE_DATAPATH_bkp_1_0__3_), .Y(AES_CORE_DATAPATH__abc_16259_n10346) );
  OR2X2 OR2X2_3628 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf5), .B(AES_CORE_DATAPATH__abc_16259_n8635), .Y(AES_CORE_DATAPATH__abc_16259_n10349) );
  OR2X2 OR2X2_3629 ( .A(AES_CORE_DATAPATH__abc_16259_n10348), .B(AES_CORE_DATAPATH__abc_16259_n10349), .Y(AES_CORE_DATAPATH__abc_16259_n10350) );
  OR2X2 OR2X2_363 ( .A(AES_CORE_DATAPATH__abc_16259_n3159), .B(AES_CORE_DATAPATH__abc_16259_n3160), .Y(AES_CORE_DATAPATH__abc_16259_n3161) );
  OR2X2 OR2X2_3630 ( .A(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf5), .B(AES_CORE_DATAPATH_bkp_0__3_), .Y(AES_CORE_DATAPATH__abc_16259_n10351) );
  OR2X2 OR2X2_3631 ( .A(AES_CORE_DATAPATH__abc_16259_n8257), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n10353) );
  OR2X2 OR2X2_3632 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf11), .B(AES_CORE_DATAPATH_bkp_1_0__4_), .Y(AES_CORE_DATAPATH__abc_16259_n10354) );
  OR2X2 OR2X2_3633 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n8644), .Y(AES_CORE_DATAPATH__abc_16259_n10357) );
  OR2X2 OR2X2_3634 ( .A(AES_CORE_DATAPATH__abc_16259_n10356), .B(AES_CORE_DATAPATH__abc_16259_n10357), .Y(AES_CORE_DATAPATH__abc_16259_n10358) );
  OR2X2 OR2X2_3635 ( .A(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf4), .B(AES_CORE_DATAPATH_bkp_0__4_), .Y(AES_CORE_DATAPATH__abc_16259_n10359) );
  OR2X2 OR2X2_3636 ( .A(AES_CORE_DATAPATH__abc_16259_n8265), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n10361) );
  OR2X2 OR2X2_3637 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf10), .B(AES_CORE_DATAPATH_bkp_1_0__5_), .Y(AES_CORE_DATAPATH__abc_16259_n10362) );
  OR2X2 OR2X2_3638 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n8653), .Y(AES_CORE_DATAPATH__abc_16259_n10365) );
  OR2X2 OR2X2_3639 ( .A(AES_CORE_DATAPATH__abc_16259_n10364), .B(AES_CORE_DATAPATH__abc_16259_n10365), .Y(AES_CORE_DATAPATH__abc_16259_n10366) );
  OR2X2 OR2X2_364 ( .A(AES_CORE_DATAPATH__abc_16259_n3161), .B(AES_CORE_DATAPATH__abc_16259_n3158_1), .Y(AES_CORE_DATAPATH__abc_16259_n3162) );
  OR2X2 OR2X2_3640 ( .A(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf3), .B(AES_CORE_DATAPATH_bkp_0__5_), .Y(AES_CORE_DATAPATH__abc_16259_n10367) );
  OR2X2 OR2X2_3641 ( .A(AES_CORE_DATAPATH__abc_16259_n8273), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n10369) );
  OR2X2 OR2X2_3642 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf9), .B(AES_CORE_DATAPATH_bkp_1_0__6_), .Y(AES_CORE_DATAPATH__abc_16259_n10370) );
  OR2X2 OR2X2_3643 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n8662), .Y(AES_CORE_DATAPATH__abc_16259_n10373) );
  OR2X2 OR2X2_3644 ( .A(AES_CORE_DATAPATH__abc_16259_n10372), .B(AES_CORE_DATAPATH__abc_16259_n10373), .Y(AES_CORE_DATAPATH__abc_16259_n10374) );
  OR2X2 OR2X2_3645 ( .A(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf2), .B(AES_CORE_DATAPATH_bkp_0__6_), .Y(AES_CORE_DATAPATH__abc_16259_n10375) );
  OR2X2 OR2X2_3646 ( .A(AES_CORE_DATAPATH__abc_16259_n8281), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n10377) );
  OR2X2 OR2X2_3647 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf8), .B(AES_CORE_DATAPATH_bkp_1_0__7_), .Y(AES_CORE_DATAPATH__abc_16259_n10378) );
  OR2X2 OR2X2_3648 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n8671), .Y(AES_CORE_DATAPATH__abc_16259_n10381) );
  OR2X2 OR2X2_3649 ( .A(AES_CORE_DATAPATH__abc_16259_n10380), .B(AES_CORE_DATAPATH__abc_16259_n10381), .Y(AES_CORE_DATAPATH__abc_16259_n10382) );
  OR2X2 OR2X2_365 ( .A(AES_CORE_DATAPATH__abc_16259_n3166), .B(AES_CORE_DATAPATH__abc_16259_n2826_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n3167) );
  OR2X2 OR2X2_3650 ( .A(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf1), .B(AES_CORE_DATAPATH_bkp_0__7_), .Y(AES_CORE_DATAPATH__abc_16259_n10383) );
  OR2X2 OR2X2_3651 ( .A(AES_CORE_DATAPATH__abc_16259_n8289), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n10385) );
  OR2X2 OR2X2_3652 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf7), .B(AES_CORE_DATAPATH_bkp_1_0__8_), .Y(AES_CORE_DATAPATH__abc_16259_n10386) );
  OR2X2 OR2X2_3653 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n8680), .Y(AES_CORE_DATAPATH__abc_16259_n10389) );
  OR2X2 OR2X2_3654 ( .A(AES_CORE_DATAPATH__abc_16259_n10388), .B(AES_CORE_DATAPATH__abc_16259_n10389), .Y(AES_CORE_DATAPATH__abc_16259_n10390) );
  OR2X2 OR2X2_3655 ( .A(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf0), .B(AES_CORE_DATAPATH_bkp_0__8_), .Y(AES_CORE_DATAPATH__abc_16259_n10391) );
  OR2X2 OR2X2_3656 ( .A(AES_CORE_DATAPATH__abc_16259_n8297), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n10393) );
  OR2X2 OR2X2_3657 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf6), .B(AES_CORE_DATAPATH_bkp_1_0__9_), .Y(AES_CORE_DATAPATH__abc_16259_n10394) );
  OR2X2 OR2X2_3658 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf6), .B(AES_CORE_DATAPATH__abc_16259_n8689), .Y(AES_CORE_DATAPATH__abc_16259_n10397) );
  OR2X2 OR2X2_3659 ( .A(AES_CORE_DATAPATH__abc_16259_n10396), .B(AES_CORE_DATAPATH__abc_16259_n10397), .Y(AES_CORE_DATAPATH__abc_16259_n10398) );
  OR2X2 OR2X2_366 ( .A(AES_CORE_DATAPATH__abc_16259_n3168), .B(AES_CORE_DATAPATH__abc_16259_n3169), .Y(AES_CORE_DATAPATH__abc_16259_n3170_1) );
  OR2X2 OR2X2_3660 ( .A(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf7), .B(AES_CORE_DATAPATH_bkp_0__9_), .Y(AES_CORE_DATAPATH__abc_16259_n10399) );
  OR2X2 OR2X2_3661 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf4), .B(AES_CORE_DATAPATH_bkp_1_0__10_), .Y(AES_CORE_DATAPATH__abc_16259_n10403) );
  OR2X2 OR2X2_3662 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf5), .B(AES_CORE_DATAPATH__abc_16259_n8699), .Y(AES_CORE_DATAPATH__abc_16259_n10406) );
  OR2X2 OR2X2_3663 ( .A(AES_CORE_DATAPATH__abc_16259_n10405), .B(AES_CORE_DATAPATH__abc_16259_n10406), .Y(AES_CORE_DATAPATH__abc_16259_n10407) );
  OR2X2 OR2X2_3664 ( .A(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf6), .B(AES_CORE_DATAPATH_bkp_0__10_), .Y(AES_CORE_DATAPATH__abc_16259_n10408) );
  OR2X2 OR2X2_3665 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf2), .B(AES_CORE_DATAPATH_bkp_1_0__11_), .Y(AES_CORE_DATAPATH__abc_16259_n10412) );
  OR2X2 OR2X2_3666 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n8709), .Y(AES_CORE_DATAPATH__abc_16259_n10415) );
  OR2X2 OR2X2_3667 ( .A(AES_CORE_DATAPATH__abc_16259_n10414), .B(AES_CORE_DATAPATH__abc_16259_n10415), .Y(AES_CORE_DATAPATH__abc_16259_n10416) );
  OR2X2 OR2X2_3668 ( .A(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf5), .B(AES_CORE_DATAPATH_bkp_0__11_), .Y(AES_CORE_DATAPATH__abc_16259_n10417) );
  OR2X2 OR2X2_3669 ( .A(AES_CORE_DATAPATH__abc_16259_n8327), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n10419) );
  OR2X2 OR2X2_367 ( .A(AES_CORE_DATAPATH__abc_16259_n3170_1), .B(AES_CORE_DATAPATH__abc_16259_n3167), .Y(AES_CORE_DATAPATH__abc_16259_n3171) );
  OR2X2 OR2X2_3670 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf1), .B(AES_CORE_DATAPATH_bkp_1_0__12_), .Y(AES_CORE_DATAPATH__abc_16259_n10420) );
  OR2X2 OR2X2_3671 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n8718), .Y(AES_CORE_DATAPATH__abc_16259_n10423) );
  OR2X2 OR2X2_3672 ( .A(AES_CORE_DATAPATH__abc_16259_n10422), .B(AES_CORE_DATAPATH__abc_16259_n10423), .Y(AES_CORE_DATAPATH__abc_16259_n10424) );
  OR2X2 OR2X2_3673 ( .A(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf4), .B(AES_CORE_DATAPATH_bkp_0__12_), .Y(AES_CORE_DATAPATH__abc_16259_n10425) );
  OR2X2 OR2X2_3674 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf11), .B(AES_CORE_DATAPATH_bkp_1_0__13_), .Y(AES_CORE_DATAPATH__abc_16259_n10429) );
  OR2X2 OR2X2_3675 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n8728), .Y(AES_CORE_DATAPATH__abc_16259_n10432) );
  OR2X2 OR2X2_3676 ( .A(AES_CORE_DATAPATH__abc_16259_n10431), .B(AES_CORE_DATAPATH__abc_16259_n10432), .Y(AES_CORE_DATAPATH__abc_16259_n10433) );
  OR2X2 OR2X2_3677 ( .A(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf3), .B(AES_CORE_DATAPATH_bkp_0__13_), .Y(AES_CORE_DATAPATH__abc_16259_n10434) );
  OR2X2 OR2X2_3678 ( .A(AES_CORE_DATAPATH__abc_16259_n8346), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n10436) );
  OR2X2 OR2X2_3679 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf10), .B(AES_CORE_DATAPATH_bkp_1_0__14_), .Y(AES_CORE_DATAPATH__abc_16259_n10437) );
  OR2X2 OR2X2_368 ( .A(AES_CORE_DATAPATH__abc_16259_n2841_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__8_), .Y(AES_CORE_DATAPATH__abc_16259_n3172_1) );
  OR2X2 OR2X2_3680 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n8737), .Y(AES_CORE_DATAPATH__abc_16259_n10440) );
  OR2X2 OR2X2_3681 ( .A(AES_CORE_DATAPATH__abc_16259_n10439), .B(AES_CORE_DATAPATH__abc_16259_n10440), .Y(AES_CORE_DATAPATH__abc_16259_n10441) );
  OR2X2 OR2X2_3682 ( .A(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf2), .B(AES_CORE_DATAPATH_bkp_0__14_), .Y(AES_CORE_DATAPATH__abc_16259_n10442) );
  OR2X2 OR2X2_3683 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf8), .B(AES_CORE_DATAPATH_bkp_1_0__15_), .Y(AES_CORE_DATAPATH__abc_16259_n10446) );
  OR2X2 OR2X2_3684 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n8747), .Y(AES_CORE_DATAPATH__abc_16259_n10449) );
  OR2X2 OR2X2_3685 ( .A(AES_CORE_DATAPATH__abc_16259_n10448), .B(AES_CORE_DATAPATH__abc_16259_n10449), .Y(AES_CORE_DATAPATH__abc_16259_n10450) );
  OR2X2 OR2X2_3686 ( .A(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf1), .B(AES_CORE_DATAPATH_bkp_0__15_), .Y(AES_CORE_DATAPATH__abc_16259_n10451) );
  OR2X2 OR2X2_3687 ( .A(AES_CORE_DATAPATH__abc_16259_n8365), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf9), .Y(AES_CORE_DATAPATH__abc_16259_n10453) );
  OR2X2 OR2X2_3688 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf7), .B(AES_CORE_DATAPATH_bkp_1_0__16_), .Y(AES_CORE_DATAPATH__abc_16259_n10454) );
  OR2X2 OR2X2_3689 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf6), .B(AES_CORE_DATAPATH__abc_16259_n8756), .Y(AES_CORE_DATAPATH__abc_16259_n10457) );
  OR2X2 OR2X2_369 ( .A(AES_CORE_DATAPATH__abc_16259_n3164), .B(AES_CORE_DATAPATH__abc_16259_n2853_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n3174) );
  OR2X2 OR2X2_3690 ( .A(AES_CORE_DATAPATH__abc_16259_n10456), .B(AES_CORE_DATAPATH__abc_16259_n10457), .Y(AES_CORE_DATAPATH__abc_16259_n10458) );
  OR2X2 OR2X2_3691 ( .A(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf0), .B(AES_CORE_DATAPATH_bkp_0__16_), .Y(AES_CORE_DATAPATH__abc_16259_n10459) );
  OR2X2 OR2X2_3692 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf5), .B(AES_CORE_DATAPATH_bkp_1_0__17_), .Y(AES_CORE_DATAPATH__abc_16259_n10463) );
  OR2X2 OR2X2_3693 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf5), .B(AES_CORE_DATAPATH__abc_16259_n8766), .Y(AES_CORE_DATAPATH__abc_16259_n10466) );
  OR2X2 OR2X2_3694 ( .A(AES_CORE_DATAPATH__abc_16259_n10465), .B(AES_CORE_DATAPATH__abc_16259_n10466), .Y(AES_CORE_DATAPATH__abc_16259_n10467) );
  OR2X2 OR2X2_3695 ( .A(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf7), .B(AES_CORE_DATAPATH_bkp_0__17_), .Y(AES_CORE_DATAPATH__abc_16259_n10468) );
  OR2X2 OR2X2_3696 ( .A(AES_CORE_DATAPATH__abc_16259_n8384), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf8), .Y(AES_CORE_DATAPATH__abc_16259_n10470) );
  OR2X2 OR2X2_3697 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf4), .B(AES_CORE_DATAPATH_bkp_1_0__18_), .Y(AES_CORE_DATAPATH__abc_16259_n10471) );
  OR2X2 OR2X2_3698 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n8775), .Y(AES_CORE_DATAPATH__abc_16259_n10474) );
  OR2X2 OR2X2_3699 ( .A(AES_CORE_DATAPATH__abc_16259_n10473), .B(AES_CORE_DATAPATH__abc_16259_n10474), .Y(AES_CORE_DATAPATH__abc_16259_n10475) );
  OR2X2 OR2X2_37 ( .A(AES_CORE_CONTROL_UNIT_state_14_), .B(AES_CORE_CONTROL_UNIT_state_1_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n188) );
  OR2X2 OR2X2_370 ( .A(AES_CORE_DATAPATH__abc_16259_n3175), .B(AES_CORE_DATAPATH__abc_16259_n3176), .Y(AES_CORE_DATAPATH__abc_16259_n3177_1) );
  OR2X2 OR2X2_3700 ( .A(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf6), .B(AES_CORE_DATAPATH_bkp_0__18_), .Y(AES_CORE_DATAPATH__abc_16259_n10476) );
  OR2X2 OR2X2_3701 ( .A(AES_CORE_DATAPATH__abc_16259_n8392), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n10478) );
  OR2X2 OR2X2_3702 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1_0__19_), .Y(AES_CORE_DATAPATH__abc_16259_n10479) );
  OR2X2 OR2X2_3703 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n8784), .Y(AES_CORE_DATAPATH__abc_16259_n10482) );
  OR2X2 OR2X2_3704 ( .A(AES_CORE_DATAPATH__abc_16259_n10481), .B(AES_CORE_DATAPATH__abc_16259_n10482), .Y(AES_CORE_DATAPATH__abc_16259_n10483) );
  OR2X2 OR2X2_3705 ( .A(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf5), .B(AES_CORE_DATAPATH_bkp_0__19_), .Y(AES_CORE_DATAPATH__abc_16259_n10484) );
  OR2X2 OR2X2_3706 ( .A(AES_CORE_DATAPATH__abc_16259_n8400), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n10486) );
  OR2X2 OR2X2_3707 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf2), .B(AES_CORE_DATAPATH_bkp_1_0__20_), .Y(AES_CORE_DATAPATH__abc_16259_n10487) );
  OR2X2 OR2X2_3708 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n8793), .Y(AES_CORE_DATAPATH__abc_16259_n10490) );
  OR2X2 OR2X2_3709 ( .A(AES_CORE_DATAPATH__abc_16259_n10489), .B(AES_CORE_DATAPATH__abc_16259_n10490), .Y(AES_CORE_DATAPATH__abc_16259_n10491) );
  OR2X2 OR2X2_371 ( .A(_auto_iopadmap_cc_313_execute_26949_8_), .B(AES_CORE_DATAPATH__abc_16259_n3179), .Y(AES_CORE_DATAPATH__abc_16259_n3180) );
  OR2X2 OR2X2_3710 ( .A(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf4), .B(AES_CORE_DATAPATH_bkp_0__20_), .Y(AES_CORE_DATAPATH__abc_16259_n10492) );
  OR2X2 OR2X2_3711 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf0), .B(AES_CORE_DATAPATH_bkp_1_0__21_), .Y(AES_CORE_DATAPATH__abc_16259_n10496) );
  OR2X2 OR2X2_3712 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n8803), .Y(AES_CORE_DATAPATH__abc_16259_n10499) );
  OR2X2 OR2X2_3713 ( .A(AES_CORE_DATAPATH__abc_16259_n10498), .B(AES_CORE_DATAPATH__abc_16259_n10499), .Y(AES_CORE_DATAPATH__abc_16259_n10500) );
  OR2X2 OR2X2_3714 ( .A(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf3), .B(AES_CORE_DATAPATH_bkp_0__21_), .Y(AES_CORE_DATAPATH__abc_16259_n10501) );
  OR2X2 OR2X2_3715 ( .A(AES_CORE_DATAPATH__abc_16259_n8419), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n10503) );
  OR2X2 OR2X2_3716 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf11), .B(AES_CORE_DATAPATH_bkp_1_0__22_), .Y(AES_CORE_DATAPATH__abc_16259_n10504) );
  OR2X2 OR2X2_3717 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n8812), .Y(AES_CORE_DATAPATH__abc_16259_n10507) );
  OR2X2 OR2X2_3718 ( .A(AES_CORE_DATAPATH__abc_16259_n10506), .B(AES_CORE_DATAPATH__abc_16259_n10507), .Y(AES_CORE_DATAPATH__abc_16259_n10508) );
  OR2X2 OR2X2_3719 ( .A(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf2), .B(AES_CORE_DATAPATH_bkp_0__22_), .Y(AES_CORE_DATAPATH__abc_16259_n10509) );
  OR2X2 OR2X2_372 ( .A(AES_CORE_DATAPATH__abc_16259_n3182), .B(AES_CORE_DATAPATH__abc_16259_n2864_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n3183_1) );
  OR2X2 OR2X2_3720 ( .A(AES_CORE_DATAPATH__abc_16259_n8427), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n10511) );
  OR2X2 OR2X2_3721 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf10), .B(AES_CORE_DATAPATH_bkp_1_0__23_), .Y(AES_CORE_DATAPATH__abc_16259_n10512) );
  OR2X2 OR2X2_3722 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf6), .B(AES_CORE_DATAPATH__abc_16259_n8821), .Y(AES_CORE_DATAPATH__abc_16259_n10515) );
  OR2X2 OR2X2_3723 ( .A(AES_CORE_DATAPATH__abc_16259_n10514), .B(AES_CORE_DATAPATH__abc_16259_n10515), .Y(AES_CORE_DATAPATH__abc_16259_n10516) );
  OR2X2 OR2X2_3724 ( .A(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf1), .B(AES_CORE_DATAPATH_bkp_0__23_), .Y(AES_CORE_DATAPATH__abc_16259_n10517) );
  OR2X2 OR2X2_3725 ( .A(AES_CORE_DATAPATH__abc_16259_n8435), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n10519) );
  OR2X2 OR2X2_3726 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf9), .B(AES_CORE_DATAPATH_bkp_1_0__24_), .Y(AES_CORE_DATAPATH__abc_16259_n10520) );
  OR2X2 OR2X2_3727 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf5), .B(AES_CORE_DATAPATH__abc_16259_n8830), .Y(AES_CORE_DATAPATH__abc_16259_n10523) );
  OR2X2 OR2X2_3728 ( .A(AES_CORE_DATAPATH__abc_16259_n10522), .B(AES_CORE_DATAPATH__abc_16259_n10523), .Y(AES_CORE_DATAPATH__abc_16259_n10524) );
  OR2X2 OR2X2_3729 ( .A(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf0), .B(AES_CORE_DATAPATH_bkp_0__24_), .Y(AES_CORE_DATAPATH__abc_16259_n10525) );
  OR2X2 OR2X2_373 ( .A(AES_CORE_DATAPATH__abc_16259_n3183_1), .B(AES_CORE_DATAPATH__abc_16259_n3181_1), .Y(AES_CORE_DATAPATH__abc_16259_n3184) );
  OR2X2 OR2X2_3730 ( .A(AES_CORE_DATAPATH__abc_16259_n8443), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n10527) );
  OR2X2 OR2X2_3731 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf8), .B(AES_CORE_DATAPATH_bkp_1_0__25_), .Y(AES_CORE_DATAPATH__abc_16259_n10528) );
  OR2X2 OR2X2_3732 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n8839), .Y(AES_CORE_DATAPATH__abc_16259_n10531) );
  OR2X2 OR2X2_3733 ( .A(AES_CORE_DATAPATH__abc_16259_n10530), .B(AES_CORE_DATAPATH__abc_16259_n10531), .Y(AES_CORE_DATAPATH__abc_16259_n10532) );
  OR2X2 OR2X2_3734 ( .A(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf7), .B(AES_CORE_DATAPATH_bkp_0__25_), .Y(AES_CORE_DATAPATH__abc_16259_n10533) );
  OR2X2 OR2X2_3735 ( .A(AES_CORE_DATAPATH__abc_16259_n8451), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n10535) );
  OR2X2 OR2X2_3736 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf7), .B(AES_CORE_DATAPATH_bkp_1_0__26_), .Y(AES_CORE_DATAPATH__abc_16259_n10536) );
  OR2X2 OR2X2_3737 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n8848), .Y(AES_CORE_DATAPATH__abc_16259_n10539) );
  OR2X2 OR2X2_3738 ( .A(AES_CORE_DATAPATH__abc_16259_n10538), .B(AES_CORE_DATAPATH__abc_16259_n10539), .Y(AES_CORE_DATAPATH__abc_16259_n10540) );
  OR2X2 OR2X2_3739 ( .A(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf6), .B(AES_CORE_DATAPATH_bkp_0__26_), .Y(AES_CORE_DATAPATH__abc_16259_n10541) );
  OR2X2 OR2X2_374 ( .A(AES_CORE_DATAPATH__abc_16259_n3186), .B(AES_CORE_DATAPATH__abc_16259_n3185_1), .Y(AES_CORE_DATAPATH__abc_16259_n3187_1) );
  OR2X2 OR2X2_3740 ( .A(AES_CORE_DATAPATH__abc_16259_n8459), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n10543) );
  OR2X2 OR2X2_3741 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf6), .B(AES_CORE_DATAPATH_bkp_1_0__27_), .Y(AES_CORE_DATAPATH__abc_16259_n10544) );
  OR2X2 OR2X2_3742 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n8857), .Y(AES_CORE_DATAPATH__abc_16259_n10547) );
  OR2X2 OR2X2_3743 ( .A(AES_CORE_DATAPATH__abc_16259_n10546), .B(AES_CORE_DATAPATH__abc_16259_n10547), .Y(AES_CORE_DATAPATH__abc_16259_n10548) );
  OR2X2 OR2X2_3744 ( .A(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf5), .B(AES_CORE_DATAPATH_bkp_0__27_), .Y(AES_CORE_DATAPATH__abc_16259_n10549) );
  OR2X2 OR2X2_3745 ( .A(AES_CORE_DATAPATH__abc_16259_n8467), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf9), .Y(AES_CORE_DATAPATH__abc_16259_n10551) );
  OR2X2 OR2X2_3746 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf5), .B(AES_CORE_DATAPATH_bkp_1_0__28_), .Y(AES_CORE_DATAPATH__abc_16259_n10552) );
  OR2X2 OR2X2_3747 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n8866), .Y(AES_CORE_DATAPATH__abc_16259_n10555) );
  OR2X2 OR2X2_3748 ( .A(AES_CORE_DATAPATH__abc_16259_n10554), .B(AES_CORE_DATAPATH__abc_16259_n10555), .Y(AES_CORE_DATAPATH__abc_16259_n10556) );
  OR2X2 OR2X2_3749 ( .A(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf4), .B(AES_CORE_DATAPATH_bkp_0__28_), .Y(AES_CORE_DATAPATH__abc_16259_n10557) );
  OR2X2 OR2X2_375 ( .A(AES_CORE_DATAPATH__abc_16259_n3187_1), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n3188) );
  OR2X2 OR2X2_3750 ( .A(AES_CORE_DATAPATH__abc_16259_n8475), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf8), .Y(AES_CORE_DATAPATH__abc_16259_n10559) );
  OR2X2 OR2X2_3751 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf4), .B(AES_CORE_DATAPATH_bkp_1_0__29_), .Y(AES_CORE_DATAPATH__abc_16259_n10560) );
  OR2X2 OR2X2_3752 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n8875), .Y(AES_CORE_DATAPATH__abc_16259_n10563) );
  OR2X2 OR2X2_3753 ( .A(AES_CORE_DATAPATH__abc_16259_n10562), .B(AES_CORE_DATAPATH__abc_16259_n10563), .Y(AES_CORE_DATAPATH__abc_16259_n10564) );
  OR2X2 OR2X2_3754 ( .A(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf3), .B(AES_CORE_DATAPATH_bkp_0__29_), .Y(AES_CORE_DATAPATH__abc_16259_n10565) );
  OR2X2 OR2X2_3755 ( .A(AES_CORE_DATAPATH__abc_16259_n8483), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n10567) );
  OR2X2 OR2X2_3756 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf3), .B(AES_CORE_DATAPATH_bkp_1_0__30_), .Y(AES_CORE_DATAPATH__abc_16259_n10568) );
  OR2X2 OR2X2_3757 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf6), .B(AES_CORE_DATAPATH__abc_16259_n8884), .Y(AES_CORE_DATAPATH__abc_16259_n10571) );
  OR2X2 OR2X2_3758 ( .A(AES_CORE_DATAPATH__abc_16259_n10570), .B(AES_CORE_DATAPATH__abc_16259_n10571), .Y(AES_CORE_DATAPATH__abc_16259_n10572) );
  OR2X2 OR2X2_3759 ( .A(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf2), .B(AES_CORE_DATAPATH_bkp_0__30_), .Y(AES_CORE_DATAPATH__abc_16259_n10573) );
  OR2X2 OR2X2_376 ( .A(AES_CORE_DATAPATH__abc_16259_n3190), .B(AES_CORE_DATAPATH__abc_16259_n3191), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_8_) );
  OR2X2 OR2X2_3760 ( .A(AES_CORE_DATAPATH__abc_16259_n8491), .B(AES_CORE_DATAPATH__abc_16259_n8603_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n10575) );
  OR2X2 OR2X2_3761 ( .A(AES_CORE_DATAPATH__abc_16259_n8496_bF_buf2), .B(AES_CORE_DATAPATH_bkp_1_0__31_), .Y(AES_CORE_DATAPATH__abc_16259_n10576) );
  OR2X2 OR2X2_3762 ( .A(AES_CORE_DATAPATH__abc_16259_n10218_bF_buf5), .B(AES_CORE_DATAPATH__abc_16259_n8893), .Y(AES_CORE_DATAPATH__abc_16259_n10579) );
  OR2X2 OR2X2_3763 ( .A(AES_CORE_DATAPATH__abc_16259_n10578), .B(AES_CORE_DATAPATH__abc_16259_n10579), .Y(AES_CORE_DATAPATH__abc_16259_n10580) );
  OR2X2 OR2X2_3764 ( .A(AES_CORE_DATAPATH__abc_16259_n10217_bF_buf1), .B(AES_CORE_DATAPATH_bkp_0__31_), .Y(AES_CORE_DATAPATH__abc_16259_n10581) );
  OR2X2 OR2X2_3765 ( .A(AES_CORE_DATAPATH_iv_0__0_), .B(iv_en_0_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n10583) );
  OR2X2 OR2X2_3766 ( .A(AES_CORE_DATAPATH__abc_16259_n10584_bF_buf4), .B(\bus_in[0] ), .Y(AES_CORE_DATAPATH__abc_16259_n10585) );
  OR2X2 OR2X2_3767 ( .A(AES_CORE_DATAPATH_iv_0__1_), .B(iv_en_0_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n10587) );
  OR2X2 OR2X2_3768 ( .A(AES_CORE_DATAPATH__abc_16259_n10584_bF_buf3), .B(\bus_in[1] ), .Y(AES_CORE_DATAPATH__abc_16259_n10588) );
  OR2X2 OR2X2_3769 ( .A(AES_CORE_DATAPATH_iv_0__2_), .B(iv_en_0_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n10590) );
  OR2X2 OR2X2_377 ( .A(AES_CORE_DATAPATH__abc_16259_n2774_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n3193), .Y(AES_CORE_DATAPATH__abc_16259_n3194) );
  OR2X2 OR2X2_3770 ( .A(AES_CORE_DATAPATH__abc_16259_n10584_bF_buf2), .B(\bus_in[2] ), .Y(AES_CORE_DATAPATH__abc_16259_n10591) );
  OR2X2 OR2X2_3771 ( .A(AES_CORE_DATAPATH_iv_0__3_), .B(iv_en_0_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n10593) );
  OR2X2 OR2X2_3772 ( .A(AES_CORE_DATAPATH__abc_16259_n10584_bF_buf1), .B(\bus_in[3] ), .Y(AES_CORE_DATAPATH__abc_16259_n10594) );
  OR2X2 OR2X2_3773 ( .A(AES_CORE_DATAPATH_iv_0__4_), .B(iv_en_0_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n10596) );
  OR2X2 OR2X2_3774 ( .A(AES_CORE_DATAPATH__abc_16259_n10584_bF_buf0), .B(\bus_in[4] ), .Y(AES_CORE_DATAPATH__abc_16259_n10597) );
  OR2X2 OR2X2_3775 ( .A(AES_CORE_DATAPATH_iv_0__5_), .B(iv_en_0_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n10599) );
  OR2X2 OR2X2_3776 ( .A(AES_CORE_DATAPATH__abc_16259_n10584_bF_buf4), .B(\bus_in[5] ), .Y(AES_CORE_DATAPATH__abc_16259_n10600) );
  OR2X2 OR2X2_3777 ( .A(AES_CORE_DATAPATH_iv_0__6_), .B(iv_en_0_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n10602) );
  OR2X2 OR2X2_3778 ( .A(AES_CORE_DATAPATH__abc_16259_n10584_bF_buf3), .B(\bus_in[6] ), .Y(AES_CORE_DATAPATH__abc_16259_n10603) );
  OR2X2 OR2X2_3779 ( .A(AES_CORE_DATAPATH_iv_0__7_), .B(iv_en_0_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n10605) );
  OR2X2 OR2X2_378 ( .A(AES_CORE_DATAPATH__abc_16259_n2778_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n3195), .Y(AES_CORE_DATAPATH__abc_16259_n3196) );
  OR2X2 OR2X2_3780 ( .A(AES_CORE_DATAPATH__abc_16259_n10584_bF_buf2), .B(\bus_in[7] ), .Y(AES_CORE_DATAPATH__abc_16259_n10606) );
  OR2X2 OR2X2_3781 ( .A(AES_CORE_DATAPATH_iv_0__8_), .B(iv_en_0_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n10608) );
  OR2X2 OR2X2_3782 ( .A(AES_CORE_DATAPATH__abc_16259_n10584_bF_buf1), .B(\bus_in[8] ), .Y(AES_CORE_DATAPATH__abc_16259_n10609) );
  OR2X2 OR2X2_3783 ( .A(AES_CORE_DATAPATH_iv_0__9_), .B(iv_en_0_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n10611) );
  OR2X2 OR2X2_3784 ( .A(AES_CORE_DATAPATH__abc_16259_n10584_bF_buf0), .B(\bus_in[9] ), .Y(AES_CORE_DATAPATH__abc_16259_n10612) );
  OR2X2 OR2X2_3785 ( .A(AES_CORE_DATAPATH_iv_0__10_), .B(iv_en_0_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n10614) );
  OR2X2 OR2X2_3786 ( .A(AES_CORE_DATAPATH__abc_16259_n10584_bF_buf4), .B(\bus_in[10] ), .Y(AES_CORE_DATAPATH__abc_16259_n10615) );
  OR2X2 OR2X2_3787 ( .A(AES_CORE_DATAPATH_iv_0__11_), .B(iv_en_0_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n10617) );
  OR2X2 OR2X2_3788 ( .A(AES_CORE_DATAPATH__abc_16259_n10584_bF_buf3), .B(\bus_in[11] ), .Y(AES_CORE_DATAPATH__abc_16259_n10618) );
  OR2X2 OR2X2_3789 ( .A(AES_CORE_DATAPATH_iv_0__12_), .B(iv_en_0_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n10620) );
  OR2X2 OR2X2_379 ( .A(AES_CORE_DATAPATH__abc_16259_n3199_1), .B(AES_CORE_DATAPATH__abc_16259_n3200), .Y(AES_CORE_DATAPATH__abc_16259_n3201_1) );
  OR2X2 OR2X2_3790 ( .A(AES_CORE_DATAPATH__abc_16259_n10584_bF_buf2), .B(\bus_in[12] ), .Y(AES_CORE_DATAPATH__abc_16259_n10621) );
  OR2X2 OR2X2_3791 ( .A(AES_CORE_DATAPATH_iv_0__13_), .B(iv_en_0_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n10623) );
  OR2X2 OR2X2_3792 ( .A(AES_CORE_DATAPATH__abc_16259_n10584_bF_buf1), .B(\bus_in[13] ), .Y(AES_CORE_DATAPATH__abc_16259_n10624) );
  OR2X2 OR2X2_3793 ( .A(AES_CORE_DATAPATH_iv_0__14_), .B(iv_en_0_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n10626) );
  OR2X2 OR2X2_3794 ( .A(AES_CORE_DATAPATH__abc_16259_n10584_bF_buf0), .B(\bus_in[14] ), .Y(AES_CORE_DATAPATH__abc_16259_n10627) );
  OR2X2 OR2X2_3795 ( .A(AES_CORE_DATAPATH_iv_0__15_), .B(iv_en_0_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n10629) );
  OR2X2 OR2X2_3796 ( .A(AES_CORE_DATAPATH__abc_16259_n10584_bF_buf4), .B(\bus_in[15] ), .Y(AES_CORE_DATAPATH__abc_16259_n10630) );
  OR2X2 OR2X2_3797 ( .A(AES_CORE_DATAPATH_iv_0__16_), .B(iv_en_0_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n10632) );
  OR2X2 OR2X2_3798 ( .A(AES_CORE_DATAPATH__abc_16259_n10584_bF_buf3), .B(\bus_in[16] ), .Y(AES_CORE_DATAPATH__abc_16259_n10633) );
  OR2X2 OR2X2_3799 ( .A(AES_CORE_DATAPATH_iv_0__17_), .B(iv_en_0_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n10635) );
  OR2X2 OR2X2_38 ( .A(AES_CORE_CONTROL_UNIT_state_9_), .B(AES_CORE_CONTROL_UNIT_state_6_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n189_1) );
  OR2X2 OR2X2_380 ( .A(AES_CORE_DATAPATH__abc_16259_n3201_1), .B(AES_CORE_DATAPATH__abc_16259_n3198), .Y(AES_CORE_DATAPATH__abc_16259_n3202) );
  OR2X2 OR2X2_3800 ( .A(AES_CORE_DATAPATH__abc_16259_n10584_bF_buf2), .B(\bus_in[17] ), .Y(AES_CORE_DATAPATH__abc_16259_n10636) );
  OR2X2 OR2X2_3801 ( .A(AES_CORE_DATAPATH_iv_0__18_), .B(iv_en_0_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n10638) );
  OR2X2 OR2X2_3802 ( .A(AES_CORE_DATAPATH__abc_16259_n10584_bF_buf1), .B(\bus_in[18] ), .Y(AES_CORE_DATAPATH__abc_16259_n10639) );
  OR2X2 OR2X2_3803 ( .A(AES_CORE_DATAPATH_iv_0__19_), .B(iv_en_0_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n10641) );
  OR2X2 OR2X2_3804 ( .A(AES_CORE_DATAPATH__abc_16259_n10584_bF_buf0), .B(\bus_in[19] ), .Y(AES_CORE_DATAPATH__abc_16259_n10642) );
  OR2X2 OR2X2_3805 ( .A(AES_CORE_DATAPATH_iv_0__20_), .B(iv_en_0_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n10644) );
  OR2X2 OR2X2_3806 ( .A(AES_CORE_DATAPATH__abc_16259_n10584_bF_buf4), .B(\bus_in[20] ), .Y(AES_CORE_DATAPATH__abc_16259_n10645) );
  OR2X2 OR2X2_3807 ( .A(AES_CORE_DATAPATH_iv_0__21_), .B(iv_en_0_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n10647) );
  OR2X2 OR2X2_3808 ( .A(AES_CORE_DATAPATH__abc_16259_n10584_bF_buf3), .B(\bus_in[21] ), .Y(AES_CORE_DATAPATH__abc_16259_n10648) );
  OR2X2 OR2X2_3809 ( .A(AES_CORE_DATAPATH_iv_0__22_), .B(iv_en_0_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n10650) );
  OR2X2 OR2X2_381 ( .A(AES_CORE_DATAPATH__abc_16259_n3206_1), .B(AES_CORE_DATAPATH__abc_16259_n2826_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n3207_1) );
  OR2X2 OR2X2_3810 ( .A(AES_CORE_DATAPATH__abc_16259_n10584_bF_buf2), .B(\bus_in[22] ), .Y(AES_CORE_DATAPATH__abc_16259_n10651) );
  OR2X2 OR2X2_3811 ( .A(AES_CORE_DATAPATH_iv_0__23_), .B(iv_en_0_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n10653) );
  OR2X2 OR2X2_3812 ( .A(AES_CORE_DATAPATH__abc_16259_n10584_bF_buf1), .B(\bus_in[23] ), .Y(AES_CORE_DATAPATH__abc_16259_n10654) );
  OR2X2 OR2X2_3813 ( .A(AES_CORE_DATAPATH_iv_0__24_), .B(iv_en_0_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n10656) );
  OR2X2 OR2X2_3814 ( .A(AES_CORE_DATAPATH__abc_16259_n10584_bF_buf0), .B(\bus_in[24] ), .Y(AES_CORE_DATAPATH__abc_16259_n10657) );
  OR2X2 OR2X2_3815 ( .A(AES_CORE_DATAPATH_iv_0__25_), .B(iv_en_0_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n10659) );
  OR2X2 OR2X2_3816 ( .A(AES_CORE_DATAPATH__abc_16259_n10584_bF_buf4), .B(\bus_in[25] ), .Y(AES_CORE_DATAPATH__abc_16259_n10660) );
  OR2X2 OR2X2_3817 ( .A(AES_CORE_DATAPATH_iv_0__26_), .B(iv_en_0_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n10662) );
  OR2X2 OR2X2_3818 ( .A(AES_CORE_DATAPATH__abc_16259_n10584_bF_buf3), .B(\bus_in[26] ), .Y(AES_CORE_DATAPATH__abc_16259_n10663) );
  OR2X2 OR2X2_3819 ( .A(AES_CORE_DATAPATH_iv_0__27_), .B(iv_en_0_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n10665) );
  OR2X2 OR2X2_382 ( .A(AES_CORE_DATAPATH__abc_16259_n3208), .B(AES_CORE_DATAPATH__abc_16259_n3209), .Y(AES_CORE_DATAPATH__abc_16259_n3210_1) );
  OR2X2 OR2X2_3820 ( .A(AES_CORE_DATAPATH__abc_16259_n10584_bF_buf2), .B(\bus_in[27] ), .Y(AES_CORE_DATAPATH__abc_16259_n10666) );
  OR2X2 OR2X2_3821 ( .A(AES_CORE_DATAPATH_iv_0__28_), .B(iv_en_0_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n10668) );
  OR2X2 OR2X2_3822 ( .A(AES_CORE_DATAPATH__abc_16259_n10584_bF_buf1), .B(\bus_in[28] ), .Y(AES_CORE_DATAPATH__abc_16259_n10669) );
  OR2X2 OR2X2_3823 ( .A(AES_CORE_DATAPATH_iv_0__29_), .B(iv_en_0_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n10671) );
  OR2X2 OR2X2_3824 ( .A(AES_CORE_DATAPATH__abc_16259_n10584_bF_buf0), .B(\bus_in[29] ), .Y(AES_CORE_DATAPATH__abc_16259_n10672) );
  OR2X2 OR2X2_3825 ( .A(AES_CORE_DATAPATH_iv_0__30_), .B(iv_en_0_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n10674) );
  OR2X2 OR2X2_3826 ( .A(AES_CORE_DATAPATH__abc_16259_n10584_bF_buf4), .B(\bus_in[30] ), .Y(AES_CORE_DATAPATH__abc_16259_n10675) );
  OR2X2 OR2X2_3827 ( .A(AES_CORE_DATAPATH_iv_0__31_), .B(iv_en_0_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n10677) );
  OR2X2 OR2X2_3828 ( .A(AES_CORE_DATAPATH__abc_16259_n10584_bF_buf3), .B(\bus_in[31] ), .Y(AES_CORE_DATAPATH__abc_16259_n10678) );
  OR2X2 OR2X2_3829 ( .A(AES_CORE_CONTROL_UNIT_bypass_key_en), .B(AES_CORE_CONTROL_UNIT_key_en_0_), .Y(AES_CORE_DATAPATH__abc_16259_n10680) );
  OR2X2 OR2X2_383 ( .A(AES_CORE_DATAPATH__abc_16259_n3210_1), .B(AES_CORE_DATAPATH__abc_16259_n3207_1), .Y(AES_CORE_DATAPATH__abc_16259_n3211) );
  OR2X2 OR2X2_3830 ( .A(AES_CORE_DATAPATH__abc_16259_n2806_1), .B(AES_CORE_DATAPATH_key_en_pp1_0_), .Y(AES_CORE_DATAPATH__abc_16259_n10681) );
  OR2X2 OR2X2_3831 ( .A(AES_CORE_CONTROL_UNIT_bypass_key_en), .B(AES_CORE_CONTROL_UNIT_key_en_1_), .Y(AES_CORE_DATAPATH__abc_16259_n10683) );
  OR2X2 OR2X2_3832 ( .A(AES_CORE_DATAPATH__abc_16259_n2806_1), .B(AES_CORE_DATAPATH_key_en_pp1_1_), .Y(AES_CORE_DATAPATH__abc_16259_n10684) );
  OR2X2 OR2X2_3833 ( .A(AES_CORE_CONTROL_UNIT_bypass_key_en), .B(AES_CORE_CONTROL_UNIT_key_en_2_), .Y(AES_CORE_DATAPATH__abc_16259_n10686) );
  OR2X2 OR2X2_3834 ( .A(AES_CORE_DATAPATH__abc_16259_n2806_1), .B(AES_CORE_DATAPATH_key_en_pp1_2_), .Y(AES_CORE_DATAPATH__abc_16259_n10687) );
  OR2X2 OR2X2_3835 ( .A(AES_CORE_CONTROL_UNIT_bypass_key_en), .B(AES_CORE_CONTROL_UNIT_key_en_3_), .Y(AES_CORE_DATAPATH__abc_16259_n10689) );
  OR2X2 OR2X2_3836 ( .A(AES_CORE_DATAPATH__abc_16259_n2806_1), .B(AES_CORE_DATAPATH_key_en_pp1_3_), .Y(AES_CORE_DATAPATH__abc_16259_n10690) );
  OR2X2 OR2X2_3837 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk_bF_buf3), .B(AES_CORE_DATAPATH_col_en_cnt_unit_pp1_0_), .Y(AES_CORE_DATAPATH__abc_16259_n10692) );
  OR2X2 OR2X2_3838 ( .A(AES_CORE_DATAPATH__abc_16259_n2457_1), .B(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_0_), .Y(AES_CORE_DATAPATH__abc_16259_n10693) );
  OR2X2 OR2X2_3839 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk_bF_buf2), .B(AES_CORE_DATAPATH_col_en_cnt_unit_pp1_1_), .Y(AES_CORE_DATAPATH__abc_16259_n10695) );
  OR2X2 OR2X2_384 ( .A(AES_CORE_DATAPATH__abc_16259_n2841_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__9_), .Y(AES_CORE_DATAPATH__abc_16259_n3212_1) );
  OR2X2 OR2X2_3840 ( .A(AES_CORE_DATAPATH__abc_16259_n2457_1), .B(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_1_), .Y(AES_CORE_DATAPATH__abc_16259_n10696) );
  OR2X2 OR2X2_3841 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk_bF_buf1), .B(AES_CORE_DATAPATH_col_en_cnt_unit_pp1_2_), .Y(AES_CORE_DATAPATH__abc_16259_n10698) );
  OR2X2 OR2X2_3842 ( .A(AES_CORE_DATAPATH__abc_16259_n2457_1), .B(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_2_), .Y(AES_CORE_DATAPATH__abc_16259_n10699) );
  OR2X2 OR2X2_3843 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk_bF_buf0), .B(AES_CORE_DATAPATH_col_en_cnt_unit_pp1_3_), .Y(AES_CORE_DATAPATH__abc_16259_n10701) );
  OR2X2 OR2X2_3844 ( .A(AES_CORE_DATAPATH__abc_16259_n2457_1), .B(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_3_), .Y(AES_CORE_DATAPATH__abc_16259_n10702) );
  OR2X2 OR2X2_3845 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk_bF_buf3), .B(AES_CORE_CONTROL_UNIT_col_en_0_), .Y(AES_CORE_DATAPATH__abc_16259_n10704) );
  OR2X2 OR2X2_3846 ( .A(AES_CORE_DATAPATH__abc_16259_n2457_1), .B(AES_CORE_DATAPATH_col_en_cnt_unit_pp1_0_), .Y(AES_CORE_DATAPATH__abc_16259_n10705) );
  OR2X2 OR2X2_3847 ( .A(AES_CORE_CONTROL_UNIT_col_en_1_), .B(AES_CORE_CONTROL_UNIT_bypass_rk_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n10707) );
  OR2X2 OR2X2_3848 ( .A(AES_CORE_DATAPATH__abc_16259_n2457_1), .B(AES_CORE_DATAPATH_col_en_cnt_unit_pp1_1_), .Y(AES_CORE_DATAPATH__abc_16259_n10708) );
  OR2X2 OR2X2_3849 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk_bF_buf1), .B(AES_CORE_CONTROL_UNIT_col_en_2_), .Y(AES_CORE_DATAPATH__abc_16259_n10710) );
  OR2X2 OR2X2_385 ( .A(AES_CORE_DATAPATH__abc_16259_n3204), .B(AES_CORE_DATAPATH__abc_16259_n2853_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n3214_1) );
  OR2X2 OR2X2_3850 ( .A(AES_CORE_DATAPATH__abc_16259_n2457_1), .B(AES_CORE_DATAPATH_col_en_cnt_unit_pp1_2_), .Y(AES_CORE_DATAPATH__abc_16259_n10711) );
  OR2X2 OR2X2_3851 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk_bF_buf0), .B(AES_CORE_CONTROL_UNIT_col_en_3_), .Y(AES_CORE_DATAPATH__abc_16259_n10713) );
  OR2X2 OR2X2_3852 ( .A(AES_CORE_DATAPATH__abc_16259_n2457_1), .B(AES_CORE_DATAPATH_col_en_cnt_unit_pp1_3_), .Y(AES_CORE_DATAPATH__abc_16259_n10714) );
  OR2X2 OR2X2_3853 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf11), .B(AES_CORE_CONTROL_UNIT_key_gen), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec) );
  OR2X2 OR2X2_3854 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n327_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__0_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n328_1) );
  OR2X2 OR2X2_3855 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n329_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__0_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n330_1) );
  OR2X2 OR2X2_3856 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n332_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n333_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n334_1) );
  OR2X2 OR2X2_3857 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n331_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n335_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n336_1) );
  OR2X2 OR2X2_3858 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n338_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__1_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n339_1) );
  OR2X2 OR2X2_3859 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n340_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__1_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n341_1) );
  OR2X2 OR2X2_386 ( .A(AES_CORE_DATAPATH__abc_16259_n3215), .B(AES_CORE_DATAPATH__abc_16259_n3216_1), .Y(AES_CORE_DATAPATH__abc_16259_n3217) );
  OR2X2 OR2X2_3860 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n343_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n344_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n345_1) );
  OR2X2 OR2X2_3861 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n342_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n346_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n347_1) );
  OR2X2 OR2X2_3862 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n349_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__2_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n350_1) );
  OR2X2 OR2X2_3863 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n351_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__2_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n352_1) );
  OR2X2 OR2X2_3864 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n354_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n355_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n356_1) );
  OR2X2 OR2X2_3865 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n353_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n357_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n358_1) );
  OR2X2 OR2X2_3866 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n360_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__3_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n361_1) );
  OR2X2 OR2X2_3867 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n362_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__3_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n363_1) );
  OR2X2 OR2X2_3868 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n365_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n366_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n367_1) );
  OR2X2 OR2X2_3869 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n364_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n368_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n369_1) );
  OR2X2 OR2X2_387 ( .A(_auto_iopadmap_cc_313_execute_26949_9_), .B(AES_CORE_DATAPATH__abc_16259_n3219), .Y(AES_CORE_DATAPATH__abc_16259_n3220) );
  OR2X2 OR2X2_3870 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n371_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__4_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n372_1) );
  OR2X2 OR2X2_3871 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n373_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__4_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n374_1) );
  OR2X2 OR2X2_3872 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n376_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n377_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n378_1) );
  OR2X2 OR2X2_3873 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n375_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n379_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n380_1) );
  OR2X2 OR2X2_3874 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n382_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__5_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n383_1) );
  OR2X2 OR2X2_3875 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n384_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__5_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n385_1) );
  OR2X2 OR2X2_3876 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n387_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n388_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n389_1) );
  OR2X2 OR2X2_3877 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n386_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n390_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n391_1) );
  OR2X2 OR2X2_3878 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n393_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__6_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n394_1) );
  OR2X2 OR2X2_3879 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n395_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__6_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n396_1) );
  OR2X2 OR2X2_388 ( .A(AES_CORE_DATAPATH__abc_16259_n3222), .B(AES_CORE_DATAPATH__abc_16259_n2864_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n3223) );
  OR2X2 OR2X2_3880 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n398_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n399_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n400_1) );
  OR2X2 OR2X2_3881 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n397_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n401_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n402_1) );
  OR2X2 OR2X2_3882 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n404_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__7_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n405_1) );
  OR2X2 OR2X2_3883 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n406_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__7_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n407_1) );
  OR2X2 OR2X2_3884 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n409_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n410_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n411_1) );
  OR2X2 OR2X2_3885 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n408_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n412_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n413_1) );
  OR2X2 OR2X2_3886 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n415_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__8_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n416_1) );
  OR2X2 OR2X2_3887 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n417_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__8_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n418_1) );
  OR2X2 OR2X2_3888 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n420_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n421_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n422_1) );
  OR2X2 OR2X2_3889 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n419_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n423_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n424_1) );
  OR2X2 OR2X2_389 ( .A(AES_CORE_DATAPATH__abc_16259_n3223), .B(AES_CORE_DATAPATH__abc_16259_n3221), .Y(AES_CORE_DATAPATH__abc_16259_n3224) );
  OR2X2 OR2X2_3890 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n426_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__9_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n427_1) );
  OR2X2 OR2X2_3891 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n428_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__9_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n429_1) );
  OR2X2 OR2X2_3892 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n431_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n432_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n433_1) );
  OR2X2 OR2X2_3893 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n430_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n434_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n435_1) );
  OR2X2 OR2X2_3894 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n437_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__10_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n438_1) );
  OR2X2 OR2X2_3895 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n439_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__10_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n440_1) );
  OR2X2 OR2X2_3896 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n442_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n443_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n444_1) );
  OR2X2 OR2X2_3897 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n441_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n445_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n446_1) );
  OR2X2 OR2X2_3898 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n448_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__11_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n449_1) );
  OR2X2 OR2X2_3899 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n450_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__11_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n451_1) );
  OR2X2 OR2X2_39 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n188), .B(AES_CORE_CONTROL_UNIT__abc_15841_n189_1), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n190) );
  OR2X2 OR2X2_390 ( .A(AES_CORE_DATAPATH__abc_16259_n3226), .B(AES_CORE_DATAPATH__abc_16259_n3225), .Y(AES_CORE_DATAPATH__abc_16259_n3227) );
  OR2X2 OR2X2_3900 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n453_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n454_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n455_1) );
  OR2X2 OR2X2_3901 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n452_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n456_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n457_1) );
  OR2X2 OR2X2_3902 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n459_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__12_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n460_1) );
  OR2X2 OR2X2_3903 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n461_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__12_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n462_1) );
  OR2X2 OR2X2_3904 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n464_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n465_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n466_1) );
  OR2X2 OR2X2_3905 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n463_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n467_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n468_1) );
  OR2X2 OR2X2_3906 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n470_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__13_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n471_1) );
  OR2X2 OR2X2_3907 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n472_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__13_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n473_1) );
  OR2X2 OR2X2_3908 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n475_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n476_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n477_1) );
  OR2X2 OR2X2_3909 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n474_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n478_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n479_1) );
  OR2X2 OR2X2_391 ( .A(AES_CORE_DATAPATH__abc_16259_n3227), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n3228_1) );
  OR2X2 OR2X2_3910 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n481_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__14_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n482_1) );
  OR2X2 OR2X2_3911 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n483_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__14_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n484_1) );
  OR2X2 OR2X2_3912 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n486_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n487_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n488_1) );
  OR2X2 OR2X2_3913 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n485_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n489_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n490_1) );
  OR2X2 OR2X2_3914 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n492_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__15_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n493_1) );
  OR2X2 OR2X2_3915 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n494_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__15_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n495_1) );
  OR2X2 OR2X2_3916 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n497_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n498_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n499_1) );
  OR2X2 OR2X2_3917 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n496_1), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n500_1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n501_1) );
  OR2X2 OR2X2_3918 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n503), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__16_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n504) );
  OR2X2 OR2X2_3919 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n505), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__16_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n506) );
  OR2X2 OR2X2_392 ( .A(AES_CORE_DATAPATH__abc_16259_n3230_1), .B(AES_CORE_DATAPATH__abc_16259_n3231), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_9_) );
  OR2X2 OR2X2_3920 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n508), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n509), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n510) );
  OR2X2 OR2X2_3921 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n507), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n511), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n512) );
  OR2X2 OR2X2_3922 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n514), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__17_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n515) );
  OR2X2 OR2X2_3923 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n516), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__17_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n517) );
  OR2X2 OR2X2_3924 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n519), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n520), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n521) );
  OR2X2 OR2X2_3925 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n518), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n522), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n523) );
  OR2X2 OR2X2_3926 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n525), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__18_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n526) );
  OR2X2 OR2X2_3927 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n527), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__18_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n528) );
  OR2X2 OR2X2_3928 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n530), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n531), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n532) );
  OR2X2 OR2X2_3929 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n529), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n533), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n534) );
  OR2X2 OR2X2_393 ( .A(AES_CORE_DATAPATH__abc_16259_n2774_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n3233), .Y(AES_CORE_DATAPATH__abc_16259_n3234) );
  OR2X2 OR2X2_3930 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n536), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__19_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n537) );
  OR2X2 OR2X2_3931 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n538), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__19_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n539) );
  OR2X2 OR2X2_3932 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n541), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n542), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n543) );
  OR2X2 OR2X2_3933 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n540), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n544), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n545) );
  OR2X2 OR2X2_3934 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n547), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__20_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n548) );
  OR2X2 OR2X2_3935 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n549), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__20_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n550) );
  OR2X2 OR2X2_3936 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n552), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n553), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n554) );
  OR2X2 OR2X2_3937 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n551), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n555), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n556) );
  OR2X2 OR2X2_3938 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n558), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__21_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n559) );
  OR2X2 OR2X2_3939 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n560), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__21_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n561) );
  OR2X2 OR2X2_394 ( .A(AES_CORE_DATAPATH__abc_16259_n2778_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n3235_1), .Y(AES_CORE_DATAPATH__abc_16259_n3236_1) );
  OR2X2 OR2X2_3940 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n563), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n564), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n565) );
  OR2X2 OR2X2_3941 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n562), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n566), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n567) );
  OR2X2 OR2X2_3942 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n569), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__22_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n570) );
  OR2X2 OR2X2_3943 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n571), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__22_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n572) );
  OR2X2 OR2X2_3944 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n574), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n575), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n576) );
  OR2X2 OR2X2_3945 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n573), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n577), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n578) );
  OR2X2 OR2X2_3946 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n580), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__23_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n581) );
  OR2X2 OR2X2_3947 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n582), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__23_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n583) );
  OR2X2 OR2X2_3948 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n585), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n586), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n587) );
  OR2X2 OR2X2_3949 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n584), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n588), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n589) );
  OR2X2 OR2X2_395 ( .A(AES_CORE_DATAPATH__abc_16259_n3239_1), .B(AES_CORE_DATAPATH__abc_16259_n3240), .Y(AES_CORE_DATAPATH__abc_16259_n3241_1) );
  OR2X2 OR2X2_3950 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__24_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__24_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n591) );
  OR2X2 OR2X2_3951 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_round_2_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_round_1_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n604) );
  OR2X2 OR2X2_3952 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n604), .B(AES_CORE_DATAPATH_KEY_EXPANDER_round_0_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n605) );
  OR2X2 OR2X2_3953 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n603), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n606), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n607) );
  OR2X2 OR2X2_3954 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n607), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_24_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n610) );
  OR2X2 OR2X2_3955 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n611), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n596), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n612) );
  OR2X2 OR2X2_3956 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n614), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n615), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_88_) );
  OR2X2 OR2X2_3957 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__25_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__25_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n617) );
  OR2X2 OR2X2_3958 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n623), .B(AES_CORE_DATAPATH_KEY_EXPANDER_round_1_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n624) );
  OR2X2 OR2X2_3959 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_round_3_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_round_2_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n625) );
  OR2X2 OR2X2_396 ( .A(AES_CORE_DATAPATH__abc_16259_n3241_1), .B(AES_CORE_DATAPATH__abc_16259_n3238), .Y(AES_CORE_DATAPATH__abc_16259_n3242) );
  OR2X2 OR2X2_3960 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n624), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n625), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n626) );
  OR2X2 OR2X2_3961 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n631), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597_bF_buf2), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n632) );
  OR2X2 OR2X2_3962 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n634), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n628), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n635) );
  OR2X2 OR2X2_3963 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n635), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n622), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n636) );
  OR2X2 OR2X2_3964 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n645), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n637), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n646) );
  OR2X2 OR2X2_3965 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n646), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n596), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n647) );
  OR2X2 OR2X2_3966 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n648), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n641), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_89_) );
  OR2X2 OR2X2_3967 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__26_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__26_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n650) );
  OR2X2 OR2X2_3968 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n604), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n656), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n657) );
  OR2X2 OR2X2_3969 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n657), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n623), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n658) );
  OR2X2 OR2X2_397 ( .A(AES_CORE_DATAPATH__abc_16259_n3246), .B(AES_CORE_DATAPATH__abc_16259_n2826_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n3247) );
  OR2X2 OR2X2_3970 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n663), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n632), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n664) );
  OR2X2 OR2X2_3971 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n665), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n668), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n669) );
  OR2X2 OR2X2_3972 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n672), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n655), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n675) );
  OR2X2 OR2X2_3973 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n681), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n661), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n682) );
  OR2X2 OR2X2_3974 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n683), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n670), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n684) );
  OR2X2 OR2X2_3975 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n685), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n673), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n686) );
  OR2X2 OR2X2_3976 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n686), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n596), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n687) );
  OR2X2 OR2X2_3977 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n688), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n678), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_90_) );
  OR2X2 OR2X2_3978 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__27_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__27_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n690) );
  OR2X2 OR2X2_3979 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n695), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf5), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n696) );
  OR2X2 OR2X2_398 ( .A(AES_CORE_DATAPATH__abc_16259_n3248), .B(AES_CORE_DATAPATH__abc_16259_n3249), .Y(AES_CORE_DATAPATH__abc_16259_n3250) );
  OR2X2 OR2X2_3980 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n696), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n697), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n698) );
  OR2X2 OR2X2_3981 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n632), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n699), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n700) );
  OR2X2 OR2X2_3982 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n701), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_27_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n704) );
  OR2X2 OR2X2_3983 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n709), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n707), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_91_) );
  OR2X2 OR2X2_3984 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__28_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__28_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n711) );
  OR2X2 OR2X2_3985 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n717), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf4), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n718) );
  OR2X2 OR2X2_3986 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n718), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n719), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n720) );
  OR2X2 OR2X2_3987 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n721), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n725), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n726) );
  OR2X2 OR2X2_3988 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n726), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n716), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n727) );
  OR2X2 OR2X2_3989 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n729), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_28_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n730) );
  OR2X2 OR2X2_399 ( .A(AES_CORE_DATAPATH__abc_16259_n3250), .B(AES_CORE_DATAPATH__abc_16259_n3247), .Y(AES_CORE_DATAPATH__abc_16259_n3251) );
  OR2X2 OR2X2_3990 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n734), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n735), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n736) );
  OR2X2 OR2X2_3991 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n736), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n596), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n737) );
  OR2X2 OR2X2_3992 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n738), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n733), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_92_) );
  OR2X2 OR2X2_3993 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__29_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__29_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n740) );
  OR2X2 OR2X2_3994 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n747), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n632), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n748) );
  OR2X2 OR2X2_3995 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n749), .B(AES_CORE_DATAPATH_KEY_EXPANDER_round_3_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n750) );
  OR2X2 OR2X2_3996 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n696), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n750), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n751) );
  OR2X2 OR2X2_3997 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n752), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n745), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n755) );
  OR2X2 OR2X2_3998 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n681), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n719), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n759) );
  OR2X2 OR2X2_3999 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n760), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n761), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n762) );
  OR2X2 OR2X2_4 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n78), .B(AES_CORE_CONTROL_UNIT_state_13_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n79_1) );
  OR2X2 OR2X2_40 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n193), .B(AES_CORE_CONTROL_UNIT__abc_15841_n140), .Y(AES_CORE_CONTROL_UNIT_col_en_0_) );
  OR2X2 OR2X2_400 ( .A(AES_CORE_DATAPATH__abc_16259_n2841_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__10_), .Y(AES_CORE_DATAPATH__abc_16259_n3252) );
  OR2X2 OR2X2_4000 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n763), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n753), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n764) );
  OR2X2 OR2X2_4001 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n764), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n596), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n765) );
  OR2X2 OR2X2_4002 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n766), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n758), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_93_) );
  OR2X2 OR2X2_4003 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__30_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__30_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n768) );
  OR2X2 OR2X2_4004 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n779), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n696), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n780) );
  OR2X2 OR2X2_4005 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n780), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n774), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n781) );
  OR2X2 OR2X2_4006 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n785), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n773), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n786) );
  OR2X2 OR2X2_4007 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n788), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n783), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n789) );
  OR2X2 OR2X2_4008 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n789), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_30_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n790) );
  OR2X2 OR2X2_4009 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n795), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n794), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n796) );
  OR2X2 OR2X2_401 ( .A(AES_CORE_DATAPATH__abc_16259_n3244), .B(AES_CORE_DATAPATH__abc_16259_n2853_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n3254) );
  OR2X2 OR2X2_4010 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n796), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n596), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n797) );
  OR2X2 OR2X2_4011 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n798), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n793), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_94_) );
  OR2X2 OR2X2_4012 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__31_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__31_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n800) );
  OR2X2 OR2X2_4013 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n780), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n806), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n807) );
  OR2X2 OR2X2_4014 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n810), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n805), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n811) );
  OR2X2 OR2X2_4015 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n812), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n808), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n813) );
  OR2X2 OR2X2_4016 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n813), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_31_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n814) );
  OR2X2 OR2X2_4017 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n819), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n818), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n820) );
  OR2X2 OR2X2_4018 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n820), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n596), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n821) );
  OR2X2 OR2X2_4019 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n822), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n817), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_95_) );
  OR2X2 OR2X2_402 ( .A(AES_CORE_DATAPATH__abc_16259_n3255), .B(AES_CORE_DATAPATH__abc_16259_n3256), .Y(AES_CORE_DATAPATH__abc_16259_n3257_1) );
  OR2X2 OR2X2_4020 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__0_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__0_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n824) );
  OR2X2 OR2X2_4021 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_0_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf2), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n828) );
  OR2X2 OR2X2_4022 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__0_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n829) );
  OR2X2 OR2X2_4023 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__1_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__1_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n831) );
  OR2X2 OR2X2_4024 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_1_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n835) );
  OR2X2 OR2X2_4025 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__1_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n836) );
  OR2X2 OR2X2_4026 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__2_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__2_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n838) );
  OR2X2 OR2X2_4027 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_2_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf0), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n842) );
  OR2X2 OR2X2_4028 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__2_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n843) );
  OR2X2 OR2X2_4029 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__3_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__3_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n845) );
  OR2X2 OR2X2_403 ( .A(_auto_iopadmap_cc_313_execute_26949_10_), .B(AES_CORE_DATAPATH__abc_16259_n3259_1), .Y(AES_CORE_DATAPATH__abc_16259_n3260) );
  OR2X2 OR2X2_4030 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_3_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf7), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n849) );
  OR2X2 OR2X2_4031 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__3_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n850) );
  OR2X2 OR2X2_4032 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__4_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__4_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n852) );
  OR2X2 OR2X2_4033 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_4_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf6), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n856) );
  OR2X2 OR2X2_4034 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__4_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n857) );
  OR2X2 OR2X2_4035 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__5_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__5_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n859) );
  OR2X2 OR2X2_4036 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_5_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf5), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n863) );
  OR2X2 OR2X2_4037 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__5_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n864) );
  OR2X2 OR2X2_4038 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__6_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__6_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n866) );
  OR2X2 OR2X2_4039 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_6_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf4), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n870) );
  OR2X2 OR2X2_404 ( .A(AES_CORE_DATAPATH__abc_16259_n3262), .B(AES_CORE_DATAPATH__abc_16259_n2864_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n3263) );
  OR2X2 OR2X2_4040 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__6_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n871) );
  OR2X2 OR2X2_4041 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__7_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__7_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n873) );
  OR2X2 OR2X2_4042 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_7_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf3), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n877) );
  OR2X2 OR2X2_4043 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__7_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n878) );
  OR2X2 OR2X2_4044 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__8_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__8_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n880) );
  OR2X2 OR2X2_4045 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_8_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf2), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n884) );
  OR2X2 OR2X2_4046 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__8_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n885) );
  OR2X2 OR2X2_4047 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__9_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__9_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n887) );
  OR2X2 OR2X2_4048 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_9_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n891) );
  OR2X2 OR2X2_4049 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__9_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n892) );
  OR2X2 OR2X2_405 ( .A(AES_CORE_DATAPATH__abc_16259_n3263), .B(AES_CORE_DATAPATH__abc_16259_n3261), .Y(AES_CORE_DATAPATH__abc_16259_n3264_1) );
  OR2X2 OR2X2_4050 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__10_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__10_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n894) );
  OR2X2 OR2X2_4051 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_10_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf0), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n898) );
  OR2X2 OR2X2_4052 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__10_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n899) );
  OR2X2 OR2X2_4053 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__11_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__11_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n901) );
  OR2X2 OR2X2_4054 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_11_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf7), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n905) );
  OR2X2 OR2X2_4055 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__11_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n906) );
  OR2X2 OR2X2_4056 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__12_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__12_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n908) );
  OR2X2 OR2X2_4057 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_12_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf6), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n912) );
  OR2X2 OR2X2_4058 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__12_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n913) );
  OR2X2 OR2X2_4059 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__13_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__13_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n915) );
  OR2X2 OR2X2_406 ( .A(AES_CORE_DATAPATH__abc_16259_n3266), .B(AES_CORE_DATAPATH__abc_16259_n3265_1), .Y(AES_CORE_DATAPATH__abc_16259_n3267) );
  OR2X2 OR2X2_4060 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_13_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf5), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n919) );
  OR2X2 OR2X2_4061 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__13_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n920) );
  OR2X2 OR2X2_4062 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__14_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__14_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n922) );
  OR2X2 OR2X2_4063 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_14_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf4), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n926) );
  OR2X2 OR2X2_4064 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__14_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n927) );
  OR2X2 OR2X2_4065 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__15_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__15_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n929) );
  OR2X2 OR2X2_4066 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_15_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf3), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n933) );
  OR2X2 OR2X2_4067 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__15_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n934) );
  OR2X2 OR2X2_4068 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__16_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__16_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n936) );
  OR2X2 OR2X2_4069 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_16_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf2), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n940) );
  OR2X2 OR2X2_407 ( .A(AES_CORE_DATAPATH__abc_16259_n3267), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n3268_1) );
  OR2X2 OR2X2_4070 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__16_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n941) );
  OR2X2 OR2X2_4071 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__17_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__17_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n943) );
  OR2X2 OR2X2_4072 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_17_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n947) );
  OR2X2 OR2X2_4073 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__17_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n948) );
  OR2X2 OR2X2_4074 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__18_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__18_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n950) );
  OR2X2 OR2X2_4075 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_18_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf0), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n954) );
  OR2X2 OR2X2_4076 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__18_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n955) );
  OR2X2 OR2X2_4077 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__19_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__19_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n957) );
  OR2X2 OR2X2_4078 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_19_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf7), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n961) );
  OR2X2 OR2X2_4079 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__19_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n962) );
  OR2X2 OR2X2_408 ( .A(AES_CORE_DATAPATH__abc_16259_n3270_1), .B(AES_CORE_DATAPATH__abc_16259_n3271), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_10_) );
  OR2X2 OR2X2_4080 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__20_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__20_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n964) );
  OR2X2 OR2X2_4081 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_20_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf6), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n968) );
  OR2X2 OR2X2_4082 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__20_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n969) );
  OR2X2 OR2X2_4083 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__21_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__21_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n971) );
  OR2X2 OR2X2_4084 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_21_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf5), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n975) );
  OR2X2 OR2X2_4085 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__21_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n976) );
  OR2X2 OR2X2_4086 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__22_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__22_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n978) );
  OR2X2 OR2X2_4087 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_22_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf4), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n982) );
  OR2X2 OR2X2_4088 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__22_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n983) );
  OR2X2 OR2X2_4089 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__23_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__23_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n985) );
  OR2X2 OR2X2_409 ( .A(AES_CORE_DATAPATH__abc_16259_n2774_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n3273), .Y(AES_CORE_DATAPATH__abc_16259_n3274_1) );
  OR2X2 OR2X2_4090 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_23_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf3), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n989) );
  OR2X2 OR2X2_4091 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__23_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n990) );
  OR2X2 OR2X2_4092 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__24_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__24_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n992) );
  OR2X2 OR2X2_4093 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_24_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf2), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n996) );
  OR2X2 OR2X2_4094 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__24_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n997) );
  OR2X2 OR2X2_4095 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__25_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__25_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n999) );
  OR2X2 OR2X2_4096 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_25_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf1), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1003) );
  OR2X2 OR2X2_4097 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__25_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1004) );
  OR2X2 OR2X2_4098 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__26_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__26_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1006) );
  OR2X2 OR2X2_4099 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_26_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf0), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1010) );
  OR2X2 OR2X2_41 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt_bF_buf9), .B(AES_CORE_CONTROL_UNIT_last_round_bF_buf1), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n195) );
  OR2X2 OR2X2_410 ( .A(AES_CORE_DATAPATH__abc_16259_n2778_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n3275), .Y(AES_CORE_DATAPATH__abc_16259_n3276) );
  OR2X2 OR2X2_4100 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__26_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1011) );
  OR2X2 OR2X2_4101 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__27_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__27_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1013) );
  OR2X2 OR2X2_4102 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_27_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf7), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1017) );
  OR2X2 OR2X2_4103 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__27_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1018) );
  OR2X2 OR2X2_4104 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__28_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__28_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1020) );
  OR2X2 OR2X2_4105 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_28_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf6), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1024) );
  OR2X2 OR2X2_4106 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__28_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1025) );
  OR2X2 OR2X2_4107 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__29_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__29_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1027) );
  OR2X2 OR2X2_4108 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_29_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf5), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1031) );
  OR2X2 OR2X2_4109 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__29_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1032) );
  OR2X2 OR2X2_411 ( .A(AES_CORE_DATAPATH__abc_16259_n3279), .B(AES_CORE_DATAPATH__abc_16259_n3280), .Y(AES_CORE_DATAPATH__abc_16259_n3281) );
  OR2X2 OR2X2_4110 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__30_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__30_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1034) );
  OR2X2 OR2X2_4111 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_30_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf4), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1038) );
  OR2X2 OR2X2_4112 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__30_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1039) );
  OR2X2 OR2X2_4113 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__31_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__31_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1041) );
  OR2X2 OR2X2_4114 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_31_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf3), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1045) );
  OR2X2 OR2X2_4115 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n597_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__31_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1046) );
  OR2X2 OR2X2_4116 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__0_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_0_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1048) );
  OR2X2 OR2X2_4117 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__1_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_1_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1052) );
  OR2X2 OR2X2_4118 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__2_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_2_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1056) );
  OR2X2 OR2X2_4119 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__3_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_3_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1060) );
  OR2X2 OR2X2_412 ( .A(AES_CORE_DATAPATH__abc_16259_n3281), .B(AES_CORE_DATAPATH__abc_16259_n3278), .Y(AES_CORE_DATAPATH__abc_16259_n3282) );
  OR2X2 OR2X2_4120 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__4_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_4_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1064) );
  OR2X2 OR2X2_4121 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__5_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_5_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1068) );
  OR2X2 OR2X2_4122 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__6_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_6_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1072) );
  OR2X2 OR2X2_4123 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__7_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_7_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1076) );
  OR2X2 OR2X2_4124 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__8_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_8_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1080) );
  OR2X2 OR2X2_4125 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__9_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_9_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1084) );
  OR2X2 OR2X2_4126 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__10_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_10_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1088) );
  OR2X2 OR2X2_4127 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__11_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_11_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1092) );
  OR2X2 OR2X2_4128 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__12_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_12_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1096) );
  OR2X2 OR2X2_4129 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__13_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_13_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1100) );
  OR2X2 OR2X2_413 ( .A(AES_CORE_DATAPATH__abc_16259_n3286_1), .B(AES_CORE_DATAPATH__abc_16259_n2826_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n3287) );
  OR2X2 OR2X2_4130 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__14_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_14_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1104) );
  OR2X2 OR2X2_4131 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__15_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_15_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1108) );
  OR2X2 OR2X2_4132 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__16_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_16_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1112) );
  OR2X2 OR2X2_4133 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__17_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_17_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1116) );
  OR2X2 OR2X2_4134 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__18_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_18_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1120) );
  OR2X2 OR2X2_4135 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__19_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_19_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1124) );
  OR2X2 OR2X2_4136 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__20_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_20_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1128) );
  OR2X2 OR2X2_4137 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__21_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_21_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1132) );
  OR2X2 OR2X2_4138 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__22_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_22_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1136) );
  OR2X2 OR2X2_4139 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__23_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_23_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1140) );
  OR2X2 OR2X2_414 ( .A(AES_CORE_DATAPATH__abc_16259_n3288_1), .B(AES_CORE_DATAPATH__abc_16259_n3289), .Y(AES_CORE_DATAPATH__abc_16259_n3290) );
  OR2X2 OR2X2_4140 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1146), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1147), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_120_) );
  OR2X2 OR2X2_4141 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n646), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1149), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1150) );
  OR2X2 OR2X2_4142 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n639), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__25_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1151) );
  OR2X2 OR2X2_4143 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1153), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1155), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_122_) );
  OR2X2 OR2X2_4144 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1158), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1157), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1159) );
  OR2X2 OR2X2_4145 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n705), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__27_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1160) );
  OR2X2 OR2X2_4146 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n736), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1162), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1163) );
  OR2X2 OR2X2_4147 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n731), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__28_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1164) );
  OR2X2 OR2X2_4148 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1166), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1168), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_125_) );
  OR2X2 OR2X2_4149 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n791), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__30_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1170) );
  OR2X2 OR2X2_415 ( .A(AES_CORE_DATAPATH__abc_16259_n3290), .B(AES_CORE_DATAPATH__abc_16259_n3287), .Y(AES_CORE_DATAPATH__abc_16259_n3291) );
  OR2X2 OR2X2_4150 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n796), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1171), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1172) );
  OR2X2 OR2X2_4151 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n815), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__31_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1174) );
  OR2X2 OR2X2_4152 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n820), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1175), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1176) );
  OR2X2 OR2X2_4153 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__0_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__0_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1178) );
  OR2X2 OR2X2_4154 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__1_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__1_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1182) );
  OR2X2 OR2X2_4155 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__2_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__2_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1186) );
  OR2X2 OR2X2_4156 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__3_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__3_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1190) );
  OR2X2 OR2X2_4157 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__4_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__4_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1194) );
  OR2X2 OR2X2_4158 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__5_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__5_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1198) );
  OR2X2 OR2X2_4159 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__6_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__6_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1202) );
  OR2X2 OR2X2_416 ( .A(AES_CORE_DATAPATH__abc_16259_n2841_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__11_), .Y(AES_CORE_DATAPATH__abc_16259_n3292) );
  OR2X2 OR2X2_4160 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__7_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__7_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1206) );
  OR2X2 OR2X2_4161 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__8_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__8_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1210) );
  OR2X2 OR2X2_4162 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__9_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__9_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1214) );
  OR2X2 OR2X2_4163 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__10_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__10_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1218) );
  OR2X2 OR2X2_4164 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__11_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__11_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1222) );
  OR2X2 OR2X2_4165 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__12_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__12_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1226) );
  OR2X2 OR2X2_4166 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__13_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__13_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1230) );
  OR2X2 OR2X2_4167 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__14_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__14_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1234) );
  OR2X2 OR2X2_4168 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__15_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__15_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1238) );
  OR2X2 OR2X2_4169 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__16_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__16_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1242) );
  OR2X2 OR2X2_417 ( .A(AES_CORE_DATAPATH__abc_16259_n3284), .B(AES_CORE_DATAPATH__abc_16259_n2853_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n3294_1) );
  OR2X2 OR2X2_4170 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__17_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__17_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1246) );
  OR2X2 OR2X2_4171 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__18_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__18_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1250) );
  OR2X2 OR2X2_4172 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__19_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__19_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1254) );
  OR2X2 OR2X2_4173 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__20_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__20_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1258) );
  OR2X2 OR2X2_4174 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__21_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__21_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1262) );
  OR2X2 OR2X2_4175 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__22_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__22_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1266) );
  OR2X2 OR2X2_4176 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__23_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__23_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1270) );
  OR2X2 OR2X2_4177 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__24_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__24_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1274) );
  OR2X2 OR2X2_4178 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__25_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__25_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1278) );
  OR2X2 OR2X2_4179 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__26_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__26_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1282) );
  OR2X2 OR2X2_418 ( .A(AES_CORE_DATAPATH__abc_16259_n3295), .B(AES_CORE_DATAPATH__abc_16259_n3296), .Y(AES_CORE_DATAPATH__abc_16259_n3297_1) );
  OR2X2 OR2X2_4180 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__27_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__27_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1286) );
  OR2X2 OR2X2_4181 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__28_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__28_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1290) );
  OR2X2 OR2X2_4182 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__29_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__29_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1294) );
  OR2X2 OR2X2_4183 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__30_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__30_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1298) );
  OR2X2 OR2X2_4184 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__31_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__31_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24521_n1302) );
  OR2X2 OR2X2_4185 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n99), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n100), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n101) );
  OR2X2 OR2X2_4186 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n102), .B(AES_CORE_DATAPATH_MIX_COL_col_0__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n103) );
  OR2X2 OR2X2_4187 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n104), .B(AES_CORE_DATAPATH_MIX_COL_col_3__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n105_1) );
  OR2X2 OR2X2_4188 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n108), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n110), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n111) );
  OR2X2 OR2X2_4189 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n111), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n101), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n112) );
  OR2X2 OR2X2_419 ( .A(_auto_iopadmap_cc_313_execute_26949_11_), .B(AES_CORE_DATAPATH__abc_16259_n3299_1), .Y(AES_CORE_DATAPATH__abc_16259_n3300) );
  OR2X2 OR2X2_4190 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__0_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n113) );
  OR2X2 OR2X2_4191 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n116), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n115_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n117) );
  OR2X2 OR2X2_4192 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n122), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n123_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n124) );
  OR2X2 OR2X2_4193 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__5_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n125) );
  OR2X2 OR2X2_4194 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__5_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n129_1) );
  OR2X2 OR2X2_4195 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n128), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n132), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n133) );
  OR2X2 OR2X2_4196 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n136_1), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n126), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n137) );
  OR2X2 OR2X2_4197 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n140_1), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n130), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n141) );
  OR2X2 OR2X2_4198 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n137), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n141), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n142_1) );
  OR2X2 OR2X2_4199 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n143), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n124), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n144) );
  OR2X2 OR2X2_42 ( .A(AES_CORE_CONTROL_UNIT_state_14_), .B(AES_CORE_CONTROL_UNIT_state_4_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n198) );
  OR2X2 OR2X2_420 ( .A(AES_CORE_DATAPATH__abc_16259_n3302), .B(AES_CORE_DATAPATH__abc_16259_n2864_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n3303_1) );
  OR2X2 OR2X2_4200 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__6_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n145) );
  OR2X2 OR2X2_4201 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n148), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n149_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n150) );
  OR2X2 OR2X2_4202 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n150), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n147_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n151) );
  OR2X2 OR2X2_4203 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n119_1), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n152), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n153) );
  OR2X2 OR2X2_4204 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n143), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n147_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n154_1) );
  OR2X2 OR2X2_4205 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n150), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n124), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n155) );
  OR2X2 OR2X2_4206 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_0_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n156_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n157) );
  OR2X2 OR2X2_4207 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n98), .B(AES_CORE_DATAPATH_MIX_COL_col_0__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n159) );
  OR2X2 OR2X2_4208 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n160_1), .B(AES_CORE_DATAPATH_MIX_COL_col_3__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n161) );
  OR2X2 OR2X2_4209 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n107), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n162_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n165) );
  OR2X2 OR2X2_421 ( .A(AES_CORE_DATAPATH__abc_16259_n3303_1), .B(AES_CORE_DATAPATH__abc_16259_n3301_1), .Y(AES_CORE_DATAPATH__abc_16259_n3304) );
  OR2X2 OR2X2_4210 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__1_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n168_1) );
  OR2X2 OR2X2_4211 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n176_1), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n169), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n177_1) );
  OR2X2 OR2X2_4212 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n178), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n172_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n179) );
  OR2X2 OR2X2_4213 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n181_1), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n182), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n183_1) );
  OR2X2 OR2X2_4214 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__7_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n185) );
  OR2X2 OR2X2_4215 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n191_1), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n186), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n192_1) );
  OR2X2 OR2X2_4216 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n189), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n193), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n194_1) );
  OR2X2 OR2X2_4217 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n197_1), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n198_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n199) );
  OR2X2 OR2X2_4218 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n152), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n199), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n200_1) );
  OR2X2 OR2X2_4219 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__6_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n201_1) );
  OR2X2 OR2X2_422 ( .A(AES_CORE_DATAPATH__abc_16259_n3306), .B(AES_CORE_DATAPATH__abc_16259_n3305), .Y(AES_CORE_DATAPATH__abc_16259_n3307) );
  OR2X2 OR2X2_4220 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n156_1), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n203_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n204_1) );
  OR2X2 OR2X2_4221 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n205), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n194_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n206) );
  OR2X2 OR2X2_4222 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n192_1), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n147_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n207_1) );
  OR2X2 OR2X2_4223 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n124), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n188_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n208_1) );
  OR2X2 OR2X2_4224 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n210_1), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n211_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n212) );
  OR2X2 OR2X2_4225 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n212), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n209), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n213) );
  OR2X2 OR2X2_4226 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n214_1), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n215_1) );
  OR2X2 OR2X2_4227 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n212), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n194_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n216) );
  OR2X2 OR2X2_4228 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n205), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n209), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n217) );
  OR2X2 OR2X2_4229 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n218_1), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n183_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n219_1) );
  OR2X2 OR2X2_423 ( .A(AES_CORE_DATAPATH__abc_16259_n3307), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n3308) );
  OR2X2 OR2X2_4230 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n175), .B(AES_CORE_DATAPATH_MIX_COL_col_0__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n221_1) );
  OR2X2 OR2X2_4231 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n222_1), .B(AES_CORE_DATAPATH_MIX_COL_col_3__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n223) );
  OR2X2 OR2X2_4232 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n224_1), .B(AES_CORE_DATAPATH_MIX_COL_col_2__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n227_1) );
  OR2X2 OR2X2_4233 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n231), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n233), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n234) );
  OR2X2 OR2X2_4234 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n236), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n237), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_2_) );
  OR2X2 OR2X2_4235 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__0_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n239) );
  OR2X2 OR2X2_4236 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n192_1), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n242), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n243) );
  OR2X2 OR2X2_4237 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n244), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n240), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n245) );
  OR2X2 OR2X2_4238 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n245), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n188_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n246) );
  OR2X2 OR2X2_4239 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n249), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n250), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n251) );
  OR2X2 OR2X2_424 ( .A(AES_CORE_DATAPATH__abc_16259_n3310), .B(AES_CORE_DATAPATH__abc_16259_n3311), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_11_) );
  OR2X2 OR2X2_4240 ( .A(AES_CORE_DATAPATH_MIX_COL_col_3__7_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n253) );
  OR2X2 OR2X2_4241 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n252), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n256), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n257) );
  OR2X2 OR2X2_4242 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n199), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n255), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n259) );
  OR2X2 OR2X2_4243 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n251), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n203_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n260) );
  OR2X2 OR2X2_4244 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n258), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n262), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n263) );
  OR2X2 OR2X2_4245 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n264), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n247), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n265) );
  OR2X2 OR2X2_4246 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n266), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n267), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n268) );
  OR2X2 OR2X2_4247 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n263), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n268), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n269) );
  OR2X2 OR2X2_4248 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n271), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n272) );
  OR2X2 OR2X2_4249 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n270), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n273), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n274) );
  OR2X2 OR2X2_425 ( .A(AES_CORE_DATAPATH__abc_16259_n2774_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n3313), .Y(AES_CORE_DATAPATH__abc_16259_n3314) );
  OR2X2 OR2X2_4250 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n230), .B(AES_CORE_DATAPATH_MIX_COL_col_0__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n276) );
  OR2X2 OR2X2_4251 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n277), .B(AES_CORE_DATAPATH_MIX_COL_col_3__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n278) );
  OR2X2 OR2X2_4252 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n107), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n279), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n282) );
  OR2X2 OR2X2_4253 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n286), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n288), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n289) );
  OR2X2 OR2X2_4254 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n293), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n290), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n294) );
  OR2X2 OR2X2_4255 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n296), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n297), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n298) );
  OR2X2 OR2X2_4256 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n101), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n255), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n300) );
  OR2X2 OR2X2_4257 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n251), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n115_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n301) );
  OR2X2 OR2X2_4258 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n247), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n302), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n303) );
  OR2X2 OR2X2_4259 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n304), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n305), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n306) );
  OR2X2 OR2X2_426 ( .A(AES_CORE_DATAPATH__abc_16259_n2778_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n3315_1), .Y(AES_CORE_DATAPATH__abc_16259_n3316) );
  OR2X2 OR2X2_4260 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n268), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n306), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n307) );
  OR2X2 OR2X2_4261 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n308), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n143), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n309) );
  OR2X2 OR2X2_4262 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n310), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n311), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n312) );
  OR2X2 OR2X2_4263 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n312), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n150), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n313) );
  OR2X2 OR2X2_4264 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__1_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n315) );
  OR2X2 OR2X2_4265 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n147_1), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n318), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n319) );
  OR2X2 OR2X2_4266 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n320), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n316), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n321) );
  OR2X2 OR2X2_4267 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n124), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n321), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n322) );
  OR2X2 OR2X2_4268 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n314), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n323), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n324) );
  OR2X2 OR2X2_4269 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n312), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n143), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n325) );
  OR2X2 OR2X2_427 ( .A(AES_CORE_DATAPATH__abc_16259_n3319), .B(AES_CORE_DATAPATH__abc_16259_n3320), .Y(AES_CORE_DATAPATH__abc_16259_n3321) );
  OR2X2 OR2X2_4270 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n308), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n150), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n326) );
  OR2X2 OR2X2_4271 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n328), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n329), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n330) );
  OR2X2 OR2X2_4272 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n327), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n330), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n331) );
  OR2X2 OR2X2_4273 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n332), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n333) );
  OR2X2 OR2X2_4274 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n314), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n330), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n334) );
  OR2X2 OR2X2_4275 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n327), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n323), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n335) );
  OR2X2 OR2X2_4276 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n336), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n298), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n337) );
  OR2X2 OR2X2_4277 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n285), .B(AES_CORE_DATAPATH_MIX_COL_col_0__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n339) );
  OR2X2 OR2X2_4278 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n340), .B(AES_CORE_DATAPATH_MIX_COL_col_3__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n341) );
  OR2X2 OR2X2_4279 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n107), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n342), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n345) );
  OR2X2 OR2X2_428 ( .A(AES_CORE_DATAPATH__abc_16259_n3321), .B(AES_CORE_DATAPATH__abc_16259_n3318), .Y(AES_CORE_DATAPATH__abc_16259_n3322_1) );
  OR2X2 OR2X2_4280 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n348), .B(AES_CORE_DATAPATH_MIX_COL_col_3__4_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n349) );
  OR2X2 OR2X2_4281 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n350), .B(AES_CORE_DATAPATH_MIX_COL_col_1__4_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n351) );
  OR2X2 OR2X2_4282 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n354), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n356), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n357) );
  OR2X2 OR2X2_4283 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n359), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n360), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n361) );
  OR2X2 OR2X2_4284 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n363), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n365), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n366) );
  OR2X2 OR2X2_4285 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n209), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n366), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n367) );
  OR2X2 OR2X2_4286 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n194_1), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n368), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n369) );
  OR2X2 OR2X2_4287 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n372), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n371), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n373) );
  OR2X2 OR2X2_4288 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n177_1), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n199), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n375) );
  OR2X2 OR2X2_4289 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n171), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n203_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n376) );
  OR2X2 OR2X2_429 ( .A(AES_CORE_DATAPATH__abc_16259_n3326_1), .B(AES_CORE_DATAPATH__abc_16259_n2826_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n3327) );
  OR2X2 OR2X2_4290 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n378), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n374), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n379) );
  OR2X2 OR2X2_4291 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n379), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n150), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n380) );
  OR2X2 OR2X2_4292 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n323), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n377), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n381) );
  OR2X2 OR2X2_4293 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n330), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n373), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n382) );
  OR2X2 OR2X2_4294 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n383), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n143), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n384) );
  OR2X2 OR2X2_4295 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n385), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n370), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n386) );
  OR2X2 OR2X2_4296 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n209), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n368), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n387) );
  OR2X2 OR2X2_4297 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n194_1), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n366), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n388) );
  OR2X2 OR2X2_4298 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n383), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n150), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n390) );
  OR2X2 OR2X2_4299 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n379), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n143), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n391) );
  OR2X2 OR2X2_43 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n193), .B(AES_CORE_CONTROL_UNIT__abc_15841_n199), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n200_1) );
  OR2X2 OR2X2_430 ( .A(AES_CORE_DATAPATH__abc_16259_n3328_1), .B(AES_CORE_DATAPATH__abc_16259_n3329), .Y(AES_CORE_DATAPATH__abc_16259_n3330_1) );
  OR2X2 OR2X2_4300 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n392), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n389), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n393) );
  OR2X2 OR2X2_4301 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n394), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n361), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n395) );
  OR2X2 OR2X2_4302 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n392), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n370), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n396) );
  OR2X2 OR2X2_4303 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n385), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n389), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n397) );
  OR2X2 OR2X2_4304 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n398), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_4_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n399) );
  OR2X2 OR2X2_4305 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n402), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n401), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n403) );
  OR2X2 OR2X2_4306 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n406), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n407), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n408) );
  OR2X2 OR2X2_4307 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n410), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n411), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n412) );
  OR2X2 OR2X2_4308 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__3_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n414) );
  OR2X2 OR2X2_4309 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n419), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n420), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n421) );
  OR2X2 OR2X2_431 ( .A(AES_CORE_DATAPATH__abc_16259_n3330_1), .B(AES_CORE_DATAPATH__abc_16259_n3327), .Y(AES_CORE_DATAPATH__abc_16259_n3331) );
  OR2X2 OR2X2_4310 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n261), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n235), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n422) );
  OR2X2 OR2X2_4311 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n257), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n234), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n423) );
  OR2X2 OR2X2_4312 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n389), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n424), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n425) );
  OR2X2 OR2X2_4313 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n426), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n427), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n428) );
  OR2X2 OR2X2_4314 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n428), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n370), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n429) );
  OR2X2 OR2X2_4315 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n430), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n421), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n431) );
  OR2X2 OR2X2_4316 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n433), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n434), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n435) );
  OR2X2 OR2X2_4317 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n435), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n432), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n436) );
  OR2X2 OR2X2_4318 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n437), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n438) );
  OR2X2 OR2X2_4319 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n439), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n440), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n441) );
  OR2X2 OR2X2_432 ( .A(AES_CORE_DATAPATH__abc_16259_n2841_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__12_), .Y(AES_CORE_DATAPATH__abc_16259_n3332_1) );
  OR2X2 OR2X2_4320 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n441), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n412), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n442) );
  OR2X2 OR2X2_4321 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n139), .B(AES_CORE_DATAPATH_MIX_COL_col_0__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n444) );
  OR2X2 OR2X2_4322 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n134_1), .B(AES_CORE_DATAPATH_MIX_COL_col_3__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n445) );
  OR2X2 OR2X2_4323 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n446), .B(AES_CORE_DATAPATH_MIX_COL_col_1__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n449) );
  OR2X2 OR2X2_4324 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n121), .B(AES_CORE_DATAPATH_MIX_COL_col_3__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n451) );
  OR2X2 OR2X2_4325 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n196), .B(AES_CORE_DATAPATH_MIX_COL_col_2__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n452) );
  OR2X2 OR2X2_4326 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n450), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n453), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n454) );
  OR2X2 OR2X2_4327 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n455), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n456), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n457) );
  OR2X2 OR2X2_4328 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n460), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n461), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n462) );
  OR2X2 OR2X2_4329 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n464), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n463), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n465) );
  OR2X2 OR2X2_433 ( .A(AES_CORE_DATAPATH__abc_16259_n3324), .B(AES_CORE_DATAPATH__abc_16259_n2853_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n3334) );
  OR2X2 OR2X2_4330 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n466), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n432), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n467) );
  OR2X2 OR2X2_4331 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n465), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n421), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n468) );
  OR2X2 OR2X2_4332 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n469), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n462), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n470) );
  OR2X2 OR2X2_4333 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n472), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n471), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n473) );
  OR2X2 OR2X2_4334 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n476), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n477), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_6_) );
  OR2X2 OR2X2_4335 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n120), .B(AES_CORE_DATAPATH_MIX_COL_col_3__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n479) );
  OR2X2 OR2X2_4336 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n196), .B(AES_CORE_DATAPATH_MIX_COL_col_0__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n480) );
  OR2X2 OR2X2_4337 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n483), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n484), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n485) );
  OR2X2 OR2X2_4338 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n485), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n251), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n486) );
  OR2X2 OR2X2_4339 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n487), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n255), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n488) );
  OR2X2 OR2X2_434 ( .A(AES_CORE_DATAPATH__abc_16259_n3335), .B(AES_CORE_DATAPATH__abc_16259_n3336), .Y(AES_CORE_DATAPATH__abc_16259_n3337) );
  OR2X2 OR2X2_4340 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n491), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n492), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n493) );
  OR2X2 OR2X2_4341 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n494), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n128), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n495) );
  OR2X2 OR2X2_4342 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n493), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n137), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n496) );
  OR2X2 OR2X2_4343 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n490), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n497), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n498) );
  OR2X2 OR2X2_4344 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n499), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n500) );
  OR2X2 OR2X2_4345 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n104), .B(AES_CORE_DATAPATH_MIX_COL_col_1__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n502) );
  OR2X2 OR2X2_4346 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n248), .B(AES_CORE_DATAPATH_MIX_COL_col_0__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n503) );
  OR2X2 OR2X2_4347 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n505), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n506), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n507) );
  OR2X2 OR2X2_4348 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n508), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n504), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n509) );
  OR2X2 OR2X2_4349 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n507), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n510), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n511) );
  OR2X2 OR2X2_435 ( .A(_auto_iopadmap_cc_313_execute_26949_12_), .B(AES_CORE_DATAPATH__abc_16259_n3339), .Y(AES_CORE_DATAPATH__abc_16259_n3340) );
  OR2X2 OR2X2_4350 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n143), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n199), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n514) );
  OR2X2 OR2X2_4351 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n150), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n203_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n515) );
  OR2X2 OR2X2_4352 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n518), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n519), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_8_) );
  OR2X2 OR2X2_4353 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n97_1), .B(AES_CORE_DATAPATH_MIX_COL_col_0__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n521) );
  OR2X2 OR2X2_4354 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n160_1), .B(AES_CORE_DATAPATH_MIX_COL_col_1__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n522) );
  OR2X2 OR2X2_4355 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n525), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n526), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n527) );
  OR2X2 OR2X2_4356 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n528), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n529), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n530) );
  OR2X2 OR2X2_4357 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n527), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n531), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n534) );
  OR2X2 OR2X2_4358 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n537), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n538), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n539) );
  OR2X2 OR2X2_4359 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n542), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n540), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_9_) );
  OR2X2 OR2X2_436 ( .A(AES_CORE_DATAPATH__abc_16259_n3342), .B(AES_CORE_DATAPATH__abc_16259_n2864_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n3343) );
  OR2X2 OR2X2_4360 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n174_1), .B(AES_CORE_DATAPATH_MIX_COL_col_0__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n544) );
  OR2X2 OR2X2_4361 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n222_1), .B(AES_CORE_DATAPATH_MIX_COL_col_1__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n545) );
  OR2X2 OR2X2_4362 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n547), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n548), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n549) );
  OR2X2 OR2X2_4363 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n550), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n546), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n551) );
  OR2X2 OR2X2_4364 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n549), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n552), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n553) );
  OR2X2 OR2X2_4365 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n264), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n302), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n556) );
  OR2X2 OR2X2_4366 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n263), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n306), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n557) );
  OR2X2 OR2X2_4367 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n558), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n555), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n559) );
  OR2X2 OR2X2_4368 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n560), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_10_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n561) );
  OR2X2 OR2X2_4369 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n563), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n564), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n565) );
  OR2X2 OR2X2_437 ( .A(AES_CORE_DATAPATH__abc_16259_n3343), .B(AES_CORE_DATAPATH__abc_16259_n3341), .Y(AES_CORE_DATAPATH__abc_16259_n3344_1) );
  OR2X2 OR2X2_4370 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n232), .B(AES_CORE_DATAPATH_MIX_COL_col_0__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n567) );
  OR2X2 OR2X2_4371 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n277), .B(AES_CORE_DATAPATH_MIX_COL_col_1__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n568) );
  OR2X2 OR2X2_4372 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n571), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n572), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n573) );
  OR2X2 OR2X2_4373 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n575), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n576), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_11_) );
  OR2X2 OR2X2_4374 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n578), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n579), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n580) );
  OR2X2 OR2X2_4375 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n314), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n377), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n583) );
  OR2X2 OR2X2_4376 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n327), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n373), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n584) );
  OR2X2 OR2X2_4377 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n581), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n586), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_11_) );
  OR2X2 OR2X2_4378 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n589), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n588), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n590) );
  OR2X2 OR2X2_4379 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n287), .B(AES_CORE_DATAPATH_MIX_COL_col_0__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n592) );
  OR2X2 OR2X2_438 ( .A(AES_CORE_DATAPATH__abc_16259_n3346_1), .B(AES_CORE_DATAPATH__abc_16259_n3345), .Y(AES_CORE_DATAPATH__abc_16259_n3347) );
  OR2X2 OR2X2_4380 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n340), .B(AES_CORE_DATAPATH_MIX_COL_col_1__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n593) );
  OR2X2 OR2X2_4381 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n596), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n597), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n598) );
  OR2X2 OR2X2_4382 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n600), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n601), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_12_) );
  OR2X2 OR2X2_4383 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n385), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n424), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n603) );
  OR2X2 OR2X2_4384 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n392), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n428), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n604) );
  OR2X2 OR2X2_4385 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n605), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_12_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n606) );
  OR2X2 OR2X2_4386 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n385), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n428), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n608) );
  OR2X2 OR2X2_4387 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n392), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n424), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n609) );
  OR2X2 OR2X2_4388 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n610), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n607), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n611) );
  OR2X2 OR2X2_4389 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n348), .B(AES_CORE_DATAPATH_MIX_COL_col_0__4_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n613) );
  OR2X2 OR2X2_439 ( .A(AES_CORE_DATAPATH__abc_16259_n3347), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n3348) );
  OR2X2 OR2X2_4390 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n405), .B(AES_CORE_DATAPATH_MIX_COL_col_1__4_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n614) );
  OR2X2 OR2X2_4391 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n616), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n617), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n618) );
  OR2X2 OR2X2_4392 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n619), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n615), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n620) );
  OR2X2 OR2X2_4393 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n618), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n621), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n622) );
  OR2X2 OR2X2_4394 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n430), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n466), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n625) );
  OR2X2 OR2X2_4395 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n435), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n465), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n626) );
  OR2X2 OR2X2_4396 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n627), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n624), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n628) );
  OR2X2 OR2X2_4397 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n435), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n466), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n629) );
  OR2X2 OR2X2_4398 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n430), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n465), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n630) );
  OR2X2 OR2X2_4399 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n631), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_13_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n632) );
  OR2X2 OR2X2_44 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n200_1), .B(AES_CORE_CONTROL_UNIT__abc_15841_n198), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n201) );
  OR2X2 OR2X2_440 ( .A(AES_CORE_DATAPATH__abc_16259_n3350), .B(AES_CORE_DATAPATH__abc_16259_n3351_1), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_12_) );
  OR2X2 OR2X2_4400 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n138), .B(AES_CORE_DATAPATH_MIX_COL_col_0__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n634) );
  OR2X2 OR2X2_4401 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n134_1), .B(AES_CORE_DATAPATH_MIX_COL_col_1__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n635) );
  OR2X2 OR2X2_4402 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n639), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n638), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n640) );
  OR2X2 OR2X2_4403 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n642), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n643), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n644) );
  OR2X2 OR2X2_4404 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n469), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n352), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n646) );
  OR2X2 OR2X2_4405 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n472), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n353), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n647) );
  OR2X2 OR2X2_4406 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n648), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n644), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n649) );
  OR2X2 OR2X2_4407 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n650), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_14_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n651) );
  OR2X2 OR2X2_4408 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n120), .B(AES_CORE_DATAPATH_MIX_COL_col_1__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n653) );
  OR2X2 OR2X2_4409 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n195_1), .B(AES_CORE_DATAPATH_MIX_COL_col_0__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n654) );
  OR2X2 OR2X2_441 ( .A(AES_CORE_DATAPATH__abc_16259_n2774_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n3353), .Y(AES_CORE_DATAPATH__abc_16259_n3354) );
  OR2X2 OR2X2_4410 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n102), .B(AES_CORE_DATAPATH_MIX_COL_col_2__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n656) );
  OR2X2 OR2X2_4411 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n190), .B(AES_CORE_DATAPATH_MIX_COL_col_3__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n657) );
  OR2X2 OR2X2_4412 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n660), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n661), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n662) );
  OR2X2 OR2X2_4413 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n663), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n655), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n664) );
  OR2X2 OR2X2_4414 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n662), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n665), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n666) );
  OR2X2 OR2X2_4415 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n494), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n132), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n669) );
  OR2X2 OR2X2_4416 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n493), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n141), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n670) );
  OR2X2 OR2X2_4417 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n671), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n667), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n672) );
  OR2X2 OR2X2_4418 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n673), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_15_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n674) );
  OR2X2 OR2X2_4419 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n676), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n677), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n678) );
  OR2X2 OR2X2_442 ( .A(AES_CORE_DATAPATH__abc_16259_n2778_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n3355_1), .Y(AES_CORE_DATAPATH__abc_16259_n3356) );
  OR2X2 OR2X2_4420 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n680), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n679), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n681) );
  OR2X2 OR2X2_4421 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n683), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n685), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_16_) );
  OR2X2 OR2X2_4422 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n688), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n689), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_16_) );
  OR2X2 OR2X2_4423 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n691), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n692), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n693) );
  OR2X2 OR2X2_4424 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n695), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n696), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n697) );
  OR2X2 OR2X2_4425 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n699), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n700), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n701) );
  OR2X2 OR2X2_4426 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n703), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n704), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n705) );
  OR2X2 OR2X2_4427 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n214_1), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_17_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n707) );
  OR2X2 OR2X2_4428 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n218_1), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n705), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n708) );
  OR2X2 OR2X2_4429 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n710), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n711), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n712) );
  OR2X2 OR2X2_443 ( .A(AES_CORE_DATAPATH__abc_16259_n3359_1), .B(AES_CORE_DATAPATH__abc_16259_n3360), .Y(AES_CORE_DATAPATH__abc_16259_n3361_1) );
  OR2X2 OR2X2_4430 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n713), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n714), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n715) );
  OR2X2 OR2X2_4431 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n715), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n712), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n716) );
  OR2X2 OR2X2_4432 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n718), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n717), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n719) );
  OR2X2 OR2X2_4433 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n270), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n721), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n722) );
  OR2X2 OR2X2_4434 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n271), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_18_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n723) );
  OR2X2 OR2X2_4435 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n725), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n726), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n727) );
  OR2X2 OR2X2_4436 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n728), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n730), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n731) );
  OR2X2 OR2X2_4437 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n594), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n285), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n732) );
  OR2X2 OR2X2_4438 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n595), .B(AES_CORE_DATAPATH_MIX_COL_col_3__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n733) );
  OR2X2 OR2X2_4439 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n731), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n734), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n737) );
  OR2X2 OR2X2_444 ( .A(AES_CORE_DATAPATH__abc_16259_n3361_1), .B(AES_CORE_DATAPATH__abc_16259_n3358), .Y(AES_CORE_DATAPATH__abc_16259_n3362) );
  OR2X2 OR2X2_4440 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n332), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_19_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n739) );
  OR2X2 OR2X2_4441 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n336), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n740), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n741) );
  OR2X2 OR2X2_4442 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n743), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n744), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n745) );
  OR2X2 OR2X2_4443 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n684), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n745), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n748) );
  OR2X2 OR2X2_4444 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n751), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n752), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n753) );
  OR2X2 OR2X2_4445 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n755), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n756), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n757) );
  OR2X2 OR2X2_4446 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n394), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n757), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n759) );
  OR2X2 OR2X2_4447 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n398), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_20_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n760) );
  OR2X2 OR2X2_4448 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n762), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n763), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n764) );
  OR2X2 OR2X2_4449 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n764), .B(AES_CORE_DATAPATH_MIX_COL_col_0__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n767) );
  OR2X2 OR2X2_445 ( .A(AES_CORE_DATAPATH__abc_16259_n3366), .B(AES_CORE_DATAPATH__abc_16259_n2826_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n3367) );
  OR2X2 OR2X2_4450 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n768), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n132), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n769) );
  OR2X2 OR2X2_4451 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n770), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n141), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n771) );
  OR2X2 OR2X2_4452 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n437), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_21_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n774) );
  OR2X2 OR2X2_4453 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n441), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n772), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n775) );
  OR2X2 OR2X2_4454 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n138), .B(AES_CORE_DATAPATH_MIX_COL_col_2__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n777) );
  OR2X2 OR2X2_4455 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n135), .B(AES_CORE_DATAPATH_MIX_COL_col_1__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n778) );
  OR2X2 OR2X2_4456 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n781), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n782), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n783) );
  OR2X2 OR2X2_4457 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n785), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n786), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_22_) );
  OR2X2 OR2X2_4458 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n789), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n790), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_22_) );
  OR2X2 OR2X2_4459 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n792), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n793), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n794) );
  OR2X2 OR2X2_446 ( .A(AES_CORE_DATAPATH__abc_16259_n3368), .B(AES_CORE_DATAPATH__abc_16259_n3369), .Y(AES_CORE_DATAPATH__abc_16259_n3370) );
  OR2X2 OR2X2_4460 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n795), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n796), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n797) );
  OR2X2 OR2X2_4461 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n798), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n794), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n801) );
  OR2X2 OR2X2_4462 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n802), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n497), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n804) );
  OR2X2 OR2X2_4463 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_23_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n499), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n805) );
  OR2X2 OR2X2_4464 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n807), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n808), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n809) );
  OR2X2 OR2X2_4465 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n811), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n812), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_24_) );
  OR2X2 OR2X2_4466 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n815), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n816), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_24_) );
  OR2X2 OR2X2_4467 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n818), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n819), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n820) );
  OR2X2 OR2X2_4468 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n659), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n820), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n823) );
  OR2X2 OR2X2_4469 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n318), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n174_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n826) );
  OR2X2 OR2X2_447 ( .A(AES_CORE_DATAPATH__abc_16259_n3370), .B(AES_CORE_DATAPATH__abc_16259_n3367), .Y(AES_CORE_DATAPATH__abc_16259_n3371) );
  OR2X2 OR2X2_4470 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n321), .B(AES_CORE_DATAPATH_MIX_COL_col_1__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n827) );
  OR2X2 OR2X2_4471 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n825), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n828), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n831) );
  OR2X2 OR2X2_4472 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n541), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n832), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n834) );
  OR2X2 OR2X2_4473 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_25_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n539), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n835) );
  OR2X2 OR2X2_4474 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n837), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n838), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n839) );
  OR2X2 OR2X2_4475 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n839), .B(AES_CORE_DATAPATH_MIX_COL_col_0__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n841) );
  OR2X2 OR2X2_4476 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n842), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n840), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n843) );
  OR2X2 OR2X2_4477 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n844), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n729), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n845) );
  OR2X2 OR2X2_4478 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n843), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n727), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n846) );
  OR2X2 OR2X2_4479 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n849), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n850), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_26_) );
  OR2X2 OR2X2_448 ( .A(AES_CORE_DATAPATH__abc_16259_n2841_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__13_), .Y(AES_CORE_DATAPATH__abc_16259_n3372) );
  OR2X2 OR2X2_4480 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n852), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n853), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n854) );
  OR2X2 OR2X2_4481 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n659), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n854), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n857) );
  OR2X2 OR2X2_4482 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n860), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n861), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n862) );
  OR2X2 OR2X2_4483 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n864), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n865), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_27_) );
  OR2X2 OR2X2_4484 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n585), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_27_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n867) );
  OR2X2 OR2X2_4485 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n580), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n868), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n869) );
  OR2X2 OR2X2_4486 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n871), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n872), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n873) );
  OR2X2 OR2X2_4487 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n875), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n876), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n877) );
  OR2X2 OR2X2_4488 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n659), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n877), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n880) );
  OR2X2 OR2X2_4489 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n883), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n884), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n885) );
  OR2X2 OR2X2_449 ( .A(AES_CORE_DATAPATH__abc_16259_n3364), .B(AES_CORE_DATAPATH__abc_16259_n2853_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n3374) );
  OR2X2 OR2X2_4490 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n605), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_28_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n887) );
  OR2X2 OR2X2_4491 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n610), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n885), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n888) );
  OR2X2 OR2X2_4492 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n890), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n891), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n892) );
  OR2X2 OR2X2_4493 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n894), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n895), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n896) );
  OR2X2 OR2X2_4494 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n896), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n893), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n897) );
  OR2X2 OR2X2_4495 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n898), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n892), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n899) );
  OR2X2 OR2X2_4496 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n627), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n900), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n902) );
  OR2X2 OR2X2_4497 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n631), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_29_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n903) );
  OR2X2 OR2X2_4498 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n905), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n906), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n907) );
  OR2X2 OR2X2_4499 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n910), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n908), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n911) );
  OR2X2 OR2X2_45 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n201), .B(AES_CORE_CONTROL_UNIT__abc_15841_n197_1), .Y(AES_CORE_CONTROL_UNIT_col_en_1_) );
  OR2X2 OR2X2_450 ( .A(AES_CORE_DATAPATH__abc_16259_n3375_1), .B(AES_CORE_DATAPATH__abc_16259_n3376), .Y(AES_CORE_DATAPATH__abc_16259_n3377) );
  OR2X2 OR2X2_4500 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n912), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n124), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n913) );
  OR2X2 OR2X2_4501 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n911), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n147_1), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n914) );
  OR2X2 OR2X2_4502 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n648), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n916), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n917) );
  OR2X2 OR2X2_4503 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n650), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_30_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n918) );
  OR2X2 OR2X2_4504 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n921), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n920), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n922) );
  OR2X2 OR2X2_4505 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n923), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n456), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n924) );
  OR2X2 OR2X2_4506 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n922), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n453), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25501_n925) );
  OR2X2 OR2X2_4507 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25501_n928), .B(AES_CORE_DATAPATH_MIX_COL__abc_25501_n929), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_31_) );
  OR2X2 OR2X2_4508 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n51_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n53_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n54_1) );
  OR2X2 OR2X2_4509 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n56), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n57) );
  OR2X2 OR2X2_451 ( .A(_auto_iopadmap_cc_313_execute_26949_13_), .B(AES_CORE_DATAPATH__abc_16259_n3379), .Y(AES_CORE_DATAPATH__abc_16259_n3380_1) );
  OR2X2 OR2X2_4510 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n58), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n59) );
  OR2X2 OR2X2_4511 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n62), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n63), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n64) );
  OR2X2 OR2X2_4512 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n69), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n68), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n70) );
  OR2X2 OR2X2_4513 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n74), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n71_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n75) );
  OR2X2 OR2X2_4514 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n76), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n65), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_4_) );
  OR2X2 OR2X2_4515 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n52), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n78) );
  OR2X2 OR2X2_4516 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n79), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n80) );
  OR2X2 OR2X2_4517 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n81), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf0), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n82) );
  OR2X2 OR2X2_4518 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n84_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n83), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n85) );
  OR2X2 OR2X2_4519 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n90), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n89), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n91) );
  OR2X2 OR2X2_452 ( .A(AES_CORE_DATAPATH__abc_16259_n3382), .B(AES_CORE_DATAPATH__abc_16259_n2864_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n3383) );
  OR2X2 OR2X2_4520 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n91), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n66_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n92) );
  OR2X2 OR2X2_4521 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n93), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n94_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n95) );
  OR2X2 OR2X2_4522 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n97_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n98), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_6_) );
  OR2X2 OR2X2_4523 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n58), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n100) );
  OR2X2 OR2X2_4524 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n79), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n101_1) );
  OR2X2 OR2X2_4525 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n105), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n106), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n107) );
  OR2X2 OR2X2_4526 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n110), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n66_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n111) );
  OR2X2 OR2X2_4527 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n111), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n108), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n112) );
  OR2X2 OR2X2_4528 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n113), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n103), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n114) );
  OR2X2 OR2X2_4529 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n75), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n118) );
  OR2X2 OR2X2_453 ( .A(AES_CORE_DATAPATH__abc_16259_n3383), .B(AES_CORE_DATAPATH__abc_16259_n3381_1), .Y(AES_CORE_DATAPATH__abc_16259_n3384_1) );
  OR2X2 OR2X2_4530 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n119), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n66_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n120) );
  OR2X2 OR2X2_4531 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n85), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n123) );
  OR2X2 OR2X2_4532 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n124), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf6), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n125) );
  OR2X2 OR2X2_4533 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n50), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n128) );
  OR2X2 OR2X2_4534 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n72), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n129) );
  OR2X2 OR2X2_4535 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n133), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf5), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n134) );
  OR2X2 OR2X2_4536 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n134), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n132), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n135) );
  OR2X2 OR2X2_4537 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n138), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n139_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n140) );
  OR2X2 OR2X2_4538 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n144), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf3), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n145_1) );
  OR2X2 OR2X2_4539 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n145_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n143_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n146_1) );
  OR2X2 OR2X2_454 ( .A(AES_CORE_DATAPATH__abc_16259_n3386_1), .B(AES_CORE_DATAPATH__abc_16259_n3385), .Y(AES_CORE_DATAPATH__abc_16259_n3387) );
  OR2X2 OR2X2_4540 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n147), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n148_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n149) );
  OR2X2 OR2X2_4541 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n152_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n66_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n153_1) );
  OR2X2 OR2X2_4542 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n153_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n151_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n154) );
  OR2X2 OR2X2_4543 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n160), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n162), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n163) );
  OR2X2 OR2X2_4544 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n165) );
  OR2X2 OR2X2_4545 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n165), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n164), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n166_1) );
  OR2X2 OR2X2_4546 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n171), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n156), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n172) );
  OR2X2 OR2X2_4547 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n178), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n167), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n179) );
  OR2X2 OR2X2_4548 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_1_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n180) );
  OR2X2 OR2X2_4549 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n179), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n181), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n182_1) );
  OR2X2 OR2X2_455 ( .A(AES_CORE_DATAPATH__abc_16259_n3387), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n3388_1) );
  OR2X2 OR2X2_4550 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n182_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n157), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n183) );
  OR2X2 OR2X2_4551 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n184), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n172), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n185) );
  OR2X2 OR2X2_4552 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n179), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n187_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n188_1) );
  OR2X2 OR2X2_4553 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n188_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n157), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n189_1) );
  OR2X2 OR2X2_4554 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n192), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n173), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n193) );
  OR2X2 OR2X2_4555 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n190_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n193), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n194) );
  OR2X2 OR2X2_4556 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n196), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n197) );
  OR2X2 OR2X2_4557 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n198), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n199) );
  OR2X2 OR2X2_4558 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n203), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n181), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n204) );
  OR2X2 OR2X2_4559 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n205), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n204), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n206) );
  OR2X2 OR2X2_456 ( .A(AES_CORE_DATAPATH__abc_16259_n3390_1), .B(AES_CORE_DATAPATH__abc_16259_n3391), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_13_) );
  OR2X2 OR2X2_4560 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n163), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n164), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n208) );
  OR2X2 OR2X2_4561 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n207), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n209), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n210) );
  OR2X2 OR2X2_4562 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n210), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n206), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n211) );
  OR2X2 OR2X2_4563 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n179), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n213), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n214) );
  OR2X2 OR2X2_4564 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n215), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n212), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n216) );
  OR2X2 OR2X2_4565 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n218), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n219) );
  OR2X2 OR2X2_4566 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n220), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n221) );
  OR2X2 OR2X2_4567 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n225), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n226), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n227) );
  OR2X2 OR2X2_4568 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n227), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n200), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n228) );
  OR2X2 OR2X2_4569 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n215), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n206), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n229) );
  OR2X2 OR2X2_457 ( .A(AES_CORE_DATAPATH__abc_16259_n2774_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n3393), .Y(AES_CORE_DATAPATH__abc_16259_n3394) );
  OR2X2 OR2X2_4570 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n210), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n212), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n230) );
  OR2X2 OR2X2_4571 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n231), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n232), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n233) );
  OR2X2 OR2X2_4572 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n217), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n201), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n234) );
  OR2X2 OR2X2_4573 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n236), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n224), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n237) );
  OR2X2 OR2X2_4574 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n238), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n239), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n240) );
  OR2X2 OR2X2_4575 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n196), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n241) );
  OR2X2 OR2X2_4576 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n218), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n242) );
  OR2X2 OR2X2_4577 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n240), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n243), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n244) );
  OR2X2 OR2X2_4578 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n245), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n244), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n248) );
  OR2X2 OR2X2_4579 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n237), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n250), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n251) );
  OR2X2 OR2X2_458 ( .A(AES_CORE_DATAPATH__abc_16259_n2778_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n3395), .Y(AES_CORE_DATAPATH__abc_16259_n3396) );
  OR2X2 OR2X2_4580 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n228), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n233), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n252) );
  OR2X2 OR2X2_4581 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n223), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n253), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n254) );
  OR2X2 OR2X2_4582 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n254), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n202), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n255) );
  OR2X2 OR2X2_4583 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n256), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n249), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n257) );
  OR2X2 OR2X2_4584 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n259), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n260) );
  OR2X2 OR2X2_4585 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n261), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n262) );
  OR2X2 OR2X2_4586 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n267), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n268) );
  OR2X2 OR2X2_4587 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n269), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n270) );
  OR2X2 OR2X2_4588 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n273), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n266), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n274) );
  OR2X2 OR2X2_4589 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n275), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n265), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n276) );
  OR2X2 OR2X2_459 ( .A(AES_CORE_DATAPATH__abc_16259_n3399), .B(AES_CORE_DATAPATH__abc_16259_n3400), .Y(AES_CORE_DATAPATH__abc_16259_n3401) );
  OR2X2 OR2X2_4590 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n278), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n181), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n279) );
  OR2X2 OR2X2_4591 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n280), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n281), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n282) );
  OR2X2 OR2X2_4592 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n279), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n282), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n283) );
  OR2X2 OR2X2_4593 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n283), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n285), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n286) );
  OR2X2 OR2X2_4594 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n184), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n206), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n287) );
  OR2X2 OR2X2_4595 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n290), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n284), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n291) );
  OR2X2 OR2X2_4596 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n277), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n293), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n294) );
  OR2X2 OR2X2_4597 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n295), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n292), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n296) );
  OR2X2 OR2X2_4598 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n269), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n298) );
  OR2X2 OR2X2_4599 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n261), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n299) );
  OR2X2 OR2X2_46 ( .A(AES_CORE_CONTROL_UNIT_state_12_), .B(AES_CORE_CONTROL_UNIT_state_1_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n203_1) );
  OR2X2 OR2X2_460 ( .A(AES_CORE_DATAPATH__abc_16259_n3401), .B(AES_CORE_DATAPATH__abc_16259_n3398), .Y(AES_CORE_DATAPATH__abc_16259_n3402_1) );
  OR2X2 OR2X2_4600 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n240), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n300), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n301) );
  OR2X2 OR2X2_4601 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n302), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n301), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n305) );
  OR2X2 OR2X2_4602 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n295), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n307), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n308) );
  OR2X2 OR2X2_4603 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n277), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n306), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n309) );
  OR2X2 OR2X2_4604 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n312), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n314), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n315) );
  OR2X2 OR2X2_4605 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n319), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n316), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_0_) );
  OR2X2 OR2X2_4606 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n322), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n324), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n325) );
  OR2X2 OR2X2_4607 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n321), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n323), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n326) );
  OR2X2 OR2X2_4608 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n329), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n244), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n332) );
  OR2X2 OR2X2_4609 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n328), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n333), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n334) );
  OR2X2 OR2X2_461 ( .A(AES_CORE_DATAPATH__abc_16259_n3406), .B(AES_CORE_DATAPATH__abc_16259_n2826_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n3407) );
  OR2X2 OR2X2_4610 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n327), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n335), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n336) );
  OR2X2 OR2X2_4611 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n339), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n340), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_5_) );
  OR2X2 OR2X2_4612 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n220), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n342) );
  OR2X2 OR2X2_4613 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n198), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n343) );
  OR2X2 OR2X2_4614 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n346), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n348), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n349) );
  OR2X2 OR2X2_4615 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n279), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n344), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n350) );
  OR2X2 OR2X2_4616 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n350), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n347), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n351) );
  OR2X2 OR2X2_4617 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n328), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n353), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n354) );
  OR2X2 OR2X2_4618 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n327), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n352), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n355) );
  OR2X2 OR2X2_4619 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n346), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n358), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n359) );
  OR2X2 OR2X2_462 ( .A(AES_CORE_DATAPATH__abc_16259_n3408), .B(AES_CORE_DATAPATH__abc_16259_n3409_1), .Y(AES_CORE_DATAPATH__abc_16259_n3410_1) );
  OR2X2 OR2X2_4620 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n350), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n360), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n361) );
  OR2X2 OR2X2_4621 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n237), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n362), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n363) );
  OR2X2 OR2X2_4622 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n346), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n360), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n364) );
  OR2X2 OR2X2_4623 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n350), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n358), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n365) );
  OR2X2 OR2X2_4624 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n256), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n366), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n367) );
  OR2X2 OR2X2_4625 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n227), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n263), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n372) );
  OR2X2 OR2X2_4626 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n231), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n272), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n373) );
  OR2X2 OR2X2_4627 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n217), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n264), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n374) );
  OR2X2 OR2X2_4628 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n376), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n371), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n377) );
  OR2X2 OR2X2_4629 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n378), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n301), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n381) );
  OR2X2 OR2X2_463 ( .A(AES_CORE_DATAPATH__abc_16259_n3410_1), .B(AES_CORE_DATAPATH__abc_16259_n3407), .Y(AES_CORE_DATAPATH__abc_16259_n3411) );
  OR2X2 OR2X2_4630 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n377), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n383), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n384) );
  OR2X2 OR2X2_4631 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n372), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n373), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n385) );
  OR2X2 OR2X2_4632 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n370), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n386), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n387) );
  OR2X2 OR2X2_4633 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n387), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n369), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n388) );
  OR2X2 OR2X2_4634 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n389), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n382), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n390) );
  OR2X2 OR2X2_4635 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n368), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n391), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n392) );
  OR2X2 OR2X2_4636 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n237), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n366), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n393) );
  OR2X2 OR2X2_4637 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n256), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n362), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n394) );
  OR2X2 OR2X2_4638 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n377), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n382), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n396) );
  OR2X2 OR2X2_4639 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n389), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n383), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n397) );
  OR2X2 OR2X2_464 ( .A(AES_CORE_DATAPATH__abc_16259_n2841_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__14_), .Y(AES_CORE_DATAPATH__abc_16259_n3412) );
  OR2X2 OR2X2_4640 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n395), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n398), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n399) );
  OR2X2 OR2X2_4641 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_7_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_1_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n402) );
  OR2X2 OR2X2_4642 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n403), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n404), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n405) );
  OR2X2 OR2X2_4643 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n405), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n356), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n406) );
  OR2X2 OR2X2_4644 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n407), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n401), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n408) );
  OR2X2 OR2X2_4645 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n409), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n410) );
  OR2X2 OR2X2_4646 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n290), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n413), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n414) );
  OR2X2 OR2X2_4647 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n283), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n412), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n415) );
  OR2X2 OR2X2_4648 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n377), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n416), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n417) );
  OR2X2 OR2X2_4649 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n290), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n412), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n418) );
  OR2X2 OR2X2_465 ( .A(AES_CORE_DATAPATH__abc_16259_n3404_1), .B(AES_CORE_DATAPATH__abc_16259_n2853_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n3414) );
  OR2X2 OR2X2_4650 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n283), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n413), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n419) );
  OR2X2 OR2X2_4651 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n389), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n420), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n421) );
  OR2X2 OR2X2_4652 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n377), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n420), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n424) );
  OR2X2 OR2X2_4653 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n389), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n416), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n425) );
  OR2X2 OR2X2_4654 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n423), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n427), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_6_) );
  OR2X2 OR2X2_4655 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_7_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n422), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n429) );
  OR2X2 OR2X2_4656 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n405), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n426), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n430) );
  OR2X2 OR2X2_4657 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n431), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n318), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n432) );
  OR2X2 OR2X2_4658 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n398), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n433) );
  OR2X2 OR2X2_4659 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n368), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n426), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n434) );
  OR2X2 OR2X2_466 ( .A(AES_CORE_DATAPATH__abc_16259_n3415_1), .B(AES_CORE_DATAPATH__abc_16259_n3416), .Y(AES_CORE_DATAPATH__abc_16259_n3417_1) );
  OR2X2 OR2X2_4660 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n395), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n422), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n435) );
  OR2X2 OR2X2_4661 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n436), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n391), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n437) );
  OR2X2 OR2X2_4662 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n315), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n439) );
  OR2X2 OR2X2_4663 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n315), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n258), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n442) );
  OR2X2 OR2X2_4664 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n443), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n407), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n444) );
  OR2X2 OR2X2_4665 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_0_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n409), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n445) );
  OR2X2 OR2X2_4666 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n431), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n401), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n447) );
  OR2X2 OR2X2_4667 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_4_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n448) );
  OR2X2 OR2X2_4668 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n449), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n356), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n450) );
  OR2X2 OR2X2_4669 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n451), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n452), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n453) );
  OR2X2 OR2X2_467 ( .A(_auto_iopadmap_cc_313_execute_26949_14_), .B(AES_CORE_DATAPATH__abc_16259_n3419_1), .Y(AES_CORE_DATAPATH__abc_16259_n3420) );
  OR2X2 OR2X2_4670 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n453), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_1_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n454) );
  OR2X2 OR2X2_4671 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n449), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n317), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n456) );
  OR2X2 OR2X2_4672 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n453), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n258), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n457) );
  OR2X2 OR2X2_4673 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n459), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n460), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n461) );
  OR2X2 OR2X2_4674 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_1_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n311), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n463) );
  OR2X2 OR2X2_4675 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n461), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n310), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n464) );
  OR2X2 OR2X2_4676 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n126_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n136), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n466) );
  OR2X2 OR2X2_4677 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_0_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n467) );
  OR2X2 OR2X2_4678 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n473), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n474), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n475) );
  OR2X2 OR2X2_4679 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n477), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n480), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n481) );
  OR2X2 OR2X2_468 ( .A(AES_CORE_DATAPATH__abc_16259_n3422), .B(AES_CORE_DATAPATH__abc_16259_n2864_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n3423) );
  OR2X2 OR2X2_4680 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n126_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n482) );
  OR2X2 OR2X2_4681 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_0_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n140), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n483) );
  OR2X2 OR2X2_4682 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n487), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n488), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n489) );
  OR2X2 OR2X2_4683 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n492) );
  OR2X2 OR2X2_4684 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n493), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n136), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n494) );
  OR2X2 OR2X2_4685 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n472), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n114), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n496) );
  OR2X2 OR2X2_4686 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n491), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n500), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n503) );
  OR2X2 OR2X2_4687 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n506), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n508), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_stage1_0_) );
  OR2X2 OR2X2_4688 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n114), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n511) );
  OR2X2 OR2X2_4689 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n516), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n517), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n518) );
  OR2X2 OR2X2_469 ( .A(AES_CORE_DATAPATH__abc_16259_n3423), .B(AES_CORE_DATAPATH__abc_16259_n3421), .Y(AES_CORE_DATAPATH__abc_16259_n3424) );
  OR2X2 OR2X2_4690 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_0_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n136), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n519) );
  OR2X2 OR2X2_4691 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n126_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n520) );
  OR2X2 OR2X2_4692 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n493), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n522) );
  OR2X2 OR2X2_4693 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n140), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n523) );
  OR2X2 OR2X2_4694 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n526), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n527), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n528) );
  OR2X2 OR2X2_4695 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n468), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n475), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n532) );
  OR2X2 OR2X2_4696 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n533), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n531), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n534) );
  OR2X2 OR2X2_4697 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n532), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n478), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n536) );
  OR2X2 OR2X2_4698 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n530), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n479), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n537) );
  OR2X2 OR2X2_4699 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n535), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n539), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n540) );
  OR2X2 OR2X2_47 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n200_1), .B(AES_CORE_CONTROL_UNIT__abc_15841_n203_1), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n204) );
  OR2X2 OR2X2_470 ( .A(AES_CORE_DATAPATH__abc_16259_n3426), .B(AES_CORE_DATAPATH__abc_16259_n3425), .Y(AES_CORE_DATAPATH__abc_16259_n3427) );
  OR2X2 OR2X2_4700 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n540), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n529), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n541) );
  OR2X2 OR2X2_4701 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n538), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n491), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n543) );
  OR2X2 OR2X2_4702 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n534), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n490), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n544) );
  OR2X2 OR2X2_4703 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n545), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n542), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n546) );
  OR2X2 OR2X2_4704 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n499), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n495), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n550) );
  OR2X2 OR2X2_4705 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n551), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n549), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n554) );
  OR2X2 OR2X2_4706 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n556), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n548), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n557) );
  OR2X2 OR2X2_4707 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n555), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n558), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n559) );
  OR2X2 OR2X2_4708 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n560), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n490), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n561) );
  OR2X2 OR2X2_4709 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n556), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n558), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n562) );
  OR2X2 OR2X2_471 ( .A(AES_CORE_DATAPATH__abc_16259_n3427), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n3428) );
  OR2X2 OR2X2_4710 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n555), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n548), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n563) );
  OR2X2 OR2X2_4711 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n564), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n491), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n565) );
  OR2X2 OR2X2_4712 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n485), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n489), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n567) );
  OR2X2 OR2X2_4713 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n571), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n572), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n573) );
  OR2X2 OR2X2_4714 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n568), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n573), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n574) );
  OR2X2 OR2X2_4715 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n575), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n567), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n576) );
  OR2X2 OR2X2_4716 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n578), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n542), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n579) );
  OR2X2 OR2X2_4717 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n577), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n529), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n580) );
  OR2X2 OR2X2_4718 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_1_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n422), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n582) );
  OR2X2 OR2X2_4719 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n583), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n426), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n584) );
  OR2X2 OR2X2_472 ( .A(AES_CORE_DATAPATH__abc_16259_n3430), .B(AES_CORE_DATAPATH__abc_16259_n3431_1), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_14_) );
  OR2X2 OR2X2_4720 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n586), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n587), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_4_) );
  OR2X2 OR2X2_4721 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n310), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n258), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n589) );
  OR2X2 OR2X2_4722 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n311), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n317), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26337_n590) );
  OR2X2 OR2X2_4723 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n51_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n53_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n54_1) );
  OR2X2 OR2X2_4724 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n56), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n57) );
  OR2X2 OR2X2_4725 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n58), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n59) );
  OR2X2 OR2X2_4726 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n62), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n63), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n64) );
  OR2X2 OR2X2_4727 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n69), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n68), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n70) );
  OR2X2 OR2X2_4728 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n74), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n71_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n75) );
  OR2X2 OR2X2_4729 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n76), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n65), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_4_) );
  OR2X2 OR2X2_473 ( .A(AES_CORE_DATAPATH__abc_16259_n2774_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n3433_1), .Y(AES_CORE_DATAPATH__abc_16259_n3434) );
  OR2X2 OR2X2_4730 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n52), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n78) );
  OR2X2 OR2X2_4731 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n79), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n80) );
  OR2X2 OR2X2_4732 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n81), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf0), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n82) );
  OR2X2 OR2X2_4733 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n84_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n83), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n85) );
  OR2X2 OR2X2_4734 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n90), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n89), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n91) );
  OR2X2 OR2X2_4735 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n91), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n66_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n92) );
  OR2X2 OR2X2_4736 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n93), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n94_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n95) );
  OR2X2 OR2X2_4737 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n97_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n98), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_6_) );
  OR2X2 OR2X2_4738 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n58), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n100) );
  OR2X2 OR2X2_4739 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n79), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n101_1) );
  OR2X2 OR2X2_474 ( .A(AES_CORE_DATAPATH__abc_16259_n2778_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n3435), .Y(AES_CORE_DATAPATH__abc_16259_n3436) );
  OR2X2 OR2X2_4740 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n105), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n106), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n107) );
  OR2X2 OR2X2_4741 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n110), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n66_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n111) );
  OR2X2 OR2X2_4742 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n111), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n108), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n112) );
  OR2X2 OR2X2_4743 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n113), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n103), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n114) );
  OR2X2 OR2X2_4744 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n75), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n118) );
  OR2X2 OR2X2_4745 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n119), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n66_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n120) );
  OR2X2 OR2X2_4746 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n85), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n123) );
  OR2X2 OR2X2_4747 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n124), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf6), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n125) );
  OR2X2 OR2X2_4748 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n50), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n128) );
  OR2X2 OR2X2_4749 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n72), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n129) );
  OR2X2 OR2X2_475 ( .A(AES_CORE_DATAPATH__abc_16259_n3439_1), .B(AES_CORE_DATAPATH__abc_16259_n3440), .Y(AES_CORE_DATAPATH__abc_16259_n3441) );
  OR2X2 OR2X2_4750 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n133), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf5), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n134) );
  OR2X2 OR2X2_4751 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n134), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n132), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n135) );
  OR2X2 OR2X2_4752 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n138), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n139_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n140) );
  OR2X2 OR2X2_4753 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n144), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf3), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n145_1) );
  OR2X2 OR2X2_4754 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n145_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n143_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n146_1) );
  OR2X2 OR2X2_4755 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n147), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n148_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n149) );
  OR2X2 OR2X2_4756 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n152_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n66_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n153_1) );
  OR2X2 OR2X2_4757 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n153_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n151_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n154) );
  OR2X2 OR2X2_4758 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n160), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n162), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n163) );
  OR2X2 OR2X2_4759 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n165) );
  OR2X2 OR2X2_476 ( .A(AES_CORE_DATAPATH__abc_16259_n3441), .B(AES_CORE_DATAPATH__abc_16259_n3438_1), .Y(AES_CORE_DATAPATH__abc_16259_n3442_1) );
  OR2X2 OR2X2_4760 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n165), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n164), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n166_1) );
  OR2X2 OR2X2_4761 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n171), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n156), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n172) );
  OR2X2 OR2X2_4762 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n178), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n167), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n179) );
  OR2X2 OR2X2_4763 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_1_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n180) );
  OR2X2 OR2X2_4764 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n179), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n181), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n182_1) );
  OR2X2 OR2X2_4765 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n182_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n157), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n183) );
  OR2X2 OR2X2_4766 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n184), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n172), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n185) );
  OR2X2 OR2X2_4767 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n179), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n187_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n188_1) );
  OR2X2 OR2X2_4768 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n188_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n157), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n189_1) );
  OR2X2 OR2X2_4769 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n192), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n173), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n193) );
  OR2X2 OR2X2_477 ( .A(AES_CORE_DATAPATH__abc_16259_n3446_1), .B(AES_CORE_DATAPATH__abc_16259_n2826_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n3447) );
  OR2X2 OR2X2_4770 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n190_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n193), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n194) );
  OR2X2 OR2X2_4771 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n196), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n197) );
  OR2X2 OR2X2_4772 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n198), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n199) );
  OR2X2 OR2X2_4773 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n203), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n181), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n204) );
  OR2X2 OR2X2_4774 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n205), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n204), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n206) );
  OR2X2 OR2X2_4775 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n163), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n164), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n208) );
  OR2X2 OR2X2_4776 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n207), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n209), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n210) );
  OR2X2 OR2X2_4777 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n210), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n206), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n211) );
  OR2X2 OR2X2_4778 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n179), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n213), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n214) );
  OR2X2 OR2X2_4779 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n215), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n212), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n216) );
  OR2X2 OR2X2_478 ( .A(AES_CORE_DATAPATH__abc_16259_n3448_1), .B(AES_CORE_DATAPATH__abc_16259_n3449), .Y(AES_CORE_DATAPATH__abc_16259_n3450) );
  OR2X2 OR2X2_4780 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n218), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n219) );
  OR2X2 OR2X2_4781 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n220), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n221) );
  OR2X2 OR2X2_4782 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n225), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n226), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n227) );
  OR2X2 OR2X2_4783 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n227), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n200), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n228) );
  OR2X2 OR2X2_4784 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n215), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n206), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n229) );
  OR2X2 OR2X2_4785 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n210), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n212), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n230) );
  OR2X2 OR2X2_4786 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n231), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n232), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n233) );
  OR2X2 OR2X2_4787 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n217), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n201), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n234) );
  OR2X2 OR2X2_4788 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n236), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n224), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n237) );
  OR2X2 OR2X2_4789 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n238), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n239), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n240) );
  OR2X2 OR2X2_479 ( .A(AES_CORE_DATAPATH__abc_16259_n3450), .B(AES_CORE_DATAPATH__abc_16259_n3447), .Y(AES_CORE_DATAPATH__abc_16259_n3451) );
  OR2X2 OR2X2_4790 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n196), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n241) );
  OR2X2 OR2X2_4791 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n218), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n242) );
  OR2X2 OR2X2_4792 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n240), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n243), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n244) );
  OR2X2 OR2X2_4793 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n245), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n244), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n248) );
  OR2X2 OR2X2_4794 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n237), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n250), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n251) );
  OR2X2 OR2X2_4795 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n228), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n233), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n252) );
  OR2X2 OR2X2_4796 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n223), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n253), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n254) );
  OR2X2 OR2X2_4797 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n254), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n202), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n255) );
  OR2X2 OR2X2_4798 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n256), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n249), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n257) );
  OR2X2 OR2X2_4799 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n259), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n260) );
  OR2X2 OR2X2_48 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n204), .B(AES_CORE_CONTROL_UNIT__abc_15841_n197_1), .Y(AES_CORE_CONTROL_UNIT_col_en_2_) );
  OR2X2 OR2X2_480 ( .A(AES_CORE_DATAPATH__abc_16259_n2841_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__15_), .Y(AES_CORE_DATAPATH__abc_16259_n3452) );
  OR2X2 OR2X2_4800 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n261), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n262) );
  OR2X2 OR2X2_4801 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n267), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n268) );
  OR2X2 OR2X2_4802 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n269), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n270) );
  OR2X2 OR2X2_4803 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n273), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n266), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n274) );
  OR2X2 OR2X2_4804 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n275), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n265), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n276) );
  OR2X2 OR2X2_4805 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n278), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n181), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n279) );
  OR2X2 OR2X2_4806 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n280), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n281), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n282) );
  OR2X2 OR2X2_4807 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n279), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n282), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n283) );
  OR2X2 OR2X2_4808 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n283), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n285), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n286) );
  OR2X2 OR2X2_4809 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n184), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n206), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n287) );
  OR2X2 OR2X2_481 ( .A(AES_CORE_DATAPATH__abc_16259_n3444_1), .B(AES_CORE_DATAPATH__abc_16259_n2853_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n3454) );
  OR2X2 OR2X2_4810 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n290), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n284), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n291) );
  OR2X2 OR2X2_4811 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n277), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n293), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n294) );
  OR2X2 OR2X2_4812 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n295), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n292), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n296) );
  OR2X2 OR2X2_4813 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n269), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n298) );
  OR2X2 OR2X2_4814 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n261), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n299) );
  OR2X2 OR2X2_4815 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n240), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n300), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n301) );
  OR2X2 OR2X2_4816 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n302), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n301), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n305) );
  OR2X2 OR2X2_4817 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n295), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n307), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n308) );
  OR2X2 OR2X2_4818 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n277), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n306), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n309) );
  OR2X2 OR2X2_4819 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n312), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n314), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n315) );
  OR2X2 OR2X2_482 ( .A(AES_CORE_DATAPATH__abc_16259_n3455), .B(AES_CORE_DATAPATH__abc_16259_n3456), .Y(AES_CORE_DATAPATH__abc_16259_n3457) );
  OR2X2 OR2X2_4820 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n319), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n316), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_8_) );
  OR2X2 OR2X2_4821 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n322), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n324), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n325) );
  OR2X2 OR2X2_4822 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n321), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n323), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n326) );
  OR2X2 OR2X2_4823 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n329), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n244), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n332) );
  OR2X2 OR2X2_4824 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n328), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n333), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n334) );
  OR2X2 OR2X2_4825 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n327), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n335), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n336) );
  OR2X2 OR2X2_4826 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n339), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n340), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_13_) );
  OR2X2 OR2X2_4827 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n220), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n342) );
  OR2X2 OR2X2_4828 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n198), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n343) );
  OR2X2 OR2X2_4829 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n346), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n348), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n349) );
  OR2X2 OR2X2_483 ( .A(_auto_iopadmap_cc_313_execute_26949_15_), .B(AES_CORE_DATAPATH__abc_16259_n3459), .Y(AES_CORE_DATAPATH__abc_16259_n3460_1) );
  OR2X2 OR2X2_4830 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n279), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n344), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n350) );
  OR2X2 OR2X2_4831 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n350), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n347), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n351) );
  OR2X2 OR2X2_4832 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n328), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n353), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n354) );
  OR2X2 OR2X2_4833 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n327), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n352), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n355) );
  OR2X2 OR2X2_4834 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n346), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n358), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n359) );
  OR2X2 OR2X2_4835 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n350), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n360), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n361) );
  OR2X2 OR2X2_4836 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n237), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n362), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n363) );
  OR2X2 OR2X2_4837 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n346), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n360), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n364) );
  OR2X2 OR2X2_4838 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n350), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n358), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n365) );
  OR2X2 OR2X2_4839 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n256), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n366), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n367) );
  OR2X2 OR2X2_484 ( .A(AES_CORE_DATAPATH__abc_16259_n3462_1), .B(AES_CORE_DATAPATH__abc_16259_n2864_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n3463) );
  OR2X2 OR2X2_4840 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n227), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n263), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n372) );
  OR2X2 OR2X2_4841 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n231), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n272), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n373) );
  OR2X2 OR2X2_4842 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n217), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n264), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n374) );
  OR2X2 OR2X2_4843 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n376), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n371), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n377) );
  OR2X2 OR2X2_4844 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n378), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n301), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n381) );
  OR2X2 OR2X2_4845 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n377), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n383), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n384) );
  OR2X2 OR2X2_4846 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n372), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n373), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n385) );
  OR2X2 OR2X2_4847 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n370), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n386), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n387) );
  OR2X2 OR2X2_4848 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n387), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n369), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n388) );
  OR2X2 OR2X2_4849 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n389), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n382), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n390) );
  OR2X2 OR2X2_485 ( .A(AES_CORE_DATAPATH__abc_16259_n3463), .B(AES_CORE_DATAPATH__abc_16259_n3461), .Y(AES_CORE_DATAPATH__abc_16259_n3464) );
  OR2X2 OR2X2_4850 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n368), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n391), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n392) );
  OR2X2 OR2X2_4851 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n237), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n366), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n393) );
  OR2X2 OR2X2_4852 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n256), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n362), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n394) );
  OR2X2 OR2X2_4853 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n377), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n382), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n396) );
  OR2X2 OR2X2_4854 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n389), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n383), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n397) );
  OR2X2 OR2X2_4855 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n395), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n398), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n399) );
  OR2X2 OR2X2_4856 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_15_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_1_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n402) );
  OR2X2 OR2X2_4857 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n403), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n404), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n405) );
  OR2X2 OR2X2_4858 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n405), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n356), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n406) );
  OR2X2 OR2X2_4859 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n407), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n401), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n408) );
  OR2X2 OR2X2_486 ( .A(AES_CORE_DATAPATH__abc_16259_n3466), .B(AES_CORE_DATAPATH__abc_16259_n3465), .Y(AES_CORE_DATAPATH__abc_16259_n3467_1) );
  OR2X2 OR2X2_4860 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n409), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_13_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n410) );
  OR2X2 OR2X2_4861 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n290), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n413), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n414) );
  OR2X2 OR2X2_4862 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n283), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n412), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n415) );
  OR2X2 OR2X2_4863 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n377), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n416), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n417) );
  OR2X2 OR2X2_4864 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n290), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n412), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n418) );
  OR2X2 OR2X2_4865 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n283), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n413), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n419) );
  OR2X2 OR2X2_4866 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n389), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n420), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n421) );
  OR2X2 OR2X2_4867 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n377), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n420), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n424) );
  OR2X2 OR2X2_4868 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n389), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n416), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n425) );
  OR2X2 OR2X2_4869 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n423), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n427), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_14_) );
  OR2X2 OR2X2_487 ( .A(AES_CORE_DATAPATH__abc_16259_n3467_1), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n3468_1) );
  OR2X2 OR2X2_4870 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_15_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n422), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n429) );
  OR2X2 OR2X2_4871 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n405), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n426), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n430) );
  OR2X2 OR2X2_4872 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n431), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n318), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n432) );
  OR2X2 OR2X2_4873 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_14_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n398), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n433) );
  OR2X2 OR2X2_4874 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n368), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n426), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n434) );
  OR2X2 OR2X2_4875 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n395), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n422), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n435) );
  OR2X2 OR2X2_4876 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n436), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n391), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n437) );
  OR2X2 OR2X2_4877 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_12_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n315), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n439) );
  OR2X2 OR2X2_4878 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n315), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n258), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n442) );
  OR2X2 OR2X2_4879 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n443), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n407), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n444) );
  OR2X2 OR2X2_488 ( .A(AES_CORE_DATAPATH__abc_16259_n3470), .B(AES_CORE_DATAPATH__abc_16259_n3471_1), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_15_) );
  OR2X2 OR2X2_4880 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_8_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n409), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n445) );
  OR2X2 OR2X2_4881 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n431), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n401), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n447) );
  OR2X2 OR2X2_4882 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_12_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_13_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n448) );
  OR2X2 OR2X2_4883 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n449), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n356), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n450) );
  OR2X2 OR2X2_4884 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n451), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n452), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n453) );
  OR2X2 OR2X2_4885 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n453), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_1_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n454) );
  OR2X2 OR2X2_4886 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n449), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n317), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n456) );
  OR2X2 OR2X2_4887 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n453), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n258), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n457) );
  OR2X2 OR2X2_4888 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n459), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n460), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n461) );
  OR2X2 OR2X2_4889 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_1_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n311), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n463) );
  OR2X2 OR2X2_489 ( .A(AES_CORE_DATAPATH__abc_16259_n2774_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n3473_1), .Y(AES_CORE_DATAPATH__abc_16259_n3474) );
  OR2X2 OR2X2_4890 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n461), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n310), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n464) );
  OR2X2 OR2X2_4891 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n126_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n136), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n466) );
  OR2X2 OR2X2_4892 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_0_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n467) );
  OR2X2 OR2X2_4893 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n473), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n474), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n475) );
  OR2X2 OR2X2_4894 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n477), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n480), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n481) );
  OR2X2 OR2X2_4895 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n126_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n482) );
  OR2X2 OR2X2_4896 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_0_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n140), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n483) );
  OR2X2 OR2X2_4897 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n487), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n488), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n489) );
  OR2X2 OR2X2_4898 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n492) );
  OR2X2 OR2X2_4899 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n493), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n136), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n494) );
  OR2X2 OR2X2_49 ( .A(AES_CORE_CONTROL_UNIT_state_9_), .B(AES_CORE_CONTROL_UNIT_state_2_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n206_1) );
  OR2X2 OR2X2_490 ( .A(AES_CORE_DATAPATH__abc_16259_n2778_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n3475_1), .Y(AES_CORE_DATAPATH__abc_16259_n3476) );
  OR2X2 OR2X2_4900 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n472), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n114), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n496) );
  OR2X2 OR2X2_4901 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n491), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n500), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n503) );
  OR2X2 OR2X2_4902 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n506), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n508), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_stage1_0_) );
  OR2X2 OR2X2_4903 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n114), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n511) );
  OR2X2 OR2X2_4904 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n516), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n517), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n518) );
  OR2X2 OR2X2_4905 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_0_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n136), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n519) );
  OR2X2 OR2X2_4906 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n126_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n520) );
  OR2X2 OR2X2_4907 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n493), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n522) );
  OR2X2 OR2X2_4908 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n140), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n523) );
  OR2X2 OR2X2_4909 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n526), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n527), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n528) );
  OR2X2 OR2X2_491 ( .A(AES_CORE_DATAPATH__abc_16259_n3479), .B(AES_CORE_DATAPATH__abc_16259_n3480), .Y(AES_CORE_DATAPATH__abc_16259_n3481) );
  OR2X2 OR2X2_4910 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n468), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n475), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n532) );
  OR2X2 OR2X2_4911 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n533), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n531), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n534) );
  OR2X2 OR2X2_4912 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n532), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n478), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n536) );
  OR2X2 OR2X2_4913 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n530), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n479), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n537) );
  OR2X2 OR2X2_4914 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n535), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n539), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n540) );
  OR2X2 OR2X2_4915 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n540), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n529), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n541) );
  OR2X2 OR2X2_4916 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n538), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n491), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n543) );
  OR2X2 OR2X2_4917 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n534), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n490), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n544) );
  OR2X2 OR2X2_4918 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n545), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n542), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n546) );
  OR2X2 OR2X2_4919 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n499), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n495), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n550) );
  OR2X2 OR2X2_492 ( .A(AES_CORE_DATAPATH__abc_16259_n3481), .B(AES_CORE_DATAPATH__abc_16259_n3478), .Y(AES_CORE_DATAPATH__abc_16259_n3482) );
  OR2X2 OR2X2_4920 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n551), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n549), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n554) );
  OR2X2 OR2X2_4921 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n556), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n548), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n557) );
  OR2X2 OR2X2_4922 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n555), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n558), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n559) );
  OR2X2 OR2X2_4923 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n560), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n490), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n561) );
  OR2X2 OR2X2_4924 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n556), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n558), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n562) );
  OR2X2 OR2X2_4925 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n555), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n548), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n563) );
  OR2X2 OR2X2_4926 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n564), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n491), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n565) );
  OR2X2 OR2X2_4927 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n485), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n489), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n567) );
  OR2X2 OR2X2_4928 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n571), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n572), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n573) );
  OR2X2 OR2X2_4929 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n568), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n573), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n574) );
  OR2X2 OR2X2_493 ( .A(AES_CORE_DATAPATH__abc_16259_n3486), .B(AES_CORE_DATAPATH__abc_16259_n2826_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n3487) );
  OR2X2 OR2X2_4930 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n575), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n567), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n576) );
  OR2X2 OR2X2_4931 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n578), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n542), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n579) );
  OR2X2 OR2X2_4932 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n577), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n529), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n580) );
  OR2X2 OR2X2_4933 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_9_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n422), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n582) );
  OR2X2 OR2X2_4934 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n583), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n426), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n584) );
  OR2X2 OR2X2_4935 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n586), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n587), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_4_) );
  OR2X2 OR2X2_4936 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n310), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n258), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n589) );
  OR2X2 OR2X2_4937 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n311), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n317), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26337_n590) );
  OR2X2 OR2X2_4938 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n51_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n53_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n54_1) );
  OR2X2 OR2X2_4939 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n56), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n57) );
  OR2X2 OR2X2_494 ( .A(AES_CORE_DATAPATH__abc_16259_n3488), .B(AES_CORE_DATAPATH__abc_16259_n3489_1), .Y(AES_CORE_DATAPATH__abc_16259_n3490) );
  OR2X2 OR2X2_4940 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n58), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n59) );
  OR2X2 OR2X2_4941 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n62), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n63), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n64) );
  OR2X2 OR2X2_4942 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n69), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n68), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n70) );
  OR2X2 OR2X2_4943 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n74), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n71_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n75) );
  OR2X2 OR2X2_4944 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n76), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n65), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_4_) );
  OR2X2 OR2X2_4945 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n52), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n78) );
  OR2X2 OR2X2_4946 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n79), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n80) );
  OR2X2 OR2X2_4947 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n81), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf0), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n82) );
  OR2X2 OR2X2_4948 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n84_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n83), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n85) );
  OR2X2 OR2X2_4949 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n90), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n89), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n91) );
  OR2X2 OR2X2_495 ( .A(AES_CORE_DATAPATH__abc_16259_n3490), .B(AES_CORE_DATAPATH__abc_16259_n3487), .Y(AES_CORE_DATAPATH__abc_16259_n3491_1) );
  OR2X2 OR2X2_4950 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n91), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n66_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n92) );
  OR2X2 OR2X2_4951 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n93), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n94_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n95) );
  OR2X2 OR2X2_4952 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n97_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n98), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_6_) );
  OR2X2 OR2X2_4953 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n58), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n100) );
  OR2X2 OR2X2_4954 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n79), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n101_1) );
  OR2X2 OR2X2_4955 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n105), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n106), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n107) );
  OR2X2 OR2X2_4956 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n110), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n66_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n111) );
  OR2X2 OR2X2_4957 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n111), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n108), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n112) );
  OR2X2 OR2X2_4958 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n113), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n103), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n114) );
  OR2X2 OR2X2_4959 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n75), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n118) );
  OR2X2 OR2X2_496 ( .A(AES_CORE_DATAPATH__abc_16259_n2841_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__16_), .Y(AES_CORE_DATAPATH__abc_16259_n3492) );
  OR2X2 OR2X2_4960 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n119), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n66_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n120) );
  OR2X2 OR2X2_4961 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n85), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n123) );
  OR2X2 OR2X2_4962 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n124), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf6), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n125) );
  OR2X2 OR2X2_4963 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n50), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n128) );
  OR2X2 OR2X2_4964 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n72), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n129) );
  OR2X2 OR2X2_4965 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n133), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf5), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n134) );
  OR2X2 OR2X2_4966 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n134), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n132), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n135) );
  OR2X2 OR2X2_4967 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n138), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n139_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n140) );
  OR2X2 OR2X2_4968 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n144), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf3), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n145_1) );
  OR2X2 OR2X2_4969 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n145_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n143_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n146_1) );
  OR2X2 OR2X2_497 ( .A(AES_CORE_DATAPATH__abc_16259_n3484), .B(AES_CORE_DATAPATH__abc_16259_n2853_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n3494) );
  OR2X2 OR2X2_4970 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n147), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n148_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n149) );
  OR2X2 OR2X2_4971 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n152_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n66_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n153_1) );
  OR2X2 OR2X2_4972 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n153_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n151_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n154) );
  OR2X2 OR2X2_4973 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n160), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n162), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n163) );
  OR2X2 OR2X2_4974 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n165) );
  OR2X2 OR2X2_4975 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n165), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n164), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n166_1) );
  OR2X2 OR2X2_4976 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n171), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n156), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n172) );
  OR2X2 OR2X2_4977 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n178), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n167), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n179) );
  OR2X2 OR2X2_4978 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_1_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n180) );
  OR2X2 OR2X2_4979 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n179), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n181), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n182_1) );
  OR2X2 OR2X2_498 ( .A(AES_CORE_DATAPATH__abc_16259_n3495), .B(AES_CORE_DATAPATH__abc_16259_n3496_1), .Y(AES_CORE_DATAPATH__abc_16259_n3497_1) );
  OR2X2 OR2X2_4980 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n182_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n157), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n183) );
  OR2X2 OR2X2_4981 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n184), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n172), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n185) );
  OR2X2 OR2X2_4982 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n179), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n187_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n188_1) );
  OR2X2 OR2X2_4983 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n188_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n157), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n189_1) );
  OR2X2 OR2X2_4984 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n192), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n173), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n193) );
  OR2X2 OR2X2_4985 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n190_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n193), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n194) );
  OR2X2 OR2X2_4986 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n196), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n197) );
  OR2X2 OR2X2_4987 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n198), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n199) );
  OR2X2 OR2X2_4988 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n203), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n181), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n204) );
  OR2X2 OR2X2_4989 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n205), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n204), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n206) );
  OR2X2 OR2X2_499 ( .A(_auto_iopadmap_cc_313_execute_26949_16_), .B(AES_CORE_DATAPATH__abc_16259_n3499), .Y(AES_CORE_DATAPATH__abc_16259_n3500_1) );
  OR2X2 OR2X2_4990 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n163), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n164), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n208) );
  OR2X2 OR2X2_4991 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n207), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n209), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n210) );
  OR2X2 OR2X2_4992 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n210), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n206), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n211) );
  OR2X2 OR2X2_4993 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n179), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n213), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n214) );
  OR2X2 OR2X2_4994 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n215), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n212), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n216) );
  OR2X2 OR2X2_4995 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n218), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n219) );
  OR2X2 OR2X2_4996 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n220), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n221) );
  OR2X2 OR2X2_4997 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n225), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n226), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n227) );
  OR2X2 OR2X2_4998 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n227), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n200), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n228) );
  OR2X2 OR2X2_4999 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n215), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n206), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n229) );
  OR2X2 OR2X2_5 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n79_1), .B(AES_CORE_CONTROL_UNIT__abc_15841_n76_1), .Y(AES_CORE_CONTROL_UNIT_encrypt_decrypt) );
  OR2X2 OR2X2_50 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n199), .B(AES_CORE_CONTROL_UNIT__abc_15841_n206_1), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n207_1) );
  OR2X2 OR2X2_500 ( .A(AES_CORE_DATAPATH__abc_16259_n3502_1), .B(AES_CORE_DATAPATH__abc_16259_n2864_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n3503) );
  OR2X2 OR2X2_5000 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n210), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n212), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n230) );
  OR2X2 OR2X2_5001 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n231), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n232), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n233) );
  OR2X2 OR2X2_5002 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n217), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n201), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n234) );
  OR2X2 OR2X2_5003 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n236), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n224), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n237) );
  OR2X2 OR2X2_5004 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n238), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n239), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n240) );
  OR2X2 OR2X2_5005 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n196), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n241) );
  OR2X2 OR2X2_5006 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n218), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n242) );
  OR2X2 OR2X2_5007 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n240), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n243), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n244) );
  OR2X2 OR2X2_5008 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n245), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n244), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n248) );
  OR2X2 OR2X2_5009 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n237), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n250), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n251) );
  OR2X2 OR2X2_501 ( .A(AES_CORE_DATAPATH__abc_16259_n3503), .B(AES_CORE_DATAPATH__abc_16259_n3501), .Y(AES_CORE_DATAPATH__abc_16259_n3504_1) );
  OR2X2 OR2X2_5010 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n228), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n233), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n252) );
  OR2X2 OR2X2_5011 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n223), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n253), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n254) );
  OR2X2 OR2X2_5012 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n254), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n202), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n255) );
  OR2X2 OR2X2_5013 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n256), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n249), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n257) );
  OR2X2 OR2X2_5014 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n259), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n260) );
  OR2X2 OR2X2_5015 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n261), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n262) );
  OR2X2 OR2X2_5016 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n267), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n268) );
  OR2X2 OR2X2_5017 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n269), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n270) );
  OR2X2 OR2X2_5018 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n273), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n266), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n274) );
  OR2X2 OR2X2_5019 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n275), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n265), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n276) );
  OR2X2 OR2X2_502 ( .A(AES_CORE_DATAPATH__abc_16259_n3506_1), .B(AES_CORE_DATAPATH__abc_16259_n3505), .Y(AES_CORE_DATAPATH__abc_16259_n3507) );
  OR2X2 OR2X2_5020 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n278), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n181), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n279) );
  OR2X2 OR2X2_5021 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n280), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n281), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n282) );
  OR2X2 OR2X2_5022 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n279), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n282), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n283) );
  OR2X2 OR2X2_5023 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n283), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n285), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n286) );
  OR2X2 OR2X2_5024 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n184), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n206), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n287) );
  OR2X2 OR2X2_5025 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n290), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n284), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n291) );
  OR2X2 OR2X2_5026 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n277), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n293), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n294) );
  OR2X2 OR2X2_5027 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n295), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n292), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n296) );
  OR2X2 OR2X2_5028 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n269), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n298) );
  OR2X2 OR2X2_5029 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n261), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n299) );
  OR2X2 OR2X2_503 ( .A(AES_CORE_DATAPATH__abc_16259_n3507), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n3508) );
  OR2X2 OR2X2_5030 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n240), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n300), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n301) );
  OR2X2 OR2X2_5031 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n302), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n301), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n305) );
  OR2X2 OR2X2_5032 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n295), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n307), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n308) );
  OR2X2 OR2X2_5033 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n277), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n306), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n309) );
  OR2X2 OR2X2_5034 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n312), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n314), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n315) );
  OR2X2 OR2X2_5035 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n319), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n316), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_16_) );
  OR2X2 OR2X2_5036 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n322), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n324), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n325) );
  OR2X2 OR2X2_5037 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n321), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n323), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n326) );
  OR2X2 OR2X2_5038 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n329), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n244), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n332) );
  OR2X2 OR2X2_5039 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n328), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n333), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n334) );
  OR2X2 OR2X2_504 ( .A(AES_CORE_DATAPATH__abc_16259_n3510), .B(AES_CORE_DATAPATH__abc_16259_n3511), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_16_) );
  OR2X2 OR2X2_5040 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n327), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n335), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n336) );
  OR2X2 OR2X2_5041 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n339), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n340), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_21_) );
  OR2X2 OR2X2_5042 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n220), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n342) );
  OR2X2 OR2X2_5043 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n198), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n343) );
  OR2X2 OR2X2_5044 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n346), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n348), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n349) );
  OR2X2 OR2X2_5045 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n279), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n344), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n350) );
  OR2X2 OR2X2_5046 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n350), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n347), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n351) );
  OR2X2 OR2X2_5047 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n328), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n353), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n354) );
  OR2X2 OR2X2_5048 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n327), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n352), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n355) );
  OR2X2 OR2X2_5049 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n346), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n358), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n359) );
  OR2X2 OR2X2_505 ( .A(AES_CORE_DATAPATH__abc_16259_n2774_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n3513), .Y(AES_CORE_DATAPATH__abc_16259_n3514) );
  OR2X2 OR2X2_5050 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n350), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n360), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n361) );
  OR2X2 OR2X2_5051 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n237), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n362), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n363) );
  OR2X2 OR2X2_5052 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n346), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n360), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n364) );
  OR2X2 OR2X2_5053 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n350), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n358), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n365) );
  OR2X2 OR2X2_5054 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n256), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n366), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n367) );
  OR2X2 OR2X2_5055 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n227), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n263), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n372) );
  OR2X2 OR2X2_5056 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n231), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n272), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n373) );
  OR2X2 OR2X2_5057 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n217), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n264), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n374) );
  OR2X2 OR2X2_5058 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n376), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n371), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n377) );
  OR2X2 OR2X2_5059 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n378), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n301), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n381) );
  OR2X2 OR2X2_506 ( .A(AES_CORE_DATAPATH__abc_16259_n2778_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n3515), .Y(AES_CORE_DATAPATH__abc_16259_n3516) );
  OR2X2 OR2X2_5060 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n377), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n383), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n384) );
  OR2X2 OR2X2_5061 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n372), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n373), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n385) );
  OR2X2 OR2X2_5062 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n370), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n386), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n387) );
  OR2X2 OR2X2_5063 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n387), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n369), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n388) );
  OR2X2 OR2X2_5064 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n389), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n382), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n390) );
  OR2X2 OR2X2_5065 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n368), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n391), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n392) );
  OR2X2 OR2X2_5066 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n237), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n366), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n393) );
  OR2X2 OR2X2_5067 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n256), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n362), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n394) );
  OR2X2 OR2X2_5068 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n377), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n382), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n396) );
  OR2X2 OR2X2_5069 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n389), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n383), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n397) );
  OR2X2 OR2X2_507 ( .A(AES_CORE_DATAPATH__abc_16259_n3519), .B(AES_CORE_DATAPATH__abc_16259_n3520_1), .Y(AES_CORE_DATAPATH__abc_16259_n3521) );
  OR2X2 OR2X2_5070 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n395), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n398), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n399) );
  OR2X2 OR2X2_5071 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_23_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_1_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n402) );
  OR2X2 OR2X2_5072 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n403), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n404), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n405) );
  OR2X2 OR2X2_5073 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n405), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n356), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n406) );
  OR2X2 OR2X2_5074 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n407), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n401), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n408) );
  OR2X2 OR2X2_5075 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n409), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_21_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n410) );
  OR2X2 OR2X2_5076 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n290), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n413), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n414) );
  OR2X2 OR2X2_5077 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n283), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n412), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n415) );
  OR2X2 OR2X2_5078 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n377), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n416), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n417) );
  OR2X2 OR2X2_5079 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n290), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n412), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n418) );
  OR2X2 OR2X2_508 ( .A(AES_CORE_DATAPATH__abc_16259_n3521), .B(AES_CORE_DATAPATH__abc_16259_n3518_1), .Y(AES_CORE_DATAPATH__abc_16259_n3522) );
  OR2X2 OR2X2_5080 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n283), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n413), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n419) );
  OR2X2 OR2X2_5081 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n389), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n420), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n421) );
  OR2X2 OR2X2_5082 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n377), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n420), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n424) );
  OR2X2 OR2X2_5083 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n389), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n416), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n425) );
  OR2X2 OR2X2_5084 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n423), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n427), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_22_) );
  OR2X2 OR2X2_5085 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_23_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n422), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n429) );
  OR2X2 OR2X2_5086 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n405), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n426), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n430) );
  OR2X2 OR2X2_5087 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n431), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n318), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n432) );
  OR2X2 OR2X2_5088 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_22_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n398), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n433) );
  OR2X2 OR2X2_5089 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n368), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n426), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n434) );
  OR2X2 OR2X2_509 ( .A(AES_CORE_DATAPATH__abc_16259_n3526_1), .B(AES_CORE_DATAPATH__abc_16259_n2826_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n3527) );
  OR2X2 OR2X2_5090 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n395), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n422), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n435) );
  OR2X2 OR2X2_5091 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n436), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n391), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n437) );
  OR2X2 OR2X2_5092 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_20_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n315), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n439) );
  OR2X2 OR2X2_5093 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n315), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n258), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n442) );
  OR2X2 OR2X2_5094 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n443), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n407), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n444) );
  OR2X2 OR2X2_5095 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_16_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n409), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n445) );
  OR2X2 OR2X2_5096 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n431), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n401), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n447) );
  OR2X2 OR2X2_5097 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_20_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_21_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n448) );
  OR2X2 OR2X2_5098 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n449), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n356), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n450) );
  OR2X2 OR2X2_5099 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n451), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n452), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n453) );
  OR2X2 OR2X2_51 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n197_1), .B(AES_CORE_CONTROL_UNIT__abc_15841_n207_1), .Y(AES_CORE_CONTROL_UNIT_col_en_3_) );
  OR2X2 OR2X2_510 ( .A(AES_CORE_DATAPATH__abc_16259_n3528), .B(AES_CORE_DATAPATH__abc_16259_n3529_1), .Y(AES_CORE_DATAPATH__abc_16259_n3530) );
  OR2X2 OR2X2_5100 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n453), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_1_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n454) );
  OR2X2 OR2X2_5101 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n449), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n317), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n456) );
  OR2X2 OR2X2_5102 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n453), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n258), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n457) );
  OR2X2 OR2X2_5103 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n459), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n460), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n461) );
  OR2X2 OR2X2_5104 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_1_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n311), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n463) );
  OR2X2 OR2X2_5105 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n461), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n310), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n464) );
  OR2X2 OR2X2_5106 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n126_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n136), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n466) );
  OR2X2 OR2X2_5107 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_0_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n467) );
  OR2X2 OR2X2_5108 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n473), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n474), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n475) );
  OR2X2 OR2X2_5109 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n477), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n480), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n481) );
  OR2X2 OR2X2_511 ( .A(AES_CORE_DATAPATH__abc_16259_n3530), .B(AES_CORE_DATAPATH__abc_16259_n3527), .Y(AES_CORE_DATAPATH__abc_16259_n3531_1) );
  OR2X2 OR2X2_5110 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n126_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n482) );
  OR2X2 OR2X2_5111 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_0_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n140), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n483) );
  OR2X2 OR2X2_5112 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n487), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n488), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n489) );
  OR2X2 OR2X2_5113 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n492) );
  OR2X2 OR2X2_5114 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n493), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n136), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n494) );
  OR2X2 OR2X2_5115 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n472), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n114), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n496) );
  OR2X2 OR2X2_5116 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n491), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n500), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n503) );
  OR2X2 OR2X2_5117 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n506), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n508), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_stage1_0_) );
  OR2X2 OR2X2_5118 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n114), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n511) );
  OR2X2 OR2X2_5119 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n516), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n517), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n518) );
  OR2X2 OR2X2_512 ( .A(AES_CORE_DATAPATH__abc_16259_n2841_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__17_), .Y(AES_CORE_DATAPATH__abc_16259_n3532) );
  OR2X2 OR2X2_5120 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_0_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n136), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n519) );
  OR2X2 OR2X2_5121 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n126_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n520) );
  OR2X2 OR2X2_5122 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n493), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n522) );
  OR2X2 OR2X2_5123 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n140), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n523) );
  OR2X2 OR2X2_5124 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n526), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n527), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n528) );
  OR2X2 OR2X2_5125 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n468), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n475), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n532) );
  OR2X2 OR2X2_5126 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n533), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n531), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n534) );
  OR2X2 OR2X2_5127 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n532), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n478), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n536) );
  OR2X2 OR2X2_5128 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n530), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n479), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n537) );
  OR2X2 OR2X2_5129 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n535), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n539), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n540) );
  OR2X2 OR2X2_513 ( .A(AES_CORE_DATAPATH__abc_16259_n3524), .B(AES_CORE_DATAPATH__abc_16259_n2853_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n3534) );
  OR2X2 OR2X2_5130 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n540), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n529), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n541) );
  OR2X2 OR2X2_5131 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n538), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n491), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n543) );
  OR2X2 OR2X2_5132 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n534), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n490), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n544) );
  OR2X2 OR2X2_5133 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n545), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n542), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n546) );
  OR2X2 OR2X2_5134 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n499), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n495), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n550) );
  OR2X2 OR2X2_5135 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n551), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n549), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n554) );
  OR2X2 OR2X2_5136 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n556), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n548), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n557) );
  OR2X2 OR2X2_5137 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n555), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n558), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n559) );
  OR2X2 OR2X2_5138 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n560), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n490), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n561) );
  OR2X2 OR2X2_5139 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n556), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n558), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n562) );
  OR2X2 OR2X2_514 ( .A(AES_CORE_DATAPATH__abc_16259_n3535_1), .B(AES_CORE_DATAPATH__abc_16259_n3536), .Y(AES_CORE_DATAPATH__abc_16259_n3537) );
  OR2X2 OR2X2_5140 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n555), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n548), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n563) );
  OR2X2 OR2X2_5141 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n564), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n491), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n565) );
  OR2X2 OR2X2_5142 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n485), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n489), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n567) );
  OR2X2 OR2X2_5143 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n571), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n572), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n573) );
  OR2X2 OR2X2_5144 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n568), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n573), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n574) );
  OR2X2 OR2X2_5145 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n575), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n567), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n576) );
  OR2X2 OR2X2_5146 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n578), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n542), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n579) );
  OR2X2 OR2X2_5147 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n577), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n529), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n580) );
  OR2X2 OR2X2_5148 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_17_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n422), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n582) );
  OR2X2 OR2X2_5149 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n583), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n426), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n584) );
  OR2X2 OR2X2_515 ( .A(_auto_iopadmap_cc_313_execute_26949_17_), .B(AES_CORE_DATAPATH__abc_16259_n3539), .Y(AES_CORE_DATAPATH__abc_16259_n3540) );
  OR2X2 OR2X2_5150 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n586), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n587), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_4_) );
  OR2X2 OR2X2_5151 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n310), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n258), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n589) );
  OR2X2 OR2X2_5152 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n311), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n317), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26337_n590) );
  OR2X2 OR2X2_5153 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n51_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n53_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n54_1) );
  OR2X2 OR2X2_5154 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n56), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n57) );
  OR2X2 OR2X2_5155 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n58), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n59) );
  OR2X2 OR2X2_5156 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n62), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n63), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n64) );
  OR2X2 OR2X2_5157 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n69), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n68), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n70) );
  OR2X2 OR2X2_5158 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n74), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n71_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n75) );
  OR2X2 OR2X2_5159 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n76), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n65), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_4_) );
  OR2X2 OR2X2_516 ( .A(AES_CORE_DATAPATH__abc_16259_n3542), .B(AES_CORE_DATAPATH__abc_16259_n2864_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n3543) );
  OR2X2 OR2X2_5160 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n52), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n78) );
  OR2X2 OR2X2_5161 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n79), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n80) );
  OR2X2 OR2X2_5162 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n81), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf0), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n82) );
  OR2X2 OR2X2_5163 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n84_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n83), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n85) );
  OR2X2 OR2X2_5164 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n90), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n89), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n91) );
  OR2X2 OR2X2_5165 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n91), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n66_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n92) );
  OR2X2 OR2X2_5166 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n93), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n94_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n95) );
  OR2X2 OR2X2_5167 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n97_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n98), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_6_) );
  OR2X2 OR2X2_5168 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n58), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n100) );
  OR2X2 OR2X2_5169 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n79), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n101_1) );
  OR2X2 OR2X2_517 ( .A(AES_CORE_DATAPATH__abc_16259_n3543), .B(AES_CORE_DATAPATH__abc_16259_n3541), .Y(AES_CORE_DATAPATH__abc_16259_n3544) );
  OR2X2 OR2X2_5170 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n105), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n106), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n107) );
  OR2X2 OR2X2_5171 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n110), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n66_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n111) );
  OR2X2 OR2X2_5172 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n111), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n108), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n112) );
  OR2X2 OR2X2_5173 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n113), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n103), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n114) );
  OR2X2 OR2X2_5174 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n75), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n118) );
  OR2X2 OR2X2_5175 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n119), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n66_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n120) );
  OR2X2 OR2X2_5176 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n85), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n123) );
  OR2X2 OR2X2_5177 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n124), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf6), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n125) );
  OR2X2 OR2X2_5178 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n50), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n128) );
  OR2X2 OR2X2_5179 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n72), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n129) );
  OR2X2 OR2X2_518 ( .A(AES_CORE_DATAPATH__abc_16259_n3546), .B(AES_CORE_DATAPATH__abc_16259_n3545), .Y(AES_CORE_DATAPATH__abc_16259_n3547_1) );
  OR2X2 OR2X2_5180 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n133), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf5), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n134) );
  OR2X2 OR2X2_5181 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n134), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n132), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n135) );
  OR2X2 OR2X2_5182 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n138), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n139_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n140) );
  OR2X2 OR2X2_5183 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n144), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec_bF_buf3), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n145_1) );
  OR2X2 OR2X2_5184 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n145_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n143_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n146_1) );
  OR2X2 OR2X2_5185 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n147), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n148_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n149) );
  OR2X2 OR2X2_5186 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n152_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n66_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n153_1) );
  OR2X2 OR2X2_5187 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n153_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n151_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n154) );
  OR2X2 OR2X2_5188 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n160), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n162), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n163) );
  OR2X2 OR2X2_5189 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n165) );
  OR2X2 OR2X2_519 ( .A(AES_CORE_DATAPATH__abc_16259_n3547_1), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n3548) );
  OR2X2 OR2X2_5190 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n165), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n164), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n166_1) );
  OR2X2 OR2X2_5191 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n171), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n156), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n172) );
  OR2X2 OR2X2_5192 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n178), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n167), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n179) );
  OR2X2 OR2X2_5193 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_1_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n180) );
  OR2X2 OR2X2_5194 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n179), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n181), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n182_1) );
  OR2X2 OR2X2_5195 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n182_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n157), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n183) );
  OR2X2 OR2X2_5196 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n184), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n172), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n185) );
  OR2X2 OR2X2_5197 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n179), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n187_1), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n188_1) );
  OR2X2 OR2X2_5198 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n188_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n157), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n189_1) );
  OR2X2 OR2X2_5199 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n192), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n173), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n193) );
  OR2X2 OR2X2_52 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n210_1), .B(AES_CORE_CONTROL_UNIT__abc_15841_n137), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n211_1) );
  OR2X2 OR2X2_520 ( .A(AES_CORE_DATAPATH__abc_16259_n3550), .B(AES_CORE_DATAPATH__abc_16259_n3551), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_17_) );
  OR2X2 OR2X2_5200 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n190_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n193), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n194) );
  OR2X2 OR2X2_5201 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n196), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n197) );
  OR2X2 OR2X2_5202 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n198), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n199) );
  OR2X2 OR2X2_5203 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n203), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n181), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n204) );
  OR2X2 OR2X2_5204 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n205), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n204), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n206) );
  OR2X2 OR2X2_5205 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n163), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n164), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n208) );
  OR2X2 OR2X2_5206 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n207), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n209), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n210) );
  OR2X2 OR2X2_5207 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n210), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n206), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n211) );
  OR2X2 OR2X2_5208 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n179), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n213), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n214) );
  OR2X2 OR2X2_5209 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n215), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n212), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n216) );
  OR2X2 OR2X2_521 ( .A(AES_CORE_DATAPATH__abc_16259_n2774_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n3553), .Y(AES_CORE_DATAPATH__abc_16259_n3554_1) );
  OR2X2 OR2X2_5210 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n218), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n219) );
  OR2X2 OR2X2_5211 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n220), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n221) );
  OR2X2 OR2X2_5212 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n225), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n226), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n227) );
  OR2X2 OR2X2_5213 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n227), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n200), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n228) );
  OR2X2 OR2X2_5214 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n215), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n206), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n229) );
  OR2X2 OR2X2_5215 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n210), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n212), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n230) );
  OR2X2 OR2X2_5216 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n231), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n232), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n233) );
  OR2X2 OR2X2_5217 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n217), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n201), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n234) );
  OR2X2 OR2X2_5218 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n236), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n224), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n237) );
  OR2X2 OR2X2_5219 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n238), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n239), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n240) );
  OR2X2 OR2X2_522 ( .A(AES_CORE_DATAPATH__abc_16259_n2778_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n3555_1), .Y(AES_CORE_DATAPATH__abc_16259_n3556) );
  OR2X2 OR2X2_5220 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n196), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n241) );
  OR2X2 OR2X2_5221 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n218), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n242) );
  OR2X2 OR2X2_5222 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n240), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n243), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n244) );
  OR2X2 OR2X2_5223 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n245), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n244), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n248) );
  OR2X2 OR2X2_5224 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n237), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n250), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n251) );
  OR2X2 OR2X2_5225 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n228), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n233), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n252) );
  OR2X2 OR2X2_5226 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n223), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n253), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n254) );
  OR2X2 OR2X2_5227 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n254), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n202), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n255) );
  OR2X2 OR2X2_5228 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n256), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n249), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n257) );
  OR2X2 OR2X2_5229 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n259), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n260) );
  OR2X2 OR2X2_523 ( .A(AES_CORE_DATAPATH__abc_16259_n3559), .B(AES_CORE_DATAPATH__abc_16259_n3560_1), .Y(AES_CORE_DATAPATH__abc_16259_n3561) );
  OR2X2 OR2X2_5230 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n261), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n262) );
  OR2X2 OR2X2_5231 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n267), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n268) );
  OR2X2 OR2X2_5232 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n269), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n270) );
  OR2X2 OR2X2_5233 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n273), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n266), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n274) );
  OR2X2 OR2X2_5234 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n275), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n265), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n276) );
  OR2X2 OR2X2_5235 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n278), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n181), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n279) );
  OR2X2 OR2X2_5236 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n280), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n281), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n282) );
  OR2X2 OR2X2_5237 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n279), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n282), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n283) );
  OR2X2 OR2X2_5238 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n283), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n285), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n286) );
  OR2X2 OR2X2_5239 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n184), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n206), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n287) );
  OR2X2 OR2X2_524 ( .A(AES_CORE_DATAPATH__abc_16259_n3561), .B(AES_CORE_DATAPATH__abc_16259_n3558_1), .Y(AES_CORE_DATAPATH__abc_16259_n3562_1) );
  OR2X2 OR2X2_5240 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n290), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n284), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n291) );
  OR2X2 OR2X2_5241 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n277), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n293), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n294) );
  OR2X2 OR2X2_5242 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n295), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n292), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n296) );
  OR2X2 OR2X2_5243 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n269), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n298) );
  OR2X2 OR2X2_5244 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n261), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n299) );
  OR2X2 OR2X2_5245 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n240), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n300), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n301) );
  OR2X2 OR2X2_5246 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n302), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n301), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n305) );
  OR2X2 OR2X2_5247 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n295), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n307), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n308) );
  OR2X2 OR2X2_5248 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n277), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n306), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n309) );
  OR2X2 OR2X2_5249 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n312), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n314), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n315) );
  OR2X2 OR2X2_525 ( .A(AES_CORE_DATAPATH__abc_16259_n3566), .B(AES_CORE_DATAPATH__abc_16259_n2826_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n3567) );
  OR2X2 OR2X2_5250 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n319), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n316), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_24_) );
  OR2X2 OR2X2_5251 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n322), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n324), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n325) );
  OR2X2 OR2X2_5252 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n321), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n323), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n326) );
  OR2X2 OR2X2_5253 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n329), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n244), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n332) );
  OR2X2 OR2X2_5254 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n328), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n333), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n334) );
  OR2X2 OR2X2_5255 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n327), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n335), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n336) );
  OR2X2 OR2X2_5256 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n339), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n340), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_29_) );
  OR2X2 OR2X2_5257 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n220), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n342) );
  OR2X2 OR2X2_5258 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n198), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n343) );
  OR2X2 OR2X2_5259 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n346), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n348), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n349) );
  OR2X2 OR2X2_526 ( .A(AES_CORE_DATAPATH__abc_16259_n3568), .B(AES_CORE_DATAPATH__abc_16259_n3569), .Y(AES_CORE_DATAPATH__abc_16259_n3570) );
  OR2X2 OR2X2_5260 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n279), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n344), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n350) );
  OR2X2 OR2X2_5261 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n350), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n347), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n351) );
  OR2X2 OR2X2_5262 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n328), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n353), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n354) );
  OR2X2 OR2X2_5263 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n327), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n352), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n355) );
  OR2X2 OR2X2_5264 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n346), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n358), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n359) );
  OR2X2 OR2X2_5265 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n350), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n360), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n361) );
  OR2X2 OR2X2_5266 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n237), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n362), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n363) );
  OR2X2 OR2X2_5267 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n346), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n360), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n364) );
  OR2X2 OR2X2_5268 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n350), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n358), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n365) );
  OR2X2 OR2X2_5269 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n256), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n366), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n367) );
  OR2X2 OR2X2_527 ( .A(AES_CORE_DATAPATH__abc_16259_n3570), .B(AES_CORE_DATAPATH__abc_16259_n3567), .Y(AES_CORE_DATAPATH__abc_16259_n3571) );
  OR2X2 OR2X2_5270 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n227), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n263), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n372) );
  OR2X2 OR2X2_5271 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n231), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n272), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n373) );
  OR2X2 OR2X2_5272 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n217), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n264), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n374) );
  OR2X2 OR2X2_5273 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n376), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n371), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n377) );
  OR2X2 OR2X2_5274 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n378), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n301), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n381) );
  OR2X2 OR2X2_5275 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n377), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n383), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n384) );
  OR2X2 OR2X2_5276 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n372), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n373), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n385) );
  OR2X2 OR2X2_5277 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n370), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n386), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n387) );
  OR2X2 OR2X2_5278 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n387), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n369), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n388) );
  OR2X2 OR2X2_5279 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n389), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n382), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n390) );
  OR2X2 OR2X2_528 ( .A(AES_CORE_DATAPATH__abc_16259_n2841_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__18_), .Y(AES_CORE_DATAPATH__abc_16259_n3572) );
  OR2X2 OR2X2_5280 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n368), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n391), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n392) );
  OR2X2 OR2X2_5281 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n237), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n366), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n393) );
  OR2X2 OR2X2_5282 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n256), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n362), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n394) );
  OR2X2 OR2X2_5283 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n377), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n382), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n396) );
  OR2X2 OR2X2_5284 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n389), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n383), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n397) );
  OR2X2 OR2X2_5285 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n395), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n398), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n399) );
  OR2X2 OR2X2_5286 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_31_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_1_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n402) );
  OR2X2 OR2X2_5287 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n403), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n404), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n405) );
  OR2X2 OR2X2_5288 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n405), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n356), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n406) );
  OR2X2 OR2X2_5289 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n407), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n401), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n408) );
  OR2X2 OR2X2_529 ( .A(AES_CORE_DATAPATH__abc_16259_n3564_1), .B(AES_CORE_DATAPATH__abc_16259_n2853_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n3574) );
  OR2X2 OR2X2_5290 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n409), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_29_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n410) );
  OR2X2 OR2X2_5291 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n290), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n413), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n414) );
  OR2X2 OR2X2_5292 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n283), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n412), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n415) );
  OR2X2 OR2X2_5293 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n377), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n416), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n417) );
  OR2X2 OR2X2_5294 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n290), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n412), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n418) );
  OR2X2 OR2X2_5295 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n283), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n413), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n419) );
  OR2X2 OR2X2_5296 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n389), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n420), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n421) );
  OR2X2 OR2X2_5297 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n377), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n420), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n424) );
  OR2X2 OR2X2_5298 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n389), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n416), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n425) );
  OR2X2 OR2X2_5299 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n423), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n427), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_30_) );
  OR2X2 OR2X2_53 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n211_1), .B(AES_CORE_CONTROL_UNIT__abc_15841_n209_1), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n212_1) );
  OR2X2 OR2X2_530 ( .A(AES_CORE_DATAPATH__abc_16259_n3575), .B(AES_CORE_DATAPATH__abc_16259_n3576_1), .Y(AES_CORE_DATAPATH__abc_16259_n3577) );
  OR2X2 OR2X2_5300 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_31_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n422), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n429) );
  OR2X2 OR2X2_5301 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n405), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n426), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n430) );
  OR2X2 OR2X2_5302 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n431), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n318), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n432) );
  OR2X2 OR2X2_5303 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_30_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n398), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n433) );
  OR2X2 OR2X2_5304 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n368), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n426), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n434) );
  OR2X2 OR2X2_5305 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n395), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n422), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n435) );
  OR2X2 OR2X2_5306 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n436), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n391), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n437) );
  OR2X2 OR2X2_5307 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_28_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n315), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n439) );
  OR2X2 OR2X2_5308 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n315), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n258), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n442) );
  OR2X2 OR2X2_5309 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n443), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n407), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n444) );
  OR2X2 OR2X2_531 ( .A(_auto_iopadmap_cc_313_execute_26949_18_), .B(AES_CORE_DATAPATH__abc_16259_n3579), .Y(AES_CORE_DATAPATH__abc_16259_n3580) );
  OR2X2 OR2X2_5310 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_24_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n409), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n445) );
  OR2X2 OR2X2_5311 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n431), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n401), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n447) );
  OR2X2 OR2X2_5312 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_28_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_29_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n448) );
  OR2X2 OR2X2_5313 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n449), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n356), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n450) );
  OR2X2 OR2X2_5314 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n451), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n452), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n453) );
  OR2X2 OR2X2_5315 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n453), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_1_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n454) );
  OR2X2 OR2X2_5316 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n449), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n317), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n456) );
  OR2X2 OR2X2_5317 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n453), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n258), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n457) );
  OR2X2 OR2X2_5318 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n459), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n460), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n461) );
  OR2X2 OR2X2_5319 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_1_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n311), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n463) );
  OR2X2 OR2X2_532 ( .A(AES_CORE_DATAPATH__abc_16259_n3582), .B(AES_CORE_DATAPATH__abc_16259_n2864_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n3583_1) );
  OR2X2 OR2X2_5320 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n461), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n310), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n464) );
  OR2X2 OR2X2_5321 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n126_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n136), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n466) );
  OR2X2 OR2X2_5322 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_0_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n467) );
  OR2X2 OR2X2_5323 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n473), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n474), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n475) );
  OR2X2 OR2X2_5324 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n477), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n480), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n481) );
  OR2X2 OR2X2_5325 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n126_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n482) );
  OR2X2 OR2X2_5326 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_0_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n140), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n483) );
  OR2X2 OR2X2_5327 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n487), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n488), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n489) );
  OR2X2 OR2X2_5328 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n492) );
  OR2X2 OR2X2_5329 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n493), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n136), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n494) );
  OR2X2 OR2X2_533 ( .A(AES_CORE_DATAPATH__abc_16259_n3583_1), .B(AES_CORE_DATAPATH__abc_16259_n3581), .Y(AES_CORE_DATAPATH__abc_16259_n3584_1) );
  OR2X2 OR2X2_5330 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n472), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n114), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n496) );
  OR2X2 OR2X2_5331 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n491), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n500), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n503) );
  OR2X2 OR2X2_5332 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n506), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n508), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_stage1_0_) );
  OR2X2 OR2X2_5333 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n114), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n511) );
  OR2X2 OR2X2_5334 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n516), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n517), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n518) );
  OR2X2 OR2X2_5335 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_0_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n136), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n519) );
  OR2X2 OR2X2_5336 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n126_1), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n520) );
  OR2X2 OR2X2_5337 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n493), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n522) );
  OR2X2 OR2X2_5338 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n140), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n523) );
  OR2X2 OR2X2_5339 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n526), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n527), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n528) );
  OR2X2 OR2X2_534 ( .A(AES_CORE_DATAPATH__abc_16259_n3586), .B(AES_CORE_DATAPATH__abc_16259_n3585), .Y(AES_CORE_DATAPATH__abc_16259_n3587_1) );
  OR2X2 OR2X2_5340 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n468), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n475), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n532) );
  OR2X2 OR2X2_5341 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n533), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n531), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n534) );
  OR2X2 OR2X2_5342 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n532), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n478), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n536) );
  OR2X2 OR2X2_5343 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n530), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n479), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n537) );
  OR2X2 OR2X2_5344 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n535), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n539), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n540) );
  OR2X2 OR2X2_5345 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n540), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n529), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n541) );
  OR2X2 OR2X2_5346 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n538), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n491), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n543) );
  OR2X2 OR2X2_5347 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n534), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n490), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n544) );
  OR2X2 OR2X2_5348 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n545), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n542), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n546) );
  OR2X2 OR2X2_5349 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n499), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n495), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n550) );
  OR2X2 OR2X2_535 ( .A(AES_CORE_DATAPATH__abc_16259_n3587_1), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n3588) );
  OR2X2 OR2X2_5350 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n551), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n549), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n554) );
  OR2X2 OR2X2_5351 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n556), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n548), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n557) );
  OR2X2 OR2X2_5352 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n555), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n558), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n559) );
  OR2X2 OR2X2_5353 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n560), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n490), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n561) );
  OR2X2 OR2X2_5354 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n556), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n558), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n562) );
  OR2X2 OR2X2_5355 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n555), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n548), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n563) );
  OR2X2 OR2X2_5356 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n564), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n491), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n565) );
  OR2X2 OR2X2_5357 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n485), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n489), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n567) );
  OR2X2 OR2X2_5358 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n571), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n572), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n573) );
  OR2X2 OR2X2_5359 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n568), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n573), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n574) );
  OR2X2 OR2X2_536 ( .A(AES_CORE_DATAPATH__abc_16259_n3590), .B(AES_CORE_DATAPATH__abc_16259_n3591_1), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_18_) );
  OR2X2 OR2X2_5360 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n575), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n567), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n576) );
  OR2X2 OR2X2_5361 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n578), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n542), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n579) );
  OR2X2 OR2X2_5362 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n577), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n529), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n580) );
  OR2X2 OR2X2_5363 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_25_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n422), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n582) );
  OR2X2 OR2X2_5364 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n583), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n426), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n584) );
  OR2X2 OR2X2_5365 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n586), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n587), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_4_) );
  OR2X2 OR2X2_5366 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n310), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n258), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n589) );
  OR2X2 OR2X2_5367 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n311), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n317), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26337_n590) );
  OR2X2 OR2X2_5368 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n71_1), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n68), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n72_1) );
  OR2X2 OR2X2_5369 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n75), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n77_1), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n78) );
  OR2X2 OR2X2_537 ( .A(AES_CORE_DATAPATH__abc_16259_n2774_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n3593_1), .Y(AES_CORE_DATAPATH__abc_16259_n3594) );
  OR2X2 OR2X2_5370 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n78), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n72_1), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_0_) );
  OR2X2 OR2X2_5371 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n81_1), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n80), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n82_1) );
  OR2X2 OR2X2_5372 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n83), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n84), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n85) );
  OR2X2 OR2X2_5373 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n85), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n82_1), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_1_) );
  OR2X2 OR2X2_5374 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n88), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n87_1), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n89) );
  OR2X2 OR2X2_5375 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n90), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n91_1), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n92_1) );
  OR2X2 OR2X2_5376 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n92_1), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n89), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_2_) );
  OR2X2 OR2X2_5377 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n95), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n94), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n96_1) );
  OR2X2 OR2X2_5378 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n97_1), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n98), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n99) );
  OR2X2 OR2X2_5379 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n99), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n96_1), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_3_) );
  OR2X2 OR2X2_538 ( .A(AES_CORE_DATAPATH__abc_16259_n2778_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n3595), .Y(AES_CORE_DATAPATH__abc_16259_n3596) );
  OR2X2 OR2X2_5380 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n102_1), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n101_1), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n103) );
  OR2X2 OR2X2_5381 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n104), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n105), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n106_1) );
  OR2X2 OR2X2_5382 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n106_1), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n103), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_4_) );
  OR2X2 OR2X2_5383 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n109), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n108), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n110_1) );
  OR2X2 OR2X2_5384 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n111), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n112), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n113) );
  OR2X2 OR2X2_5385 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n113), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n110_1), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_5_) );
  OR2X2 OR2X2_5386 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n116), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n115), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n117) );
  OR2X2 OR2X2_5387 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n118_1), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n119), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n120) );
  OR2X2 OR2X2_5388 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n120), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n117), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_6_) );
  OR2X2 OR2X2_5389 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n123), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n122_1), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n124) );
  OR2X2 OR2X2_539 ( .A(AES_CORE_DATAPATH__abc_16259_n3599), .B(AES_CORE_DATAPATH__abc_16259_n3600), .Y(AES_CORE_DATAPATH__abc_16259_n3601) );
  OR2X2 OR2X2_5390 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n125), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n126_1), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n127) );
  OR2X2 OR2X2_5391 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n127), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n124), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_7_) );
  OR2X2 OR2X2_5392 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n130_1), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n129), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n131) );
  OR2X2 OR2X2_5393 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n132), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n133), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n134_1) );
  OR2X2 OR2X2_5394 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n134_1), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n131), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_8_) );
  OR2X2 OR2X2_5395 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n137), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n136), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n138_1) );
  OR2X2 OR2X2_5396 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n139), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n140), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n141) );
  OR2X2 OR2X2_5397 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n141), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n138_1), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_9_) );
  OR2X2 OR2X2_5398 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n144), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n143), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n145) );
  OR2X2 OR2X2_5399 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n146_1), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n147), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n148) );
  OR2X2 OR2X2_54 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n215), .B(AES_CORE_CONTROL_UNIT__abc_15841_n213), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n216) );
  OR2X2 OR2X2_540 ( .A(AES_CORE_DATAPATH__abc_16259_n3601), .B(AES_CORE_DATAPATH__abc_16259_n3598), .Y(AES_CORE_DATAPATH__abc_16259_n3602) );
  OR2X2 OR2X2_5400 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n148), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n145), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_10_) );
  OR2X2 OR2X2_5401 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n151), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n150_1), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n152) );
  OR2X2 OR2X2_5402 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n153), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n154_1), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n155) );
  OR2X2 OR2X2_5403 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n155), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n152), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_11_) );
  OR2X2 OR2X2_5404 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n158_1), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n157), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n159) );
  OR2X2 OR2X2_5405 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n160), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n161), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n162_1) );
  OR2X2 OR2X2_5406 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n162_1), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n159), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_12_) );
  OR2X2 OR2X2_5407 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n165), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n164), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n166_1) );
  OR2X2 OR2X2_5408 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n167), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n168), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n169) );
  OR2X2 OR2X2_5409 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n169), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n166_1), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_13_) );
  OR2X2 OR2X2_541 ( .A(AES_CORE_DATAPATH__abc_16259_n3606), .B(AES_CORE_DATAPATH__abc_16259_n2826_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n3607_1) );
  OR2X2 OR2X2_5410 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n172), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n171), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n173) );
  OR2X2 OR2X2_5411 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n174), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n175), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n176) );
  OR2X2 OR2X2_5412 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n176), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n173), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_14_) );
  OR2X2 OR2X2_5413 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n179), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n178), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n180) );
  OR2X2 OR2X2_5414 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n181), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n182), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n183) );
  OR2X2 OR2X2_5415 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n183), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n180), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_15_) );
  OR2X2 OR2X2_5416 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n186), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n185), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n187) );
  OR2X2 OR2X2_5417 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n188), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n189), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n190) );
  OR2X2 OR2X2_5418 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n190), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n187), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_16_) );
  OR2X2 OR2X2_5419 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n193), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n192), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n194) );
  OR2X2 OR2X2_542 ( .A(AES_CORE_DATAPATH__abc_16259_n3608), .B(AES_CORE_DATAPATH__abc_16259_n3609), .Y(AES_CORE_DATAPATH__abc_16259_n3610) );
  OR2X2 OR2X2_5420 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n195), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n196), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n197) );
  OR2X2 OR2X2_5421 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n197), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n194), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_17_) );
  OR2X2 OR2X2_5422 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n200), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n199), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n201) );
  OR2X2 OR2X2_5423 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n202), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n203), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n204) );
  OR2X2 OR2X2_5424 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n204), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n201), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_18_) );
  OR2X2 OR2X2_5425 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n207), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n206), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n208) );
  OR2X2 OR2X2_5426 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n209), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n210), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n211) );
  OR2X2 OR2X2_5427 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n211), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n208), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_19_) );
  OR2X2 OR2X2_5428 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n214), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n213), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n215) );
  OR2X2 OR2X2_5429 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n216), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n217), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n218) );
  OR2X2 OR2X2_543 ( .A(AES_CORE_DATAPATH__abc_16259_n3610), .B(AES_CORE_DATAPATH__abc_16259_n3607_1), .Y(AES_CORE_DATAPATH__abc_16259_n3611) );
  OR2X2 OR2X2_5430 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n218), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n215), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_20_) );
  OR2X2 OR2X2_5431 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n221), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n220), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n222) );
  OR2X2 OR2X2_5432 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n223), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n224), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n225) );
  OR2X2 OR2X2_5433 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n225), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n222), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_21_) );
  OR2X2 OR2X2_5434 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n228), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n227), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n229) );
  OR2X2 OR2X2_5435 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n230), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n231), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n232) );
  OR2X2 OR2X2_5436 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n232), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n229), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_22_) );
  OR2X2 OR2X2_5437 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n235), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n234), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n236) );
  OR2X2 OR2X2_5438 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n237), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n238), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n239) );
  OR2X2 OR2X2_5439 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n239), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n236), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_23_) );
  OR2X2 OR2X2_544 ( .A(AES_CORE_DATAPATH__abc_16259_n2841_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__19_), .Y(AES_CORE_DATAPATH__abc_16259_n3612_1) );
  OR2X2 OR2X2_5440 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n242), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n241), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n243) );
  OR2X2 OR2X2_5441 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n244), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n245), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n246) );
  OR2X2 OR2X2_5442 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n246), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n243), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_24_) );
  OR2X2 OR2X2_5443 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n249), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n248), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n250) );
  OR2X2 OR2X2_5444 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n251), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n252), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n253) );
  OR2X2 OR2X2_5445 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n253), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n250), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_25_) );
  OR2X2 OR2X2_5446 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n256), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n255), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n257) );
  OR2X2 OR2X2_5447 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n258), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n259), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n260) );
  OR2X2 OR2X2_5448 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n260), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n257), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_26_) );
  OR2X2 OR2X2_5449 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n263), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n262), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n264) );
  OR2X2 OR2X2_545 ( .A(AES_CORE_DATAPATH__abc_16259_n3604), .B(AES_CORE_DATAPATH__abc_16259_n2853_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n3614) );
  OR2X2 OR2X2_5450 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n265), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n266), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n267) );
  OR2X2 OR2X2_5451 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n267), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n264), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_27_) );
  OR2X2 OR2X2_5452 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n270), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n269), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n271) );
  OR2X2 OR2X2_5453 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n272), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n273), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n274) );
  OR2X2 OR2X2_5454 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n274), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n271), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_28_) );
  OR2X2 OR2X2_5455 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n277), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n276), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n278) );
  OR2X2 OR2X2_5456 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n279), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n280), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n281) );
  OR2X2 OR2X2_5457 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n281), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n278), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_29_) );
  OR2X2 OR2X2_5458 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n284), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n283), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n285) );
  OR2X2 OR2X2_5459 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n286), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n287), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n288) );
  OR2X2 OR2X2_546 ( .A(AES_CORE_DATAPATH__abc_16259_n3615), .B(AES_CORE_DATAPATH__abc_16259_n3616_1), .Y(AES_CORE_DATAPATH__abc_16259_n3617) );
  OR2X2 OR2X2_5460 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n288), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n285), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_30_) );
  OR2X2 OR2X2_5461 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n291), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n290), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n292) );
  OR2X2 OR2X2_5462 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n293), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n294), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n295) );
  OR2X2 OR2X2_5463 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n295), .B(AES_CORE_DATAPATH_SWAP_IN__abc_16028_n292), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_31_) );
  OR2X2 OR2X2_5464 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n71_1), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n68), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n72_1) );
  OR2X2 OR2X2_5465 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n75), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n77_1), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n78) );
  OR2X2 OR2X2_5466 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n78), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n72_1), .Y(_auto_iopadmap_cc_313_execute_26881_0_) );
  OR2X2 OR2X2_5467 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n81_1), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n80), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n82_1) );
  OR2X2 OR2X2_5468 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n83), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n84), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n85) );
  OR2X2 OR2X2_5469 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n85), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n82_1), .Y(_auto_iopadmap_cc_313_execute_26881_1_) );
  OR2X2 OR2X2_547 ( .A(_auto_iopadmap_cc_313_execute_26949_19_), .B(AES_CORE_DATAPATH__abc_16259_n3619), .Y(AES_CORE_DATAPATH__abc_16259_n3620_1) );
  OR2X2 OR2X2_5470 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n88), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n87_1), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n89) );
  OR2X2 OR2X2_5471 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n90), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n91_1), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n92_1) );
  OR2X2 OR2X2_5472 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n92_1), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n89), .Y(_auto_iopadmap_cc_313_execute_26881_2_) );
  OR2X2 OR2X2_5473 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n95), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n94), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n96_1) );
  OR2X2 OR2X2_5474 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n97_1), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n98), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n99) );
  OR2X2 OR2X2_5475 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n99), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n96_1), .Y(_auto_iopadmap_cc_313_execute_26881_3_) );
  OR2X2 OR2X2_5476 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n102_1), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n101_1), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n103) );
  OR2X2 OR2X2_5477 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n104), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n105), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n106_1) );
  OR2X2 OR2X2_5478 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n106_1), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n103), .Y(_auto_iopadmap_cc_313_execute_26881_4_) );
  OR2X2 OR2X2_5479 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n109), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n108), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n110_1) );
  OR2X2 OR2X2_548 ( .A(AES_CORE_DATAPATH__abc_16259_n3622_1), .B(AES_CORE_DATAPATH__abc_16259_n2864_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n3623) );
  OR2X2 OR2X2_5480 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n111), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n112), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n113) );
  OR2X2 OR2X2_5481 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n113), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n110_1), .Y(_auto_iopadmap_cc_313_execute_26881_5_) );
  OR2X2 OR2X2_5482 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n116), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n115), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n117) );
  OR2X2 OR2X2_5483 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n118_1), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n119), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n120) );
  OR2X2 OR2X2_5484 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n120), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n117), .Y(_auto_iopadmap_cc_313_execute_26881_6_) );
  OR2X2 OR2X2_5485 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n123), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n122_1), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n124) );
  OR2X2 OR2X2_5486 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n125), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n126_1), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n127) );
  OR2X2 OR2X2_5487 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n127), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n124), .Y(_auto_iopadmap_cc_313_execute_26881_7_) );
  OR2X2 OR2X2_5488 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n130_1), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n129), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n131) );
  OR2X2 OR2X2_5489 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n132), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n133), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n134_1) );
  OR2X2 OR2X2_549 ( .A(AES_CORE_DATAPATH__abc_16259_n3623), .B(AES_CORE_DATAPATH__abc_16259_n3621), .Y(AES_CORE_DATAPATH__abc_16259_n3624) );
  OR2X2 OR2X2_5490 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n134_1), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n131), .Y(_auto_iopadmap_cc_313_execute_26881_8_) );
  OR2X2 OR2X2_5491 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n137), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n136), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n138_1) );
  OR2X2 OR2X2_5492 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n139), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n140), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n141) );
  OR2X2 OR2X2_5493 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n141), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n138_1), .Y(_auto_iopadmap_cc_313_execute_26881_9_) );
  OR2X2 OR2X2_5494 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n144), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n143), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n145) );
  OR2X2 OR2X2_5495 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n146_1), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n147), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n148) );
  OR2X2 OR2X2_5496 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n148), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n145), .Y(_auto_iopadmap_cc_313_execute_26881_10_) );
  OR2X2 OR2X2_5497 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n151), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n150_1), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n152) );
  OR2X2 OR2X2_5498 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n153), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n154_1), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n155) );
  OR2X2 OR2X2_5499 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n155), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n152), .Y(_auto_iopadmap_cc_313_execute_26881_11_) );
  OR2X2 OR2X2_55 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n219), .B(AES_CORE_CONTROL_UNIT__abc_15841_n188), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n220) );
  OR2X2 OR2X2_550 ( .A(AES_CORE_DATAPATH__abc_16259_n3626), .B(AES_CORE_DATAPATH__abc_16259_n3625), .Y(AES_CORE_DATAPATH__abc_16259_n3627) );
  OR2X2 OR2X2_5500 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n158_1), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n157), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n159) );
  OR2X2 OR2X2_5501 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n160), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n161), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n162_1) );
  OR2X2 OR2X2_5502 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n162_1), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n159), .Y(_auto_iopadmap_cc_313_execute_26881_12_) );
  OR2X2 OR2X2_5503 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n165), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n164), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n166_1) );
  OR2X2 OR2X2_5504 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n167), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n168), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n169) );
  OR2X2 OR2X2_5505 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n169), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n166_1), .Y(_auto_iopadmap_cc_313_execute_26881_13_) );
  OR2X2 OR2X2_5506 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n172), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n171), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n173) );
  OR2X2 OR2X2_5507 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n174), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n175), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n176) );
  OR2X2 OR2X2_5508 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n176), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n173), .Y(_auto_iopadmap_cc_313_execute_26881_14_) );
  OR2X2 OR2X2_5509 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n179), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n178), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n180) );
  OR2X2 OR2X2_551 ( .A(AES_CORE_DATAPATH__abc_16259_n3627), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n3628) );
  OR2X2 OR2X2_5510 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n181), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n182), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n183) );
  OR2X2 OR2X2_5511 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n183), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n180), .Y(_auto_iopadmap_cc_313_execute_26881_15_) );
  OR2X2 OR2X2_5512 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n186), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n185), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n187) );
  OR2X2 OR2X2_5513 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n188), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n189), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n190) );
  OR2X2 OR2X2_5514 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n190), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n187), .Y(_auto_iopadmap_cc_313_execute_26881_16_) );
  OR2X2 OR2X2_5515 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n193), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n192), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n194) );
  OR2X2 OR2X2_5516 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n195), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n196), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n197) );
  OR2X2 OR2X2_5517 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n197), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n194), .Y(_auto_iopadmap_cc_313_execute_26881_17_) );
  OR2X2 OR2X2_5518 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n200), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n199), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n201) );
  OR2X2 OR2X2_5519 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n202), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n203), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n204) );
  OR2X2 OR2X2_552 ( .A(AES_CORE_DATAPATH__abc_16259_n3630), .B(AES_CORE_DATAPATH__abc_16259_n3631), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_19_) );
  OR2X2 OR2X2_5520 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n204), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n201), .Y(_auto_iopadmap_cc_313_execute_26881_18_) );
  OR2X2 OR2X2_5521 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n207), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n206), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n208) );
  OR2X2 OR2X2_5522 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n209), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n210), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n211) );
  OR2X2 OR2X2_5523 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n211), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n208), .Y(_auto_iopadmap_cc_313_execute_26881_19_) );
  OR2X2 OR2X2_5524 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n214), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n213), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n215) );
  OR2X2 OR2X2_5525 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n216), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n217), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n218) );
  OR2X2 OR2X2_5526 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n218), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n215), .Y(_auto_iopadmap_cc_313_execute_26881_20_) );
  OR2X2 OR2X2_5527 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n221), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n220), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n222) );
  OR2X2 OR2X2_5528 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n223), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n224), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n225) );
  OR2X2 OR2X2_5529 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n225), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n222), .Y(_auto_iopadmap_cc_313_execute_26881_21_) );
  OR2X2 OR2X2_553 ( .A(AES_CORE_DATAPATH__abc_16259_n2774_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n3633), .Y(AES_CORE_DATAPATH__abc_16259_n3634_1) );
  OR2X2 OR2X2_5530 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n228), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n227), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n229) );
  OR2X2 OR2X2_5531 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n230), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n231), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n232) );
  OR2X2 OR2X2_5532 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n232), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n229), .Y(_auto_iopadmap_cc_313_execute_26881_22_) );
  OR2X2 OR2X2_5533 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n235), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n234), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n236) );
  OR2X2 OR2X2_5534 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n237), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n238), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n239) );
  OR2X2 OR2X2_5535 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n239), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n236), .Y(_auto_iopadmap_cc_313_execute_26881_23_) );
  OR2X2 OR2X2_5536 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n242), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n241), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n243) );
  OR2X2 OR2X2_5537 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n244), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n245), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n246) );
  OR2X2 OR2X2_5538 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n246), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n243), .Y(_auto_iopadmap_cc_313_execute_26881_24_) );
  OR2X2 OR2X2_5539 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n249), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n248), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n250) );
  OR2X2 OR2X2_554 ( .A(AES_CORE_DATAPATH__abc_16259_n2778_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n3635), .Y(AES_CORE_DATAPATH__abc_16259_n3636_1) );
  OR2X2 OR2X2_5540 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n251), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n252), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n253) );
  OR2X2 OR2X2_5541 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n253), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n250), .Y(_auto_iopadmap_cc_313_execute_26881_25_) );
  OR2X2 OR2X2_5542 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n256), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n255), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n257) );
  OR2X2 OR2X2_5543 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n258), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n259), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n260) );
  OR2X2 OR2X2_5544 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n260), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n257), .Y(_auto_iopadmap_cc_313_execute_26881_26_) );
  OR2X2 OR2X2_5545 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n263), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n262), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n264) );
  OR2X2 OR2X2_5546 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n265), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n266), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n267) );
  OR2X2 OR2X2_5547 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n267), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n264), .Y(_auto_iopadmap_cc_313_execute_26881_27_) );
  OR2X2 OR2X2_5548 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n270), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n269), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n271) );
  OR2X2 OR2X2_5549 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n272), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n273), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n274) );
  OR2X2 OR2X2_555 ( .A(AES_CORE_DATAPATH__abc_16259_n3639), .B(AES_CORE_DATAPATH__abc_16259_n3640), .Y(AES_CORE_DATAPATH__abc_16259_n3641_1) );
  OR2X2 OR2X2_5550 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n274), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n271), .Y(_auto_iopadmap_cc_313_execute_26881_28_) );
  OR2X2 OR2X2_5551 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n277), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n276), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n278) );
  OR2X2 OR2X2_5552 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n279), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n280), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n281) );
  OR2X2 OR2X2_5553 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n281), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n278), .Y(_auto_iopadmap_cc_313_execute_26881_29_) );
  OR2X2 OR2X2_5554 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n284), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n283), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n285) );
  OR2X2 OR2X2_5555 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n286), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n287), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n288) );
  OR2X2 OR2X2_5556 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n288), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n285), .Y(_auto_iopadmap_cc_313_execute_26881_30_) );
  OR2X2 OR2X2_5557 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n291), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n290), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n292) );
  OR2X2 OR2X2_5558 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n293), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n294), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n295) );
  OR2X2 OR2X2_5559 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n295), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_16028_n292), .Y(_auto_iopadmap_cc_313_execute_26881_31_) );
  OR2X2 OR2X2_556 ( .A(AES_CORE_DATAPATH__abc_16259_n3641_1), .B(AES_CORE_DATAPATH__abc_16259_n3638), .Y(AES_CORE_DATAPATH__abc_16259_n3642_1) );
  OR2X2 OR2X2_557 ( .A(AES_CORE_DATAPATH__abc_16259_n3646), .B(AES_CORE_DATAPATH__abc_16259_n2826_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n3647_1) );
  OR2X2 OR2X2_558 ( .A(AES_CORE_DATAPATH__abc_16259_n3648), .B(AES_CORE_DATAPATH__abc_16259_n3649_1), .Y(AES_CORE_DATAPATH__abc_16259_n3650) );
  OR2X2 OR2X2_559 ( .A(AES_CORE_DATAPATH__abc_16259_n3650), .B(AES_CORE_DATAPATH__abc_16259_n3647_1), .Y(AES_CORE_DATAPATH__abc_16259_n3651_1) );
  OR2X2 OR2X2_56 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n118), .B(AES_CORE_CONTROL_UNIT__abc_15841_n220), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n221) );
  OR2X2 OR2X2_560 ( .A(AES_CORE_DATAPATH__abc_16259_n2841_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__20_), .Y(AES_CORE_DATAPATH__abc_16259_n3652) );
  OR2X2 OR2X2_561 ( .A(AES_CORE_DATAPATH__abc_16259_n3644), .B(AES_CORE_DATAPATH__abc_16259_n2853_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n3654) );
  OR2X2 OR2X2_562 ( .A(AES_CORE_DATAPATH__abc_16259_n3655), .B(AES_CORE_DATAPATH__abc_16259_n3656), .Y(AES_CORE_DATAPATH__abc_16259_n3657) );
  OR2X2 OR2X2_563 ( .A(_auto_iopadmap_cc_313_execute_26949_20_), .B(AES_CORE_DATAPATH__abc_16259_n3659), .Y(AES_CORE_DATAPATH__abc_16259_n3660) );
  OR2X2 OR2X2_564 ( .A(AES_CORE_DATAPATH__abc_16259_n3662), .B(AES_CORE_DATAPATH__abc_16259_n2864_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n3663_1) );
  OR2X2 OR2X2_565 ( .A(AES_CORE_DATAPATH__abc_16259_n3663_1), .B(AES_CORE_DATAPATH__abc_16259_n3661), .Y(AES_CORE_DATAPATH__abc_16259_n3664) );
  OR2X2 OR2X2_566 ( .A(AES_CORE_DATAPATH__abc_16259_n3666), .B(AES_CORE_DATAPATH__abc_16259_n3665_1), .Y(AES_CORE_DATAPATH__abc_16259_n3667) );
  OR2X2 OR2X2_567 ( .A(AES_CORE_DATAPATH__abc_16259_n3667), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n3668) );
  OR2X2 OR2X2_568 ( .A(AES_CORE_DATAPATH__abc_16259_n3670_1), .B(AES_CORE_DATAPATH__abc_16259_n3671_1), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_20_) );
  OR2X2 OR2X2_569 ( .A(AES_CORE_DATAPATH__abc_16259_n2774_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n3673_1), .Y(AES_CORE_DATAPATH__abc_16259_n3674) );
  OR2X2 OR2X2_57 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n218), .B(AES_CORE_CONTROL_UNIT__abc_15841_n221), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n222) );
  OR2X2 OR2X2_570 ( .A(AES_CORE_DATAPATH__abc_16259_n2778_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n3675), .Y(AES_CORE_DATAPATH__abc_16259_n3676) );
  OR2X2 OR2X2_571 ( .A(AES_CORE_DATAPATH__abc_16259_n3679_1), .B(AES_CORE_DATAPATH__abc_16259_n3680), .Y(AES_CORE_DATAPATH__abc_16259_n3681_1) );
  OR2X2 OR2X2_572 ( .A(AES_CORE_DATAPATH__abc_16259_n3681_1), .B(AES_CORE_DATAPATH__abc_16259_n3678_1), .Y(AES_CORE_DATAPATH__abc_16259_n3682) );
  OR2X2 OR2X2_573 ( .A(AES_CORE_DATAPATH__abc_16259_n3686_1), .B(AES_CORE_DATAPATH__abc_16259_n2826_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n3687_1) );
  OR2X2 OR2X2_574 ( .A(AES_CORE_DATAPATH__abc_16259_n3688), .B(AES_CORE_DATAPATH__abc_16259_n3689_1), .Y(AES_CORE_DATAPATH__abc_16259_n3690) );
  OR2X2 OR2X2_575 ( .A(AES_CORE_DATAPATH__abc_16259_n3690), .B(AES_CORE_DATAPATH__abc_16259_n3687_1), .Y(AES_CORE_DATAPATH__abc_16259_n3691) );
  OR2X2 OR2X2_576 ( .A(AES_CORE_DATAPATH__abc_16259_n2841_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__21_), .Y(AES_CORE_DATAPATH__abc_16259_n3692) );
  OR2X2 OR2X2_577 ( .A(AES_CORE_DATAPATH__abc_16259_n3684), .B(AES_CORE_DATAPATH__abc_16259_n2853_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n3694_1) );
  OR2X2 OR2X2_578 ( .A(AES_CORE_DATAPATH__abc_16259_n3695_1), .B(AES_CORE_DATAPATH__abc_16259_n3696), .Y(AES_CORE_DATAPATH__abc_16259_n3697_1) );
  OR2X2 OR2X2_579 ( .A(_auto_iopadmap_cc_313_execute_26949_21_), .B(AES_CORE_DATAPATH__abc_16259_n3699), .Y(AES_CORE_DATAPATH__abc_16259_n3700) );
  OR2X2 OR2X2_58 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n223), .B(AES_CORE_CONTROL_UNIT__abc_15841_n212_1), .Y(AES_CORE_CONTROL_UNIT_col_sel_0_) );
  OR2X2 OR2X2_580 ( .A(AES_CORE_DATAPATH__abc_16259_n3702_1), .B(AES_CORE_DATAPATH__abc_16259_n2864_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n3703_1) );
  OR2X2 OR2X2_581 ( .A(AES_CORE_DATAPATH__abc_16259_n3703_1), .B(AES_CORE_DATAPATH__abc_16259_n3701), .Y(AES_CORE_DATAPATH__abc_16259_n3704) );
  OR2X2 OR2X2_582 ( .A(AES_CORE_DATAPATH__abc_16259_n3706), .B(AES_CORE_DATAPATH__abc_16259_n3705_1), .Y(AES_CORE_DATAPATH__abc_16259_n3707) );
  OR2X2 OR2X2_583 ( .A(AES_CORE_DATAPATH__abc_16259_n3707), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n3708) );
  OR2X2 OR2X2_584 ( .A(AES_CORE_DATAPATH__abc_16259_n3710_1), .B(AES_CORE_DATAPATH__abc_16259_n3711_1), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_21_) );
  OR2X2 OR2X2_585 ( .A(AES_CORE_DATAPATH__abc_16259_n2774_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n3713_1), .Y(AES_CORE_DATAPATH__abc_16259_n3714) );
  OR2X2 OR2X2_586 ( .A(AES_CORE_DATAPATH__abc_16259_n2778_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n3715), .Y(AES_CORE_DATAPATH__abc_16259_n3716) );
  OR2X2 OR2X2_587 ( .A(AES_CORE_DATAPATH__abc_16259_n3719_1), .B(AES_CORE_DATAPATH__abc_16259_n3720), .Y(AES_CORE_DATAPATH__abc_16259_n3721_1) );
  OR2X2 OR2X2_588 ( .A(AES_CORE_DATAPATH__abc_16259_n3721_1), .B(AES_CORE_DATAPATH__abc_16259_n3718_1), .Y(AES_CORE_DATAPATH__abc_16259_n3722) );
  OR2X2 OR2X2_589 ( .A(AES_CORE_DATAPATH__abc_16259_n3726_1), .B(AES_CORE_DATAPATH__abc_16259_n2826_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n3727_1) );
  OR2X2 OR2X2_59 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n225), .B(AES_CORE_CONTROL_UNIT__abc_15841_n232), .Y(AES_CORE_CONTROL_UNIT_col_sel_1_) );
  OR2X2 OR2X2_590 ( .A(AES_CORE_DATAPATH__abc_16259_n3728), .B(AES_CORE_DATAPATH__abc_16259_n3729_1), .Y(AES_CORE_DATAPATH__abc_16259_n3730) );
  OR2X2 OR2X2_591 ( .A(AES_CORE_DATAPATH__abc_16259_n3730), .B(AES_CORE_DATAPATH__abc_16259_n3727_1), .Y(AES_CORE_DATAPATH__abc_16259_n3731) );
  OR2X2 OR2X2_592 ( .A(AES_CORE_DATAPATH__abc_16259_n2841_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__22_), .Y(AES_CORE_DATAPATH__abc_16259_n3732) );
  OR2X2 OR2X2_593 ( .A(AES_CORE_DATAPATH__abc_16259_n3724), .B(AES_CORE_DATAPATH__abc_16259_n2853_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n3734_1) );
  OR2X2 OR2X2_594 ( .A(AES_CORE_DATAPATH__abc_16259_n3735_1), .B(AES_CORE_DATAPATH__abc_16259_n3736), .Y(AES_CORE_DATAPATH__abc_16259_n3737_1) );
  OR2X2 OR2X2_595 ( .A(_auto_iopadmap_cc_313_execute_26949_22_), .B(AES_CORE_DATAPATH__abc_16259_n3739), .Y(AES_CORE_DATAPATH__abc_16259_n3740) );
  OR2X2 OR2X2_596 ( .A(AES_CORE_DATAPATH__abc_16259_n3742_1), .B(AES_CORE_DATAPATH__abc_16259_n2864_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n3743_1) );
  OR2X2 OR2X2_597 ( .A(AES_CORE_DATAPATH__abc_16259_n3743_1), .B(AES_CORE_DATAPATH__abc_16259_n3741), .Y(AES_CORE_DATAPATH__abc_16259_n3744) );
  OR2X2 OR2X2_598 ( .A(AES_CORE_DATAPATH__abc_16259_n3746), .B(AES_CORE_DATAPATH__abc_16259_n3745_1), .Y(AES_CORE_DATAPATH__abc_16259_n3747) );
  OR2X2 OR2X2_599 ( .A(AES_CORE_DATAPATH__abc_16259_n3747), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n3748) );
  OR2X2 OR2X2_6 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n88), .B(\aes_mode[0] ), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n89_1) );
  OR2X2 OR2X2_60 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n198), .B(AES_CORE_CONTROL_UNIT__abc_15841_n206_1), .Y(AES_CORE_CONTROL_UNIT_key_out_sel_0_) );
  OR2X2 OR2X2_600 ( .A(AES_CORE_DATAPATH__abc_16259_n3750_1), .B(AES_CORE_DATAPATH__abc_16259_n3751_1), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_22_) );
  OR2X2 OR2X2_601 ( .A(AES_CORE_DATAPATH__abc_16259_n2774_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n3753_1), .Y(AES_CORE_DATAPATH__abc_16259_n3754) );
  OR2X2 OR2X2_602 ( .A(AES_CORE_DATAPATH__abc_16259_n2778_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n3755), .Y(AES_CORE_DATAPATH__abc_16259_n3756) );
  OR2X2 OR2X2_603 ( .A(AES_CORE_DATAPATH__abc_16259_n3759_1), .B(AES_CORE_DATAPATH__abc_16259_n3760), .Y(AES_CORE_DATAPATH__abc_16259_n3761_1) );
  OR2X2 OR2X2_604 ( .A(AES_CORE_DATAPATH__abc_16259_n3761_1), .B(AES_CORE_DATAPATH__abc_16259_n3758_1), .Y(AES_CORE_DATAPATH__abc_16259_n3762) );
  OR2X2 OR2X2_605 ( .A(AES_CORE_DATAPATH__abc_16259_n3766_1), .B(AES_CORE_DATAPATH__abc_16259_n2826_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n3767_1) );
  OR2X2 OR2X2_606 ( .A(AES_CORE_DATAPATH__abc_16259_n3768), .B(AES_CORE_DATAPATH__abc_16259_n3769_1), .Y(AES_CORE_DATAPATH__abc_16259_n3770) );
  OR2X2 OR2X2_607 ( .A(AES_CORE_DATAPATH__abc_16259_n3770), .B(AES_CORE_DATAPATH__abc_16259_n3767_1), .Y(AES_CORE_DATAPATH__abc_16259_n3771) );
  OR2X2 OR2X2_608 ( .A(AES_CORE_DATAPATH__abc_16259_n2841_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__23_), .Y(AES_CORE_DATAPATH__abc_16259_n3772) );
  OR2X2 OR2X2_609 ( .A(AES_CORE_DATAPATH__abc_16259_n3764), .B(AES_CORE_DATAPATH__abc_16259_n2853_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n3774_1) );
  OR2X2 OR2X2_61 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n203_1), .B(AES_CORE_CONTROL_UNIT__abc_15841_n206_1), .Y(AES_CORE_CONTROL_UNIT_key_out_sel_1_) );
  OR2X2 OR2X2_610 ( .A(AES_CORE_DATAPATH__abc_16259_n3775_1), .B(AES_CORE_DATAPATH__abc_16259_n3776), .Y(AES_CORE_DATAPATH__abc_16259_n3777_1) );
  OR2X2 OR2X2_611 ( .A(_auto_iopadmap_cc_313_execute_26949_23_), .B(AES_CORE_DATAPATH__abc_16259_n3779), .Y(AES_CORE_DATAPATH__abc_16259_n3780) );
  OR2X2 OR2X2_612 ( .A(AES_CORE_DATAPATH__abc_16259_n3782_1), .B(AES_CORE_DATAPATH__abc_16259_n2864_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n3783_1) );
  OR2X2 OR2X2_613 ( .A(AES_CORE_DATAPATH__abc_16259_n3783_1), .B(AES_CORE_DATAPATH__abc_16259_n3781), .Y(AES_CORE_DATAPATH__abc_16259_n3784) );
  OR2X2 OR2X2_614 ( .A(AES_CORE_DATAPATH__abc_16259_n3786), .B(AES_CORE_DATAPATH__abc_16259_n3785_1), .Y(AES_CORE_DATAPATH__abc_16259_n3787) );
  OR2X2 OR2X2_615 ( .A(AES_CORE_DATAPATH__abc_16259_n3787), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n3788) );
  OR2X2 OR2X2_616 ( .A(AES_CORE_DATAPATH__abc_16259_n3790_1), .B(AES_CORE_DATAPATH__abc_16259_n3791_1), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_23_) );
  OR2X2 OR2X2_617 ( .A(AES_CORE_DATAPATH__abc_16259_n2774_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n3793_1), .Y(AES_CORE_DATAPATH__abc_16259_n3794) );
  OR2X2 OR2X2_618 ( .A(AES_CORE_DATAPATH__abc_16259_n2778_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n3795), .Y(AES_CORE_DATAPATH__abc_16259_n3796) );
  OR2X2 OR2X2_619 ( .A(AES_CORE_DATAPATH__abc_16259_n3799_1), .B(AES_CORE_DATAPATH__abc_16259_n3800), .Y(AES_CORE_DATAPATH__abc_16259_n3801_1) );
  OR2X2 OR2X2_62 ( .A(AES_CORE_CONTROL_UNIT_state_3_), .B(AES_CORE_CONTROL_UNIT_key_gen), .Y(AES_CORE_CONTROL_UNIT_key_en_0_) );
  OR2X2 OR2X2_620 ( .A(AES_CORE_DATAPATH__abc_16259_n3801_1), .B(AES_CORE_DATAPATH__abc_16259_n3798_1), .Y(AES_CORE_DATAPATH__abc_16259_n3802) );
  OR2X2 OR2X2_621 ( .A(AES_CORE_DATAPATH__abc_16259_n3806_1), .B(AES_CORE_DATAPATH__abc_16259_n2826_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n3807_1) );
  OR2X2 OR2X2_622 ( .A(AES_CORE_DATAPATH__abc_16259_n3808), .B(AES_CORE_DATAPATH__abc_16259_n3809_1), .Y(AES_CORE_DATAPATH__abc_16259_n3810) );
  OR2X2 OR2X2_623 ( .A(AES_CORE_DATAPATH__abc_16259_n3810), .B(AES_CORE_DATAPATH__abc_16259_n3807_1), .Y(AES_CORE_DATAPATH__abc_16259_n3811) );
  OR2X2 OR2X2_624 ( .A(AES_CORE_DATAPATH__abc_16259_n2841_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__24_), .Y(AES_CORE_DATAPATH__abc_16259_n3812) );
  OR2X2 OR2X2_625 ( .A(AES_CORE_DATAPATH__abc_16259_n3804), .B(AES_CORE_DATAPATH__abc_16259_n2853_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n3814_1) );
  OR2X2 OR2X2_626 ( .A(AES_CORE_DATAPATH__abc_16259_n3815_1), .B(AES_CORE_DATAPATH__abc_16259_n3816), .Y(AES_CORE_DATAPATH__abc_16259_n3817_1) );
  OR2X2 OR2X2_627 ( .A(_auto_iopadmap_cc_313_execute_26949_24_), .B(AES_CORE_DATAPATH__abc_16259_n3819), .Y(AES_CORE_DATAPATH__abc_16259_n3820) );
  OR2X2 OR2X2_628 ( .A(AES_CORE_DATAPATH__abc_16259_n3822_1), .B(AES_CORE_DATAPATH__abc_16259_n2864_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n3823_1) );
  OR2X2 OR2X2_629 ( .A(AES_CORE_DATAPATH__abc_16259_n3823_1), .B(AES_CORE_DATAPATH__abc_16259_n3821), .Y(AES_CORE_DATAPATH__abc_16259_n3824) );
  OR2X2 OR2X2_63 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n75), .B(AES_CORE_CONTROL_UNIT_key_en_0_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n238) );
  OR2X2 OR2X2_630 ( .A(AES_CORE_DATAPATH__abc_16259_n3826), .B(AES_CORE_DATAPATH__abc_16259_n3825_1), .Y(AES_CORE_DATAPATH__abc_16259_n3827) );
  OR2X2 OR2X2_631 ( .A(AES_CORE_DATAPATH__abc_16259_n3827), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf6), .Y(AES_CORE_DATAPATH__abc_16259_n3828) );
  OR2X2 OR2X2_632 ( .A(AES_CORE_DATAPATH__abc_16259_n3830_1), .B(AES_CORE_DATAPATH__abc_16259_n3831_1), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_24_) );
  OR2X2 OR2X2_633 ( .A(AES_CORE_DATAPATH__abc_16259_n2774_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n3833_1), .Y(AES_CORE_DATAPATH__abc_16259_n3834) );
  OR2X2 OR2X2_634 ( .A(AES_CORE_DATAPATH__abc_16259_n2778_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n3835), .Y(AES_CORE_DATAPATH__abc_16259_n3836) );
  OR2X2 OR2X2_635 ( .A(AES_CORE_DATAPATH__abc_16259_n3839_1), .B(AES_CORE_DATAPATH__abc_16259_n3840), .Y(AES_CORE_DATAPATH__abc_16259_n3841_1) );
  OR2X2 OR2X2_636 ( .A(AES_CORE_DATAPATH__abc_16259_n3841_1), .B(AES_CORE_DATAPATH__abc_16259_n3838_1), .Y(AES_CORE_DATAPATH__abc_16259_n3842) );
  OR2X2 OR2X2_637 ( .A(AES_CORE_DATAPATH__abc_16259_n3846_1), .B(AES_CORE_DATAPATH__abc_16259_n2826_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n3847_1) );
  OR2X2 OR2X2_638 ( .A(AES_CORE_DATAPATH__abc_16259_n3848), .B(AES_CORE_DATAPATH__abc_16259_n3849_1), .Y(AES_CORE_DATAPATH__abc_16259_n3850) );
  OR2X2 OR2X2_639 ( .A(AES_CORE_DATAPATH__abc_16259_n3850), .B(AES_CORE_DATAPATH__abc_16259_n3847_1), .Y(AES_CORE_DATAPATH__abc_16259_n3851) );
  OR2X2 OR2X2_64 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n190), .B(AES_CORE_CONTROL_UNIT__abc_15841_n238), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n239) );
  OR2X2 OR2X2_640 ( .A(AES_CORE_DATAPATH__abc_16259_n2841_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__25_), .Y(AES_CORE_DATAPATH__abc_16259_n3852) );
  OR2X2 OR2X2_641 ( .A(AES_CORE_DATAPATH__abc_16259_n3844), .B(AES_CORE_DATAPATH__abc_16259_n2853_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n3854_1) );
  OR2X2 OR2X2_642 ( .A(AES_CORE_DATAPATH__abc_16259_n3855_1), .B(AES_CORE_DATAPATH__abc_16259_n3856), .Y(AES_CORE_DATAPATH__abc_16259_n3857_1) );
  OR2X2 OR2X2_643 ( .A(_auto_iopadmap_cc_313_execute_26949_25_), .B(AES_CORE_DATAPATH__abc_16259_n3859), .Y(AES_CORE_DATAPATH__abc_16259_n3860) );
  OR2X2 OR2X2_644 ( .A(AES_CORE_DATAPATH__abc_16259_n3862_1), .B(AES_CORE_DATAPATH__abc_16259_n2864_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n3863_1) );
  OR2X2 OR2X2_645 ( .A(AES_CORE_DATAPATH__abc_16259_n3863_1), .B(AES_CORE_DATAPATH__abc_16259_n3861), .Y(AES_CORE_DATAPATH__abc_16259_n3864) );
  OR2X2 OR2X2_646 ( .A(AES_CORE_DATAPATH__abc_16259_n3866), .B(AES_CORE_DATAPATH__abc_16259_n3865_1), .Y(AES_CORE_DATAPATH__abc_16259_n3867) );
  OR2X2 OR2X2_647 ( .A(AES_CORE_DATAPATH__abc_16259_n3867), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n3868) );
  OR2X2 OR2X2_648 ( .A(AES_CORE_DATAPATH__abc_16259_n3870_1), .B(AES_CORE_DATAPATH__abc_16259_n3871_1), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_25_) );
  OR2X2 OR2X2_649 ( .A(AES_CORE_DATAPATH__abc_16259_n2774_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n3873_1), .Y(AES_CORE_DATAPATH__abc_16259_n3874) );
  OR2X2 OR2X2_65 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n236), .B(AES_CORE_CONTROL_UNIT__abc_15841_n239), .Y(AES_CORE_CONTROL_UNIT_key_sel) );
  OR2X2 OR2X2_650 ( .A(AES_CORE_DATAPATH__abc_16259_n2778_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n3875), .Y(AES_CORE_DATAPATH__abc_16259_n3876) );
  OR2X2 OR2X2_651 ( .A(AES_CORE_DATAPATH__abc_16259_n3879_1), .B(AES_CORE_DATAPATH__abc_16259_n3880), .Y(AES_CORE_DATAPATH__abc_16259_n3881_1) );
  OR2X2 OR2X2_652 ( .A(AES_CORE_DATAPATH__abc_16259_n3881_1), .B(AES_CORE_DATAPATH__abc_16259_n3878_1), .Y(AES_CORE_DATAPATH__abc_16259_n3882) );
  OR2X2 OR2X2_653 ( .A(AES_CORE_DATAPATH__abc_16259_n3886_1), .B(AES_CORE_DATAPATH__abc_16259_n2826_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n3887_1) );
  OR2X2 OR2X2_654 ( .A(AES_CORE_DATAPATH__abc_16259_n3888), .B(AES_CORE_DATAPATH__abc_16259_n3889_1), .Y(AES_CORE_DATAPATH__abc_16259_n3890) );
  OR2X2 OR2X2_655 ( .A(AES_CORE_DATAPATH__abc_16259_n3890), .B(AES_CORE_DATAPATH__abc_16259_n3887_1), .Y(AES_CORE_DATAPATH__abc_16259_n3891) );
  OR2X2 OR2X2_656 ( .A(AES_CORE_DATAPATH__abc_16259_n2841_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__26_), .Y(AES_CORE_DATAPATH__abc_16259_n3892) );
  OR2X2 OR2X2_657 ( .A(AES_CORE_DATAPATH__abc_16259_n3884), .B(AES_CORE_DATAPATH__abc_16259_n2853_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n3894_1) );
  OR2X2 OR2X2_658 ( .A(AES_CORE_DATAPATH__abc_16259_n3895_1), .B(AES_CORE_DATAPATH__abc_16259_n3896), .Y(AES_CORE_DATAPATH__abc_16259_n3897_1) );
  OR2X2 OR2X2_659 ( .A(_auto_iopadmap_cc_313_execute_26949_26_), .B(AES_CORE_DATAPATH__abc_16259_n3899), .Y(AES_CORE_DATAPATH__abc_16259_n3900) );
  OR2X2 OR2X2_66 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n158), .B(AES_CORE_CONTROL_UNIT_state_3_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n242) );
  OR2X2 OR2X2_660 ( .A(AES_CORE_DATAPATH__abc_16259_n3902_1), .B(AES_CORE_DATAPATH__abc_16259_n2864_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n3903_1) );
  OR2X2 OR2X2_661 ( .A(AES_CORE_DATAPATH__abc_16259_n3903_1), .B(AES_CORE_DATAPATH__abc_16259_n3901), .Y(AES_CORE_DATAPATH__abc_16259_n3904) );
  OR2X2 OR2X2_662 ( .A(AES_CORE_DATAPATH__abc_16259_n3906), .B(AES_CORE_DATAPATH__abc_16259_n3905_1), .Y(AES_CORE_DATAPATH__abc_16259_n3907) );
  OR2X2 OR2X2_663 ( .A(AES_CORE_DATAPATH__abc_16259_n3907), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n3908) );
  OR2X2 OR2X2_664 ( .A(AES_CORE_DATAPATH__abc_16259_n3910_1), .B(AES_CORE_DATAPATH__abc_16259_n3911_1), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_26_) );
  OR2X2 OR2X2_665 ( .A(AES_CORE_DATAPATH__abc_16259_n2774_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n3913_1), .Y(AES_CORE_DATAPATH__abc_16259_n3914) );
  OR2X2 OR2X2_666 ( .A(AES_CORE_DATAPATH__abc_16259_n2778_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n3915), .Y(AES_CORE_DATAPATH__abc_16259_n3916) );
  OR2X2 OR2X2_667 ( .A(AES_CORE_DATAPATH__abc_16259_n3919_1), .B(AES_CORE_DATAPATH__abc_16259_n3920), .Y(AES_CORE_DATAPATH__abc_16259_n3921_1) );
  OR2X2 OR2X2_668 ( .A(AES_CORE_DATAPATH__abc_16259_n3921_1), .B(AES_CORE_DATAPATH__abc_16259_n3918_1), .Y(AES_CORE_DATAPATH__abc_16259_n3922) );
  OR2X2 OR2X2_669 ( .A(AES_CORE_DATAPATH__abc_16259_n3926_1), .B(AES_CORE_DATAPATH__abc_16259_n2826_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n3927_1) );
  OR2X2 OR2X2_67 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n242), .B(AES_CORE_CONTROL_UNIT__abc_15841_n241), .Y(AES_CORE_CONTROL_UNIT_key_en_1_) );
  OR2X2 OR2X2_670 ( .A(AES_CORE_DATAPATH__abc_16259_n3928), .B(AES_CORE_DATAPATH__abc_16259_n3929_1), .Y(AES_CORE_DATAPATH__abc_16259_n3930) );
  OR2X2 OR2X2_671 ( .A(AES_CORE_DATAPATH__abc_16259_n3930), .B(AES_CORE_DATAPATH__abc_16259_n3927_1), .Y(AES_CORE_DATAPATH__abc_16259_n3931) );
  OR2X2 OR2X2_672 ( .A(AES_CORE_DATAPATH__abc_16259_n2841_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__27_), .Y(AES_CORE_DATAPATH__abc_16259_n3932) );
  OR2X2 OR2X2_673 ( .A(AES_CORE_DATAPATH__abc_16259_n3924), .B(AES_CORE_DATAPATH__abc_16259_n2853_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n3934_1) );
  OR2X2 OR2X2_674 ( .A(AES_CORE_DATAPATH__abc_16259_n3935_1), .B(AES_CORE_DATAPATH__abc_16259_n3936), .Y(AES_CORE_DATAPATH__abc_16259_n3937_1) );
  OR2X2 OR2X2_675 ( .A(_auto_iopadmap_cc_313_execute_26949_27_), .B(AES_CORE_DATAPATH__abc_16259_n3939), .Y(AES_CORE_DATAPATH__abc_16259_n3940) );
  OR2X2 OR2X2_676 ( .A(AES_CORE_DATAPATH__abc_16259_n3942_1), .B(AES_CORE_DATAPATH__abc_16259_n2864_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n3943_1) );
  OR2X2 OR2X2_677 ( .A(AES_CORE_DATAPATH__abc_16259_n3943_1), .B(AES_CORE_DATAPATH__abc_16259_n3941), .Y(AES_CORE_DATAPATH__abc_16259_n3944) );
  OR2X2 OR2X2_678 ( .A(AES_CORE_DATAPATH__abc_16259_n3946), .B(AES_CORE_DATAPATH__abc_16259_n3945_1), .Y(AES_CORE_DATAPATH__abc_16259_n3947) );
  OR2X2 OR2X2_679 ( .A(AES_CORE_DATAPATH__abc_16259_n3947), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n3948) );
  OR2X2 OR2X2_68 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n117_1), .B(AES_CORE_CONTROL_UNIT_state_11_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n245) );
  OR2X2 OR2X2_680 ( .A(AES_CORE_DATAPATH__abc_16259_n3950_1), .B(AES_CORE_DATAPATH__abc_16259_n3951_1), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_27_) );
  OR2X2 OR2X2_681 ( .A(AES_CORE_DATAPATH__abc_16259_n2774_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n3953_1), .Y(AES_CORE_DATAPATH__abc_16259_n3954) );
  OR2X2 OR2X2_682 ( .A(AES_CORE_DATAPATH__abc_16259_n2778_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n3955), .Y(AES_CORE_DATAPATH__abc_16259_n3956) );
  OR2X2 OR2X2_683 ( .A(AES_CORE_DATAPATH__abc_16259_n3959_1), .B(AES_CORE_DATAPATH__abc_16259_n3960), .Y(AES_CORE_DATAPATH__abc_16259_n3961_1) );
  OR2X2 OR2X2_684 ( .A(AES_CORE_DATAPATH__abc_16259_n3961_1), .B(AES_CORE_DATAPATH__abc_16259_n3958_1), .Y(AES_CORE_DATAPATH__abc_16259_n3962) );
  OR2X2 OR2X2_685 ( .A(AES_CORE_DATAPATH__abc_16259_n3966_1), .B(AES_CORE_DATAPATH__abc_16259_n2826_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n3967_1) );
  OR2X2 OR2X2_686 ( .A(AES_CORE_DATAPATH__abc_16259_n3968), .B(AES_CORE_DATAPATH__abc_16259_n3969_1), .Y(AES_CORE_DATAPATH__abc_16259_n3970) );
  OR2X2 OR2X2_687 ( .A(AES_CORE_DATAPATH__abc_16259_n3970), .B(AES_CORE_DATAPATH__abc_16259_n3967_1), .Y(AES_CORE_DATAPATH__abc_16259_n3971) );
  OR2X2 OR2X2_688 ( .A(AES_CORE_DATAPATH__abc_16259_n2841_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__28_), .Y(AES_CORE_DATAPATH__abc_16259_n3972) );
  OR2X2 OR2X2_689 ( .A(AES_CORE_DATAPATH__abc_16259_n3964), .B(AES_CORE_DATAPATH__abc_16259_n2853_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n3974_1) );
  OR2X2 OR2X2_69 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n245), .B(AES_CORE_CONTROL_UNIT__abc_15841_n244), .Y(AES_CORE_CONTROL_UNIT_key_en_2_) );
  OR2X2 OR2X2_690 ( .A(AES_CORE_DATAPATH__abc_16259_n3975_1), .B(AES_CORE_DATAPATH__abc_16259_n3976), .Y(AES_CORE_DATAPATH__abc_16259_n3977_1) );
  OR2X2 OR2X2_691 ( .A(_auto_iopadmap_cc_313_execute_26949_28_), .B(AES_CORE_DATAPATH__abc_16259_n3979), .Y(AES_CORE_DATAPATH__abc_16259_n3980) );
  OR2X2 OR2X2_692 ( .A(AES_CORE_DATAPATH__abc_16259_n3982_1), .B(AES_CORE_DATAPATH__abc_16259_n2864_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n3983_1) );
  OR2X2 OR2X2_693 ( .A(AES_CORE_DATAPATH__abc_16259_n3983_1), .B(AES_CORE_DATAPATH__abc_16259_n3981), .Y(AES_CORE_DATAPATH__abc_16259_n3984) );
  OR2X2 OR2X2_694 ( .A(AES_CORE_DATAPATH__abc_16259_n3986), .B(AES_CORE_DATAPATH__abc_16259_n3985_1), .Y(AES_CORE_DATAPATH__abc_16259_n3987) );
  OR2X2 OR2X2_695 ( .A(AES_CORE_DATAPATH__abc_16259_n3987), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n3988) );
  OR2X2 OR2X2_696 ( .A(AES_CORE_DATAPATH__abc_16259_n3990_1), .B(AES_CORE_DATAPATH__abc_16259_n3991_1), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_28_) );
  OR2X2 OR2X2_697 ( .A(AES_CORE_DATAPATH__abc_16259_n2774_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n3993_1), .Y(AES_CORE_DATAPATH__abc_16259_n3994) );
  OR2X2 OR2X2_698 ( .A(AES_CORE_DATAPATH__abc_16259_n2778_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n3995), .Y(AES_CORE_DATAPATH__abc_16259_n3996) );
  OR2X2 OR2X2_699 ( .A(AES_CORE_DATAPATH__abc_16259_n3999_1), .B(AES_CORE_DATAPATH__abc_16259_n4000), .Y(AES_CORE_DATAPATH__abc_16259_n4001_1) );
  OR2X2 OR2X2_7 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n94), .B(AES_CORE_CONTROL_UNIT__abc_15841_n100), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n101_1) );
  OR2X2 OR2X2_70 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n248), .B(AES_CORE_CONTROL_UNIT_state_7_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n249) );
  OR2X2 OR2X2_700 ( .A(AES_CORE_DATAPATH__abc_16259_n4001_1), .B(AES_CORE_DATAPATH__abc_16259_n3998_1), .Y(AES_CORE_DATAPATH__abc_16259_n4002) );
  OR2X2 OR2X2_701 ( .A(AES_CORE_DATAPATH__abc_16259_n4006_1), .B(AES_CORE_DATAPATH__abc_16259_n2826_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n4007_1) );
  OR2X2 OR2X2_702 ( .A(AES_CORE_DATAPATH__abc_16259_n4008), .B(AES_CORE_DATAPATH__abc_16259_n4009_1), .Y(AES_CORE_DATAPATH__abc_16259_n4010) );
  OR2X2 OR2X2_703 ( .A(AES_CORE_DATAPATH__abc_16259_n4010), .B(AES_CORE_DATAPATH__abc_16259_n4007_1), .Y(AES_CORE_DATAPATH__abc_16259_n4011) );
  OR2X2 OR2X2_704 ( .A(AES_CORE_DATAPATH__abc_16259_n2841_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__29_), .Y(AES_CORE_DATAPATH__abc_16259_n4012) );
  OR2X2 OR2X2_705 ( .A(AES_CORE_DATAPATH__abc_16259_n4004), .B(AES_CORE_DATAPATH__abc_16259_n2853_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n4014_1) );
  OR2X2 OR2X2_706 ( .A(AES_CORE_DATAPATH__abc_16259_n4015_1), .B(AES_CORE_DATAPATH__abc_16259_n4016), .Y(AES_CORE_DATAPATH__abc_16259_n4017_1) );
  OR2X2 OR2X2_707 ( .A(_auto_iopadmap_cc_313_execute_26949_29_), .B(AES_CORE_DATAPATH__abc_16259_n4019), .Y(AES_CORE_DATAPATH__abc_16259_n4020) );
  OR2X2 OR2X2_708 ( .A(AES_CORE_DATAPATH__abc_16259_n4022_1), .B(AES_CORE_DATAPATH__abc_16259_n2864_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n4023_1) );
  OR2X2 OR2X2_709 ( .A(AES_CORE_DATAPATH__abc_16259_n4023_1), .B(AES_CORE_DATAPATH__abc_16259_n4021), .Y(AES_CORE_DATAPATH__abc_16259_n4024) );
  OR2X2 OR2X2_71 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n249), .B(AES_CORE_CONTROL_UNIT__abc_15841_n247), .Y(AES_CORE_CONTROL_UNIT_key_en_3_) );
  OR2X2 OR2X2_710 ( .A(AES_CORE_DATAPATH__abc_16259_n4026), .B(AES_CORE_DATAPATH__abc_16259_n4025_1), .Y(AES_CORE_DATAPATH__abc_16259_n4027) );
  OR2X2 OR2X2_711 ( .A(AES_CORE_DATAPATH__abc_16259_n4027), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n4028) );
  OR2X2 OR2X2_712 ( .A(AES_CORE_DATAPATH__abc_16259_n4030_1), .B(AES_CORE_DATAPATH__abc_16259_n4031_1), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_29_) );
  OR2X2 OR2X2_713 ( .A(AES_CORE_DATAPATH__abc_16259_n2774_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n4033_1), .Y(AES_CORE_DATAPATH__abc_16259_n4034) );
  OR2X2 OR2X2_714 ( .A(AES_CORE_DATAPATH__abc_16259_n2778_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n4035), .Y(AES_CORE_DATAPATH__abc_16259_n4036) );
  OR2X2 OR2X2_715 ( .A(AES_CORE_DATAPATH__abc_16259_n4039_1), .B(AES_CORE_DATAPATH__abc_16259_n4040), .Y(AES_CORE_DATAPATH__abc_16259_n4041_1) );
  OR2X2 OR2X2_716 ( .A(AES_CORE_DATAPATH__abc_16259_n4041_1), .B(AES_CORE_DATAPATH__abc_16259_n4038_1), .Y(AES_CORE_DATAPATH__abc_16259_n4042) );
  OR2X2 OR2X2_717 ( .A(AES_CORE_DATAPATH__abc_16259_n4046_1), .B(AES_CORE_DATAPATH__abc_16259_n2826_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n4047_1) );
  OR2X2 OR2X2_718 ( .A(AES_CORE_DATAPATH__abc_16259_n4048), .B(AES_CORE_DATAPATH__abc_16259_n4049_1), .Y(AES_CORE_DATAPATH__abc_16259_n4050) );
  OR2X2 OR2X2_719 ( .A(AES_CORE_DATAPATH__abc_16259_n4050), .B(AES_CORE_DATAPATH__abc_16259_n4047_1), .Y(AES_CORE_DATAPATH__abc_16259_n4051) );
  OR2X2 OR2X2_72 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n198), .B(AES_CORE_CONTROL_UNIT__abc_15841_n206_1), .Y(AES_CORE_CONTROL_UNIT_sbox_sel_0_) );
  OR2X2 OR2X2_720 ( .A(AES_CORE_DATAPATH__abc_16259_n2841_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__30_), .Y(AES_CORE_DATAPATH__abc_16259_n4052) );
  OR2X2 OR2X2_721 ( .A(AES_CORE_DATAPATH__abc_16259_n4044), .B(AES_CORE_DATAPATH__abc_16259_n2853_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n4054_1) );
  OR2X2 OR2X2_722 ( .A(AES_CORE_DATAPATH__abc_16259_n4055_1), .B(AES_CORE_DATAPATH__abc_16259_n4056), .Y(AES_CORE_DATAPATH__abc_16259_n4057_1) );
  OR2X2 OR2X2_723 ( .A(_auto_iopadmap_cc_313_execute_26949_30_), .B(AES_CORE_DATAPATH__abc_16259_n4059), .Y(AES_CORE_DATAPATH__abc_16259_n4060) );
  OR2X2 OR2X2_724 ( .A(AES_CORE_DATAPATH__abc_16259_n4062_1), .B(AES_CORE_DATAPATH__abc_16259_n2864_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n4063_1) );
  OR2X2 OR2X2_725 ( .A(AES_CORE_DATAPATH__abc_16259_n4063_1), .B(AES_CORE_DATAPATH__abc_16259_n4061), .Y(AES_CORE_DATAPATH__abc_16259_n4064) );
  OR2X2 OR2X2_726 ( .A(AES_CORE_DATAPATH__abc_16259_n4066), .B(AES_CORE_DATAPATH__abc_16259_n4065_1), .Y(AES_CORE_DATAPATH__abc_16259_n4067) );
  OR2X2 OR2X2_727 ( .A(AES_CORE_DATAPATH__abc_16259_n4067), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n4068) );
  OR2X2 OR2X2_728 ( .A(AES_CORE_DATAPATH__abc_16259_n4070_1), .B(AES_CORE_DATAPATH__abc_16259_n4071_1), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_30_) );
  OR2X2 OR2X2_729 ( .A(AES_CORE_DATAPATH__abc_16259_n2774_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n4073_1), .Y(AES_CORE_DATAPATH__abc_16259_n4074) );
  OR2X2 OR2X2_73 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n203_1), .B(AES_CORE_CONTROL_UNIT__abc_15841_n206_1), .Y(AES_CORE_CONTROL_UNIT_sbox_sel_1_) );
  OR2X2 OR2X2_730 ( .A(AES_CORE_DATAPATH__abc_16259_n2778_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n4075), .Y(AES_CORE_DATAPATH__abc_16259_n4076) );
  OR2X2 OR2X2_731 ( .A(AES_CORE_DATAPATH__abc_16259_n4079_1), .B(AES_CORE_DATAPATH__abc_16259_n4080), .Y(AES_CORE_DATAPATH__abc_16259_n4081_1) );
  OR2X2 OR2X2_732 ( .A(AES_CORE_DATAPATH__abc_16259_n4081_1), .B(AES_CORE_DATAPATH__abc_16259_n4078_1), .Y(AES_CORE_DATAPATH__abc_16259_n4082) );
  OR2X2 OR2X2_733 ( .A(AES_CORE_DATAPATH__abc_16259_n4086_1), .B(AES_CORE_DATAPATH__abc_16259_n2826_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n4087_1) );
  OR2X2 OR2X2_734 ( .A(AES_CORE_DATAPATH__abc_16259_n4088), .B(AES_CORE_DATAPATH__abc_16259_n4089_1), .Y(AES_CORE_DATAPATH__abc_16259_n4090) );
  OR2X2 OR2X2_735 ( .A(AES_CORE_DATAPATH__abc_16259_n4090), .B(AES_CORE_DATAPATH__abc_16259_n4087_1), .Y(AES_CORE_DATAPATH__abc_16259_n4091) );
  OR2X2 OR2X2_736 ( .A(AES_CORE_DATAPATH__abc_16259_n2841_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__31_), .Y(AES_CORE_DATAPATH__abc_16259_n4092) );
  OR2X2 OR2X2_737 ( .A(AES_CORE_DATAPATH__abc_16259_n4084), .B(AES_CORE_DATAPATH__abc_16259_n2853_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n4094_1) );
  OR2X2 OR2X2_738 ( .A(AES_CORE_DATAPATH__abc_16259_n4095_1), .B(AES_CORE_DATAPATH__abc_16259_n4096), .Y(AES_CORE_DATAPATH__abc_16259_n4097_1) );
  OR2X2 OR2X2_739 ( .A(_auto_iopadmap_cc_313_execute_26949_31_), .B(AES_CORE_DATAPATH__abc_16259_n4099), .Y(AES_CORE_DATAPATH__abc_16259_n4100) );
  OR2X2 OR2X2_74 ( .A(AES_CORE_DATAPATH__abc_16259_n2459_1), .B(AES_CORE_DATAPATH_col_en_host_1_), .Y(AES_CORE_DATAPATH__abc_16259_n2460) );
  OR2X2 OR2X2_740 ( .A(AES_CORE_DATAPATH__abc_16259_n4102_1), .B(AES_CORE_DATAPATH__abc_16259_n2864_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n4103_1) );
  OR2X2 OR2X2_741 ( .A(AES_CORE_DATAPATH__abc_16259_n4103_1), .B(AES_CORE_DATAPATH__abc_16259_n4101), .Y(AES_CORE_DATAPATH__abc_16259_n4104) );
  OR2X2 OR2X2_742 ( .A(AES_CORE_DATAPATH__abc_16259_n4106), .B(AES_CORE_DATAPATH__abc_16259_n4105_1), .Y(AES_CORE_DATAPATH__abc_16259_n4107) );
  OR2X2 OR2X2_743 ( .A(AES_CORE_DATAPATH__abc_16259_n4107), .B(AES_CORE_DATAPATH__abc_16259_n2796_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n4108) );
  OR2X2 OR2X2_744 ( .A(AES_CORE_DATAPATH__abc_16259_n4110_1), .B(AES_CORE_DATAPATH__abc_16259_n4111_1), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_31_) );
  OR2X2 OR2X2_745 ( .A(AES_CORE_DATAPATH__abc_16259_n4114), .B(AES_CORE_DATAPATH__abc_16259_n4113_1), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_96_) );
  OR2X2 OR2X2_746 ( .A(AES_CORE_DATAPATH__abc_16259_n4117), .B(AES_CORE_DATAPATH__abc_16259_n4116), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_97_) );
  OR2X2 OR2X2_747 ( .A(AES_CORE_DATAPATH__abc_16259_n4120), .B(AES_CORE_DATAPATH__abc_16259_n4119_1), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_98_) );
  OR2X2 OR2X2_748 ( .A(AES_CORE_DATAPATH__abc_16259_n4123), .B(AES_CORE_DATAPATH__abc_16259_n4122), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_99_) );
  OR2X2 OR2X2_749 ( .A(AES_CORE_DATAPATH__abc_16259_n4126_1), .B(AES_CORE_DATAPATH__abc_16259_n4125), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_100_) );
  OR2X2 OR2X2_75 ( .A(AES_CORE_DATAPATH__abc_16259_n2460), .B(AES_CORE_DATAPATH__abc_16259_n2458), .Y(AES_CORE_DATAPATH__abc_16259_n2461_1) );
  OR2X2 OR2X2_750 ( .A(AES_CORE_DATAPATH__abc_16259_n4129_1), .B(AES_CORE_DATAPATH__abc_16259_n4128), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_101_) );
  OR2X2 OR2X2_751 ( .A(AES_CORE_DATAPATH__abc_16259_n4132), .B(AES_CORE_DATAPATH__abc_16259_n4131), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_102_) );
  OR2X2 OR2X2_752 ( .A(AES_CORE_DATAPATH__abc_16259_n4135_1), .B(AES_CORE_DATAPATH__abc_16259_n4134_1), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_103_) );
  OR2X2 OR2X2_753 ( .A(AES_CORE_DATAPATH__abc_16259_n4138), .B(AES_CORE_DATAPATH__abc_16259_n4137_1), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_104_) );
  OR2X2 OR2X2_754 ( .A(AES_CORE_DATAPATH__abc_16259_n4141), .B(AES_CORE_DATAPATH__abc_16259_n4140), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_105_) );
  OR2X2 OR2X2_755 ( .A(AES_CORE_DATAPATH__abc_16259_n4144), .B(AES_CORE_DATAPATH__abc_16259_n4143_1), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_106_) );
  OR2X2 OR2X2_756 ( .A(AES_CORE_DATAPATH__abc_16259_n4147), .B(AES_CORE_DATAPATH__abc_16259_n4146), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_107_) );
  OR2X2 OR2X2_757 ( .A(AES_CORE_DATAPATH__abc_16259_n4150_1), .B(AES_CORE_DATAPATH__abc_16259_n4149), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_108_) );
  OR2X2 OR2X2_758 ( .A(AES_CORE_DATAPATH__abc_16259_n4153_1), .B(AES_CORE_DATAPATH__abc_16259_n4152), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_109_) );
  OR2X2 OR2X2_759 ( .A(AES_CORE_DATAPATH__abc_16259_n4156), .B(AES_CORE_DATAPATH__abc_16259_n4155), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_110_) );
  OR2X2 OR2X2_76 ( .A(AES_CORE_DATAPATH__abc_16259_n2461_1_bF_buf5), .B(\iv_sel_rd[1] ), .Y(AES_CORE_DATAPATH__abc_16259_n2462) );
  OR2X2 OR2X2_760 ( .A(AES_CORE_DATAPATH__abc_16259_n4159_1), .B(AES_CORE_DATAPATH__abc_16259_n4158_1), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_111_) );
  OR2X2 OR2X2_761 ( .A(AES_CORE_DATAPATH__abc_16259_n4162), .B(AES_CORE_DATAPATH__abc_16259_n4161_1), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_112_) );
  OR2X2 OR2X2_762 ( .A(AES_CORE_DATAPATH__abc_16259_n4165), .B(AES_CORE_DATAPATH__abc_16259_n4164), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_113_) );
  OR2X2 OR2X2_763 ( .A(AES_CORE_DATAPATH__abc_16259_n4168), .B(AES_CORE_DATAPATH__abc_16259_n4167_1), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_114_) );
  OR2X2 OR2X2_764 ( .A(AES_CORE_DATAPATH__abc_16259_n4171), .B(AES_CORE_DATAPATH__abc_16259_n4170), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_115_) );
  OR2X2 OR2X2_765 ( .A(AES_CORE_DATAPATH__abc_16259_n4174_1), .B(AES_CORE_DATAPATH__abc_16259_n4173), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_116_) );
  OR2X2 OR2X2_766 ( .A(AES_CORE_DATAPATH__abc_16259_n4177_1), .B(AES_CORE_DATAPATH__abc_16259_n4176), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_117_) );
  OR2X2 OR2X2_767 ( .A(AES_CORE_DATAPATH__abc_16259_n4180), .B(AES_CORE_DATAPATH__abc_16259_n4179), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_118_) );
  OR2X2 OR2X2_768 ( .A(AES_CORE_DATAPATH__abc_16259_n4183_1), .B(AES_CORE_DATAPATH__abc_16259_n4182_1), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_119_) );
  OR2X2 OR2X2_769 ( .A(AES_CORE_DATAPATH__abc_16259_n4186), .B(AES_CORE_DATAPATH__abc_16259_n4185_1), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_120_) );
  OR2X2 OR2X2_77 ( .A(AES_CORE_DATAPATH__abc_16259_n2465_1), .B(AES_CORE_DATAPATH_col_en_host_0_), .Y(AES_CORE_DATAPATH__abc_16259_n2466) );
  OR2X2 OR2X2_770 ( .A(AES_CORE_DATAPATH__abc_16259_n4189), .B(AES_CORE_DATAPATH__abc_16259_n4188), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_121_) );
  OR2X2 OR2X2_771 ( .A(AES_CORE_DATAPATH__abc_16259_n4192), .B(AES_CORE_DATAPATH__abc_16259_n4191_1), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_122_) );
  OR2X2 OR2X2_772 ( .A(AES_CORE_DATAPATH__abc_16259_n4195), .B(AES_CORE_DATAPATH__abc_16259_n4194), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_123_) );
  OR2X2 OR2X2_773 ( .A(AES_CORE_DATAPATH__abc_16259_n4198_1), .B(AES_CORE_DATAPATH__abc_16259_n4197), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_124_) );
  OR2X2 OR2X2_774 ( .A(AES_CORE_DATAPATH__abc_16259_n4201_1), .B(AES_CORE_DATAPATH__abc_16259_n4200), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_125_) );
  OR2X2 OR2X2_775 ( .A(AES_CORE_DATAPATH__abc_16259_n4204), .B(AES_CORE_DATAPATH__abc_16259_n4203), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_126_) );
  OR2X2 OR2X2_776 ( .A(AES_CORE_DATAPATH__abc_16259_n4207_1), .B(AES_CORE_DATAPATH__abc_16259_n4206_1), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_127_) );
  OR2X2 OR2X2_777 ( .A(AES_CORE_DATAPATH__abc_16259_n2804_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_0_), .Y(AES_CORE_DATAPATH__abc_16259_n4209_1) );
  OR2X2 OR2X2_778 ( .A(AES_CORE_DATAPATH__abc_16259_n4213), .B(AES_CORE_DATAPATH__abc_16259_n4211), .Y(AES_CORE_DATAPATH__abc_16259_n4214_1) );
  OR2X2 OR2X2_779 ( .A(AES_CORE_DATAPATH__abc_16259_n4214_1), .B(AES_CORE_DATAPATH__abc_16259_n2807_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n4215_1) );
  OR2X2 OR2X2_78 ( .A(AES_CORE_DATAPATH__abc_16259_n2466), .B(AES_CORE_DATAPATH__abc_16259_n2464), .Y(AES_CORE_DATAPATH__abc_16259_n2467_1) );
  OR2X2 OR2X2_780 ( .A(AES_CORE_DATAPATH__abc_16259_n2804_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_1_), .Y(AES_CORE_DATAPATH__abc_16259_n4217_1) );
  OR2X2 OR2X2_781 ( .A(AES_CORE_DATAPATH__abc_16259_n4221), .B(AES_CORE_DATAPATH__abc_16259_n4219), .Y(AES_CORE_DATAPATH__abc_16259_n4222_1) );
  OR2X2 OR2X2_782 ( .A(AES_CORE_DATAPATH__abc_16259_n4222_1), .B(AES_CORE_DATAPATH__abc_16259_n2807_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n4223_1) );
  OR2X2 OR2X2_783 ( .A(AES_CORE_DATAPATH__abc_16259_n2804_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_2_), .Y(AES_CORE_DATAPATH__abc_16259_n4225_1) );
  OR2X2 OR2X2_784 ( .A(AES_CORE_DATAPATH__abc_16259_n4229), .B(AES_CORE_DATAPATH__abc_16259_n4227), .Y(AES_CORE_DATAPATH__abc_16259_n4230_1) );
  OR2X2 OR2X2_785 ( .A(AES_CORE_DATAPATH__abc_16259_n4230_1), .B(AES_CORE_DATAPATH__abc_16259_n2807_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n4231_1) );
  OR2X2 OR2X2_786 ( .A(AES_CORE_DATAPATH__abc_16259_n2804_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_3_), .Y(AES_CORE_DATAPATH__abc_16259_n4233_1) );
  OR2X2 OR2X2_787 ( .A(AES_CORE_DATAPATH__abc_16259_n4237), .B(AES_CORE_DATAPATH__abc_16259_n4235), .Y(AES_CORE_DATAPATH__abc_16259_n4238_1) );
  OR2X2 OR2X2_788 ( .A(AES_CORE_DATAPATH__abc_16259_n4238_1), .B(AES_CORE_DATAPATH__abc_16259_n2807_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n4239_1) );
  OR2X2 OR2X2_789 ( .A(AES_CORE_DATAPATH__abc_16259_n2804_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_4_), .Y(AES_CORE_DATAPATH__abc_16259_n4241_1) );
  OR2X2 OR2X2_79 ( .A(AES_CORE_DATAPATH__abc_16259_n2467_1_bF_buf5), .B(\iv_sel_rd[0] ), .Y(AES_CORE_DATAPATH__abc_16259_n2468) );
  OR2X2 OR2X2_790 ( .A(AES_CORE_DATAPATH__abc_16259_n4245), .B(AES_CORE_DATAPATH__abc_16259_n4243), .Y(AES_CORE_DATAPATH__abc_16259_n4246_1) );
  OR2X2 OR2X2_791 ( .A(AES_CORE_DATAPATH__abc_16259_n4246_1), .B(AES_CORE_DATAPATH__abc_16259_n2807_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n4247_1) );
  OR2X2 OR2X2_792 ( .A(AES_CORE_DATAPATH__abc_16259_n2804_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_5_), .Y(AES_CORE_DATAPATH__abc_16259_n4249_1) );
  OR2X2 OR2X2_793 ( .A(AES_CORE_DATAPATH__abc_16259_n4253), .B(AES_CORE_DATAPATH__abc_16259_n4251), .Y(AES_CORE_DATAPATH__abc_16259_n4254_1) );
  OR2X2 OR2X2_794 ( .A(AES_CORE_DATAPATH__abc_16259_n4254_1), .B(AES_CORE_DATAPATH__abc_16259_n2807_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n4255_1) );
  OR2X2 OR2X2_795 ( .A(AES_CORE_DATAPATH__abc_16259_n2804_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_6_), .Y(AES_CORE_DATAPATH__abc_16259_n4257_1) );
  OR2X2 OR2X2_796 ( .A(AES_CORE_DATAPATH__abc_16259_n4261), .B(AES_CORE_DATAPATH__abc_16259_n2807_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n4262_1) );
  OR2X2 OR2X2_797 ( .A(AES_CORE_DATAPATH__abc_16259_n4262_1), .B(AES_CORE_DATAPATH__abc_16259_n4259), .Y(AES_CORE_DATAPATH__abc_16259_n4263_1) );
  OR2X2 OR2X2_798 ( .A(AES_CORE_DATAPATH__abc_16259_n2804_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_7_), .Y(AES_CORE_DATAPATH__abc_16259_n4265_1) );
  OR2X2 OR2X2_799 ( .A(AES_CORE_DATAPATH__abc_16259_n4269), .B(AES_CORE_DATAPATH__abc_16259_n2807_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n4270_1) );
  OR2X2 OR2X2_8 ( .A(AES_CORE_CONTROL_UNIT__abc_15841_n101_1), .B(AES_CORE_CONTROL_UNIT__abc_15841_n86_1), .Y(AES_CORE_CONTROL_UNIT__abc_10818_n4) );
  OR2X2 OR2X2_80 ( .A(AES_CORE_DATAPATH__abc_16259_n2472), .B(AES_CORE_DATAPATH_col_en_host_2_), .Y(AES_CORE_DATAPATH__abc_16259_n2473_1) );
  OR2X2 OR2X2_800 ( .A(AES_CORE_DATAPATH__abc_16259_n4270_1), .B(AES_CORE_DATAPATH__abc_16259_n4267), .Y(AES_CORE_DATAPATH__abc_16259_n4271_1) );
  OR2X2 OR2X2_801 ( .A(AES_CORE_DATAPATH__abc_16259_n2804_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_8_), .Y(AES_CORE_DATAPATH__abc_16259_n4273_1) );
  OR2X2 OR2X2_802 ( .A(AES_CORE_DATAPATH__abc_16259_n4277), .B(AES_CORE_DATAPATH__abc_16259_n4275), .Y(AES_CORE_DATAPATH__abc_16259_n4278_1) );
  OR2X2 OR2X2_803 ( .A(AES_CORE_DATAPATH__abc_16259_n4278_1), .B(AES_CORE_DATAPATH__abc_16259_n2807_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n4279_1) );
  OR2X2 OR2X2_804 ( .A(AES_CORE_DATAPATH__abc_16259_n2804_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_9_), .Y(AES_CORE_DATAPATH__abc_16259_n4281_1) );
  OR2X2 OR2X2_805 ( .A(AES_CORE_DATAPATH__abc_16259_n4285), .B(AES_CORE_DATAPATH__abc_16259_n4283), .Y(AES_CORE_DATAPATH__abc_16259_n4286_1) );
  OR2X2 OR2X2_806 ( .A(AES_CORE_DATAPATH__abc_16259_n4286_1), .B(AES_CORE_DATAPATH__abc_16259_n2807_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n4287_1) );
  OR2X2 OR2X2_807 ( .A(AES_CORE_DATAPATH__abc_16259_n2804_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_10_), .Y(AES_CORE_DATAPATH__abc_16259_n4289_1) );
  OR2X2 OR2X2_808 ( .A(AES_CORE_DATAPATH__abc_16259_n4293), .B(AES_CORE_DATAPATH__abc_16259_n4291), .Y(AES_CORE_DATAPATH__abc_16259_n4294_1) );
  OR2X2 OR2X2_809 ( .A(AES_CORE_DATAPATH__abc_16259_n4294_1), .B(AES_CORE_DATAPATH__abc_16259_n2807_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n4295_1) );
  OR2X2 OR2X2_81 ( .A(AES_CORE_DATAPATH__abc_16259_n2473_1), .B(AES_CORE_DATAPATH__abc_16259_n2471_1), .Y(AES_CORE_DATAPATH__abc_16259_n2474) );
  OR2X2 OR2X2_810 ( .A(AES_CORE_DATAPATH__abc_16259_n2804_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_11_), .Y(AES_CORE_DATAPATH__abc_16259_n4297_1) );
  OR2X2 OR2X2_811 ( .A(AES_CORE_DATAPATH__abc_16259_n4301), .B(AES_CORE_DATAPATH__abc_16259_n4299), .Y(AES_CORE_DATAPATH__abc_16259_n4302_1) );
  OR2X2 OR2X2_812 ( .A(AES_CORE_DATAPATH__abc_16259_n4302_1), .B(AES_CORE_DATAPATH__abc_16259_n2807_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n4303_1) );
  OR2X2 OR2X2_813 ( .A(AES_CORE_DATAPATH__abc_16259_n2804_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_12_), .Y(AES_CORE_DATAPATH__abc_16259_n4305_1) );
  OR2X2 OR2X2_814 ( .A(AES_CORE_DATAPATH__abc_16259_n4309), .B(AES_CORE_DATAPATH__abc_16259_n4307), .Y(AES_CORE_DATAPATH__abc_16259_n4310_1) );
  OR2X2 OR2X2_815 ( .A(AES_CORE_DATAPATH__abc_16259_n4310_1), .B(AES_CORE_DATAPATH__abc_16259_n2807_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n4311_1) );
  OR2X2 OR2X2_816 ( .A(AES_CORE_DATAPATH__abc_16259_n4315), .B(AES_CORE_DATAPATH__abc_16259_n4314), .Y(AES_CORE_DATAPATH__abc_16259_n4316) );
  OR2X2 OR2X2_817 ( .A(_auto_iopadmap_cc_313_execute_26949_13_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_5_), .Y(AES_CORE_DATAPATH__abc_16259_n4317) );
  OR2X2 OR2X2_818 ( .A(AES_CORE_DATAPATH__abc_16259_n4319_1), .B(AES_CORE_DATAPATH__abc_16259_n4313_1), .Y(AES_CORE_DATAPATH_sbox_pp2_13__FF_INPUT) );
  OR2X2 OR2X2_819 ( .A(AES_CORE_DATAPATH__abc_16259_n2804_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_14_), .Y(AES_CORE_DATAPATH__abc_16259_n4321_1) );
  OR2X2 OR2X2_82 ( .A(AES_CORE_DATAPATH__abc_16259_n2474_bF_buf5), .B(\iv_sel_rd[2] ), .Y(AES_CORE_DATAPATH__abc_16259_n2475_1) );
  OR2X2 OR2X2_820 ( .A(AES_CORE_DATAPATH__abc_16259_n4325), .B(AES_CORE_DATAPATH__abc_16259_n4323), .Y(AES_CORE_DATAPATH__abc_16259_n4326_1) );
  OR2X2 OR2X2_821 ( .A(AES_CORE_DATAPATH__abc_16259_n4326_1), .B(AES_CORE_DATAPATH__abc_16259_n2807_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n4327_1) );
  OR2X2 OR2X2_822 ( .A(AES_CORE_DATAPATH__abc_16259_n2804_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_15_), .Y(AES_CORE_DATAPATH__abc_16259_n4329_1) );
  OR2X2 OR2X2_823 ( .A(AES_CORE_DATAPATH__abc_16259_n4333), .B(AES_CORE_DATAPATH__abc_16259_n2807_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n4334_1) );
  OR2X2 OR2X2_824 ( .A(AES_CORE_DATAPATH__abc_16259_n4334_1), .B(AES_CORE_DATAPATH__abc_16259_n4331), .Y(AES_CORE_DATAPATH__abc_16259_n4335_1) );
  OR2X2 OR2X2_825 ( .A(AES_CORE_DATAPATH__abc_16259_n2804_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_16_), .Y(AES_CORE_DATAPATH__abc_16259_n4337_1) );
  OR2X2 OR2X2_826 ( .A(AES_CORE_DATAPATH__abc_16259_n4341), .B(AES_CORE_DATAPATH__abc_16259_n4339), .Y(AES_CORE_DATAPATH__abc_16259_n4342_1) );
  OR2X2 OR2X2_827 ( .A(AES_CORE_DATAPATH__abc_16259_n4342_1), .B(AES_CORE_DATAPATH__abc_16259_n2807_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n4343_1) );
  OR2X2 OR2X2_828 ( .A(AES_CORE_DATAPATH__abc_16259_n2804_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_17_), .Y(AES_CORE_DATAPATH__abc_16259_n4345_1) );
  OR2X2 OR2X2_829 ( .A(AES_CORE_DATAPATH__abc_16259_n4349), .B(AES_CORE_DATAPATH__abc_16259_n4347), .Y(AES_CORE_DATAPATH__abc_16259_n4350_1) );
  OR2X2 OR2X2_83 ( .A(AES_CORE_DATAPATH__abc_16259_n2476), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf7), .Y(AES_CORE_DATAPATH__abc_16259_n2477_1) );
  OR2X2 OR2X2_830 ( .A(AES_CORE_DATAPATH__abc_16259_n4350_1), .B(AES_CORE_DATAPATH__abc_16259_n2807_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n4351_1) );
  OR2X2 OR2X2_831 ( .A(AES_CORE_DATAPATH__abc_16259_n2804_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_18_), .Y(AES_CORE_DATAPATH__abc_16259_n4353_1) );
  OR2X2 OR2X2_832 ( .A(AES_CORE_DATAPATH__abc_16259_n4357), .B(AES_CORE_DATAPATH__abc_16259_n4355), .Y(AES_CORE_DATAPATH__abc_16259_n4358_1) );
  OR2X2 OR2X2_833 ( .A(AES_CORE_DATAPATH__abc_16259_n4358_1), .B(AES_CORE_DATAPATH__abc_16259_n2807_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n4359_1) );
  OR2X2 OR2X2_834 ( .A(AES_CORE_DATAPATH__abc_16259_n2804_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_19_), .Y(AES_CORE_DATAPATH__abc_16259_n4361_1) );
  OR2X2 OR2X2_835 ( .A(AES_CORE_DATAPATH__abc_16259_n4365), .B(AES_CORE_DATAPATH__abc_16259_n4363), .Y(AES_CORE_DATAPATH__abc_16259_n4366_1) );
  OR2X2 OR2X2_836 ( .A(AES_CORE_DATAPATH__abc_16259_n4366_1), .B(AES_CORE_DATAPATH__abc_16259_n2807_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n4367_1) );
  OR2X2 OR2X2_837 ( .A(AES_CORE_DATAPATH__abc_16259_n2804_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_20_), .Y(AES_CORE_DATAPATH__abc_16259_n4369_1) );
  OR2X2 OR2X2_838 ( .A(AES_CORE_DATAPATH__abc_16259_n4373), .B(AES_CORE_DATAPATH__abc_16259_n4371), .Y(AES_CORE_DATAPATH__abc_16259_n4374_1) );
  OR2X2 OR2X2_839 ( .A(AES_CORE_DATAPATH__abc_16259_n4374_1), .B(AES_CORE_DATAPATH__abc_16259_n2807_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n4375_1) );
  OR2X2 OR2X2_84 ( .A(AES_CORE_DATAPATH__abc_16259_n2470), .B(AES_CORE_DATAPATH__abc_16259_n2477_1), .Y(AES_CORE_DATAPATH__abc_16259_n2478) );
  OR2X2 OR2X2_840 ( .A(AES_CORE_DATAPATH__abc_16259_n2804_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_21_), .Y(AES_CORE_DATAPATH__abc_16259_n4377_1) );
  OR2X2 OR2X2_841 ( .A(AES_CORE_DATAPATH__abc_16259_n4381), .B(AES_CORE_DATAPATH__abc_16259_n4379), .Y(AES_CORE_DATAPATH__abc_16259_n4382_1) );
  OR2X2 OR2X2_842 ( .A(AES_CORE_DATAPATH__abc_16259_n4382_1), .B(AES_CORE_DATAPATH__abc_16259_n2807_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n4383_1) );
  OR2X2 OR2X2_843 ( .A(AES_CORE_DATAPATH__abc_16259_n2804_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_22_), .Y(AES_CORE_DATAPATH__abc_16259_n4385_1) );
  OR2X2 OR2X2_844 ( .A(AES_CORE_DATAPATH__abc_16259_n4389), .B(AES_CORE_DATAPATH__abc_16259_n4387), .Y(AES_CORE_DATAPATH__abc_16259_n4390_1) );
  OR2X2 OR2X2_845 ( .A(AES_CORE_DATAPATH__abc_16259_n4390_1), .B(AES_CORE_DATAPATH__abc_16259_n2807_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n4391_1) );
  OR2X2 OR2X2_846 ( .A(AES_CORE_DATAPATH__abc_16259_n2804_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_23_), .Y(AES_CORE_DATAPATH__abc_16259_n4393_1) );
  OR2X2 OR2X2_847 ( .A(AES_CORE_DATAPATH__abc_16259_n4397), .B(AES_CORE_DATAPATH__abc_16259_n4395), .Y(AES_CORE_DATAPATH__abc_16259_n4398_1) );
  OR2X2 OR2X2_848 ( .A(AES_CORE_DATAPATH__abc_16259_n4398_1), .B(AES_CORE_DATAPATH__abc_16259_n2807_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n4399_1) );
  OR2X2 OR2X2_849 ( .A(AES_CORE_DATAPATH__abc_16259_n2804_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_24_), .Y(AES_CORE_DATAPATH__abc_16259_n4401_1) );
  OR2X2 OR2X2_85 ( .A(AES_CORE_DATAPATH__abc_16259_n2480), .B(AES_CORE_DATAPATH_col_en_host_3_), .Y(AES_CORE_DATAPATH__abc_16259_n2481_1) );
  OR2X2 OR2X2_850 ( .A(AES_CORE_DATAPATH__abc_16259_n4405), .B(AES_CORE_DATAPATH__abc_16259_n4403), .Y(AES_CORE_DATAPATH__abc_16259_n4406_1) );
  OR2X2 OR2X2_851 ( .A(AES_CORE_DATAPATH__abc_16259_n4406_1), .B(AES_CORE_DATAPATH__abc_16259_n2807_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n4407_1) );
  OR2X2 OR2X2_852 ( .A(AES_CORE_DATAPATH__abc_16259_n2804_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_25_), .Y(AES_CORE_DATAPATH__abc_16259_n4409_1) );
  OR2X2 OR2X2_853 ( .A(AES_CORE_DATAPATH__abc_16259_n4413), .B(AES_CORE_DATAPATH__abc_16259_n4411), .Y(AES_CORE_DATAPATH__abc_16259_n4414_1) );
  OR2X2 OR2X2_854 ( .A(AES_CORE_DATAPATH__abc_16259_n4414_1), .B(AES_CORE_DATAPATH__abc_16259_n2807_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n4415_1) );
  OR2X2 OR2X2_855 ( .A(AES_CORE_DATAPATH__abc_16259_n4419), .B(AES_CORE_DATAPATH__abc_16259_n4418), .Y(AES_CORE_DATAPATH__abc_16259_n4420) );
  OR2X2 OR2X2_856 ( .A(_auto_iopadmap_cc_313_execute_26949_26_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_2_), .Y(AES_CORE_DATAPATH__abc_16259_n4421) );
  OR2X2 OR2X2_857 ( .A(AES_CORE_DATAPATH__abc_16259_n4423_1), .B(AES_CORE_DATAPATH__abc_16259_n4417_1), .Y(AES_CORE_DATAPATH_sbox_pp2_26__FF_INPUT) );
  OR2X2 OR2X2_858 ( .A(AES_CORE_DATAPATH__abc_16259_n2804_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_27_), .Y(AES_CORE_DATAPATH__abc_16259_n4425_1) );
  OR2X2 OR2X2_859 ( .A(AES_CORE_DATAPATH__abc_16259_n4429), .B(AES_CORE_DATAPATH__abc_16259_n4427), .Y(AES_CORE_DATAPATH__abc_16259_n4430_1) );
  OR2X2 OR2X2_86 ( .A(AES_CORE_DATAPATH__abc_16259_n2481_1), .B(AES_CORE_DATAPATH__abc_16259_n2479_1), .Y(AES_CORE_DATAPATH__abc_16259_n2482) );
  OR2X2 OR2X2_860 ( .A(AES_CORE_DATAPATH__abc_16259_n4430_1), .B(AES_CORE_DATAPATH__abc_16259_n2807_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n4431_1) );
  OR2X2 OR2X2_861 ( .A(AES_CORE_DATAPATH__abc_16259_n2804_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_28_), .Y(AES_CORE_DATAPATH__abc_16259_n4433_1) );
  OR2X2 OR2X2_862 ( .A(AES_CORE_DATAPATH__abc_16259_n4437), .B(AES_CORE_DATAPATH__abc_16259_n4435), .Y(AES_CORE_DATAPATH__abc_16259_n4438_1) );
  OR2X2 OR2X2_863 ( .A(AES_CORE_DATAPATH__abc_16259_n4438_1), .B(AES_CORE_DATAPATH__abc_16259_n2807_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n4439) );
  OR2X2 OR2X2_864 ( .A(AES_CORE_DATAPATH__abc_16259_n2804_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_29_), .Y(AES_CORE_DATAPATH__abc_16259_n4441) );
  OR2X2 OR2X2_865 ( .A(AES_CORE_DATAPATH__abc_16259_n4445_1), .B(AES_CORE_DATAPATH__abc_16259_n4443_1), .Y(AES_CORE_DATAPATH__abc_16259_n4446_1) );
  OR2X2 OR2X2_866 ( .A(AES_CORE_DATAPATH__abc_16259_n4446_1), .B(AES_CORE_DATAPATH__abc_16259_n2807_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n4447_1) );
  OR2X2 OR2X2_867 ( .A(AES_CORE_DATAPATH__abc_16259_n2804_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_30_), .Y(AES_CORE_DATAPATH__abc_16259_n4449_1) );
  OR2X2 OR2X2_868 ( .A(AES_CORE_DATAPATH__abc_16259_n4453_1), .B(AES_CORE_DATAPATH__abc_16259_n4451_1), .Y(AES_CORE_DATAPATH__abc_16259_n4454_1) );
  OR2X2 OR2X2_869 ( .A(AES_CORE_DATAPATH__abc_16259_n4454_1), .B(AES_CORE_DATAPATH__abc_16259_n2807_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n4455_1) );
  OR2X2 OR2X2_87 ( .A(AES_CORE_DATAPATH__abc_16259_n2482_bF_buf5), .B(\iv_sel_rd[3] ), .Y(AES_CORE_DATAPATH__abc_16259_n2483_1) );
  OR2X2 OR2X2_870 ( .A(AES_CORE_DATAPATH__abc_16259_n2804_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_31_), .Y(AES_CORE_DATAPATH__abc_16259_n4457_1) );
  OR2X2 OR2X2_871 ( .A(AES_CORE_DATAPATH__abc_16259_n4461_1), .B(AES_CORE_DATAPATH__abc_16259_n2807_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n4462_1) );
  OR2X2 OR2X2_872 ( .A(AES_CORE_DATAPATH__abc_16259_n4462_1), .B(AES_CORE_DATAPATH__abc_16259_n4459_1), .Y(AES_CORE_DATAPATH__abc_16259_n4463_1) );
  OR2X2 OR2X2_873 ( .A(AES_CORE_DATAPATH__abc_16259_n2807_bF_buf0), .B(AES_CORE_CONTROL_UNIT_bypass_rk_bF_buf2), .Y(AES_CORE_DATAPATH_rk_out_sel) );
  OR2X2 OR2X2_874 ( .A(AES_CORE_DATAPATH__abc_16259_n4476_1), .B(AES_CORE_DATAPATH__abc_16259_n4477_1), .Y(AES_CORE_DATAPATH__abc_16259_n4478_1) );
  OR2X2 OR2X2_875 ( .A(AES_CORE_DATAPATH__abc_16259_n4482_1), .B(AES_CORE_DATAPATH__abc_16259_n4481_1), .Y(AES_CORE_DATAPATH__abc_16259_n4483_1) );
  OR2X2 OR2X2_876 ( .A(AES_CORE_DATAPATH__abc_16259_n4484_1), .B(AES_CORE_DATAPATH__abc_16259_n4479_1), .Y(AES_CORE_DATAPATH__abc_16259_n4485_1) );
  OR2X2 OR2X2_877 ( .A(AES_CORE_DATAPATH__abc_16259_n4486_1), .B(AES_CORE_DATAPATH__abc_16259_n4487_1), .Y(AES_CORE_DATAPATH__0key_0__31_0__0_) );
  OR2X2 OR2X2_878 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf9), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_97_), .Y(AES_CORE_DATAPATH__abc_16259_n4489_1) );
  OR2X2 OR2X2_879 ( .A(AES_CORE_DATAPATH__abc_16259_n4490_1), .B(AES_CORE_DATAPATH__abc_16259_n4491_1), .Y(AES_CORE_DATAPATH__abc_16259_n4492_1) );
  OR2X2 OR2X2_88 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf7), .B(AES_CORE_DATAPATH_iv_2__0_), .Y(AES_CORE_DATAPATH__abc_16259_n2486) );
  OR2X2 OR2X2_880 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf8), .B(AES_CORE_DATAPATH__abc_16259_n4492_1), .Y(AES_CORE_DATAPATH__abc_16259_n4493_1) );
  OR2X2 OR2X2_881 ( .A(AES_CORE_DATAPATH__abc_16259_n4495_1), .B(AES_CORE_DATAPATH__abc_16259_n4496_1), .Y(AES_CORE_DATAPATH__0key_0__31_0__1_) );
  OR2X2 OR2X2_882 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf8), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_98_), .Y(AES_CORE_DATAPATH__abc_16259_n4498_1) );
  OR2X2 OR2X2_883 ( .A(AES_CORE_DATAPATH__abc_16259_n4499_1), .B(AES_CORE_DATAPATH__abc_16259_n4500_1), .Y(AES_CORE_DATAPATH__abc_16259_n4501_1) );
  OR2X2 OR2X2_884 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf7), .B(AES_CORE_DATAPATH__abc_16259_n4501_1), .Y(AES_CORE_DATAPATH__abc_16259_n4502_1) );
  OR2X2 OR2X2_885 ( .A(AES_CORE_DATAPATH__abc_16259_n4504_1), .B(AES_CORE_DATAPATH__abc_16259_n4505_1), .Y(AES_CORE_DATAPATH__0key_0__31_0__2_) );
  OR2X2 OR2X2_886 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf7), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_99_), .Y(AES_CORE_DATAPATH__abc_16259_n4507) );
  OR2X2 OR2X2_887 ( .A(AES_CORE_DATAPATH__abc_16259_n4508), .B(AES_CORE_DATAPATH__abc_16259_n4509), .Y(AES_CORE_DATAPATH__abc_16259_n4510_1) );
  OR2X2 OR2X2_888 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf6), .B(AES_CORE_DATAPATH__abc_16259_n4510_1), .Y(AES_CORE_DATAPATH__abc_16259_n4511) );
  OR2X2 OR2X2_889 ( .A(AES_CORE_DATAPATH__abc_16259_n4513_1), .B(AES_CORE_DATAPATH__abc_16259_n4514), .Y(AES_CORE_DATAPATH__0key_0__31_0__3_) );
  OR2X2 OR2X2_89 ( .A(AES_CORE_DATAPATH__abc_16259_n2488), .B(AES_CORE_DATAPATH__abc_16259_n2489_1), .Y(_auto_iopadmap_cc_313_execute_26916_0_) );
  OR2X2 OR2X2_890 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf6), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_100_), .Y(AES_CORE_DATAPATH__abc_16259_n4516_1) );
  OR2X2 OR2X2_891 ( .A(AES_CORE_DATAPATH__abc_16259_n4517), .B(AES_CORE_DATAPATH__abc_16259_n4518), .Y(AES_CORE_DATAPATH__abc_16259_n4519_1) );
  OR2X2 OR2X2_892 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf5), .B(AES_CORE_DATAPATH__abc_16259_n4519_1), .Y(AES_CORE_DATAPATH__abc_16259_n4520) );
  OR2X2 OR2X2_893 ( .A(AES_CORE_DATAPATH__abc_16259_n4521), .B(AES_CORE_DATAPATH__abc_16259_n4474_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n4522_1) );
  OR2X2 OR2X2_894 ( .A(AES_CORE_DATAPATH__abc_16259_n4475_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__4_), .Y(AES_CORE_DATAPATH__abc_16259_n4523) );
  OR2X2 OR2X2_895 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf5), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_101_), .Y(AES_CORE_DATAPATH__abc_16259_n4525_1) );
  OR2X2 OR2X2_896 ( .A(AES_CORE_DATAPATH__abc_16259_n4526), .B(AES_CORE_DATAPATH__abc_16259_n4527), .Y(AES_CORE_DATAPATH__abc_16259_n4528_1) );
  OR2X2 OR2X2_897 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n4528_1), .Y(AES_CORE_DATAPATH__abc_16259_n4529) );
  OR2X2 OR2X2_898 ( .A(AES_CORE_DATAPATH__abc_16259_n4530), .B(AES_CORE_DATAPATH__abc_16259_n4474_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n4531_1) );
  OR2X2 OR2X2_899 ( .A(AES_CORE_DATAPATH__abc_16259_n4475_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__5_), .Y(AES_CORE_DATAPATH__abc_16259_n4532) );
  OR2X2 OR2X2_9 ( .A(AES_CORE_CONTROL_UNIT_rd_count_0_), .B(AES_CORE_CONTROL_UNIT_rd_count_1_), .Y(AES_CORE_CONTROL_UNIT__abc_15841_n109_1) );
  OR2X2 OR2X2_90 ( .A(AES_CORE_DATAPATH__abc_16259_n2492_1), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf5), .Y(AES_CORE_DATAPATH__abc_16259_n2493) );
  OR2X2 OR2X2_900 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_102_), .Y(AES_CORE_DATAPATH__abc_16259_n4534_1) );
  OR2X2 OR2X2_901 ( .A(AES_CORE_DATAPATH__abc_16259_n4535), .B(AES_CORE_DATAPATH__abc_16259_n4536), .Y(AES_CORE_DATAPATH__abc_16259_n4537_1) );
  OR2X2 OR2X2_902 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n4537_1), .Y(AES_CORE_DATAPATH__abc_16259_n4538) );
  OR2X2 OR2X2_903 ( .A(AES_CORE_DATAPATH__abc_16259_n4540_1), .B(AES_CORE_DATAPATH__abc_16259_n4541), .Y(AES_CORE_DATAPATH__0key_0__31_0__6_) );
  OR2X2 OR2X2_904 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_103_), .Y(AES_CORE_DATAPATH__abc_16259_n4543_1) );
  OR2X2 OR2X2_905 ( .A(AES_CORE_DATAPATH__abc_16259_n4544), .B(AES_CORE_DATAPATH__abc_16259_n4545), .Y(AES_CORE_DATAPATH__abc_16259_n4546_1) );
  OR2X2 OR2X2_906 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n4546_1), .Y(AES_CORE_DATAPATH__abc_16259_n4547) );
  OR2X2 OR2X2_907 ( .A(AES_CORE_DATAPATH__abc_16259_n4549_1), .B(AES_CORE_DATAPATH__abc_16259_n4550), .Y(AES_CORE_DATAPATH__0key_0__31_0__7_) );
  OR2X2 OR2X2_908 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_104_), .Y(AES_CORE_DATAPATH__abc_16259_n4552_1) );
  OR2X2 OR2X2_909 ( .A(AES_CORE_DATAPATH__abc_16259_n4553), .B(AES_CORE_DATAPATH__abc_16259_n4554), .Y(AES_CORE_DATAPATH__abc_16259_n4555_1) );
  OR2X2 OR2X2_91 ( .A(AES_CORE_DATAPATH__abc_16259_n2491_1), .B(AES_CORE_DATAPATH__abc_16259_n2493), .Y(AES_CORE_DATAPATH__abc_16259_n2494_1) );
  OR2X2 OR2X2_910 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n4555_1), .Y(AES_CORE_DATAPATH__abc_16259_n4556) );
  OR2X2 OR2X2_911 ( .A(AES_CORE_DATAPATH__abc_16259_n4558_1), .B(AES_CORE_DATAPATH__abc_16259_n4559), .Y(AES_CORE_DATAPATH__0key_0__31_0__8_) );
  OR2X2 OR2X2_912 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_105_), .Y(AES_CORE_DATAPATH__abc_16259_n4561_1) );
  OR2X2 OR2X2_913 ( .A(AES_CORE_DATAPATH__abc_16259_n4562), .B(AES_CORE_DATAPATH__abc_16259_n4563), .Y(AES_CORE_DATAPATH__abc_16259_n4564_1) );
  OR2X2 OR2X2_914 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n4564_1), .Y(AES_CORE_DATAPATH__abc_16259_n4565) );
  OR2X2 OR2X2_915 ( .A(AES_CORE_DATAPATH__abc_16259_n4567_1), .B(AES_CORE_DATAPATH__abc_16259_n4568), .Y(AES_CORE_DATAPATH__0key_0__31_0__9_) );
  OR2X2 OR2X2_916 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_106_), .Y(AES_CORE_DATAPATH__abc_16259_n4570_1) );
  OR2X2 OR2X2_917 ( .A(AES_CORE_DATAPATH__abc_16259_n4571), .B(AES_CORE_DATAPATH__abc_16259_n4572), .Y(AES_CORE_DATAPATH__abc_16259_n4573_1) );
  OR2X2 OR2X2_918 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf10), .B(AES_CORE_DATAPATH__abc_16259_n4573_1), .Y(AES_CORE_DATAPATH__abc_16259_n4574) );
  OR2X2 OR2X2_919 ( .A(AES_CORE_DATAPATH__abc_16259_n4575), .B(AES_CORE_DATAPATH__abc_16259_n4474_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n4576_1) );
  OR2X2 OR2X2_92 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf6), .B(AES_CORE_DATAPATH_iv_2__1_), .Y(AES_CORE_DATAPATH__abc_16259_n2495) );
  OR2X2 OR2X2_920 ( .A(AES_CORE_DATAPATH__abc_16259_n4475_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__10_), .Y(AES_CORE_DATAPATH__abc_16259_n4577) );
  OR2X2 OR2X2_921 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf10), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_107_), .Y(AES_CORE_DATAPATH__abc_16259_n4579_1) );
  OR2X2 OR2X2_922 ( .A(AES_CORE_DATAPATH__abc_16259_n4580), .B(AES_CORE_DATAPATH__abc_16259_n4581), .Y(AES_CORE_DATAPATH__abc_16259_n4582_1) );
  OR2X2 OR2X2_923 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf9), .B(AES_CORE_DATAPATH__abc_16259_n4582_1), .Y(AES_CORE_DATAPATH__abc_16259_n4583) );
  OR2X2 OR2X2_924 ( .A(AES_CORE_DATAPATH__abc_16259_n4585_1), .B(AES_CORE_DATAPATH__abc_16259_n4586), .Y(AES_CORE_DATAPATH__0key_0__31_0__11_) );
  OR2X2 OR2X2_925 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf9), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_108_), .Y(AES_CORE_DATAPATH__abc_16259_n4588_1) );
  OR2X2 OR2X2_926 ( .A(AES_CORE_DATAPATH__abc_16259_n4589), .B(AES_CORE_DATAPATH__abc_16259_n4590), .Y(AES_CORE_DATAPATH__abc_16259_n4591_1) );
  OR2X2 OR2X2_927 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf8), .B(AES_CORE_DATAPATH__abc_16259_n4591_1), .Y(AES_CORE_DATAPATH__abc_16259_n4592) );
  OR2X2 OR2X2_928 ( .A(AES_CORE_DATAPATH__abc_16259_n4594_1), .B(AES_CORE_DATAPATH__abc_16259_n4595), .Y(AES_CORE_DATAPATH__0key_0__31_0__12_) );
  OR2X2 OR2X2_929 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf8), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_109_), .Y(AES_CORE_DATAPATH__abc_16259_n4597_1) );
  OR2X2 OR2X2_93 ( .A(AES_CORE_DATAPATH__abc_16259_n2497_1), .B(AES_CORE_DATAPATH__abc_16259_n2498), .Y(_auto_iopadmap_cc_313_execute_26916_1_) );
  OR2X2 OR2X2_930 ( .A(AES_CORE_DATAPATH__abc_16259_n4598), .B(AES_CORE_DATAPATH__abc_16259_n4599), .Y(AES_CORE_DATAPATH__abc_16259_n4600_1) );
  OR2X2 OR2X2_931 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf7), .B(AES_CORE_DATAPATH__abc_16259_n4600_1), .Y(AES_CORE_DATAPATH__abc_16259_n4601) );
  OR2X2 OR2X2_932 ( .A(AES_CORE_DATAPATH__abc_16259_n4602), .B(AES_CORE_DATAPATH__abc_16259_n4474_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n4603_1) );
  OR2X2 OR2X2_933 ( .A(AES_CORE_DATAPATH__abc_16259_n4475_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__13_), .Y(AES_CORE_DATAPATH__abc_16259_n4604_1) );
  OR2X2 OR2X2_934 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf7), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_110_), .Y(AES_CORE_DATAPATH__abc_16259_n4606) );
  OR2X2 OR2X2_935 ( .A(AES_CORE_DATAPATH__abc_16259_n4607_1), .B(AES_CORE_DATAPATH__abc_16259_n4608), .Y(AES_CORE_DATAPATH__abc_16259_n4609) );
  OR2X2 OR2X2_936 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf6), .B(AES_CORE_DATAPATH__abc_16259_n4609), .Y(AES_CORE_DATAPATH__abc_16259_n4610) );
  OR2X2 OR2X2_937 ( .A(AES_CORE_DATAPATH__abc_16259_n4611_1), .B(AES_CORE_DATAPATH__abc_16259_n4474_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n4612) );
  OR2X2 OR2X2_938 ( .A(AES_CORE_DATAPATH__abc_16259_n4475_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__14_), .Y(AES_CORE_DATAPATH__abc_16259_n4613) );
  OR2X2 OR2X2_939 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf6), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_111_), .Y(AES_CORE_DATAPATH__abc_16259_n4615) );
  OR2X2 OR2X2_94 ( .A(AES_CORE_DATAPATH__abc_16259_n2501_1), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf4), .Y(AES_CORE_DATAPATH__abc_16259_n2502) );
  OR2X2 OR2X2_940 ( .A(AES_CORE_DATAPATH__abc_16259_n4616_1), .B(AES_CORE_DATAPATH__abc_16259_n4617), .Y(AES_CORE_DATAPATH__abc_16259_n4618) );
  OR2X2 OR2X2_941 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf5), .B(AES_CORE_DATAPATH__abc_16259_n4618), .Y(AES_CORE_DATAPATH__abc_16259_n4619) );
  OR2X2 OR2X2_942 ( .A(AES_CORE_DATAPATH__abc_16259_n4621), .B(AES_CORE_DATAPATH__abc_16259_n4622_1), .Y(AES_CORE_DATAPATH__0key_0__31_0__15_) );
  OR2X2 OR2X2_943 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf5), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_112_), .Y(AES_CORE_DATAPATH__abc_16259_n4624) );
  OR2X2 OR2X2_944 ( .A(AES_CORE_DATAPATH__abc_16259_n4625), .B(AES_CORE_DATAPATH__abc_16259_n4626), .Y(AES_CORE_DATAPATH__abc_16259_n4627) );
  OR2X2 OR2X2_945 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n4627), .Y(AES_CORE_DATAPATH__abc_16259_n4628_1) );
  OR2X2 OR2X2_946 ( .A(AES_CORE_DATAPATH__abc_16259_n4630), .B(AES_CORE_DATAPATH__abc_16259_n4631), .Y(AES_CORE_DATAPATH__0key_0__31_0__16_) );
  OR2X2 OR2X2_947 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_113_), .Y(AES_CORE_DATAPATH__abc_16259_n4633) );
  OR2X2 OR2X2_948 ( .A(AES_CORE_DATAPATH__abc_16259_n4634), .B(AES_CORE_DATAPATH__abc_16259_n4635_1), .Y(AES_CORE_DATAPATH__abc_16259_n4636) );
  OR2X2 OR2X2_949 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n4636), .Y(AES_CORE_DATAPATH__abc_16259_n4637) );
  OR2X2 OR2X2_95 ( .A(AES_CORE_DATAPATH__abc_16259_n2500), .B(AES_CORE_DATAPATH__abc_16259_n2502), .Y(AES_CORE_DATAPATH__abc_16259_n2503_1) );
  OR2X2 OR2X2_950 ( .A(AES_CORE_DATAPATH__abc_16259_n4639), .B(AES_CORE_DATAPATH__abc_16259_n4640), .Y(AES_CORE_DATAPATH__0key_0__31_0__17_) );
  OR2X2 OR2X2_951 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_114_), .Y(AES_CORE_DATAPATH__abc_16259_n4642) );
  OR2X2 OR2X2_952 ( .A(AES_CORE_DATAPATH__abc_16259_n4643), .B(AES_CORE_DATAPATH__abc_16259_n4644), .Y(AES_CORE_DATAPATH__abc_16259_n4645) );
  OR2X2 OR2X2_953 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf2), .B(AES_CORE_DATAPATH__abc_16259_n4645), .Y(AES_CORE_DATAPATH__abc_16259_n4646) );
  OR2X2 OR2X2_954 ( .A(AES_CORE_DATAPATH__abc_16259_n4647), .B(AES_CORE_DATAPATH__abc_16259_n4474_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n4648_1) );
  OR2X2 OR2X2_955 ( .A(AES_CORE_DATAPATH__abc_16259_n4475_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__18_), .Y(AES_CORE_DATAPATH__abc_16259_n4649) );
  OR2X2 OR2X2_956 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_115_), .Y(AES_CORE_DATAPATH__abc_16259_n4651) );
  OR2X2 OR2X2_957 ( .A(AES_CORE_DATAPATH__abc_16259_n4652), .B(AES_CORE_DATAPATH__abc_16259_n4653), .Y(AES_CORE_DATAPATH__abc_16259_n4654_1) );
  OR2X2 OR2X2_958 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf1), .B(AES_CORE_DATAPATH__abc_16259_n4654_1), .Y(AES_CORE_DATAPATH__abc_16259_n4655) );
  OR2X2 OR2X2_959 ( .A(AES_CORE_DATAPATH__abc_16259_n4657), .B(AES_CORE_DATAPATH__abc_16259_n4658), .Y(AES_CORE_DATAPATH__0key_0__31_0__19_) );
  OR2X2 OR2X2_96 ( .A(AES_CORE_DATAPATH__abc_16259_n2485_1_bF_buf5), .B(AES_CORE_DATAPATH_iv_2__2_), .Y(AES_CORE_DATAPATH__abc_16259_n2504_1) );
  OR2X2 OR2X2_960 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_116_), .Y(AES_CORE_DATAPATH__abc_16259_n4660) );
  OR2X2 OR2X2_961 ( .A(AES_CORE_DATAPATH__abc_16259_n4661), .B(AES_CORE_DATAPATH__abc_16259_n4662_1), .Y(AES_CORE_DATAPATH__abc_16259_n4663) );
  OR2X2 OR2X2_962 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf0), .B(AES_CORE_DATAPATH__abc_16259_n4663), .Y(AES_CORE_DATAPATH__abc_16259_n4664) );
  OR2X2 OR2X2_963 ( .A(AES_CORE_DATAPATH__abc_16259_n4666), .B(AES_CORE_DATAPATH__abc_16259_n4667), .Y(AES_CORE_DATAPATH__0key_0__31_0__20_) );
  OR2X2 OR2X2_964 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf0), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_117_), .Y(AES_CORE_DATAPATH__abc_16259_n4669) );
  OR2X2 OR2X2_965 ( .A(AES_CORE_DATAPATH__abc_16259_n4670), .B(AES_CORE_DATAPATH__abc_16259_n4671), .Y(AES_CORE_DATAPATH__abc_16259_n4672) );
  OR2X2 OR2X2_966 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf10), .B(AES_CORE_DATAPATH__abc_16259_n4672), .Y(AES_CORE_DATAPATH__abc_16259_n4673) );
  OR2X2 OR2X2_967 ( .A(AES_CORE_DATAPATH__abc_16259_n4674), .B(AES_CORE_DATAPATH__abc_16259_n4474_1_bF_buf2), .Y(AES_CORE_DATAPATH__abc_16259_n4675_1) );
  OR2X2 OR2X2_968 ( .A(AES_CORE_DATAPATH__abc_16259_n4475_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__21_), .Y(AES_CORE_DATAPATH__abc_16259_n4676) );
  OR2X2 OR2X2_969 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf10), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_118_), .Y(AES_CORE_DATAPATH__abc_16259_n4678) );
  OR2X2 OR2X2_97 ( .A(AES_CORE_DATAPATH__abc_16259_n2506_1), .B(AES_CORE_DATAPATH__abc_16259_n2507), .Y(_auto_iopadmap_cc_313_execute_26916_2_) );
  OR2X2 OR2X2_970 ( .A(AES_CORE_DATAPATH__abc_16259_n4679), .B(AES_CORE_DATAPATH__abc_16259_n4680), .Y(AES_CORE_DATAPATH__abc_16259_n4681_1) );
  OR2X2 OR2X2_971 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf9), .B(AES_CORE_DATAPATH__abc_16259_n4681_1), .Y(AES_CORE_DATAPATH__abc_16259_n4682) );
  OR2X2 OR2X2_972 ( .A(AES_CORE_DATAPATH__abc_16259_n4683), .B(AES_CORE_DATAPATH__abc_16259_n4474_1_bF_buf1), .Y(AES_CORE_DATAPATH__abc_16259_n4684) );
  OR2X2 OR2X2_973 ( .A(AES_CORE_DATAPATH__abc_16259_n4475_1_bF_buf2), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__22_), .Y(AES_CORE_DATAPATH__abc_16259_n4685) );
  OR2X2 OR2X2_974 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf9), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_119_), .Y(AES_CORE_DATAPATH__abc_16259_n4687) );
  OR2X2 OR2X2_975 ( .A(AES_CORE_DATAPATH__abc_16259_n4688), .B(AES_CORE_DATAPATH__abc_16259_n4689_1), .Y(AES_CORE_DATAPATH__abc_16259_n4690) );
  OR2X2 OR2X2_976 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf8), .B(AES_CORE_DATAPATH__abc_16259_n4690), .Y(AES_CORE_DATAPATH__abc_16259_n4691) );
  OR2X2 OR2X2_977 ( .A(AES_CORE_DATAPATH__abc_16259_n4693), .B(AES_CORE_DATAPATH__abc_16259_n4694), .Y(AES_CORE_DATAPATH__0key_0__31_0__23_) );
  OR2X2 OR2X2_978 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf8), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_120_), .Y(AES_CORE_DATAPATH__abc_16259_n4696) );
  OR2X2 OR2X2_979 ( .A(AES_CORE_DATAPATH__abc_16259_n4697), .B(AES_CORE_DATAPATH__abc_16259_n4698), .Y(AES_CORE_DATAPATH__abc_16259_n4699) );
  OR2X2 OR2X2_98 ( .A(AES_CORE_DATAPATH__abc_16259_n2510), .B(AES_CORE_DATAPATH__abc_16259_n2475_1_bF_buf3), .Y(AES_CORE_DATAPATH__abc_16259_n2511_1) );
  OR2X2 OR2X2_980 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf7), .B(AES_CORE_DATAPATH__abc_16259_n4699), .Y(AES_CORE_DATAPATH__abc_16259_n4700) );
  OR2X2 OR2X2_981 ( .A(AES_CORE_DATAPATH__abc_16259_n4702_1), .B(AES_CORE_DATAPATH__abc_16259_n4703), .Y(AES_CORE_DATAPATH__0key_0__31_0__24_) );
  OR2X2 OR2X2_982 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf7), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_121_), .Y(AES_CORE_DATAPATH__abc_16259_n4705) );
  OR2X2 OR2X2_983 ( .A(AES_CORE_DATAPATH__abc_16259_n4706), .B(AES_CORE_DATAPATH__abc_16259_n4707), .Y(AES_CORE_DATAPATH__abc_16259_n4708_1) );
  OR2X2 OR2X2_984 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf6), .B(AES_CORE_DATAPATH__abc_16259_n4708_1), .Y(AES_CORE_DATAPATH__abc_16259_n4709) );
  OR2X2 OR2X2_985 ( .A(AES_CORE_DATAPATH__abc_16259_n4711), .B(AES_CORE_DATAPATH__abc_16259_n4712), .Y(AES_CORE_DATAPATH__0key_0__31_0__25_) );
  OR2X2 OR2X2_986 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf6), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_122_), .Y(AES_CORE_DATAPATH__abc_16259_n4714) );
  OR2X2 OR2X2_987 ( .A(AES_CORE_DATAPATH__abc_16259_n4715), .B(AES_CORE_DATAPATH__abc_16259_n4716), .Y(AES_CORE_DATAPATH__abc_16259_n4717_1) );
  OR2X2 OR2X2_988 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf5), .B(AES_CORE_DATAPATH__abc_16259_n4717_1), .Y(AES_CORE_DATAPATH__abc_16259_n4718) );
  OR2X2 OR2X2_989 ( .A(AES_CORE_DATAPATH__abc_16259_n4720), .B(AES_CORE_DATAPATH__abc_16259_n4721), .Y(AES_CORE_DATAPATH__0key_0__31_0__26_) );
  OR2X2 OR2X2_99 ( .A(AES_CORE_DATAPATH__abc_16259_n2509_1), .B(AES_CORE_DATAPATH__abc_16259_n2511_1), .Y(AES_CORE_DATAPATH__abc_16259_n2512) );
  OR2X2 OR2X2_990 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf5), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_123_), .Y(AES_CORE_DATAPATH__abc_16259_n4723_1) );
  OR2X2 OR2X2_991 ( .A(AES_CORE_DATAPATH__abc_16259_n4724), .B(AES_CORE_DATAPATH__abc_16259_n4725), .Y(AES_CORE_DATAPATH__abc_16259_n4726) );
  OR2X2 OR2X2_992 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf4), .B(AES_CORE_DATAPATH__abc_16259_n4726), .Y(AES_CORE_DATAPATH__abc_16259_n4727) );
  OR2X2 OR2X2_993 ( .A(AES_CORE_DATAPATH__abc_16259_n4729), .B(AES_CORE_DATAPATH__abc_16259_n4730_1), .Y(AES_CORE_DATAPATH__0key_0__31_0__27_) );
  OR2X2 OR2X2_994 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf4), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_124_), .Y(AES_CORE_DATAPATH__abc_16259_n4732) );
  OR2X2 OR2X2_995 ( .A(AES_CORE_DATAPATH__abc_16259_n4733), .B(AES_CORE_DATAPATH__abc_16259_n4734), .Y(AES_CORE_DATAPATH__abc_16259_n4735) );
  OR2X2 OR2X2_996 ( .A(AES_CORE_DATAPATH__abc_16259_n4478_1_bF_buf3), .B(AES_CORE_DATAPATH__abc_16259_n4735), .Y(AES_CORE_DATAPATH__abc_16259_n4736_1) );
  OR2X2 OR2X2_997 ( .A(AES_CORE_DATAPATH__abc_16259_n4737), .B(AES_CORE_DATAPATH__abc_16259_n4474_1_bF_buf0), .Y(AES_CORE_DATAPATH__abc_16259_n4738) );
  OR2X2 OR2X2_998 ( .A(AES_CORE_DATAPATH__abc_16259_n4475_1_bF_buf1), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__28_), .Y(AES_CORE_DATAPATH__abc_16259_n4739) );
  OR2X2 OR2X2_999 ( .A(AES_CORE_DATAPATH__abc_16259_n4480_1_bF_buf3), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_125_), .Y(AES_CORE_DATAPATH__abc_16259_n4741) );
endmodule
