module b09_reset(clock, RESET_G, nRESET_G, X, Y_REG);

wire D_IN_REG_0_; 
wire D_IN_REG_1_; 
wire D_IN_REG_2_; 
wire D_IN_REG_3_; 
wire D_IN_REG_4_; 
wire D_IN_REG_5_; 
wire D_IN_REG_6_; 
wire D_IN_REG_7_; 
wire D_IN_REG_8_; 
wire D_OUT_REG_0_; 
wire D_OUT_REG_1_; 
wire D_OUT_REG_2_; 
wire D_OUT_REG_3_; 
wire D_OUT_REG_4_; 
wire D_OUT_REG_5_; 
wire D_OUT_REG_6_; 
wire D_OUT_REG_7_; 
wire OLD_REG_0_; 
wire OLD_REG_1_; 
wire OLD_REG_2_; 
wire OLD_REG_3_; 
wire OLD_REG_4_; 
wire OLD_REG_5_; 
wire OLD_REG_6_; 
wire OLD_REG_7_; 
input RESET_G;
wire STATO_REG_0_; 
wire STATO_REG_1_; 
input X;
output Y_REG;
wire _abc_898_new_n100_; 
wire _abc_898_new_n101_; 
wire _abc_898_new_n102_; 
wire _abc_898_new_n103_; 
wire _abc_898_new_n104_; 
wire _abc_898_new_n105_; 
wire _abc_898_new_n106_; 
wire _abc_898_new_n107_; 
wire _abc_898_new_n108_; 
wire _abc_898_new_n109_; 
wire _abc_898_new_n110_; 
wire _abc_898_new_n111_; 
wire _abc_898_new_n112_; 
wire _abc_898_new_n113_; 
wire _abc_898_new_n114_; 
wire _abc_898_new_n115_; 
wire _abc_898_new_n116_; 
wire _abc_898_new_n117_; 
wire _abc_898_new_n118_; 
wire _abc_898_new_n120_; 
wire _abc_898_new_n121_; 
wire _abc_898_new_n122_; 
wire _abc_898_new_n123_; 
wire _abc_898_new_n124_; 
wire _abc_898_new_n125_; 
wire _abc_898_new_n126_; 
wire _abc_898_new_n127_; 
wire _abc_898_new_n129_; 
wire _abc_898_new_n130_; 
wire _abc_898_new_n131_; 
wire _abc_898_new_n140_; 
wire _abc_898_new_n141_; 
wire _abc_898_new_n142_; 
wire _abc_898_new_n143_; 
wire _abc_898_new_n144_; 
wire _abc_898_new_n145_; 
wire _abc_898_new_n146_; 
wire _abc_898_new_n147_; 
wire _abc_898_new_n148_; 
wire _abc_898_new_n150_; 
wire _abc_898_new_n151_; 
wire _abc_898_new_n152_; 
wire _abc_898_new_n154_; 
wire _abc_898_new_n155_; 
wire _abc_898_new_n156_; 
wire _abc_898_new_n158_; 
wire _abc_898_new_n159_; 
wire _abc_898_new_n160_; 
wire _abc_898_new_n162_; 
wire _abc_898_new_n163_; 
wire _abc_898_new_n164_; 
wire _abc_898_new_n166_; 
wire _abc_898_new_n167_; 
wire _abc_898_new_n168_; 
wire _abc_898_new_n170_; 
wire _abc_898_new_n171_; 
wire _abc_898_new_n172_; 
wire _abc_898_new_n174_; 
wire _abc_898_new_n175_; 
wire _abc_898_new_n176_; 
wire _abc_898_new_n178_; 
wire _abc_898_new_n179_; 
wire _abc_898_new_n180_; 
wire _abc_898_new_n182_; 
wire _abc_898_new_n183_; 
wire _abc_898_new_n184_; 
wire _abc_898_new_n185_; 
wire _abc_898_new_n186_; 
wire _abc_898_new_n187_; 
wire _abc_898_new_n188_; 
wire _abc_898_new_n189_; 
wire _abc_898_new_n191_; 
wire _abc_898_new_n192_; 
wire _abc_898_new_n193_; 
wire _abc_898_new_n194_; 
wire _abc_898_new_n195_; 
wire _abc_898_new_n197_; 
wire _abc_898_new_n198_; 
wire _abc_898_new_n199_; 
wire _abc_898_new_n200_; 
wire _abc_898_new_n201_; 
wire _abc_898_new_n203_; 
wire _abc_898_new_n204_; 
wire _abc_898_new_n205_; 
wire _abc_898_new_n206_; 
wire _abc_898_new_n207_; 
wire _abc_898_new_n209_; 
wire _abc_898_new_n210_; 
wire _abc_898_new_n211_; 
wire _abc_898_new_n212_; 
wire _abc_898_new_n213_; 
wire _abc_898_new_n215_; 
wire _abc_898_new_n216_; 
wire _abc_898_new_n217_; 
wire _abc_898_new_n218_; 
wire _abc_898_new_n219_; 
wire _abc_898_new_n221_; 
wire _abc_898_new_n222_; 
wire _abc_898_new_n223_; 
wire _abc_898_new_n225_; 
wire _abc_898_new_n226_; 
wire _abc_898_new_n227_; 
wire _abc_898_new_n228_; 
wire _abc_898_new_n229_; 
wire _abc_898_new_n59_; 
wire _abc_898_new_n60_; 
wire _abc_898_new_n61_; 
wire _abc_898_new_n63_; 
wire _abc_898_new_n64_; 
wire _abc_898_new_n65_; 
wire _abc_898_new_n66_; 
wire _abc_898_new_n67_; 
wire _abc_898_new_n68_; 
wire _abc_898_new_n69_; 
wire _abc_898_new_n70_; 
wire _abc_898_new_n71_; 
wire _abc_898_new_n72_; 
wire _abc_898_new_n73_; 
wire _abc_898_new_n74_; 
wire _abc_898_new_n75_; 
wire _abc_898_new_n76_; 
wire _abc_898_new_n77_; 
wire _abc_898_new_n78_; 
wire _abc_898_new_n79_; 
wire _abc_898_new_n80_; 
wire _abc_898_new_n81_; 
wire _abc_898_new_n82_; 
wire _abc_898_new_n83_; 
wire _abc_898_new_n84_; 
wire _abc_898_new_n85_; 
wire _abc_898_new_n86_; 
wire _abc_898_new_n87_; 
wire _abc_898_new_n88_; 
wire _abc_898_new_n89_; 
wire _abc_898_new_n90_; 
wire _abc_898_new_n91_; 
wire _abc_898_new_n92_; 
wire _abc_898_new_n93_; 
wire _abc_898_new_n94_; 
wire _abc_898_new_n95_; 
wire _abc_898_new_n96_; 
wire _abc_898_new_n97_; 
wire _abc_898_new_n98_; 
wire _abc_898_new_n99_; 
input clock;
wire n10; 
wire n104; 
wire n109; 
wire n114; 
wire n119; 
wire n124; 
wire n129; 
wire n134; 
wire n139; 
wire n144; 
wire n15; 
wire n20; 
wire n25; 
wire n30; 
wire n35; 
wire n40; 
wire n45; 
wire n50; 
wire n55; 
wire n60; 
wire n65; 
wire n70; 
wire n75; 
wire n80; 
wire n85; 
wire n90; 
wire n95; 
wire n99; 
input nRESET_G;
AND2X2 AND2X2_1 ( .A(_abc_898_new_n130_), .B(OLD_REG_3_), .Y(_abc_898_new_n162_));
AND2X2 AND2X2_10 ( .A(_abc_898_new_n59_), .B(D_IN_REG_8_), .Y(_abc_898_new_n179_));
AND2X2 AND2X2_11 ( .A(_abc_898_new_n129_), .B(_abc_898_new_n182_), .Y(_abc_898_new_n183_));
AND2X2 AND2X2_12 ( .A(_abc_898_new_n140_), .B(_abc_898_new_n183_), .Y(_abc_898_new_n184_));
AND2X2 AND2X2_13 ( .A(_abc_898_new_n184_), .B(D_OUT_REG_0_), .Y(_abc_898_new_n185_));
AND2X2 AND2X2_14 ( .A(_abc_898_new_n120_), .B(_abc_898_new_n151_), .Y(_abc_898_new_n186_));
AND2X2 AND2X2_15 ( .A(_abc_898_new_n143_), .B(D_OUT_REG_1_), .Y(_abc_898_new_n187_));
AND2X2 AND2X2_16 ( .A(_abc_898_new_n184_), .B(D_OUT_REG_1_), .Y(_abc_898_new_n191_));
AND2X2 AND2X2_17 ( .A(_abc_898_new_n120_), .B(_abc_898_new_n155_), .Y(_abc_898_new_n192_));
AND2X2 AND2X2_18 ( .A(_abc_898_new_n143_), .B(D_OUT_REG_2_), .Y(_abc_898_new_n193_));
AND2X2 AND2X2_19 ( .A(_abc_898_new_n184_), .B(D_OUT_REG_2_), .Y(_abc_898_new_n197_));
AND2X2 AND2X2_2 ( .A(_abc_898_new_n59_), .B(D_IN_REG_4_), .Y(_abc_898_new_n163_));
AND2X2 AND2X2_20 ( .A(_abc_898_new_n120_), .B(_abc_898_new_n159_), .Y(_abc_898_new_n198_));
AND2X2 AND2X2_21 ( .A(_abc_898_new_n143_), .B(D_OUT_REG_3_), .Y(_abc_898_new_n199_));
AND2X2 AND2X2_22 ( .A(_abc_898_new_n184_), .B(D_OUT_REG_3_), .Y(_abc_898_new_n203_));
AND2X2 AND2X2_23 ( .A(_abc_898_new_n120_), .B(_abc_898_new_n163_), .Y(_abc_898_new_n204_));
AND2X2 AND2X2_24 ( .A(_abc_898_new_n143_), .B(D_OUT_REG_4_), .Y(_abc_898_new_n205_));
AND2X2 AND2X2_25 ( .A(_abc_898_new_n184_), .B(D_OUT_REG_4_), .Y(_abc_898_new_n209_));
AND2X2 AND2X2_26 ( .A(_abc_898_new_n120_), .B(_abc_898_new_n167_), .Y(_abc_898_new_n210_));
AND2X2 AND2X2_27 ( .A(_abc_898_new_n143_), .B(D_OUT_REG_5_), .Y(_abc_898_new_n211_));
AND2X2 AND2X2_28 ( .A(_abc_898_new_n184_), .B(D_OUT_REG_5_), .Y(_abc_898_new_n215_));
AND2X2 AND2X2_29 ( .A(_abc_898_new_n120_), .B(_abc_898_new_n171_), .Y(_abc_898_new_n216_));
AND2X2 AND2X2_3 ( .A(_abc_898_new_n130_), .B(OLD_REG_4_), .Y(_abc_898_new_n166_));
AND2X2 AND2X2_30 ( .A(_abc_898_new_n143_), .B(D_OUT_REG_6_), .Y(_abc_898_new_n217_));
AND2X2 AND2X2_31 ( .A(_abc_898_new_n184_), .B(D_OUT_REG_7_), .Y(_abc_898_new_n221_));
AND2X2 AND2X2_32 ( .A(_abc_898_new_n120_), .B(_abc_898_new_n179_), .Y(_abc_898_new_n222_));
AND2X2 AND2X2_33 ( .A(_abc_898_new_n184_), .B(D_OUT_REG_6_), .Y(_abc_898_new_n225_));
AND2X2 AND2X2_34 ( .A(_abc_898_new_n120_), .B(_abc_898_new_n175_), .Y(_abc_898_new_n226_));
AND2X2 AND2X2_35 ( .A(_abc_898_new_n143_), .B(D_OUT_REG_7_), .Y(_abc_898_new_n227_));
AND2X2 AND2X2_36 ( .A(D_IN_REG_0_), .B(STATO_REG_0_), .Y(_abc_898_new_n59_));
AND2X2 AND2X2_37 ( .A(_abc_898_new_n65_), .B(_abc_898_new_n67_), .Y(_abc_898_new_n68_));
AND2X2 AND2X2_38 ( .A(_abc_898_new_n70_), .B(_abc_898_new_n72_), .Y(_abc_898_new_n73_));
AND2X2 AND2X2_39 ( .A(_abc_898_new_n68_), .B(_abc_898_new_n73_), .Y(_abc_898_new_n74_));
AND2X2 AND2X2_4 ( .A(_abc_898_new_n59_), .B(D_IN_REG_5_), .Y(_abc_898_new_n167_));
AND2X2 AND2X2_40 ( .A(_abc_898_new_n76_), .B(_abc_898_new_n78_), .Y(_abc_898_new_n79_));
AND2X2 AND2X2_41 ( .A(_abc_898_new_n81_), .B(_abc_898_new_n83_), .Y(_abc_898_new_n84_));
AND2X2 AND2X2_42 ( .A(_abc_898_new_n79_), .B(_abc_898_new_n84_), .Y(_abc_898_new_n85_));
AND2X2 AND2X2_43 ( .A(_abc_898_new_n74_), .B(_abc_898_new_n85_), .Y(_abc_898_new_n86_));
AND2X2 AND2X2_44 ( .A(_abc_898_new_n88_), .B(_abc_898_new_n90_), .Y(_abc_898_new_n91_));
AND2X2 AND2X2_45 ( .A(_abc_898_new_n93_), .B(_abc_898_new_n95_), .Y(_abc_898_new_n96_));
AND2X2 AND2X2_46 ( .A(_abc_898_new_n91_), .B(_abc_898_new_n96_), .Y(_abc_898_new_n97_));
AND2X2 AND2X2_47 ( .A(_abc_898_new_n99_), .B(_abc_898_new_n101_), .Y(_abc_898_new_n102_));
AND2X2 AND2X2_48 ( .A(_abc_898_new_n104_), .B(_abc_898_new_n106_), .Y(_abc_898_new_n107_));
AND2X2 AND2X2_49 ( .A(_abc_898_new_n102_), .B(_abc_898_new_n107_), .Y(_abc_898_new_n108_));
AND2X2 AND2X2_5 ( .A(_abc_898_new_n130_), .B(OLD_REG_5_), .Y(_abc_898_new_n170_));
AND2X2 AND2X2_50 ( .A(_abc_898_new_n97_), .B(_abc_898_new_n108_), .Y(_abc_898_new_n109_));
AND2X2 AND2X2_51 ( .A(_abc_898_new_n86_), .B(_abc_898_new_n109_), .Y(_abc_898_new_n110_));
AND2X2 AND2X2_52 ( .A(_abc_898_new_n110_), .B(STATO_REG_1_), .Y(_abc_898_new_n111_));
AND2X2 AND2X2_53 ( .A(_abc_898_new_n112_), .B(STATO_REG_0_), .Y(_abc_898_new_n113_));
AND2X2 AND2X2_54 ( .A(_abc_898_new_n116_), .B(_abc_898_new_n114_), .Y(_abc_898_new_n117_));
AND2X2 AND2X2_55 ( .A(_abc_898_new_n120_), .B(_abc_898_new_n59_), .Y(_abc_898_new_n121_));
AND2X2 AND2X2_56 ( .A(_abc_898_new_n115_), .B(STATO_REG_0_), .Y(_abc_898_new_n122_));
AND2X2 AND2X2_57 ( .A(_abc_898_new_n123_), .B(STATO_REG_1_), .Y(_abc_898_new_n124_));
AND2X2 AND2X2_58 ( .A(_abc_898_new_n125_), .B(X), .Y(_abc_898_new_n126_));
AND2X2 AND2X2_59 ( .A(_abc_898_new_n125_), .B(_abc_898_new_n129_), .Y(_abc_898_new_n130_));
AND2X2 AND2X2_6 ( .A(_abc_898_new_n59_), .B(D_IN_REG_6_), .Y(_abc_898_new_n171_));
AND2X2 AND2X2_60 ( .A(_abc_898_new_n130_), .B(nRESET_G), .Y(_abc_898_new_n131_));
AND2X2 AND2X2_61 ( .A(_abc_898_new_n131_), .B(D_IN_REG_1_), .Y(n10));
AND2X2 AND2X2_62 ( .A(_abc_898_new_n131_), .B(D_IN_REG_2_), .Y(n144));
AND2X2 AND2X2_63 ( .A(_abc_898_new_n131_), .B(D_IN_REG_3_), .Y(n139));
AND2X2 AND2X2_64 ( .A(_abc_898_new_n131_), .B(D_IN_REG_4_), .Y(n134));
AND2X2 AND2X2_65 ( .A(_abc_898_new_n131_), .B(D_IN_REG_5_), .Y(n129));
AND2X2 AND2X2_66 ( .A(_abc_898_new_n131_), .B(D_IN_REG_6_), .Y(n124));
AND2X2 AND2X2_67 ( .A(_abc_898_new_n131_), .B(D_IN_REG_7_), .Y(n119));
AND2X2 AND2X2_68 ( .A(_abc_898_new_n131_), .B(D_IN_REG_8_), .Y(n114));
AND2X2 AND2X2_69 ( .A(_abc_898_new_n114_), .B(STATO_REG_1_), .Y(_abc_898_new_n142_));
AND2X2 AND2X2_7 ( .A(_abc_898_new_n130_), .B(OLD_REG_6_), .Y(_abc_898_new_n174_));
AND2X2 AND2X2_70 ( .A(_abc_898_new_n142_), .B(_abc_898_new_n63_), .Y(_abc_898_new_n143_));
AND2X2 AND2X2_71 ( .A(_abc_898_new_n143_), .B(D_OUT_REG_0_), .Y(_abc_898_new_n144_));
AND2X2 AND2X2_72 ( .A(_abc_898_new_n122_), .B(_abc_898_new_n145_), .Y(_abc_898_new_n146_));
AND2X2 AND2X2_73 ( .A(_abc_898_new_n130_), .B(OLD_REG_0_), .Y(_abc_898_new_n150_));
AND2X2 AND2X2_74 ( .A(_abc_898_new_n59_), .B(D_IN_REG_1_), .Y(_abc_898_new_n151_));
AND2X2 AND2X2_75 ( .A(_abc_898_new_n130_), .B(OLD_REG_1_), .Y(_abc_898_new_n154_));
AND2X2 AND2X2_76 ( .A(_abc_898_new_n59_), .B(D_IN_REG_2_), .Y(_abc_898_new_n155_));
AND2X2 AND2X2_77 ( .A(_abc_898_new_n130_), .B(OLD_REG_2_), .Y(_abc_898_new_n158_));
AND2X2 AND2X2_78 ( .A(_abc_898_new_n59_), .B(D_IN_REG_3_), .Y(_abc_898_new_n159_));
AND2X2 AND2X2_8 ( .A(_abc_898_new_n59_), .B(D_IN_REG_7_), .Y(_abc_898_new_n175_));
AND2X2 AND2X2_9 ( .A(_abc_898_new_n130_), .B(OLD_REG_7_), .Y(_abc_898_new_n178_));
DFFPOSX1 DFFPOSX1_1 ( .CLK(clock), .D(n25), .Q(D_OUT_REG_5_));
DFFPOSX1 DFFPOSX1_10 ( .CLK(clock), .D(n50), .Q(D_OUT_REG_0_));
DFFPOSX1 DFFPOSX1_11 ( .CLK(clock), .D(n55), .Q(OLD_REG_7_));
DFFPOSX1 DFFPOSX1_12 ( .CLK(clock), .D(n60), .Q(OLD_REG_6_));
DFFPOSX1 DFFPOSX1_13 ( .CLK(clock), .D(n65), .Q(OLD_REG_5_));
DFFPOSX1 DFFPOSX1_14 ( .CLK(clock), .D(n70), .Q(OLD_REG_4_));
DFFPOSX1 DFFPOSX1_15 ( .CLK(clock), .D(n75), .Q(OLD_REG_3_));
DFFPOSX1 DFFPOSX1_16 ( .CLK(clock), .D(n80), .Q(OLD_REG_2_));
DFFPOSX1 DFFPOSX1_17 ( .CLK(clock), .D(n85), .Q(OLD_REG_1_));
DFFPOSX1 DFFPOSX1_18 ( .CLK(clock), .D(n90), .Q(OLD_REG_0_));
DFFPOSX1 DFFPOSX1_19 ( .CLK(clock), .D(n99), .Q(STATO_REG_1_));
DFFPOSX1 DFFPOSX1_2 ( .CLK(clock), .D(n15), .Q(D_OUT_REG_7_));
DFFPOSX1 DFFPOSX1_20 ( .CLK(clock), .D(n104), .Q(STATO_REG_0_));
DFFPOSX1 DFFPOSX1_21 ( .CLK(clock), .D(n109), .Q(D_IN_REG_8_));
DFFPOSX1 DFFPOSX1_22 ( .CLK(clock), .D(n114), .Q(D_IN_REG_7_));
DFFPOSX1 DFFPOSX1_23 ( .CLK(clock), .D(n119), .Q(D_IN_REG_6_));
DFFPOSX1 DFFPOSX1_24 ( .CLK(clock), .D(n124), .Q(D_IN_REG_5_));
DFFPOSX1 DFFPOSX1_25 ( .CLK(clock), .D(n129), .Q(D_IN_REG_4_));
DFFPOSX1 DFFPOSX1_26 ( .CLK(clock), .D(n134), .Q(D_IN_REG_3_));
DFFPOSX1 DFFPOSX1_27 ( .CLK(clock), .D(n139), .Q(D_IN_REG_2_));
DFFPOSX1 DFFPOSX1_28 ( .CLK(clock), .D(n144), .Q(D_IN_REG_1_));
DFFPOSX1 DFFPOSX1_3 ( .CLK(clock), .D(n10), .Q(D_IN_REG_0_));
DFFPOSX1 DFFPOSX1_4 ( .CLK(clock), .D(n20), .Q(D_OUT_REG_6_));
DFFPOSX1 DFFPOSX1_5 ( .CLK(clock), .D(n95), .Q(Y_REG));
DFFPOSX1 DFFPOSX1_6 ( .CLK(clock), .D(n30), .Q(D_OUT_REG_4_));
DFFPOSX1 DFFPOSX1_7 ( .CLK(clock), .D(n35), .Q(D_OUT_REG_3_));
DFFPOSX1 DFFPOSX1_8 ( .CLK(clock), .D(n40), .Q(D_OUT_REG_2_));
DFFPOSX1 DFFPOSX1_9 ( .CLK(clock), .D(n45), .Q(D_OUT_REG_1_));
INVX1 INVX1_1 ( .A(nRESET_G), .Y(_abc_898_new_n60_));
INVX1 INVX1_10 ( .A(OLD_REG_3_), .Y(_abc_898_new_n82_));
INVX1 INVX1_11 ( .A(OLD_REG_4_), .Y(_abc_898_new_n87_));
INVX1 INVX1_12 ( .A(D_IN_REG_5_), .Y(_abc_898_new_n89_));
INVX1 INVX1_13 ( .A(D_IN_REG_6_), .Y(_abc_898_new_n92_));
INVX1 INVX1_14 ( .A(OLD_REG_5_), .Y(_abc_898_new_n94_));
INVX1 INVX1_15 ( .A(OLD_REG_0_), .Y(_abc_898_new_n98_));
INVX1 INVX1_16 ( .A(D_IN_REG_1_), .Y(_abc_898_new_n100_));
INVX1 INVX1_17 ( .A(D_IN_REG_2_), .Y(_abc_898_new_n103_));
INVX1 INVX1_18 ( .A(OLD_REG_1_), .Y(_abc_898_new_n105_));
INVX1 INVX1_19 ( .A(STATO_REG_0_), .Y(_abc_898_new_n114_));
INVX1 INVX1_2 ( .A(D_IN_REG_0_), .Y(_abc_898_new_n63_));
INVX1 INVX1_20 ( .A(STATO_REG_1_), .Y(_abc_898_new_n115_));
INVX1 INVX1_21 ( .A(_abc_898_new_n111_), .Y(_abc_898_new_n120_));
INVX1 INVX1_22 ( .A(_abc_898_new_n59_), .Y(_abc_898_new_n123_));
INVX1 INVX1_23 ( .A(_abc_898_new_n140_), .Y(_abc_898_new_n141_));
INVX1 INVX1_3 ( .A(OLD_REG_7_), .Y(_abc_898_new_n64_));
INVX1 INVX1_4 ( .A(D_IN_REG_8_), .Y(_abc_898_new_n66_));
INVX1 INVX1_5 ( .A(D_IN_REG_7_), .Y(_abc_898_new_n69_));
INVX1 INVX1_6 ( .A(OLD_REG_6_), .Y(_abc_898_new_n71_));
INVX1 INVX1_7 ( .A(OLD_REG_2_), .Y(_abc_898_new_n75_));
INVX1 INVX1_8 ( .A(D_IN_REG_3_), .Y(_abc_898_new_n77_));
INVX1 INVX1_9 ( .A(D_IN_REG_4_), .Y(_abc_898_new_n80_));
OR2X2 OR2X2_1 ( .A(_abc_898_new_n159_), .B(_abc_898_new_n60_), .Y(_abc_898_new_n160_));
OR2X2 OR2X2_10 ( .A(_abc_898_new_n174_), .B(_abc_898_new_n176_), .Y(n60));
OR2X2 OR2X2_11 ( .A(_abc_898_new_n179_), .B(_abc_898_new_n60_), .Y(_abc_898_new_n180_));
OR2X2 OR2X2_12 ( .A(_abc_898_new_n178_), .B(_abc_898_new_n180_), .Y(n55));
OR2X2 OR2X2_13 ( .A(D_IN_REG_0_), .B(STATO_REG_0_), .Y(_abc_898_new_n182_));
OR2X2 OR2X2_14 ( .A(_abc_898_new_n187_), .B(_abc_898_new_n60_), .Y(_abc_898_new_n188_));
OR2X2 OR2X2_15 ( .A(_abc_898_new_n186_), .B(_abc_898_new_n188_), .Y(_abc_898_new_n189_));
OR2X2 OR2X2_16 ( .A(_abc_898_new_n189_), .B(_abc_898_new_n185_), .Y(n50));
OR2X2 OR2X2_17 ( .A(_abc_898_new_n193_), .B(_abc_898_new_n60_), .Y(_abc_898_new_n194_));
OR2X2 OR2X2_18 ( .A(_abc_898_new_n192_), .B(_abc_898_new_n194_), .Y(_abc_898_new_n195_));
OR2X2 OR2X2_19 ( .A(_abc_898_new_n195_), .B(_abc_898_new_n191_), .Y(n45));
OR2X2 OR2X2_2 ( .A(_abc_898_new_n158_), .B(_abc_898_new_n160_), .Y(n80));
OR2X2 OR2X2_20 ( .A(_abc_898_new_n199_), .B(_abc_898_new_n60_), .Y(_abc_898_new_n200_));
OR2X2 OR2X2_21 ( .A(_abc_898_new_n198_), .B(_abc_898_new_n200_), .Y(_abc_898_new_n201_));
OR2X2 OR2X2_22 ( .A(_abc_898_new_n201_), .B(_abc_898_new_n197_), .Y(n40));
OR2X2 OR2X2_23 ( .A(_abc_898_new_n205_), .B(_abc_898_new_n60_), .Y(_abc_898_new_n206_));
OR2X2 OR2X2_24 ( .A(_abc_898_new_n204_), .B(_abc_898_new_n206_), .Y(_abc_898_new_n207_));
OR2X2 OR2X2_25 ( .A(_abc_898_new_n207_), .B(_abc_898_new_n203_), .Y(n35));
OR2X2 OR2X2_26 ( .A(_abc_898_new_n211_), .B(_abc_898_new_n60_), .Y(_abc_898_new_n212_));
OR2X2 OR2X2_27 ( .A(_abc_898_new_n210_), .B(_abc_898_new_n212_), .Y(_abc_898_new_n213_));
OR2X2 OR2X2_28 ( .A(_abc_898_new_n213_), .B(_abc_898_new_n209_), .Y(n30));
OR2X2 OR2X2_29 ( .A(_abc_898_new_n217_), .B(_abc_898_new_n60_), .Y(_abc_898_new_n218_));
OR2X2 OR2X2_3 ( .A(_abc_898_new_n163_), .B(_abc_898_new_n60_), .Y(_abc_898_new_n164_));
OR2X2 OR2X2_30 ( .A(_abc_898_new_n216_), .B(_abc_898_new_n218_), .Y(_abc_898_new_n219_));
OR2X2 OR2X2_31 ( .A(_abc_898_new_n219_), .B(_abc_898_new_n215_), .Y(n25));
OR2X2 OR2X2_32 ( .A(_abc_898_new_n222_), .B(_abc_898_new_n60_), .Y(_abc_898_new_n223_));
OR2X2 OR2X2_33 ( .A(_abc_898_new_n223_), .B(_abc_898_new_n221_), .Y(n15));
OR2X2 OR2X2_34 ( .A(_abc_898_new_n227_), .B(_abc_898_new_n60_), .Y(_abc_898_new_n228_));
OR2X2 OR2X2_35 ( .A(_abc_898_new_n226_), .B(_abc_898_new_n228_), .Y(_abc_898_new_n229_));
OR2X2 OR2X2_36 ( .A(_abc_898_new_n229_), .B(_abc_898_new_n225_), .Y(n20));
OR2X2 OR2X2_37 ( .A(_abc_898_new_n60_), .B(STATO_REG_1_), .Y(_abc_898_new_n61_));
OR2X2 OR2X2_38 ( .A(_abc_898_new_n61_), .B(_abc_898_new_n59_), .Y(n99));
OR2X2 OR2X2_39 ( .A(_abc_898_new_n64_), .B(D_IN_REG_8_), .Y(_abc_898_new_n65_));
OR2X2 OR2X2_4 ( .A(_abc_898_new_n162_), .B(_abc_898_new_n164_), .Y(n75));
OR2X2 OR2X2_40 ( .A(_abc_898_new_n66_), .B(OLD_REG_7_), .Y(_abc_898_new_n67_));
OR2X2 OR2X2_41 ( .A(_abc_898_new_n69_), .B(OLD_REG_6_), .Y(_abc_898_new_n70_));
OR2X2 OR2X2_42 ( .A(_abc_898_new_n71_), .B(D_IN_REG_7_), .Y(_abc_898_new_n72_));
OR2X2 OR2X2_43 ( .A(_abc_898_new_n75_), .B(D_IN_REG_3_), .Y(_abc_898_new_n76_));
OR2X2 OR2X2_44 ( .A(_abc_898_new_n77_), .B(OLD_REG_2_), .Y(_abc_898_new_n78_));
OR2X2 OR2X2_45 ( .A(_abc_898_new_n80_), .B(OLD_REG_3_), .Y(_abc_898_new_n81_));
OR2X2 OR2X2_46 ( .A(_abc_898_new_n82_), .B(D_IN_REG_4_), .Y(_abc_898_new_n83_));
OR2X2 OR2X2_47 ( .A(_abc_898_new_n87_), .B(D_IN_REG_5_), .Y(_abc_898_new_n88_));
OR2X2 OR2X2_48 ( .A(_abc_898_new_n89_), .B(OLD_REG_4_), .Y(_abc_898_new_n90_));
OR2X2 OR2X2_49 ( .A(_abc_898_new_n92_), .B(OLD_REG_5_), .Y(_abc_898_new_n93_));
OR2X2 OR2X2_5 ( .A(_abc_898_new_n167_), .B(_abc_898_new_n60_), .Y(_abc_898_new_n168_));
OR2X2 OR2X2_50 ( .A(_abc_898_new_n94_), .B(D_IN_REG_6_), .Y(_abc_898_new_n95_));
OR2X2 OR2X2_51 ( .A(_abc_898_new_n98_), .B(D_IN_REG_1_), .Y(_abc_898_new_n99_));
OR2X2 OR2X2_52 ( .A(_abc_898_new_n100_), .B(OLD_REG_0_), .Y(_abc_898_new_n101_));
OR2X2 OR2X2_53 ( .A(_abc_898_new_n103_), .B(OLD_REG_1_), .Y(_abc_898_new_n104_));
OR2X2 OR2X2_54 ( .A(_abc_898_new_n105_), .B(D_IN_REG_2_), .Y(_abc_898_new_n106_));
OR2X2 OR2X2_55 ( .A(_abc_898_new_n111_), .B(_abc_898_new_n63_), .Y(_abc_898_new_n112_));
OR2X2 OR2X2_56 ( .A(_abc_898_new_n115_), .B(D_IN_REG_0_), .Y(_abc_898_new_n116_));
OR2X2 OR2X2_57 ( .A(_abc_898_new_n117_), .B(_abc_898_new_n60_), .Y(_abc_898_new_n118_));
OR2X2 OR2X2_58 ( .A(_abc_898_new_n113_), .B(_abc_898_new_n118_), .Y(n104));
OR2X2 OR2X2_59 ( .A(_abc_898_new_n124_), .B(_abc_898_new_n122_), .Y(_abc_898_new_n125_));
OR2X2 OR2X2_6 ( .A(_abc_898_new_n166_), .B(_abc_898_new_n168_), .Y(n70));
OR2X2 OR2X2_60 ( .A(_abc_898_new_n126_), .B(_abc_898_new_n60_), .Y(_abc_898_new_n127_));
OR2X2 OR2X2_61 ( .A(_abc_898_new_n121_), .B(_abc_898_new_n127_), .Y(n109));
OR2X2 OR2X2_62 ( .A(_abc_898_new_n63_), .B(STATO_REG_1_), .Y(_abc_898_new_n129_));
OR2X2 OR2X2_63 ( .A(_abc_898_new_n110_), .B(_abc_898_new_n123_), .Y(_abc_898_new_n140_));
OR2X2 OR2X2_64 ( .A(D_IN_REG_0_), .B(Y_REG), .Y(_abc_898_new_n145_));
OR2X2 OR2X2_65 ( .A(_abc_898_new_n146_), .B(_abc_898_new_n60_), .Y(_abc_898_new_n147_));
OR2X2 OR2X2_66 ( .A(_abc_898_new_n147_), .B(_abc_898_new_n144_), .Y(_abc_898_new_n148_));
OR2X2 OR2X2_67 ( .A(_abc_898_new_n141_), .B(_abc_898_new_n148_), .Y(n95));
OR2X2 OR2X2_68 ( .A(_abc_898_new_n151_), .B(_abc_898_new_n60_), .Y(_abc_898_new_n152_));
OR2X2 OR2X2_69 ( .A(_abc_898_new_n150_), .B(_abc_898_new_n152_), .Y(n90));
OR2X2 OR2X2_7 ( .A(_abc_898_new_n171_), .B(_abc_898_new_n60_), .Y(_abc_898_new_n172_));
OR2X2 OR2X2_70 ( .A(_abc_898_new_n155_), .B(_abc_898_new_n60_), .Y(_abc_898_new_n156_));
OR2X2 OR2X2_71 ( .A(_abc_898_new_n154_), .B(_abc_898_new_n156_), .Y(n85));
OR2X2 OR2X2_8 ( .A(_abc_898_new_n170_), .B(_abc_898_new_n172_), .Y(n65));
OR2X2 OR2X2_9 ( .A(_abc_898_new_n175_), .B(_abc_898_new_n60_), .Y(_abc_898_new_n176_));


endmodule