module FSM(clk, reset, \codif[0] , \codif[1] , \codif[2] , \codif[3] , \codif[4] , \codif[5] , \codif[6] , \codif[7] , \codif[8] , \codif[9] , \codif[10] , \codif[11] , busy_mem, done_mem, aligned_mem, done_exec, is_exec, \W_R_mem[0] , \W_R_mem[1] , \wordsize_mem[0] , \wordsize_mem[1] , sign_mem, en_mem, enable_exec, enable_exec_mem, trap, enable_pc);

output \W_R_mem[0] ;
output \W_R_mem[1] ;
wire _0W_R_mem_1_0__0_; 
wire _0W_R_mem_1_0__1_; 
wire _0en_mem_0_0_; 
wire _0enable_exec_0_0_; 
wire _0enable_exec_mem_0_0_; 
wire _0enable_pc_aux_0_0_; 
wire _0enable_pc_fsm_0_0_; 
wire _0trap_0_0_; 
wire _abc_801_auto_fsm_map_cc_170_map_fsm_238_0_; 
wire _abc_801_auto_fsm_map_cc_170_map_fsm_238_1_; 
wire _abc_801_auto_fsm_map_cc_170_map_fsm_238_2_; 
wire _abc_801_auto_fsm_map_cc_170_map_fsm_238_3_; 
wire _abc_801_auto_fsm_map_cc_170_map_fsm_238_4_; 
wire _abc_801_auto_fsm_map_cc_170_map_fsm_238_5_; 
wire _abc_801_auto_fsm_map_cc_170_map_fsm_238_6_; 
wire _abc_934_new_n100_; 
wire _abc_934_new_n102_; 
wire _abc_934_new_n103_; 
wire _abc_934_new_n104_; 
wire _abc_934_new_n105_; 
wire _abc_934_new_n106_; 
wire _abc_934_new_n107_; 
wire _abc_934_new_n108_; 
wire _abc_934_new_n109_; 
wire _abc_934_new_n110_; 
wire _abc_934_new_n111_; 
wire _abc_934_new_n112_; 
wire _abc_934_new_n113_; 
wire _abc_934_new_n114_; 
wire _abc_934_new_n116_; 
wire _abc_934_new_n117_; 
wire _abc_934_new_n118_; 
wire _abc_934_new_n119_; 
wire _abc_934_new_n120_; 
wire _abc_934_new_n123_; 
wire _abc_934_new_n124_; 
wire _abc_934_new_n125_; 
wire _abc_934_new_n126_; 
wire _abc_934_new_n127_; 
wire _abc_934_new_n129_; 
wire _abc_934_new_n131_; 
wire _abc_934_new_n132_; 
wire _abc_934_new_n133_; 
wire _abc_934_new_n134_; 
wire _abc_934_new_n136_; 
wire _abc_934_new_n137_; 
wire _abc_934_new_n138_; 
wire _abc_934_new_n139_; 
wire _abc_934_new_n141_; 
wire _abc_934_new_n49_; 
wire _abc_934_new_n50_; 
wire _abc_934_new_n51_; 
wire _abc_934_new_n52_; 
wire _abc_934_new_n53_; 
wire _abc_934_new_n54_; 
wire _abc_934_new_n55_; 
wire _abc_934_new_n56_; 
wire _abc_934_new_n57_; 
wire _abc_934_new_n58_; 
wire _abc_934_new_n59_; 
wire _abc_934_new_n60_; 
wire _abc_934_new_n61_; 
wire _abc_934_new_n62_; 
wire _abc_934_new_n63_; 
wire _abc_934_new_n64_; 
wire _abc_934_new_n65_; 
wire _abc_934_new_n66_; 
wire _abc_934_new_n67_; 
wire _abc_934_new_n68_; 
wire _abc_934_new_n69_; 
wire _abc_934_new_n70_; 
wire _abc_934_new_n71_; 
wire _abc_934_new_n72_; 
wire _abc_934_new_n73_; 
wire _abc_934_new_n74_; 
wire _abc_934_new_n76_; 
wire _abc_934_new_n77_; 
wire _abc_934_new_n78_; 
wire _abc_934_new_n80_; 
wire _abc_934_new_n81_; 
wire _abc_934_new_n82_; 
wire _abc_934_new_n83_; 
wire _abc_934_new_n85_; 
wire _abc_934_new_n86_; 
wire _abc_934_new_n87_; 
wire _abc_934_new_n88_; 
wire _abc_934_new_n89_; 
wire _abc_934_new_n90_; 
wire _abc_934_new_n91_; 
wire _abc_934_new_n92_; 
wire _abc_934_new_n94_; 
wire _abc_934_new_n95_; 
wire _abc_934_new_n97_; 
wire _auto_iopadmap_cc_368_execute_1030_0_; 
wire _auto_iopadmap_cc_368_execute_1030_1_; 
wire _auto_iopadmap_cc_368_execute_1033; 
wire _auto_iopadmap_cc_368_execute_1035; 
wire _auto_iopadmap_cc_368_execute_1037; 
wire _auto_iopadmap_cc_368_execute_1039; 
wire _auto_iopadmap_cc_368_execute_1041; 
wire _auto_iopadmap_cc_368_execute_1043; 
input aligned_mem;
input busy_mem;
input clk;
input \codif[0] ;
input \codif[10] ;
input \codif[11] ;
input \codif[1] ;
input \codif[2] ;
input \codif[3] ;
input \codif[4] ;
input \codif[5] ;
input \codif[6] ;
input \codif[7] ;
input \codif[8] ;
input \codif[9] ;
input done_exec;
input done_mem;
output en_mem;
output enable_exec;
output enable_exec_mem;
output enable_pc;
wire enable_pc_aux; 
wire enable_pc_fsm; 
input is_exec;
input reset;
output sign_mem;
wire state_0_; 
wire state_1_; 
wire state_2_; 
wire state_3_; 
wire state_4_; 
wire state_5_; 
wire state_6_; 
output trap;
output \wordsize_mem[0] ;
output \wordsize_mem[1] ;
AND2X2 AND2X2_1 ( .A(\codif[0] ), .B(\codif[1] ), .Y(_abc_934_new_n53_));
AND2X2 AND2X2_2 ( .A(_abc_934_new_n57_), .B(state_2_), .Y(_abc_934_new_n58_));
AND2X2 AND2X2_3 ( .A(\codif[2] ), .B(\codif[3] ), .Y(_abc_934_new_n63_));
AND2X2 AND2X2_4 ( .A(_abc_934_new_n53_), .B(_abc_934_new_n63_), .Y(_abc_934_new_n64_));
AND2X2 AND2X2_5 ( .A(_abc_934_new_n53_), .B(_abc_934_new_n54_), .Y(_abc_934_new_n69_));
AND2X2 AND2X2_6 ( .A(_abc_934_new_n70_), .B(_abc_934_new_n71_), .Y(_abc_934_new_n72_));
AOI21X1 AOI21X1_1 ( .A(_abc_934_new_n107_), .B(_abc_934_new_n114_), .C(_abc_934_new_n49_), .Y(_0W_R_mem_1_0__0_));
AOI21X1 AOI21X1_10 ( .A(_abc_934_new_n80_), .B(_abc_934_new_n83_), .C(_abc_934_new_n82_), .Y(_abc_801_auto_fsm_map_cc_170_map_fsm_238_3_));
AOI21X1 AOI21X1_11 ( .A(aligned_mem), .B(_abc_934_new_n89_), .C(_abc_934_new_n91_), .Y(_abc_934_new_n92_));
AOI21X1 AOI21X1_12 ( .A(_auto_iopadmap_cc_368_execute_1033), .B(state_0_), .C(state_5_), .Y(_abc_934_new_n97_));
AOI21X1 AOI21X1_2 ( .A(_abc_934_new_n118_), .B(_abc_934_new_n120_), .C(_abc_934_new_n49_), .Y(_0W_R_mem_1_0__1_));
AOI21X1 AOI21X1_3 ( .A(_abc_934_new_n56_), .B(_abc_934_new_n58_), .C(state_4_), .Y(_abc_934_new_n125_));
AOI21X1 AOI21X1_4 ( .A(_abc_934_new_n100_), .B(_abc_934_new_n74_), .C(_abc_934_new_n127_), .Y(_0enable_pc_fsm_0_0_));
AOI21X1 AOI21X1_5 ( .A(_abc_934_new_n76_), .B(_abc_934_new_n129_), .C(_abc_934_new_n49_), .Y(_0trap_0_0_));
AOI21X1 AOI21X1_6 ( .A(_abc_934_new_n131_), .B(_abc_934_new_n81_), .C(_abc_934_new_n132_), .Y(_abc_934_new_n133_));
AOI21X1 AOI21X1_7 ( .A(_abc_934_new_n136_), .B(_abc_934_new_n74_), .C(_abc_934_new_n139_), .Y(_0enable_exec_0_0_));
AOI21X1 AOI21X1_8 ( .A(_abc_934_new_n74_), .B(_abc_934_new_n59_), .C(_abc_934_new_n52_), .Y(_abc_801_auto_fsm_map_cc_170_map_fsm_238_2_));
AOI21X1 AOI21X1_9 ( .A(_abc_934_new_n78_), .B(_abc_934_new_n76_), .C(_abc_934_new_n49_), .Y(_abc_801_auto_fsm_map_cc_170_map_fsm_238_1_));
AOI22X1 AOI22X1_1 ( .A(_auto_iopadmap_cc_368_execute_1033), .B(done_mem), .C(_abc_934_new_n88_), .D(_abc_934_new_n83_), .Y(_abc_934_new_n116_));
AOI22X1 AOI22X1_2 ( .A(_abc_934_new_n94_), .B(_abc_934_new_n104_), .C(_auto_iopadmap_cc_368_execute_1033), .D(_abc_934_new_n117_), .Y(_abc_934_new_n141_));
BUFX2 BUFX2_1 ( .A(_auto_iopadmap_cc_368_execute_1030_0_), .Y(\W_R_mem[0] ));
BUFX2 BUFX2_10 ( .A(\codif[8] ), .Y(\wordsize_mem[1] ));
BUFX2 BUFX2_2 ( .A(_auto_iopadmap_cc_368_execute_1030_1_), .Y(\W_R_mem[1] ));
BUFX2 BUFX2_3 ( .A(_auto_iopadmap_cc_368_execute_1033), .Y(en_mem));
BUFX2 BUFX2_4 ( .A(_auto_iopadmap_cc_368_execute_1035), .Y(enable_exec));
BUFX2 BUFX2_5 ( .A(_auto_iopadmap_cc_368_execute_1037), .Y(enable_exec_mem));
BUFX2 BUFX2_6 ( .A(_auto_iopadmap_cc_368_execute_1039), .Y(enable_pc));
BUFX2 BUFX2_7 ( .A(_auto_iopadmap_cc_368_execute_1041), .Y(sign_mem));
BUFX2 BUFX2_8 ( .A(_auto_iopadmap_cc_368_execute_1043), .Y(trap));
BUFX2 BUFX2_9 ( .A(\codif[7] ), .Y(\wordsize_mem[0] ));
DFFPOSX1 DFFPOSX1_1 ( .CLK(clk), .D(_abc_801_auto_fsm_map_cc_170_map_fsm_238_0_), .Q(state_0_));
DFFPOSX1 DFFPOSX1_10 ( .CLK(clk), .D(_0en_mem_0_0_), .Q(_auto_iopadmap_cc_368_execute_1033));
DFFPOSX1 DFFPOSX1_11 ( .CLK(clk), .D(_0enable_exec_0_0_), .Q(_auto_iopadmap_cc_368_execute_1035));
DFFPOSX1 DFFPOSX1_12 ( .CLK(clk), .D(_0enable_exec_mem_0_0_), .Q(_auto_iopadmap_cc_368_execute_1037));
DFFPOSX1 DFFPOSX1_13 ( .CLK(clk), .D(_0trap_0_0_), .Q(_auto_iopadmap_cc_368_execute_1043));
DFFPOSX1 DFFPOSX1_14 ( .CLK(clk), .D(_0enable_pc_fsm_0_0_), .Q(enable_pc_fsm));
DFFPOSX1 DFFPOSX1_15 ( .CLK(clk), .D(_0enable_pc_aux_0_0_), .Q(enable_pc_aux));
DFFPOSX1 DFFPOSX1_2 ( .CLK(clk), .D(_abc_801_auto_fsm_map_cc_170_map_fsm_238_1_), .Q(state_1_));
DFFPOSX1 DFFPOSX1_3 ( .CLK(clk), .D(_abc_801_auto_fsm_map_cc_170_map_fsm_238_2_), .Q(state_2_));
DFFPOSX1 DFFPOSX1_4 ( .CLK(clk), .D(_abc_801_auto_fsm_map_cc_170_map_fsm_238_3_), .Q(state_3_));
DFFPOSX1 DFFPOSX1_5 ( .CLK(clk), .D(_abc_801_auto_fsm_map_cc_170_map_fsm_238_4_), .Q(state_4_));
DFFPOSX1 DFFPOSX1_6 ( .CLK(clk), .D(_abc_801_auto_fsm_map_cc_170_map_fsm_238_5_), .Q(state_5_));
DFFPOSX1 DFFPOSX1_7 ( .CLK(clk), .D(_abc_801_auto_fsm_map_cc_170_map_fsm_238_6_), .Q(state_6_));
DFFPOSX1 DFFPOSX1_8 ( .CLK(clk), .D(_0W_R_mem_1_0__0_), .Q(_auto_iopadmap_cc_368_execute_1030_0_));
DFFPOSX1 DFFPOSX1_9 ( .CLK(clk), .D(_0W_R_mem_1_0__1_), .Q(_auto_iopadmap_cc_368_execute_1030_1_));
INVX1 INVX1_1 ( .A(\codif[9] ), .Y(_auto_iopadmap_cc_368_execute_1041));
INVX1 INVX1_10 ( .A(_abc_934_new_n105_), .Y(_abc_934_new_n106_));
INVX1 INVX1_11 ( .A(_auto_iopadmap_cc_368_execute_1030_0_), .Y(_abc_934_new_n108_));
INVX1 INVX1_2 ( .A(_auto_iopadmap_cc_368_execute_1043), .Y(_abc_934_new_n129_));
INVX1 INVX1_3 ( .A(_auto_iopadmap_cc_368_execute_1035), .Y(_abc_934_new_n136_));
INVX1 INVX1_4 ( .A(_abc_934_new_n51_), .Y(_abc_934_new_n52_));
INVX1 INVX1_5 ( .A(done_exec), .Y(_abc_934_new_n57_));
INVX1 INVX1_6 ( .A(state_3_), .Y(_abc_934_new_n80_));
INVX1 INVX1_7 ( .A(_abc_934_new_n56_), .Y(_abc_934_new_n85_));
INVX1 INVX1_8 ( .A(enable_pc_fsm), .Y(_abc_934_new_n100_));
INVX1 INVX1_9 ( .A(state_6_), .Y(_abc_934_new_n103_));
INVX2 INVX2_1 ( .A(reset), .Y(_abc_934_new_n49_));
INVX2 INVX2_2 ( .A(done_mem), .Y(_abc_934_new_n81_));
INVX2 INVX2_3 ( .A(state_0_), .Y(_abc_934_new_n88_));
INVX4 INVX4_1 ( .A(aligned_mem), .Y(_abc_934_new_n50_));
NAND2X1 NAND2X1_1 ( .A(aligned_mem), .B(_abc_934_new_n113_), .Y(_abc_934_new_n114_));
NAND2X1 NAND2X1_10 ( .A(_abc_934_new_n68_), .B(_abc_934_new_n73_), .Y(_abc_934_new_n77_));
NAND2X1 NAND2X1_11 ( .A(state_4_), .B(_abc_934_new_n77_), .Y(_abc_934_new_n78_));
NAND2X1 NAND2X1_12 ( .A(_abc_934_new_n81_), .B(_abc_934_new_n51_), .Y(_abc_934_new_n82_));
NAND2X1 NAND2X1_13 ( .A(state_6_), .B(_auto_iopadmap_cc_368_execute_1033), .Y(_abc_934_new_n83_));
NAND2X1 NAND2X1_14 ( .A(state_2_), .B(_abc_934_new_n51_), .Y(_abc_934_new_n86_));
NAND2X1 NAND2X1_15 ( .A(done_mem), .B(_abc_934_new_n51_), .Y(_abc_934_new_n90_));
NAND2X1 NAND2X1_16 ( .A(_abc_934_new_n103_), .B(_abc_934_new_n88_), .Y(_abc_934_new_n104_));
NAND2X1 NAND2X1_2 ( .A(reset), .B(_abc_934_new_n126_), .Y(_abc_934_new_n127_));
NAND2X1 NAND2X1_3 ( .A(reset), .B(_auto_iopadmap_cc_368_execute_1037), .Y(_abc_934_new_n134_));
NAND2X1 NAND2X1_4 ( .A(reset), .B(_abc_934_new_n138_), .Y(_abc_934_new_n139_));
NAND2X1 NAND2X1_5 ( .A(_abc_934_new_n58_), .B(_abc_934_new_n56_), .Y(_abc_934_new_n59_));
NAND2X1 NAND2X1_6 ( .A(\codif[4] ), .B(\codif[5] ), .Y(_abc_934_new_n60_));
NAND2X1 NAND2X1_7 ( .A(\codif[6] ), .B(\codif[7] ), .Y(_abc_934_new_n61_));
NAND2X1 NAND2X1_8 ( .A(\codif[10] ), .B(\codif[11] ), .Y(_abc_934_new_n65_));
NAND2X1 NAND2X1_9 ( .A(\codif[8] ), .B(\codif[9] ), .Y(_abc_934_new_n66_));
NAND3X1 NAND3X1_1 ( .A(aligned_mem), .B(_abc_934_new_n109_), .C(_abc_934_new_n105_), .Y(_abc_934_new_n117_));
NAND3X1 NAND3X1_2 ( .A(aligned_mem), .B(_abc_934_new_n119_), .C(_abc_934_new_n105_), .Y(_abc_934_new_n120_));
NAND3X1 NAND3X1_3 ( .A(_abc_934_new_n54_), .B(_abc_934_new_n55_), .C(_abc_934_new_n53_), .Y(_abc_934_new_n56_));
NAND3X1 NAND3X1_4 ( .A(_abc_934_new_n62_), .B(_abc_934_new_n67_), .C(_abc_934_new_n64_), .Y(_abc_934_new_n68_));
NAND3X1 NAND3X1_5 ( .A(_abc_934_new_n62_), .B(_abc_934_new_n72_), .C(_abc_934_new_n69_), .Y(_abc_934_new_n73_));
NAND3X1 NAND3X1_6 ( .A(state_4_), .B(_abc_934_new_n68_), .C(_abc_934_new_n73_), .Y(_abc_934_new_n74_));
NAND3X1 NAND3X1_7 ( .A(reset), .B(state_6_), .C(_abc_934_new_n94_), .Y(_abc_934_new_n95_));
NOR2X1 NOR2X1_1 ( .A(_auto_iopadmap_cc_368_execute_1033), .B(_abc_934_new_n88_), .Y(_abc_934_new_n119_));
NOR2X1 NOR2X1_10 ( .A(\codif[10] ), .B(\codif[11] ), .Y(_abc_934_new_n70_));
NOR2X1 NOR2X1_11 ( .A(\codif[8] ), .B(\codif[9] ), .Y(_abc_934_new_n71_));
NOR2X1 NOR2X1_12 ( .A(state_1_), .B(_abc_934_new_n50_), .Y(_abc_934_new_n76_));
NOR2X1 NOR2X1_13 ( .A(_auto_iopadmap_cc_368_execute_1033), .B(_abc_934_new_n50_), .Y(_abc_934_new_n94_));
NOR2X1 NOR2X1_14 ( .A(_abc_934_new_n97_), .B(_abc_934_new_n90_), .Y(_abc_801_auto_fsm_map_cc_170_map_fsm_238_4_));
NOR2X1 NOR2X1_15 ( .A(_abc_934_new_n97_), .B(_abc_934_new_n82_), .Y(_abc_801_auto_fsm_map_cc_170_map_fsm_238_5_));
NOR2X1 NOR2X1_16 ( .A(enable_pc_aux), .B(_abc_934_new_n100_), .Y(_auto_iopadmap_cc_368_execute_1039));
NOR2X1 NOR2X1_2 ( .A(state_2_), .B(state_4_), .Y(_abc_934_new_n123_));
NOR2X1 NOR2X1_3 ( .A(_abc_934_new_n49_), .B(_abc_934_new_n141_), .Y(_0en_mem_0_0_));
NOR2X1 NOR2X1_4 ( .A(_abc_934_new_n49_), .B(_abc_934_new_n100_), .Y(_0enable_pc_aux_0_0_));
NOR2X1 NOR2X1_5 ( .A(_abc_934_new_n49_), .B(_abc_934_new_n50_), .Y(_abc_934_new_n51_));
NOR2X1 NOR2X1_6 ( .A(\codif[2] ), .B(\codif[3] ), .Y(_abc_934_new_n54_));
NOR2X1 NOR2X1_7 ( .A(\codif[4] ), .B(\codif[6] ), .Y(_abc_934_new_n55_));
NOR2X1 NOR2X1_8 ( .A(_abc_934_new_n60_), .B(_abc_934_new_n61_), .Y(_abc_934_new_n62_));
NOR2X1 NOR2X1_9 ( .A(_abc_934_new_n65_), .B(_abc_934_new_n66_), .Y(_abc_934_new_n67_));
OAI21X1 OAI21X1_1 ( .A(_abc_934_new_n116_), .B(_abc_934_new_n117_), .C(_auto_iopadmap_cc_368_execute_1030_1_), .Y(_abc_934_new_n118_));
OAI21X1 OAI21X1_10 ( .A(_abc_934_new_n50_), .B(_abc_934_new_n106_), .C(_auto_iopadmap_cc_368_execute_1030_0_), .Y(_abc_934_new_n107_));
OAI21X1 OAI21X1_11 ( .A(state_3_), .B(state_5_), .C(_abc_934_new_n81_), .Y(_abc_934_new_n109_));
OAI21X1 OAI21X1_12 ( .A(done_mem), .B(_abc_934_new_n108_), .C(_auto_iopadmap_cc_368_execute_1033), .Y(_abc_934_new_n110_));
OAI21X1 OAI21X1_13 ( .A(\codif[5] ), .B(_abc_934_new_n103_), .C(_abc_934_new_n83_), .Y(_abc_934_new_n111_));
OAI21X1 OAI21X1_14 ( .A(state_0_), .B(_abc_934_new_n111_), .C(_abc_934_new_n110_), .Y(_abc_934_new_n112_));
OAI21X1 OAI21X1_15 ( .A(_abc_934_new_n108_), .B(_abc_934_new_n109_), .C(_abc_934_new_n112_), .Y(_abc_934_new_n113_));
OAI21X1 OAI21X1_2 ( .A(_abc_934_new_n50_), .B(_abc_934_new_n123_), .C(enable_pc_fsm), .Y(_abc_934_new_n124_));
OAI21X1 OAI21X1_3 ( .A(_abc_934_new_n50_), .B(_abc_934_new_n125_), .C(_abc_934_new_n124_), .Y(_abc_934_new_n126_));
OAI21X1 OAI21X1_4 ( .A(state_3_), .B(state_6_), .C(aligned_mem), .Y(_abc_934_new_n132_));
OAI21X1 OAI21X1_5 ( .A(_abc_934_new_n50_), .B(_abc_934_new_n123_), .C(_auto_iopadmap_cc_368_execute_1035), .Y(_abc_934_new_n137_));
OAI21X1 OAI21X1_6 ( .A(_abc_934_new_n50_), .B(_abc_934_new_n125_), .C(_abc_934_new_n137_), .Y(_abc_934_new_n138_));
OAI21X1 OAI21X1_7 ( .A(_abc_934_new_n80_), .B(_abc_934_new_n90_), .C(reset), .Y(_abc_934_new_n91_));
OAI21X1 OAI21X1_8 ( .A(_abc_934_new_n85_), .B(_abc_934_new_n87_), .C(_abc_934_new_n92_), .Y(_abc_801_auto_fsm_map_cc_170_map_fsm_238_0_));
OAI21X1 OAI21X1_9 ( .A(_abc_934_new_n56_), .B(_abc_934_new_n86_), .C(_abc_934_new_n95_), .Y(_abc_801_auto_fsm_map_cc_170_map_fsm_238_6_));
OAI22X1 OAI22X1_1 ( .A(\codif[5] ), .B(_abc_934_new_n95_), .C(_abc_934_new_n134_), .D(_abc_934_new_n133_), .Y(_0enable_exec_mem_0_0_));
OAI22X1 OAI22X1_2 ( .A(_auto_iopadmap_cc_368_execute_1033), .B(_abc_934_new_n88_), .C(_abc_934_new_n81_), .D(_abc_934_new_n83_), .Y(_abc_934_new_n89_));
OR2X2 OR2X2_1 ( .A(_abc_934_new_n111_), .B(state_3_), .Y(_abc_934_new_n131_));
OR2X2 OR2X2_2 ( .A(_abc_934_new_n86_), .B(_abc_934_new_n57_), .Y(_abc_934_new_n87_));
OR2X2 OR2X2_3 ( .A(state_3_), .B(state_5_), .Y(_abc_934_new_n102_));
OR2X2 OR2X2_4 ( .A(_abc_934_new_n104_), .B(_abc_934_new_n102_), .Y(_abc_934_new_n105_));


endmodule