module siphash(clk, reset_n, cs, we, \addr[0] , \addr[1] , \addr[2] , \addr[3] , \addr[4] , \addr[5] , \addr[6] , \addr[7] , \write_data[0] , \write_data[1] , \write_data[2] , \write_data[3] , \write_data[4] , \write_data[5] , \write_data[6] , \write_data[7] , \write_data[8] , \write_data[9] , \write_data[10] , \write_data[11] , \write_data[12] , \write_data[13] , \write_data[14] , \write_data[15] , \write_data[16] , \write_data[17] , \write_data[18] , \write_data[19] , \write_data[20] , \write_data[21] , \write_data[22] , \write_data[23] , \write_data[24] , \write_data[25] , \write_data[26] , \write_data[27] , \write_data[28] , \write_data[29] , \write_data[30] , \write_data[31] , \read_data[0] , \read_data[1] , \read_data[2] , \read_data[3] , \read_data[4] , \read_data[5] , \read_data[6] , \read_data[7] , \read_data[8] , \read_data[9] , \read_data[10] , \read_data[11] , \read_data[12] , \read_data[13] , \read_data[14] , \read_data[15] , \read_data[16] , \read_data[17] , \read_data[18] , \read_data[19] , \read_data[20] , \read_data[21] , \read_data[22] , \read_data[23] , \read_data[24] , \read_data[25] , \read_data[26] , \read_data[27] , \read_data[28] , \read_data[29] , \read_data[30] , \read_data[31] );

wire _0ctrl_reg_2_0__0_; 
wire _0ctrl_reg_2_0__1_; 
wire _0ctrl_reg_2_0__2_; 
wire _0key0_reg_31_0__0_; 
wire _0key0_reg_31_0__10_; 
wire _0key0_reg_31_0__11_; 
wire _0key0_reg_31_0__12_; 
wire _0key0_reg_31_0__13_; 
wire _0key0_reg_31_0__14_; 
wire _0key0_reg_31_0__15_; 
wire _0key0_reg_31_0__16_; 
wire _0key0_reg_31_0__17_; 
wire _0key0_reg_31_0__18_; 
wire _0key0_reg_31_0__19_; 
wire _0key0_reg_31_0__1_; 
wire _0key0_reg_31_0__20_; 
wire _0key0_reg_31_0__21_; 
wire _0key0_reg_31_0__22_; 
wire _0key0_reg_31_0__23_; 
wire _0key0_reg_31_0__24_; 
wire _0key0_reg_31_0__25_; 
wire _0key0_reg_31_0__26_; 
wire _0key0_reg_31_0__27_; 
wire _0key0_reg_31_0__28_; 
wire _0key0_reg_31_0__29_; 
wire _0key0_reg_31_0__2_; 
wire _0key0_reg_31_0__30_; 
wire _0key0_reg_31_0__31_; 
wire _0key0_reg_31_0__3_; 
wire _0key0_reg_31_0__4_; 
wire _0key0_reg_31_0__5_; 
wire _0key0_reg_31_0__6_; 
wire _0key0_reg_31_0__7_; 
wire _0key0_reg_31_0__8_; 
wire _0key0_reg_31_0__9_; 
wire _0key1_reg_31_0__0_; 
wire _0key1_reg_31_0__10_; 
wire _0key1_reg_31_0__11_; 
wire _0key1_reg_31_0__12_; 
wire _0key1_reg_31_0__13_; 
wire _0key1_reg_31_0__14_; 
wire _0key1_reg_31_0__15_; 
wire _0key1_reg_31_0__16_; 
wire _0key1_reg_31_0__17_; 
wire _0key1_reg_31_0__18_; 
wire _0key1_reg_31_0__19_; 
wire _0key1_reg_31_0__1_; 
wire _0key1_reg_31_0__20_; 
wire _0key1_reg_31_0__21_; 
wire _0key1_reg_31_0__22_; 
wire _0key1_reg_31_0__23_; 
wire _0key1_reg_31_0__24_; 
wire _0key1_reg_31_0__25_; 
wire _0key1_reg_31_0__26_; 
wire _0key1_reg_31_0__27_; 
wire _0key1_reg_31_0__28_; 
wire _0key1_reg_31_0__29_; 
wire _0key1_reg_31_0__2_; 
wire _0key1_reg_31_0__30_; 
wire _0key1_reg_31_0__31_; 
wire _0key1_reg_31_0__3_; 
wire _0key1_reg_31_0__4_; 
wire _0key1_reg_31_0__5_; 
wire _0key1_reg_31_0__6_; 
wire _0key1_reg_31_0__7_; 
wire _0key1_reg_31_0__8_; 
wire _0key1_reg_31_0__9_; 
wire _0key2_reg_31_0__0_; 
wire _0key2_reg_31_0__10_; 
wire _0key2_reg_31_0__11_; 
wire _0key2_reg_31_0__12_; 
wire _0key2_reg_31_0__13_; 
wire _0key2_reg_31_0__14_; 
wire _0key2_reg_31_0__15_; 
wire _0key2_reg_31_0__16_; 
wire _0key2_reg_31_0__17_; 
wire _0key2_reg_31_0__18_; 
wire _0key2_reg_31_0__19_; 
wire _0key2_reg_31_0__1_; 
wire _0key2_reg_31_0__20_; 
wire _0key2_reg_31_0__21_; 
wire _0key2_reg_31_0__22_; 
wire _0key2_reg_31_0__23_; 
wire _0key2_reg_31_0__24_; 
wire _0key2_reg_31_0__25_; 
wire _0key2_reg_31_0__26_; 
wire _0key2_reg_31_0__27_; 
wire _0key2_reg_31_0__28_; 
wire _0key2_reg_31_0__29_; 
wire _0key2_reg_31_0__2_; 
wire _0key2_reg_31_0__30_; 
wire _0key2_reg_31_0__31_; 
wire _0key2_reg_31_0__3_; 
wire _0key2_reg_31_0__4_; 
wire _0key2_reg_31_0__5_; 
wire _0key2_reg_31_0__6_; 
wire _0key2_reg_31_0__7_; 
wire _0key2_reg_31_0__8_; 
wire _0key2_reg_31_0__9_; 
wire _0key3_reg_31_0__0_; 
wire _0key3_reg_31_0__10_; 
wire _0key3_reg_31_0__11_; 
wire _0key3_reg_31_0__12_; 
wire _0key3_reg_31_0__13_; 
wire _0key3_reg_31_0__14_; 
wire _0key3_reg_31_0__15_; 
wire _0key3_reg_31_0__16_; 
wire _0key3_reg_31_0__17_; 
wire _0key3_reg_31_0__18_; 
wire _0key3_reg_31_0__19_; 
wire _0key3_reg_31_0__1_; 
wire _0key3_reg_31_0__20_; 
wire _0key3_reg_31_0__21_; 
wire _0key3_reg_31_0__22_; 
wire _0key3_reg_31_0__23_; 
wire _0key3_reg_31_0__24_; 
wire _0key3_reg_31_0__25_; 
wire _0key3_reg_31_0__26_; 
wire _0key3_reg_31_0__27_; 
wire _0key3_reg_31_0__28_; 
wire _0key3_reg_31_0__29_; 
wire _0key3_reg_31_0__2_; 
wire _0key3_reg_31_0__30_; 
wire _0key3_reg_31_0__31_; 
wire _0key3_reg_31_0__3_; 
wire _0key3_reg_31_0__4_; 
wire _0key3_reg_31_0__5_; 
wire _0key3_reg_31_0__6_; 
wire _0key3_reg_31_0__7_; 
wire _0key3_reg_31_0__8_; 
wire _0key3_reg_31_0__9_; 
wire _0long_reg_0_0_; 
wire _0mi0_reg_31_0__0_; 
wire _0mi0_reg_31_0__10_; 
wire _0mi0_reg_31_0__11_; 
wire _0mi0_reg_31_0__12_; 
wire _0mi0_reg_31_0__13_; 
wire _0mi0_reg_31_0__14_; 
wire _0mi0_reg_31_0__15_; 
wire _0mi0_reg_31_0__16_; 
wire _0mi0_reg_31_0__17_; 
wire _0mi0_reg_31_0__18_; 
wire _0mi0_reg_31_0__19_; 
wire _0mi0_reg_31_0__1_; 
wire _0mi0_reg_31_0__20_; 
wire _0mi0_reg_31_0__21_; 
wire _0mi0_reg_31_0__22_; 
wire _0mi0_reg_31_0__23_; 
wire _0mi0_reg_31_0__24_; 
wire _0mi0_reg_31_0__25_; 
wire _0mi0_reg_31_0__26_; 
wire _0mi0_reg_31_0__27_; 
wire _0mi0_reg_31_0__28_; 
wire _0mi0_reg_31_0__29_; 
wire _0mi0_reg_31_0__2_; 
wire _0mi0_reg_31_0__30_; 
wire _0mi0_reg_31_0__31_; 
wire _0mi0_reg_31_0__3_; 
wire _0mi0_reg_31_0__4_; 
wire _0mi0_reg_31_0__5_; 
wire _0mi0_reg_31_0__6_; 
wire _0mi0_reg_31_0__7_; 
wire _0mi0_reg_31_0__8_; 
wire _0mi0_reg_31_0__9_; 
wire _0mi1_reg_31_0__0_; 
wire _0mi1_reg_31_0__10_; 
wire _0mi1_reg_31_0__11_; 
wire _0mi1_reg_31_0__12_; 
wire _0mi1_reg_31_0__13_; 
wire _0mi1_reg_31_0__14_; 
wire _0mi1_reg_31_0__15_; 
wire _0mi1_reg_31_0__16_; 
wire _0mi1_reg_31_0__17_; 
wire _0mi1_reg_31_0__18_; 
wire _0mi1_reg_31_0__19_; 
wire _0mi1_reg_31_0__1_; 
wire _0mi1_reg_31_0__20_; 
wire _0mi1_reg_31_0__21_; 
wire _0mi1_reg_31_0__22_; 
wire _0mi1_reg_31_0__23_; 
wire _0mi1_reg_31_0__24_; 
wire _0mi1_reg_31_0__25_; 
wire _0mi1_reg_31_0__26_; 
wire _0mi1_reg_31_0__27_; 
wire _0mi1_reg_31_0__28_; 
wire _0mi1_reg_31_0__29_; 
wire _0mi1_reg_31_0__2_; 
wire _0mi1_reg_31_0__30_; 
wire _0mi1_reg_31_0__31_; 
wire _0mi1_reg_31_0__3_; 
wire _0mi1_reg_31_0__4_; 
wire _0mi1_reg_31_0__5_; 
wire _0mi1_reg_31_0__6_; 
wire _0mi1_reg_31_0__7_; 
wire _0mi1_reg_31_0__8_; 
wire _0mi1_reg_31_0__9_; 
wire _0param_reg_7_0__0_; 
wire _0param_reg_7_0__1_; 
wire _0param_reg_7_0__2_; 
wire _0param_reg_7_0__3_; 
wire _0param_reg_7_0__4_; 
wire _0param_reg_7_0__5_; 
wire _0param_reg_7_0__6_; 
wire _0param_reg_7_0__7_; 
wire _0word0_reg_31_0__0_; 
wire _0word0_reg_31_0__10_; 
wire _0word0_reg_31_0__11_; 
wire _0word0_reg_31_0__12_; 
wire _0word0_reg_31_0__13_; 
wire _0word0_reg_31_0__14_; 
wire _0word0_reg_31_0__15_; 
wire _0word0_reg_31_0__16_; 
wire _0word0_reg_31_0__17_; 
wire _0word0_reg_31_0__18_; 
wire _0word0_reg_31_0__19_; 
wire _0word0_reg_31_0__1_; 
wire _0word0_reg_31_0__20_; 
wire _0word0_reg_31_0__21_; 
wire _0word0_reg_31_0__22_; 
wire _0word0_reg_31_0__23_; 
wire _0word0_reg_31_0__24_; 
wire _0word0_reg_31_0__25_; 
wire _0word0_reg_31_0__26_; 
wire _0word0_reg_31_0__27_; 
wire _0word0_reg_31_0__28_; 
wire _0word0_reg_31_0__29_; 
wire _0word0_reg_31_0__2_; 
wire _0word0_reg_31_0__30_; 
wire _0word0_reg_31_0__31_; 
wire _0word0_reg_31_0__3_; 
wire _0word0_reg_31_0__4_; 
wire _0word0_reg_31_0__5_; 
wire _0word0_reg_31_0__6_; 
wire _0word0_reg_31_0__7_; 
wire _0word0_reg_31_0__8_; 
wire _0word0_reg_31_0__9_; 
wire _0word1_reg_31_0__0_; 
wire _0word1_reg_31_0__10_; 
wire _0word1_reg_31_0__11_; 
wire _0word1_reg_31_0__12_; 
wire _0word1_reg_31_0__13_; 
wire _0word1_reg_31_0__14_; 
wire _0word1_reg_31_0__15_; 
wire _0word1_reg_31_0__16_; 
wire _0word1_reg_31_0__17_; 
wire _0word1_reg_31_0__18_; 
wire _0word1_reg_31_0__19_; 
wire _0word1_reg_31_0__1_; 
wire _0word1_reg_31_0__20_; 
wire _0word1_reg_31_0__21_; 
wire _0word1_reg_31_0__22_; 
wire _0word1_reg_31_0__23_; 
wire _0word1_reg_31_0__24_; 
wire _0word1_reg_31_0__25_; 
wire _0word1_reg_31_0__26_; 
wire _0word1_reg_31_0__27_; 
wire _0word1_reg_31_0__28_; 
wire _0word1_reg_31_0__29_; 
wire _0word1_reg_31_0__2_; 
wire _0word1_reg_31_0__30_; 
wire _0word1_reg_31_0__31_; 
wire _0word1_reg_31_0__3_; 
wire _0word1_reg_31_0__4_; 
wire _0word1_reg_31_0__5_; 
wire _0word1_reg_31_0__6_; 
wire _0word1_reg_31_0__7_; 
wire _0word1_reg_31_0__8_; 
wire _0word1_reg_31_0__9_; 
wire _0word2_reg_31_0__0_; 
wire _0word2_reg_31_0__10_; 
wire _0word2_reg_31_0__11_; 
wire _0word2_reg_31_0__12_; 
wire _0word2_reg_31_0__13_; 
wire _0word2_reg_31_0__14_; 
wire _0word2_reg_31_0__15_; 
wire _0word2_reg_31_0__16_; 
wire _0word2_reg_31_0__17_; 
wire _0word2_reg_31_0__18_; 
wire _0word2_reg_31_0__19_; 
wire _0word2_reg_31_0__1_; 
wire _0word2_reg_31_0__20_; 
wire _0word2_reg_31_0__21_; 
wire _0word2_reg_31_0__22_; 
wire _0word2_reg_31_0__23_; 
wire _0word2_reg_31_0__24_; 
wire _0word2_reg_31_0__25_; 
wire _0word2_reg_31_0__26_; 
wire _0word2_reg_31_0__27_; 
wire _0word2_reg_31_0__28_; 
wire _0word2_reg_31_0__29_; 
wire _0word2_reg_31_0__2_; 
wire _0word2_reg_31_0__30_; 
wire _0word2_reg_31_0__31_; 
wire _0word2_reg_31_0__3_; 
wire _0word2_reg_31_0__4_; 
wire _0word2_reg_31_0__5_; 
wire _0word2_reg_31_0__6_; 
wire _0word2_reg_31_0__7_; 
wire _0word2_reg_31_0__8_; 
wire _0word2_reg_31_0__9_; 
wire _0word3_reg_31_0__0_; 
wire _0word3_reg_31_0__10_; 
wire _0word3_reg_31_0__11_; 
wire _0word3_reg_31_0__12_; 
wire _0word3_reg_31_0__13_; 
wire _0word3_reg_31_0__14_; 
wire _0word3_reg_31_0__15_; 
wire _0word3_reg_31_0__16_; 
wire _0word3_reg_31_0__17_; 
wire _0word3_reg_31_0__18_; 
wire _0word3_reg_31_0__19_; 
wire _0word3_reg_31_0__1_; 
wire _0word3_reg_31_0__20_; 
wire _0word3_reg_31_0__21_; 
wire _0word3_reg_31_0__22_; 
wire _0word3_reg_31_0__23_; 
wire _0word3_reg_31_0__24_; 
wire _0word3_reg_31_0__25_; 
wire _0word3_reg_31_0__26_; 
wire _0word3_reg_31_0__27_; 
wire _0word3_reg_31_0__28_; 
wire _0word3_reg_31_0__29_; 
wire _0word3_reg_31_0__2_; 
wire _0word3_reg_31_0__30_; 
wire _0word3_reg_31_0__31_; 
wire _0word3_reg_31_0__3_; 
wire _0word3_reg_31_0__4_; 
wire _0word3_reg_31_0__5_; 
wire _0word3_reg_31_0__6_; 
wire _0word3_reg_31_0__7_; 
wire _0word3_reg_31_0__8_; 
wire _0word3_reg_31_0__9_; 
wire _abc_19873_new_n1000_; 
wire _abc_19873_new_n1001_; 
wire _abc_19873_new_n1002_; 
wire _abc_19873_new_n1003_; 
wire _abc_19873_new_n1004_; 
wire _abc_19873_new_n1005_; 
wire _abc_19873_new_n1006_; 
wire _abc_19873_new_n1007_; 
wire _abc_19873_new_n1008_; 
wire _abc_19873_new_n1009_; 
wire _abc_19873_new_n1010_; 
wire _abc_19873_new_n1011_; 
wire _abc_19873_new_n1013_; 
wire _abc_19873_new_n1014_; 
wire _abc_19873_new_n1015_; 
wire _abc_19873_new_n1016_; 
wire _abc_19873_new_n1017_; 
wire _abc_19873_new_n1018_; 
wire _abc_19873_new_n1019_; 
wire _abc_19873_new_n1020_; 
wire _abc_19873_new_n1021_; 
wire _abc_19873_new_n1022_; 
wire _abc_19873_new_n1023_; 
wire _abc_19873_new_n1024_; 
wire _abc_19873_new_n1025_; 
wire _abc_19873_new_n1026_; 
wire _abc_19873_new_n1027_; 
wire _abc_19873_new_n1028_; 
wire _abc_19873_new_n1029_; 
wire _abc_19873_new_n1030_; 
wire _abc_19873_new_n1031_; 
wire _abc_19873_new_n1032_; 
wire _abc_19873_new_n1033_; 
wire _abc_19873_new_n1034_; 
wire _abc_19873_new_n1035_; 
wire _abc_19873_new_n1037_; 
wire _abc_19873_new_n1038_; 
wire _abc_19873_new_n1039_; 
wire _abc_19873_new_n1040_; 
wire _abc_19873_new_n1041_; 
wire _abc_19873_new_n1042_; 
wire _abc_19873_new_n1043_; 
wire _abc_19873_new_n1044_; 
wire _abc_19873_new_n1045_; 
wire _abc_19873_new_n1046_; 
wire _abc_19873_new_n1047_; 
wire _abc_19873_new_n1048_; 
wire _abc_19873_new_n1049_; 
wire _abc_19873_new_n1050_; 
wire _abc_19873_new_n1051_; 
wire _abc_19873_new_n1052_; 
wire _abc_19873_new_n1053_; 
wire _abc_19873_new_n1054_; 
wire _abc_19873_new_n1055_; 
wire _abc_19873_new_n1056_; 
wire _abc_19873_new_n1057_; 
wire _abc_19873_new_n1058_; 
wire _abc_19873_new_n1059_; 
wire _abc_19873_new_n1060_; 
wire _abc_19873_new_n1061_; 
wire _abc_19873_new_n1063_; 
wire _abc_19873_new_n1064_; 
wire _abc_19873_new_n1065_; 
wire _abc_19873_new_n1066_; 
wire _abc_19873_new_n1067_; 
wire _abc_19873_new_n1068_; 
wire _abc_19873_new_n1069_; 
wire _abc_19873_new_n1070_; 
wire _abc_19873_new_n1071_; 
wire _abc_19873_new_n1072_; 
wire _abc_19873_new_n1073_; 
wire _abc_19873_new_n1074_; 
wire _abc_19873_new_n1075_; 
wire _abc_19873_new_n1076_; 
wire _abc_19873_new_n1077_; 
wire _abc_19873_new_n1078_; 
wire _abc_19873_new_n1079_; 
wire _abc_19873_new_n1080_; 
wire _abc_19873_new_n1081_; 
wire _abc_19873_new_n1082_; 
wire _abc_19873_new_n1083_; 
wire _abc_19873_new_n1084_; 
wire _abc_19873_new_n1086_; 
wire _abc_19873_new_n1087_; 
wire _abc_19873_new_n1088_; 
wire _abc_19873_new_n1089_; 
wire _abc_19873_new_n1090_; 
wire _abc_19873_new_n1091_; 
wire _abc_19873_new_n1092_; 
wire _abc_19873_new_n1093_; 
wire _abc_19873_new_n1094_; 
wire _abc_19873_new_n1095_; 
wire _abc_19873_new_n1096_; 
wire _abc_19873_new_n1097_; 
wire _abc_19873_new_n1098_; 
wire _abc_19873_new_n1099_; 
wire _abc_19873_new_n1100_; 
wire _abc_19873_new_n1101_; 
wire _abc_19873_new_n1102_; 
wire _abc_19873_new_n1103_; 
wire _abc_19873_new_n1104_; 
wire _abc_19873_new_n1105_; 
wire _abc_19873_new_n1106_; 
wire _abc_19873_new_n1108_; 
wire _abc_19873_new_n1109_; 
wire _abc_19873_new_n1110_; 
wire _abc_19873_new_n1111_; 
wire _abc_19873_new_n1112_; 
wire _abc_19873_new_n1113_; 
wire _abc_19873_new_n1114_; 
wire _abc_19873_new_n1115_; 
wire _abc_19873_new_n1116_; 
wire _abc_19873_new_n1117_; 
wire _abc_19873_new_n1118_; 
wire _abc_19873_new_n1119_; 
wire _abc_19873_new_n1120_; 
wire _abc_19873_new_n1121_; 
wire _abc_19873_new_n1122_; 
wire _abc_19873_new_n1123_; 
wire _abc_19873_new_n1124_; 
wire _abc_19873_new_n1125_; 
wire _abc_19873_new_n1126_; 
wire _abc_19873_new_n1128_; 
wire _abc_19873_new_n1129_; 
wire _abc_19873_new_n1130_; 
wire _abc_19873_new_n1131_; 
wire _abc_19873_new_n1132_; 
wire _abc_19873_new_n1133_; 
wire _abc_19873_new_n1134_; 
wire _abc_19873_new_n1135_; 
wire _abc_19873_new_n1136_; 
wire _abc_19873_new_n1137_; 
wire _abc_19873_new_n1138_; 
wire _abc_19873_new_n1139_; 
wire _abc_19873_new_n1140_; 
wire _abc_19873_new_n1141_; 
wire _abc_19873_new_n1142_; 
wire _abc_19873_new_n1143_; 
wire _abc_19873_new_n1144_; 
wire _abc_19873_new_n1145_; 
wire _abc_19873_new_n1146_; 
wire _abc_19873_new_n1148_; 
wire _abc_19873_new_n1149_; 
wire _abc_19873_new_n1150_; 
wire _abc_19873_new_n1151_; 
wire _abc_19873_new_n1152_; 
wire _abc_19873_new_n1153_; 
wire _abc_19873_new_n1154_; 
wire _abc_19873_new_n1155_; 
wire _abc_19873_new_n1156_; 
wire _abc_19873_new_n1157_; 
wire _abc_19873_new_n1158_; 
wire _abc_19873_new_n1159_; 
wire _abc_19873_new_n1160_; 
wire _abc_19873_new_n1161_; 
wire _abc_19873_new_n1162_; 
wire _abc_19873_new_n1163_; 
wire _abc_19873_new_n1164_; 
wire _abc_19873_new_n1165_; 
wire _abc_19873_new_n1166_; 
wire _abc_19873_new_n1168_; 
wire _abc_19873_new_n1169_; 
wire _abc_19873_new_n1170_; 
wire _abc_19873_new_n1171_; 
wire _abc_19873_new_n1172_; 
wire _abc_19873_new_n1173_; 
wire _abc_19873_new_n1174_; 
wire _abc_19873_new_n1175_; 
wire _abc_19873_new_n1176_; 
wire _abc_19873_new_n1177_; 
wire _abc_19873_new_n1178_; 
wire _abc_19873_new_n1179_; 
wire _abc_19873_new_n1180_; 
wire _abc_19873_new_n1181_; 
wire _abc_19873_new_n1182_; 
wire _abc_19873_new_n1183_; 
wire _abc_19873_new_n1184_; 
wire _abc_19873_new_n1185_; 
wire _abc_19873_new_n1186_; 
wire _abc_19873_new_n1187_; 
wire _abc_19873_new_n1189_; 
wire _abc_19873_new_n1190_; 
wire _abc_19873_new_n1191_; 
wire _abc_19873_new_n1192_; 
wire _abc_19873_new_n1193_; 
wire _abc_19873_new_n1194_; 
wire _abc_19873_new_n1195_; 
wire _abc_19873_new_n1196_; 
wire _abc_19873_new_n1197_; 
wire _abc_19873_new_n1198_; 
wire _abc_19873_new_n1199_; 
wire _abc_19873_new_n1200_; 
wire _abc_19873_new_n1201_; 
wire _abc_19873_new_n1202_; 
wire _abc_19873_new_n1203_; 
wire _abc_19873_new_n1204_; 
wire _abc_19873_new_n1205_; 
wire _abc_19873_new_n1206_; 
wire _abc_19873_new_n1207_; 
wire _abc_19873_new_n1208_; 
wire _abc_19873_new_n1209_; 
wire _abc_19873_new_n1211_; 
wire _abc_19873_new_n1212_; 
wire _abc_19873_new_n1213_; 
wire _abc_19873_new_n1214_; 
wire _abc_19873_new_n1215_; 
wire _abc_19873_new_n1216_; 
wire _abc_19873_new_n1217_; 
wire _abc_19873_new_n1218_; 
wire _abc_19873_new_n1219_; 
wire _abc_19873_new_n1220_; 
wire _abc_19873_new_n1221_; 
wire _abc_19873_new_n1222_; 
wire _abc_19873_new_n1223_; 
wire _abc_19873_new_n1224_; 
wire _abc_19873_new_n1225_; 
wire _abc_19873_new_n1226_; 
wire _abc_19873_new_n1227_; 
wire _abc_19873_new_n1228_; 
wire _abc_19873_new_n1229_; 
wire _abc_19873_new_n1230_; 
wire _abc_19873_new_n1232_; 
wire _abc_19873_new_n1233_; 
wire _abc_19873_new_n1234_; 
wire _abc_19873_new_n1235_; 
wire _abc_19873_new_n1236_; 
wire _abc_19873_new_n1237_; 
wire _abc_19873_new_n1238_; 
wire _abc_19873_new_n1239_; 
wire _abc_19873_new_n1240_; 
wire _abc_19873_new_n1241_; 
wire _abc_19873_new_n1242_; 
wire _abc_19873_new_n1243_; 
wire _abc_19873_new_n1244_; 
wire _abc_19873_new_n1245_; 
wire _abc_19873_new_n1246_; 
wire _abc_19873_new_n1247_; 
wire _abc_19873_new_n1248_; 
wire _abc_19873_new_n1249_; 
wire _abc_19873_new_n1250_; 
wire _abc_19873_new_n1251_; 
wire _abc_19873_new_n1253_; 
wire _abc_19873_new_n1254_; 
wire _abc_19873_new_n1255_; 
wire _abc_19873_new_n1256_; 
wire _abc_19873_new_n1257_; 
wire _abc_19873_new_n1258_; 
wire _abc_19873_new_n1259_; 
wire _abc_19873_new_n1260_; 
wire _abc_19873_new_n1261_; 
wire _abc_19873_new_n1262_; 
wire _abc_19873_new_n1263_; 
wire _abc_19873_new_n1264_; 
wire _abc_19873_new_n1265_; 
wire _abc_19873_new_n1266_; 
wire _abc_19873_new_n1267_; 
wire _abc_19873_new_n1268_; 
wire _abc_19873_new_n1269_; 
wire _abc_19873_new_n1270_; 
wire _abc_19873_new_n1271_; 
wire _abc_19873_new_n1273_; 
wire _abc_19873_new_n1274_; 
wire _abc_19873_new_n1275_; 
wire _abc_19873_new_n1276_; 
wire _abc_19873_new_n1277_; 
wire _abc_19873_new_n1278_; 
wire _abc_19873_new_n1279_; 
wire _abc_19873_new_n1280_; 
wire _abc_19873_new_n1281_; 
wire _abc_19873_new_n1282_; 
wire _abc_19873_new_n1283_; 
wire _abc_19873_new_n1284_; 
wire _abc_19873_new_n1285_; 
wire _abc_19873_new_n1286_; 
wire _abc_19873_new_n1287_; 
wire _abc_19873_new_n1288_; 
wire _abc_19873_new_n1289_; 
wire _abc_19873_new_n1290_; 
wire _abc_19873_new_n1291_; 
wire _abc_19873_new_n1292_; 
wire _abc_19873_new_n1294_; 
wire _abc_19873_new_n1295_; 
wire _abc_19873_new_n1296_; 
wire _abc_19873_new_n1297_; 
wire _abc_19873_new_n1298_; 
wire _abc_19873_new_n1299_; 
wire _abc_19873_new_n1300_; 
wire _abc_19873_new_n1301_; 
wire _abc_19873_new_n1302_; 
wire _abc_19873_new_n1303_; 
wire _abc_19873_new_n1304_; 
wire _abc_19873_new_n1305_; 
wire _abc_19873_new_n1306_; 
wire _abc_19873_new_n1307_; 
wire _abc_19873_new_n1308_; 
wire _abc_19873_new_n1309_; 
wire _abc_19873_new_n1310_; 
wire _abc_19873_new_n1311_; 
wire _abc_19873_new_n1312_; 
wire _abc_19873_new_n1313_; 
wire _abc_19873_new_n1314_; 
wire _abc_19873_new_n1316_; 
wire _abc_19873_new_n1317_; 
wire _abc_19873_new_n1318_; 
wire _abc_19873_new_n1319_; 
wire _abc_19873_new_n1320_; 
wire _abc_19873_new_n1321_; 
wire _abc_19873_new_n1322_; 
wire _abc_19873_new_n1323_; 
wire _abc_19873_new_n1324_; 
wire _abc_19873_new_n1325_; 
wire _abc_19873_new_n1326_; 
wire _abc_19873_new_n1327_; 
wire _abc_19873_new_n1328_; 
wire _abc_19873_new_n1329_; 
wire _abc_19873_new_n1330_; 
wire _abc_19873_new_n1331_; 
wire _abc_19873_new_n1332_; 
wire _abc_19873_new_n1333_; 
wire _abc_19873_new_n1334_; 
wire _abc_19873_new_n1335_; 
wire _abc_19873_new_n1337_; 
wire _abc_19873_new_n1338_; 
wire _abc_19873_new_n1339_; 
wire _abc_19873_new_n1340_; 
wire _abc_19873_new_n1341_; 
wire _abc_19873_new_n1342_; 
wire _abc_19873_new_n1343_; 
wire _abc_19873_new_n1344_; 
wire _abc_19873_new_n1345_; 
wire _abc_19873_new_n1346_; 
wire _abc_19873_new_n1347_; 
wire _abc_19873_new_n1348_; 
wire _abc_19873_new_n1349_; 
wire _abc_19873_new_n1350_; 
wire _abc_19873_new_n1351_; 
wire _abc_19873_new_n1352_; 
wire _abc_19873_new_n1353_; 
wire _abc_19873_new_n1354_; 
wire _abc_19873_new_n1355_; 
wire _abc_19873_new_n1356_; 
wire _abc_19873_new_n1358_; 
wire _abc_19873_new_n1359_; 
wire _abc_19873_new_n1360_; 
wire _abc_19873_new_n1361_; 
wire _abc_19873_new_n1362_; 
wire _abc_19873_new_n1363_; 
wire _abc_19873_new_n1364_; 
wire _abc_19873_new_n1365_; 
wire _abc_19873_new_n1366_; 
wire _abc_19873_new_n1367_; 
wire _abc_19873_new_n1368_; 
wire _abc_19873_new_n1369_; 
wire _abc_19873_new_n1370_; 
wire _abc_19873_new_n1371_; 
wire _abc_19873_new_n1372_; 
wire _abc_19873_new_n1373_; 
wire _abc_19873_new_n1374_; 
wire _abc_19873_new_n1375_; 
wire _abc_19873_new_n1376_; 
wire _abc_19873_new_n1377_; 
wire _abc_19873_new_n1379_; 
wire _abc_19873_new_n1380_; 
wire _abc_19873_new_n1381_; 
wire _abc_19873_new_n1382_; 
wire _abc_19873_new_n1383_; 
wire _abc_19873_new_n1384_; 
wire _abc_19873_new_n1385_; 
wire _abc_19873_new_n1386_; 
wire _abc_19873_new_n1387_; 
wire _abc_19873_new_n1388_; 
wire _abc_19873_new_n1389_; 
wire _abc_19873_new_n1390_; 
wire _abc_19873_new_n1391_; 
wire _abc_19873_new_n1392_; 
wire _abc_19873_new_n1393_; 
wire _abc_19873_new_n1394_; 
wire _abc_19873_new_n1395_; 
wire _abc_19873_new_n1396_; 
wire _abc_19873_new_n1397_; 
wire _abc_19873_new_n1398_; 
wire _abc_19873_new_n1400_; 
wire _abc_19873_new_n1401_; 
wire _abc_19873_new_n1402_; 
wire _abc_19873_new_n1403_; 
wire _abc_19873_new_n1404_; 
wire _abc_19873_new_n1405_; 
wire _abc_19873_new_n1406_; 
wire _abc_19873_new_n1407_; 
wire _abc_19873_new_n1408_; 
wire _abc_19873_new_n1409_; 
wire _abc_19873_new_n1410_; 
wire _abc_19873_new_n1411_; 
wire _abc_19873_new_n1412_; 
wire _abc_19873_new_n1413_; 
wire _abc_19873_new_n1414_; 
wire _abc_19873_new_n1415_; 
wire _abc_19873_new_n1416_; 
wire _abc_19873_new_n1417_; 
wire _abc_19873_new_n1418_; 
wire _abc_19873_new_n1419_; 
wire _abc_19873_new_n1421_; 
wire _abc_19873_new_n1422_; 
wire _abc_19873_new_n1423_; 
wire _abc_19873_new_n1424_; 
wire _abc_19873_new_n1425_; 
wire _abc_19873_new_n1426_; 
wire _abc_19873_new_n1427_; 
wire _abc_19873_new_n1428_; 
wire _abc_19873_new_n1429_; 
wire _abc_19873_new_n1430_; 
wire _abc_19873_new_n1431_; 
wire _abc_19873_new_n1432_; 
wire _abc_19873_new_n1433_; 
wire _abc_19873_new_n1434_; 
wire _abc_19873_new_n1435_; 
wire _abc_19873_new_n1436_; 
wire _abc_19873_new_n1437_; 
wire _abc_19873_new_n1438_; 
wire _abc_19873_new_n1439_; 
wire _abc_19873_new_n1441_; 
wire _abc_19873_new_n1442_; 
wire _abc_19873_new_n1443_; 
wire _abc_19873_new_n1444_; 
wire _abc_19873_new_n1445_; 
wire _abc_19873_new_n1446_; 
wire _abc_19873_new_n1447_; 
wire _abc_19873_new_n1448_; 
wire _abc_19873_new_n1449_; 
wire _abc_19873_new_n1450_; 
wire _abc_19873_new_n1451_; 
wire _abc_19873_new_n1452_; 
wire _abc_19873_new_n1453_; 
wire _abc_19873_new_n1454_; 
wire _abc_19873_new_n1455_; 
wire _abc_19873_new_n1456_; 
wire _abc_19873_new_n1457_; 
wire _abc_19873_new_n1458_; 
wire _abc_19873_new_n1459_; 
wire _abc_19873_new_n1460_; 
wire _abc_19873_new_n1462_; 
wire _abc_19873_new_n1463_; 
wire _abc_19873_new_n1464_; 
wire _abc_19873_new_n1465_; 
wire _abc_19873_new_n1466_; 
wire _abc_19873_new_n1467_; 
wire _abc_19873_new_n1468_; 
wire _abc_19873_new_n1469_; 
wire _abc_19873_new_n1470_; 
wire _abc_19873_new_n1471_; 
wire _abc_19873_new_n1472_; 
wire _abc_19873_new_n1473_; 
wire _abc_19873_new_n1474_; 
wire _abc_19873_new_n1475_; 
wire _abc_19873_new_n1476_; 
wire _abc_19873_new_n1477_; 
wire _abc_19873_new_n1478_; 
wire _abc_19873_new_n1479_; 
wire _abc_19873_new_n1480_; 
wire _abc_19873_new_n1481_; 
wire _abc_19873_new_n1483_; 
wire _abc_19873_new_n1484_; 
wire _abc_19873_new_n1485_; 
wire _abc_19873_new_n1486_; 
wire _abc_19873_new_n1487_; 
wire _abc_19873_new_n1488_; 
wire _abc_19873_new_n1489_; 
wire _abc_19873_new_n1490_; 
wire _abc_19873_new_n1491_; 
wire _abc_19873_new_n1492_; 
wire _abc_19873_new_n1493_; 
wire _abc_19873_new_n1494_; 
wire _abc_19873_new_n1495_; 
wire _abc_19873_new_n1496_; 
wire _abc_19873_new_n1497_; 
wire _abc_19873_new_n1498_; 
wire _abc_19873_new_n1499_; 
wire _abc_19873_new_n1500_; 
wire _abc_19873_new_n1501_; 
wire _abc_19873_new_n1503_; 
wire _abc_19873_new_n1504_; 
wire _abc_19873_new_n1505_; 
wire _abc_19873_new_n1506_; 
wire _abc_19873_new_n1507_; 
wire _abc_19873_new_n1508_; 
wire _abc_19873_new_n1509_; 
wire _abc_19873_new_n1510_; 
wire _abc_19873_new_n1511_; 
wire _abc_19873_new_n1512_; 
wire _abc_19873_new_n1513_; 
wire _abc_19873_new_n1514_; 
wire _abc_19873_new_n1515_; 
wire _abc_19873_new_n1516_; 
wire _abc_19873_new_n1517_; 
wire _abc_19873_new_n1518_; 
wire _abc_19873_new_n1519_; 
wire _abc_19873_new_n1520_; 
wire _abc_19873_new_n1521_; 
wire _abc_19873_new_n1523_; 
wire _abc_19873_new_n1524_; 
wire _abc_19873_new_n1525_; 
wire _abc_19873_new_n1526_; 
wire _abc_19873_new_n1527_; 
wire _abc_19873_new_n1528_; 
wire _abc_19873_new_n1529_; 
wire _abc_19873_new_n1530_; 
wire _abc_19873_new_n1531_; 
wire _abc_19873_new_n1532_; 
wire _abc_19873_new_n1533_; 
wire _abc_19873_new_n1534_; 
wire _abc_19873_new_n1535_; 
wire _abc_19873_new_n1536_; 
wire _abc_19873_new_n1537_; 
wire _abc_19873_new_n1538_; 
wire _abc_19873_new_n1539_; 
wire _abc_19873_new_n1540_; 
wire _abc_19873_new_n1541_; 
wire _abc_19873_new_n1542_; 
wire _abc_19873_new_n1544_; 
wire _abc_19873_new_n1545_; 
wire _abc_19873_new_n1546_; 
wire _abc_19873_new_n1547_; 
wire _abc_19873_new_n1548_; 
wire _abc_19873_new_n1549_; 
wire _abc_19873_new_n1550_; 
wire _abc_19873_new_n1551_; 
wire _abc_19873_new_n1552_; 
wire _abc_19873_new_n1553_; 
wire _abc_19873_new_n1554_; 
wire _abc_19873_new_n1555_; 
wire _abc_19873_new_n1556_; 
wire _abc_19873_new_n1557_; 
wire _abc_19873_new_n1558_; 
wire _abc_19873_new_n1559_; 
wire _abc_19873_new_n1560_; 
wire _abc_19873_new_n1561_; 
wire _abc_19873_new_n1562_; 
wire _abc_19873_new_n1563_; 
wire _abc_19873_new_n1565_; 
wire _abc_19873_new_n1566_; 
wire _abc_19873_new_n1567_; 
wire _abc_19873_new_n1568_; 
wire _abc_19873_new_n1569_; 
wire _abc_19873_new_n1570_; 
wire _abc_19873_new_n1571_; 
wire _abc_19873_new_n1572_; 
wire _abc_19873_new_n1573_; 
wire _abc_19873_new_n1574_; 
wire _abc_19873_new_n1575_; 
wire _abc_19873_new_n1576_; 
wire _abc_19873_new_n1577_; 
wire _abc_19873_new_n1578_; 
wire _abc_19873_new_n1579_; 
wire _abc_19873_new_n1580_; 
wire _abc_19873_new_n1581_; 
wire _abc_19873_new_n1582_; 
wire _abc_19873_new_n1583_; 
wire _abc_19873_new_n1584_; 
wire _abc_19873_new_n1586_; 
wire _abc_19873_new_n1587_; 
wire _abc_19873_new_n1588_; 
wire _abc_19873_new_n1589_; 
wire _abc_19873_new_n1590_; 
wire _abc_19873_new_n1591_; 
wire _abc_19873_new_n1592_; 
wire _abc_19873_new_n1593_; 
wire _abc_19873_new_n1594_; 
wire _abc_19873_new_n1595_; 
wire _abc_19873_new_n1596_; 
wire _abc_19873_new_n1597_; 
wire _abc_19873_new_n1598_; 
wire _abc_19873_new_n1599_; 
wire _abc_19873_new_n1600_; 
wire _abc_19873_new_n1601_; 
wire _abc_19873_new_n1602_; 
wire _abc_19873_new_n1603_; 
wire _abc_19873_new_n1604_; 
wire _abc_19873_new_n1606_; 
wire _abc_19873_new_n1607_; 
wire _abc_19873_new_n1608_; 
wire _abc_19873_new_n1609_; 
wire _abc_19873_new_n1611_; 
wire _abc_19873_new_n1612_; 
wire _abc_19873_new_n1613_; 
wire _abc_19873_new_n1615_; 
wire _abc_19873_new_n1616_; 
wire _abc_19873_new_n1617_; 
wire _abc_19873_new_n1619_; 
wire _abc_19873_new_n1620_; 
wire _abc_19873_new_n1621_; 
wire _abc_19873_new_n1623_; 
wire _abc_19873_new_n1624_; 
wire _abc_19873_new_n1625_; 
wire _abc_19873_new_n1627_; 
wire _abc_19873_new_n1628_; 
wire _abc_19873_new_n1629_; 
wire _abc_19873_new_n1631_; 
wire _abc_19873_new_n1632_; 
wire _abc_19873_new_n1633_; 
wire _abc_19873_new_n1635_; 
wire _abc_19873_new_n1636_; 
wire _abc_19873_new_n1637_; 
wire _abc_19873_new_n1639_; 
wire _abc_19873_new_n1640_; 
wire _abc_19873_new_n1641_; 
wire _abc_19873_new_n1643_; 
wire _abc_19873_new_n1644_; 
wire _abc_19873_new_n1645_; 
wire _abc_19873_new_n1647_; 
wire _abc_19873_new_n1648_; 
wire _abc_19873_new_n1649_; 
wire _abc_19873_new_n1651_; 
wire _abc_19873_new_n1652_; 
wire _abc_19873_new_n1653_; 
wire _abc_19873_new_n1655_; 
wire _abc_19873_new_n1656_; 
wire _abc_19873_new_n1657_; 
wire _abc_19873_new_n1659_; 
wire _abc_19873_new_n1660_; 
wire _abc_19873_new_n1661_; 
wire _abc_19873_new_n1663_; 
wire _abc_19873_new_n1664_; 
wire _abc_19873_new_n1665_; 
wire _abc_19873_new_n1667_; 
wire _abc_19873_new_n1668_; 
wire _abc_19873_new_n1669_; 
wire _abc_19873_new_n1671_; 
wire _abc_19873_new_n1672_; 
wire _abc_19873_new_n1673_; 
wire _abc_19873_new_n1675_; 
wire _abc_19873_new_n1676_; 
wire _abc_19873_new_n1677_; 
wire _abc_19873_new_n1679_; 
wire _abc_19873_new_n1680_; 
wire _abc_19873_new_n1681_; 
wire _abc_19873_new_n1683_; 
wire _abc_19873_new_n1684_; 
wire _abc_19873_new_n1685_; 
wire _abc_19873_new_n1687_; 
wire _abc_19873_new_n1688_; 
wire _abc_19873_new_n1689_; 
wire _abc_19873_new_n1691_; 
wire _abc_19873_new_n1692_; 
wire _abc_19873_new_n1693_; 
wire _abc_19873_new_n1695_; 
wire _abc_19873_new_n1696_; 
wire _abc_19873_new_n1697_; 
wire _abc_19873_new_n1699_; 
wire _abc_19873_new_n1700_; 
wire _abc_19873_new_n1701_; 
wire _abc_19873_new_n1703_; 
wire _abc_19873_new_n1704_; 
wire _abc_19873_new_n1705_; 
wire _abc_19873_new_n1707_; 
wire _abc_19873_new_n1708_; 
wire _abc_19873_new_n1709_; 
wire _abc_19873_new_n1711_; 
wire _abc_19873_new_n1712_; 
wire _abc_19873_new_n1713_; 
wire _abc_19873_new_n1715_; 
wire _abc_19873_new_n1716_; 
wire _abc_19873_new_n1717_; 
wire _abc_19873_new_n1719_; 
wire _abc_19873_new_n1720_; 
wire _abc_19873_new_n1721_; 
wire _abc_19873_new_n1723_; 
wire _abc_19873_new_n1724_; 
wire _abc_19873_new_n1725_; 
wire _abc_19873_new_n1727_; 
wire _abc_19873_new_n1728_; 
wire _abc_19873_new_n1729_; 
wire _abc_19873_new_n1731_; 
wire _abc_19873_new_n1732_; 
wire _abc_19873_new_n1733_; 
wire _abc_19873_new_n1735_; 
wire _abc_19873_new_n1736_; 
wire _abc_19873_new_n1737_; 
wire _abc_19873_new_n1739_; 
wire _abc_19873_new_n1740_; 
wire _abc_19873_new_n1741_; 
wire _abc_19873_new_n1743_; 
wire _abc_19873_new_n1744_; 
wire _abc_19873_new_n1745_; 
wire _abc_19873_new_n1747_; 
wire _abc_19873_new_n1748_; 
wire _abc_19873_new_n1749_; 
wire _abc_19873_new_n1751_; 
wire _abc_19873_new_n1752_; 
wire _abc_19873_new_n1753_; 
wire _abc_19873_new_n1755_; 
wire _abc_19873_new_n1756_; 
wire _abc_19873_new_n1757_; 
wire _abc_19873_new_n1759_; 
wire _abc_19873_new_n1760_; 
wire _abc_19873_new_n1761_; 
wire _abc_19873_new_n1763_; 
wire _abc_19873_new_n1764_; 
wire _abc_19873_new_n1765_; 
wire _abc_19873_new_n1767_; 
wire _abc_19873_new_n1768_; 
wire _abc_19873_new_n1769_; 
wire _abc_19873_new_n1771_; 
wire _abc_19873_new_n1772_; 
wire _abc_19873_new_n1773_; 
wire _abc_19873_new_n1775_; 
wire _abc_19873_new_n1776_; 
wire _abc_19873_new_n1777_; 
wire _abc_19873_new_n1779_; 
wire _abc_19873_new_n1780_; 
wire _abc_19873_new_n1781_; 
wire _abc_19873_new_n1783_; 
wire _abc_19873_new_n1784_; 
wire _abc_19873_new_n1785_; 
wire _abc_19873_new_n1787_; 
wire _abc_19873_new_n1788_; 
wire _abc_19873_new_n1789_; 
wire _abc_19873_new_n1791_; 
wire _abc_19873_new_n1792_; 
wire _abc_19873_new_n1793_; 
wire _abc_19873_new_n1795_; 
wire _abc_19873_new_n1796_; 
wire _abc_19873_new_n1797_; 
wire _abc_19873_new_n1799_; 
wire _abc_19873_new_n1800_; 
wire _abc_19873_new_n1801_; 
wire _abc_19873_new_n1803_; 
wire _abc_19873_new_n1804_; 
wire _abc_19873_new_n1805_; 
wire _abc_19873_new_n1807_; 
wire _abc_19873_new_n1808_; 
wire _abc_19873_new_n1809_; 
wire _abc_19873_new_n1811_; 
wire _abc_19873_new_n1812_; 
wire _abc_19873_new_n1813_; 
wire _abc_19873_new_n1815_; 
wire _abc_19873_new_n1816_; 
wire _abc_19873_new_n1817_; 
wire _abc_19873_new_n1819_; 
wire _abc_19873_new_n1820_; 
wire _abc_19873_new_n1821_; 
wire _abc_19873_new_n1823_; 
wire _abc_19873_new_n1824_; 
wire _abc_19873_new_n1825_; 
wire _abc_19873_new_n1827_; 
wire _abc_19873_new_n1828_; 
wire _abc_19873_new_n1829_; 
wire _abc_19873_new_n1831_; 
wire _abc_19873_new_n1832_; 
wire _abc_19873_new_n1833_; 
wire _abc_19873_new_n1835_; 
wire _abc_19873_new_n1836_; 
wire _abc_19873_new_n1837_; 
wire _abc_19873_new_n1839_; 
wire _abc_19873_new_n1840_; 
wire _abc_19873_new_n1841_; 
wire _abc_19873_new_n1843_; 
wire _abc_19873_new_n1844_; 
wire _abc_19873_new_n1845_; 
wire _abc_19873_new_n1847_; 
wire _abc_19873_new_n1848_; 
wire _abc_19873_new_n1849_; 
wire _abc_19873_new_n1851_; 
wire _abc_19873_new_n1852_; 
wire _abc_19873_new_n1853_; 
wire _abc_19873_new_n1855_; 
wire _abc_19873_new_n1856_; 
wire _abc_19873_new_n1857_; 
wire _abc_19873_new_n1859_; 
wire _abc_19873_new_n1860_; 
wire _abc_19873_new_n1861_; 
wire _abc_19873_new_n1863_; 
wire _abc_19873_new_n1864_; 
wire _abc_19873_new_n1865_; 
wire _abc_19873_new_n1867_; 
wire _abc_19873_new_n1868_; 
wire _abc_19873_new_n1869_; 
wire _abc_19873_new_n1871_; 
wire _abc_19873_new_n1872_; 
wire _abc_19873_new_n1873_; 
wire _abc_19873_new_n1875_; 
wire _abc_19873_new_n1876_; 
wire _abc_19873_new_n1877_; 
wire _abc_19873_new_n1879_; 
wire _abc_19873_new_n1880_; 
wire _abc_19873_new_n1881_; 
wire _abc_19873_new_n1883_; 
wire _abc_19873_new_n1884_; 
wire _abc_19873_new_n1885_; 
wire _abc_19873_new_n1887_; 
wire _abc_19873_new_n1888_; 
wire _abc_19873_new_n1889_; 
wire _abc_19873_new_n1891_; 
wire _abc_19873_new_n1892_; 
wire _abc_19873_new_n1893_; 
wire _abc_19873_new_n1895_; 
wire _abc_19873_new_n1896_; 
wire _abc_19873_new_n1897_; 
wire _abc_19873_new_n1899_; 
wire _abc_19873_new_n1900_; 
wire _abc_19873_new_n1901_; 
wire _abc_19873_new_n1903_; 
wire _abc_19873_new_n1904_; 
wire _abc_19873_new_n1905_; 
wire _abc_19873_new_n1907_; 
wire _abc_19873_new_n1908_; 
wire _abc_19873_new_n1909_; 
wire _abc_19873_new_n1911_; 
wire _abc_19873_new_n1912_; 
wire _abc_19873_new_n1913_; 
wire _abc_19873_new_n1915_; 
wire _abc_19873_new_n1916_; 
wire _abc_19873_new_n1917_; 
wire _abc_19873_new_n1919_; 
wire _abc_19873_new_n1920_; 
wire _abc_19873_new_n1921_; 
wire _abc_19873_new_n1923_; 
wire _abc_19873_new_n1924_; 
wire _abc_19873_new_n1925_; 
wire _abc_19873_new_n1927_; 
wire _abc_19873_new_n1928_; 
wire _abc_19873_new_n1929_; 
wire _abc_19873_new_n1931_; 
wire _abc_19873_new_n1932_; 
wire _abc_19873_new_n1933_; 
wire _abc_19873_new_n1935_; 
wire _abc_19873_new_n1936_; 
wire _abc_19873_new_n1937_; 
wire _abc_19873_new_n1939_; 
wire _abc_19873_new_n1940_; 
wire _abc_19873_new_n1941_; 
wire _abc_19873_new_n1943_; 
wire _abc_19873_new_n1944_; 
wire _abc_19873_new_n1945_; 
wire _abc_19873_new_n1947_; 
wire _abc_19873_new_n1948_; 
wire _abc_19873_new_n1949_; 
wire _abc_19873_new_n1951_; 
wire _abc_19873_new_n1952_; 
wire _abc_19873_new_n1953_; 
wire _abc_19873_new_n1955_; 
wire _abc_19873_new_n1956_; 
wire _abc_19873_new_n1957_; 
wire _abc_19873_new_n1959_; 
wire _abc_19873_new_n1960_; 
wire _abc_19873_new_n1961_; 
wire _abc_19873_new_n1963_; 
wire _abc_19873_new_n1964_; 
wire _abc_19873_new_n1965_; 
wire _abc_19873_new_n1967_; 
wire _abc_19873_new_n1968_; 
wire _abc_19873_new_n1969_; 
wire _abc_19873_new_n1971_; 
wire _abc_19873_new_n1972_; 
wire _abc_19873_new_n1973_; 
wire _abc_19873_new_n1975_; 
wire _abc_19873_new_n1976_; 
wire _abc_19873_new_n1977_; 
wire _abc_19873_new_n1979_; 
wire _abc_19873_new_n1980_; 
wire _abc_19873_new_n1981_; 
wire _abc_19873_new_n1983_; 
wire _abc_19873_new_n1984_; 
wire _abc_19873_new_n1985_; 
wire _abc_19873_new_n1987_; 
wire _abc_19873_new_n1988_; 
wire _abc_19873_new_n1989_; 
wire _abc_19873_new_n1991_; 
wire _abc_19873_new_n1992_; 
wire _abc_19873_new_n1993_; 
wire _abc_19873_new_n1995_; 
wire _abc_19873_new_n1996_; 
wire _abc_19873_new_n1997_; 
wire _abc_19873_new_n1999_; 
wire _abc_19873_new_n2000_; 
wire _abc_19873_new_n2001_; 
wire _abc_19873_new_n2003_; 
wire _abc_19873_new_n2004_; 
wire _abc_19873_new_n2005_; 
wire _abc_19873_new_n2007_; 
wire _abc_19873_new_n2008_; 
wire _abc_19873_new_n2009_; 
wire _abc_19873_new_n2011_; 
wire _abc_19873_new_n2012_; 
wire _abc_19873_new_n2013_; 
wire _abc_19873_new_n2015_; 
wire _abc_19873_new_n2016_; 
wire _abc_19873_new_n2017_; 
wire _abc_19873_new_n2019_; 
wire _abc_19873_new_n2020_; 
wire _abc_19873_new_n2021_; 
wire _abc_19873_new_n2023_; 
wire _abc_19873_new_n2024_; 
wire _abc_19873_new_n2025_; 
wire _abc_19873_new_n2027_; 
wire _abc_19873_new_n2028_; 
wire _abc_19873_new_n2029_; 
wire _abc_19873_new_n2031_; 
wire _abc_19873_new_n2032_; 
wire _abc_19873_new_n2033_; 
wire _abc_19873_new_n2035_; 
wire _abc_19873_new_n2036_; 
wire _abc_19873_new_n2037_; 
wire _abc_19873_new_n2039_; 
wire _abc_19873_new_n2040_; 
wire _abc_19873_new_n2041_; 
wire _abc_19873_new_n2043_; 
wire _abc_19873_new_n2044_; 
wire _abc_19873_new_n2045_; 
wire _abc_19873_new_n2047_; 
wire _abc_19873_new_n2048_; 
wire _abc_19873_new_n2049_; 
wire _abc_19873_new_n2051_; 
wire _abc_19873_new_n2052_; 
wire _abc_19873_new_n2053_; 
wire _abc_19873_new_n2055_; 
wire _abc_19873_new_n2056_; 
wire _abc_19873_new_n2057_; 
wire _abc_19873_new_n2059_; 
wire _abc_19873_new_n2060_; 
wire _abc_19873_new_n2061_; 
wire _abc_19873_new_n2063_; 
wire _abc_19873_new_n2064_; 
wire _abc_19873_new_n2065_; 
wire _abc_19873_new_n2067_; 
wire _abc_19873_new_n2068_; 
wire _abc_19873_new_n2069_; 
wire _abc_19873_new_n2071_; 
wire _abc_19873_new_n2072_; 
wire _abc_19873_new_n2073_; 
wire _abc_19873_new_n2075_; 
wire _abc_19873_new_n2076_; 
wire _abc_19873_new_n2077_; 
wire _abc_19873_new_n2079_; 
wire _abc_19873_new_n2080_; 
wire _abc_19873_new_n2081_; 
wire _abc_19873_new_n2083_; 
wire _abc_19873_new_n2084_; 
wire _abc_19873_new_n2085_; 
wire _abc_19873_new_n2087_; 
wire _abc_19873_new_n2088_; 
wire _abc_19873_new_n2089_; 
wire _abc_19873_new_n2091_; 
wire _abc_19873_new_n2092_; 
wire _abc_19873_new_n2093_; 
wire _abc_19873_new_n2095_; 
wire _abc_19873_new_n2096_; 
wire _abc_19873_new_n2097_; 
wire _abc_19873_new_n2099_; 
wire _abc_19873_new_n2100_; 
wire _abc_19873_new_n2101_; 
wire _abc_19873_new_n2103_; 
wire _abc_19873_new_n2104_; 
wire _abc_19873_new_n2105_; 
wire _abc_19873_new_n2107_; 
wire _abc_19873_new_n2108_; 
wire _abc_19873_new_n2109_; 
wire _abc_19873_new_n2111_; 
wire _abc_19873_new_n2112_; 
wire _abc_19873_new_n2113_; 
wire _abc_19873_new_n2115_; 
wire _abc_19873_new_n2116_; 
wire _abc_19873_new_n2117_; 
wire _abc_19873_new_n2119_; 
wire _abc_19873_new_n2120_; 
wire _abc_19873_new_n2121_; 
wire _abc_19873_new_n2122_; 
wire _abc_19873_new_n2123_; 
wire _abc_19873_new_n2124_; 
wire _abc_19873_new_n2125_; 
wire _abc_19873_new_n2127_; 
wire _abc_19873_new_n2128_; 
wire _abc_19873_new_n2129_; 
wire _abc_19873_new_n2130_; 
wire _abc_19873_new_n2131_; 
wire _abc_19873_new_n2133_; 
wire _abc_19873_new_n2134_; 
wire _abc_19873_new_n2135_; 
wire _abc_19873_new_n2136_; 
wire _abc_19873_new_n2137_; 
wire _abc_19873_new_n2139_; 
wire _abc_19873_new_n2140_; 
wire _abc_19873_new_n2141_; 
wire _abc_19873_new_n2142_; 
wire _abc_19873_new_n2143_; 
wire _abc_19873_new_n2145_; 
wire _abc_19873_new_n2146_; 
wire _abc_19873_new_n2147_; 
wire _abc_19873_new_n2148_; 
wire _abc_19873_new_n2149_; 
wire _abc_19873_new_n2151_; 
wire _abc_19873_new_n2152_; 
wire _abc_19873_new_n2153_; 
wire _abc_19873_new_n2154_; 
wire _abc_19873_new_n2155_; 
wire _abc_19873_new_n2157_; 
wire _abc_19873_new_n2158_; 
wire _abc_19873_new_n2159_; 
wire _abc_19873_new_n2160_; 
wire _abc_19873_new_n2161_; 
wire _abc_19873_new_n2163_; 
wire _abc_19873_new_n2164_; 
wire _abc_19873_new_n2165_; 
wire _abc_19873_new_n2166_; 
wire _abc_19873_new_n2167_; 
wire _abc_19873_new_n2169_; 
wire _abc_19873_new_n2170_; 
wire _abc_19873_new_n2171_; 
wire _abc_19873_new_n2172_; 
wire _abc_19873_new_n2173_; 
wire _abc_19873_new_n2175_; 
wire _abc_19873_new_n2176_; 
wire _abc_19873_new_n2177_; 
wire _abc_19873_new_n2178_; 
wire _abc_19873_new_n2179_; 
wire _abc_19873_new_n2181_; 
wire _abc_19873_new_n2182_; 
wire _abc_19873_new_n2183_; 
wire _abc_19873_new_n2184_; 
wire _abc_19873_new_n2185_; 
wire _abc_19873_new_n2187_; 
wire _abc_19873_new_n2188_; 
wire _abc_19873_new_n2189_; 
wire _abc_19873_new_n2190_; 
wire _abc_19873_new_n2191_; 
wire _abc_19873_new_n2193_; 
wire _abc_19873_new_n2194_; 
wire _abc_19873_new_n2195_; 
wire _abc_19873_new_n2196_; 
wire _abc_19873_new_n2197_; 
wire _abc_19873_new_n2199_; 
wire _abc_19873_new_n2200_; 
wire _abc_19873_new_n2201_; 
wire _abc_19873_new_n2202_; 
wire _abc_19873_new_n2203_; 
wire _abc_19873_new_n2205_; 
wire _abc_19873_new_n2206_; 
wire _abc_19873_new_n2207_; 
wire _abc_19873_new_n2208_; 
wire _abc_19873_new_n2209_; 
wire _abc_19873_new_n2211_; 
wire _abc_19873_new_n2212_; 
wire _abc_19873_new_n2213_; 
wire _abc_19873_new_n2214_; 
wire _abc_19873_new_n2215_; 
wire _abc_19873_new_n2217_; 
wire _abc_19873_new_n2218_; 
wire _abc_19873_new_n2219_; 
wire _abc_19873_new_n2220_; 
wire _abc_19873_new_n2221_; 
wire _abc_19873_new_n2223_; 
wire _abc_19873_new_n2224_; 
wire _abc_19873_new_n2225_; 
wire _abc_19873_new_n2226_; 
wire _abc_19873_new_n2227_; 
wire _abc_19873_new_n2229_; 
wire _abc_19873_new_n2230_; 
wire _abc_19873_new_n2231_; 
wire _abc_19873_new_n2232_; 
wire _abc_19873_new_n2233_; 
wire _abc_19873_new_n2235_; 
wire _abc_19873_new_n2236_; 
wire _abc_19873_new_n2237_; 
wire _abc_19873_new_n2238_; 
wire _abc_19873_new_n2239_; 
wire _abc_19873_new_n2241_; 
wire _abc_19873_new_n2242_; 
wire _abc_19873_new_n2243_; 
wire _abc_19873_new_n2244_; 
wire _abc_19873_new_n2245_; 
wire _abc_19873_new_n2247_; 
wire _abc_19873_new_n2248_; 
wire _abc_19873_new_n2249_; 
wire _abc_19873_new_n2250_; 
wire _abc_19873_new_n2251_; 
wire _abc_19873_new_n2253_; 
wire _abc_19873_new_n2254_; 
wire _abc_19873_new_n2255_; 
wire _abc_19873_new_n2256_; 
wire _abc_19873_new_n2257_; 
wire _abc_19873_new_n2259_; 
wire _abc_19873_new_n2260_; 
wire _abc_19873_new_n2261_; 
wire _abc_19873_new_n2262_; 
wire _abc_19873_new_n2263_; 
wire _abc_19873_new_n2265_; 
wire _abc_19873_new_n2266_; 
wire _abc_19873_new_n2267_; 
wire _abc_19873_new_n2268_; 
wire _abc_19873_new_n2269_; 
wire _abc_19873_new_n2271_; 
wire _abc_19873_new_n2272_; 
wire _abc_19873_new_n2273_; 
wire _abc_19873_new_n2274_; 
wire _abc_19873_new_n2275_; 
wire _abc_19873_new_n2277_; 
wire _abc_19873_new_n2278_; 
wire _abc_19873_new_n2279_; 
wire _abc_19873_new_n2280_; 
wire _abc_19873_new_n2281_; 
wire _abc_19873_new_n2283_; 
wire _abc_19873_new_n2284_; 
wire _abc_19873_new_n2285_; 
wire _abc_19873_new_n2286_; 
wire _abc_19873_new_n2287_; 
wire _abc_19873_new_n2289_; 
wire _abc_19873_new_n2290_; 
wire _abc_19873_new_n2291_; 
wire _abc_19873_new_n2292_; 
wire _abc_19873_new_n2293_; 
wire _abc_19873_new_n2295_; 
wire _abc_19873_new_n2296_; 
wire _abc_19873_new_n2297_; 
wire _abc_19873_new_n2298_; 
wire _abc_19873_new_n2299_; 
wire _abc_19873_new_n2301_; 
wire _abc_19873_new_n2302_; 
wire _abc_19873_new_n2303_; 
wire _abc_19873_new_n2304_; 
wire _abc_19873_new_n2305_; 
wire _abc_19873_new_n2307_; 
wire _abc_19873_new_n2308_; 
wire _abc_19873_new_n2309_; 
wire _abc_19873_new_n2310_; 
wire _abc_19873_new_n2311_; 
wire _abc_19873_new_n2313_; 
wire _abc_19873_new_n2314_; 
wire _abc_19873_new_n2315_; 
wire _abc_19873_new_n2316_; 
wire _abc_19873_new_n2317_; 
wire _abc_19873_new_n2319_; 
wire _abc_19873_new_n2320_; 
wire _abc_19873_new_n2321_; 
wire _abc_19873_new_n2322_; 
wire _abc_19873_new_n2324_; 
wire _abc_19873_new_n2325_; 
wire _abc_19873_new_n2326_; 
wire _abc_19873_new_n2327_; 
wire _abc_19873_new_n2329_; 
wire _abc_19873_new_n2330_; 
wire _abc_19873_new_n2331_; 
wire _abc_19873_new_n2332_; 
wire _abc_19873_new_n2334_; 
wire _abc_19873_new_n2335_; 
wire _abc_19873_new_n2336_; 
wire _abc_19873_new_n2337_; 
wire _abc_19873_new_n2339_; 
wire _abc_19873_new_n2340_; 
wire _abc_19873_new_n2341_; 
wire _abc_19873_new_n2342_; 
wire _abc_19873_new_n2344_; 
wire _abc_19873_new_n2345_; 
wire _abc_19873_new_n2346_; 
wire _abc_19873_new_n2347_; 
wire _abc_19873_new_n2349_; 
wire _abc_19873_new_n2350_; 
wire _abc_19873_new_n2351_; 
wire _abc_19873_new_n2352_; 
wire _abc_19873_new_n2354_; 
wire _abc_19873_new_n2355_; 
wire _abc_19873_new_n2356_; 
wire _abc_19873_new_n2357_; 
wire _abc_19873_new_n2359_; 
wire _abc_19873_new_n2360_; 
wire _abc_19873_new_n2361_; 
wire _abc_19873_new_n2362_; 
wire _abc_19873_new_n2364_; 
wire _abc_19873_new_n2365_; 
wire _abc_19873_new_n2366_; 
wire _abc_19873_new_n2367_; 
wire _abc_19873_new_n2369_; 
wire _abc_19873_new_n2370_; 
wire _abc_19873_new_n2371_; 
wire _abc_19873_new_n2372_; 
wire _abc_19873_new_n2374_; 
wire _abc_19873_new_n2375_; 
wire _abc_19873_new_n2376_; 
wire _abc_19873_new_n2377_; 
wire _abc_19873_new_n2379_; 
wire _abc_19873_new_n2380_; 
wire _abc_19873_new_n2381_; 
wire _abc_19873_new_n2382_; 
wire _abc_19873_new_n2384_; 
wire _abc_19873_new_n2385_; 
wire _abc_19873_new_n2386_; 
wire _abc_19873_new_n2387_; 
wire _abc_19873_new_n2389_; 
wire _abc_19873_new_n2390_; 
wire _abc_19873_new_n2391_; 
wire _abc_19873_new_n2392_; 
wire _abc_19873_new_n2394_; 
wire _abc_19873_new_n2395_; 
wire _abc_19873_new_n2396_; 
wire _abc_19873_new_n2397_; 
wire _abc_19873_new_n2399_; 
wire _abc_19873_new_n2400_; 
wire _abc_19873_new_n2401_; 
wire _abc_19873_new_n2402_; 
wire _abc_19873_new_n2404_; 
wire _abc_19873_new_n2405_; 
wire _abc_19873_new_n2406_; 
wire _abc_19873_new_n2407_; 
wire _abc_19873_new_n2409_; 
wire _abc_19873_new_n2410_; 
wire _abc_19873_new_n2411_; 
wire _abc_19873_new_n2412_; 
wire _abc_19873_new_n2414_; 
wire _abc_19873_new_n2415_; 
wire _abc_19873_new_n2416_; 
wire _abc_19873_new_n2417_; 
wire _abc_19873_new_n2419_; 
wire _abc_19873_new_n2420_; 
wire _abc_19873_new_n2421_; 
wire _abc_19873_new_n2422_; 
wire _abc_19873_new_n2424_; 
wire _abc_19873_new_n2425_; 
wire _abc_19873_new_n2426_; 
wire _abc_19873_new_n2427_; 
wire _abc_19873_new_n2429_; 
wire _abc_19873_new_n2430_; 
wire _abc_19873_new_n2431_; 
wire _abc_19873_new_n2432_; 
wire _abc_19873_new_n2434_; 
wire _abc_19873_new_n2435_; 
wire _abc_19873_new_n2436_; 
wire _abc_19873_new_n2437_; 
wire _abc_19873_new_n2439_; 
wire _abc_19873_new_n2440_; 
wire _abc_19873_new_n2441_; 
wire _abc_19873_new_n2442_; 
wire _abc_19873_new_n2444_; 
wire _abc_19873_new_n2445_; 
wire _abc_19873_new_n2446_; 
wire _abc_19873_new_n2447_; 
wire _abc_19873_new_n2449_; 
wire _abc_19873_new_n2450_; 
wire _abc_19873_new_n2451_; 
wire _abc_19873_new_n2452_; 
wire _abc_19873_new_n2454_; 
wire _abc_19873_new_n2455_; 
wire _abc_19873_new_n2456_; 
wire _abc_19873_new_n2457_; 
wire _abc_19873_new_n2459_; 
wire _abc_19873_new_n2460_; 
wire _abc_19873_new_n2461_; 
wire _abc_19873_new_n2462_; 
wire _abc_19873_new_n2464_; 
wire _abc_19873_new_n2465_; 
wire _abc_19873_new_n2466_; 
wire _abc_19873_new_n2467_; 
wire _abc_19873_new_n2469_; 
wire _abc_19873_new_n2470_; 
wire _abc_19873_new_n2471_; 
wire _abc_19873_new_n2472_; 
wire _abc_19873_new_n2474_; 
wire _abc_19873_new_n2475_; 
wire _abc_19873_new_n2476_; 
wire _abc_19873_new_n2477_; 
wire _abc_19873_new_n2478_; 
wire _abc_19873_new_n2480_; 
wire _abc_19873_new_n2481_; 
wire _abc_19873_new_n2482_; 
wire _abc_19873_new_n2483_; 
wire _abc_19873_new_n2485_; 
wire _abc_19873_new_n2486_; 
wire _abc_19873_new_n2487_; 
wire _abc_19873_new_n2488_; 
wire _abc_19873_new_n2490_; 
wire _abc_19873_new_n2491_; 
wire _abc_19873_new_n2492_; 
wire _abc_19873_new_n2493_; 
wire _abc_19873_new_n2495_; 
wire _abc_19873_new_n2496_; 
wire _abc_19873_new_n2497_; 
wire _abc_19873_new_n2498_; 
wire _abc_19873_new_n2500_; 
wire _abc_19873_new_n2501_; 
wire _abc_19873_new_n2502_; 
wire _abc_19873_new_n2503_; 
wire _abc_19873_new_n2505_; 
wire _abc_19873_new_n2506_; 
wire _abc_19873_new_n2507_; 
wire _abc_19873_new_n2508_; 
wire _abc_19873_new_n2510_; 
wire _abc_19873_new_n2511_; 
wire _abc_19873_new_n2512_; 
wire _abc_19873_new_n2513_; 
wire _abc_19873_new_n2515_; 
wire _abc_19873_new_n2516_; 
wire _abc_19873_new_n2517_; 
wire _abc_19873_new_n2518_; 
wire _abc_19873_new_n2520_; 
wire _abc_19873_new_n2521_; 
wire _abc_19873_new_n2522_; 
wire _abc_19873_new_n2523_; 
wire _abc_19873_new_n2525_; 
wire _abc_19873_new_n2526_; 
wire _abc_19873_new_n2527_; 
wire _abc_19873_new_n2528_; 
wire _abc_19873_new_n2530_; 
wire _abc_19873_new_n2531_; 
wire _abc_19873_new_n2532_; 
wire _abc_19873_new_n2533_; 
wire _abc_19873_new_n2535_; 
wire _abc_19873_new_n2536_; 
wire _abc_19873_new_n2537_; 
wire _abc_19873_new_n2538_; 
wire _abc_19873_new_n2540_; 
wire _abc_19873_new_n2541_; 
wire _abc_19873_new_n2542_; 
wire _abc_19873_new_n2543_; 
wire _abc_19873_new_n2545_; 
wire _abc_19873_new_n2546_; 
wire _abc_19873_new_n2547_; 
wire _abc_19873_new_n2548_; 
wire _abc_19873_new_n2550_; 
wire _abc_19873_new_n2551_; 
wire _abc_19873_new_n2552_; 
wire _abc_19873_new_n2553_; 
wire _abc_19873_new_n2555_; 
wire _abc_19873_new_n2556_; 
wire _abc_19873_new_n2557_; 
wire _abc_19873_new_n2558_; 
wire _abc_19873_new_n2560_; 
wire _abc_19873_new_n2561_; 
wire _abc_19873_new_n2562_; 
wire _abc_19873_new_n2563_; 
wire _abc_19873_new_n2565_; 
wire _abc_19873_new_n2566_; 
wire _abc_19873_new_n2567_; 
wire _abc_19873_new_n2568_; 
wire _abc_19873_new_n2570_; 
wire _abc_19873_new_n2571_; 
wire _abc_19873_new_n2572_; 
wire _abc_19873_new_n2573_; 
wire _abc_19873_new_n2575_; 
wire _abc_19873_new_n2576_; 
wire _abc_19873_new_n2577_; 
wire _abc_19873_new_n2578_; 
wire _abc_19873_new_n2580_; 
wire _abc_19873_new_n2581_; 
wire _abc_19873_new_n2582_; 
wire _abc_19873_new_n2583_; 
wire _abc_19873_new_n2585_; 
wire _abc_19873_new_n2586_; 
wire _abc_19873_new_n2587_; 
wire _abc_19873_new_n2588_; 
wire _abc_19873_new_n2590_; 
wire _abc_19873_new_n2591_; 
wire _abc_19873_new_n2592_; 
wire _abc_19873_new_n2593_; 
wire _abc_19873_new_n2595_; 
wire _abc_19873_new_n2596_; 
wire _abc_19873_new_n2597_; 
wire _abc_19873_new_n2598_; 
wire _abc_19873_new_n2600_; 
wire _abc_19873_new_n2601_; 
wire _abc_19873_new_n2602_; 
wire _abc_19873_new_n2603_; 
wire _abc_19873_new_n2605_; 
wire _abc_19873_new_n2606_; 
wire _abc_19873_new_n2607_; 
wire _abc_19873_new_n2608_; 
wire _abc_19873_new_n2610_; 
wire _abc_19873_new_n2611_; 
wire _abc_19873_new_n2612_; 
wire _abc_19873_new_n2613_; 
wire _abc_19873_new_n2615_; 
wire _abc_19873_new_n2616_; 
wire _abc_19873_new_n2617_; 
wire _abc_19873_new_n2618_; 
wire _abc_19873_new_n2620_; 
wire _abc_19873_new_n2621_; 
wire _abc_19873_new_n2622_; 
wire _abc_19873_new_n2623_; 
wire _abc_19873_new_n2625_; 
wire _abc_19873_new_n2626_; 
wire _abc_19873_new_n2627_; 
wire _abc_19873_new_n2628_; 
wire _abc_19873_new_n2630_; 
wire _abc_19873_new_n2631_; 
wire _abc_19873_new_n2632_; 
wire _abc_19873_new_n2633_; 
wire _abc_19873_new_n2635_; 
wire _abc_19873_new_n2636_; 
wire _abc_19873_new_n2637_; 
wire _abc_19873_new_n2638_; 
wire _abc_19873_new_n2639_; 
wire _abc_19873_new_n2641_; 
wire _abc_19873_new_n2642_; 
wire _abc_19873_new_n2643_; 
wire _abc_19873_new_n2644_; 
wire _abc_19873_new_n2646_; 
wire _abc_19873_new_n2647_; 
wire _abc_19873_new_n2648_; 
wire _abc_19873_new_n2649_; 
wire _abc_19873_new_n2651_; 
wire _abc_19873_new_n2652_; 
wire _abc_19873_new_n2653_; 
wire _abc_19873_new_n2654_; 
wire _abc_19873_new_n2656_; 
wire _abc_19873_new_n2657_; 
wire _abc_19873_new_n2658_; 
wire _abc_19873_new_n2659_; 
wire _abc_19873_new_n2661_; 
wire _abc_19873_new_n2662_; 
wire _abc_19873_new_n2663_; 
wire _abc_19873_new_n2664_; 
wire _abc_19873_new_n2666_; 
wire _abc_19873_new_n2667_; 
wire _abc_19873_new_n2668_; 
wire _abc_19873_new_n2669_; 
wire _abc_19873_new_n2671_; 
wire _abc_19873_new_n2672_; 
wire _abc_19873_new_n2673_; 
wire _abc_19873_new_n2674_; 
wire _abc_19873_new_n2676_; 
wire _abc_19873_new_n2677_; 
wire _abc_19873_new_n2678_; 
wire _abc_19873_new_n2679_; 
wire _abc_19873_new_n2681_; 
wire _abc_19873_new_n2682_; 
wire _abc_19873_new_n2683_; 
wire _abc_19873_new_n2684_; 
wire _abc_19873_new_n2686_; 
wire _abc_19873_new_n2687_; 
wire _abc_19873_new_n2688_; 
wire _abc_19873_new_n2689_; 
wire _abc_19873_new_n2691_; 
wire _abc_19873_new_n2692_; 
wire _abc_19873_new_n2693_; 
wire _abc_19873_new_n2694_; 
wire _abc_19873_new_n2696_; 
wire _abc_19873_new_n2697_; 
wire _abc_19873_new_n2698_; 
wire _abc_19873_new_n2699_; 
wire _abc_19873_new_n2701_; 
wire _abc_19873_new_n2702_; 
wire _abc_19873_new_n2703_; 
wire _abc_19873_new_n2704_; 
wire _abc_19873_new_n2706_; 
wire _abc_19873_new_n2707_; 
wire _abc_19873_new_n2708_; 
wire _abc_19873_new_n2709_; 
wire _abc_19873_new_n2711_; 
wire _abc_19873_new_n2712_; 
wire _abc_19873_new_n2713_; 
wire _abc_19873_new_n2714_; 
wire _abc_19873_new_n2716_; 
wire _abc_19873_new_n2717_; 
wire _abc_19873_new_n2718_; 
wire _abc_19873_new_n2719_; 
wire _abc_19873_new_n2721_; 
wire _abc_19873_new_n2722_; 
wire _abc_19873_new_n2723_; 
wire _abc_19873_new_n2724_; 
wire _abc_19873_new_n2726_; 
wire _abc_19873_new_n2727_; 
wire _abc_19873_new_n2728_; 
wire _abc_19873_new_n2729_; 
wire _abc_19873_new_n2731_; 
wire _abc_19873_new_n2732_; 
wire _abc_19873_new_n2733_; 
wire _abc_19873_new_n2734_; 
wire _abc_19873_new_n2736_; 
wire _abc_19873_new_n2737_; 
wire _abc_19873_new_n2738_; 
wire _abc_19873_new_n2739_; 
wire _abc_19873_new_n2741_; 
wire _abc_19873_new_n2742_; 
wire _abc_19873_new_n2743_; 
wire _abc_19873_new_n2744_; 
wire _abc_19873_new_n2746_; 
wire _abc_19873_new_n2747_; 
wire _abc_19873_new_n2748_; 
wire _abc_19873_new_n2749_; 
wire _abc_19873_new_n2751_; 
wire _abc_19873_new_n2752_; 
wire _abc_19873_new_n2753_; 
wire _abc_19873_new_n2754_; 
wire _abc_19873_new_n2756_; 
wire _abc_19873_new_n2757_; 
wire _abc_19873_new_n2758_; 
wire _abc_19873_new_n2759_; 
wire _abc_19873_new_n2761_; 
wire _abc_19873_new_n2762_; 
wire _abc_19873_new_n2763_; 
wire _abc_19873_new_n2764_; 
wire _abc_19873_new_n2766_; 
wire _abc_19873_new_n2767_; 
wire _abc_19873_new_n2768_; 
wire _abc_19873_new_n2769_; 
wire _abc_19873_new_n2771_; 
wire _abc_19873_new_n2772_; 
wire _abc_19873_new_n2773_; 
wire _abc_19873_new_n2774_; 
wire _abc_19873_new_n2776_; 
wire _abc_19873_new_n2777_; 
wire _abc_19873_new_n2778_; 
wire _abc_19873_new_n2779_; 
wire _abc_19873_new_n2781_; 
wire _abc_19873_new_n2782_; 
wire _abc_19873_new_n2783_; 
wire _abc_19873_new_n2784_; 
wire _abc_19873_new_n2786_; 
wire _abc_19873_new_n2787_; 
wire _abc_19873_new_n2788_; 
wire _abc_19873_new_n2789_; 
wire _abc_19873_new_n2791_; 
wire _abc_19873_new_n2792_; 
wire _abc_19873_new_n2793_; 
wire _abc_19873_new_n2794_; 
wire _abc_19873_new_n2796_; 
wire _abc_19873_new_n2797_; 
wire _abc_19873_new_n2798_; 
wire _abc_19873_new_n2799_; 
wire _abc_19873_new_n2800_; 
wire _abc_19873_new_n2802_; 
wire _abc_19873_new_n2803_; 
wire _abc_19873_new_n2804_; 
wire _abc_19873_new_n2805_; 
wire _abc_19873_new_n2807_; 
wire _abc_19873_new_n2808_; 
wire _abc_19873_new_n2809_; 
wire _abc_19873_new_n2810_; 
wire _abc_19873_new_n2812_; 
wire _abc_19873_new_n2813_; 
wire _abc_19873_new_n2814_; 
wire _abc_19873_new_n2815_; 
wire _abc_19873_new_n2817_; 
wire _abc_19873_new_n2818_; 
wire _abc_19873_new_n2819_; 
wire _abc_19873_new_n2820_; 
wire _abc_19873_new_n2822_; 
wire _abc_19873_new_n2823_; 
wire _abc_19873_new_n2824_; 
wire _abc_19873_new_n2825_; 
wire _abc_19873_new_n2827_; 
wire _abc_19873_new_n2828_; 
wire _abc_19873_new_n2829_; 
wire _abc_19873_new_n2830_; 
wire _abc_19873_new_n2832_; 
wire _abc_19873_new_n2833_; 
wire _abc_19873_new_n2834_; 
wire _abc_19873_new_n2835_; 
wire _abc_19873_new_n2837_; 
wire _abc_19873_new_n2838_; 
wire _abc_19873_new_n2839_; 
wire _abc_19873_new_n2840_; 
wire _abc_19873_new_n2842_; 
wire _abc_19873_new_n2843_; 
wire _abc_19873_new_n2844_; 
wire _abc_19873_new_n2845_; 
wire _abc_19873_new_n2847_; 
wire _abc_19873_new_n2848_; 
wire _abc_19873_new_n2849_; 
wire _abc_19873_new_n2850_; 
wire _abc_19873_new_n2852_; 
wire _abc_19873_new_n2853_; 
wire _abc_19873_new_n2854_; 
wire _abc_19873_new_n2855_; 
wire _abc_19873_new_n2857_; 
wire _abc_19873_new_n2858_; 
wire _abc_19873_new_n2859_; 
wire _abc_19873_new_n2860_; 
wire _abc_19873_new_n2862_; 
wire _abc_19873_new_n2863_; 
wire _abc_19873_new_n2864_; 
wire _abc_19873_new_n2865_; 
wire _abc_19873_new_n2867_; 
wire _abc_19873_new_n2868_; 
wire _abc_19873_new_n2869_; 
wire _abc_19873_new_n2870_; 
wire _abc_19873_new_n2872_; 
wire _abc_19873_new_n2873_; 
wire _abc_19873_new_n2874_; 
wire _abc_19873_new_n2875_; 
wire _abc_19873_new_n2877_; 
wire _abc_19873_new_n2878_; 
wire _abc_19873_new_n2879_; 
wire _abc_19873_new_n2880_; 
wire _abc_19873_new_n2882_; 
wire _abc_19873_new_n2883_; 
wire _abc_19873_new_n2884_; 
wire _abc_19873_new_n2885_; 
wire _abc_19873_new_n2887_; 
wire _abc_19873_new_n2888_; 
wire _abc_19873_new_n2889_; 
wire _abc_19873_new_n2890_; 
wire _abc_19873_new_n2892_; 
wire _abc_19873_new_n2893_; 
wire _abc_19873_new_n2894_; 
wire _abc_19873_new_n2895_; 
wire _abc_19873_new_n2897_; 
wire _abc_19873_new_n2898_; 
wire _abc_19873_new_n2899_; 
wire _abc_19873_new_n2900_; 
wire _abc_19873_new_n2902_; 
wire _abc_19873_new_n2903_; 
wire _abc_19873_new_n2904_; 
wire _abc_19873_new_n2905_; 
wire _abc_19873_new_n2907_; 
wire _abc_19873_new_n2908_; 
wire _abc_19873_new_n2909_; 
wire _abc_19873_new_n2910_; 
wire _abc_19873_new_n2912_; 
wire _abc_19873_new_n2913_; 
wire _abc_19873_new_n2914_; 
wire _abc_19873_new_n2915_; 
wire _abc_19873_new_n2917_; 
wire _abc_19873_new_n2918_; 
wire _abc_19873_new_n2919_; 
wire _abc_19873_new_n2920_; 
wire _abc_19873_new_n2922_; 
wire _abc_19873_new_n2923_; 
wire _abc_19873_new_n2924_; 
wire _abc_19873_new_n2925_; 
wire _abc_19873_new_n2927_; 
wire _abc_19873_new_n2928_; 
wire _abc_19873_new_n2929_; 
wire _abc_19873_new_n2930_; 
wire _abc_19873_new_n2932_; 
wire _abc_19873_new_n2933_; 
wire _abc_19873_new_n2934_; 
wire _abc_19873_new_n2935_; 
wire _abc_19873_new_n2937_; 
wire _abc_19873_new_n2938_; 
wire _abc_19873_new_n2939_; 
wire _abc_19873_new_n2940_; 
wire _abc_19873_new_n2942_; 
wire _abc_19873_new_n2943_; 
wire _abc_19873_new_n2944_; 
wire _abc_19873_new_n2945_; 
wire _abc_19873_new_n2947_; 
wire _abc_19873_new_n2948_; 
wire _abc_19873_new_n2949_; 
wire _abc_19873_new_n2950_; 
wire _abc_19873_new_n2952_; 
wire _abc_19873_new_n2953_; 
wire _abc_19873_new_n2954_; 
wire _abc_19873_new_n2955_; 
wire _abc_19873_new_n2957_; 
wire _abc_19873_new_n2958_; 
wire _abc_19873_new_n2959_; 
wire _abc_19873_new_n2960_; 
wire _abc_19873_new_n2961_; 
wire _abc_19873_new_n2963_; 
wire _abc_19873_new_n2964_; 
wire _abc_19873_new_n2965_; 
wire _abc_19873_new_n2966_; 
wire _abc_19873_new_n2968_; 
wire _abc_19873_new_n2969_; 
wire _abc_19873_new_n2970_; 
wire _abc_19873_new_n2971_; 
wire _abc_19873_new_n2973_; 
wire _abc_19873_new_n2974_; 
wire _abc_19873_new_n2975_; 
wire _abc_19873_new_n2976_; 
wire _abc_19873_new_n2978_; 
wire _abc_19873_new_n2979_; 
wire _abc_19873_new_n2980_; 
wire _abc_19873_new_n2981_; 
wire _abc_19873_new_n2983_; 
wire _abc_19873_new_n2984_; 
wire _abc_19873_new_n2985_; 
wire _abc_19873_new_n2986_; 
wire _abc_19873_new_n2988_; 
wire _abc_19873_new_n2989_; 
wire _abc_19873_new_n2990_; 
wire _abc_19873_new_n2991_; 
wire _abc_19873_new_n2993_; 
wire _abc_19873_new_n2994_; 
wire _abc_19873_new_n2995_; 
wire _abc_19873_new_n2996_; 
wire _abc_19873_new_n2998_; 
wire _abc_19873_new_n2999_; 
wire _abc_19873_new_n3000_; 
wire _abc_19873_new_n3001_; 
wire _abc_19873_new_n3003_; 
wire _abc_19873_new_n3004_; 
wire _abc_19873_new_n3005_; 
wire _abc_19873_new_n3006_; 
wire _abc_19873_new_n3008_; 
wire _abc_19873_new_n3009_; 
wire _abc_19873_new_n3010_; 
wire _abc_19873_new_n3011_; 
wire _abc_19873_new_n3013_; 
wire _abc_19873_new_n3014_; 
wire _abc_19873_new_n3015_; 
wire _abc_19873_new_n3016_; 
wire _abc_19873_new_n3018_; 
wire _abc_19873_new_n3019_; 
wire _abc_19873_new_n3020_; 
wire _abc_19873_new_n3021_; 
wire _abc_19873_new_n3023_; 
wire _abc_19873_new_n3024_; 
wire _abc_19873_new_n3025_; 
wire _abc_19873_new_n3026_; 
wire _abc_19873_new_n3028_; 
wire _abc_19873_new_n3029_; 
wire _abc_19873_new_n3030_; 
wire _abc_19873_new_n3031_; 
wire _abc_19873_new_n3033_; 
wire _abc_19873_new_n3034_; 
wire _abc_19873_new_n3035_; 
wire _abc_19873_new_n3036_; 
wire _abc_19873_new_n3038_; 
wire _abc_19873_new_n3039_; 
wire _abc_19873_new_n3040_; 
wire _abc_19873_new_n3041_; 
wire _abc_19873_new_n3043_; 
wire _abc_19873_new_n3044_; 
wire _abc_19873_new_n3045_; 
wire _abc_19873_new_n3046_; 
wire _abc_19873_new_n3048_; 
wire _abc_19873_new_n3049_; 
wire _abc_19873_new_n3050_; 
wire _abc_19873_new_n3051_; 
wire _abc_19873_new_n3053_; 
wire _abc_19873_new_n3054_; 
wire _abc_19873_new_n3055_; 
wire _abc_19873_new_n3056_; 
wire _abc_19873_new_n3058_; 
wire _abc_19873_new_n3059_; 
wire _abc_19873_new_n3060_; 
wire _abc_19873_new_n3061_; 
wire _abc_19873_new_n3063_; 
wire _abc_19873_new_n3064_; 
wire _abc_19873_new_n3065_; 
wire _abc_19873_new_n3066_; 
wire _abc_19873_new_n3068_; 
wire _abc_19873_new_n3069_; 
wire _abc_19873_new_n3070_; 
wire _abc_19873_new_n3071_; 
wire _abc_19873_new_n3073_; 
wire _abc_19873_new_n3074_; 
wire _abc_19873_new_n3075_; 
wire _abc_19873_new_n3076_; 
wire _abc_19873_new_n3078_; 
wire _abc_19873_new_n3079_; 
wire _abc_19873_new_n3080_; 
wire _abc_19873_new_n3081_; 
wire _abc_19873_new_n3083_; 
wire _abc_19873_new_n3084_; 
wire _abc_19873_new_n3085_; 
wire _abc_19873_new_n3086_; 
wire _abc_19873_new_n3088_; 
wire _abc_19873_new_n3089_; 
wire _abc_19873_new_n3090_; 
wire _abc_19873_new_n3091_; 
wire _abc_19873_new_n3093_; 
wire _abc_19873_new_n3094_; 
wire _abc_19873_new_n3095_; 
wire _abc_19873_new_n3096_; 
wire _abc_19873_new_n3098_; 
wire _abc_19873_new_n3099_; 
wire _abc_19873_new_n3100_; 
wire _abc_19873_new_n3101_; 
wire _abc_19873_new_n3103_; 
wire _abc_19873_new_n3104_; 
wire _abc_19873_new_n3105_; 
wire _abc_19873_new_n3106_; 
wire _abc_19873_new_n3108_; 
wire _abc_19873_new_n3109_; 
wire _abc_19873_new_n3110_; 
wire _abc_19873_new_n3111_; 
wire _abc_19873_new_n3113_; 
wire _abc_19873_new_n3114_; 
wire _abc_19873_new_n3115_; 
wire _abc_19873_new_n3116_; 
wire _abc_19873_new_n3118_; 
wire _abc_19873_new_n3119_; 
wire _abc_19873_new_n3120_; 
wire _abc_19873_new_n3121_; 
wire _abc_19873_new_n3122_; 
wire _abc_19873_new_n3124_; 
wire _abc_19873_new_n3125_; 
wire _abc_19873_new_n3126_; 
wire _abc_19873_new_n3127_; 
wire _abc_19873_new_n3129_; 
wire _abc_19873_new_n3130_; 
wire _abc_19873_new_n3131_; 
wire _abc_19873_new_n3133_; 
wire _abc_19873_new_n3134_; 
wire _abc_19873_new_n3135_; 
wire _abc_19873_new_n3137_; 
wire _abc_19873_new_n3138_; 
wire _abc_19873_new_n3139_; 
wire _abc_19873_new_n3141_; 
wire _abc_19873_new_n3142_; 
wire _abc_19873_new_n3143_; 
wire _abc_19873_new_n3145_; 
wire _abc_19873_new_n3146_; 
wire _abc_19873_new_n3147_; 
wire _abc_19873_new_n3149_; 
wire _abc_19873_new_n3150_; 
wire _abc_19873_new_n3151_; 
wire _abc_19873_new_n3153_; 
wire _abc_19873_new_n3154_; 
wire _abc_19873_new_n3156_; 
wire _abc_19873_new_n3158_; 
wire _abc_19873_new_n3160_; 
wire _abc_19873_new_n3161_; 
wire _abc_19873_new_n3162_; 
wire _abc_19873_new_n3163_; 
wire _abc_19873_new_n3164_; 
wire _abc_19873_new_n3165_; 
wire _abc_19873_new_n3166_; 
wire _abc_19873_new_n870_; 
wire _abc_19873_new_n871_; 
wire _abc_19873_new_n872_; 
wire _abc_19873_new_n873_; 
wire _abc_19873_new_n874_; 
wire _abc_19873_new_n875_; 
wire _abc_19873_new_n876_; 
wire _abc_19873_new_n877_; 
wire _abc_19873_new_n878_; 
wire _abc_19873_new_n879_; 
wire _abc_19873_new_n880_; 
wire _abc_19873_new_n881_; 
wire _abc_19873_new_n882_; 
wire _abc_19873_new_n883_; 
wire _abc_19873_new_n884_; 
wire _abc_19873_new_n885_; 
wire _abc_19873_new_n886_; 
wire _abc_19873_new_n887_; 
wire _abc_19873_new_n888_; 
wire _abc_19873_new_n889_; 
wire _abc_19873_new_n890_; 
wire _abc_19873_new_n891_; 
wire _abc_19873_new_n892_; 
wire _abc_19873_new_n893_; 
wire _abc_19873_new_n894_; 
wire _abc_19873_new_n895_; 
wire _abc_19873_new_n896_; 
wire _abc_19873_new_n897_; 
wire _abc_19873_new_n898_; 
wire _abc_19873_new_n899_; 
wire _abc_19873_new_n900_; 
wire _abc_19873_new_n901_; 
wire _abc_19873_new_n902_; 
wire _abc_19873_new_n903_; 
wire _abc_19873_new_n904_; 
wire _abc_19873_new_n905_; 
wire _abc_19873_new_n906_; 
wire _abc_19873_new_n907_; 
wire _abc_19873_new_n908_; 
wire _abc_19873_new_n909_; 
wire _abc_19873_new_n910_; 
wire _abc_19873_new_n911_; 
wire _abc_19873_new_n912_; 
wire _abc_19873_new_n913_; 
wire _abc_19873_new_n914_; 
wire _abc_19873_new_n915_; 
wire _abc_19873_new_n916_; 
wire _abc_19873_new_n917_; 
wire _abc_19873_new_n918_; 
wire _abc_19873_new_n919_; 
wire _abc_19873_new_n920_; 
wire _abc_19873_new_n921_; 
wire _abc_19873_new_n922_; 
wire _abc_19873_new_n923_; 
wire _abc_19873_new_n924_; 
wire _abc_19873_new_n925_; 
wire _abc_19873_new_n926_; 
wire _abc_19873_new_n927_; 
wire _abc_19873_new_n928_; 
wire _abc_19873_new_n929_; 
wire _abc_19873_new_n930_; 
wire _abc_19873_new_n931_; 
wire _abc_19873_new_n932_; 
wire _abc_19873_new_n933_; 
wire _abc_19873_new_n934_; 
wire _abc_19873_new_n935_; 
wire _abc_19873_new_n936_; 
wire _abc_19873_new_n937_; 
wire _abc_19873_new_n939_; 
wire _abc_19873_new_n940_; 
wire _abc_19873_new_n941_; 
wire _abc_19873_new_n942_; 
wire _abc_19873_new_n943_; 
wire _abc_19873_new_n944_; 
wire _abc_19873_new_n945_; 
wire _abc_19873_new_n946_; 
wire _abc_19873_new_n947_; 
wire _abc_19873_new_n948_; 
wire _abc_19873_new_n949_; 
wire _abc_19873_new_n950_; 
wire _abc_19873_new_n951_; 
wire _abc_19873_new_n952_; 
wire _abc_19873_new_n953_; 
wire _abc_19873_new_n954_; 
wire _abc_19873_new_n955_; 
wire _abc_19873_new_n956_; 
wire _abc_19873_new_n957_; 
wire _abc_19873_new_n958_; 
wire _abc_19873_new_n959_; 
wire _abc_19873_new_n960_; 
wire _abc_19873_new_n961_; 
wire _abc_19873_new_n962_; 
wire _abc_19873_new_n963_; 
wire _abc_19873_new_n965_; 
wire _abc_19873_new_n966_; 
wire _abc_19873_new_n967_; 
wire _abc_19873_new_n968_; 
wire _abc_19873_new_n969_; 
wire _abc_19873_new_n970_; 
wire _abc_19873_new_n971_; 
wire _abc_19873_new_n972_; 
wire _abc_19873_new_n973_; 
wire _abc_19873_new_n974_; 
wire _abc_19873_new_n975_; 
wire _abc_19873_new_n976_; 
wire _abc_19873_new_n977_; 
wire _abc_19873_new_n978_; 
wire _abc_19873_new_n979_; 
wire _abc_19873_new_n980_; 
wire _abc_19873_new_n981_; 
wire _abc_19873_new_n982_; 
wire _abc_19873_new_n983_; 
wire _abc_19873_new_n984_; 
wire _abc_19873_new_n985_; 
wire _abc_19873_new_n986_; 
wire _abc_19873_new_n987_; 
wire _abc_19873_new_n989_; 
wire _abc_19873_new_n990_; 
wire _abc_19873_new_n991_; 
wire _abc_19873_new_n992_; 
wire _abc_19873_new_n993_; 
wire _abc_19873_new_n994_; 
wire _abc_19873_new_n995_; 
wire _abc_19873_new_n996_; 
wire _abc_19873_new_n997_; 
wire _abc_19873_new_n998_; 
wire _abc_19873_new_n999_; 
input \addr[0] ;
input \addr[1] ;
input \addr[2] ;
input \addr[3] ;
input \addr[4] ;
input \addr[5] ;
input \addr[6] ;
input \addr[7] ;
input clk;
wire core__0loop_ctr_reg_3_0__0_; 
wire core__0loop_ctr_reg_3_0__1_; 
wire core__0loop_ctr_reg_3_0__2_; 
wire core__0loop_ctr_reg_3_0__3_; 
wire core__0mi_reg_63_0__0_; 
wire core__0mi_reg_63_0__10_; 
wire core__0mi_reg_63_0__11_; 
wire core__0mi_reg_63_0__12_; 
wire core__0mi_reg_63_0__13_; 
wire core__0mi_reg_63_0__14_; 
wire core__0mi_reg_63_0__15_; 
wire core__0mi_reg_63_0__16_; 
wire core__0mi_reg_63_0__17_; 
wire core__0mi_reg_63_0__18_; 
wire core__0mi_reg_63_0__19_; 
wire core__0mi_reg_63_0__1_; 
wire core__0mi_reg_63_0__20_; 
wire core__0mi_reg_63_0__21_; 
wire core__0mi_reg_63_0__22_; 
wire core__0mi_reg_63_0__23_; 
wire core__0mi_reg_63_0__24_; 
wire core__0mi_reg_63_0__25_; 
wire core__0mi_reg_63_0__26_; 
wire core__0mi_reg_63_0__27_; 
wire core__0mi_reg_63_0__28_; 
wire core__0mi_reg_63_0__29_; 
wire core__0mi_reg_63_0__2_; 
wire core__0mi_reg_63_0__30_; 
wire core__0mi_reg_63_0__31_; 
wire core__0mi_reg_63_0__32_; 
wire core__0mi_reg_63_0__33_; 
wire core__0mi_reg_63_0__34_; 
wire core__0mi_reg_63_0__35_; 
wire core__0mi_reg_63_0__36_; 
wire core__0mi_reg_63_0__37_; 
wire core__0mi_reg_63_0__38_; 
wire core__0mi_reg_63_0__39_; 
wire core__0mi_reg_63_0__3_; 
wire core__0mi_reg_63_0__40_; 
wire core__0mi_reg_63_0__41_; 
wire core__0mi_reg_63_0__42_; 
wire core__0mi_reg_63_0__43_; 
wire core__0mi_reg_63_0__44_; 
wire core__0mi_reg_63_0__45_; 
wire core__0mi_reg_63_0__46_; 
wire core__0mi_reg_63_0__47_; 
wire core__0mi_reg_63_0__48_; 
wire core__0mi_reg_63_0__49_; 
wire core__0mi_reg_63_0__4_; 
wire core__0mi_reg_63_0__50_; 
wire core__0mi_reg_63_0__51_; 
wire core__0mi_reg_63_0__52_; 
wire core__0mi_reg_63_0__53_; 
wire core__0mi_reg_63_0__54_; 
wire core__0mi_reg_63_0__55_; 
wire core__0mi_reg_63_0__56_; 
wire core__0mi_reg_63_0__57_; 
wire core__0mi_reg_63_0__58_; 
wire core__0mi_reg_63_0__59_; 
wire core__0mi_reg_63_0__5_; 
wire core__0mi_reg_63_0__60_; 
wire core__0mi_reg_63_0__61_; 
wire core__0mi_reg_63_0__62_; 
wire core__0mi_reg_63_0__63_; 
wire core__0mi_reg_63_0__6_; 
wire core__0mi_reg_63_0__7_; 
wire core__0mi_reg_63_0__8_; 
wire core__0mi_reg_63_0__9_; 
wire core__0ready_reg_0_0_; 
wire core__0siphash_valid_reg_0_0_; 
wire core__0siphash_word0_reg_63_0__0_; 
wire core__0siphash_word0_reg_63_0__10_; 
wire core__0siphash_word0_reg_63_0__11_; 
wire core__0siphash_word0_reg_63_0__12_; 
wire core__0siphash_word0_reg_63_0__13_; 
wire core__0siphash_word0_reg_63_0__14_; 
wire core__0siphash_word0_reg_63_0__15_; 
wire core__0siphash_word0_reg_63_0__16_; 
wire core__0siphash_word0_reg_63_0__17_; 
wire core__0siphash_word0_reg_63_0__18_; 
wire core__0siphash_word0_reg_63_0__19_; 
wire core__0siphash_word0_reg_63_0__1_; 
wire core__0siphash_word0_reg_63_0__20_; 
wire core__0siphash_word0_reg_63_0__21_; 
wire core__0siphash_word0_reg_63_0__22_; 
wire core__0siphash_word0_reg_63_0__23_; 
wire core__0siphash_word0_reg_63_0__24_; 
wire core__0siphash_word0_reg_63_0__25_; 
wire core__0siphash_word0_reg_63_0__26_; 
wire core__0siphash_word0_reg_63_0__27_; 
wire core__0siphash_word0_reg_63_0__28_; 
wire core__0siphash_word0_reg_63_0__29_; 
wire core__0siphash_word0_reg_63_0__2_; 
wire core__0siphash_word0_reg_63_0__30_; 
wire core__0siphash_word0_reg_63_0__31_; 
wire core__0siphash_word0_reg_63_0__32_; 
wire core__0siphash_word0_reg_63_0__33_; 
wire core__0siphash_word0_reg_63_0__34_; 
wire core__0siphash_word0_reg_63_0__35_; 
wire core__0siphash_word0_reg_63_0__36_; 
wire core__0siphash_word0_reg_63_0__37_; 
wire core__0siphash_word0_reg_63_0__38_; 
wire core__0siphash_word0_reg_63_0__39_; 
wire core__0siphash_word0_reg_63_0__3_; 
wire core__0siphash_word0_reg_63_0__40_; 
wire core__0siphash_word0_reg_63_0__41_; 
wire core__0siphash_word0_reg_63_0__42_; 
wire core__0siphash_word0_reg_63_0__43_; 
wire core__0siphash_word0_reg_63_0__44_; 
wire core__0siphash_word0_reg_63_0__45_; 
wire core__0siphash_word0_reg_63_0__46_; 
wire core__0siphash_word0_reg_63_0__47_; 
wire core__0siphash_word0_reg_63_0__48_; 
wire core__0siphash_word0_reg_63_0__49_; 
wire core__0siphash_word0_reg_63_0__4_; 
wire core__0siphash_word0_reg_63_0__50_; 
wire core__0siphash_word0_reg_63_0__51_; 
wire core__0siphash_word0_reg_63_0__52_; 
wire core__0siphash_word0_reg_63_0__53_; 
wire core__0siphash_word0_reg_63_0__54_; 
wire core__0siphash_word0_reg_63_0__55_; 
wire core__0siphash_word0_reg_63_0__56_; 
wire core__0siphash_word0_reg_63_0__57_; 
wire core__0siphash_word0_reg_63_0__58_; 
wire core__0siphash_word0_reg_63_0__59_; 
wire core__0siphash_word0_reg_63_0__5_; 
wire core__0siphash_word0_reg_63_0__60_; 
wire core__0siphash_word0_reg_63_0__61_; 
wire core__0siphash_word0_reg_63_0__62_; 
wire core__0siphash_word0_reg_63_0__63_; 
wire core__0siphash_word0_reg_63_0__6_; 
wire core__0siphash_word0_reg_63_0__7_; 
wire core__0siphash_word0_reg_63_0__8_; 
wire core__0siphash_word0_reg_63_0__9_; 
wire core__0siphash_word1_reg_63_0__0_; 
wire core__0siphash_word1_reg_63_0__10_; 
wire core__0siphash_word1_reg_63_0__11_; 
wire core__0siphash_word1_reg_63_0__12_; 
wire core__0siphash_word1_reg_63_0__13_; 
wire core__0siphash_word1_reg_63_0__14_; 
wire core__0siphash_word1_reg_63_0__15_; 
wire core__0siphash_word1_reg_63_0__16_; 
wire core__0siphash_word1_reg_63_0__17_; 
wire core__0siphash_word1_reg_63_0__18_; 
wire core__0siphash_word1_reg_63_0__19_; 
wire core__0siphash_word1_reg_63_0__1_; 
wire core__0siphash_word1_reg_63_0__20_; 
wire core__0siphash_word1_reg_63_0__21_; 
wire core__0siphash_word1_reg_63_0__22_; 
wire core__0siphash_word1_reg_63_0__23_; 
wire core__0siphash_word1_reg_63_0__24_; 
wire core__0siphash_word1_reg_63_0__25_; 
wire core__0siphash_word1_reg_63_0__26_; 
wire core__0siphash_word1_reg_63_0__27_; 
wire core__0siphash_word1_reg_63_0__28_; 
wire core__0siphash_word1_reg_63_0__29_; 
wire core__0siphash_word1_reg_63_0__2_; 
wire core__0siphash_word1_reg_63_0__30_; 
wire core__0siphash_word1_reg_63_0__31_; 
wire core__0siphash_word1_reg_63_0__32_; 
wire core__0siphash_word1_reg_63_0__33_; 
wire core__0siphash_word1_reg_63_0__34_; 
wire core__0siphash_word1_reg_63_0__35_; 
wire core__0siphash_word1_reg_63_0__36_; 
wire core__0siphash_word1_reg_63_0__37_; 
wire core__0siphash_word1_reg_63_0__38_; 
wire core__0siphash_word1_reg_63_0__39_; 
wire core__0siphash_word1_reg_63_0__3_; 
wire core__0siphash_word1_reg_63_0__40_; 
wire core__0siphash_word1_reg_63_0__41_; 
wire core__0siphash_word1_reg_63_0__42_; 
wire core__0siphash_word1_reg_63_0__43_; 
wire core__0siphash_word1_reg_63_0__44_; 
wire core__0siphash_word1_reg_63_0__45_; 
wire core__0siphash_word1_reg_63_0__46_; 
wire core__0siphash_word1_reg_63_0__47_; 
wire core__0siphash_word1_reg_63_0__48_; 
wire core__0siphash_word1_reg_63_0__49_; 
wire core__0siphash_word1_reg_63_0__4_; 
wire core__0siphash_word1_reg_63_0__50_; 
wire core__0siphash_word1_reg_63_0__51_; 
wire core__0siphash_word1_reg_63_0__52_; 
wire core__0siphash_word1_reg_63_0__53_; 
wire core__0siphash_word1_reg_63_0__54_; 
wire core__0siphash_word1_reg_63_0__55_; 
wire core__0siphash_word1_reg_63_0__56_; 
wire core__0siphash_word1_reg_63_0__57_; 
wire core__0siphash_word1_reg_63_0__58_; 
wire core__0siphash_word1_reg_63_0__59_; 
wire core__0siphash_word1_reg_63_0__5_; 
wire core__0siphash_word1_reg_63_0__60_; 
wire core__0siphash_word1_reg_63_0__61_; 
wire core__0siphash_word1_reg_63_0__62_; 
wire core__0siphash_word1_reg_63_0__63_; 
wire core__0siphash_word1_reg_63_0__6_; 
wire core__0siphash_word1_reg_63_0__7_; 
wire core__0siphash_word1_reg_63_0__8_; 
wire core__0siphash_word1_reg_63_0__9_; 
wire core__0v0_reg_63_0__0_; 
wire core__0v0_reg_63_0__10_; 
wire core__0v0_reg_63_0__11_; 
wire core__0v0_reg_63_0__12_; 
wire core__0v0_reg_63_0__13_; 
wire core__0v0_reg_63_0__14_; 
wire core__0v0_reg_63_0__15_; 
wire core__0v0_reg_63_0__16_; 
wire core__0v0_reg_63_0__17_; 
wire core__0v0_reg_63_0__18_; 
wire core__0v0_reg_63_0__19_; 
wire core__0v0_reg_63_0__1_; 
wire core__0v0_reg_63_0__20_; 
wire core__0v0_reg_63_0__21_; 
wire core__0v0_reg_63_0__22_; 
wire core__0v0_reg_63_0__23_; 
wire core__0v0_reg_63_0__24_; 
wire core__0v0_reg_63_0__25_; 
wire core__0v0_reg_63_0__26_; 
wire core__0v0_reg_63_0__27_; 
wire core__0v0_reg_63_0__28_; 
wire core__0v0_reg_63_0__29_; 
wire core__0v0_reg_63_0__2_; 
wire core__0v0_reg_63_0__30_; 
wire core__0v0_reg_63_0__31_; 
wire core__0v0_reg_63_0__32_; 
wire core__0v0_reg_63_0__33_; 
wire core__0v0_reg_63_0__34_; 
wire core__0v0_reg_63_0__35_; 
wire core__0v0_reg_63_0__36_; 
wire core__0v0_reg_63_0__37_; 
wire core__0v0_reg_63_0__38_; 
wire core__0v0_reg_63_0__39_; 
wire core__0v0_reg_63_0__3_; 
wire core__0v0_reg_63_0__40_; 
wire core__0v0_reg_63_0__41_; 
wire core__0v0_reg_63_0__42_; 
wire core__0v0_reg_63_0__43_; 
wire core__0v0_reg_63_0__44_; 
wire core__0v0_reg_63_0__45_; 
wire core__0v0_reg_63_0__46_; 
wire core__0v0_reg_63_0__47_; 
wire core__0v0_reg_63_0__48_; 
wire core__0v0_reg_63_0__49_; 
wire core__0v0_reg_63_0__4_; 
wire core__0v0_reg_63_0__50_; 
wire core__0v0_reg_63_0__51_; 
wire core__0v0_reg_63_0__52_; 
wire core__0v0_reg_63_0__53_; 
wire core__0v0_reg_63_0__54_; 
wire core__0v0_reg_63_0__55_; 
wire core__0v0_reg_63_0__56_; 
wire core__0v0_reg_63_0__57_; 
wire core__0v0_reg_63_0__58_; 
wire core__0v0_reg_63_0__59_; 
wire core__0v0_reg_63_0__5_; 
wire core__0v0_reg_63_0__60_; 
wire core__0v0_reg_63_0__61_; 
wire core__0v0_reg_63_0__62_; 
wire core__0v0_reg_63_0__63_; 
wire core__0v0_reg_63_0__6_; 
wire core__0v0_reg_63_0__7_; 
wire core__0v0_reg_63_0__8_; 
wire core__0v0_reg_63_0__9_; 
wire core__0v1_reg_63_0__0_; 
wire core__0v1_reg_63_0__10_; 
wire core__0v1_reg_63_0__11_; 
wire core__0v1_reg_63_0__12_; 
wire core__0v1_reg_63_0__13_; 
wire core__0v1_reg_63_0__14_; 
wire core__0v1_reg_63_0__15_; 
wire core__0v1_reg_63_0__16_; 
wire core__0v1_reg_63_0__17_; 
wire core__0v1_reg_63_0__18_; 
wire core__0v1_reg_63_0__19_; 
wire core__0v1_reg_63_0__1_; 
wire core__0v1_reg_63_0__20_; 
wire core__0v1_reg_63_0__21_; 
wire core__0v1_reg_63_0__22_; 
wire core__0v1_reg_63_0__23_; 
wire core__0v1_reg_63_0__24_; 
wire core__0v1_reg_63_0__25_; 
wire core__0v1_reg_63_0__26_; 
wire core__0v1_reg_63_0__27_; 
wire core__0v1_reg_63_0__28_; 
wire core__0v1_reg_63_0__29_; 
wire core__0v1_reg_63_0__2_; 
wire core__0v1_reg_63_0__30_; 
wire core__0v1_reg_63_0__31_; 
wire core__0v1_reg_63_0__32_; 
wire core__0v1_reg_63_0__33_; 
wire core__0v1_reg_63_0__34_; 
wire core__0v1_reg_63_0__35_; 
wire core__0v1_reg_63_0__36_; 
wire core__0v1_reg_63_0__37_; 
wire core__0v1_reg_63_0__38_; 
wire core__0v1_reg_63_0__39_; 
wire core__0v1_reg_63_0__3_; 
wire core__0v1_reg_63_0__40_; 
wire core__0v1_reg_63_0__41_; 
wire core__0v1_reg_63_0__42_; 
wire core__0v1_reg_63_0__43_; 
wire core__0v1_reg_63_0__44_; 
wire core__0v1_reg_63_0__45_; 
wire core__0v1_reg_63_0__46_; 
wire core__0v1_reg_63_0__47_; 
wire core__0v1_reg_63_0__48_; 
wire core__0v1_reg_63_0__49_; 
wire core__0v1_reg_63_0__4_; 
wire core__0v1_reg_63_0__50_; 
wire core__0v1_reg_63_0__51_; 
wire core__0v1_reg_63_0__52_; 
wire core__0v1_reg_63_0__53_; 
wire core__0v1_reg_63_0__54_; 
wire core__0v1_reg_63_0__55_; 
wire core__0v1_reg_63_0__56_; 
wire core__0v1_reg_63_0__57_; 
wire core__0v1_reg_63_0__58_; 
wire core__0v1_reg_63_0__59_; 
wire core__0v1_reg_63_0__5_; 
wire core__0v1_reg_63_0__60_; 
wire core__0v1_reg_63_0__61_; 
wire core__0v1_reg_63_0__62_; 
wire core__0v1_reg_63_0__63_; 
wire core__0v1_reg_63_0__6_; 
wire core__0v1_reg_63_0__7_; 
wire core__0v1_reg_63_0__8_; 
wire core__0v1_reg_63_0__9_; 
wire core__0v2_reg_63_0__0_; 
wire core__0v2_reg_63_0__10_; 
wire core__0v2_reg_63_0__11_; 
wire core__0v2_reg_63_0__12_; 
wire core__0v2_reg_63_0__13_; 
wire core__0v2_reg_63_0__14_; 
wire core__0v2_reg_63_0__15_; 
wire core__0v2_reg_63_0__16_; 
wire core__0v2_reg_63_0__17_; 
wire core__0v2_reg_63_0__18_; 
wire core__0v2_reg_63_0__19_; 
wire core__0v2_reg_63_0__1_; 
wire core__0v2_reg_63_0__20_; 
wire core__0v2_reg_63_0__21_; 
wire core__0v2_reg_63_0__22_; 
wire core__0v2_reg_63_0__23_; 
wire core__0v2_reg_63_0__24_; 
wire core__0v2_reg_63_0__25_; 
wire core__0v2_reg_63_0__26_; 
wire core__0v2_reg_63_0__27_; 
wire core__0v2_reg_63_0__28_; 
wire core__0v2_reg_63_0__29_; 
wire core__0v2_reg_63_0__2_; 
wire core__0v2_reg_63_0__30_; 
wire core__0v2_reg_63_0__31_; 
wire core__0v2_reg_63_0__32_; 
wire core__0v2_reg_63_0__33_; 
wire core__0v2_reg_63_0__34_; 
wire core__0v2_reg_63_0__35_; 
wire core__0v2_reg_63_0__36_; 
wire core__0v2_reg_63_0__37_; 
wire core__0v2_reg_63_0__38_; 
wire core__0v2_reg_63_0__39_; 
wire core__0v2_reg_63_0__3_; 
wire core__0v2_reg_63_0__40_; 
wire core__0v2_reg_63_0__41_; 
wire core__0v2_reg_63_0__42_; 
wire core__0v2_reg_63_0__43_; 
wire core__0v2_reg_63_0__44_; 
wire core__0v2_reg_63_0__45_; 
wire core__0v2_reg_63_0__46_; 
wire core__0v2_reg_63_0__47_; 
wire core__0v2_reg_63_0__48_; 
wire core__0v2_reg_63_0__49_; 
wire core__0v2_reg_63_0__4_; 
wire core__0v2_reg_63_0__50_; 
wire core__0v2_reg_63_0__51_; 
wire core__0v2_reg_63_0__52_; 
wire core__0v2_reg_63_0__53_; 
wire core__0v2_reg_63_0__54_; 
wire core__0v2_reg_63_0__55_; 
wire core__0v2_reg_63_0__56_; 
wire core__0v2_reg_63_0__57_; 
wire core__0v2_reg_63_0__58_; 
wire core__0v2_reg_63_0__59_; 
wire core__0v2_reg_63_0__5_; 
wire core__0v2_reg_63_0__60_; 
wire core__0v2_reg_63_0__61_; 
wire core__0v2_reg_63_0__62_; 
wire core__0v2_reg_63_0__63_; 
wire core__0v2_reg_63_0__6_; 
wire core__0v2_reg_63_0__7_; 
wire core__0v2_reg_63_0__8_; 
wire core__0v2_reg_63_0__9_; 
wire core__0v3_reg_63_0__0_; 
wire core__0v3_reg_63_0__10_; 
wire core__0v3_reg_63_0__11_; 
wire core__0v3_reg_63_0__12_; 
wire core__0v3_reg_63_0__13_; 
wire core__0v3_reg_63_0__14_; 
wire core__0v3_reg_63_0__15_; 
wire core__0v3_reg_63_0__16_; 
wire core__0v3_reg_63_0__17_; 
wire core__0v3_reg_63_0__18_; 
wire core__0v3_reg_63_0__19_; 
wire core__0v3_reg_63_0__1_; 
wire core__0v3_reg_63_0__20_; 
wire core__0v3_reg_63_0__21_; 
wire core__0v3_reg_63_0__22_; 
wire core__0v3_reg_63_0__23_; 
wire core__0v3_reg_63_0__24_; 
wire core__0v3_reg_63_0__25_; 
wire core__0v3_reg_63_0__26_; 
wire core__0v3_reg_63_0__27_; 
wire core__0v3_reg_63_0__28_; 
wire core__0v3_reg_63_0__29_; 
wire core__0v3_reg_63_0__2_; 
wire core__0v3_reg_63_0__30_; 
wire core__0v3_reg_63_0__31_; 
wire core__0v3_reg_63_0__32_; 
wire core__0v3_reg_63_0__33_; 
wire core__0v3_reg_63_0__34_; 
wire core__0v3_reg_63_0__35_; 
wire core__0v3_reg_63_0__36_; 
wire core__0v3_reg_63_0__37_; 
wire core__0v3_reg_63_0__38_; 
wire core__0v3_reg_63_0__39_; 
wire core__0v3_reg_63_0__3_; 
wire core__0v3_reg_63_0__40_; 
wire core__0v3_reg_63_0__41_; 
wire core__0v3_reg_63_0__42_; 
wire core__0v3_reg_63_0__43_; 
wire core__0v3_reg_63_0__44_; 
wire core__0v3_reg_63_0__45_; 
wire core__0v3_reg_63_0__46_; 
wire core__0v3_reg_63_0__47_; 
wire core__0v3_reg_63_0__48_; 
wire core__0v3_reg_63_0__49_; 
wire core__0v3_reg_63_0__4_; 
wire core__0v3_reg_63_0__50_; 
wire core__0v3_reg_63_0__51_; 
wire core__0v3_reg_63_0__52_; 
wire core__0v3_reg_63_0__53_; 
wire core__0v3_reg_63_0__54_; 
wire core__0v3_reg_63_0__55_; 
wire core__0v3_reg_63_0__56_; 
wire core__0v3_reg_63_0__57_; 
wire core__0v3_reg_63_0__58_; 
wire core__0v3_reg_63_0__59_; 
wire core__0v3_reg_63_0__5_; 
wire core__0v3_reg_63_0__60_; 
wire core__0v3_reg_63_0__61_; 
wire core__0v3_reg_63_0__62_; 
wire core__0v3_reg_63_0__63_; 
wire core__0v3_reg_63_0__6_; 
wire core__0v3_reg_63_0__7_; 
wire core__0v3_reg_63_0__8_; 
wire core__0v3_reg_63_0__9_; 
wire core__abc_15204_auto_fsm_map_cc_118_implement_pattern_cache_1470; 
wire core__abc_15204_auto_fsm_map_cc_118_implement_pattern_cache_1474; 
wire core__abc_15204_auto_fsm_map_cc_118_implement_pattern_cache_1496; 
wire core__abc_15204_auto_fsm_map_cc_118_implement_pattern_cache_1509; 
wire core__abc_15204_auto_fsm_map_cc_170_map_fsm_1439_0_; 
wire core__abc_15204_auto_fsm_map_cc_170_map_fsm_1439_3_; 
wire core__abc_15204_auto_fsm_map_cc_170_map_fsm_1439_4_; 
wire core__abc_15204_auto_fsm_map_cc_170_map_fsm_1439_6_; 
wire core__abc_22172_new_n1130_; 
wire core__abc_22172_new_n1131_; 
wire core__abc_22172_new_n1132_; 
wire core__abc_22172_new_n1133_; 
wire core__abc_22172_new_n1134_; 
wire core__abc_22172_new_n1135_; 
wire core__abc_22172_new_n1136_; 
wire core__abc_22172_new_n1137_; 
wire core__abc_22172_new_n1138_; 
wire core__abc_22172_new_n1139_; 
wire core__abc_22172_new_n1140_; 
wire core__abc_22172_new_n1141_; 
wire core__abc_22172_new_n1142_; 
wire core__abc_22172_new_n1143_; 
wire core__abc_22172_new_n1144_; 
wire core__abc_22172_new_n1145_; 
wire core__abc_22172_new_n1146_; 
wire core__abc_22172_new_n1147_; 
wire core__abc_22172_new_n1148_; 
wire core__abc_22172_new_n1149_; 
wire core__abc_22172_new_n1150_; 
wire core__abc_22172_new_n1151_; 
wire core__abc_22172_new_n1152_; 
wire core__abc_22172_new_n1153_; 
wire core__abc_22172_new_n1154_; 
wire core__abc_22172_new_n1155_; 
wire core__abc_22172_new_n1156_; 
wire core__abc_22172_new_n1157_; 
wire core__abc_22172_new_n1158_; 
wire core__abc_22172_new_n1159_; 
wire core__abc_22172_new_n1160_; 
wire core__abc_22172_new_n1161_; 
wire core__abc_22172_new_n1162_; 
wire core__abc_22172_new_n1163_; 
wire core__abc_22172_new_n1164_; 
wire core__abc_22172_new_n1165_; 
wire core__abc_22172_new_n1166_; 
wire core__abc_22172_new_n1167_; 
wire core__abc_22172_new_n1168_; 
wire core__abc_22172_new_n1169_; 
wire core__abc_22172_new_n1170_; 
wire core__abc_22172_new_n1171_; 
wire core__abc_22172_new_n1172_; 
wire core__abc_22172_new_n1173_; 
wire core__abc_22172_new_n1174_; 
wire core__abc_22172_new_n1175_; 
wire core__abc_22172_new_n1176_; 
wire core__abc_22172_new_n1177_; 
wire core__abc_22172_new_n1178_; 
wire core__abc_22172_new_n1179_; 
wire core__abc_22172_new_n1180_; 
wire core__abc_22172_new_n1181_; 
wire core__abc_22172_new_n1182_; 
wire core__abc_22172_new_n1183_; 
wire core__abc_22172_new_n1184_; 
wire core__abc_22172_new_n1185_; 
wire core__abc_22172_new_n1186_; 
wire core__abc_22172_new_n1187_; 
wire core__abc_22172_new_n1188_; 
wire core__abc_22172_new_n1189_; 
wire core__abc_22172_new_n1190_; 
wire core__abc_22172_new_n1191_; 
wire core__abc_22172_new_n1192_; 
wire core__abc_22172_new_n1193_; 
wire core__abc_22172_new_n1194_; 
wire core__abc_22172_new_n1195_; 
wire core__abc_22172_new_n1196_; 
wire core__abc_22172_new_n1197_; 
wire core__abc_22172_new_n1198_; 
wire core__abc_22172_new_n1199_; 
wire core__abc_22172_new_n1200_; 
wire core__abc_22172_new_n1201_; 
wire core__abc_22172_new_n1202_; 
wire core__abc_22172_new_n1203_; 
wire core__abc_22172_new_n1204_; 
wire core__abc_22172_new_n1205_; 
wire core__abc_22172_new_n1206_; 
wire core__abc_22172_new_n1207_; 
wire core__abc_22172_new_n1208_; 
wire core__abc_22172_new_n1209_; 
wire core__abc_22172_new_n1210_; 
wire core__abc_22172_new_n1211_; 
wire core__abc_22172_new_n1212_; 
wire core__abc_22172_new_n1213_; 
wire core__abc_22172_new_n1214_; 
wire core__abc_22172_new_n1215_; 
wire core__abc_22172_new_n1216_; 
wire core__abc_22172_new_n1217_; 
wire core__abc_22172_new_n1218_; 
wire core__abc_22172_new_n1219_; 
wire core__abc_22172_new_n1220_; 
wire core__abc_22172_new_n1221_; 
wire core__abc_22172_new_n1222_; 
wire core__abc_22172_new_n1223_; 
wire core__abc_22172_new_n1224_; 
wire core__abc_22172_new_n1225_; 
wire core__abc_22172_new_n1226_; 
wire core__abc_22172_new_n1227_; 
wire core__abc_22172_new_n1228_; 
wire core__abc_22172_new_n1229_; 
wire core__abc_22172_new_n1230_; 
wire core__abc_22172_new_n1231_; 
wire core__abc_22172_new_n1232_; 
wire core__abc_22172_new_n1233_; 
wire core__abc_22172_new_n1234_; 
wire core__abc_22172_new_n1235_; 
wire core__abc_22172_new_n1236_; 
wire core__abc_22172_new_n1237_; 
wire core__abc_22172_new_n1238_; 
wire core__abc_22172_new_n1239_; 
wire core__abc_22172_new_n1240_; 
wire core__abc_22172_new_n1241_; 
wire core__abc_22172_new_n1243_; 
wire core__abc_22172_new_n1244_; 
wire core__abc_22172_new_n1245_; 
wire core__abc_22172_new_n1247_; 
wire core__abc_22172_new_n1248_; 
wire core__abc_22172_new_n1249_; 
wire core__abc_22172_new_n1251_; 
wire core__abc_22172_new_n1252_; 
wire core__abc_22172_new_n1253_; 
wire core__abc_22172_new_n1254_; 
wire core__abc_22172_new_n1256_; 
wire core__abc_22172_new_n1257_; 
wire core__abc_22172_new_n1258_; 
wire core__abc_22172_new_n1259_; 
wire core__abc_22172_new_n1260_; 
wire core__abc_22172_new_n1261_; 
wire core__abc_22172_new_n1262_; 
wire core__abc_22172_new_n1263_; 
wire core__abc_22172_new_n1264_; 
wire core__abc_22172_new_n1265_; 
wire core__abc_22172_new_n1266_; 
wire core__abc_22172_new_n1267_; 
wire core__abc_22172_new_n1268_; 
wire core__abc_22172_new_n1269_; 
wire core__abc_22172_new_n1270_; 
wire core__abc_22172_new_n1271_; 
wire core__abc_22172_new_n1272_; 
wire core__abc_22172_new_n1273_; 
wire core__abc_22172_new_n1275_; 
wire core__abc_22172_new_n1276_; 
wire core__abc_22172_new_n1277_; 
wire core__abc_22172_new_n1278_; 
wire core__abc_22172_new_n1279_; 
wire core__abc_22172_new_n1280_; 
wire core__abc_22172_new_n1281_; 
wire core__abc_22172_new_n1282_; 
wire core__abc_22172_new_n1283_; 
wire core__abc_22172_new_n1284_; 
wire core__abc_22172_new_n1285_; 
wire core__abc_22172_new_n1286_; 
wire core__abc_22172_new_n1287_; 
wire core__abc_22172_new_n1288_; 
wire core__abc_22172_new_n1289_; 
wire core__abc_22172_new_n1290_; 
wire core__abc_22172_new_n1291_; 
wire core__abc_22172_new_n1292_; 
wire core__abc_22172_new_n1293_; 
wire core__abc_22172_new_n1294_; 
wire core__abc_22172_new_n1296_; 
wire core__abc_22172_new_n1297_; 
wire core__abc_22172_new_n1298_; 
wire core__abc_22172_new_n1299_; 
wire core__abc_22172_new_n1300_; 
wire core__abc_22172_new_n1301_; 
wire core__abc_22172_new_n1302_; 
wire core__abc_22172_new_n1303_; 
wire core__abc_22172_new_n1304_; 
wire core__abc_22172_new_n1305_; 
wire core__abc_22172_new_n1306_; 
wire core__abc_22172_new_n1307_; 
wire core__abc_22172_new_n1308_; 
wire core__abc_22172_new_n1309_; 
wire core__abc_22172_new_n1310_; 
wire core__abc_22172_new_n1311_; 
wire core__abc_22172_new_n1312_; 
wire core__abc_22172_new_n1314_; 
wire core__abc_22172_new_n1315_; 
wire core__abc_22172_new_n1316_; 
wire core__abc_22172_new_n1317_; 
wire core__abc_22172_new_n1318_; 
wire core__abc_22172_new_n1319_; 
wire core__abc_22172_new_n1320_; 
wire core__abc_22172_new_n1321_; 
wire core__abc_22172_new_n1322_; 
wire core__abc_22172_new_n1323_; 
wire core__abc_22172_new_n1324_; 
wire core__abc_22172_new_n1325_; 
wire core__abc_22172_new_n1326_; 
wire core__abc_22172_new_n1327_; 
wire core__abc_22172_new_n1328_; 
wire core__abc_22172_new_n1329_; 
wire core__abc_22172_new_n1330_; 
wire core__abc_22172_new_n1332_; 
wire core__abc_22172_new_n1333_; 
wire core__abc_22172_new_n1334_; 
wire core__abc_22172_new_n1335_; 
wire core__abc_22172_new_n1336_; 
wire core__abc_22172_new_n1337_; 
wire core__abc_22172_new_n1338_; 
wire core__abc_22172_new_n1339_; 
wire core__abc_22172_new_n1340_; 
wire core__abc_22172_new_n1341_; 
wire core__abc_22172_new_n1342_; 
wire core__abc_22172_new_n1343_; 
wire core__abc_22172_new_n1344_; 
wire core__abc_22172_new_n1345_; 
wire core__abc_22172_new_n1346_; 
wire core__abc_22172_new_n1347_; 
wire core__abc_22172_new_n1348_; 
wire core__abc_22172_new_n1350_; 
wire core__abc_22172_new_n1351_; 
wire core__abc_22172_new_n1352_; 
wire core__abc_22172_new_n1353_; 
wire core__abc_22172_new_n1354_; 
wire core__abc_22172_new_n1355_; 
wire core__abc_22172_new_n1356_; 
wire core__abc_22172_new_n1357_; 
wire core__abc_22172_new_n1358_; 
wire core__abc_22172_new_n1359_; 
wire core__abc_22172_new_n1360_; 
wire core__abc_22172_new_n1361_; 
wire core__abc_22172_new_n1362_; 
wire core__abc_22172_new_n1363_; 
wire core__abc_22172_new_n1364_; 
wire core__abc_22172_new_n1365_; 
wire core__abc_22172_new_n1366_; 
wire core__abc_22172_new_n1367_; 
wire core__abc_22172_new_n1368_; 
wire core__abc_22172_new_n1370_; 
wire core__abc_22172_new_n1371_; 
wire core__abc_22172_new_n1372_; 
wire core__abc_22172_new_n1373_; 
wire core__abc_22172_new_n1374_; 
wire core__abc_22172_new_n1375_; 
wire core__abc_22172_new_n1376_; 
wire core__abc_22172_new_n1377_; 
wire core__abc_22172_new_n1378_; 
wire core__abc_22172_new_n1379_; 
wire core__abc_22172_new_n1380_; 
wire core__abc_22172_new_n1381_; 
wire core__abc_22172_new_n1382_; 
wire core__abc_22172_new_n1383_; 
wire core__abc_22172_new_n1384_; 
wire core__abc_22172_new_n1385_; 
wire core__abc_22172_new_n1386_; 
wire core__abc_22172_new_n1388_; 
wire core__abc_22172_new_n1389_; 
wire core__abc_22172_new_n1390_; 
wire core__abc_22172_new_n1391_; 
wire core__abc_22172_new_n1392_; 
wire core__abc_22172_new_n1393_; 
wire core__abc_22172_new_n1394_; 
wire core__abc_22172_new_n1395_; 
wire core__abc_22172_new_n1396_; 
wire core__abc_22172_new_n1397_; 
wire core__abc_22172_new_n1398_; 
wire core__abc_22172_new_n1399_; 
wire core__abc_22172_new_n1400_; 
wire core__abc_22172_new_n1401_; 
wire core__abc_22172_new_n1402_; 
wire core__abc_22172_new_n1403_; 
wire core__abc_22172_new_n1404_; 
wire core__abc_22172_new_n1405_; 
wire core__abc_22172_new_n1406_; 
wire core__abc_22172_new_n1408_; 
wire core__abc_22172_new_n1409_; 
wire core__abc_22172_new_n1410_; 
wire core__abc_22172_new_n1411_; 
wire core__abc_22172_new_n1412_; 
wire core__abc_22172_new_n1413_; 
wire core__abc_22172_new_n1414_; 
wire core__abc_22172_new_n1415_; 
wire core__abc_22172_new_n1416_; 
wire core__abc_22172_new_n1417_; 
wire core__abc_22172_new_n1418_; 
wire core__abc_22172_new_n1419_; 
wire core__abc_22172_new_n1420_; 
wire core__abc_22172_new_n1421_; 
wire core__abc_22172_new_n1422_; 
wire core__abc_22172_new_n1423_; 
wire core__abc_22172_new_n1425_; 
wire core__abc_22172_new_n1426_; 
wire core__abc_22172_new_n1427_; 
wire core__abc_22172_new_n1428_; 
wire core__abc_22172_new_n1429_; 
wire core__abc_22172_new_n1430_; 
wire core__abc_22172_new_n1431_; 
wire core__abc_22172_new_n1432_; 
wire core__abc_22172_new_n1433_; 
wire core__abc_22172_new_n1434_; 
wire core__abc_22172_new_n1435_; 
wire core__abc_22172_new_n1436_; 
wire core__abc_22172_new_n1437_; 
wire core__abc_22172_new_n1438_; 
wire core__abc_22172_new_n1439_; 
wire core__abc_22172_new_n1440_; 
wire core__abc_22172_new_n1442_; 
wire core__abc_22172_new_n1443_; 
wire core__abc_22172_new_n1444_; 
wire core__abc_22172_new_n1445_; 
wire core__abc_22172_new_n1446_; 
wire core__abc_22172_new_n1447_; 
wire core__abc_22172_new_n1448_; 
wire core__abc_22172_new_n1449_; 
wire core__abc_22172_new_n1450_; 
wire core__abc_22172_new_n1451_; 
wire core__abc_22172_new_n1452_; 
wire core__abc_22172_new_n1453_; 
wire core__abc_22172_new_n1454_; 
wire core__abc_22172_new_n1455_; 
wire core__abc_22172_new_n1456_; 
wire core__abc_22172_new_n1457_; 
wire core__abc_22172_new_n1459_; 
wire core__abc_22172_new_n1460_; 
wire core__abc_22172_new_n1461_; 
wire core__abc_22172_new_n1462_; 
wire core__abc_22172_new_n1463_; 
wire core__abc_22172_new_n1464_; 
wire core__abc_22172_new_n1465_; 
wire core__abc_22172_new_n1466_; 
wire core__abc_22172_new_n1467_; 
wire core__abc_22172_new_n1468_; 
wire core__abc_22172_new_n1469_; 
wire core__abc_22172_new_n1470_; 
wire core__abc_22172_new_n1471_; 
wire core__abc_22172_new_n1472_; 
wire core__abc_22172_new_n1473_; 
wire core__abc_22172_new_n1474_; 
wire core__abc_22172_new_n1476_; 
wire core__abc_22172_new_n1477_; 
wire core__abc_22172_new_n1478_; 
wire core__abc_22172_new_n1479_; 
wire core__abc_22172_new_n1480_; 
wire core__abc_22172_new_n1481_; 
wire core__abc_22172_new_n1482_; 
wire core__abc_22172_new_n1483_; 
wire core__abc_22172_new_n1484_; 
wire core__abc_22172_new_n1485_; 
wire core__abc_22172_new_n1486_; 
wire core__abc_22172_new_n1487_; 
wire core__abc_22172_new_n1488_; 
wire core__abc_22172_new_n1489_; 
wire core__abc_22172_new_n1490_; 
wire core__abc_22172_new_n1491_; 
wire core__abc_22172_new_n1493_; 
wire core__abc_22172_new_n1494_; 
wire core__abc_22172_new_n1495_; 
wire core__abc_22172_new_n1496_; 
wire core__abc_22172_new_n1497_; 
wire core__abc_22172_new_n1498_; 
wire core__abc_22172_new_n1499_; 
wire core__abc_22172_new_n1500_; 
wire core__abc_22172_new_n1501_; 
wire core__abc_22172_new_n1502_; 
wire core__abc_22172_new_n1503_; 
wire core__abc_22172_new_n1504_; 
wire core__abc_22172_new_n1505_; 
wire core__abc_22172_new_n1506_; 
wire core__abc_22172_new_n1507_; 
wire core__abc_22172_new_n1508_; 
wire core__abc_22172_new_n1510_; 
wire core__abc_22172_new_n1511_; 
wire core__abc_22172_new_n1512_; 
wire core__abc_22172_new_n1513_; 
wire core__abc_22172_new_n1514_; 
wire core__abc_22172_new_n1515_; 
wire core__abc_22172_new_n1516_; 
wire core__abc_22172_new_n1517_; 
wire core__abc_22172_new_n1518_; 
wire core__abc_22172_new_n1519_; 
wire core__abc_22172_new_n1520_; 
wire core__abc_22172_new_n1521_; 
wire core__abc_22172_new_n1522_; 
wire core__abc_22172_new_n1523_; 
wire core__abc_22172_new_n1524_; 
wire core__abc_22172_new_n1525_; 
wire core__abc_22172_new_n1527_; 
wire core__abc_22172_new_n1528_; 
wire core__abc_22172_new_n1529_; 
wire core__abc_22172_new_n1530_; 
wire core__abc_22172_new_n1531_; 
wire core__abc_22172_new_n1532_; 
wire core__abc_22172_new_n1533_; 
wire core__abc_22172_new_n1534_; 
wire core__abc_22172_new_n1535_; 
wire core__abc_22172_new_n1536_; 
wire core__abc_22172_new_n1537_; 
wire core__abc_22172_new_n1538_; 
wire core__abc_22172_new_n1539_; 
wire core__abc_22172_new_n1540_; 
wire core__abc_22172_new_n1541_; 
wire core__abc_22172_new_n1542_; 
wire core__abc_22172_new_n1544_; 
wire core__abc_22172_new_n1545_; 
wire core__abc_22172_new_n1546_; 
wire core__abc_22172_new_n1547_; 
wire core__abc_22172_new_n1548_; 
wire core__abc_22172_new_n1549_; 
wire core__abc_22172_new_n1550_; 
wire core__abc_22172_new_n1551_; 
wire core__abc_22172_new_n1552_; 
wire core__abc_22172_new_n1553_; 
wire core__abc_22172_new_n1554_; 
wire core__abc_22172_new_n1555_; 
wire core__abc_22172_new_n1556_; 
wire core__abc_22172_new_n1557_; 
wire core__abc_22172_new_n1558_; 
wire core__abc_22172_new_n1559_; 
wire core__abc_22172_new_n1561_; 
wire core__abc_22172_new_n1562_; 
wire core__abc_22172_new_n1563_; 
wire core__abc_22172_new_n1564_; 
wire core__abc_22172_new_n1565_; 
wire core__abc_22172_new_n1566_; 
wire core__abc_22172_new_n1567_; 
wire core__abc_22172_new_n1568_; 
wire core__abc_22172_new_n1569_; 
wire core__abc_22172_new_n1570_; 
wire core__abc_22172_new_n1571_; 
wire core__abc_22172_new_n1572_; 
wire core__abc_22172_new_n1573_; 
wire core__abc_22172_new_n1574_; 
wire core__abc_22172_new_n1575_; 
wire core__abc_22172_new_n1576_; 
wire core__abc_22172_new_n1578_; 
wire core__abc_22172_new_n1579_; 
wire core__abc_22172_new_n1580_; 
wire core__abc_22172_new_n1581_; 
wire core__abc_22172_new_n1582_; 
wire core__abc_22172_new_n1583_; 
wire core__abc_22172_new_n1584_; 
wire core__abc_22172_new_n1585_; 
wire core__abc_22172_new_n1586_; 
wire core__abc_22172_new_n1587_; 
wire core__abc_22172_new_n1588_; 
wire core__abc_22172_new_n1589_; 
wire core__abc_22172_new_n1590_; 
wire core__abc_22172_new_n1591_; 
wire core__abc_22172_new_n1592_; 
wire core__abc_22172_new_n1593_; 
wire core__abc_22172_new_n1595_; 
wire core__abc_22172_new_n1596_; 
wire core__abc_22172_new_n1597_; 
wire core__abc_22172_new_n1598_; 
wire core__abc_22172_new_n1599_; 
wire core__abc_22172_new_n1600_; 
wire core__abc_22172_new_n1601_; 
wire core__abc_22172_new_n1602_; 
wire core__abc_22172_new_n1603_; 
wire core__abc_22172_new_n1604_; 
wire core__abc_22172_new_n1605_; 
wire core__abc_22172_new_n1606_; 
wire core__abc_22172_new_n1607_; 
wire core__abc_22172_new_n1608_; 
wire core__abc_22172_new_n1609_; 
wire core__abc_22172_new_n1610_; 
wire core__abc_22172_new_n1612_; 
wire core__abc_22172_new_n1613_; 
wire core__abc_22172_new_n1614_; 
wire core__abc_22172_new_n1615_; 
wire core__abc_22172_new_n1616_; 
wire core__abc_22172_new_n1617_; 
wire core__abc_22172_new_n1618_; 
wire core__abc_22172_new_n1619_; 
wire core__abc_22172_new_n1620_; 
wire core__abc_22172_new_n1621_; 
wire core__abc_22172_new_n1622_; 
wire core__abc_22172_new_n1623_; 
wire core__abc_22172_new_n1624_; 
wire core__abc_22172_new_n1625_; 
wire core__abc_22172_new_n1626_; 
wire core__abc_22172_new_n1627_; 
wire core__abc_22172_new_n1629_; 
wire core__abc_22172_new_n1630_; 
wire core__abc_22172_new_n1631_; 
wire core__abc_22172_new_n1632_; 
wire core__abc_22172_new_n1633_; 
wire core__abc_22172_new_n1634_; 
wire core__abc_22172_new_n1635_; 
wire core__abc_22172_new_n1636_; 
wire core__abc_22172_new_n1637_; 
wire core__abc_22172_new_n1638_; 
wire core__abc_22172_new_n1639_; 
wire core__abc_22172_new_n1640_; 
wire core__abc_22172_new_n1641_; 
wire core__abc_22172_new_n1642_; 
wire core__abc_22172_new_n1643_; 
wire core__abc_22172_new_n1644_; 
wire core__abc_22172_new_n1646_; 
wire core__abc_22172_new_n1647_; 
wire core__abc_22172_new_n1648_; 
wire core__abc_22172_new_n1649_; 
wire core__abc_22172_new_n1650_; 
wire core__abc_22172_new_n1651_; 
wire core__abc_22172_new_n1652_; 
wire core__abc_22172_new_n1653_; 
wire core__abc_22172_new_n1654_; 
wire core__abc_22172_new_n1655_; 
wire core__abc_22172_new_n1656_; 
wire core__abc_22172_new_n1657_; 
wire core__abc_22172_new_n1658_; 
wire core__abc_22172_new_n1659_; 
wire core__abc_22172_new_n1660_; 
wire core__abc_22172_new_n1661_; 
wire core__abc_22172_new_n1663_; 
wire core__abc_22172_new_n1664_; 
wire core__abc_22172_new_n1665_; 
wire core__abc_22172_new_n1666_; 
wire core__abc_22172_new_n1667_; 
wire core__abc_22172_new_n1668_; 
wire core__abc_22172_new_n1669_; 
wire core__abc_22172_new_n1670_; 
wire core__abc_22172_new_n1671_; 
wire core__abc_22172_new_n1672_; 
wire core__abc_22172_new_n1673_; 
wire core__abc_22172_new_n1674_; 
wire core__abc_22172_new_n1675_; 
wire core__abc_22172_new_n1676_; 
wire core__abc_22172_new_n1677_; 
wire core__abc_22172_new_n1678_; 
wire core__abc_22172_new_n1680_; 
wire core__abc_22172_new_n1681_; 
wire core__abc_22172_new_n1682_; 
wire core__abc_22172_new_n1683_; 
wire core__abc_22172_new_n1684_; 
wire core__abc_22172_new_n1685_; 
wire core__abc_22172_new_n1686_; 
wire core__abc_22172_new_n1687_; 
wire core__abc_22172_new_n1688_; 
wire core__abc_22172_new_n1689_; 
wire core__abc_22172_new_n1690_; 
wire core__abc_22172_new_n1691_; 
wire core__abc_22172_new_n1692_; 
wire core__abc_22172_new_n1693_; 
wire core__abc_22172_new_n1694_; 
wire core__abc_22172_new_n1695_; 
wire core__abc_22172_new_n1697_; 
wire core__abc_22172_new_n1698_; 
wire core__abc_22172_new_n1699_; 
wire core__abc_22172_new_n1700_; 
wire core__abc_22172_new_n1701_; 
wire core__abc_22172_new_n1702_; 
wire core__abc_22172_new_n1703_; 
wire core__abc_22172_new_n1704_; 
wire core__abc_22172_new_n1705_; 
wire core__abc_22172_new_n1706_; 
wire core__abc_22172_new_n1707_; 
wire core__abc_22172_new_n1708_; 
wire core__abc_22172_new_n1709_; 
wire core__abc_22172_new_n1710_; 
wire core__abc_22172_new_n1711_; 
wire core__abc_22172_new_n1712_; 
wire core__abc_22172_new_n1714_; 
wire core__abc_22172_new_n1715_; 
wire core__abc_22172_new_n1716_; 
wire core__abc_22172_new_n1717_; 
wire core__abc_22172_new_n1718_; 
wire core__abc_22172_new_n1719_; 
wire core__abc_22172_new_n1720_; 
wire core__abc_22172_new_n1721_; 
wire core__abc_22172_new_n1722_; 
wire core__abc_22172_new_n1723_; 
wire core__abc_22172_new_n1724_; 
wire core__abc_22172_new_n1725_; 
wire core__abc_22172_new_n1726_; 
wire core__abc_22172_new_n1727_; 
wire core__abc_22172_new_n1728_; 
wire core__abc_22172_new_n1729_; 
wire core__abc_22172_new_n1731_; 
wire core__abc_22172_new_n1732_; 
wire core__abc_22172_new_n1733_; 
wire core__abc_22172_new_n1734_; 
wire core__abc_22172_new_n1735_; 
wire core__abc_22172_new_n1736_; 
wire core__abc_22172_new_n1737_; 
wire core__abc_22172_new_n1738_; 
wire core__abc_22172_new_n1739_; 
wire core__abc_22172_new_n1740_; 
wire core__abc_22172_new_n1741_; 
wire core__abc_22172_new_n1742_; 
wire core__abc_22172_new_n1743_; 
wire core__abc_22172_new_n1744_; 
wire core__abc_22172_new_n1745_; 
wire core__abc_22172_new_n1746_; 
wire core__abc_22172_new_n1748_; 
wire core__abc_22172_new_n1749_; 
wire core__abc_22172_new_n1750_; 
wire core__abc_22172_new_n1751_; 
wire core__abc_22172_new_n1752_; 
wire core__abc_22172_new_n1753_; 
wire core__abc_22172_new_n1754_; 
wire core__abc_22172_new_n1755_; 
wire core__abc_22172_new_n1756_; 
wire core__abc_22172_new_n1757_; 
wire core__abc_22172_new_n1758_; 
wire core__abc_22172_new_n1759_; 
wire core__abc_22172_new_n1760_; 
wire core__abc_22172_new_n1761_; 
wire core__abc_22172_new_n1762_; 
wire core__abc_22172_new_n1763_; 
wire core__abc_22172_new_n1765_; 
wire core__abc_22172_new_n1766_; 
wire core__abc_22172_new_n1767_; 
wire core__abc_22172_new_n1768_; 
wire core__abc_22172_new_n1769_; 
wire core__abc_22172_new_n1770_; 
wire core__abc_22172_new_n1771_; 
wire core__abc_22172_new_n1772_; 
wire core__abc_22172_new_n1773_; 
wire core__abc_22172_new_n1774_; 
wire core__abc_22172_new_n1775_; 
wire core__abc_22172_new_n1776_; 
wire core__abc_22172_new_n1777_; 
wire core__abc_22172_new_n1778_; 
wire core__abc_22172_new_n1779_; 
wire core__abc_22172_new_n1780_; 
wire core__abc_22172_new_n1782_; 
wire core__abc_22172_new_n1783_; 
wire core__abc_22172_new_n1784_; 
wire core__abc_22172_new_n1785_; 
wire core__abc_22172_new_n1786_; 
wire core__abc_22172_new_n1787_; 
wire core__abc_22172_new_n1788_; 
wire core__abc_22172_new_n1789_; 
wire core__abc_22172_new_n1790_; 
wire core__abc_22172_new_n1791_; 
wire core__abc_22172_new_n1792_; 
wire core__abc_22172_new_n1793_; 
wire core__abc_22172_new_n1794_; 
wire core__abc_22172_new_n1795_; 
wire core__abc_22172_new_n1796_; 
wire core__abc_22172_new_n1797_; 
wire core__abc_22172_new_n1799_; 
wire core__abc_22172_new_n1800_; 
wire core__abc_22172_new_n1801_; 
wire core__abc_22172_new_n1802_; 
wire core__abc_22172_new_n1803_; 
wire core__abc_22172_new_n1804_; 
wire core__abc_22172_new_n1805_; 
wire core__abc_22172_new_n1806_; 
wire core__abc_22172_new_n1807_; 
wire core__abc_22172_new_n1808_; 
wire core__abc_22172_new_n1809_; 
wire core__abc_22172_new_n1810_; 
wire core__abc_22172_new_n1811_; 
wire core__abc_22172_new_n1812_; 
wire core__abc_22172_new_n1813_; 
wire core__abc_22172_new_n1814_; 
wire core__abc_22172_new_n1816_; 
wire core__abc_22172_new_n1817_; 
wire core__abc_22172_new_n1818_; 
wire core__abc_22172_new_n1819_; 
wire core__abc_22172_new_n1820_; 
wire core__abc_22172_new_n1821_; 
wire core__abc_22172_new_n1822_; 
wire core__abc_22172_new_n1823_; 
wire core__abc_22172_new_n1824_; 
wire core__abc_22172_new_n1825_; 
wire core__abc_22172_new_n1826_; 
wire core__abc_22172_new_n1827_; 
wire core__abc_22172_new_n1828_; 
wire core__abc_22172_new_n1829_; 
wire core__abc_22172_new_n1830_; 
wire core__abc_22172_new_n1831_; 
wire core__abc_22172_new_n1833_; 
wire core__abc_22172_new_n1834_; 
wire core__abc_22172_new_n1835_; 
wire core__abc_22172_new_n1836_; 
wire core__abc_22172_new_n1837_; 
wire core__abc_22172_new_n1838_; 
wire core__abc_22172_new_n1839_; 
wire core__abc_22172_new_n1840_; 
wire core__abc_22172_new_n1841_; 
wire core__abc_22172_new_n1842_; 
wire core__abc_22172_new_n1843_; 
wire core__abc_22172_new_n1844_; 
wire core__abc_22172_new_n1845_; 
wire core__abc_22172_new_n1846_; 
wire core__abc_22172_new_n1847_; 
wire core__abc_22172_new_n1848_; 
wire core__abc_22172_new_n1850_; 
wire core__abc_22172_new_n1851_; 
wire core__abc_22172_new_n1852_; 
wire core__abc_22172_new_n1853_; 
wire core__abc_22172_new_n1854_; 
wire core__abc_22172_new_n1855_; 
wire core__abc_22172_new_n1856_; 
wire core__abc_22172_new_n1857_; 
wire core__abc_22172_new_n1858_; 
wire core__abc_22172_new_n1859_; 
wire core__abc_22172_new_n1860_; 
wire core__abc_22172_new_n1861_; 
wire core__abc_22172_new_n1862_; 
wire core__abc_22172_new_n1863_; 
wire core__abc_22172_new_n1864_; 
wire core__abc_22172_new_n1865_; 
wire core__abc_22172_new_n1867_; 
wire core__abc_22172_new_n1868_; 
wire core__abc_22172_new_n1869_; 
wire core__abc_22172_new_n1870_; 
wire core__abc_22172_new_n1871_; 
wire core__abc_22172_new_n1872_; 
wire core__abc_22172_new_n1873_; 
wire core__abc_22172_new_n1874_; 
wire core__abc_22172_new_n1875_; 
wire core__abc_22172_new_n1876_; 
wire core__abc_22172_new_n1877_; 
wire core__abc_22172_new_n1878_; 
wire core__abc_22172_new_n1879_; 
wire core__abc_22172_new_n1880_; 
wire core__abc_22172_new_n1881_; 
wire core__abc_22172_new_n1882_; 
wire core__abc_22172_new_n1884_; 
wire core__abc_22172_new_n1885_; 
wire core__abc_22172_new_n1886_; 
wire core__abc_22172_new_n1887_; 
wire core__abc_22172_new_n1888_; 
wire core__abc_22172_new_n1889_; 
wire core__abc_22172_new_n1890_; 
wire core__abc_22172_new_n1891_; 
wire core__abc_22172_new_n1892_; 
wire core__abc_22172_new_n1893_; 
wire core__abc_22172_new_n1894_; 
wire core__abc_22172_new_n1895_; 
wire core__abc_22172_new_n1896_; 
wire core__abc_22172_new_n1897_; 
wire core__abc_22172_new_n1898_; 
wire core__abc_22172_new_n1899_; 
wire core__abc_22172_new_n1901_; 
wire core__abc_22172_new_n1902_; 
wire core__abc_22172_new_n1903_; 
wire core__abc_22172_new_n1904_; 
wire core__abc_22172_new_n1905_; 
wire core__abc_22172_new_n1906_; 
wire core__abc_22172_new_n1907_; 
wire core__abc_22172_new_n1908_; 
wire core__abc_22172_new_n1909_; 
wire core__abc_22172_new_n1910_; 
wire core__abc_22172_new_n1911_; 
wire core__abc_22172_new_n1912_; 
wire core__abc_22172_new_n1913_; 
wire core__abc_22172_new_n1914_; 
wire core__abc_22172_new_n1915_; 
wire core__abc_22172_new_n1916_; 
wire core__abc_22172_new_n1918_; 
wire core__abc_22172_new_n1919_; 
wire core__abc_22172_new_n1920_; 
wire core__abc_22172_new_n1921_; 
wire core__abc_22172_new_n1922_; 
wire core__abc_22172_new_n1923_; 
wire core__abc_22172_new_n1924_; 
wire core__abc_22172_new_n1925_; 
wire core__abc_22172_new_n1926_; 
wire core__abc_22172_new_n1927_; 
wire core__abc_22172_new_n1928_; 
wire core__abc_22172_new_n1929_; 
wire core__abc_22172_new_n1930_; 
wire core__abc_22172_new_n1931_; 
wire core__abc_22172_new_n1932_; 
wire core__abc_22172_new_n1933_; 
wire core__abc_22172_new_n1935_; 
wire core__abc_22172_new_n1936_; 
wire core__abc_22172_new_n1937_; 
wire core__abc_22172_new_n1938_; 
wire core__abc_22172_new_n1939_; 
wire core__abc_22172_new_n1940_; 
wire core__abc_22172_new_n1941_; 
wire core__abc_22172_new_n1942_; 
wire core__abc_22172_new_n1943_; 
wire core__abc_22172_new_n1944_; 
wire core__abc_22172_new_n1945_; 
wire core__abc_22172_new_n1946_; 
wire core__abc_22172_new_n1947_; 
wire core__abc_22172_new_n1948_; 
wire core__abc_22172_new_n1949_; 
wire core__abc_22172_new_n1950_; 
wire core__abc_22172_new_n1952_; 
wire core__abc_22172_new_n1953_; 
wire core__abc_22172_new_n1954_; 
wire core__abc_22172_new_n1955_; 
wire core__abc_22172_new_n1956_; 
wire core__abc_22172_new_n1957_; 
wire core__abc_22172_new_n1958_; 
wire core__abc_22172_new_n1959_; 
wire core__abc_22172_new_n1960_; 
wire core__abc_22172_new_n1961_; 
wire core__abc_22172_new_n1962_; 
wire core__abc_22172_new_n1963_; 
wire core__abc_22172_new_n1964_; 
wire core__abc_22172_new_n1965_; 
wire core__abc_22172_new_n1966_; 
wire core__abc_22172_new_n1967_; 
wire core__abc_22172_new_n1969_; 
wire core__abc_22172_new_n1970_; 
wire core__abc_22172_new_n1971_; 
wire core__abc_22172_new_n1972_; 
wire core__abc_22172_new_n1973_; 
wire core__abc_22172_new_n1974_; 
wire core__abc_22172_new_n1975_; 
wire core__abc_22172_new_n1976_; 
wire core__abc_22172_new_n1977_; 
wire core__abc_22172_new_n1978_; 
wire core__abc_22172_new_n1979_; 
wire core__abc_22172_new_n1980_; 
wire core__abc_22172_new_n1981_; 
wire core__abc_22172_new_n1982_; 
wire core__abc_22172_new_n1983_; 
wire core__abc_22172_new_n1984_; 
wire core__abc_22172_new_n1986_; 
wire core__abc_22172_new_n1987_; 
wire core__abc_22172_new_n1988_; 
wire core__abc_22172_new_n1989_; 
wire core__abc_22172_new_n1990_; 
wire core__abc_22172_new_n1991_; 
wire core__abc_22172_new_n1992_; 
wire core__abc_22172_new_n1993_; 
wire core__abc_22172_new_n1994_; 
wire core__abc_22172_new_n1995_; 
wire core__abc_22172_new_n1996_; 
wire core__abc_22172_new_n1997_; 
wire core__abc_22172_new_n1998_; 
wire core__abc_22172_new_n1999_; 
wire core__abc_22172_new_n2000_; 
wire core__abc_22172_new_n2001_; 
wire core__abc_22172_new_n2003_; 
wire core__abc_22172_new_n2004_; 
wire core__abc_22172_new_n2005_; 
wire core__abc_22172_new_n2006_; 
wire core__abc_22172_new_n2007_; 
wire core__abc_22172_new_n2008_; 
wire core__abc_22172_new_n2009_; 
wire core__abc_22172_new_n2010_; 
wire core__abc_22172_new_n2011_; 
wire core__abc_22172_new_n2012_; 
wire core__abc_22172_new_n2013_; 
wire core__abc_22172_new_n2014_; 
wire core__abc_22172_new_n2015_; 
wire core__abc_22172_new_n2016_; 
wire core__abc_22172_new_n2017_; 
wire core__abc_22172_new_n2018_; 
wire core__abc_22172_new_n2020_; 
wire core__abc_22172_new_n2021_; 
wire core__abc_22172_new_n2022_; 
wire core__abc_22172_new_n2023_; 
wire core__abc_22172_new_n2024_; 
wire core__abc_22172_new_n2025_; 
wire core__abc_22172_new_n2026_; 
wire core__abc_22172_new_n2027_; 
wire core__abc_22172_new_n2028_; 
wire core__abc_22172_new_n2029_; 
wire core__abc_22172_new_n2030_; 
wire core__abc_22172_new_n2031_; 
wire core__abc_22172_new_n2032_; 
wire core__abc_22172_new_n2033_; 
wire core__abc_22172_new_n2034_; 
wire core__abc_22172_new_n2035_; 
wire core__abc_22172_new_n2037_; 
wire core__abc_22172_new_n2038_; 
wire core__abc_22172_new_n2039_; 
wire core__abc_22172_new_n2040_; 
wire core__abc_22172_new_n2041_; 
wire core__abc_22172_new_n2042_; 
wire core__abc_22172_new_n2043_; 
wire core__abc_22172_new_n2044_; 
wire core__abc_22172_new_n2045_; 
wire core__abc_22172_new_n2046_; 
wire core__abc_22172_new_n2047_; 
wire core__abc_22172_new_n2048_; 
wire core__abc_22172_new_n2049_; 
wire core__abc_22172_new_n2050_; 
wire core__abc_22172_new_n2051_; 
wire core__abc_22172_new_n2052_; 
wire core__abc_22172_new_n2054_; 
wire core__abc_22172_new_n2055_; 
wire core__abc_22172_new_n2056_; 
wire core__abc_22172_new_n2057_; 
wire core__abc_22172_new_n2058_; 
wire core__abc_22172_new_n2059_; 
wire core__abc_22172_new_n2060_; 
wire core__abc_22172_new_n2061_; 
wire core__abc_22172_new_n2062_; 
wire core__abc_22172_new_n2063_; 
wire core__abc_22172_new_n2064_; 
wire core__abc_22172_new_n2065_; 
wire core__abc_22172_new_n2066_; 
wire core__abc_22172_new_n2067_; 
wire core__abc_22172_new_n2068_; 
wire core__abc_22172_new_n2069_; 
wire core__abc_22172_new_n2071_; 
wire core__abc_22172_new_n2072_; 
wire core__abc_22172_new_n2073_; 
wire core__abc_22172_new_n2074_; 
wire core__abc_22172_new_n2075_; 
wire core__abc_22172_new_n2076_; 
wire core__abc_22172_new_n2077_; 
wire core__abc_22172_new_n2078_; 
wire core__abc_22172_new_n2079_; 
wire core__abc_22172_new_n2080_; 
wire core__abc_22172_new_n2081_; 
wire core__abc_22172_new_n2082_; 
wire core__abc_22172_new_n2083_; 
wire core__abc_22172_new_n2084_; 
wire core__abc_22172_new_n2085_; 
wire core__abc_22172_new_n2086_; 
wire core__abc_22172_new_n2088_; 
wire core__abc_22172_new_n2089_; 
wire core__abc_22172_new_n2090_; 
wire core__abc_22172_new_n2091_; 
wire core__abc_22172_new_n2092_; 
wire core__abc_22172_new_n2093_; 
wire core__abc_22172_new_n2094_; 
wire core__abc_22172_new_n2095_; 
wire core__abc_22172_new_n2096_; 
wire core__abc_22172_new_n2097_; 
wire core__abc_22172_new_n2098_; 
wire core__abc_22172_new_n2099_; 
wire core__abc_22172_new_n2100_; 
wire core__abc_22172_new_n2101_; 
wire core__abc_22172_new_n2102_; 
wire core__abc_22172_new_n2103_; 
wire core__abc_22172_new_n2105_; 
wire core__abc_22172_new_n2106_; 
wire core__abc_22172_new_n2107_; 
wire core__abc_22172_new_n2108_; 
wire core__abc_22172_new_n2109_; 
wire core__abc_22172_new_n2110_; 
wire core__abc_22172_new_n2111_; 
wire core__abc_22172_new_n2112_; 
wire core__abc_22172_new_n2113_; 
wire core__abc_22172_new_n2114_; 
wire core__abc_22172_new_n2115_; 
wire core__abc_22172_new_n2116_; 
wire core__abc_22172_new_n2117_; 
wire core__abc_22172_new_n2118_; 
wire core__abc_22172_new_n2119_; 
wire core__abc_22172_new_n2120_; 
wire core__abc_22172_new_n2122_; 
wire core__abc_22172_new_n2123_; 
wire core__abc_22172_new_n2124_; 
wire core__abc_22172_new_n2125_; 
wire core__abc_22172_new_n2126_; 
wire core__abc_22172_new_n2127_; 
wire core__abc_22172_new_n2128_; 
wire core__abc_22172_new_n2129_; 
wire core__abc_22172_new_n2130_; 
wire core__abc_22172_new_n2131_; 
wire core__abc_22172_new_n2132_; 
wire core__abc_22172_new_n2133_; 
wire core__abc_22172_new_n2134_; 
wire core__abc_22172_new_n2135_; 
wire core__abc_22172_new_n2136_; 
wire core__abc_22172_new_n2137_; 
wire core__abc_22172_new_n2139_; 
wire core__abc_22172_new_n2140_; 
wire core__abc_22172_new_n2141_; 
wire core__abc_22172_new_n2142_; 
wire core__abc_22172_new_n2143_; 
wire core__abc_22172_new_n2144_; 
wire core__abc_22172_new_n2145_; 
wire core__abc_22172_new_n2146_; 
wire core__abc_22172_new_n2147_; 
wire core__abc_22172_new_n2148_; 
wire core__abc_22172_new_n2149_; 
wire core__abc_22172_new_n2150_; 
wire core__abc_22172_new_n2151_; 
wire core__abc_22172_new_n2152_; 
wire core__abc_22172_new_n2153_; 
wire core__abc_22172_new_n2154_; 
wire core__abc_22172_new_n2156_; 
wire core__abc_22172_new_n2157_; 
wire core__abc_22172_new_n2158_; 
wire core__abc_22172_new_n2159_; 
wire core__abc_22172_new_n2160_; 
wire core__abc_22172_new_n2161_; 
wire core__abc_22172_new_n2162_; 
wire core__abc_22172_new_n2163_; 
wire core__abc_22172_new_n2164_; 
wire core__abc_22172_new_n2165_; 
wire core__abc_22172_new_n2166_; 
wire core__abc_22172_new_n2167_; 
wire core__abc_22172_new_n2168_; 
wire core__abc_22172_new_n2169_; 
wire core__abc_22172_new_n2170_; 
wire core__abc_22172_new_n2171_; 
wire core__abc_22172_new_n2173_; 
wire core__abc_22172_new_n2174_; 
wire core__abc_22172_new_n2175_; 
wire core__abc_22172_new_n2176_; 
wire core__abc_22172_new_n2177_; 
wire core__abc_22172_new_n2178_; 
wire core__abc_22172_new_n2179_; 
wire core__abc_22172_new_n2180_; 
wire core__abc_22172_new_n2181_; 
wire core__abc_22172_new_n2182_; 
wire core__abc_22172_new_n2183_; 
wire core__abc_22172_new_n2184_; 
wire core__abc_22172_new_n2185_; 
wire core__abc_22172_new_n2186_; 
wire core__abc_22172_new_n2187_; 
wire core__abc_22172_new_n2188_; 
wire core__abc_22172_new_n2190_; 
wire core__abc_22172_new_n2191_; 
wire core__abc_22172_new_n2192_; 
wire core__abc_22172_new_n2193_; 
wire core__abc_22172_new_n2194_; 
wire core__abc_22172_new_n2195_; 
wire core__abc_22172_new_n2196_; 
wire core__abc_22172_new_n2197_; 
wire core__abc_22172_new_n2198_; 
wire core__abc_22172_new_n2199_; 
wire core__abc_22172_new_n2200_; 
wire core__abc_22172_new_n2201_; 
wire core__abc_22172_new_n2202_; 
wire core__abc_22172_new_n2203_; 
wire core__abc_22172_new_n2204_; 
wire core__abc_22172_new_n2205_; 
wire core__abc_22172_new_n2207_; 
wire core__abc_22172_new_n2208_; 
wire core__abc_22172_new_n2209_; 
wire core__abc_22172_new_n2210_; 
wire core__abc_22172_new_n2211_; 
wire core__abc_22172_new_n2212_; 
wire core__abc_22172_new_n2213_; 
wire core__abc_22172_new_n2214_; 
wire core__abc_22172_new_n2215_; 
wire core__abc_22172_new_n2216_; 
wire core__abc_22172_new_n2217_; 
wire core__abc_22172_new_n2218_; 
wire core__abc_22172_new_n2219_; 
wire core__abc_22172_new_n2220_; 
wire core__abc_22172_new_n2221_; 
wire core__abc_22172_new_n2222_; 
wire core__abc_22172_new_n2224_; 
wire core__abc_22172_new_n2225_; 
wire core__abc_22172_new_n2226_; 
wire core__abc_22172_new_n2227_; 
wire core__abc_22172_new_n2228_; 
wire core__abc_22172_new_n2229_; 
wire core__abc_22172_new_n2230_; 
wire core__abc_22172_new_n2231_; 
wire core__abc_22172_new_n2232_; 
wire core__abc_22172_new_n2233_; 
wire core__abc_22172_new_n2234_; 
wire core__abc_22172_new_n2235_; 
wire core__abc_22172_new_n2236_; 
wire core__abc_22172_new_n2237_; 
wire core__abc_22172_new_n2238_; 
wire core__abc_22172_new_n2239_; 
wire core__abc_22172_new_n2241_; 
wire core__abc_22172_new_n2242_; 
wire core__abc_22172_new_n2243_; 
wire core__abc_22172_new_n2244_; 
wire core__abc_22172_new_n2245_; 
wire core__abc_22172_new_n2246_; 
wire core__abc_22172_new_n2247_; 
wire core__abc_22172_new_n2248_; 
wire core__abc_22172_new_n2249_; 
wire core__abc_22172_new_n2250_; 
wire core__abc_22172_new_n2251_; 
wire core__abc_22172_new_n2252_; 
wire core__abc_22172_new_n2253_; 
wire core__abc_22172_new_n2254_; 
wire core__abc_22172_new_n2255_; 
wire core__abc_22172_new_n2256_; 
wire core__abc_22172_new_n2258_; 
wire core__abc_22172_new_n2259_; 
wire core__abc_22172_new_n2260_; 
wire core__abc_22172_new_n2261_; 
wire core__abc_22172_new_n2262_; 
wire core__abc_22172_new_n2263_; 
wire core__abc_22172_new_n2264_; 
wire core__abc_22172_new_n2265_; 
wire core__abc_22172_new_n2266_; 
wire core__abc_22172_new_n2267_; 
wire core__abc_22172_new_n2268_; 
wire core__abc_22172_new_n2269_; 
wire core__abc_22172_new_n2270_; 
wire core__abc_22172_new_n2271_; 
wire core__abc_22172_new_n2272_; 
wire core__abc_22172_new_n2273_; 
wire core__abc_22172_new_n2275_; 
wire core__abc_22172_new_n2276_; 
wire core__abc_22172_new_n2277_; 
wire core__abc_22172_new_n2278_; 
wire core__abc_22172_new_n2279_; 
wire core__abc_22172_new_n2280_; 
wire core__abc_22172_new_n2281_; 
wire core__abc_22172_new_n2282_; 
wire core__abc_22172_new_n2283_; 
wire core__abc_22172_new_n2284_; 
wire core__abc_22172_new_n2285_; 
wire core__abc_22172_new_n2286_; 
wire core__abc_22172_new_n2287_; 
wire core__abc_22172_new_n2288_; 
wire core__abc_22172_new_n2289_; 
wire core__abc_22172_new_n2290_; 
wire core__abc_22172_new_n2292_; 
wire core__abc_22172_new_n2293_; 
wire core__abc_22172_new_n2294_; 
wire core__abc_22172_new_n2295_; 
wire core__abc_22172_new_n2296_; 
wire core__abc_22172_new_n2297_; 
wire core__abc_22172_new_n2298_; 
wire core__abc_22172_new_n2299_; 
wire core__abc_22172_new_n2300_; 
wire core__abc_22172_new_n2301_; 
wire core__abc_22172_new_n2302_; 
wire core__abc_22172_new_n2303_; 
wire core__abc_22172_new_n2304_; 
wire core__abc_22172_new_n2305_; 
wire core__abc_22172_new_n2306_; 
wire core__abc_22172_new_n2307_; 
wire core__abc_22172_new_n2309_; 
wire core__abc_22172_new_n2310_; 
wire core__abc_22172_new_n2311_; 
wire core__abc_22172_new_n2312_; 
wire core__abc_22172_new_n2313_; 
wire core__abc_22172_new_n2314_; 
wire core__abc_22172_new_n2315_; 
wire core__abc_22172_new_n2316_; 
wire core__abc_22172_new_n2317_; 
wire core__abc_22172_new_n2318_; 
wire core__abc_22172_new_n2319_; 
wire core__abc_22172_new_n2320_; 
wire core__abc_22172_new_n2321_; 
wire core__abc_22172_new_n2322_; 
wire core__abc_22172_new_n2323_; 
wire core__abc_22172_new_n2324_; 
wire core__abc_22172_new_n2326_; 
wire core__abc_22172_new_n2327_; 
wire core__abc_22172_new_n2328_; 
wire core__abc_22172_new_n2329_; 
wire core__abc_22172_new_n2330_; 
wire core__abc_22172_new_n2331_; 
wire core__abc_22172_new_n2332_; 
wire core__abc_22172_new_n2333_; 
wire core__abc_22172_new_n2334_; 
wire core__abc_22172_new_n2335_; 
wire core__abc_22172_new_n2336_; 
wire core__abc_22172_new_n2337_; 
wire core__abc_22172_new_n2338_; 
wire core__abc_22172_new_n2339_; 
wire core__abc_22172_new_n2340_; 
wire core__abc_22172_new_n2341_; 
wire core__abc_22172_new_n2343_; 
wire core__abc_22172_new_n2344_; 
wire core__abc_22172_new_n2345_; 
wire core__abc_22172_new_n2346_; 
wire core__abc_22172_new_n2347_; 
wire core__abc_22172_new_n2348_; 
wire core__abc_22172_new_n2349_; 
wire core__abc_22172_new_n2350_; 
wire core__abc_22172_new_n2351_; 
wire core__abc_22172_new_n2352_; 
wire core__abc_22172_new_n2353_; 
wire core__abc_22172_new_n2354_; 
wire core__abc_22172_new_n2355_; 
wire core__abc_22172_new_n2356_; 
wire core__abc_22172_new_n2357_; 
wire core__abc_22172_new_n2358_; 
wire core__abc_22172_new_n2359_; 
wire core__abc_22172_new_n2361_; 
wire core__abc_22172_new_n2362_; 
wire core__abc_22172_new_n2363_; 
wire core__abc_22172_new_n2364_; 
wire core__abc_22172_new_n2365_; 
wire core__abc_22172_new_n2366_; 
wire core__abc_22172_new_n2367_; 
wire core__abc_22172_new_n2368_; 
wire core__abc_22172_new_n2370_; 
wire core__abc_22172_new_n2371_; 
wire core__abc_22172_new_n2372_; 
wire core__abc_22172_new_n2374_; 
wire core__abc_22172_new_n2375_; 
wire core__abc_22172_new_n2376_; 
wire core__abc_22172_new_n2378_; 
wire core__abc_22172_new_n2379_; 
wire core__abc_22172_new_n2380_; 
wire core__abc_22172_new_n2382_; 
wire core__abc_22172_new_n2383_; 
wire core__abc_22172_new_n2384_; 
wire core__abc_22172_new_n2386_; 
wire core__abc_22172_new_n2387_; 
wire core__abc_22172_new_n2388_; 
wire core__abc_22172_new_n2390_; 
wire core__abc_22172_new_n2391_; 
wire core__abc_22172_new_n2392_; 
wire core__abc_22172_new_n2394_; 
wire core__abc_22172_new_n2395_; 
wire core__abc_22172_new_n2396_; 
wire core__abc_22172_new_n2398_; 
wire core__abc_22172_new_n2399_; 
wire core__abc_22172_new_n2400_; 
wire core__abc_22172_new_n2402_; 
wire core__abc_22172_new_n2403_; 
wire core__abc_22172_new_n2404_; 
wire core__abc_22172_new_n2406_; 
wire core__abc_22172_new_n2407_; 
wire core__abc_22172_new_n2408_; 
wire core__abc_22172_new_n2410_; 
wire core__abc_22172_new_n2411_; 
wire core__abc_22172_new_n2412_; 
wire core__abc_22172_new_n2414_; 
wire core__abc_22172_new_n2415_; 
wire core__abc_22172_new_n2416_; 
wire core__abc_22172_new_n2418_; 
wire core__abc_22172_new_n2419_; 
wire core__abc_22172_new_n2420_; 
wire core__abc_22172_new_n2422_; 
wire core__abc_22172_new_n2423_; 
wire core__abc_22172_new_n2424_; 
wire core__abc_22172_new_n2426_; 
wire core__abc_22172_new_n2427_; 
wire core__abc_22172_new_n2428_; 
wire core__abc_22172_new_n2430_; 
wire core__abc_22172_new_n2431_; 
wire core__abc_22172_new_n2432_; 
wire core__abc_22172_new_n2434_; 
wire core__abc_22172_new_n2435_; 
wire core__abc_22172_new_n2436_; 
wire core__abc_22172_new_n2438_; 
wire core__abc_22172_new_n2439_; 
wire core__abc_22172_new_n2440_; 
wire core__abc_22172_new_n2442_; 
wire core__abc_22172_new_n2443_; 
wire core__abc_22172_new_n2444_; 
wire core__abc_22172_new_n2446_; 
wire core__abc_22172_new_n2447_; 
wire core__abc_22172_new_n2448_; 
wire core__abc_22172_new_n2450_; 
wire core__abc_22172_new_n2451_; 
wire core__abc_22172_new_n2452_; 
wire core__abc_22172_new_n2454_; 
wire core__abc_22172_new_n2455_; 
wire core__abc_22172_new_n2456_; 
wire core__abc_22172_new_n2458_; 
wire core__abc_22172_new_n2459_; 
wire core__abc_22172_new_n2460_; 
wire core__abc_22172_new_n2462_; 
wire core__abc_22172_new_n2463_; 
wire core__abc_22172_new_n2464_; 
wire core__abc_22172_new_n2466_; 
wire core__abc_22172_new_n2467_; 
wire core__abc_22172_new_n2468_; 
wire core__abc_22172_new_n2470_; 
wire core__abc_22172_new_n2471_; 
wire core__abc_22172_new_n2472_; 
wire core__abc_22172_new_n2474_; 
wire core__abc_22172_new_n2475_; 
wire core__abc_22172_new_n2476_; 
wire core__abc_22172_new_n2478_; 
wire core__abc_22172_new_n2479_; 
wire core__abc_22172_new_n2480_; 
wire core__abc_22172_new_n2482_; 
wire core__abc_22172_new_n2483_; 
wire core__abc_22172_new_n2484_; 
wire core__abc_22172_new_n2486_; 
wire core__abc_22172_new_n2487_; 
wire core__abc_22172_new_n2488_; 
wire core__abc_22172_new_n2490_; 
wire core__abc_22172_new_n2491_; 
wire core__abc_22172_new_n2492_; 
wire core__abc_22172_new_n2494_; 
wire core__abc_22172_new_n2495_; 
wire core__abc_22172_new_n2496_; 
wire core__abc_22172_new_n2498_; 
wire core__abc_22172_new_n2499_; 
wire core__abc_22172_new_n2500_; 
wire core__abc_22172_new_n2502_; 
wire core__abc_22172_new_n2503_; 
wire core__abc_22172_new_n2504_; 
wire core__abc_22172_new_n2506_; 
wire core__abc_22172_new_n2507_; 
wire core__abc_22172_new_n2508_; 
wire core__abc_22172_new_n2510_; 
wire core__abc_22172_new_n2511_; 
wire core__abc_22172_new_n2512_; 
wire core__abc_22172_new_n2514_; 
wire core__abc_22172_new_n2515_; 
wire core__abc_22172_new_n2516_; 
wire core__abc_22172_new_n2518_; 
wire core__abc_22172_new_n2519_; 
wire core__abc_22172_new_n2520_; 
wire core__abc_22172_new_n2522_; 
wire core__abc_22172_new_n2523_; 
wire core__abc_22172_new_n2524_; 
wire core__abc_22172_new_n2526_; 
wire core__abc_22172_new_n2527_; 
wire core__abc_22172_new_n2528_; 
wire core__abc_22172_new_n2530_; 
wire core__abc_22172_new_n2531_; 
wire core__abc_22172_new_n2532_; 
wire core__abc_22172_new_n2534_; 
wire core__abc_22172_new_n2535_; 
wire core__abc_22172_new_n2536_; 
wire core__abc_22172_new_n2538_; 
wire core__abc_22172_new_n2539_; 
wire core__abc_22172_new_n2540_; 
wire core__abc_22172_new_n2542_; 
wire core__abc_22172_new_n2543_; 
wire core__abc_22172_new_n2544_; 
wire core__abc_22172_new_n2546_; 
wire core__abc_22172_new_n2547_; 
wire core__abc_22172_new_n2548_; 
wire core__abc_22172_new_n2550_; 
wire core__abc_22172_new_n2551_; 
wire core__abc_22172_new_n2552_; 
wire core__abc_22172_new_n2554_; 
wire core__abc_22172_new_n2555_; 
wire core__abc_22172_new_n2556_; 
wire core__abc_22172_new_n2558_; 
wire core__abc_22172_new_n2559_; 
wire core__abc_22172_new_n2560_; 
wire core__abc_22172_new_n2562_; 
wire core__abc_22172_new_n2563_; 
wire core__abc_22172_new_n2564_; 
wire core__abc_22172_new_n2566_; 
wire core__abc_22172_new_n2567_; 
wire core__abc_22172_new_n2568_; 
wire core__abc_22172_new_n2570_; 
wire core__abc_22172_new_n2571_; 
wire core__abc_22172_new_n2572_; 
wire core__abc_22172_new_n2574_; 
wire core__abc_22172_new_n2575_; 
wire core__abc_22172_new_n2576_; 
wire core__abc_22172_new_n2578_; 
wire core__abc_22172_new_n2579_; 
wire core__abc_22172_new_n2580_; 
wire core__abc_22172_new_n2582_; 
wire core__abc_22172_new_n2583_; 
wire core__abc_22172_new_n2584_; 
wire core__abc_22172_new_n2586_; 
wire core__abc_22172_new_n2587_; 
wire core__abc_22172_new_n2588_; 
wire core__abc_22172_new_n2590_; 
wire core__abc_22172_new_n2591_; 
wire core__abc_22172_new_n2592_; 
wire core__abc_22172_new_n2594_; 
wire core__abc_22172_new_n2595_; 
wire core__abc_22172_new_n2596_; 
wire core__abc_22172_new_n2598_; 
wire core__abc_22172_new_n2599_; 
wire core__abc_22172_new_n2600_; 
wire core__abc_22172_new_n2602_; 
wire core__abc_22172_new_n2603_; 
wire core__abc_22172_new_n2604_; 
wire core__abc_22172_new_n2606_; 
wire core__abc_22172_new_n2607_; 
wire core__abc_22172_new_n2608_; 
wire core__abc_22172_new_n2610_; 
wire core__abc_22172_new_n2611_; 
wire core__abc_22172_new_n2612_; 
wire core__abc_22172_new_n2614_; 
wire core__abc_22172_new_n2615_; 
wire core__abc_22172_new_n2616_; 
wire core__abc_22172_new_n2618_; 
wire core__abc_22172_new_n2619_; 
wire core__abc_22172_new_n2620_; 
wire core__abc_22172_new_n2622_; 
wire core__abc_22172_new_n2623_; 
wire core__abc_22172_new_n2624_; 
wire core__abc_22172_new_n2625_; 
wire core__abc_22172_new_n2626_; 
wire core__abc_22172_new_n2628_; 
wire core__abc_22172_new_n2629_; 
wire core__abc_22172_new_n2630_; 
wire core__abc_22172_new_n2631_; 
wire core__abc_22172_new_n2632_; 
wire core__abc_22172_new_n2633_; 
wire core__abc_22172_new_n2634_; 
wire core__abc_22172_new_n2635_; 
wire core__abc_22172_new_n2636_; 
wire core__abc_22172_new_n2637_; 
wire core__abc_22172_new_n2639_; 
wire core__abc_22172_new_n2640_; 
wire core__abc_22172_new_n2641_; 
wire core__abc_22172_new_n2642_; 
wire core__abc_22172_new_n2643_; 
wire core__abc_22172_new_n2644_; 
wire core__abc_22172_new_n2646_; 
wire core__abc_22172_new_n2647_; 
wire core__abc_22172_new_n2648_; 
wire core__abc_22172_new_n2649_; 
wire core__abc_22172_new_n2650_; 
wire core__abc_22172_new_n2651_; 
wire core__abc_22172_new_n2652_; 
wire core__abc_22172_new_n2654_; 
wire core__abc_22172_new_n2655_; 
wire core__abc_22172_new_n2656_; 
wire core__abc_22172_new_n2657_; 
wire core__abc_22172_new_n2659_; 
wire core__abc_22172_new_n2660_; 
wire core__abc_22172_new_n2661_; 
wire core__abc_22172_new_n2662_; 
wire core__abc_22172_new_n2663_; 
wire core__abc_22172_new_n2664_; 
wire core__abc_22172_new_n2666_; 
wire core__abc_22172_new_n2667_; 
wire core__abc_22172_new_n2668_; 
wire core__abc_22172_new_n2670_; 
wire core__abc_22172_new_n2671_; 
wire core__abc_22172_new_n2672_; 
wire core__abc_22172_new_n2674_; 
wire core__abc_22172_new_n2675_; 
wire core__abc_22172_new_n2676_; 
wire core__abc_22172_new_n2678_; 
wire core__abc_22172_new_n2679_; 
wire core__abc_22172_new_n2680_; 
wire core__abc_22172_new_n2682_; 
wire core__abc_22172_new_n2683_; 
wire core__abc_22172_new_n2684_; 
wire core__abc_22172_new_n2686_; 
wire core__abc_22172_new_n2687_; 
wire core__abc_22172_new_n2688_; 
wire core__abc_22172_new_n2690_; 
wire core__abc_22172_new_n2691_; 
wire core__abc_22172_new_n2692_; 
wire core__abc_22172_new_n2694_; 
wire core__abc_22172_new_n2695_; 
wire core__abc_22172_new_n2696_; 
wire core__abc_22172_new_n2698_; 
wire core__abc_22172_new_n2699_; 
wire core__abc_22172_new_n2700_; 
wire core__abc_22172_new_n2702_; 
wire core__abc_22172_new_n2703_; 
wire core__abc_22172_new_n2704_; 
wire core__abc_22172_new_n2706_; 
wire core__abc_22172_new_n2707_; 
wire core__abc_22172_new_n2708_; 
wire core__abc_22172_new_n2710_; 
wire core__abc_22172_new_n2711_; 
wire core__abc_22172_new_n2712_; 
wire core__abc_22172_new_n2714_; 
wire core__abc_22172_new_n2715_; 
wire core__abc_22172_new_n2716_; 
wire core__abc_22172_new_n2718_; 
wire core__abc_22172_new_n2719_; 
wire core__abc_22172_new_n2720_; 
wire core__abc_22172_new_n2722_; 
wire core__abc_22172_new_n2723_; 
wire core__abc_22172_new_n2724_; 
wire core__abc_22172_new_n2726_; 
wire core__abc_22172_new_n2727_; 
wire core__abc_22172_new_n2728_; 
wire core__abc_22172_new_n2730_; 
wire core__abc_22172_new_n2731_; 
wire core__abc_22172_new_n2732_; 
wire core__abc_22172_new_n2734_; 
wire core__abc_22172_new_n2735_; 
wire core__abc_22172_new_n2736_; 
wire core__abc_22172_new_n2738_; 
wire core__abc_22172_new_n2739_; 
wire core__abc_22172_new_n2740_; 
wire core__abc_22172_new_n2742_; 
wire core__abc_22172_new_n2743_; 
wire core__abc_22172_new_n2744_; 
wire core__abc_22172_new_n2746_; 
wire core__abc_22172_new_n2747_; 
wire core__abc_22172_new_n2748_; 
wire core__abc_22172_new_n2750_; 
wire core__abc_22172_new_n2751_; 
wire core__abc_22172_new_n2752_; 
wire core__abc_22172_new_n2754_; 
wire core__abc_22172_new_n2755_; 
wire core__abc_22172_new_n2756_; 
wire core__abc_22172_new_n2758_; 
wire core__abc_22172_new_n2759_; 
wire core__abc_22172_new_n2760_; 
wire core__abc_22172_new_n2762_; 
wire core__abc_22172_new_n2763_; 
wire core__abc_22172_new_n2764_; 
wire core__abc_22172_new_n2766_; 
wire core__abc_22172_new_n2767_; 
wire core__abc_22172_new_n2768_; 
wire core__abc_22172_new_n2770_; 
wire core__abc_22172_new_n2771_; 
wire core__abc_22172_new_n2772_; 
wire core__abc_22172_new_n2774_; 
wire core__abc_22172_new_n2775_; 
wire core__abc_22172_new_n2776_; 
wire core__abc_22172_new_n2778_; 
wire core__abc_22172_new_n2779_; 
wire core__abc_22172_new_n2780_; 
wire core__abc_22172_new_n2782_; 
wire core__abc_22172_new_n2783_; 
wire core__abc_22172_new_n2784_; 
wire core__abc_22172_new_n2786_; 
wire core__abc_22172_new_n2787_; 
wire core__abc_22172_new_n2788_; 
wire core__abc_22172_new_n2790_; 
wire core__abc_22172_new_n2791_; 
wire core__abc_22172_new_n2792_; 
wire core__abc_22172_new_n2794_; 
wire core__abc_22172_new_n2795_; 
wire core__abc_22172_new_n2796_; 
wire core__abc_22172_new_n2798_; 
wire core__abc_22172_new_n2799_; 
wire core__abc_22172_new_n2800_; 
wire core__abc_22172_new_n2802_; 
wire core__abc_22172_new_n2803_; 
wire core__abc_22172_new_n2804_; 
wire core__abc_22172_new_n2806_; 
wire core__abc_22172_new_n2807_; 
wire core__abc_22172_new_n2808_; 
wire core__abc_22172_new_n2810_; 
wire core__abc_22172_new_n2811_; 
wire core__abc_22172_new_n2812_; 
wire core__abc_22172_new_n2814_; 
wire core__abc_22172_new_n2815_; 
wire core__abc_22172_new_n2816_; 
wire core__abc_22172_new_n2818_; 
wire core__abc_22172_new_n2819_; 
wire core__abc_22172_new_n2820_; 
wire core__abc_22172_new_n2822_; 
wire core__abc_22172_new_n2823_; 
wire core__abc_22172_new_n2824_; 
wire core__abc_22172_new_n2826_; 
wire core__abc_22172_new_n2827_; 
wire core__abc_22172_new_n2828_; 
wire core__abc_22172_new_n2830_; 
wire core__abc_22172_new_n2831_; 
wire core__abc_22172_new_n2832_; 
wire core__abc_22172_new_n2834_; 
wire core__abc_22172_new_n2835_; 
wire core__abc_22172_new_n2836_; 
wire core__abc_22172_new_n2838_; 
wire core__abc_22172_new_n2839_; 
wire core__abc_22172_new_n2840_; 
wire core__abc_22172_new_n2842_; 
wire core__abc_22172_new_n2843_; 
wire core__abc_22172_new_n2844_; 
wire core__abc_22172_new_n2846_; 
wire core__abc_22172_new_n2847_; 
wire core__abc_22172_new_n2848_; 
wire core__abc_22172_new_n2850_; 
wire core__abc_22172_new_n2851_; 
wire core__abc_22172_new_n2852_; 
wire core__abc_22172_new_n2854_; 
wire core__abc_22172_new_n2855_; 
wire core__abc_22172_new_n2856_; 
wire core__abc_22172_new_n2858_; 
wire core__abc_22172_new_n2859_; 
wire core__abc_22172_new_n2860_; 
wire core__abc_22172_new_n2862_; 
wire core__abc_22172_new_n2863_; 
wire core__abc_22172_new_n2864_; 
wire core__abc_22172_new_n2866_; 
wire core__abc_22172_new_n2867_; 
wire core__abc_22172_new_n2868_; 
wire core__abc_22172_new_n2870_; 
wire core__abc_22172_new_n2871_; 
wire core__abc_22172_new_n2872_; 
wire core__abc_22172_new_n2874_; 
wire core__abc_22172_new_n2875_; 
wire core__abc_22172_new_n2876_; 
wire core__abc_22172_new_n2878_; 
wire core__abc_22172_new_n2879_; 
wire core__abc_22172_new_n2880_; 
wire core__abc_22172_new_n2882_; 
wire core__abc_22172_new_n2883_; 
wire core__abc_22172_new_n2884_; 
wire core__abc_22172_new_n2886_; 
wire core__abc_22172_new_n2887_; 
wire core__abc_22172_new_n2888_; 
wire core__abc_22172_new_n2890_; 
wire core__abc_22172_new_n2891_; 
wire core__abc_22172_new_n2892_; 
wire core__abc_22172_new_n2894_; 
wire core__abc_22172_new_n2895_; 
wire core__abc_22172_new_n2896_; 
wire core__abc_22172_new_n2898_; 
wire core__abc_22172_new_n2899_; 
wire core__abc_22172_new_n2900_; 
wire core__abc_22172_new_n2902_; 
wire core__abc_22172_new_n2903_; 
wire core__abc_22172_new_n2904_; 
wire core__abc_22172_new_n2906_; 
wire core__abc_22172_new_n2907_; 
wire core__abc_22172_new_n2908_; 
wire core__abc_22172_new_n2910_; 
wire core__abc_22172_new_n2911_; 
wire core__abc_22172_new_n2912_; 
wire core__abc_22172_new_n2914_; 
wire core__abc_22172_new_n2915_; 
wire core__abc_22172_new_n2916_; 
wire core__abc_22172_new_n2918_; 
wire core__abc_22172_new_n2919_; 
wire core__abc_22172_new_n2920_; 
wire core__abc_22172_new_n2921_; 
wire core__abc_22172_new_n2922_; 
wire core__abc_22172_new_n2923_; 
wire core__abc_22172_new_n2924_; 
wire core__abc_22172_new_n2925_; 
wire core__abc_22172_new_n2926_; 
wire core__abc_22172_new_n2927_; 
wire core__abc_22172_new_n2928_; 
wire core__abc_22172_new_n2929_; 
wire core__abc_22172_new_n2930_; 
wire core__abc_22172_new_n2931_; 
wire core__abc_22172_new_n2932_; 
wire core__abc_22172_new_n2933_; 
wire core__abc_22172_new_n2934_; 
wire core__abc_22172_new_n2935_; 
wire core__abc_22172_new_n2936_; 
wire core__abc_22172_new_n2937_; 
wire core__abc_22172_new_n2938_; 
wire core__abc_22172_new_n2939_; 
wire core__abc_22172_new_n2940_; 
wire core__abc_22172_new_n2941_; 
wire core__abc_22172_new_n2942_; 
wire core__abc_22172_new_n2943_; 
wire core__abc_22172_new_n2944_; 
wire core__abc_22172_new_n2945_; 
wire core__abc_22172_new_n2946_; 
wire core__abc_22172_new_n2947_; 
wire core__abc_22172_new_n2948_; 
wire core__abc_22172_new_n2949_; 
wire core__abc_22172_new_n2950_; 
wire core__abc_22172_new_n2951_; 
wire core__abc_22172_new_n2952_; 
wire core__abc_22172_new_n2953_; 
wire core__abc_22172_new_n2954_; 
wire core__abc_22172_new_n2955_; 
wire core__abc_22172_new_n2956_; 
wire core__abc_22172_new_n2957_; 
wire core__abc_22172_new_n2958_; 
wire core__abc_22172_new_n2959_; 
wire core__abc_22172_new_n2960_; 
wire core__abc_22172_new_n2961_; 
wire core__abc_22172_new_n2962_; 
wire core__abc_22172_new_n2963_; 
wire core__abc_22172_new_n2964_; 
wire core__abc_22172_new_n2965_; 
wire core__abc_22172_new_n2966_; 
wire core__abc_22172_new_n2967_; 
wire core__abc_22172_new_n2968_; 
wire core__abc_22172_new_n2969_; 
wire core__abc_22172_new_n2970_; 
wire core__abc_22172_new_n2971_; 
wire core__abc_22172_new_n2972_; 
wire core__abc_22172_new_n2973_; 
wire core__abc_22172_new_n2974_; 
wire core__abc_22172_new_n2975_; 
wire core__abc_22172_new_n2976_; 
wire core__abc_22172_new_n2977_; 
wire core__abc_22172_new_n2978_; 
wire core__abc_22172_new_n2979_; 
wire core__abc_22172_new_n2980_; 
wire core__abc_22172_new_n2981_; 
wire core__abc_22172_new_n2982_; 
wire core__abc_22172_new_n2983_; 
wire core__abc_22172_new_n2984_; 
wire core__abc_22172_new_n2985_; 
wire core__abc_22172_new_n2986_; 
wire core__abc_22172_new_n2987_; 
wire core__abc_22172_new_n2988_; 
wire core__abc_22172_new_n2989_; 
wire core__abc_22172_new_n2990_; 
wire core__abc_22172_new_n2991_; 
wire core__abc_22172_new_n2992_; 
wire core__abc_22172_new_n2993_; 
wire core__abc_22172_new_n2994_; 
wire core__abc_22172_new_n2995_; 
wire core__abc_22172_new_n2996_; 
wire core__abc_22172_new_n2997_; 
wire core__abc_22172_new_n2998_; 
wire core__abc_22172_new_n2999_; 
wire core__abc_22172_new_n3000_; 
wire core__abc_22172_new_n3001_; 
wire core__abc_22172_new_n3002_; 
wire core__abc_22172_new_n3003_; 
wire core__abc_22172_new_n3004_; 
wire core__abc_22172_new_n3005_; 
wire core__abc_22172_new_n3006_; 
wire core__abc_22172_new_n3007_; 
wire core__abc_22172_new_n3008_; 
wire core__abc_22172_new_n3009_; 
wire core__abc_22172_new_n3010_; 
wire core__abc_22172_new_n3011_; 
wire core__abc_22172_new_n3012_; 
wire core__abc_22172_new_n3013_; 
wire core__abc_22172_new_n3014_; 
wire core__abc_22172_new_n3015_; 
wire core__abc_22172_new_n3016_; 
wire core__abc_22172_new_n3017_; 
wire core__abc_22172_new_n3018_; 
wire core__abc_22172_new_n3019_; 
wire core__abc_22172_new_n3020_; 
wire core__abc_22172_new_n3021_; 
wire core__abc_22172_new_n3022_; 
wire core__abc_22172_new_n3023_; 
wire core__abc_22172_new_n3024_; 
wire core__abc_22172_new_n3025_; 
wire core__abc_22172_new_n3026_; 
wire core__abc_22172_new_n3027_; 
wire core__abc_22172_new_n3028_; 
wire core__abc_22172_new_n3029_; 
wire core__abc_22172_new_n3030_; 
wire core__abc_22172_new_n3031_; 
wire core__abc_22172_new_n3032_; 
wire core__abc_22172_new_n3033_; 
wire core__abc_22172_new_n3034_; 
wire core__abc_22172_new_n3035_; 
wire core__abc_22172_new_n3036_; 
wire core__abc_22172_new_n3037_; 
wire core__abc_22172_new_n3038_; 
wire core__abc_22172_new_n3039_; 
wire core__abc_22172_new_n3040_; 
wire core__abc_22172_new_n3041_; 
wire core__abc_22172_new_n3042_; 
wire core__abc_22172_new_n3043_; 
wire core__abc_22172_new_n3044_; 
wire core__abc_22172_new_n3045_; 
wire core__abc_22172_new_n3046_; 
wire core__abc_22172_new_n3047_; 
wire core__abc_22172_new_n3048_; 
wire core__abc_22172_new_n3049_; 
wire core__abc_22172_new_n3050_; 
wire core__abc_22172_new_n3051_; 
wire core__abc_22172_new_n3052_; 
wire core__abc_22172_new_n3053_; 
wire core__abc_22172_new_n3054_; 
wire core__abc_22172_new_n3055_; 
wire core__abc_22172_new_n3056_; 
wire core__abc_22172_new_n3057_; 
wire core__abc_22172_new_n3058_; 
wire core__abc_22172_new_n3059_; 
wire core__abc_22172_new_n3060_; 
wire core__abc_22172_new_n3061_; 
wire core__abc_22172_new_n3062_; 
wire core__abc_22172_new_n3063_; 
wire core__abc_22172_new_n3064_; 
wire core__abc_22172_new_n3065_; 
wire core__abc_22172_new_n3066_; 
wire core__abc_22172_new_n3067_; 
wire core__abc_22172_new_n3068_; 
wire core__abc_22172_new_n3069_; 
wire core__abc_22172_new_n3070_; 
wire core__abc_22172_new_n3071_; 
wire core__abc_22172_new_n3072_; 
wire core__abc_22172_new_n3073_; 
wire core__abc_22172_new_n3074_; 
wire core__abc_22172_new_n3075_; 
wire core__abc_22172_new_n3076_; 
wire core__abc_22172_new_n3077_; 
wire core__abc_22172_new_n3078_; 
wire core__abc_22172_new_n3079_; 
wire core__abc_22172_new_n3080_; 
wire core__abc_22172_new_n3081_; 
wire core__abc_22172_new_n3082_; 
wire core__abc_22172_new_n3083_; 
wire core__abc_22172_new_n3084_; 
wire core__abc_22172_new_n3085_; 
wire core__abc_22172_new_n3086_; 
wire core__abc_22172_new_n3087_; 
wire core__abc_22172_new_n3088_; 
wire core__abc_22172_new_n3089_; 
wire core__abc_22172_new_n3090_; 
wire core__abc_22172_new_n3091_; 
wire core__abc_22172_new_n3092_; 
wire core__abc_22172_new_n3093_; 
wire core__abc_22172_new_n3094_; 
wire core__abc_22172_new_n3095_; 
wire core__abc_22172_new_n3096_; 
wire core__abc_22172_new_n3097_; 
wire core__abc_22172_new_n3098_; 
wire core__abc_22172_new_n3099_; 
wire core__abc_22172_new_n3100_; 
wire core__abc_22172_new_n3101_; 
wire core__abc_22172_new_n3102_; 
wire core__abc_22172_new_n3103_; 
wire core__abc_22172_new_n3104_; 
wire core__abc_22172_new_n3105_; 
wire core__abc_22172_new_n3106_; 
wire core__abc_22172_new_n3107_; 
wire core__abc_22172_new_n3108_; 
wire core__abc_22172_new_n3109_; 
wire core__abc_22172_new_n3110_; 
wire core__abc_22172_new_n3111_; 
wire core__abc_22172_new_n3112_; 
wire core__abc_22172_new_n3113_; 
wire core__abc_22172_new_n3114_; 
wire core__abc_22172_new_n3115_; 
wire core__abc_22172_new_n3116_; 
wire core__abc_22172_new_n3117_; 
wire core__abc_22172_new_n3118_; 
wire core__abc_22172_new_n3119_; 
wire core__abc_22172_new_n3120_; 
wire core__abc_22172_new_n3121_; 
wire core__abc_22172_new_n3122_; 
wire core__abc_22172_new_n3123_; 
wire core__abc_22172_new_n3124_; 
wire core__abc_22172_new_n3125_; 
wire core__abc_22172_new_n3126_; 
wire core__abc_22172_new_n3127_; 
wire core__abc_22172_new_n3128_; 
wire core__abc_22172_new_n3129_; 
wire core__abc_22172_new_n3130_; 
wire core__abc_22172_new_n3131_; 
wire core__abc_22172_new_n3132_; 
wire core__abc_22172_new_n3133_; 
wire core__abc_22172_new_n3134_; 
wire core__abc_22172_new_n3135_; 
wire core__abc_22172_new_n3136_; 
wire core__abc_22172_new_n3137_; 
wire core__abc_22172_new_n3138_; 
wire core__abc_22172_new_n3139_; 
wire core__abc_22172_new_n3140_; 
wire core__abc_22172_new_n3141_; 
wire core__abc_22172_new_n3142_; 
wire core__abc_22172_new_n3143_; 
wire core__abc_22172_new_n3144_; 
wire core__abc_22172_new_n3145_; 
wire core__abc_22172_new_n3146_; 
wire core__abc_22172_new_n3147_; 
wire core__abc_22172_new_n3148_; 
wire core__abc_22172_new_n3149_; 
wire core__abc_22172_new_n3150_; 
wire core__abc_22172_new_n3151_; 
wire core__abc_22172_new_n3152_; 
wire core__abc_22172_new_n3153_; 
wire core__abc_22172_new_n3154_; 
wire core__abc_22172_new_n3155_; 
wire core__abc_22172_new_n3156_; 
wire core__abc_22172_new_n3157_; 
wire core__abc_22172_new_n3158_; 
wire core__abc_22172_new_n3159_; 
wire core__abc_22172_new_n3160_; 
wire core__abc_22172_new_n3161_; 
wire core__abc_22172_new_n3162_; 
wire core__abc_22172_new_n3163_; 
wire core__abc_22172_new_n3164_; 
wire core__abc_22172_new_n3165_; 
wire core__abc_22172_new_n3166_; 
wire core__abc_22172_new_n3167_; 
wire core__abc_22172_new_n3168_; 
wire core__abc_22172_new_n3169_; 
wire core__abc_22172_new_n3170_; 
wire core__abc_22172_new_n3171_; 
wire core__abc_22172_new_n3172_; 
wire core__abc_22172_new_n3173_; 
wire core__abc_22172_new_n3174_; 
wire core__abc_22172_new_n3175_; 
wire core__abc_22172_new_n3176_; 
wire core__abc_22172_new_n3177_; 
wire core__abc_22172_new_n3178_; 
wire core__abc_22172_new_n3179_; 
wire core__abc_22172_new_n3180_; 
wire core__abc_22172_new_n3181_; 
wire core__abc_22172_new_n3182_; 
wire core__abc_22172_new_n3183_; 
wire core__abc_22172_new_n3184_; 
wire core__abc_22172_new_n3185_; 
wire core__abc_22172_new_n3186_; 
wire core__abc_22172_new_n3187_; 
wire core__abc_22172_new_n3188_; 
wire core__abc_22172_new_n3189_; 
wire core__abc_22172_new_n3190_; 
wire core__abc_22172_new_n3191_; 
wire core__abc_22172_new_n3192_; 
wire core__abc_22172_new_n3193_; 
wire core__abc_22172_new_n3194_; 
wire core__abc_22172_new_n3195_; 
wire core__abc_22172_new_n3196_; 
wire core__abc_22172_new_n3197_; 
wire core__abc_22172_new_n3198_; 
wire core__abc_22172_new_n3199_; 
wire core__abc_22172_new_n3200_; 
wire core__abc_22172_new_n3201_; 
wire core__abc_22172_new_n3202_; 
wire core__abc_22172_new_n3203_; 
wire core__abc_22172_new_n3204_; 
wire core__abc_22172_new_n3205_; 
wire core__abc_22172_new_n3206_; 
wire core__abc_22172_new_n3207_; 
wire core__abc_22172_new_n3208_; 
wire core__abc_22172_new_n3209_; 
wire core__abc_22172_new_n3210_; 
wire core__abc_22172_new_n3211_; 
wire core__abc_22172_new_n3212_; 
wire core__abc_22172_new_n3213_; 
wire core__abc_22172_new_n3214_; 
wire core__abc_22172_new_n3215_; 
wire core__abc_22172_new_n3216_; 
wire core__abc_22172_new_n3217_; 
wire core__abc_22172_new_n3218_; 
wire core__abc_22172_new_n3219_; 
wire core__abc_22172_new_n3220_; 
wire core__abc_22172_new_n3221_; 
wire core__abc_22172_new_n3222_; 
wire core__abc_22172_new_n3223_; 
wire core__abc_22172_new_n3224_; 
wire core__abc_22172_new_n3225_; 
wire core__abc_22172_new_n3226_; 
wire core__abc_22172_new_n3227_; 
wire core__abc_22172_new_n3228_; 
wire core__abc_22172_new_n3229_; 
wire core__abc_22172_new_n3230_; 
wire core__abc_22172_new_n3232_; 
wire core__abc_22172_new_n3233_; 
wire core__abc_22172_new_n3234_; 
wire core__abc_22172_new_n3235_; 
wire core__abc_22172_new_n3236_; 
wire core__abc_22172_new_n3237_; 
wire core__abc_22172_new_n3238_; 
wire core__abc_22172_new_n3239_; 
wire core__abc_22172_new_n3240_; 
wire core__abc_22172_new_n3241_; 
wire core__abc_22172_new_n3242_; 
wire core__abc_22172_new_n3243_; 
wire core__abc_22172_new_n3244_; 
wire core__abc_22172_new_n3245_; 
wire core__abc_22172_new_n3246_; 
wire core__abc_22172_new_n3247_; 
wire core__abc_22172_new_n3248_; 
wire core__abc_22172_new_n3249_; 
wire core__abc_22172_new_n3250_; 
wire core__abc_22172_new_n3251_; 
wire core__abc_22172_new_n3252_; 
wire core__abc_22172_new_n3253_; 
wire core__abc_22172_new_n3254_; 
wire core__abc_22172_new_n3255_; 
wire core__abc_22172_new_n3256_; 
wire core__abc_22172_new_n3257_; 
wire core__abc_22172_new_n3258_; 
wire core__abc_22172_new_n3259_; 
wire core__abc_22172_new_n3260_; 
wire core__abc_22172_new_n3261_; 
wire core__abc_22172_new_n3262_; 
wire core__abc_22172_new_n3263_; 
wire core__abc_22172_new_n3264_; 
wire core__abc_22172_new_n3265_; 
wire core__abc_22172_new_n3266_; 
wire core__abc_22172_new_n3267_; 
wire core__abc_22172_new_n3268_; 
wire core__abc_22172_new_n3269_; 
wire core__abc_22172_new_n3270_; 
wire core__abc_22172_new_n3271_; 
wire core__abc_22172_new_n3272_; 
wire core__abc_22172_new_n3273_; 
wire core__abc_22172_new_n3274_; 
wire core__abc_22172_new_n3275_; 
wire core__abc_22172_new_n3276_; 
wire core__abc_22172_new_n3277_; 
wire core__abc_22172_new_n3278_; 
wire core__abc_22172_new_n3279_; 
wire core__abc_22172_new_n3280_; 
wire core__abc_22172_new_n3281_; 
wire core__abc_22172_new_n3282_; 
wire core__abc_22172_new_n3283_; 
wire core__abc_22172_new_n3284_; 
wire core__abc_22172_new_n3285_; 
wire core__abc_22172_new_n3286_; 
wire core__abc_22172_new_n3287_; 
wire core__abc_22172_new_n3288_; 
wire core__abc_22172_new_n3289_; 
wire core__abc_22172_new_n3290_; 
wire core__abc_22172_new_n3292_; 
wire core__abc_22172_new_n3293_; 
wire core__abc_22172_new_n3294_; 
wire core__abc_22172_new_n3295_; 
wire core__abc_22172_new_n3296_; 
wire core__abc_22172_new_n3297_; 
wire core__abc_22172_new_n3298_; 
wire core__abc_22172_new_n3299_; 
wire core__abc_22172_new_n3300_; 
wire core__abc_22172_new_n3301_; 
wire core__abc_22172_new_n3302_; 
wire core__abc_22172_new_n3303_; 
wire core__abc_22172_new_n3304_; 
wire core__abc_22172_new_n3305_; 
wire core__abc_22172_new_n3306_; 
wire core__abc_22172_new_n3307_; 
wire core__abc_22172_new_n3308_; 
wire core__abc_22172_new_n3309_; 
wire core__abc_22172_new_n3310_; 
wire core__abc_22172_new_n3311_; 
wire core__abc_22172_new_n3312_; 
wire core__abc_22172_new_n3313_; 
wire core__abc_22172_new_n3314_; 
wire core__abc_22172_new_n3315_; 
wire core__abc_22172_new_n3316_; 
wire core__abc_22172_new_n3317_; 
wire core__abc_22172_new_n3318_; 
wire core__abc_22172_new_n3319_; 
wire core__abc_22172_new_n3320_; 
wire core__abc_22172_new_n3321_; 
wire core__abc_22172_new_n3322_; 
wire core__abc_22172_new_n3323_; 
wire core__abc_22172_new_n3324_; 
wire core__abc_22172_new_n3325_; 
wire core__abc_22172_new_n3326_; 
wire core__abc_22172_new_n3327_; 
wire core__abc_22172_new_n3328_; 
wire core__abc_22172_new_n3329_; 
wire core__abc_22172_new_n3330_; 
wire core__abc_22172_new_n3331_; 
wire core__abc_22172_new_n3332_; 
wire core__abc_22172_new_n3333_; 
wire core__abc_22172_new_n3334_; 
wire core__abc_22172_new_n3335_; 
wire core__abc_22172_new_n3336_; 
wire core__abc_22172_new_n3337_; 
wire core__abc_22172_new_n3338_; 
wire core__abc_22172_new_n3339_; 
wire core__abc_22172_new_n3340_; 
wire core__abc_22172_new_n3341_; 
wire core__abc_22172_new_n3342_; 
wire core__abc_22172_new_n3343_; 
wire core__abc_22172_new_n3344_; 
wire core__abc_22172_new_n3345_; 
wire core__abc_22172_new_n3346_; 
wire core__abc_22172_new_n3348_; 
wire core__abc_22172_new_n3349_; 
wire core__abc_22172_new_n3350_; 
wire core__abc_22172_new_n3351_; 
wire core__abc_22172_new_n3352_; 
wire core__abc_22172_new_n3353_; 
wire core__abc_22172_new_n3354_; 
wire core__abc_22172_new_n3355_; 
wire core__abc_22172_new_n3356_; 
wire core__abc_22172_new_n3357_; 
wire core__abc_22172_new_n3358_; 
wire core__abc_22172_new_n3359_; 
wire core__abc_22172_new_n3360_; 
wire core__abc_22172_new_n3361_; 
wire core__abc_22172_new_n3362_; 
wire core__abc_22172_new_n3363_; 
wire core__abc_22172_new_n3364_; 
wire core__abc_22172_new_n3365_; 
wire core__abc_22172_new_n3366_; 
wire core__abc_22172_new_n3367_; 
wire core__abc_22172_new_n3368_; 
wire core__abc_22172_new_n3369_; 
wire core__abc_22172_new_n3370_; 
wire core__abc_22172_new_n3371_; 
wire core__abc_22172_new_n3372_; 
wire core__abc_22172_new_n3373_; 
wire core__abc_22172_new_n3374_; 
wire core__abc_22172_new_n3375_; 
wire core__abc_22172_new_n3376_; 
wire core__abc_22172_new_n3377_; 
wire core__abc_22172_new_n3378_; 
wire core__abc_22172_new_n3379_; 
wire core__abc_22172_new_n3380_; 
wire core__abc_22172_new_n3381_; 
wire core__abc_22172_new_n3382_; 
wire core__abc_22172_new_n3383_; 
wire core__abc_22172_new_n3384_; 
wire core__abc_22172_new_n3385_; 
wire core__abc_22172_new_n3386_; 
wire core__abc_22172_new_n3387_; 
wire core__abc_22172_new_n3388_; 
wire core__abc_22172_new_n3389_; 
wire core__abc_22172_new_n3390_; 
wire core__abc_22172_new_n3391_; 
wire core__abc_22172_new_n3392_; 
wire core__abc_22172_new_n3393_; 
wire core__abc_22172_new_n3394_; 
wire core__abc_22172_new_n3395_; 
wire core__abc_22172_new_n3396_; 
wire core__abc_22172_new_n3397_; 
wire core__abc_22172_new_n3398_; 
wire core__abc_22172_new_n3399_; 
wire core__abc_22172_new_n3400_; 
wire core__abc_22172_new_n3401_; 
wire core__abc_22172_new_n3402_; 
wire core__abc_22172_new_n3403_; 
wire core__abc_22172_new_n3404_; 
wire core__abc_22172_new_n3405_; 
wire core__abc_22172_new_n3406_; 
wire core__abc_22172_new_n3407_; 
wire core__abc_22172_new_n3408_; 
wire core__abc_22172_new_n3409_; 
wire core__abc_22172_new_n3411_; 
wire core__abc_22172_new_n3412_; 
wire core__abc_22172_new_n3413_; 
wire core__abc_22172_new_n3414_; 
wire core__abc_22172_new_n3415_; 
wire core__abc_22172_new_n3416_; 
wire core__abc_22172_new_n3417_; 
wire core__abc_22172_new_n3418_; 
wire core__abc_22172_new_n3419_; 
wire core__abc_22172_new_n3420_; 
wire core__abc_22172_new_n3421_; 
wire core__abc_22172_new_n3422_; 
wire core__abc_22172_new_n3423_; 
wire core__abc_22172_new_n3424_; 
wire core__abc_22172_new_n3425_; 
wire core__abc_22172_new_n3426_; 
wire core__abc_22172_new_n3427_; 
wire core__abc_22172_new_n3428_; 
wire core__abc_22172_new_n3429_; 
wire core__abc_22172_new_n3430_; 
wire core__abc_22172_new_n3431_; 
wire core__abc_22172_new_n3432_; 
wire core__abc_22172_new_n3433_; 
wire core__abc_22172_new_n3434_; 
wire core__abc_22172_new_n3435_; 
wire core__abc_22172_new_n3436_; 
wire core__abc_22172_new_n3437_; 
wire core__abc_22172_new_n3438_; 
wire core__abc_22172_new_n3439_; 
wire core__abc_22172_new_n3440_; 
wire core__abc_22172_new_n3441_; 
wire core__abc_22172_new_n3442_; 
wire core__abc_22172_new_n3443_; 
wire core__abc_22172_new_n3444_; 
wire core__abc_22172_new_n3445_; 
wire core__abc_22172_new_n3446_; 
wire core__abc_22172_new_n3447_; 
wire core__abc_22172_new_n3448_; 
wire core__abc_22172_new_n3449_; 
wire core__abc_22172_new_n3450_; 
wire core__abc_22172_new_n3451_; 
wire core__abc_22172_new_n3452_; 
wire core__abc_22172_new_n3453_; 
wire core__abc_22172_new_n3454_; 
wire core__abc_22172_new_n3455_; 
wire core__abc_22172_new_n3456_; 
wire core__abc_22172_new_n3457_; 
wire core__abc_22172_new_n3458_; 
wire core__abc_22172_new_n3459_; 
wire core__abc_22172_new_n3460_; 
wire core__abc_22172_new_n3461_; 
wire core__abc_22172_new_n3462_; 
wire core__abc_22172_new_n3463_; 
wire core__abc_22172_new_n3464_; 
wire core__abc_22172_new_n3465_; 
wire core__abc_22172_new_n3466_; 
wire core__abc_22172_new_n3467_; 
wire core__abc_22172_new_n3468_; 
wire core__abc_22172_new_n3469_; 
wire core__abc_22172_new_n3470_; 
wire core__abc_22172_new_n3471_; 
wire core__abc_22172_new_n3472_; 
wire core__abc_22172_new_n3474_; 
wire core__abc_22172_new_n3475_; 
wire core__abc_22172_new_n3476_; 
wire core__abc_22172_new_n3477_; 
wire core__abc_22172_new_n3478_; 
wire core__abc_22172_new_n3479_; 
wire core__abc_22172_new_n3480_; 
wire core__abc_22172_new_n3481_; 
wire core__abc_22172_new_n3482_; 
wire core__abc_22172_new_n3483_; 
wire core__abc_22172_new_n3484_; 
wire core__abc_22172_new_n3485_; 
wire core__abc_22172_new_n3486_; 
wire core__abc_22172_new_n3487_; 
wire core__abc_22172_new_n3488_; 
wire core__abc_22172_new_n3489_; 
wire core__abc_22172_new_n3490_; 
wire core__abc_22172_new_n3491_; 
wire core__abc_22172_new_n3492_; 
wire core__abc_22172_new_n3493_; 
wire core__abc_22172_new_n3494_; 
wire core__abc_22172_new_n3495_; 
wire core__abc_22172_new_n3496_; 
wire core__abc_22172_new_n3497_; 
wire core__abc_22172_new_n3498_; 
wire core__abc_22172_new_n3499_; 
wire core__abc_22172_new_n3500_; 
wire core__abc_22172_new_n3501_; 
wire core__abc_22172_new_n3502_; 
wire core__abc_22172_new_n3503_; 
wire core__abc_22172_new_n3504_; 
wire core__abc_22172_new_n3505_; 
wire core__abc_22172_new_n3506_; 
wire core__abc_22172_new_n3507_; 
wire core__abc_22172_new_n3508_; 
wire core__abc_22172_new_n3509_; 
wire core__abc_22172_new_n3510_; 
wire core__abc_22172_new_n3511_; 
wire core__abc_22172_new_n3512_; 
wire core__abc_22172_new_n3513_; 
wire core__abc_22172_new_n3514_; 
wire core__abc_22172_new_n3515_; 
wire core__abc_22172_new_n3516_; 
wire core__abc_22172_new_n3517_; 
wire core__abc_22172_new_n3518_; 
wire core__abc_22172_new_n3519_; 
wire core__abc_22172_new_n3520_; 
wire core__abc_22172_new_n3521_; 
wire core__abc_22172_new_n3522_; 
wire core__abc_22172_new_n3523_; 
wire core__abc_22172_new_n3524_; 
wire core__abc_22172_new_n3525_; 
wire core__abc_22172_new_n3526_; 
wire core__abc_22172_new_n3527_; 
wire core__abc_22172_new_n3528_; 
wire core__abc_22172_new_n3529_; 
wire core__abc_22172_new_n3530_; 
wire core__abc_22172_new_n3531_; 
wire core__abc_22172_new_n3532_; 
wire core__abc_22172_new_n3533_; 
wire core__abc_22172_new_n3534_; 
wire core__abc_22172_new_n3535_; 
wire core__abc_22172_new_n3536_; 
wire core__abc_22172_new_n3538_; 
wire core__abc_22172_new_n3539_; 
wire core__abc_22172_new_n3540_; 
wire core__abc_22172_new_n3541_; 
wire core__abc_22172_new_n3542_; 
wire core__abc_22172_new_n3543_; 
wire core__abc_22172_new_n3544_; 
wire core__abc_22172_new_n3545_; 
wire core__abc_22172_new_n3546_; 
wire core__abc_22172_new_n3547_; 
wire core__abc_22172_new_n3548_; 
wire core__abc_22172_new_n3549_; 
wire core__abc_22172_new_n3550_; 
wire core__abc_22172_new_n3551_; 
wire core__abc_22172_new_n3552_; 
wire core__abc_22172_new_n3553_; 
wire core__abc_22172_new_n3554_; 
wire core__abc_22172_new_n3555_; 
wire core__abc_22172_new_n3556_; 
wire core__abc_22172_new_n3557_; 
wire core__abc_22172_new_n3558_; 
wire core__abc_22172_new_n3559_; 
wire core__abc_22172_new_n3560_; 
wire core__abc_22172_new_n3561_; 
wire core__abc_22172_new_n3562_; 
wire core__abc_22172_new_n3563_; 
wire core__abc_22172_new_n3564_; 
wire core__abc_22172_new_n3565_; 
wire core__abc_22172_new_n3566_; 
wire core__abc_22172_new_n3567_; 
wire core__abc_22172_new_n3568_; 
wire core__abc_22172_new_n3569_; 
wire core__abc_22172_new_n3570_; 
wire core__abc_22172_new_n3571_; 
wire core__abc_22172_new_n3572_; 
wire core__abc_22172_new_n3573_; 
wire core__abc_22172_new_n3574_; 
wire core__abc_22172_new_n3575_; 
wire core__abc_22172_new_n3576_; 
wire core__abc_22172_new_n3577_; 
wire core__abc_22172_new_n3578_; 
wire core__abc_22172_new_n3579_; 
wire core__abc_22172_new_n3580_; 
wire core__abc_22172_new_n3581_; 
wire core__abc_22172_new_n3582_; 
wire core__abc_22172_new_n3583_; 
wire core__abc_22172_new_n3584_; 
wire core__abc_22172_new_n3585_; 
wire core__abc_22172_new_n3586_; 
wire core__abc_22172_new_n3587_; 
wire core__abc_22172_new_n3588_; 
wire core__abc_22172_new_n3589_; 
wire core__abc_22172_new_n3590_; 
wire core__abc_22172_new_n3591_; 
wire core__abc_22172_new_n3592_; 
wire core__abc_22172_new_n3593_; 
wire core__abc_22172_new_n3594_; 
wire core__abc_22172_new_n3595_; 
wire core__abc_22172_new_n3596_; 
wire core__abc_22172_new_n3597_; 
wire core__abc_22172_new_n3598_; 
wire core__abc_22172_new_n3599_; 
wire core__abc_22172_new_n3600_; 
wire core__abc_22172_new_n3601_; 
wire core__abc_22172_new_n3602_; 
wire core__abc_22172_new_n3603_; 
wire core__abc_22172_new_n3605_; 
wire core__abc_22172_new_n3606_; 
wire core__abc_22172_new_n3607_; 
wire core__abc_22172_new_n3608_; 
wire core__abc_22172_new_n3609_; 
wire core__abc_22172_new_n3610_; 
wire core__abc_22172_new_n3611_; 
wire core__abc_22172_new_n3612_; 
wire core__abc_22172_new_n3613_; 
wire core__abc_22172_new_n3614_; 
wire core__abc_22172_new_n3615_; 
wire core__abc_22172_new_n3616_; 
wire core__abc_22172_new_n3617_; 
wire core__abc_22172_new_n3618_; 
wire core__abc_22172_new_n3619_; 
wire core__abc_22172_new_n3620_; 
wire core__abc_22172_new_n3621_; 
wire core__abc_22172_new_n3622_; 
wire core__abc_22172_new_n3623_; 
wire core__abc_22172_new_n3624_; 
wire core__abc_22172_new_n3625_; 
wire core__abc_22172_new_n3626_; 
wire core__abc_22172_new_n3627_; 
wire core__abc_22172_new_n3628_; 
wire core__abc_22172_new_n3629_; 
wire core__abc_22172_new_n3630_; 
wire core__abc_22172_new_n3631_; 
wire core__abc_22172_new_n3632_; 
wire core__abc_22172_new_n3633_; 
wire core__abc_22172_new_n3634_; 
wire core__abc_22172_new_n3635_; 
wire core__abc_22172_new_n3636_; 
wire core__abc_22172_new_n3637_; 
wire core__abc_22172_new_n3638_; 
wire core__abc_22172_new_n3639_; 
wire core__abc_22172_new_n3640_; 
wire core__abc_22172_new_n3641_; 
wire core__abc_22172_new_n3642_; 
wire core__abc_22172_new_n3643_; 
wire core__abc_22172_new_n3644_; 
wire core__abc_22172_new_n3645_; 
wire core__abc_22172_new_n3646_; 
wire core__abc_22172_new_n3647_; 
wire core__abc_22172_new_n3648_; 
wire core__abc_22172_new_n3649_; 
wire core__abc_22172_new_n3650_; 
wire core__abc_22172_new_n3651_; 
wire core__abc_22172_new_n3652_; 
wire core__abc_22172_new_n3653_; 
wire core__abc_22172_new_n3654_; 
wire core__abc_22172_new_n3655_; 
wire core__abc_22172_new_n3656_; 
wire core__abc_22172_new_n3657_; 
wire core__abc_22172_new_n3658_; 
wire core__abc_22172_new_n3660_; 
wire core__abc_22172_new_n3661_; 
wire core__abc_22172_new_n3662_; 
wire core__abc_22172_new_n3663_; 
wire core__abc_22172_new_n3664_; 
wire core__abc_22172_new_n3665_; 
wire core__abc_22172_new_n3666_; 
wire core__abc_22172_new_n3667_; 
wire core__abc_22172_new_n3668_; 
wire core__abc_22172_new_n3669_; 
wire core__abc_22172_new_n3670_; 
wire core__abc_22172_new_n3671_; 
wire core__abc_22172_new_n3672_; 
wire core__abc_22172_new_n3673_; 
wire core__abc_22172_new_n3674_; 
wire core__abc_22172_new_n3675_; 
wire core__abc_22172_new_n3676_; 
wire core__abc_22172_new_n3677_; 
wire core__abc_22172_new_n3678_; 
wire core__abc_22172_new_n3679_; 
wire core__abc_22172_new_n3680_; 
wire core__abc_22172_new_n3681_; 
wire core__abc_22172_new_n3682_; 
wire core__abc_22172_new_n3683_; 
wire core__abc_22172_new_n3684_; 
wire core__abc_22172_new_n3685_; 
wire core__abc_22172_new_n3686_; 
wire core__abc_22172_new_n3687_; 
wire core__abc_22172_new_n3688_; 
wire core__abc_22172_new_n3689_; 
wire core__abc_22172_new_n3690_; 
wire core__abc_22172_new_n3691_; 
wire core__abc_22172_new_n3692_; 
wire core__abc_22172_new_n3693_; 
wire core__abc_22172_new_n3694_; 
wire core__abc_22172_new_n3695_; 
wire core__abc_22172_new_n3696_; 
wire core__abc_22172_new_n3697_; 
wire core__abc_22172_new_n3698_; 
wire core__abc_22172_new_n3699_; 
wire core__abc_22172_new_n3700_; 
wire core__abc_22172_new_n3701_; 
wire core__abc_22172_new_n3702_; 
wire core__abc_22172_new_n3703_; 
wire core__abc_22172_new_n3704_; 
wire core__abc_22172_new_n3705_; 
wire core__abc_22172_new_n3706_; 
wire core__abc_22172_new_n3707_; 
wire core__abc_22172_new_n3708_; 
wire core__abc_22172_new_n3709_; 
wire core__abc_22172_new_n3710_; 
wire core__abc_22172_new_n3711_; 
wire core__abc_22172_new_n3712_; 
wire core__abc_22172_new_n3713_; 
wire core__abc_22172_new_n3714_; 
wire core__abc_22172_new_n3715_; 
wire core__abc_22172_new_n3716_; 
wire core__abc_22172_new_n3717_; 
wire core__abc_22172_new_n3718_; 
wire core__abc_22172_new_n3719_; 
wire core__abc_22172_new_n3720_; 
wire core__abc_22172_new_n3721_; 
wire core__abc_22172_new_n3722_; 
wire core__abc_22172_new_n3723_; 
wire core__abc_22172_new_n3724_; 
wire core__abc_22172_new_n3725_; 
wire core__abc_22172_new_n3726_; 
wire core__abc_22172_new_n3727_; 
wire core__abc_22172_new_n3728_; 
wire core__abc_22172_new_n3729_; 
wire core__abc_22172_new_n3730_; 
wire core__abc_22172_new_n3731_; 
wire core__abc_22172_new_n3732_; 
wire core__abc_22172_new_n3733_; 
wire core__abc_22172_new_n3735_; 
wire core__abc_22172_new_n3736_; 
wire core__abc_22172_new_n3737_; 
wire core__abc_22172_new_n3738_; 
wire core__abc_22172_new_n3739_; 
wire core__abc_22172_new_n3740_; 
wire core__abc_22172_new_n3741_; 
wire core__abc_22172_new_n3742_; 
wire core__abc_22172_new_n3743_; 
wire core__abc_22172_new_n3744_; 
wire core__abc_22172_new_n3745_; 
wire core__abc_22172_new_n3746_; 
wire core__abc_22172_new_n3747_; 
wire core__abc_22172_new_n3748_; 
wire core__abc_22172_new_n3749_; 
wire core__abc_22172_new_n3750_; 
wire core__abc_22172_new_n3751_; 
wire core__abc_22172_new_n3752_; 
wire core__abc_22172_new_n3753_; 
wire core__abc_22172_new_n3754_; 
wire core__abc_22172_new_n3755_; 
wire core__abc_22172_new_n3756_; 
wire core__abc_22172_new_n3757_; 
wire core__abc_22172_new_n3758_; 
wire core__abc_22172_new_n3759_; 
wire core__abc_22172_new_n3760_; 
wire core__abc_22172_new_n3761_; 
wire core__abc_22172_new_n3762_; 
wire core__abc_22172_new_n3763_; 
wire core__abc_22172_new_n3764_; 
wire core__abc_22172_new_n3765_; 
wire core__abc_22172_new_n3766_; 
wire core__abc_22172_new_n3767_; 
wire core__abc_22172_new_n3768_; 
wire core__abc_22172_new_n3769_; 
wire core__abc_22172_new_n3770_; 
wire core__abc_22172_new_n3771_; 
wire core__abc_22172_new_n3772_; 
wire core__abc_22172_new_n3773_; 
wire core__abc_22172_new_n3774_; 
wire core__abc_22172_new_n3775_; 
wire core__abc_22172_new_n3776_; 
wire core__abc_22172_new_n3777_; 
wire core__abc_22172_new_n3778_; 
wire core__abc_22172_new_n3779_; 
wire core__abc_22172_new_n3780_; 
wire core__abc_22172_new_n3781_; 
wire core__abc_22172_new_n3782_; 
wire core__abc_22172_new_n3783_; 
wire core__abc_22172_new_n3784_; 
wire core__abc_22172_new_n3785_; 
wire core__abc_22172_new_n3786_; 
wire core__abc_22172_new_n3787_; 
wire core__abc_22172_new_n3788_; 
wire core__abc_22172_new_n3789_; 
wire core__abc_22172_new_n3790_; 
wire core__abc_22172_new_n3791_; 
wire core__abc_22172_new_n3792_; 
wire core__abc_22172_new_n3793_; 
wire core__abc_22172_new_n3794_; 
wire core__abc_22172_new_n3795_; 
wire core__abc_22172_new_n3796_; 
wire core__abc_22172_new_n3797_; 
wire core__abc_22172_new_n3798_; 
wire core__abc_22172_new_n3799_; 
wire core__abc_22172_new_n3800_; 
wire core__abc_22172_new_n3801_; 
wire core__abc_22172_new_n3802_; 
wire core__abc_22172_new_n3804_; 
wire core__abc_22172_new_n3805_; 
wire core__abc_22172_new_n3806_; 
wire core__abc_22172_new_n3807_; 
wire core__abc_22172_new_n3808_; 
wire core__abc_22172_new_n3809_; 
wire core__abc_22172_new_n3810_; 
wire core__abc_22172_new_n3811_; 
wire core__abc_22172_new_n3812_; 
wire core__abc_22172_new_n3813_; 
wire core__abc_22172_new_n3814_; 
wire core__abc_22172_new_n3815_; 
wire core__abc_22172_new_n3816_; 
wire core__abc_22172_new_n3817_; 
wire core__abc_22172_new_n3818_; 
wire core__abc_22172_new_n3819_; 
wire core__abc_22172_new_n3820_; 
wire core__abc_22172_new_n3821_; 
wire core__abc_22172_new_n3822_; 
wire core__abc_22172_new_n3823_; 
wire core__abc_22172_new_n3824_; 
wire core__abc_22172_new_n3825_; 
wire core__abc_22172_new_n3826_; 
wire core__abc_22172_new_n3827_; 
wire core__abc_22172_new_n3828_; 
wire core__abc_22172_new_n3829_; 
wire core__abc_22172_new_n3830_; 
wire core__abc_22172_new_n3831_; 
wire core__abc_22172_new_n3832_; 
wire core__abc_22172_new_n3833_; 
wire core__abc_22172_new_n3834_; 
wire core__abc_22172_new_n3835_; 
wire core__abc_22172_new_n3836_; 
wire core__abc_22172_new_n3837_; 
wire core__abc_22172_new_n3838_; 
wire core__abc_22172_new_n3839_; 
wire core__abc_22172_new_n3840_; 
wire core__abc_22172_new_n3841_; 
wire core__abc_22172_new_n3842_; 
wire core__abc_22172_new_n3843_; 
wire core__abc_22172_new_n3844_; 
wire core__abc_22172_new_n3845_; 
wire core__abc_22172_new_n3846_; 
wire core__abc_22172_new_n3847_; 
wire core__abc_22172_new_n3848_; 
wire core__abc_22172_new_n3849_; 
wire core__abc_22172_new_n3850_; 
wire core__abc_22172_new_n3851_; 
wire core__abc_22172_new_n3852_; 
wire core__abc_22172_new_n3853_; 
wire core__abc_22172_new_n3854_; 
wire core__abc_22172_new_n3855_; 
wire core__abc_22172_new_n3856_; 
wire core__abc_22172_new_n3857_; 
wire core__abc_22172_new_n3858_; 
wire core__abc_22172_new_n3859_; 
wire core__abc_22172_new_n3860_; 
wire core__abc_22172_new_n3861_; 
wire core__abc_22172_new_n3862_; 
wire core__abc_22172_new_n3863_; 
wire core__abc_22172_new_n3864_; 
wire core__abc_22172_new_n3865_; 
wire core__abc_22172_new_n3866_; 
wire core__abc_22172_new_n3868_; 
wire core__abc_22172_new_n3869_; 
wire core__abc_22172_new_n3870_; 
wire core__abc_22172_new_n3871_; 
wire core__abc_22172_new_n3872_; 
wire core__abc_22172_new_n3873_; 
wire core__abc_22172_new_n3874_; 
wire core__abc_22172_new_n3875_; 
wire core__abc_22172_new_n3876_; 
wire core__abc_22172_new_n3877_; 
wire core__abc_22172_new_n3878_; 
wire core__abc_22172_new_n3879_; 
wire core__abc_22172_new_n3880_; 
wire core__abc_22172_new_n3881_; 
wire core__abc_22172_new_n3882_; 
wire core__abc_22172_new_n3883_; 
wire core__abc_22172_new_n3884_; 
wire core__abc_22172_new_n3885_; 
wire core__abc_22172_new_n3886_; 
wire core__abc_22172_new_n3887_; 
wire core__abc_22172_new_n3888_; 
wire core__abc_22172_new_n3889_; 
wire core__abc_22172_new_n3890_; 
wire core__abc_22172_new_n3891_; 
wire core__abc_22172_new_n3892_; 
wire core__abc_22172_new_n3893_; 
wire core__abc_22172_new_n3894_; 
wire core__abc_22172_new_n3895_; 
wire core__abc_22172_new_n3896_; 
wire core__abc_22172_new_n3897_; 
wire core__abc_22172_new_n3898_; 
wire core__abc_22172_new_n3899_; 
wire core__abc_22172_new_n3900_; 
wire core__abc_22172_new_n3901_; 
wire core__abc_22172_new_n3902_; 
wire core__abc_22172_new_n3903_; 
wire core__abc_22172_new_n3904_; 
wire core__abc_22172_new_n3905_; 
wire core__abc_22172_new_n3906_; 
wire core__abc_22172_new_n3907_; 
wire core__abc_22172_new_n3908_; 
wire core__abc_22172_new_n3909_; 
wire core__abc_22172_new_n3910_; 
wire core__abc_22172_new_n3911_; 
wire core__abc_22172_new_n3912_; 
wire core__abc_22172_new_n3913_; 
wire core__abc_22172_new_n3914_; 
wire core__abc_22172_new_n3915_; 
wire core__abc_22172_new_n3916_; 
wire core__abc_22172_new_n3917_; 
wire core__abc_22172_new_n3918_; 
wire core__abc_22172_new_n3919_; 
wire core__abc_22172_new_n3920_; 
wire core__abc_22172_new_n3921_; 
wire core__abc_22172_new_n3922_; 
wire core__abc_22172_new_n3923_; 
wire core__abc_22172_new_n3924_; 
wire core__abc_22172_new_n3926_; 
wire core__abc_22172_new_n3927_; 
wire core__abc_22172_new_n3928_; 
wire core__abc_22172_new_n3929_; 
wire core__abc_22172_new_n3930_; 
wire core__abc_22172_new_n3931_; 
wire core__abc_22172_new_n3932_; 
wire core__abc_22172_new_n3933_; 
wire core__abc_22172_new_n3934_; 
wire core__abc_22172_new_n3935_; 
wire core__abc_22172_new_n3936_; 
wire core__abc_22172_new_n3937_; 
wire core__abc_22172_new_n3938_; 
wire core__abc_22172_new_n3939_; 
wire core__abc_22172_new_n3940_; 
wire core__abc_22172_new_n3941_; 
wire core__abc_22172_new_n3942_; 
wire core__abc_22172_new_n3943_; 
wire core__abc_22172_new_n3944_; 
wire core__abc_22172_new_n3945_; 
wire core__abc_22172_new_n3946_; 
wire core__abc_22172_new_n3947_; 
wire core__abc_22172_new_n3948_; 
wire core__abc_22172_new_n3949_; 
wire core__abc_22172_new_n3950_; 
wire core__abc_22172_new_n3951_; 
wire core__abc_22172_new_n3952_; 
wire core__abc_22172_new_n3953_; 
wire core__abc_22172_new_n3954_; 
wire core__abc_22172_new_n3955_; 
wire core__abc_22172_new_n3956_; 
wire core__abc_22172_new_n3957_; 
wire core__abc_22172_new_n3958_; 
wire core__abc_22172_new_n3959_; 
wire core__abc_22172_new_n3960_; 
wire core__abc_22172_new_n3961_; 
wire core__abc_22172_new_n3962_; 
wire core__abc_22172_new_n3963_; 
wire core__abc_22172_new_n3964_; 
wire core__abc_22172_new_n3965_; 
wire core__abc_22172_new_n3966_; 
wire core__abc_22172_new_n3967_; 
wire core__abc_22172_new_n3968_; 
wire core__abc_22172_new_n3969_; 
wire core__abc_22172_new_n3970_; 
wire core__abc_22172_new_n3971_; 
wire core__abc_22172_new_n3972_; 
wire core__abc_22172_new_n3973_; 
wire core__abc_22172_new_n3974_; 
wire core__abc_22172_new_n3975_; 
wire core__abc_22172_new_n3976_; 
wire core__abc_22172_new_n3977_; 
wire core__abc_22172_new_n3978_; 
wire core__abc_22172_new_n3979_; 
wire core__abc_22172_new_n3980_; 
wire core__abc_22172_new_n3981_; 
wire core__abc_22172_new_n3982_; 
wire core__abc_22172_new_n3983_; 
wire core__abc_22172_new_n3984_; 
wire core__abc_22172_new_n3985_; 
wire core__abc_22172_new_n3986_; 
wire core__abc_22172_new_n3987_; 
wire core__abc_22172_new_n3988_; 
wire core__abc_22172_new_n3989_; 
wire core__abc_22172_new_n3990_; 
wire core__abc_22172_new_n3991_; 
wire core__abc_22172_new_n3992_; 
wire core__abc_22172_new_n3993_; 
wire core__abc_22172_new_n3994_; 
wire core__abc_22172_new_n3996_; 
wire core__abc_22172_new_n3997_; 
wire core__abc_22172_new_n3998_; 
wire core__abc_22172_new_n3999_; 
wire core__abc_22172_new_n4000_; 
wire core__abc_22172_new_n4001_; 
wire core__abc_22172_new_n4002_; 
wire core__abc_22172_new_n4003_; 
wire core__abc_22172_new_n4004_; 
wire core__abc_22172_new_n4005_; 
wire core__abc_22172_new_n4006_; 
wire core__abc_22172_new_n4007_; 
wire core__abc_22172_new_n4008_; 
wire core__abc_22172_new_n4009_; 
wire core__abc_22172_new_n4010_; 
wire core__abc_22172_new_n4011_; 
wire core__abc_22172_new_n4012_; 
wire core__abc_22172_new_n4013_; 
wire core__abc_22172_new_n4014_; 
wire core__abc_22172_new_n4015_; 
wire core__abc_22172_new_n4016_; 
wire core__abc_22172_new_n4017_; 
wire core__abc_22172_new_n4018_; 
wire core__abc_22172_new_n4019_; 
wire core__abc_22172_new_n4020_; 
wire core__abc_22172_new_n4021_; 
wire core__abc_22172_new_n4022_; 
wire core__abc_22172_new_n4023_; 
wire core__abc_22172_new_n4024_; 
wire core__abc_22172_new_n4025_; 
wire core__abc_22172_new_n4026_; 
wire core__abc_22172_new_n4027_; 
wire core__abc_22172_new_n4028_; 
wire core__abc_22172_new_n4029_; 
wire core__abc_22172_new_n4030_; 
wire core__abc_22172_new_n4031_; 
wire core__abc_22172_new_n4032_; 
wire core__abc_22172_new_n4033_; 
wire core__abc_22172_new_n4034_; 
wire core__abc_22172_new_n4035_; 
wire core__abc_22172_new_n4036_; 
wire core__abc_22172_new_n4037_; 
wire core__abc_22172_new_n4038_; 
wire core__abc_22172_new_n4039_; 
wire core__abc_22172_new_n4040_; 
wire core__abc_22172_new_n4041_; 
wire core__abc_22172_new_n4042_; 
wire core__abc_22172_new_n4043_; 
wire core__abc_22172_new_n4044_; 
wire core__abc_22172_new_n4045_; 
wire core__abc_22172_new_n4046_; 
wire core__abc_22172_new_n4047_; 
wire core__abc_22172_new_n4048_; 
wire core__abc_22172_new_n4049_; 
wire core__abc_22172_new_n4050_; 
wire core__abc_22172_new_n4051_; 
wire core__abc_22172_new_n4052_; 
wire core__abc_22172_new_n4053_; 
wire core__abc_22172_new_n4054_; 
wire core__abc_22172_new_n4055_; 
wire core__abc_22172_new_n4056_; 
wire core__abc_22172_new_n4057_; 
wire core__abc_22172_new_n4058_; 
wire core__abc_22172_new_n4059_; 
wire core__abc_22172_new_n4060_; 
wire core__abc_22172_new_n4061_; 
wire core__abc_22172_new_n4063_; 
wire core__abc_22172_new_n4064_; 
wire core__abc_22172_new_n4065_; 
wire core__abc_22172_new_n4066_; 
wire core__abc_22172_new_n4067_; 
wire core__abc_22172_new_n4068_; 
wire core__abc_22172_new_n4069_; 
wire core__abc_22172_new_n4070_; 
wire core__abc_22172_new_n4071_; 
wire core__abc_22172_new_n4072_; 
wire core__abc_22172_new_n4073_; 
wire core__abc_22172_new_n4074_; 
wire core__abc_22172_new_n4075_; 
wire core__abc_22172_new_n4076_; 
wire core__abc_22172_new_n4077_; 
wire core__abc_22172_new_n4078_; 
wire core__abc_22172_new_n4079_; 
wire core__abc_22172_new_n4080_; 
wire core__abc_22172_new_n4081_; 
wire core__abc_22172_new_n4082_; 
wire core__abc_22172_new_n4083_; 
wire core__abc_22172_new_n4084_; 
wire core__abc_22172_new_n4085_; 
wire core__abc_22172_new_n4086_; 
wire core__abc_22172_new_n4087_; 
wire core__abc_22172_new_n4088_; 
wire core__abc_22172_new_n4089_; 
wire core__abc_22172_new_n4090_; 
wire core__abc_22172_new_n4091_; 
wire core__abc_22172_new_n4092_; 
wire core__abc_22172_new_n4093_; 
wire core__abc_22172_new_n4094_; 
wire core__abc_22172_new_n4095_; 
wire core__abc_22172_new_n4096_; 
wire core__abc_22172_new_n4097_; 
wire core__abc_22172_new_n4098_; 
wire core__abc_22172_new_n4099_; 
wire core__abc_22172_new_n4100_; 
wire core__abc_22172_new_n4101_; 
wire core__abc_22172_new_n4102_; 
wire core__abc_22172_new_n4103_; 
wire core__abc_22172_new_n4104_; 
wire core__abc_22172_new_n4105_; 
wire core__abc_22172_new_n4106_; 
wire core__abc_22172_new_n4107_; 
wire core__abc_22172_new_n4108_; 
wire core__abc_22172_new_n4109_; 
wire core__abc_22172_new_n4110_; 
wire core__abc_22172_new_n4111_; 
wire core__abc_22172_new_n4112_; 
wire core__abc_22172_new_n4113_; 
wire core__abc_22172_new_n4114_; 
wire core__abc_22172_new_n4115_; 
wire core__abc_22172_new_n4116_; 
wire core__abc_22172_new_n4117_; 
wire core__abc_22172_new_n4118_; 
wire core__abc_22172_new_n4119_; 
wire core__abc_22172_new_n4120_; 
wire core__abc_22172_new_n4121_; 
wire core__abc_22172_new_n4122_; 
wire core__abc_22172_new_n4123_; 
wire core__abc_22172_new_n4124_; 
wire core__abc_22172_new_n4125_; 
wire core__abc_22172_new_n4127_; 
wire core__abc_22172_new_n4128_; 
wire core__abc_22172_new_n4129_; 
wire core__abc_22172_new_n4130_; 
wire core__abc_22172_new_n4131_; 
wire core__abc_22172_new_n4132_; 
wire core__abc_22172_new_n4133_; 
wire core__abc_22172_new_n4134_; 
wire core__abc_22172_new_n4135_; 
wire core__abc_22172_new_n4136_; 
wire core__abc_22172_new_n4137_; 
wire core__abc_22172_new_n4138_; 
wire core__abc_22172_new_n4139_; 
wire core__abc_22172_new_n4140_; 
wire core__abc_22172_new_n4141_; 
wire core__abc_22172_new_n4142_; 
wire core__abc_22172_new_n4143_; 
wire core__abc_22172_new_n4144_; 
wire core__abc_22172_new_n4145_; 
wire core__abc_22172_new_n4146_; 
wire core__abc_22172_new_n4147_; 
wire core__abc_22172_new_n4148_; 
wire core__abc_22172_new_n4149_; 
wire core__abc_22172_new_n4150_; 
wire core__abc_22172_new_n4151_; 
wire core__abc_22172_new_n4152_; 
wire core__abc_22172_new_n4153_; 
wire core__abc_22172_new_n4154_; 
wire core__abc_22172_new_n4155_; 
wire core__abc_22172_new_n4156_; 
wire core__abc_22172_new_n4157_; 
wire core__abc_22172_new_n4158_; 
wire core__abc_22172_new_n4159_; 
wire core__abc_22172_new_n4160_; 
wire core__abc_22172_new_n4161_; 
wire core__abc_22172_new_n4162_; 
wire core__abc_22172_new_n4163_; 
wire core__abc_22172_new_n4164_; 
wire core__abc_22172_new_n4165_; 
wire core__abc_22172_new_n4166_; 
wire core__abc_22172_new_n4167_; 
wire core__abc_22172_new_n4168_; 
wire core__abc_22172_new_n4169_; 
wire core__abc_22172_new_n4170_; 
wire core__abc_22172_new_n4171_; 
wire core__abc_22172_new_n4172_; 
wire core__abc_22172_new_n4173_; 
wire core__abc_22172_new_n4174_; 
wire core__abc_22172_new_n4175_; 
wire core__abc_22172_new_n4176_; 
wire core__abc_22172_new_n4177_; 
wire core__abc_22172_new_n4178_; 
wire core__abc_22172_new_n4179_; 
wire core__abc_22172_new_n4180_; 
wire core__abc_22172_new_n4181_; 
wire core__abc_22172_new_n4182_; 
wire core__abc_22172_new_n4183_; 
wire core__abc_22172_new_n4184_; 
wire core__abc_22172_new_n4186_; 
wire core__abc_22172_new_n4187_; 
wire core__abc_22172_new_n4188_; 
wire core__abc_22172_new_n4189_; 
wire core__abc_22172_new_n4190_; 
wire core__abc_22172_new_n4191_; 
wire core__abc_22172_new_n4192_; 
wire core__abc_22172_new_n4193_; 
wire core__abc_22172_new_n4194_; 
wire core__abc_22172_new_n4195_; 
wire core__abc_22172_new_n4196_; 
wire core__abc_22172_new_n4197_; 
wire core__abc_22172_new_n4198_; 
wire core__abc_22172_new_n4199_; 
wire core__abc_22172_new_n4200_; 
wire core__abc_22172_new_n4201_; 
wire core__abc_22172_new_n4202_; 
wire core__abc_22172_new_n4203_; 
wire core__abc_22172_new_n4204_; 
wire core__abc_22172_new_n4205_; 
wire core__abc_22172_new_n4206_; 
wire core__abc_22172_new_n4207_; 
wire core__abc_22172_new_n4208_; 
wire core__abc_22172_new_n4209_; 
wire core__abc_22172_new_n4210_; 
wire core__abc_22172_new_n4211_; 
wire core__abc_22172_new_n4212_; 
wire core__abc_22172_new_n4213_; 
wire core__abc_22172_new_n4214_; 
wire core__abc_22172_new_n4215_; 
wire core__abc_22172_new_n4216_; 
wire core__abc_22172_new_n4217_; 
wire core__abc_22172_new_n4218_; 
wire core__abc_22172_new_n4219_; 
wire core__abc_22172_new_n4220_; 
wire core__abc_22172_new_n4221_; 
wire core__abc_22172_new_n4222_; 
wire core__abc_22172_new_n4223_; 
wire core__abc_22172_new_n4224_; 
wire core__abc_22172_new_n4225_; 
wire core__abc_22172_new_n4226_; 
wire core__abc_22172_new_n4227_; 
wire core__abc_22172_new_n4228_; 
wire core__abc_22172_new_n4229_; 
wire core__abc_22172_new_n4230_; 
wire core__abc_22172_new_n4231_; 
wire core__abc_22172_new_n4232_; 
wire core__abc_22172_new_n4233_; 
wire core__abc_22172_new_n4234_; 
wire core__abc_22172_new_n4235_; 
wire core__abc_22172_new_n4236_; 
wire core__abc_22172_new_n4237_; 
wire core__abc_22172_new_n4238_; 
wire core__abc_22172_new_n4239_; 
wire core__abc_22172_new_n4240_; 
wire core__abc_22172_new_n4241_; 
wire core__abc_22172_new_n4242_; 
wire core__abc_22172_new_n4243_; 
wire core__abc_22172_new_n4244_; 
wire core__abc_22172_new_n4245_; 
wire core__abc_22172_new_n4246_; 
wire core__abc_22172_new_n4247_; 
wire core__abc_22172_new_n4248_; 
wire core__abc_22172_new_n4249_; 
wire core__abc_22172_new_n4250_; 
wire core__abc_22172_new_n4251_; 
wire core__abc_22172_new_n4252_; 
wire core__abc_22172_new_n4253_; 
wire core__abc_22172_new_n4254_; 
wire core__abc_22172_new_n4255_; 
wire core__abc_22172_new_n4256_; 
wire core__abc_22172_new_n4257_; 
wire core__abc_22172_new_n4258_; 
wire core__abc_22172_new_n4259_; 
wire core__abc_22172_new_n4260_; 
wire core__abc_22172_new_n4261_; 
wire core__abc_22172_new_n4262_; 
wire core__abc_22172_new_n4263_; 
wire core__abc_22172_new_n4264_; 
wire core__abc_22172_new_n4265_; 
wire core__abc_22172_new_n4266_; 
wire core__abc_22172_new_n4267_; 
wire core__abc_22172_new_n4268_; 
wire core__abc_22172_new_n4270_; 
wire core__abc_22172_new_n4271_; 
wire core__abc_22172_new_n4272_; 
wire core__abc_22172_new_n4273_; 
wire core__abc_22172_new_n4274_; 
wire core__abc_22172_new_n4275_; 
wire core__abc_22172_new_n4276_; 
wire core__abc_22172_new_n4277_; 
wire core__abc_22172_new_n4278_; 
wire core__abc_22172_new_n4279_; 
wire core__abc_22172_new_n4280_; 
wire core__abc_22172_new_n4281_; 
wire core__abc_22172_new_n4282_; 
wire core__abc_22172_new_n4283_; 
wire core__abc_22172_new_n4284_; 
wire core__abc_22172_new_n4285_; 
wire core__abc_22172_new_n4286_; 
wire core__abc_22172_new_n4287_; 
wire core__abc_22172_new_n4288_; 
wire core__abc_22172_new_n4289_; 
wire core__abc_22172_new_n4290_; 
wire core__abc_22172_new_n4291_; 
wire core__abc_22172_new_n4292_; 
wire core__abc_22172_new_n4293_; 
wire core__abc_22172_new_n4294_; 
wire core__abc_22172_new_n4295_; 
wire core__abc_22172_new_n4296_; 
wire core__abc_22172_new_n4297_; 
wire core__abc_22172_new_n4298_; 
wire core__abc_22172_new_n4299_; 
wire core__abc_22172_new_n4300_; 
wire core__abc_22172_new_n4301_; 
wire core__abc_22172_new_n4302_; 
wire core__abc_22172_new_n4303_; 
wire core__abc_22172_new_n4304_; 
wire core__abc_22172_new_n4305_; 
wire core__abc_22172_new_n4306_; 
wire core__abc_22172_new_n4307_; 
wire core__abc_22172_new_n4308_; 
wire core__abc_22172_new_n4309_; 
wire core__abc_22172_new_n4310_; 
wire core__abc_22172_new_n4311_; 
wire core__abc_22172_new_n4312_; 
wire core__abc_22172_new_n4313_; 
wire core__abc_22172_new_n4314_; 
wire core__abc_22172_new_n4315_; 
wire core__abc_22172_new_n4316_; 
wire core__abc_22172_new_n4317_; 
wire core__abc_22172_new_n4318_; 
wire core__abc_22172_new_n4319_; 
wire core__abc_22172_new_n4320_; 
wire core__abc_22172_new_n4321_; 
wire core__abc_22172_new_n4322_; 
wire core__abc_22172_new_n4323_; 
wire core__abc_22172_new_n4324_; 
wire core__abc_22172_new_n4325_; 
wire core__abc_22172_new_n4326_; 
wire core__abc_22172_new_n4327_; 
wire core__abc_22172_new_n4328_; 
wire core__abc_22172_new_n4329_; 
wire core__abc_22172_new_n4330_; 
wire core__abc_22172_new_n4331_; 
wire core__abc_22172_new_n4332_; 
wire core__abc_22172_new_n4333_; 
wire core__abc_22172_new_n4334_; 
wire core__abc_22172_new_n4335_; 
wire core__abc_22172_new_n4336_; 
wire core__abc_22172_new_n4338_; 
wire core__abc_22172_new_n4339_; 
wire core__abc_22172_new_n4340_; 
wire core__abc_22172_new_n4341_; 
wire core__abc_22172_new_n4342_; 
wire core__abc_22172_new_n4343_; 
wire core__abc_22172_new_n4344_; 
wire core__abc_22172_new_n4345_; 
wire core__abc_22172_new_n4346_; 
wire core__abc_22172_new_n4347_; 
wire core__abc_22172_new_n4348_; 
wire core__abc_22172_new_n4349_; 
wire core__abc_22172_new_n4350_; 
wire core__abc_22172_new_n4351_; 
wire core__abc_22172_new_n4352_; 
wire core__abc_22172_new_n4353_; 
wire core__abc_22172_new_n4354_; 
wire core__abc_22172_new_n4355_; 
wire core__abc_22172_new_n4356_; 
wire core__abc_22172_new_n4357_; 
wire core__abc_22172_new_n4358_; 
wire core__abc_22172_new_n4359_; 
wire core__abc_22172_new_n4360_; 
wire core__abc_22172_new_n4361_; 
wire core__abc_22172_new_n4362_; 
wire core__abc_22172_new_n4363_; 
wire core__abc_22172_new_n4364_; 
wire core__abc_22172_new_n4365_; 
wire core__abc_22172_new_n4366_; 
wire core__abc_22172_new_n4367_; 
wire core__abc_22172_new_n4368_; 
wire core__abc_22172_new_n4369_; 
wire core__abc_22172_new_n4370_; 
wire core__abc_22172_new_n4371_; 
wire core__abc_22172_new_n4372_; 
wire core__abc_22172_new_n4373_; 
wire core__abc_22172_new_n4374_; 
wire core__abc_22172_new_n4375_; 
wire core__abc_22172_new_n4376_; 
wire core__abc_22172_new_n4377_; 
wire core__abc_22172_new_n4378_; 
wire core__abc_22172_new_n4379_; 
wire core__abc_22172_new_n4380_; 
wire core__abc_22172_new_n4381_; 
wire core__abc_22172_new_n4382_; 
wire core__abc_22172_new_n4383_; 
wire core__abc_22172_new_n4384_; 
wire core__abc_22172_new_n4385_; 
wire core__abc_22172_new_n4386_; 
wire core__abc_22172_new_n4387_; 
wire core__abc_22172_new_n4388_; 
wire core__abc_22172_new_n4389_; 
wire core__abc_22172_new_n4390_; 
wire core__abc_22172_new_n4391_; 
wire core__abc_22172_new_n4392_; 
wire core__abc_22172_new_n4393_; 
wire core__abc_22172_new_n4394_; 
wire core__abc_22172_new_n4395_; 
wire core__abc_22172_new_n4396_; 
wire core__abc_22172_new_n4398_; 
wire core__abc_22172_new_n4399_; 
wire core__abc_22172_new_n4400_; 
wire core__abc_22172_new_n4401_; 
wire core__abc_22172_new_n4402_; 
wire core__abc_22172_new_n4403_; 
wire core__abc_22172_new_n4404_; 
wire core__abc_22172_new_n4405_; 
wire core__abc_22172_new_n4406_; 
wire core__abc_22172_new_n4407_; 
wire core__abc_22172_new_n4408_; 
wire core__abc_22172_new_n4409_; 
wire core__abc_22172_new_n4410_; 
wire core__abc_22172_new_n4411_; 
wire core__abc_22172_new_n4412_; 
wire core__abc_22172_new_n4413_; 
wire core__abc_22172_new_n4414_; 
wire core__abc_22172_new_n4415_; 
wire core__abc_22172_new_n4416_; 
wire core__abc_22172_new_n4417_; 
wire core__abc_22172_new_n4418_; 
wire core__abc_22172_new_n4419_; 
wire core__abc_22172_new_n4420_; 
wire core__abc_22172_new_n4421_; 
wire core__abc_22172_new_n4422_; 
wire core__abc_22172_new_n4423_; 
wire core__abc_22172_new_n4424_; 
wire core__abc_22172_new_n4425_; 
wire core__abc_22172_new_n4426_; 
wire core__abc_22172_new_n4427_; 
wire core__abc_22172_new_n4428_; 
wire core__abc_22172_new_n4429_; 
wire core__abc_22172_new_n4430_; 
wire core__abc_22172_new_n4431_; 
wire core__abc_22172_new_n4432_; 
wire core__abc_22172_new_n4433_; 
wire core__abc_22172_new_n4434_; 
wire core__abc_22172_new_n4435_; 
wire core__abc_22172_new_n4436_; 
wire core__abc_22172_new_n4437_; 
wire core__abc_22172_new_n4438_; 
wire core__abc_22172_new_n4439_; 
wire core__abc_22172_new_n4440_; 
wire core__abc_22172_new_n4441_; 
wire core__abc_22172_new_n4442_; 
wire core__abc_22172_new_n4443_; 
wire core__abc_22172_new_n4444_; 
wire core__abc_22172_new_n4445_; 
wire core__abc_22172_new_n4446_; 
wire core__abc_22172_new_n4447_; 
wire core__abc_22172_new_n4448_; 
wire core__abc_22172_new_n4450_; 
wire core__abc_22172_new_n4451_; 
wire core__abc_22172_new_n4452_; 
wire core__abc_22172_new_n4453_; 
wire core__abc_22172_new_n4454_; 
wire core__abc_22172_new_n4455_; 
wire core__abc_22172_new_n4456_; 
wire core__abc_22172_new_n4457_; 
wire core__abc_22172_new_n4458_; 
wire core__abc_22172_new_n4459_; 
wire core__abc_22172_new_n4460_; 
wire core__abc_22172_new_n4461_; 
wire core__abc_22172_new_n4462_; 
wire core__abc_22172_new_n4463_; 
wire core__abc_22172_new_n4464_; 
wire core__abc_22172_new_n4465_; 
wire core__abc_22172_new_n4466_; 
wire core__abc_22172_new_n4467_; 
wire core__abc_22172_new_n4468_; 
wire core__abc_22172_new_n4469_; 
wire core__abc_22172_new_n4470_; 
wire core__abc_22172_new_n4471_; 
wire core__abc_22172_new_n4472_; 
wire core__abc_22172_new_n4473_; 
wire core__abc_22172_new_n4474_; 
wire core__abc_22172_new_n4475_; 
wire core__abc_22172_new_n4476_; 
wire core__abc_22172_new_n4477_; 
wire core__abc_22172_new_n4478_; 
wire core__abc_22172_new_n4479_; 
wire core__abc_22172_new_n4480_; 
wire core__abc_22172_new_n4481_; 
wire core__abc_22172_new_n4482_; 
wire core__abc_22172_new_n4483_; 
wire core__abc_22172_new_n4484_; 
wire core__abc_22172_new_n4485_; 
wire core__abc_22172_new_n4486_; 
wire core__abc_22172_new_n4487_; 
wire core__abc_22172_new_n4488_; 
wire core__abc_22172_new_n4489_; 
wire core__abc_22172_new_n4490_; 
wire core__abc_22172_new_n4491_; 
wire core__abc_22172_new_n4492_; 
wire core__abc_22172_new_n4493_; 
wire core__abc_22172_new_n4494_; 
wire core__abc_22172_new_n4495_; 
wire core__abc_22172_new_n4496_; 
wire core__abc_22172_new_n4497_; 
wire core__abc_22172_new_n4498_; 
wire core__abc_22172_new_n4499_; 
wire core__abc_22172_new_n4500_; 
wire core__abc_22172_new_n4501_; 
wire core__abc_22172_new_n4502_; 
wire core__abc_22172_new_n4503_; 
wire core__abc_22172_new_n4504_; 
wire core__abc_22172_new_n4505_; 
wire core__abc_22172_new_n4506_; 
wire core__abc_22172_new_n4507_; 
wire core__abc_22172_new_n4508_; 
wire core__abc_22172_new_n4509_; 
wire core__abc_22172_new_n4510_; 
wire core__abc_22172_new_n4511_; 
wire core__abc_22172_new_n4512_; 
wire core__abc_22172_new_n4513_; 
wire core__abc_22172_new_n4514_; 
wire core__abc_22172_new_n4515_; 
wire core__abc_22172_new_n4516_; 
wire core__abc_22172_new_n4517_; 
wire core__abc_22172_new_n4518_; 
wire core__abc_22172_new_n4519_; 
wire core__abc_22172_new_n4520_; 
wire core__abc_22172_new_n4522_; 
wire core__abc_22172_new_n4523_; 
wire core__abc_22172_new_n4524_; 
wire core__abc_22172_new_n4525_; 
wire core__abc_22172_new_n4526_; 
wire core__abc_22172_new_n4527_; 
wire core__abc_22172_new_n4528_; 
wire core__abc_22172_new_n4529_; 
wire core__abc_22172_new_n4530_; 
wire core__abc_22172_new_n4531_; 
wire core__abc_22172_new_n4532_; 
wire core__abc_22172_new_n4533_; 
wire core__abc_22172_new_n4534_; 
wire core__abc_22172_new_n4535_; 
wire core__abc_22172_new_n4536_; 
wire core__abc_22172_new_n4537_; 
wire core__abc_22172_new_n4538_; 
wire core__abc_22172_new_n4539_; 
wire core__abc_22172_new_n4540_; 
wire core__abc_22172_new_n4541_; 
wire core__abc_22172_new_n4542_; 
wire core__abc_22172_new_n4543_; 
wire core__abc_22172_new_n4544_; 
wire core__abc_22172_new_n4545_; 
wire core__abc_22172_new_n4546_; 
wire core__abc_22172_new_n4547_; 
wire core__abc_22172_new_n4548_; 
wire core__abc_22172_new_n4549_; 
wire core__abc_22172_new_n4550_; 
wire core__abc_22172_new_n4551_; 
wire core__abc_22172_new_n4552_; 
wire core__abc_22172_new_n4553_; 
wire core__abc_22172_new_n4554_; 
wire core__abc_22172_new_n4555_; 
wire core__abc_22172_new_n4556_; 
wire core__abc_22172_new_n4557_; 
wire core__abc_22172_new_n4558_; 
wire core__abc_22172_new_n4559_; 
wire core__abc_22172_new_n4560_; 
wire core__abc_22172_new_n4561_; 
wire core__abc_22172_new_n4562_; 
wire core__abc_22172_new_n4563_; 
wire core__abc_22172_new_n4564_; 
wire core__abc_22172_new_n4566_; 
wire core__abc_22172_new_n4567_; 
wire core__abc_22172_new_n4568_; 
wire core__abc_22172_new_n4569_; 
wire core__abc_22172_new_n4570_; 
wire core__abc_22172_new_n4571_; 
wire core__abc_22172_new_n4572_; 
wire core__abc_22172_new_n4573_; 
wire core__abc_22172_new_n4574_; 
wire core__abc_22172_new_n4575_; 
wire core__abc_22172_new_n4576_; 
wire core__abc_22172_new_n4577_; 
wire core__abc_22172_new_n4578_; 
wire core__abc_22172_new_n4579_; 
wire core__abc_22172_new_n4580_; 
wire core__abc_22172_new_n4581_; 
wire core__abc_22172_new_n4582_; 
wire core__abc_22172_new_n4583_; 
wire core__abc_22172_new_n4584_; 
wire core__abc_22172_new_n4585_; 
wire core__abc_22172_new_n4586_; 
wire core__abc_22172_new_n4587_; 
wire core__abc_22172_new_n4588_; 
wire core__abc_22172_new_n4589_; 
wire core__abc_22172_new_n4590_; 
wire core__abc_22172_new_n4591_; 
wire core__abc_22172_new_n4592_; 
wire core__abc_22172_new_n4593_; 
wire core__abc_22172_new_n4594_; 
wire core__abc_22172_new_n4595_; 
wire core__abc_22172_new_n4596_; 
wire core__abc_22172_new_n4597_; 
wire core__abc_22172_new_n4598_; 
wire core__abc_22172_new_n4599_; 
wire core__abc_22172_new_n4600_; 
wire core__abc_22172_new_n4601_; 
wire core__abc_22172_new_n4602_; 
wire core__abc_22172_new_n4603_; 
wire core__abc_22172_new_n4604_; 
wire core__abc_22172_new_n4605_; 
wire core__abc_22172_new_n4606_; 
wire core__abc_22172_new_n4607_; 
wire core__abc_22172_new_n4608_; 
wire core__abc_22172_new_n4609_; 
wire core__abc_22172_new_n4610_; 
wire core__abc_22172_new_n4611_; 
wire core__abc_22172_new_n4612_; 
wire core__abc_22172_new_n4613_; 
wire core__abc_22172_new_n4614_; 
wire core__abc_22172_new_n4615_; 
wire core__abc_22172_new_n4616_; 
wire core__abc_22172_new_n4617_; 
wire core__abc_22172_new_n4618_; 
wire core__abc_22172_new_n4619_; 
wire core__abc_22172_new_n4621_; 
wire core__abc_22172_new_n4622_; 
wire core__abc_22172_new_n4623_; 
wire core__abc_22172_new_n4624_; 
wire core__abc_22172_new_n4625_; 
wire core__abc_22172_new_n4626_; 
wire core__abc_22172_new_n4627_; 
wire core__abc_22172_new_n4628_; 
wire core__abc_22172_new_n4629_; 
wire core__abc_22172_new_n4630_; 
wire core__abc_22172_new_n4631_; 
wire core__abc_22172_new_n4632_; 
wire core__abc_22172_new_n4633_; 
wire core__abc_22172_new_n4634_; 
wire core__abc_22172_new_n4635_; 
wire core__abc_22172_new_n4636_; 
wire core__abc_22172_new_n4637_; 
wire core__abc_22172_new_n4638_; 
wire core__abc_22172_new_n4639_; 
wire core__abc_22172_new_n4640_; 
wire core__abc_22172_new_n4641_; 
wire core__abc_22172_new_n4642_; 
wire core__abc_22172_new_n4643_; 
wire core__abc_22172_new_n4644_; 
wire core__abc_22172_new_n4645_; 
wire core__abc_22172_new_n4646_; 
wire core__abc_22172_new_n4647_; 
wire core__abc_22172_new_n4648_; 
wire core__abc_22172_new_n4649_; 
wire core__abc_22172_new_n4650_; 
wire core__abc_22172_new_n4651_; 
wire core__abc_22172_new_n4652_; 
wire core__abc_22172_new_n4653_; 
wire core__abc_22172_new_n4654_; 
wire core__abc_22172_new_n4655_; 
wire core__abc_22172_new_n4656_; 
wire core__abc_22172_new_n4657_; 
wire core__abc_22172_new_n4658_; 
wire core__abc_22172_new_n4659_; 
wire core__abc_22172_new_n4660_; 
wire core__abc_22172_new_n4661_; 
wire core__abc_22172_new_n4662_; 
wire core__abc_22172_new_n4664_; 
wire core__abc_22172_new_n4665_; 
wire core__abc_22172_new_n4666_; 
wire core__abc_22172_new_n4667_; 
wire core__abc_22172_new_n4668_; 
wire core__abc_22172_new_n4669_; 
wire core__abc_22172_new_n4670_; 
wire core__abc_22172_new_n4671_; 
wire core__abc_22172_new_n4672_; 
wire core__abc_22172_new_n4673_; 
wire core__abc_22172_new_n4674_; 
wire core__abc_22172_new_n4675_; 
wire core__abc_22172_new_n4676_; 
wire core__abc_22172_new_n4677_; 
wire core__abc_22172_new_n4678_; 
wire core__abc_22172_new_n4679_; 
wire core__abc_22172_new_n4680_; 
wire core__abc_22172_new_n4681_; 
wire core__abc_22172_new_n4682_; 
wire core__abc_22172_new_n4683_; 
wire core__abc_22172_new_n4684_; 
wire core__abc_22172_new_n4685_; 
wire core__abc_22172_new_n4686_; 
wire core__abc_22172_new_n4687_; 
wire core__abc_22172_new_n4688_; 
wire core__abc_22172_new_n4689_; 
wire core__abc_22172_new_n4690_; 
wire core__abc_22172_new_n4691_; 
wire core__abc_22172_new_n4692_; 
wire core__abc_22172_new_n4693_; 
wire core__abc_22172_new_n4694_; 
wire core__abc_22172_new_n4695_; 
wire core__abc_22172_new_n4696_; 
wire core__abc_22172_new_n4697_; 
wire core__abc_22172_new_n4698_; 
wire core__abc_22172_new_n4699_; 
wire core__abc_22172_new_n4700_; 
wire core__abc_22172_new_n4701_; 
wire core__abc_22172_new_n4702_; 
wire core__abc_22172_new_n4703_; 
wire core__abc_22172_new_n4704_; 
wire core__abc_22172_new_n4705_; 
wire core__abc_22172_new_n4706_; 
wire core__abc_22172_new_n4707_; 
wire core__abc_22172_new_n4708_; 
wire core__abc_22172_new_n4709_; 
wire core__abc_22172_new_n4710_; 
wire core__abc_22172_new_n4711_; 
wire core__abc_22172_new_n4712_; 
wire core__abc_22172_new_n4713_; 
wire core__abc_22172_new_n4714_; 
wire core__abc_22172_new_n4715_; 
wire core__abc_22172_new_n4716_; 
wire core__abc_22172_new_n4717_; 
wire core__abc_22172_new_n4718_; 
wire core__abc_22172_new_n4719_; 
wire core__abc_22172_new_n4720_; 
wire core__abc_22172_new_n4721_; 
wire core__abc_22172_new_n4722_; 
wire core__abc_22172_new_n4723_; 
wire core__abc_22172_new_n4724_; 
wire core__abc_22172_new_n4725_; 
wire core__abc_22172_new_n4726_; 
wire core__abc_22172_new_n4727_; 
wire core__abc_22172_new_n4728_; 
wire core__abc_22172_new_n4729_; 
wire core__abc_22172_new_n4730_; 
wire core__abc_22172_new_n4731_; 
wire core__abc_22172_new_n4732_; 
wire core__abc_22172_new_n4734_; 
wire core__abc_22172_new_n4735_; 
wire core__abc_22172_new_n4736_; 
wire core__abc_22172_new_n4737_; 
wire core__abc_22172_new_n4738_; 
wire core__abc_22172_new_n4739_; 
wire core__abc_22172_new_n4740_; 
wire core__abc_22172_new_n4741_; 
wire core__abc_22172_new_n4742_; 
wire core__abc_22172_new_n4743_; 
wire core__abc_22172_new_n4744_; 
wire core__abc_22172_new_n4745_; 
wire core__abc_22172_new_n4746_; 
wire core__abc_22172_new_n4747_; 
wire core__abc_22172_new_n4748_; 
wire core__abc_22172_new_n4749_; 
wire core__abc_22172_new_n4750_; 
wire core__abc_22172_new_n4751_; 
wire core__abc_22172_new_n4752_; 
wire core__abc_22172_new_n4753_; 
wire core__abc_22172_new_n4754_; 
wire core__abc_22172_new_n4755_; 
wire core__abc_22172_new_n4756_; 
wire core__abc_22172_new_n4757_; 
wire core__abc_22172_new_n4758_; 
wire core__abc_22172_new_n4759_; 
wire core__abc_22172_new_n4760_; 
wire core__abc_22172_new_n4761_; 
wire core__abc_22172_new_n4762_; 
wire core__abc_22172_new_n4763_; 
wire core__abc_22172_new_n4764_; 
wire core__abc_22172_new_n4765_; 
wire core__abc_22172_new_n4766_; 
wire core__abc_22172_new_n4767_; 
wire core__abc_22172_new_n4768_; 
wire core__abc_22172_new_n4769_; 
wire core__abc_22172_new_n4770_; 
wire core__abc_22172_new_n4771_; 
wire core__abc_22172_new_n4772_; 
wire core__abc_22172_new_n4773_; 
wire core__abc_22172_new_n4774_; 
wire core__abc_22172_new_n4775_; 
wire core__abc_22172_new_n4777_; 
wire core__abc_22172_new_n4778_; 
wire core__abc_22172_new_n4779_; 
wire core__abc_22172_new_n4780_; 
wire core__abc_22172_new_n4781_; 
wire core__abc_22172_new_n4782_; 
wire core__abc_22172_new_n4783_; 
wire core__abc_22172_new_n4784_; 
wire core__abc_22172_new_n4785_; 
wire core__abc_22172_new_n4786_; 
wire core__abc_22172_new_n4787_; 
wire core__abc_22172_new_n4788_; 
wire core__abc_22172_new_n4789_; 
wire core__abc_22172_new_n4790_; 
wire core__abc_22172_new_n4791_; 
wire core__abc_22172_new_n4792_; 
wire core__abc_22172_new_n4793_; 
wire core__abc_22172_new_n4794_; 
wire core__abc_22172_new_n4795_; 
wire core__abc_22172_new_n4796_; 
wire core__abc_22172_new_n4797_; 
wire core__abc_22172_new_n4798_; 
wire core__abc_22172_new_n4799_; 
wire core__abc_22172_new_n4800_; 
wire core__abc_22172_new_n4801_; 
wire core__abc_22172_new_n4802_; 
wire core__abc_22172_new_n4803_; 
wire core__abc_22172_new_n4804_; 
wire core__abc_22172_new_n4805_; 
wire core__abc_22172_new_n4806_; 
wire core__abc_22172_new_n4807_; 
wire core__abc_22172_new_n4808_; 
wire core__abc_22172_new_n4809_; 
wire core__abc_22172_new_n4810_; 
wire core__abc_22172_new_n4811_; 
wire core__abc_22172_new_n4812_; 
wire core__abc_22172_new_n4813_; 
wire core__abc_22172_new_n4814_; 
wire core__abc_22172_new_n4815_; 
wire core__abc_22172_new_n4816_; 
wire core__abc_22172_new_n4817_; 
wire core__abc_22172_new_n4818_; 
wire core__abc_22172_new_n4819_; 
wire core__abc_22172_new_n4820_; 
wire core__abc_22172_new_n4821_; 
wire core__abc_22172_new_n4822_; 
wire core__abc_22172_new_n4823_; 
wire core__abc_22172_new_n4824_; 
wire core__abc_22172_new_n4825_; 
wire core__abc_22172_new_n4826_; 
wire core__abc_22172_new_n4827_; 
wire core__abc_22172_new_n4828_; 
wire core__abc_22172_new_n4829_; 
wire core__abc_22172_new_n4831_; 
wire core__abc_22172_new_n4832_; 
wire core__abc_22172_new_n4833_; 
wire core__abc_22172_new_n4834_; 
wire core__abc_22172_new_n4835_; 
wire core__abc_22172_new_n4836_; 
wire core__abc_22172_new_n4837_; 
wire core__abc_22172_new_n4838_; 
wire core__abc_22172_new_n4839_; 
wire core__abc_22172_new_n4840_; 
wire core__abc_22172_new_n4841_; 
wire core__abc_22172_new_n4842_; 
wire core__abc_22172_new_n4843_; 
wire core__abc_22172_new_n4844_; 
wire core__abc_22172_new_n4845_; 
wire core__abc_22172_new_n4846_; 
wire core__abc_22172_new_n4847_; 
wire core__abc_22172_new_n4848_; 
wire core__abc_22172_new_n4849_; 
wire core__abc_22172_new_n4850_; 
wire core__abc_22172_new_n4851_; 
wire core__abc_22172_new_n4852_; 
wire core__abc_22172_new_n4853_; 
wire core__abc_22172_new_n4854_; 
wire core__abc_22172_new_n4855_; 
wire core__abc_22172_new_n4856_; 
wire core__abc_22172_new_n4857_; 
wire core__abc_22172_new_n4858_; 
wire core__abc_22172_new_n4859_; 
wire core__abc_22172_new_n4860_; 
wire core__abc_22172_new_n4861_; 
wire core__abc_22172_new_n4862_; 
wire core__abc_22172_new_n4863_; 
wire core__abc_22172_new_n4864_; 
wire core__abc_22172_new_n4865_; 
wire core__abc_22172_new_n4866_; 
wire core__abc_22172_new_n4867_; 
wire core__abc_22172_new_n4868_; 
wire core__abc_22172_new_n4869_; 
wire core__abc_22172_new_n4870_; 
wire core__abc_22172_new_n4871_; 
wire core__abc_22172_new_n4872_; 
wire core__abc_22172_new_n4874_; 
wire core__abc_22172_new_n4875_; 
wire core__abc_22172_new_n4876_; 
wire core__abc_22172_new_n4877_; 
wire core__abc_22172_new_n4878_; 
wire core__abc_22172_new_n4879_; 
wire core__abc_22172_new_n4880_; 
wire core__abc_22172_new_n4881_; 
wire core__abc_22172_new_n4882_; 
wire core__abc_22172_new_n4883_; 
wire core__abc_22172_new_n4884_; 
wire core__abc_22172_new_n4885_; 
wire core__abc_22172_new_n4886_; 
wire core__abc_22172_new_n4887_; 
wire core__abc_22172_new_n4888_; 
wire core__abc_22172_new_n4889_; 
wire core__abc_22172_new_n4890_; 
wire core__abc_22172_new_n4891_; 
wire core__abc_22172_new_n4892_; 
wire core__abc_22172_new_n4893_; 
wire core__abc_22172_new_n4894_; 
wire core__abc_22172_new_n4895_; 
wire core__abc_22172_new_n4896_; 
wire core__abc_22172_new_n4897_; 
wire core__abc_22172_new_n4898_; 
wire core__abc_22172_new_n4899_; 
wire core__abc_22172_new_n4900_; 
wire core__abc_22172_new_n4901_; 
wire core__abc_22172_new_n4902_; 
wire core__abc_22172_new_n4903_; 
wire core__abc_22172_new_n4904_; 
wire core__abc_22172_new_n4905_; 
wire core__abc_22172_new_n4906_; 
wire core__abc_22172_new_n4907_; 
wire core__abc_22172_new_n4908_; 
wire core__abc_22172_new_n4909_; 
wire core__abc_22172_new_n4910_; 
wire core__abc_22172_new_n4911_; 
wire core__abc_22172_new_n4912_; 
wire core__abc_22172_new_n4913_; 
wire core__abc_22172_new_n4914_; 
wire core__abc_22172_new_n4915_; 
wire core__abc_22172_new_n4916_; 
wire core__abc_22172_new_n4917_; 
wire core__abc_22172_new_n4918_; 
wire core__abc_22172_new_n4919_; 
wire core__abc_22172_new_n4920_; 
wire core__abc_22172_new_n4921_; 
wire core__abc_22172_new_n4922_; 
wire core__abc_22172_new_n4923_; 
wire core__abc_22172_new_n4924_; 
wire core__abc_22172_new_n4925_; 
wire core__abc_22172_new_n4926_; 
wire core__abc_22172_new_n4927_; 
wire core__abc_22172_new_n4928_; 
wire core__abc_22172_new_n4929_; 
wire core__abc_22172_new_n4930_; 
wire core__abc_22172_new_n4931_; 
wire core__abc_22172_new_n4932_; 
wire core__abc_22172_new_n4933_; 
wire core__abc_22172_new_n4934_; 
wire core__abc_22172_new_n4935_; 
wire core__abc_22172_new_n4936_; 
wire core__abc_22172_new_n4937_; 
wire core__abc_22172_new_n4939_; 
wire core__abc_22172_new_n4940_; 
wire core__abc_22172_new_n4941_; 
wire core__abc_22172_new_n4942_; 
wire core__abc_22172_new_n4943_; 
wire core__abc_22172_new_n4944_; 
wire core__abc_22172_new_n4945_; 
wire core__abc_22172_new_n4946_; 
wire core__abc_22172_new_n4947_; 
wire core__abc_22172_new_n4948_; 
wire core__abc_22172_new_n4949_; 
wire core__abc_22172_new_n4950_; 
wire core__abc_22172_new_n4951_; 
wire core__abc_22172_new_n4952_; 
wire core__abc_22172_new_n4953_; 
wire core__abc_22172_new_n4954_; 
wire core__abc_22172_new_n4955_; 
wire core__abc_22172_new_n4956_; 
wire core__abc_22172_new_n4957_; 
wire core__abc_22172_new_n4958_; 
wire core__abc_22172_new_n4959_; 
wire core__abc_22172_new_n4960_; 
wire core__abc_22172_new_n4961_; 
wire core__abc_22172_new_n4962_; 
wire core__abc_22172_new_n4963_; 
wire core__abc_22172_new_n4964_; 
wire core__abc_22172_new_n4965_; 
wire core__abc_22172_new_n4966_; 
wire core__abc_22172_new_n4967_; 
wire core__abc_22172_new_n4968_; 
wire core__abc_22172_new_n4969_; 
wire core__abc_22172_new_n4970_; 
wire core__abc_22172_new_n4971_; 
wire core__abc_22172_new_n4972_; 
wire core__abc_22172_new_n4973_; 
wire core__abc_22172_new_n4974_; 
wire core__abc_22172_new_n4975_; 
wire core__abc_22172_new_n4976_; 
wire core__abc_22172_new_n4977_; 
wire core__abc_22172_new_n4978_; 
wire core__abc_22172_new_n4979_; 
wire core__abc_22172_new_n4980_; 
wire core__abc_22172_new_n4981_; 
wire core__abc_22172_new_n4982_; 
wire core__abc_22172_new_n4983_; 
wire core__abc_22172_new_n4985_; 
wire core__abc_22172_new_n4986_; 
wire core__abc_22172_new_n4987_; 
wire core__abc_22172_new_n4988_; 
wire core__abc_22172_new_n4989_; 
wire core__abc_22172_new_n4990_; 
wire core__abc_22172_new_n4991_; 
wire core__abc_22172_new_n4992_; 
wire core__abc_22172_new_n4993_; 
wire core__abc_22172_new_n4994_; 
wire core__abc_22172_new_n4995_; 
wire core__abc_22172_new_n4996_; 
wire core__abc_22172_new_n4997_; 
wire core__abc_22172_new_n4998_; 
wire core__abc_22172_new_n4999_; 
wire core__abc_22172_new_n5000_; 
wire core__abc_22172_new_n5001_; 
wire core__abc_22172_new_n5002_; 
wire core__abc_22172_new_n5003_; 
wire core__abc_22172_new_n5004_; 
wire core__abc_22172_new_n5005_; 
wire core__abc_22172_new_n5006_; 
wire core__abc_22172_new_n5007_; 
wire core__abc_22172_new_n5008_; 
wire core__abc_22172_new_n5009_; 
wire core__abc_22172_new_n5010_; 
wire core__abc_22172_new_n5011_; 
wire core__abc_22172_new_n5012_; 
wire core__abc_22172_new_n5013_; 
wire core__abc_22172_new_n5014_; 
wire core__abc_22172_new_n5015_; 
wire core__abc_22172_new_n5016_; 
wire core__abc_22172_new_n5017_; 
wire core__abc_22172_new_n5018_; 
wire core__abc_22172_new_n5019_; 
wire core__abc_22172_new_n5020_; 
wire core__abc_22172_new_n5021_; 
wire core__abc_22172_new_n5022_; 
wire core__abc_22172_new_n5023_; 
wire core__abc_22172_new_n5024_; 
wire core__abc_22172_new_n5025_; 
wire core__abc_22172_new_n5026_; 
wire core__abc_22172_new_n5027_; 
wire core__abc_22172_new_n5028_; 
wire core__abc_22172_new_n5029_; 
wire core__abc_22172_new_n5030_; 
wire core__abc_22172_new_n5031_; 
wire core__abc_22172_new_n5032_; 
wire core__abc_22172_new_n5033_; 
wire core__abc_22172_new_n5034_; 
wire core__abc_22172_new_n5035_; 
wire core__abc_22172_new_n5036_; 
wire core__abc_22172_new_n5037_; 
wire core__abc_22172_new_n5039_; 
wire core__abc_22172_new_n5040_; 
wire core__abc_22172_new_n5041_; 
wire core__abc_22172_new_n5042_; 
wire core__abc_22172_new_n5043_; 
wire core__abc_22172_new_n5044_; 
wire core__abc_22172_new_n5045_; 
wire core__abc_22172_new_n5046_; 
wire core__abc_22172_new_n5047_; 
wire core__abc_22172_new_n5048_; 
wire core__abc_22172_new_n5049_; 
wire core__abc_22172_new_n5050_; 
wire core__abc_22172_new_n5051_; 
wire core__abc_22172_new_n5052_; 
wire core__abc_22172_new_n5053_; 
wire core__abc_22172_new_n5054_; 
wire core__abc_22172_new_n5055_; 
wire core__abc_22172_new_n5056_; 
wire core__abc_22172_new_n5057_; 
wire core__abc_22172_new_n5058_; 
wire core__abc_22172_new_n5059_; 
wire core__abc_22172_new_n5060_; 
wire core__abc_22172_new_n5061_; 
wire core__abc_22172_new_n5062_; 
wire core__abc_22172_new_n5063_; 
wire core__abc_22172_new_n5064_; 
wire core__abc_22172_new_n5065_; 
wire core__abc_22172_new_n5066_; 
wire core__abc_22172_new_n5067_; 
wire core__abc_22172_new_n5068_; 
wire core__abc_22172_new_n5069_; 
wire core__abc_22172_new_n5070_; 
wire core__abc_22172_new_n5071_; 
wire core__abc_22172_new_n5072_; 
wire core__abc_22172_new_n5073_; 
wire core__abc_22172_new_n5074_; 
wire core__abc_22172_new_n5075_; 
wire core__abc_22172_new_n5076_; 
wire core__abc_22172_new_n5077_; 
wire core__abc_22172_new_n5078_; 
wire core__abc_22172_new_n5079_; 
wire core__abc_22172_new_n5080_; 
wire core__abc_22172_new_n5081_; 
wire core__abc_22172_new_n5082_; 
wire core__abc_22172_new_n5083_; 
wire core__abc_22172_new_n5084_; 
wire core__abc_22172_new_n5086_; 
wire core__abc_22172_new_n5087_; 
wire core__abc_22172_new_n5088_; 
wire core__abc_22172_new_n5089_; 
wire core__abc_22172_new_n5090_; 
wire core__abc_22172_new_n5091_; 
wire core__abc_22172_new_n5092_; 
wire core__abc_22172_new_n5093_; 
wire core__abc_22172_new_n5094_; 
wire core__abc_22172_new_n5095_; 
wire core__abc_22172_new_n5096_; 
wire core__abc_22172_new_n5097_; 
wire core__abc_22172_new_n5098_; 
wire core__abc_22172_new_n5099_; 
wire core__abc_22172_new_n5100_; 
wire core__abc_22172_new_n5101_; 
wire core__abc_22172_new_n5102_; 
wire core__abc_22172_new_n5103_; 
wire core__abc_22172_new_n5104_; 
wire core__abc_22172_new_n5105_; 
wire core__abc_22172_new_n5106_; 
wire core__abc_22172_new_n5107_; 
wire core__abc_22172_new_n5108_; 
wire core__abc_22172_new_n5109_; 
wire core__abc_22172_new_n5110_; 
wire core__abc_22172_new_n5111_; 
wire core__abc_22172_new_n5112_; 
wire core__abc_22172_new_n5113_; 
wire core__abc_22172_new_n5114_; 
wire core__abc_22172_new_n5115_; 
wire core__abc_22172_new_n5116_; 
wire core__abc_22172_new_n5117_; 
wire core__abc_22172_new_n5118_; 
wire core__abc_22172_new_n5119_; 
wire core__abc_22172_new_n5120_; 
wire core__abc_22172_new_n5121_; 
wire core__abc_22172_new_n5122_; 
wire core__abc_22172_new_n5123_; 
wire core__abc_22172_new_n5124_; 
wire core__abc_22172_new_n5125_; 
wire core__abc_22172_new_n5126_; 
wire core__abc_22172_new_n5127_; 
wire core__abc_22172_new_n5128_; 
wire core__abc_22172_new_n5129_; 
wire core__abc_22172_new_n5130_; 
wire core__abc_22172_new_n5131_; 
wire core__abc_22172_new_n5132_; 
wire core__abc_22172_new_n5133_; 
wire core__abc_22172_new_n5134_; 
wire core__abc_22172_new_n5135_; 
wire core__abc_22172_new_n5136_; 
wire core__abc_22172_new_n5137_; 
wire core__abc_22172_new_n5138_; 
wire core__abc_22172_new_n5139_; 
wire core__abc_22172_new_n5140_; 
wire core__abc_22172_new_n5141_; 
wire core__abc_22172_new_n5142_; 
wire core__abc_22172_new_n5143_; 
wire core__abc_22172_new_n5144_; 
wire core__abc_22172_new_n5145_; 
wire core__abc_22172_new_n5146_; 
wire core__abc_22172_new_n5147_; 
wire core__abc_22172_new_n5148_; 
wire core__abc_22172_new_n5149_; 
wire core__abc_22172_new_n5150_; 
wire core__abc_22172_new_n5151_; 
wire core__abc_22172_new_n5152_; 
wire core__abc_22172_new_n5153_; 
wire core__abc_22172_new_n5154_; 
wire core__abc_22172_new_n5155_; 
wire core__abc_22172_new_n5156_; 
wire core__abc_22172_new_n5158_; 
wire core__abc_22172_new_n5159_; 
wire core__abc_22172_new_n5160_; 
wire core__abc_22172_new_n5161_; 
wire core__abc_22172_new_n5162_; 
wire core__abc_22172_new_n5163_; 
wire core__abc_22172_new_n5164_; 
wire core__abc_22172_new_n5165_; 
wire core__abc_22172_new_n5166_; 
wire core__abc_22172_new_n5167_; 
wire core__abc_22172_new_n5168_; 
wire core__abc_22172_new_n5169_; 
wire core__abc_22172_new_n5170_; 
wire core__abc_22172_new_n5171_; 
wire core__abc_22172_new_n5172_; 
wire core__abc_22172_new_n5173_; 
wire core__abc_22172_new_n5174_; 
wire core__abc_22172_new_n5175_; 
wire core__abc_22172_new_n5176_; 
wire core__abc_22172_new_n5177_; 
wire core__abc_22172_new_n5178_; 
wire core__abc_22172_new_n5179_; 
wire core__abc_22172_new_n5180_; 
wire core__abc_22172_new_n5181_; 
wire core__abc_22172_new_n5182_; 
wire core__abc_22172_new_n5183_; 
wire core__abc_22172_new_n5184_; 
wire core__abc_22172_new_n5185_; 
wire core__abc_22172_new_n5186_; 
wire core__abc_22172_new_n5187_; 
wire core__abc_22172_new_n5188_; 
wire core__abc_22172_new_n5189_; 
wire core__abc_22172_new_n5190_; 
wire core__abc_22172_new_n5191_; 
wire core__abc_22172_new_n5192_; 
wire core__abc_22172_new_n5193_; 
wire core__abc_22172_new_n5194_; 
wire core__abc_22172_new_n5195_; 
wire core__abc_22172_new_n5196_; 
wire core__abc_22172_new_n5197_; 
wire core__abc_22172_new_n5198_; 
wire core__abc_22172_new_n5200_; 
wire core__abc_22172_new_n5201_; 
wire core__abc_22172_new_n5202_; 
wire core__abc_22172_new_n5203_; 
wire core__abc_22172_new_n5204_; 
wire core__abc_22172_new_n5205_; 
wire core__abc_22172_new_n5206_; 
wire core__abc_22172_new_n5207_; 
wire core__abc_22172_new_n5208_; 
wire core__abc_22172_new_n5209_; 
wire core__abc_22172_new_n5210_; 
wire core__abc_22172_new_n5211_; 
wire core__abc_22172_new_n5212_; 
wire core__abc_22172_new_n5213_; 
wire core__abc_22172_new_n5214_; 
wire core__abc_22172_new_n5215_; 
wire core__abc_22172_new_n5216_; 
wire core__abc_22172_new_n5217_; 
wire core__abc_22172_new_n5218_; 
wire core__abc_22172_new_n5219_; 
wire core__abc_22172_new_n5220_; 
wire core__abc_22172_new_n5221_; 
wire core__abc_22172_new_n5222_; 
wire core__abc_22172_new_n5223_; 
wire core__abc_22172_new_n5224_; 
wire core__abc_22172_new_n5225_; 
wire core__abc_22172_new_n5226_; 
wire core__abc_22172_new_n5227_; 
wire core__abc_22172_new_n5228_; 
wire core__abc_22172_new_n5229_; 
wire core__abc_22172_new_n5230_; 
wire core__abc_22172_new_n5231_; 
wire core__abc_22172_new_n5232_; 
wire core__abc_22172_new_n5233_; 
wire core__abc_22172_new_n5234_; 
wire core__abc_22172_new_n5235_; 
wire core__abc_22172_new_n5236_; 
wire core__abc_22172_new_n5237_; 
wire core__abc_22172_new_n5238_; 
wire core__abc_22172_new_n5239_; 
wire core__abc_22172_new_n5240_; 
wire core__abc_22172_new_n5241_; 
wire core__abc_22172_new_n5242_; 
wire core__abc_22172_new_n5243_; 
wire core__abc_22172_new_n5244_; 
wire core__abc_22172_new_n5245_; 
wire core__abc_22172_new_n5247_; 
wire core__abc_22172_new_n5248_; 
wire core__abc_22172_new_n5249_; 
wire core__abc_22172_new_n5250_; 
wire core__abc_22172_new_n5251_; 
wire core__abc_22172_new_n5252_; 
wire core__abc_22172_new_n5253_; 
wire core__abc_22172_new_n5254_; 
wire core__abc_22172_new_n5255_; 
wire core__abc_22172_new_n5256_; 
wire core__abc_22172_new_n5257_; 
wire core__abc_22172_new_n5258_; 
wire core__abc_22172_new_n5259_; 
wire core__abc_22172_new_n5260_; 
wire core__abc_22172_new_n5261_; 
wire core__abc_22172_new_n5262_; 
wire core__abc_22172_new_n5263_; 
wire core__abc_22172_new_n5264_; 
wire core__abc_22172_new_n5265_; 
wire core__abc_22172_new_n5266_; 
wire core__abc_22172_new_n5267_; 
wire core__abc_22172_new_n5268_; 
wire core__abc_22172_new_n5269_; 
wire core__abc_22172_new_n5270_; 
wire core__abc_22172_new_n5271_; 
wire core__abc_22172_new_n5272_; 
wire core__abc_22172_new_n5273_; 
wire core__abc_22172_new_n5274_; 
wire core__abc_22172_new_n5275_; 
wire core__abc_22172_new_n5276_; 
wire core__abc_22172_new_n5277_; 
wire core__abc_22172_new_n5278_; 
wire core__abc_22172_new_n5279_; 
wire core__abc_22172_new_n5280_; 
wire core__abc_22172_new_n5281_; 
wire core__abc_22172_new_n5282_; 
wire core__abc_22172_new_n5283_; 
wire core__abc_22172_new_n5284_; 
wire core__abc_22172_new_n5285_; 
wire core__abc_22172_new_n5286_; 
wire core__abc_22172_new_n5287_; 
wire core__abc_22172_new_n5288_; 
wire core__abc_22172_new_n5289_; 
wire core__abc_22172_new_n5290_; 
wire core__abc_22172_new_n5292_; 
wire core__abc_22172_new_n5293_; 
wire core__abc_22172_new_n5294_; 
wire core__abc_22172_new_n5295_; 
wire core__abc_22172_new_n5296_; 
wire core__abc_22172_new_n5297_; 
wire core__abc_22172_new_n5298_; 
wire core__abc_22172_new_n5299_; 
wire core__abc_22172_new_n5300_; 
wire core__abc_22172_new_n5301_; 
wire core__abc_22172_new_n5302_; 
wire core__abc_22172_new_n5303_; 
wire core__abc_22172_new_n5304_; 
wire core__abc_22172_new_n5305_; 
wire core__abc_22172_new_n5306_; 
wire core__abc_22172_new_n5307_; 
wire core__abc_22172_new_n5308_; 
wire core__abc_22172_new_n5309_; 
wire core__abc_22172_new_n5310_; 
wire core__abc_22172_new_n5311_; 
wire core__abc_22172_new_n5312_; 
wire core__abc_22172_new_n5313_; 
wire core__abc_22172_new_n5314_; 
wire core__abc_22172_new_n5315_; 
wire core__abc_22172_new_n5316_; 
wire core__abc_22172_new_n5317_; 
wire core__abc_22172_new_n5318_; 
wire core__abc_22172_new_n5319_; 
wire core__abc_22172_new_n5320_; 
wire core__abc_22172_new_n5321_; 
wire core__abc_22172_new_n5322_; 
wire core__abc_22172_new_n5323_; 
wire core__abc_22172_new_n5324_; 
wire core__abc_22172_new_n5325_; 
wire core__abc_22172_new_n5326_; 
wire core__abc_22172_new_n5327_; 
wire core__abc_22172_new_n5328_; 
wire core__abc_22172_new_n5329_; 
wire core__abc_22172_new_n5330_; 
wire core__abc_22172_new_n5331_; 
wire core__abc_22172_new_n5332_; 
wire core__abc_22172_new_n5333_; 
wire core__abc_22172_new_n5334_; 
wire core__abc_22172_new_n5335_; 
wire core__abc_22172_new_n5336_; 
wire core__abc_22172_new_n5337_; 
wire core__abc_22172_new_n5338_; 
wire core__abc_22172_new_n5339_; 
wire core__abc_22172_new_n5340_; 
wire core__abc_22172_new_n5342_; 
wire core__abc_22172_new_n5343_; 
wire core__abc_22172_new_n5344_; 
wire core__abc_22172_new_n5345_; 
wire core__abc_22172_new_n5346_; 
wire core__abc_22172_new_n5347_; 
wire core__abc_22172_new_n5348_; 
wire core__abc_22172_new_n5349_; 
wire core__abc_22172_new_n5350_; 
wire core__abc_22172_new_n5351_; 
wire core__abc_22172_new_n5352_; 
wire core__abc_22172_new_n5353_; 
wire core__abc_22172_new_n5354_; 
wire core__abc_22172_new_n5355_; 
wire core__abc_22172_new_n5356_; 
wire core__abc_22172_new_n5357_; 
wire core__abc_22172_new_n5358_; 
wire core__abc_22172_new_n5359_; 
wire core__abc_22172_new_n5360_; 
wire core__abc_22172_new_n5361_; 
wire core__abc_22172_new_n5362_; 
wire core__abc_22172_new_n5363_; 
wire core__abc_22172_new_n5364_; 
wire core__abc_22172_new_n5365_; 
wire core__abc_22172_new_n5366_; 
wire core__abc_22172_new_n5367_; 
wire core__abc_22172_new_n5368_; 
wire core__abc_22172_new_n5369_; 
wire core__abc_22172_new_n5370_; 
wire core__abc_22172_new_n5371_; 
wire core__abc_22172_new_n5372_; 
wire core__abc_22172_new_n5373_; 
wire core__abc_22172_new_n5374_; 
wire core__abc_22172_new_n5375_; 
wire core__abc_22172_new_n5376_; 
wire core__abc_22172_new_n5377_; 
wire core__abc_22172_new_n5378_; 
wire core__abc_22172_new_n5379_; 
wire core__abc_22172_new_n5380_; 
wire core__abc_22172_new_n5381_; 
wire core__abc_22172_new_n5382_; 
wire core__abc_22172_new_n5383_; 
wire core__abc_22172_new_n5384_; 
wire core__abc_22172_new_n5385_; 
wire core__abc_22172_new_n5386_; 
wire core__abc_22172_new_n5387_; 
wire core__abc_22172_new_n5388_; 
wire core__abc_22172_new_n5390_; 
wire core__abc_22172_new_n5391_; 
wire core__abc_22172_new_n5392_; 
wire core__abc_22172_new_n5393_; 
wire core__abc_22172_new_n5394_; 
wire core__abc_22172_new_n5395_; 
wire core__abc_22172_new_n5396_; 
wire core__abc_22172_new_n5397_; 
wire core__abc_22172_new_n5398_; 
wire core__abc_22172_new_n5399_; 
wire core__abc_22172_new_n5400_; 
wire core__abc_22172_new_n5401_; 
wire core__abc_22172_new_n5402_; 
wire core__abc_22172_new_n5403_; 
wire core__abc_22172_new_n5404_; 
wire core__abc_22172_new_n5405_; 
wire core__abc_22172_new_n5406_; 
wire core__abc_22172_new_n5407_; 
wire core__abc_22172_new_n5408_; 
wire core__abc_22172_new_n5409_; 
wire core__abc_22172_new_n5410_; 
wire core__abc_22172_new_n5411_; 
wire core__abc_22172_new_n5412_; 
wire core__abc_22172_new_n5413_; 
wire core__abc_22172_new_n5414_; 
wire core__abc_22172_new_n5415_; 
wire core__abc_22172_new_n5416_; 
wire core__abc_22172_new_n5417_; 
wire core__abc_22172_new_n5418_; 
wire core__abc_22172_new_n5419_; 
wire core__abc_22172_new_n5420_; 
wire core__abc_22172_new_n5421_; 
wire core__abc_22172_new_n5422_; 
wire core__abc_22172_new_n5423_; 
wire core__abc_22172_new_n5424_; 
wire core__abc_22172_new_n5425_; 
wire core__abc_22172_new_n5426_; 
wire core__abc_22172_new_n5427_; 
wire core__abc_22172_new_n5428_; 
wire core__abc_22172_new_n5429_; 
wire core__abc_22172_new_n5430_; 
wire core__abc_22172_new_n5431_; 
wire core__abc_22172_new_n5432_; 
wire core__abc_22172_new_n5433_; 
wire core__abc_22172_new_n5434_; 
wire core__abc_22172_new_n5435_; 
wire core__abc_22172_new_n5436_; 
wire core__abc_22172_new_n5437_; 
wire core__abc_22172_new_n5439_; 
wire core__abc_22172_new_n5440_; 
wire core__abc_22172_new_n5441_; 
wire core__abc_22172_new_n5442_; 
wire core__abc_22172_new_n5443_; 
wire core__abc_22172_new_n5444_; 
wire core__abc_22172_new_n5445_; 
wire core__abc_22172_new_n5446_; 
wire core__abc_22172_new_n5447_; 
wire core__abc_22172_new_n5448_; 
wire core__abc_22172_new_n5449_; 
wire core__abc_22172_new_n5450_; 
wire core__abc_22172_new_n5451_; 
wire core__abc_22172_new_n5452_; 
wire core__abc_22172_new_n5453_; 
wire core__abc_22172_new_n5454_; 
wire core__abc_22172_new_n5455_; 
wire core__abc_22172_new_n5456_; 
wire core__abc_22172_new_n5457_; 
wire core__abc_22172_new_n5458_; 
wire core__abc_22172_new_n5459_; 
wire core__abc_22172_new_n5460_; 
wire core__abc_22172_new_n5461_; 
wire core__abc_22172_new_n5462_; 
wire core__abc_22172_new_n5463_; 
wire core__abc_22172_new_n5464_; 
wire core__abc_22172_new_n5465_; 
wire core__abc_22172_new_n5466_; 
wire core__abc_22172_new_n5467_; 
wire core__abc_22172_new_n5468_; 
wire core__abc_22172_new_n5469_; 
wire core__abc_22172_new_n5470_; 
wire core__abc_22172_new_n5471_; 
wire core__abc_22172_new_n5472_; 
wire core__abc_22172_new_n5473_; 
wire core__abc_22172_new_n5474_; 
wire core__abc_22172_new_n5475_; 
wire core__abc_22172_new_n5476_; 
wire core__abc_22172_new_n5477_; 
wire core__abc_22172_new_n5478_; 
wire core__abc_22172_new_n5479_; 
wire core__abc_22172_new_n5480_; 
wire core__abc_22172_new_n5482_; 
wire core__abc_22172_new_n5483_; 
wire core__abc_22172_new_n5484_; 
wire core__abc_22172_new_n5485_; 
wire core__abc_22172_new_n5486_; 
wire core__abc_22172_new_n5487_; 
wire core__abc_22172_new_n5488_; 
wire core__abc_22172_new_n5489_; 
wire core__abc_22172_new_n5490_; 
wire core__abc_22172_new_n5491_; 
wire core__abc_22172_new_n5492_; 
wire core__abc_22172_new_n5493_; 
wire core__abc_22172_new_n5494_; 
wire core__abc_22172_new_n5495_; 
wire core__abc_22172_new_n5496_; 
wire core__abc_22172_new_n5497_; 
wire core__abc_22172_new_n5498_; 
wire core__abc_22172_new_n5499_; 
wire core__abc_22172_new_n5500_; 
wire core__abc_22172_new_n5501_; 
wire core__abc_22172_new_n5502_; 
wire core__abc_22172_new_n5503_; 
wire core__abc_22172_new_n5504_; 
wire core__abc_22172_new_n5505_; 
wire core__abc_22172_new_n5506_; 
wire core__abc_22172_new_n5507_; 
wire core__abc_22172_new_n5508_; 
wire core__abc_22172_new_n5509_; 
wire core__abc_22172_new_n5510_; 
wire core__abc_22172_new_n5511_; 
wire core__abc_22172_new_n5512_; 
wire core__abc_22172_new_n5513_; 
wire core__abc_22172_new_n5514_; 
wire core__abc_22172_new_n5515_; 
wire core__abc_22172_new_n5516_; 
wire core__abc_22172_new_n5517_; 
wire core__abc_22172_new_n5518_; 
wire core__abc_22172_new_n5519_; 
wire core__abc_22172_new_n5520_; 
wire core__abc_22172_new_n5521_; 
wire core__abc_22172_new_n5522_; 
wire core__abc_22172_new_n5523_; 
wire core__abc_22172_new_n5524_; 
wire core__abc_22172_new_n5525_; 
wire core__abc_22172_new_n5526_; 
wire core__abc_22172_new_n5527_; 
wire core__abc_22172_new_n5528_; 
wire core__abc_22172_new_n5529_; 
wire core__abc_22172_new_n5530_; 
wire core__abc_22172_new_n5531_; 
wire core__abc_22172_new_n5532_; 
wire core__abc_22172_new_n5533_; 
wire core__abc_22172_new_n5534_; 
wire core__abc_22172_new_n5536_; 
wire core__abc_22172_new_n5537_; 
wire core__abc_22172_new_n5538_; 
wire core__abc_22172_new_n5539_; 
wire core__abc_22172_new_n5540_; 
wire core__abc_22172_new_n5541_; 
wire core__abc_22172_new_n5542_; 
wire core__abc_22172_new_n5543_; 
wire core__abc_22172_new_n5544_; 
wire core__abc_22172_new_n5545_; 
wire core__abc_22172_new_n5546_; 
wire core__abc_22172_new_n5547_; 
wire core__abc_22172_new_n5548_; 
wire core__abc_22172_new_n5549_; 
wire core__abc_22172_new_n5550_; 
wire core__abc_22172_new_n5551_; 
wire core__abc_22172_new_n5552_; 
wire core__abc_22172_new_n5553_; 
wire core__abc_22172_new_n5554_; 
wire core__abc_22172_new_n5555_; 
wire core__abc_22172_new_n5556_; 
wire core__abc_22172_new_n5557_; 
wire core__abc_22172_new_n5558_; 
wire core__abc_22172_new_n5559_; 
wire core__abc_22172_new_n5560_; 
wire core__abc_22172_new_n5561_; 
wire core__abc_22172_new_n5562_; 
wire core__abc_22172_new_n5563_; 
wire core__abc_22172_new_n5564_; 
wire core__abc_22172_new_n5565_; 
wire core__abc_22172_new_n5566_; 
wire core__abc_22172_new_n5567_; 
wire core__abc_22172_new_n5568_; 
wire core__abc_22172_new_n5569_; 
wire core__abc_22172_new_n5570_; 
wire core__abc_22172_new_n5571_; 
wire core__abc_22172_new_n5572_; 
wire core__abc_22172_new_n5573_; 
wire core__abc_22172_new_n5574_; 
wire core__abc_22172_new_n5575_; 
wire core__abc_22172_new_n5576_; 
wire core__abc_22172_new_n5577_; 
wire core__abc_22172_new_n5578_; 
wire core__abc_22172_new_n5579_; 
wire core__abc_22172_new_n5580_; 
wire core__abc_22172_new_n5581_; 
wire core__abc_22172_new_n5583_; 
wire core__abc_22172_new_n5584_; 
wire core__abc_22172_new_n5585_; 
wire core__abc_22172_new_n5586_; 
wire core__abc_22172_new_n5587_; 
wire core__abc_22172_new_n5588_; 
wire core__abc_22172_new_n5589_; 
wire core__abc_22172_new_n5590_; 
wire core__abc_22172_new_n5591_; 
wire core__abc_22172_new_n5592_; 
wire core__abc_22172_new_n5593_; 
wire core__abc_22172_new_n5594_; 
wire core__abc_22172_new_n5595_; 
wire core__abc_22172_new_n5596_; 
wire core__abc_22172_new_n5597_; 
wire core__abc_22172_new_n5598_; 
wire core__abc_22172_new_n5599_; 
wire core__abc_22172_new_n5600_; 
wire core__abc_22172_new_n5601_; 
wire core__abc_22172_new_n5602_; 
wire core__abc_22172_new_n5603_; 
wire core__abc_22172_new_n5604_; 
wire core__abc_22172_new_n5605_; 
wire core__abc_22172_new_n5606_; 
wire core__abc_22172_new_n5607_; 
wire core__abc_22172_new_n5608_; 
wire core__abc_22172_new_n5609_; 
wire core__abc_22172_new_n5610_; 
wire core__abc_22172_new_n5611_; 
wire core__abc_22172_new_n5612_; 
wire core__abc_22172_new_n5613_; 
wire core__abc_22172_new_n5614_; 
wire core__abc_22172_new_n5615_; 
wire core__abc_22172_new_n5616_; 
wire core__abc_22172_new_n5617_; 
wire core__abc_22172_new_n5618_; 
wire core__abc_22172_new_n5619_; 
wire core__abc_22172_new_n5620_; 
wire core__abc_22172_new_n5621_; 
wire core__abc_22172_new_n5622_; 
wire core__abc_22172_new_n5623_; 
wire core__abc_22172_new_n5624_; 
wire core__abc_22172_new_n5625_; 
wire core__abc_22172_new_n5626_; 
wire core__abc_22172_new_n5628_; 
wire core__abc_22172_new_n5629_; 
wire core__abc_22172_new_n5630_; 
wire core__abc_22172_new_n5631_; 
wire core__abc_22172_new_n5632_; 
wire core__abc_22172_new_n5633_; 
wire core__abc_22172_new_n5634_; 
wire core__abc_22172_new_n5635_; 
wire core__abc_22172_new_n5636_; 
wire core__abc_22172_new_n5637_; 
wire core__abc_22172_new_n5638_; 
wire core__abc_22172_new_n5639_; 
wire core__abc_22172_new_n5640_; 
wire core__abc_22172_new_n5641_; 
wire core__abc_22172_new_n5642_; 
wire core__abc_22172_new_n5643_; 
wire core__abc_22172_new_n5644_; 
wire core__abc_22172_new_n5645_; 
wire core__abc_22172_new_n5646_; 
wire core__abc_22172_new_n5647_; 
wire core__abc_22172_new_n5648_; 
wire core__abc_22172_new_n5649_; 
wire core__abc_22172_new_n5650_; 
wire core__abc_22172_new_n5651_; 
wire core__abc_22172_new_n5652_; 
wire core__abc_22172_new_n5653_; 
wire core__abc_22172_new_n5654_; 
wire core__abc_22172_new_n5655_; 
wire core__abc_22172_new_n5656_; 
wire core__abc_22172_new_n5657_; 
wire core__abc_22172_new_n5658_; 
wire core__abc_22172_new_n5659_; 
wire core__abc_22172_new_n5661_; 
wire core__abc_22172_new_n5662_; 
wire core__abc_22172_new_n5663_; 
wire core__abc_22172_new_n5664_; 
wire core__abc_22172_new_n5665_; 
wire core__abc_22172_new_n5666_; 
wire core__abc_22172_new_n5667_; 
wire core__abc_22172_new_n5668_; 
wire core__abc_22172_new_n5669_; 
wire core__abc_22172_new_n5670_; 
wire core__abc_22172_new_n5671_; 
wire core__abc_22172_new_n5672_; 
wire core__abc_22172_new_n5673_; 
wire core__abc_22172_new_n5674_; 
wire core__abc_22172_new_n5675_; 
wire core__abc_22172_new_n5676_; 
wire core__abc_22172_new_n5677_; 
wire core__abc_22172_new_n5678_; 
wire core__abc_22172_new_n5679_; 
wire core__abc_22172_new_n5680_; 
wire core__abc_22172_new_n5681_; 
wire core__abc_22172_new_n5682_; 
wire core__abc_22172_new_n5683_; 
wire core__abc_22172_new_n5684_; 
wire core__abc_22172_new_n5685_; 
wire core__abc_22172_new_n5686_; 
wire core__abc_22172_new_n5687_; 
wire core__abc_22172_new_n5688_; 
wire core__abc_22172_new_n5689_; 
wire core__abc_22172_new_n5690_; 
wire core__abc_22172_new_n5691_; 
wire core__abc_22172_new_n5692_; 
wire core__abc_22172_new_n5693_; 
wire core__abc_22172_new_n5694_; 
wire core__abc_22172_new_n5695_; 
wire core__abc_22172_new_n5696_; 
wire core__abc_22172_new_n5697_; 
wire core__abc_22172_new_n5698_; 
wire core__abc_22172_new_n5699_; 
wire core__abc_22172_new_n5700_; 
wire core__abc_22172_new_n5701_; 
wire core__abc_22172_new_n5702_; 
wire core__abc_22172_new_n5703_; 
wire core__abc_22172_new_n5704_; 
wire core__abc_22172_new_n5705_; 
wire core__abc_22172_new_n5706_; 
wire core__abc_22172_new_n5707_; 
wire core__abc_22172_new_n5708_; 
wire core__abc_22172_new_n5710_; 
wire core__abc_22172_new_n5711_; 
wire core__abc_22172_new_n5712_; 
wire core__abc_22172_new_n5713_; 
wire core__abc_22172_new_n5714_; 
wire core__abc_22172_new_n5715_; 
wire core__abc_22172_new_n5716_; 
wire core__abc_22172_new_n5717_; 
wire core__abc_22172_new_n5718_; 
wire core__abc_22172_new_n5719_; 
wire core__abc_22172_new_n5720_; 
wire core__abc_22172_new_n5721_; 
wire core__abc_22172_new_n5722_; 
wire core__abc_22172_new_n5723_; 
wire core__abc_22172_new_n5724_; 
wire core__abc_22172_new_n5725_; 
wire core__abc_22172_new_n5726_; 
wire core__abc_22172_new_n5727_; 
wire core__abc_22172_new_n5728_; 
wire core__abc_22172_new_n5729_; 
wire core__abc_22172_new_n5730_; 
wire core__abc_22172_new_n5731_; 
wire core__abc_22172_new_n5732_; 
wire core__abc_22172_new_n5733_; 
wire core__abc_22172_new_n5734_; 
wire core__abc_22172_new_n5735_; 
wire core__abc_22172_new_n5736_; 
wire core__abc_22172_new_n5737_; 
wire core__abc_22172_new_n5738_; 
wire core__abc_22172_new_n5739_; 
wire core__abc_22172_new_n5740_; 
wire core__abc_22172_new_n5741_; 
wire core__abc_22172_new_n5743_; 
wire core__abc_22172_new_n5744_; 
wire core__abc_22172_new_n5745_; 
wire core__abc_22172_new_n5746_; 
wire core__abc_22172_new_n5747_; 
wire core__abc_22172_new_n5748_; 
wire core__abc_22172_new_n5749_; 
wire core__abc_22172_new_n5750_; 
wire core__abc_22172_new_n5751_; 
wire core__abc_22172_new_n5752_; 
wire core__abc_22172_new_n5753_; 
wire core__abc_22172_new_n5754_; 
wire core__abc_22172_new_n5755_; 
wire core__abc_22172_new_n5756_; 
wire core__abc_22172_new_n5757_; 
wire core__abc_22172_new_n5758_; 
wire core__abc_22172_new_n5759_; 
wire core__abc_22172_new_n5760_; 
wire core__abc_22172_new_n5761_; 
wire core__abc_22172_new_n5762_; 
wire core__abc_22172_new_n5763_; 
wire core__abc_22172_new_n5764_; 
wire core__abc_22172_new_n5765_; 
wire core__abc_22172_new_n5766_; 
wire core__abc_22172_new_n5767_; 
wire core__abc_22172_new_n5768_; 
wire core__abc_22172_new_n5769_; 
wire core__abc_22172_new_n5770_; 
wire core__abc_22172_new_n5771_; 
wire core__abc_22172_new_n5772_; 
wire core__abc_22172_new_n5773_; 
wire core__abc_22172_new_n5774_; 
wire core__abc_22172_new_n5775_; 
wire core__abc_22172_new_n5776_; 
wire core__abc_22172_new_n5777_; 
wire core__abc_22172_new_n5778_; 
wire core__abc_22172_new_n5779_; 
wire core__abc_22172_new_n5780_; 
wire core__abc_22172_new_n5781_; 
wire core__abc_22172_new_n5782_; 
wire core__abc_22172_new_n5783_; 
wire core__abc_22172_new_n5785_; 
wire core__abc_22172_new_n5786_; 
wire core__abc_22172_new_n5787_; 
wire core__abc_22172_new_n5788_; 
wire core__abc_22172_new_n5789_; 
wire core__abc_22172_new_n5790_; 
wire core__abc_22172_new_n5791_; 
wire core__abc_22172_new_n5792_; 
wire core__abc_22172_new_n5793_; 
wire core__abc_22172_new_n5794_; 
wire core__abc_22172_new_n5795_; 
wire core__abc_22172_new_n5796_; 
wire core__abc_22172_new_n5797_; 
wire core__abc_22172_new_n5798_; 
wire core__abc_22172_new_n5799_; 
wire core__abc_22172_new_n5800_; 
wire core__abc_22172_new_n5801_; 
wire core__abc_22172_new_n5802_; 
wire core__abc_22172_new_n5803_; 
wire core__abc_22172_new_n5804_; 
wire core__abc_22172_new_n5805_; 
wire core__abc_22172_new_n5806_; 
wire core__abc_22172_new_n5807_; 
wire core__abc_22172_new_n5808_; 
wire core__abc_22172_new_n5809_; 
wire core__abc_22172_new_n5810_; 
wire core__abc_22172_new_n5811_; 
wire core__abc_22172_new_n5812_; 
wire core__abc_22172_new_n5813_; 
wire core__abc_22172_new_n5814_; 
wire core__abc_22172_new_n5815_; 
wire core__abc_22172_new_n5816_; 
wire core__abc_22172_new_n5817_; 
wire core__abc_22172_new_n5818_; 
wire core__abc_22172_new_n5819_; 
wire core__abc_22172_new_n5820_; 
wire core__abc_22172_new_n5821_; 
wire core__abc_22172_new_n5823_; 
wire core__abc_22172_new_n5824_; 
wire core__abc_22172_new_n5825_; 
wire core__abc_22172_new_n5826_; 
wire core__abc_22172_new_n5827_; 
wire core__abc_22172_new_n5828_; 
wire core__abc_22172_new_n5829_; 
wire core__abc_22172_new_n5830_; 
wire core__abc_22172_new_n5831_; 
wire core__abc_22172_new_n5832_; 
wire core__abc_22172_new_n5833_; 
wire core__abc_22172_new_n5834_; 
wire core__abc_22172_new_n5835_; 
wire core__abc_22172_new_n5836_; 
wire core__abc_22172_new_n5837_; 
wire core__abc_22172_new_n5838_; 
wire core__abc_22172_new_n5839_; 
wire core__abc_22172_new_n5840_; 
wire core__abc_22172_new_n5841_; 
wire core__abc_22172_new_n5842_; 
wire core__abc_22172_new_n5843_; 
wire core__abc_22172_new_n5844_; 
wire core__abc_22172_new_n5845_; 
wire core__abc_22172_new_n5846_; 
wire core__abc_22172_new_n5847_; 
wire core__abc_22172_new_n5848_; 
wire core__abc_22172_new_n5849_; 
wire core__abc_22172_new_n5850_; 
wire core__abc_22172_new_n5851_; 
wire core__abc_22172_new_n5852_; 
wire core__abc_22172_new_n5853_; 
wire core__abc_22172_new_n5854_; 
wire core__abc_22172_new_n5855_; 
wire core__abc_22172_new_n5856_; 
wire core__abc_22172_new_n5857_; 
wire core__abc_22172_new_n5858_; 
wire core__abc_22172_new_n5859_; 
wire core__abc_22172_new_n5860_; 
wire core__abc_22172_new_n5861_; 
wire core__abc_22172_new_n5862_; 
wire core__abc_22172_new_n5863_; 
wire core__abc_22172_new_n5864_; 
wire core__abc_22172_new_n5865_; 
wire core__abc_22172_new_n5866_; 
wire core__abc_22172_new_n5867_; 
wire core__abc_22172_new_n5868_; 
wire core__abc_22172_new_n5869_; 
wire core__abc_22172_new_n5870_; 
wire core__abc_22172_new_n5871_; 
wire core__abc_22172_new_n5872_; 
wire core__abc_22172_new_n5874_; 
wire core__abc_22172_new_n5875_; 
wire core__abc_22172_new_n5876_; 
wire core__abc_22172_new_n5877_; 
wire core__abc_22172_new_n5878_; 
wire core__abc_22172_new_n5879_; 
wire core__abc_22172_new_n5880_; 
wire core__abc_22172_new_n5881_; 
wire core__abc_22172_new_n5882_; 
wire core__abc_22172_new_n5883_; 
wire core__abc_22172_new_n5884_; 
wire core__abc_22172_new_n5885_; 
wire core__abc_22172_new_n5886_; 
wire core__abc_22172_new_n5887_; 
wire core__abc_22172_new_n5888_; 
wire core__abc_22172_new_n5889_; 
wire core__abc_22172_new_n5890_; 
wire core__abc_22172_new_n5891_; 
wire core__abc_22172_new_n5892_; 
wire core__abc_22172_new_n5893_; 
wire core__abc_22172_new_n5894_; 
wire core__abc_22172_new_n5895_; 
wire core__abc_22172_new_n5896_; 
wire core__abc_22172_new_n5897_; 
wire core__abc_22172_new_n5898_; 
wire core__abc_22172_new_n5899_; 
wire core__abc_22172_new_n5900_; 
wire core__abc_22172_new_n5901_; 
wire core__abc_22172_new_n5902_; 
wire core__abc_22172_new_n5903_; 
wire core__abc_22172_new_n5904_; 
wire core__abc_22172_new_n5905_; 
wire core__abc_22172_new_n5906_; 
wire core__abc_22172_new_n5907_; 
wire core__abc_22172_new_n5908_; 
wire core__abc_22172_new_n5909_; 
wire core__abc_22172_new_n5910_; 
wire core__abc_22172_new_n5911_; 
wire core__abc_22172_new_n5913_; 
wire core__abc_22172_new_n5914_; 
wire core__abc_22172_new_n5915_; 
wire core__abc_22172_new_n5916_; 
wire core__abc_22172_new_n5917_; 
wire core__abc_22172_new_n5918_; 
wire core__abc_22172_new_n5919_; 
wire core__abc_22172_new_n5920_; 
wire core__abc_22172_new_n5921_; 
wire core__abc_22172_new_n5922_; 
wire core__abc_22172_new_n5923_; 
wire core__abc_22172_new_n5924_; 
wire core__abc_22172_new_n5925_; 
wire core__abc_22172_new_n5926_; 
wire core__abc_22172_new_n5927_; 
wire core__abc_22172_new_n5928_; 
wire core__abc_22172_new_n5929_; 
wire core__abc_22172_new_n5930_; 
wire core__abc_22172_new_n5931_; 
wire core__abc_22172_new_n5932_; 
wire core__abc_22172_new_n5933_; 
wire core__abc_22172_new_n5934_; 
wire core__abc_22172_new_n5935_; 
wire core__abc_22172_new_n5936_; 
wire core__abc_22172_new_n5937_; 
wire core__abc_22172_new_n5938_; 
wire core__abc_22172_new_n5939_; 
wire core__abc_22172_new_n5940_; 
wire core__abc_22172_new_n5941_; 
wire core__abc_22172_new_n5942_; 
wire core__abc_22172_new_n5943_; 
wire core__abc_22172_new_n5944_; 
wire core__abc_22172_new_n5945_; 
wire core__abc_22172_new_n5947_; 
wire core__abc_22172_new_n5948_; 
wire core__abc_22172_new_n5949_; 
wire core__abc_22172_new_n5950_; 
wire core__abc_22172_new_n5951_; 
wire core__abc_22172_new_n5952_; 
wire core__abc_22172_new_n5953_; 
wire core__abc_22172_new_n5954_; 
wire core__abc_22172_new_n5955_; 
wire core__abc_22172_new_n5956_; 
wire core__abc_22172_new_n5957_; 
wire core__abc_22172_new_n5958_; 
wire core__abc_22172_new_n5959_; 
wire core__abc_22172_new_n5960_; 
wire core__abc_22172_new_n5961_; 
wire core__abc_22172_new_n5962_; 
wire core__abc_22172_new_n5963_; 
wire core__abc_22172_new_n5964_; 
wire core__abc_22172_new_n5965_; 
wire core__abc_22172_new_n5966_; 
wire core__abc_22172_new_n5967_; 
wire core__abc_22172_new_n5968_; 
wire core__abc_22172_new_n5969_; 
wire core__abc_22172_new_n5970_; 
wire core__abc_22172_new_n5971_; 
wire core__abc_22172_new_n5972_; 
wire core__abc_22172_new_n5973_; 
wire core__abc_22172_new_n5974_; 
wire core__abc_22172_new_n5975_; 
wire core__abc_22172_new_n5976_; 
wire core__abc_22172_new_n5977_; 
wire core__abc_22172_new_n5978_; 
wire core__abc_22172_new_n5979_; 
wire core__abc_22172_new_n5981_; 
wire core__abc_22172_new_n5982_; 
wire core__abc_22172_new_n5983_; 
wire core__abc_22172_new_n5984_; 
wire core__abc_22172_new_n5985_; 
wire core__abc_22172_new_n5986_; 
wire core__abc_22172_new_n5987_; 
wire core__abc_22172_new_n5988_; 
wire core__abc_22172_new_n5989_; 
wire core__abc_22172_new_n5990_; 
wire core__abc_22172_new_n5991_; 
wire core__abc_22172_new_n5992_; 
wire core__abc_22172_new_n5993_; 
wire core__abc_22172_new_n5994_; 
wire core__abc_22172_new_n5995_; 
wire core__abc_22172_new_n5996_; 
wire core__abc_22172_new_n5997_; 
wire core__abc_22172_new_n5998_; 
wire core__abc_22172_new_n5999_; 
wire core__abc_22172_new_n6000_; 
wire core__abc_22172_new_n6001_; 
wire core__abc_22172_new_n6002_; 
wire core__abc_22172_new_n6003_; 
wire core__abc_22172_new_n6004_; 
wire core__abc_22172_new_n6005_; 
wire core__abc_22172_new_n6006_; 
wire core__abc_22172_new_n6007_; 
wire core__abc_22172_new_n6008_; 
wire core__abc_22172_new_n6009_; 
wire core__abc_22172_new_n6010_; 
wire core__abc_22172_new_n6011_; 
wire core__abc_22172_new_n6012_; 
wire core__abc_22172_new_n6013_; 
wire core__abc_22172_new_n6014_; 
wire core__abc_22172_new_n6015_; 
wire core__abc_22172_new_n6016_; 
wire core__abc_22172_new_n6017_; 
wire core__abc_22172_new_n6018_; 
wire core__abc_22172_new_n6019_; 
wire core__abc_22172_new_n6020_; 
wire core__abc_22172_new_n6021_; 
wire core__abc_22172_new_n6022_; 
wire core__abc_22172_new_n6023_; 
wire core__abc_22172_new_n6024_; 
wire core__abc_22172_new_n6025_; 
wire core__abc_22172_new_n6027_; 
wire core__abc_22172_new_n6028_; 
wire core__abc_22172_new_n6029_; 
wire core__abc_22172_new_n6030_; 
wire core__abc_22172_new_n6031_; 
wire core__abc_22172_new_n6032_; 
wire core__abc_22172_new_n6033_; 
wire core__abc_22172_new_n6034_; 
wire core__abc_22172_new_n6035_; 
wire core__abc_22172_new_n6036_; 
wire core__abc_22172_new_n6037_; 
wire core__abc_22172_new_n6038_; 
wire core__abc_22172_new_n6039_; 
wire core__abc_22172_new_n6040_; 
wire core__abc_22172_new_n6041_; 
wire core__abc_22172_new_n6042_; 
wire core__abc_22172_new_n6043_; 
wire core__abc_22172_new_n6044_; 
wire core__abc_22172_new_n6045_; 
wire core__abc_22172_new_n6046_; 
wire core__abc_22172_new_n6047_; 
wire core__abc_22172_new_n6048_; 
wire core__abc_22172_new_n6049_; 
wire core__abc_22172_new_n6050_; 
wire core__abc_22172_new_n6051_; 
wire core__abc_22172_new_n6052_; 
wire core__abc_22172_new_n6053_; 
wire core__abc_22172_new_n6054_; 
wire core__abc_22172_new_n6055_; 
wire core__abc_22172_new_n6056_; 
wire core__abc_22172_new_n6057_; 
wire core__abc_22172_new_n6058_; 
wire core__abc_22172_new_n6060_; 
wire core__abc_22172_new_n6061_; 
wire core__abc_22172_new_n6062_; 
wire core__abc_22172_new_n6063_; 
wire core__abc_22172_new_n6064_; 
wire core__abc_22172_new_n6065_; 
wire core__abc_22172_new_n6066_; 
wire core__abc_22172_new_n6067_; 
wire core__abc_22172_new_n6068_; 
wire core__abc_22172_new_n6069_; 
wire core__abc_22172_new_n6070_; 
wire core__abc_22172_new_n6071_; 
wire core__abc_22172_new_n6072_; 
wire core__abc_22172_new_n6073_; 
wire core__abc_22172_new_n6074_; 
wire core__abc_22172_new_n6075_; 
wire core__abc_22172_new_n6076_; 
wire core__abc_22172_new_n6077_; 
wire core__abc_22172_new_n6078_; 
wire core__abc_22172_new_n6079_; 
wire core__abc_22172_new_n6080_; 
wire core__abc_22172_new_n6081_; 
wire core__abc_22172_new_n6082_; 
wire core__abc_22172_new_n6083_; 
wire core__abc_22172_new_n6084_; 
wire core__abc_22172_new_n6085_; 
wire core__abc_22172_new_n6086_; 
wire core__abc_22172_new_n6087_; 
wire core__abc_22172_new_n6088_; 
wire core__abc_22172_new_n6089_; 
wire core__abc_22172_new_n6090_; 
wire core__abc_22172_new_n6091_; 
wire core__abc_22172_new_n6092_; 
wire core__abc_22172_new_n6093_; 
wire core__abc_22172_new_n6094_; 
wire core__abc_22172_new_n6095_; 
wire core__abc_22172_new_n6096_; 
wire core__abc_22172_new_n6097_; 
wire core__abc_22172_new_n6098_; 
wire core__abc_22172_new_n6099_; 
wire core__abc_22172_new_n6100_; 
wire core__abc_22172_new_n6102_; 
wire core__abc_22172_new_n6103_; 
wire core__abc_22172_new_n6104_; 
wire core__abc_22172_new_n6105_; 
wire core__abc_22172_new_n6106_; 
wire core__abc_22172_new_n6107_; 
wire core__abc_22172_new_n6108_; 
wire core__abc_22172_new_n6109_; 
wire core__abc_22172_new_n6110_; 
wire core__abc_22172_new_n6111_; 
wire core__abc_22172_new_n6112_; 
wire core__abc_22172_new_n6113_; 
wire core__abc_22172_new_n6114_; 
wire core__abc_22172_new_n6115_; 
wire core__abc_22172_new_n6116_; 
wire core__abc_22172_new_n6117_; 
wire core__abc_22172_new_n6118_; 
wire core__abc_22172_new_n6119_; 
wire core__abc_22172_new_n6120_; 
wire core__abc_22172_new_n6121_; 
wire core__abc_22172_new_n6122_; 
wire core__abc_22172_new_n6123_; 
wire core__abc_22172_new_n6124_; 
wire core__abc_22172_new_n6125_; 
wire core__abc_22172_new_n6126_; 
wire core__abc_22172_new_n6127_; 
wire core__abc_22172_new_n6128_; 
wire core__abc_22172_new_n6129_; 
wire core__abc_22172_new_n6130_; 
wire core__abc_22172_new_n6131_; 
wire core__abc_22172_new_n6132_; 
wire core__abc_22172_new_n6133_; 
wire core__abc_22172_new_n6134_; 
wire core__abc_22172_new_n6135_; 
wire core__abc_22172_new_n6136_; 
wire core__abc_22172_new_n6137_; 
wire core__abc_22172_new_n6138_; 
wire core__abc_22172_new_n6140_; 
wire core__abc_22172_new_n6141_; 
wire core__abc_22172_new_n6142_; 
wire core__abc_22172_new_n6143_; 
wire core__abc_22172_new_n6144_; 
wire core__abc_22172_new_n6145_; 
wire core__abc_22172_new_n6146_; 
wire core__abc_22172_new_n6147_; 
wire core__abc_22172_new_n6148_; 
wire core__abc_22172_new_n6149_; 
wire core__abc_22172_new_n6150_; 
wire core__abc_22172_new_n6151_; 
wire core__abc_22172_new_n6152_; 
wire core__abc_22172_new_n6153_; 
wire core__abc_22172_new_n6154_; 
wire core__abc_22172_new_n6155_; 
wire core__abc_22172_new_n6156_; 
wire core__abc_22172_new_n6157_; 
wire core__abc_22172_new_n6158_; 
wire core__abc_22172_new_n6159_; 
wire core__abc_22172_new_n6160_; 
wire core__abc_22172_new_n6161_; 
wire core__abc_22172_new_n6162_; 
wire core__abc_22172_new_n6163_; 
wire core__abc_22172_new_n6164_; 
wire core__abc_22172_new_n6165_; 
wire core__abc_22172_new_n6166_; 
wire core__abc_22172_new_n6167_; 
wire core__abc_22172_new_n6168_; 
wire core__abc_22172_new_n6169_; 
wire core__abc_22172_new_n6170_; 
wire core__abc_22172_new_n6171_; 
wire core__abc_22172_new_n6172_; 
wire core__abc_22172_new_n6173_; 
wire core__abc_22172_new_n6174_; 
wire core__abc_22172_new_n6175_; 
wire core__abc_22172_new_n6176_; 
wire core__abc_22172_new_n6177_; 
wire core__abc_22172_new_n6178_; 
wire core__abc_22172_new_n6179_; 
wire core__abc_22172_new_n6180_; 
wire core__abc_22172_new_n6181_; 
wire core__abc_22172_new_n6182_; 
wire core__abc_22172_new_n6183_; 
wire core__abc_22172_new_n6184_; 
wire core__abc_22172_new_n6185_; 
wire core__abc_22172_new_n6186_; 
wire core__abc_22172_new_n6187_; 
wire core__abc_22172_new_n6188_; 
wire core__abc_22172_new_n6189_; 
wire core__abc_22172_new_n6190_; 
wire core__abc_22172_new_n6191_; 
wire core__abc_22172_new_n6193_; 
wire core__abc_22172_new_n6194_; 
wire core__abc_22172_new_n6195_; 
wire core__abc_22172_new_n6196_; 
wire core__abc_22172_new_n6197_; 
wire core__abc_22172_new_n6198_; 
wire core__abc_22172_new_n6199_; 
wire core__abc_22172_new_n6200_; 
wire core__abc_22172_new_n6201_; 
wire core__abc_22172_new_n6202_; 
wire core__abc_22172_new_n6203_; 
wire core__abc_22172_new_n6204_; 
wire core__abc_22172_new_n6205_; 
wire core__abc_22172_new_n6206_; 
wire core__abc_22172_new_n6207_; 
wire core__abc_22172_new_n6208_; 
wire core__abc_22172_new_n6209_; 
wire core__abc_22172_new_n6210_; 
wire core__abc_22172_new_n6211_; 
wire core__abc_22172_new_n6212_; 
wire core__abc_22172_new_n6213_; 
wire core__abc_22172_new_n6214_; 
wire core__abc_22172_new_n6215_; 
wire core__abc_22172_new_n6216_; 
wire core__abc_22172_new_n6217_; 
wire core__abc_22172_new_n6218_; 
wire core__abc_22172_new_n6219_; 
wire core__abc_22172_new_n6220_; 
wire core__abc_22172_new_n6221_; 
wire core__abc_22172_new_n6222_; 
wire core__abc_22172_new_n6223_; 
wire core__abc_22172_new_n6225_; 
wire core__abc_22172_new_n6226_; 
wire core__abc_22172_new_n6227_; 
wire core__abc_22172_new_n6228_; 
wire core__abc_22172_new_n6229_; 
wire core__abc_22172_new_n6230_; 
wire core__abc_22172_new_n6231_; 
wire core__abc_22172_new_n6232_; 
wire core__abc_22172_new_n6233_; 
wire core__abc_22172_new_n6234_; 
wire core__abc_22172_new_n6235_; 
wire core__abc_22172_new_n6236_; 
wire core__abc_22172_new_n6237_; 
wire core__abc_22172_new_n6238_; 
wire core__abc_22172_new_n6239_; 
wire core__abc_22172_new_n6240_; 
wire core__abc_22172_new_n6241_; 
wire core__abc_22172_new_n6242_; 
wire core__abc_22172_new_n6243_; 
wire core__abc_22172_new_n6244_; 
wire core__abc_22172_new_n6245_; 
wire core__abc_22172_new_n6246_; 
wire core__abc_22172_new_n6247_; 
wire core__abc_22172_new_n6248_; 
wire core__abc_22172_new_n6249_; 
wire core__abc_22172_new_n6250_; 
wire core__abc_22172_new_n6251_; 
wire core__abc_22172_new_n6252_; 
wire core__abc_22172_new_n6253_; 
wire core__abc_22172_new_n6254_; 
wire core__abc_22172_new_n6255_; 
wire core__abc_22172_new_n6256_; 
wire core__abc_22172_new_n6257_; 
wire core__abc_22172_new_n6258_; 
wire core__abc_22172_new_n6259_; 
wire core__abc_22172_new_n6260_; 
wire core__abc_22172_new_n6261_; 
wire core__abc_22172_new_n6262_; 
wire core__abc_22172_new_n6263_; 
wire core__abc_22172_new_n6264_; 
wire core__abc_22172_new_n6265_; 
wire core__abc_22172_new_n6266_; 
wire core__abc_22172_new_n6268_; 
wire core__abc_22172_new_n6269_; 
wire core__abc_22172_new_n6270_; 
wire core__abc_22172_new_n6271_; 
wire core__abc_22172_new_n6272_; 
wire core__abc_22172_new_n6273_; 
wire core__abc_22172_new_n6274_; 
wire core__abc_22172_new_n6275_; 
wire core__abc_22172_new_n6276_; 
wire core__abc_22172_new_n6277_; 
wire core__abc_22172_new_n6278_; 
wire core__abc_22172_new_n6279_; 
wire core__abc_22172_new_n6280_; 
wire core__abc_22172_new_n6281_; 
wire core__abc_22172_new_n6282_; 
wire core__abc_22172_new_n6283_; 
wire core__abc_22172_new_n6284_; 
wire core__abc_22172_new_n6285_; 
wire core__abc_22172_new_n6286_; 
wire core__abc_22172_new_n6287_; 
wire core__abc_22172_new_n6288_; 
wire core__abc_22172_new_n6289_; 
wire core__abc_22172_new_n6290_; 
wire core__abc_22172_new_n6291_; 
wire core__abc_22172_new_n6292_; 
wire core__abc_22172_new_n6293_; 
wire core__abc_22172_new_n6294_; 
wire core__abc_22172_new_n6295_; 
wire core__abc_22172_new_n6296_; 
wire core__abc_22172_new_n6297_; 
wire core__abc_22172_new_n6298_; 
wire core__abc_22172_new_n6299_; 
wire core__abc_22172_new_n6300_; 
wire core__abc_22172_new_n6301_; 
wire core__abc_22172_new_n6303_; 
wire core__abc_22172_new_n6304_; 
wire core__abc_22172_new_n6305_; 
wire core__abc_22172_new_n6306_; 
wire core__abc_22172_new_n6307_; 
wire core__abc_22172_new_n6308_; 
wire core__abc_22172_new_n6309_; 
wire core__abc_22172_new_n6310_; 
wire core__abc_22172_new_n6311_; 
wire core__abc_22172_new_n6312_; 
wire core__abc_22172_new_n6313_; 
wire core__abc_22172_new_n6314_; 
wire core__abc_22172_new_n6315_; 
wire core__abc_22172_new_n6316_; 
wire core__abc_22172_new_n6317_; 
wire core__abc_22172_new_n6318_; 
wire core__abc_22172_new_n6319_; 
wire core__abc_22172_new_n6320_; 
wire core__abc_22172_new_n6321_; 
wire core__abc_22172_new_n6322_; 
wire core__abc_22172_new_n6323_; 
wire core__abc_22172_new_n6324_; 
wire core__abc_22172_new_n6325_; 
wire core__abc_22172_new_n6326_; 
wire core__abc_22172_new_n6327_; 
wire core__abc_22172_new_n6328_; 
wire core__abc_22172_new_n6329_; 
wire core__abc_22172_new_n6330_; 
wire core__abc_22172_new_n6331_; 
wire core__abc_22172_new_n6332_; 
wire core__abc_22172_new_n6333_; 
wire core__abc_22172_new_n6334_; 
wire core__abc_22172_new_n6335_; 
wire core__abc_22172_new_n6336_; 
wire core__abc_22172_new_n6337_; 
wire core__abc_22172_new_n6338_; 
wire core__abc_22172_new_n6339_; 
wire core__abc_22172_new_n6340_; 
wire core__abc_22172_new_n6341_; 
wire core__abc_22172_new_n6342_; 
wire core__abc_22172_new_n6343_; 
wire core__abc_22172_new_n6344_; 
wire core__abc_22172_new_n6345_; 
wire core__abc_22172_new_n6346_; 
wire core__abc_22172_new_n6347_; 
wire core__abc_22172_new_n6348_; 
wire core__abc_22172_new_n6349_; 
wire core__abc_22172_new_n6351_; 
wire core__abc_22172_new_n6352_; 
wire core__abc_22172_new_n6353_; 
wire core__abc_22172_new_n6354_; 
wire core__abc_22172_new_n6355_; 
wire core__abc_22172_new_n6356_; 
wire core__abc_22172_new_n6357_; 
wire core__abc_22172_new_n6358_; 
wire core__abc_22172_new_n6359_; 
wire core__abc_22172_new_n6360_; 
wire core__abc_22172_new_n6361_; 
wire core__abc_22172_new_n6362_; 
wire core__abc_22172_new_n6363_; 
wire core__abc_22172_new_n6364_; 
wire core__abc_22172_new_n6365_; 
wire core__abc_22172_new_n6366_; 
wire core__abc_22172_new_n6367_; 
wire core__abc_22172_new_n6368_; 
wire core__abc_22172_new_n6369_; 
wire core__abc_22172_new_n6370_; 
wire core__abc_22172_new_n6371_; 
wire core__abc_22172_new_n6372_; 
wire core__abc_22172_new_n6373_; 
wire core__abc_22172_new_n6374_; 
wire core__abc_22172_new_n6375_; 
wire core__abc_22172_new_n6376_; 
wire core__abc_22172_new_n6377_; 
wire core__abc_22172_new_n6378_; 
wire core__abc_22172_new_n6379_; 
wire core__abc_22172_new_n6380_; 
wire core__abc_22172_new_n6381_; 
wire core__abc_22172_new_n6382_; 
wire core__abc_22172_new_n6383_; 
wire core__abc_22172_new_n6384_; 
wire core__abc_22172_new_n6385_; 
wire core__abc_22172_new_n6386_; 
wire core__abc_22172_new_n6387_; 
wire core__abc_22172_new_n6388_; 
wire core__abc_22172_new_n6390_; 
wire core__abc_22172_new_n6391_; 
wire core__abc_22172_new_n6392_; 
wire core__abc_22172_new_n6393_; 
wire core__abc_22172_new_n6394_; 
wire core__abc_22172_new_n6395_; 
wire core__abc_22172_new_n6396_; 
wire core__abc_22172_new_n6397_; 
wire core__abc_22172_new_n6398_; 
wire core__abc_22172_new_n6399_; 
wire core__abc_22172_new_n6400_; 
wire core__abc_22172_new_n6401_; 
wire core__abc_22172_new_n6402_; 
wire core__abc_22172_new_n6403_; 
wire core__abc_22172_new_n6404_; 
wire core__abc_22172_new_n6405_; 
wire core__abc_22172_new_n6406_; 
wire core__abc_22172_new_n6407_; 
wire core__abc_22172_new_n6408_; 
wire core__abc_22172_new_n6409_; 
wire core__abc_22172_new_n6410_; 
wire core__abc_22172_new_n6411_; 
wire core__abc_22172_new_n6412_; 
wire core__abc_22172_new_n6413_; 
wire core__abc_22172_new_n6414_; 
wire core__abc_22172_new_n6415_; 
wire core__abc_22172_new_n6416_; 
wire core__abc_22172_new_n6417_; 
wire core__abc_22172_new_n6418_; 
wire core__abc_22172_new_n6419_; 
wire core__abc_22172_new_n6420_; 
wire core__abc_22172_new_n6421_; 
wire core__abc_22172_new_n6422_; 
wire core__abc_22172_new_n6423_; 
wire core__abc_22172_new_n6424_; 
wire core__abc_22172_new_n6425_; 
wire core__abc_22172_new_n6426_; 
wire core__abc_22172_new_n6427_; 
wire core__abc_22172_new_n6428_; 
wire core__abc_22172_new_n6429_; 
wire core__abc_22172_new_n6430_; 
wire core__abc_22172_new_n6431_; 
wire core__abc_22172_new_n6433_; 
wire core__abc_22172_new_n6434_; 
wire core__abc_22172_new_n6435_; 
wire core__abc_22172_new_n6436_; 
wire core__abc_22172_new_n6437_; 
wire core__abc_22172_new_n6438_; 
wire core__abc_22172_new_n6439_; 
wire core__abc_22172_new_n6440_; 
wire core__abc_22172_new_n6441_; 
wire core__abc_22172_new_n6442_; 
wire core__abc_22172_new_n6443_; 
wire core__abc_22172_new_n6444_; 
wire core__abc_22172_new_n6445_; 
wire core__abc_22172_new_n6446_; 
wire core__abc_22172_new_n6447_; 
wire core__abc_22172_new_n6448_; 
wire core__abc_22172_new_n6449_; 
wire core__abc_22172_new_n6450_; 
wire core__abc_22172_new_n6451_; 
wire core__abc_22172_new_n6452_; 
wire core__abc_22172_new_n6453_; 
wire core__abc_22172_new_n6454_; 
wire core__abc_22172_new_n6455_; 
wire core__abc_22172_new_n6456_; 
wire core__abc_22172_new_n6457_; 
wire core__abc_22172_new_n6458_; 
wire core__abc_22172_new_n6459_; 
wire core__abc_22172_new_n6460_; 
wire core__abc_22172_new_n6461_; 
wire core__abc_22172_new_n6462_; 
wire core__abc_22172_new_n6463_; 
wire core__abc_22172_new_n6464_; 
wire core__abc_22172_new_n6465_; 
wire core__abc_22172_new_n6466_; 
wire core__abc_22172_new_n6468_; 
wire core__abc_22172_new_n6469_; 
wire core__abc_22172_new_n6470_; 
wire core__abc_22172_new_n6471_; 
wire core__abc_22172_new_n6472_; 
wire core__abc_22172_new_n6473_; 
wire core__abc_22172_new_n6474_; 
wire core__abc_22172_new_n6475_; 
wire core__abc_22172_new_n6476_; 
wire core__abc_22172_new_n6477_; 
wire core__abc_22172_new_n6478_; 
wire core__abc_22172_new_n6479_; 
wire core__abc_22172_new_n6480_; 
wire core__abc_22172_new_n6481_; 
wire core__abc_22172_new_n6482_; 
wire core__abc_22172_new_n6483_; 
wire core__abc_22172_new_n6484_; 
wire core__abc_22172_new_n6485_; 
wire core__abc_22172_new_n6486_; 
wire core__abc_22172_new_n6487_; 
wire core__abc_22172_new_n6488_; 
wire core__abc_22172_new_n6489_; 
wire core__abc_22172_new_n6490_; 
wire core__abc_22172_new_n6491_; 
wire core__abc_22172_new_n6492_; 
wire core__abc_22172_new_n6493_; 
wire core__abc_22172_new_n6494_; 
wire core__abc_22172_new_n6495_; 
wire core__abc_22172_new_n6496_; 
wire core__abc_22172_new_n6497_; 
wire core__abc_22172_new_n6498_; 
wire core__abc_22172_new_n6499_; 
wire core__abc_22172_new_n6500_; 
wire core__abc_22172_new_n6501_; 
wire core__abc_22172_new_n6502_; 
wire core__abc_22172_new_n6503_; 
wire core__abc_22172_new_n6504_; 
wire core__abc_22172_new_n6505_; 
wire core__abc_22172_new_n6506_; 
wire core__abc_22172_new_n6507_; 
wire core__abc_22172_new_n6508_; 
wire core__abc_22172_new_n6509_; 
wire core__abc_22172_new_n6510_; 
wire core__abc_22172_new_n6511_; 
wire core__abc_22172_new_n6512_; 
wire core__abc_22172_new_n6513_; 
wire core__abc_22172_new_n6514_; 
wire core__abc_22172_new_n6515_; 
wire core__abc_22172_new_n6516_; 
wire core__abc_22172_new_n6517_; 
wire core__abc_22172_new_n6518_; 
wire core__abc_22172_new_n6519_; 
wire core__abc_22172_new_n6520_; 
wire core__abc_22172_new_n6521_; 
wire core__abc_22172_new_n6522_; 
wire core__abc_22172_new_n6523_; 
wire core__abc_22172_new_n6524_; 
wire core__abc_22172_new_n6525_; 
wire core__abc_22172_new_n6526_; 
wire core__abc_22172_new_n6527_; 
wire core__abc_22172_new_n6528_; 
wire core__abc_22172_new_n6529_; 
wire core__abc_22172_new_n6530_; 
wire core__abc_22172_new_n6531_; 
wire core__abc_22172_new_n6532_; 
wire core__abc_22172_new_n6533_; 
wire core__abc_22172_new_n6534_; 
wire core__abc_22172_new_n6535_; 
wire core__abc_22172_new_n6536_; 
wire core__abc_22172_new_n6537_; 
wire core__abc_22172_new_n6538_; 
wire core__abc_22172_new_n6539_; 
wire core__abc_22172_new_n6540_; 
wire core__abc_22172_new_n6541_; 
wire core__abc_22172_new_n6542_; 
wire core__abc_22172_new_n6543_; 
wire core__abc_22172_new_n6544_; 
wire core__abc_22172_new_n6545_; 
wire core__abc_22172_new_n6546_; 
wire core__abc_22172_new_n6547_; 
wire core__abc_22172_new_n6548_; 
wire core__abc_22172_new_n6549_; 
wire core__abc_22172_new_n6550_; 
wire core__abc_22172_new_n6551_; 
wire core__abc_22172_new_n6552_; 
wire core__abc_22172_new_n6553_; 
wire core__abc_22172_new_n6554_; 
wire core__abc_22172_new_n6555_; 
wire core__abc_22172_new_n6556_; 
wire core__abc_22172_new_n6557_; 
wire core__abc_22172_new_n6558_; 
wire core__abc_22172_new_n6559_; 
wire core__abc_22172_new_n6560_; 
wire core__abc_22172_new_n6561_; 
wire core__abc_22172_new_n6562_; 
wire core__abc_22172_new_n6563_; 
wire core__abc_22172_new_n6564_; 
wire core__abc_22172_new_n6565_; 
wire core__abc_22172_new_n6566_; 
wire core__abc_22172_new_n6567_; 
wire core__abc_22172_new_n6568_; 
wire core__abc_22172_new_n6569_; 
wire core__abc_22172_new_n6570_; 
wire core__abc_22172_new_n6571_; 
wire core__abc_22172_new_n6572_; 
wire core__abc_22172_new_n6573_; 
wire core__abc_22172_new_n6574_; 
wire core__abc_22172_new_n6575_; 
wire core__abc_22172_new_n6576_; 
wire core__abc_22172_new_n6577_; 
wire core__abc_22172_new_n6578_; 
wire core__abc_22172_new_n6579_; 
wire core__abc_22172_new_n6580_; 
wire core__abc_22172_new_n6581_; 
wire core__abc_22172_new_n6582_; 
wire core__abc_22172_new_n6583_; 
wire core__abc_22172_new_n6584_; 
wire core__abc_22172_new_n6585_; 
wire core__abc_22172_new_n6586_; 
wire core__abc_22172_new_n6587_; 
wire core__abc_22172_new_n6588_; 
wire core__abc_22172_new_n6589_; 
wire core__abc_22172_new_n6590_; 
wire core__abc_22172_new_n6591_; 
wire core__abc_22172_new_n6592_; 
wire core__abc_22172_new_n6593_; 
wire core__abc_22172_new_n6594_; 
wire core__abc_22172_new_n6595_; 
wire core__abc_22172_new_n6596_; 
wire core__abc_22172_new_n6597_; 
wire core__abc_22172_new_n6598_; 
wire core__abc_22172_new_n6599_; 
wire core__abc_22172_new_n6600_; 
wire core__abc_22172_new_n6601_; 
wire core__abc_22172_new_n6602_; 
wire core__abc_22172_new_n6603_; 
wire core__abc_22172_new_n6604_; 
wire core__abc_22172_new_n6605_; 
wire core__abc_22172_new_n6606_; 
wire core__abc_22172_new_n6607_; 
wire core__abc_22172_new_n6608_; 
wire core__abc_22172_new_n6609_; 
wire core__abc_22172_new_n6610_; 
wire core__abc_22172_new_n6611_; 
wire core__abc_22172_new_n6612_; 
wire core__abc_22172_new_n6613_; 
wire core__abc_22172_new_n6614_; 
wire core__abc_22172_new_n6615_; 
wire core__abc_22172_new_n6616_; 
wire core__abc_22172_new_n6617_; 
wire core__abc_22172_new_n6618_; 
wire core__abc_22172_new_n6619_; 
wire core__abc_22172_new_n6620_; 
wire core__abc_22172_new_n6621_; 
wire core__abc_22172_new_n6622_; 
wire core__abc_22172_new_n6623_; 
wire core__abc_22172_new_n6624_; 
wire core__abc_22172_new_n6625_; 
wire core__abc_22172_new_n6626_; 
wire core__abc_22172_new_n6627_; 
wire core__abc_22172_new_n6628_; 
wire core__abc_22172_new_n6629_; 
wire core__abc_22172_new_n6630_; 
wire core__abc_22172_new_n6631_; 
wire core__abc_22172_new_n6632_; 
wire core__abc_22172_new_n6633_; 
wire core__abc_22172_new_n6634_; 
wire core__abc_22172_new_n6635_; 
wire core__abc_22172_new_n6636_; 
wire core__abc_22172_new_n6637_; 
wire core__abc_22172_new_n6638_; 
wire core__abc_22172_new_n6639_; 
wire core__abc_22172_new_n6640_; 
wire core__abc_22172_new_n6641_; 
wire core__abc_22172_new_n6642_; 
wire core__abc_22172_new_n6643_; 
wire core__abc_22172_new_n6644_; 
wire core__abc_22172_new_n6645_; 
wire core__abc_22172_new_n6646_; 
wire core__abc_22172_new_n6647_; 
wire core__abc_22172_new_n6648_; 
wire core__abc_22172_new_n6649_; 
wire core__abc_22172_new_n6650_; 
wire core__abc_22172_new_n6651_; 
wire core__abc_22172_new_n6652_; 
wire core__abc_22172_new_n6653_; 
wire core__abc_22172_new_n6654_; 
wire core__abc_22172_new_n6655_; 
wire core__abc_22172_new_n6656_; 
wire core__abc_22172_new_n6657_; 
wire core__abc_22172_new_n6658_; 
wire core__abc_22172_new_n6659_; 
wire core__abc_22172_new_n6660_; 
wire core__abc_22172_new_n6661_; 
wire core__abc_22172_new_n6662_; 
wire core__abc_22172_new_n6663_; 
wire core__abc_22172_new_n6664_; 
wire core__abc_22172_new_n6665_; 
wire core__abc_22172_new_n6666_; 
wire core__abc_22172_new_n6667_; 
wire core__abc_22172_new_n6668_; 
wire core__abc_22172_new_n6669_; 
wire core__abc_22172_new_n6670_; 
wire core__abc_22172_new_n6671_; 
wire core__abc_22172_new_n6672_; 
wire core__abc_22172_new_n6673_; 
wire core__abc_22172_new_n6674_; 
wire core__abc_22172_new_n6675_; 
wire core__abc_22172_new_n6676_; 
wire core__abc_22172_new_n6677_; 
wire core__abc_22172_new_n6678_; 
wire core__abc_22172_new_n6679_; 
wire core__abc_22172_new_n6680_; 
wire core__abc_22172_new_n6681_; 
wire core__abc_22172_new_n6682_; 
wire core__abc_22172_new_n6683_; 
wire core__abc_22172_new_n6684_; 
wire core__abc_22172_new_n6685_; 
wire core__abc_22172_new_n6686_; 
wire core__abc_22172_new_n6687_; 
wire core__abc_22172_new_n6688_; 
wire core__abc_22172_new_n6689_; 
wire core__abc_22172_new_n6690_; 
wire core__abc_22172_new_n6691_; 
wire core__abc_22172_new_n6692_; 
wire core__abc_22172_new_n6693_; 
wire core__abc_22172_new_n6694_; 
wire core__abc_22172_new_n6695_; 
wire core__abc_22172_new_n6696_; 
wire core__abc_22172_new_n6697_; 
wire core__abc_22172_new_n6698_; 
wire core__abc_22172_new_n6699_; 
wire core__abc_22172_new_n6700_; 
wire core__abc_22172_new_n6701_; 
wire core__abc_22172_new_n6702_; 
wire core__abc_22172_new_n6703_; 
wire core__abc_22172_new_n6704_; 
wire core__abc_22172_new_n6705_; 
wire core__abc_22172_new_n6706_; 
wire core__abc_22172_new_n6707_; 
wire core__abc_22172_new_n6708_; 
wire core__abc_22172_new_n6709_; 
wire core__abc_22172_new_n6710_; 
wire core__abc_22172_new_n6711_; 
wire core__abc_22172_new_n6712_; 
wire core__abc_22172_new_n6713_; 
wire core__abc_22172_new_n6714_; 
wire core__abc_22172_new_n6715_; 
wire core__abc_22172_new_n6716_; 
wire core__abc_22172_new_n6717_; 
wire core__abc_22172_new_n6718_; 
wire core__abc_22172_new_n6719_; 
wire core__abc_22172_new_n6720_; 
wire core__abc_22172_new_n6721_; 
wire core__abc_22172_new_n6722_; 
wire core__abc_22172_new_n6723_; 
wire core__abc_22172_new_n6724_; 
wire core__abc_22172_new_n6725_; 
wire core__abc_22172_new_n6726_; 
wire core__abc_22172_new_n6727_; 
wire core__abc_22172_new_n6728_; 
wire core__abc_22172_new_n6729_; 
wire core__abc_22172_new_n6730_; 
wire core__abc_22172_new_n6731_; 
wire core__abc_22172_new_n6732_; 
wire core__abc_22172_new_n6733_; 
wire core__abc_22172_new_n6734_; 
wire core__abc_22172_new_n6735_; 
wire core__abc_22172_new_n6736_; 
wire core__abc_22172_new_n6737_; 
wire core__abc_22172_new_n6738_; 
wire core__abc_22172_new_n6739_; 
wire core__abc_22172_new_n6740_; 
wire core__abc_22172_new_n6741_; 
wire core__abc_22172_new_n6742_; 
wire core__abc_22172_new_n6743_; 
wire core__abc_22172_new_n6744_; 
wire core__abc_22172_new_n6745_; 
wire core__abc_22172_new_n6746_; 
wire core__abc_22172_new_n6747_; 
wire core__abc_22172_new_n6748_; 
wire core__abc_22172_new_n6749_; 
wire core__abc_22172_new_n6750_; 
wire core__abc_22172_new_n6751_; 
wire core__abc_22172_new_n6752_; 
wire core__abc_22172_new_n6753_; 
wire core__abc_22172_new_n6754_; 
wire core__abc_22172_new_n6755_; 
wire core__abc_22172_new_n6756_; 
wire core__abc_22172_new_n6757_; 
wire core__abc_22172_new_n6758_; 
wire core__abc_22172_new_n6759_; 
wire core__abc_22172_new_n6760_; 
wire core__abc_22172_new_n6761_; 
wire core__abc_22172_new_n6762_; 
wire core__abc_22172_new_n6763_; 
wire core__abc_22172_new_n6764_; 
wire core__abc_22172_new_n6765_; 
wire core__abc_22172_new_n6766_; 
wire core__abc_22172_new_n6767_; 
wire core__abc_22172_new_n6768_; 
wire core__abc_22172_new_n6769_; 
wire core__abc_22172_new_n6770_; 
wire core__abc_22172_new_n6771_; 
wire core__abc_22172_new_n6772_; 
wire core__abc_22172_new_n6773_; 
wire core__abc_22172_new_n6774_; 
wire core__abc_22172_new_n6775_; 
wire core__abc_22172_new_n6776_; 
wire core__abc_22172_new_n6777_; 
wire core__abc_22172_new_n6778_; 
wire core__abc_22172_new_n6779_; 
wire core__abc_22172_new_n6780_; 
wire core__abc_22172_new_n6781_; 
wire core__abc_22172_new_n6782_; 
wire core__abc_22172_new_n6783_; 
wire core__abc_22172_new_n6784_; 
wire core__abc_22172_new_n6785_; 
wire core__abc_22172_new_n6786_; 
wire core__abc_22172_new_n6787_; 
wire core__abc_22172_new_n6788_; 
wire core__abc_22172_new_n6789_; 
wire core__abc_22172_new_n6790_; 
wire core__abc_22172_new_n6791_; 
wire core__abc_22172_new_n6792_; 
wire core__abc_22172_new_n6793_; 
wire core__abc_22172_new_n6794_; 
wire core__abc_22172_new_n6795_; 
wire core__abc_22172_new_n6796_; 
wire core__abc_22172_new_n6797_; 
wire core__abc_22172_new_n6798_; 
wire core__abc_22172_new_n6799_; 
wire core__abc_22172_new_n6800_; 
wire core__abc_22172_new_n6801_; 
wire core__abc_22172_new_n6802_; 
wire core__abc_22172_new_n6803_; 
wire core__abc_22172_new_n6804_; 
wire core__abc_22172_new_n6805_; 
wire core__abc_22172_new_n6806_; 
wire core__abc_22172_new_n6807_; 
wire core__abc_22172_new_n6808_; 
wire core__abc_22172_new_n6809_; 
wire core__abc_22172_new_n6810_; 
wire core__abc_22172_new_n6811_; 
wire core__abc_22172_new_n6812_; 
wire core__abc_22172_new_n6813_; 
wire core__abc_22172_new_n6814_; 
wire core__abc_22172_new_n6815_; 
wire core__abc_22172_new_n6816_; 
wire core__abc_22172_new_n6817_; 
wire core__abc_22172_new_n6818_; 
wire core__abc_22172_new_n6819_; 
wire core__abc_22172_new_n6820_; 
wire core__abc_22172_new_n6821_; 
wire core__abc_22172_new_n6822_; 
wire core__abc_22172_new_n6823_; 
wire core__abc_22172_new_n6824_; 
wire core__abc_22172_new_n6825_; 
wire core__abc_22172_new_n6826_; 
wire core__abc_22172_new_n6827_; 
wire core__abc_22172_new_n6828_; 
wire core__abc_22172_new_n6829_; 
wire core__abc_22172_new_n6830_; 
wire core__abc_22172_new_n6831_; 
wire core__abc_22172_new_n6832_; 
wire core__abc_22172_new_n6833_; 
wire core__abc_22172_new_n6834_; 
wire core__abc_22172_new_n6835_; 
wire core__abc_22172_new_n6836_; 
wire core__abc_22172_new_n6837_; 
wire core__abc_22172_new_n6838_; 
wire core__abc_22172_new_n6839_; 
wire core__abc_22172_new_n6840_; 
wire core__abc_22172_new_n6841_; 
wire core__abc_22172_new_n6842_; 
wire core__abc_22172_new_n6843_; 
wire core__abc_22172_new_n6844_; 
wire core__abc_22172_new_n6845_; 
wire core__abc_22172_new_n6846_; 
wire core__abc_22172_new_n6847_; 
wire core__abc_22172_new_n6848_; 
wire core__abc_22172_new_n6849_; 
wire core__abc_22172_new_n6850_; 
wire core__abc_22172_new_n6851_; 
wire core__abc_22172_new_n6852_; 
wire core__abc_22172_new_n6853_; 
wire core__abc_22172_new_n6854_; 
wire core__abc_22172_new_n6855_; 
wire core__abc_22172_new_n6856_; 
wire core__abc_22172_new_n6857_; 
wire core__abc_22172_new_n6858_; 
wire core__abc_22172_new_n6859_; 
wire core__abc_22172_new_n6860_; 
wire core__abc_22172_new_n6861_; 
wire core__abc_22172_new_n6862_; 
wire core__abc_22172_new_n6863_; 
wire core__abc_22172_new_n6864_; 
wire core__abc_22172_new_n6865_; 
wire core__abc_22172_new_n6866_; 
wire core__abc_22172_new_n6867_; 
wire core__abc_22172_new_n6868_; 
wire core__abc_22172_new_n6869_; 
wire core__abc_22172_new_n6870_; 
wire core__abc_22172_new_n6871_; 
wire core__abc_22172_new_n6872_; 
wire core__abc_22172_new_n6873_; 
wire core__abc_22172_new_n6874_; 
wire core__abc_22172_new_n6875_; 
wire core__abc_22172_new_n6876_; 
wire core__abc_22172_new_n6877_; 
wire core__abc_22172_new_n6878_; 
wire core__abc_22172_new_n6879_; 
wire core__abc_22172_new_n6880_; 
wire core__abc_22172_new_n6881_; 
wire core__abc_22172_new_n6882_; 
wire core__abc_22172_new_n6884_; 
wire core__abc_22172_new_n6885_; 
wire core__abc_22172_new_n6886_; 
wire core__abc_22172_new_n6887_; 
wire core__abc_22172_new_n6888_; 
wire core__abc_22172_new_n6889_; 
wire core__abc_22172_new_n6890_; 
wire core__abc_22172_new_n6891_; 
wire core__abc_22172_new_n6892_; 
wire core__abc_22172_new_n6893_; 
wire core__abc_22172_new_n6894_; 
wire core__abc_22172_new_n6895_; 
wire core__abc_22172_new_n6896_; 
wire core__abc_22172_new_n6897_; 
wire core__abc_22172_new_n6898_; 
wire core__abc_22172_new_n6899_; 
wire core__abc_22172_new_n6900_; 
wire core__abc_22172_new_n6901_; 
wire core__abc_22172_new_n6902_; 
wire core__abc_22172_new_n6903_; 
wire core__abc_22172_new_n6904_; 
wire core__abc_22172_new_n6905_; 
wire core__abc_22172_new_n6906_; 
wire core__abc_22172_new_n6907_; 
wire core__abc_22172_new_n6908_; 
wire core__abc_22172_new_n6909_; 
wire core__abc_22172_new_n6911_; 
wire core__abc_22172_new_n6912_; 
wire core__abc_22172_new_n6913_; 
wire core__abc_22172_new_n6914_; 
wire core__abc_22172_new_n6915_; 
wire core__abc_22172_new_n6916_; 
wire core__abc_22172_new_n6917_; 
wire core__abc_22172_new_n6918_; 
wire core__abc_22172_new_n6919_; 
wire core__abc_22172_new_n6920_; 
wire core__abc_22172_new_n6921_; 
wire core__abc_22172_new_n6922_; 
wire core__abc_22172_new_n6923_; 
wire core__abc_22172_new_n6924_; 
wire core__abc_22172_new_n6925_; 
wire core__abc_22172_new_n6926_; 
wire core__abc_22172_new_n6927_; 
wire core__abc_22172_new_n6928_; 
wire core__abc_22172_new_n6929_; 
wire core__abc_22172_new_n6930_; 
wire core__abc_22172_new_n6931_; 
wire core__abc_22172_new_n6932_; 
wire core__abc_22172_new_n6933_; 
wire core__abc_22172_new_n6934_; 
wire core__abc_22172_new_n6935_; 
wire core__abc_22172_new_n6936_; 
wire core__abc_22172_new_n6937_; 
wire core__abc_22172_new_n6939_; 
wire core__abc_22172_new_n6940_; 
wire core__abc_22172_new_n6941_; 
wire core__abc_22172_new_n6942_; 
wire core__abc_22172_new_n6943_; 
wire core__abc_22172_new_n6944_; 
wire core__abc_22172_new_n6945_; 
wire core__abc_22172_new_n6946_; 
wire core__abc_22172_new_n6947_; 
wire core__abc_22172_new_n6948_; 
wire core__abc_22172_new_n6949_; 
wire core__abc_22172_new_n6950_; 
wire core__abc_22172_new_n6951_; 
wire core__abc_22172_new_n6952_; 
wire core__abc_22172_new_n6953_; 
wire core__abc_22172_new_n6954_; 
wire core__abc_22172_new_n6955_; 
wire core__abc_22172_new_n6956_; 
wire core__abc_22172_new_n6957_; 
wire core__abc_22172_new_n6958_; 
wire core__abc_22172_new_n6959_; 
wire core__abc_22172_new_n6960_; 
wire core__abc_22172_new_n6962_; 
wire core__abc_22172_new_n6963_; 
wire core__abc_22172_new_n6964_; 
wire core__abc_22172_new_n6965_; 
wire core__abc_22172_new_n6966_; 
wire core__abc_22172_new_n6967_; 
wire core__abc_22172_new_n6968_; 
wire core__abc_22172_new_n6969_; 
wire core__abc_22172_new_n6970_; 
wire core__abc_22172_new_n6971_; 
wire core__abc_22172_new_n6972_; 
wire core__abc_22172_new_n6973_; 
wire core__abc_22172_new_n6974_; 
wire core__abc_22172_new_n6975_; 
wire core__abc_22172_new_n6976_; 
wire core__abc_22172_new_n6977_; 
wire core__abc_22172_new_n6978_; 
wire core__abc_22172_new_n6979_; 
wire core__abc_22172_new_n6980_; 
wire core__abc_22172_new_n6981_; 
wire core__abc_22172_new_n6982_; 
wire core__abc_22172_new_n6983_; 
wire core__abc_22172_new_n6984_; 
wire core__abc_22172_new_n6985_; 
wire core__abc_22172_new_n6986_; 
wire core__abc_22172_new_n6987_; 
wire core__abc_22172_new_n6988_; 
wire core__abc_22172_new_n6989_; 
wire core__abc_22172_new_n6990_; 
wire core__abc_22172_new_n6992_; 
wire core__abc_22172_new_n6993_; 
wire core__abc_22172_new_n6994_; 
wire core__abc_22172_new_n6995_; 
wire core__abc_22172_new_n6996_; 
wire core__abc_22172_new_n6997_; 
wire core__abc_22172_new_n6998_; 
wire core__abc_22172_new_n6999_; 
wire core__abc_22172_new_n7000_; 
wire core__abc_22172_new_n7001_; 
wire core__abc_22172_new_n7002_; 
wire core__abc_22172_new_n7003_; 
wire core__abc_22172_new_n7004_; 
wire core__abc_22172_new_n7005_; 
wire core__abc_22172_new_n7006_; 
wire core__abc_22172_new_n7007_; 
wire core__abc_22172_new_n7008_; 
wire core__abc_22172_new_n7009_; 
wire core__abc_22172_new_n7010_; 
wire core__abc_22172_new_n7011_; 
wire core__abc_22172_new_n7012_; 
wire core__abc_22172_new_n7013_; 
wire core__abc_22172_new_n7014_; 
wire core__abc_22172_new_n7015_; 
wire core__abc_22172_new_n7016_; 
wire core__abc_22172_new_n7018_; 
wire core__abc_22172_new_n7019_; 
wire core__abc_22172_new_n7020_; 
wire core__abc_22172_new_n7021_; 
wire core__abc_22172_new_n7022_; 
wire core__abc_22172_new_n7023_; 
wire core__abc_22172_new_n7024_; 
wire core__abc_22172_new_n7025_; 
wire core__abc_22172_new_n7026_; 
wire core__abc_22172_new_n7027_; 
wire core__abc_22172_new_n7028_; 
wire core__abc_22172_new_n7029_; 
wire core__abc_22172_new_n7030_; 
wire core__abc_22172_new_n7031_; 
wire core__abc_22172_new_n7032_; 
wire core__abc_22172_new_n7033_; 
wire core__abc_22172_new_n7034_; 
wire core__abc_22172_new_n7035_; 
wire core__abc_22172_new_n7036_; 
wire core__abc_22172_new_n7037_; 
wire core__abc_22172_new_n7038_; 
wire core__abc_22172_new_n7039_; 
wire core__abc_22172_new_n7040_; 
wire core__abc_22172_new_n7041_; 
wire core__abc_22172_new_n7042_; 
wire core__abc_22172_new_n7043_; 
wire core__abc_22172_new_n7044_; 
wire core__abc_22172_new_n7045_; 
wire core__abc_22172_new_n7046_; 
wire core__abc_22172_new_n7048_; 
wire core__abc_22172_new_n7049_; 
wire core__abc_22172_new_n7050_; 
wire core__abc_22172_new_n7051_; 
wire core__abc_22172_new_n7052_; 
wire core__abc_22172_new_n7053_; 
wire core__abc_22172_new_n7054_; 
wire core__abc_22172_new_n7055_; 
wire core__abc_22172_new_n7056_; 
wire core__abc_22172_new_n7057_; 
wire core__abc_22172_new_n7058_; 
wire core__abc_22172_new_n7059_; 
wire core__abc_22172_new_n7060_; 
wire core__abc_22172_new_n7061_; 
wire core__abc_22172_new_n7062_; 
wire core__abc_22172_new_n7063_; 
wire core__abc_22172_new_n7064_; 
wire core__abc_22172_new_n7065_; 
wire core__abc_22172_new_n7066_; 
wire core__abc_22172_new_n7067_; 
wire core__abc_22172_new_n7068_; 
wire core__abc_22172_new_n7069_; 
wire core__abc_22172_new_n7070_; 
wire core__abc_22172_new_n7072_; 
wire core__abc_22172_new_n7073_; 
wire core__abc_22172_new_n7074_; 
wire core__abc_22172_new_n7075_; 
wire core__abc_22172_new_n7076_; 
wire core__abc_22172_new_n7077_; 
wire core__abc_22172_new_n7078_; 
wire core__abc_22172_new_n7079_; 
wire core__abc_22172_new_n7080_; 
wire core__abc_22172_new_n7081_; 
wire core__abc_22172_new_n7082_; 
wire core__abc_22172_new_n7083_; 
wire core__abc_22172_new_n7084_; 
wire core__abc_22172_new_n7085_; 
wire core__abc_22172_new_n7086_; 
wire core__abc_22172_new_n7087_; 
wire core__abc_22172_new_n7088_; 
wire core__abc_22172_new_n7089_; 
wire core__abc_22172_new_n7090_; 
wire core__abc_22172_new_n7091_; 
wire core__abc_22172_new_n7092_; 
wire core__abc_22172_new_n7093_; 
wire core__abc_22172_new_n7094_; 
wire core__abc_22172_new_n7095_; 
wire core__abc_22172_new_n7096_; 
wire core__abc_22172_new_n7097_; 
wire core__abc_22172_new_n7098_; 
wire core__abc_22172_new_n7099_; 
wire core__abc_22172_new_n7100_; 
wire core__abc_22172_new_n7101_; 
wire core__abc_22172_new_n7102_; 
wire core__abc_22172_new_n7103_; 
wire core__abc_22172_new_n7104_; 
wire core__abc_22172_new_n7105_; 
wire core__abc_22172_new_n7106_; 
wire core__abc_22172_new_n7107_; 
wire core__abc_22172_new_n7108_; 
wire core__abc_22172_new_n7109_; 
wire core__abc_22172_new_n7110_; 
wire core__abc_22172_new_n7111_; 
wire core__abc_22172_new_n7112_; 
wire core__abc_22172_new_n7113_; 
wire core__abc_22172_new_n7114_; 
wire core__abc_22172_new_n7115_; 
wire core__abc_22172_new_n7116_; 
wire core__abc_22172_new_n7118_; 
wire core__abc_22172_new_n7119_; 
wire core__abc_22172_new_n7120_; 
wire core__abc_22172_new_n7121_; 
wire core__abc_22172_new_n7122_; 
wire core__abc_22172_new_n7123_; 
wire core__abc_22172_new_n7124_; 
wire core__abc_22172_new_n7125_; 
wire core__abc_22172_new_n7126_; 
wire core__abc_22172_new_n7127_; 
wire core__abc_22172_new_n7128_; 
wire core__abc_22172_new_n7129_; 
wire core__abc_22172_new_n7130_; 
wire core__abc_22172_new_n7131_; 
wire core__abc_22172_new_n7132_; 
wire core__abc_22172_new_n7133_; 
wire core__abc_22172_new_n7134_; 
wire core__abc_22172_new_n7135_; 
wire core__abc_22172_new_n7136_; 
wire core__abc_22172_new_n7137_; 
wire core__abc_22172_new_n7138_; 
wire core__abc_22172_new_n7139_; 
wire core__abc_22172_new_n7140_; 
wire core__abc_22172_new_n7141_; 
wire core__abc_22172_new_n7142_; 
wire core__abc_22172_new_n7143_; 
wire core__abc_22172_new_n7144_; 
wire core__abc_22172_new_n7146_; 
wire core__abc_22172_new_n7147_; 
wire core__abc_22172_new_n7148_; 
wire core__abc_22172_new_n7149_; 
wire core__abc_22172_new_n7150_; 
wire core__abc_22172_new_n7151_; 
wire core__abc_22172_new_n7152_; 
wire core__abc_22172_new_n7153_; 
wire core__abc_22172_new_n7154_; 
wire core__abc_22172_new_n7155_; 
wire core__abc_22172_new_n7156_; 
wire core__abc_22172_new_n7157_; 
wire core__abc_22172_new_n7158_; 
wire core__abc_22172_new_n7159_; 
wire core__abc_22172_new_n7160_; 
wire core__abc_22172_new_n7161_; 
wire core__abc_22172_new_n7162_; 
wire core__abc_22172_new_n7163_; 
wire core__abc_22172_new_n7164_; 
wire core__abc_22172_new_n7165_; 
wire core__abc_22172_new_n7166_; 
wire core__abc_22172_new_n7167_; 
wire core__abc_22172_new_n7168_; 
wire core__abc_22172_new_n7169_; 
wire core__abc_22172_new_n7170_; 
wire core__abc_22172_new_n7171_; 
wire core__abc_22172_new_n7172_; 
wire core__abc_22172_new_n7174_; 
wire core__abc_22172_new_n7175_; 
wire core__abc_22172_new_n7176_; 
wire core__abc_22172_new_n7177_; 
wire core__abc_22172_new_n7178_; 
wire core__abc_22172_new_n7179_; 
wire core__abc_22172_new_n7180_; 
wire core__abc_22172_new_n7181_; 
wire core__abc_22172_new_n7182_; 
wire core__abc_22172_new_n7183_; 
wire core__abc_22172_new_n7184_; 
wire core__abc_22172_new_n7185_; 
wire core__abc_22172_new_n7186_; 
wire core__abc_22172_new_n7187_; 
wire core__abc_22172_new_n7188_; 
wire core__abc_22172_new_n7189_; 
wire core__abc_22172_new_n7190_; 
wire core__abc_22172_new_n7191_; 
wire core__abc_22172_new_n7192_; 
wire core__abc_22172_new_n7193_; 
wire core__abc_22172_new_n7194_; 
wire core__abc_22172_new_n7195_; 
wire core__abc_22172_new_n7196_; 
wire core__abc_22172_new_n7198_; 
wire core__abc_22172_new_n7199_; 
wire core__abc_22172_new_n7200_; 
wire core__abc_22172_new_n7201_; 
wire core__abc_22172_new_n7202_; 
wire core__abc_22172_new_n7203_; 
wire core__abc_22172_new_n7204_; 
wire core__abc_22172_new_n7205_; 
wire core__abc_22172_new_n7206_; 
wire core__abc_22172_new_n7207_; 
wire core__abc_22172_new_n7208_; 
wire core__abc_22172_new_n7209_; 
wire core__abc_22172_new_n7210_; 
wire core__abc_22172_new_n7211_; 
wire core__abc_22172_new_n7212_; 
wire core__abc_22172_new_n7213_; 
wire core__abc_22172_new_n7214_; 
wire core__abc_22172_new_n7215_; 
wire core__abc_22172_new_n7216_; 
wire core__abc_22172_new_n7217_; 
wire core__abc_22172_new_n7218_; 
wire core__abc_22172_new_n7219_; 
wire core__abc_22172_new_n7220_; 
wire core__abc_22172_new_n7221_; 
wire core__abc_22172_new_n7222_; 
wire core__abc_22172_new_n7223_; 
wire core__abc_22172_new_n7224_; 
wire core__abc_22172_new_n7225_; 
wire core__abc_22172_new_n7226_; 
wire core__abc_22172_new_n7227_; 
wire core__abc_22172_new_n7228_; 
wire core__abc_22172_new_n7229_; 
wire core__abc_22172_new_n7231_; 
wire core__abc_22172_new_n7232_; 
wire core__abc_22172_new_n7233_; 
wire core__abc_22172_new_n7234_; 
wire core__abc_22172_new_n7235_; 
wire core__abc_22172_new_n7236_; 
wire core__abc_22172_new_n7237_; 
wire core__abc_22172_new_n7238_; 
wire core__abc_22172_new_n7239_; 
wire core__abc_22172_new_n7240_; 
wire core__abc_22172_new_n7241_; 
wire core__abc_22172_new_n7242_; 
wire core__abc_22172_new_n7243_; 
wire core__abc_22172_new_n7244_; 
wire core__abc_22172_new_n7245_; 
wire core__abc_22172_new_n7246_; 
wire core__abc_22172_new_n7247_; 
wire core__abc_22172_new_n7248_; 
wire core__abc_22172_new_n7249_; 
wire core__abc_22172_new_n7250_; 
wire core__abc_22172_new_n7251_; 
wire core__abc_22172_new_n7252_; 
wire core__abc_22172_new_n7253_; 
wire core__abc_22172_new_n7254_; 
wire core__abc_22172_new_n7256_; 
wire core__abc_22172_new_n7257_; 
wire core__abc_22172_new_n7258_; 
wire core__abc_22172_new_n7259_; 
wire core__abc_22172_new_n7260_; 
wire core__abc_22172_new_n7261_; 
wire core__abc_22172_new_n7262_; 
wire core__abc_22172_new_n7263_; 
wire core__abc_22172_new_n7264_; 
wire core__abc_22172_new_n7265_; 
wire core__abc_22172_new_n7266_; 
wire core__abc_22172_new_n7267_; 
wire core__abc_22172_new_n7268_; 
wire core__abc_22172_new_n7269_; 
wire core__abc_22172_new_n7270_; 
wire core__abc_22172_new_n7271_; 
wire core__abc_22172_new_n7272_; 
wire core__abc_22172_new_n7273_; 
wire core__abc_22172_new_n7274_; 
wire core__abc_22172_new_n7275_; 
wire core__abc_22172_new_n7276_; 
wire core__abc_22172_new_n7277_; 
wire core__abc_22172_new_n7278_; 
wire core__abc_22172_new_n7279_; 
wire core__abc_22172_new_n7280_; 
wire core__abc_22172_new_n7281_; 
wire core__abc_22172_new_n7282_; 
wire core__abc_22172_new_n7283_; 
wire core__abc_22172_new_n7284_; 
wire core__abc_22172_new_n7285_; 
wire core__abc_22172_new_n7286_; 
wire core__abc_22172_new_n7287_; 
wire core__abc_22172_new_n7289_; 
wire core__abc_22172_new_n7290_; 
wire core__abc_22172_new_n7291_; 
wire core__abc_22172_new_n7292_; 
wire core__abc_22172_new_n7293_; 
wire core__abc_22172_new_n7294_; 
wire core__abc_22172_new_n7295_; 
wire core__abc_22172_new_n7296_; 
wire core__abc_22172_new_n7297_; 
wire core__abc_22172_new_n7298_; 
wire core__abc_22172_new_n7299_; 
wire core__abc_22172_new_n7300_; 
wire core__abc_22172_new_n7301_; 
wire core__abc_22172_new_n7302_; 
wire core__abc_22172_new_n7303_; 
wire core__abc_22172_new_n7304_; 
wire core__abc_22172_new_n7305_; 
wire core__abc_22172_new_n7306_; 
wire core__abc_22172_new_n7307_; 
wire core__abc_22172_new_n7308_; 
wire core__abc_22172_new_n7309_; 
wire core__abc_22172_new_n7310_; 
wire core__abc_22172_new_n7311_; 
wire core__abc_22172_new_n7312_; 
wire core__abc_22172_new_n7313_; 
wire core__abc_22172_new_n7314_; 
wire core__abc_22172_new_n7316_; 
wire core__abc_22172_new_n7317_; 
wire core__abc_22172_new_n7318_; 
wire core__abc_22172_new_n7319_; 
wire core__abc_22172_new_n7320_; 
wire core__abc_22172_new_n7321_; 
wire core__abc_22172_new_n7322_; 
wire core__abc_22172_new_n7323_; 
wire core__abc_22172_new_n7324_; 
wire core__abc_22172_new_n7325_; 
wire core__abc_22172_new_n7326_; 
wire core__abc_22172_new_n7327_; 
wire core__abc_22172_new_n7328_; 
wire core__abc_22172_new_n7329_; 
wire core__abc_22172_new_n7330_; 
wire core__abc_22172_new_n7331_; 
wire core__abc_22172_new_n7332_; 
wire core__abc_22172_new_n7333_; 
wire core__abc_22172_new_n7334_; 
wire core__abc_22172_new_n7335_; 
wire core__abc_22172_new_n7336_; 
wire core__abc_22172_new_n7337_; 
wire core__abc_22172_new_n7338_; 
wire core__abc_22172_new_n7339_; 
wire core__abc_22172_new_n7340_; 
wire core__abc_22172_new_n7341_; 
wire core__abc_22172_new_n7342_; 
wire core__abc_22172_new_n7343_; 
wire core__abc_22172_new_n7344_; 
wire core__abc_22172_new_n7345_; 
wire core__abc_22172_new_n7346_; 
wire core__abc_22172_new_n7347_; 
wire core__abc_22172_new_n7348_; 
wire core__abc_22172_new_n7349_; 
wire core__abc_22172_new_n7350_; 
wire core__abc_22172_new_n7351_; 
wire core__abc_22172_new_n7352_; 
wire core__abc_22172_new_n7353_; 
wire core__abc_22172_new_n7354_; 
wire core__abc_22172_new_n7355_; 
wire core__abc_22172_new_n7356_; 
wire core__abc_22172_new_n7357_; 
wire core__abc_22172_new_n7358_; 
wire core__abc_22172_new_n7359_; 
wire core__abc_22172_new_n7361_; 
wire core__abc_22172_new_n7362_; 
wire core__abc_22172_new_n7363_; 
wire core__abc_22172_new_n7364_; 
wire core__abc_22172_new_n7365_; 
wire core__abc_22172_new_n7366_; 
wire core__abc_22172_new_n7367_; 
wire core__abc_22172_new_n7368_; 
wire core__abc_22172_new_n7369_; 
wire core__abc_22172_new_n7370_; 
wire core__abc_22172_new_n7371_; 
wire core__abc_22172_new_n7372_; 
wire core__abc_22172_new_n7373_; 
wire core__abc_22172_new_n7374_; 
wire core__abc_22172_new_n7375_; 
wire core__abc_22172_new_n7376_; 
wire core__abc_22172_new_n7377_; 
wire core__abc_22172_new_n7378_; 
wire core__abc_22172_new_n7379_; 
wire core__abc_22172_new_n7380_; 
wire core__abc_22172_new_n7381_; 
wire core__abc_22172_new_n7382_; 
wire core__abc_22172_new_n7383_; 
wire core__abc_22172_new_n7384_; 
wire core__abc_22172_new_n7385_; 
wire core__abc_22172_new_n7386_; 
wire core__abc_22172_new_n7387_; 
wire core__abc_22172_new_n7388_; 
wire core__abc_22172_new_n7390_; 
wire core__abc_22172_new_n7391_; 
wire core__abc_22172_new_n7392_; 
wire core__abc_22172_new_n7393_; 
wire core__abc_22172_new_n7394_; 
wire core__abc_22172_new_n7395_; 
wire core__abc_22172_new_n7396_; 
wire core__abc_22172_new_n7397_; 
wire core__abc_22172_new_n7398_; 
wire core__abc_22172_new_n7399_; 
wire core__abc_22172_new_n7400_; 
wire core__abc_22172_new_n7401_; 
wire core__abc_22172_new_n7402_; 
wire core__abc_22172_new_n7403_; 
wire core__abc_22172_new_n7404_; 
wire core__abc_22172_new_n7405_; 
wire core__abc_22172_new_n7406_; 
wire core__abc_22172_new_n7407_; 
wire core__abc_22172_new_n7408_; 
wire core__abc_22172_new_n7409_; 
wire core__abc_22172_new_n7410_; 
wire core__abc_22172_new_n7411_; 
wire core__abc_22172_new_n7412_; 
wire core__abc_22172_new_n7413_; 
wire core__abc_22172_new_n7414_; 
wire core__abc_22172_new_n7415_; 
wire core__abc_22172_new_n7417_; 
wire core__abc_22172_new_n7418_; 
wire core__abc_22172_new_n7419_; 
wire core__abc_22172_new_n7420_; 
wire core__abc_22172_new_n7421_; 
wire core__abc_22172_new_n7422_; 
wire core__abc_22172_new_n7423_; 
wire core__abc_22172_new_n7424_; 
wire core__abc_22172_new_n7425_; 
wire core__abc_22172_new_n7426_; 
wire core__abc_22172_new_n7427_; 
wire core__abc_22172_new_n7428_; 
wire core__abc_22172_new_n7429_; 
wire core__abc_22172_new_n7430_; 
wire core__abc_22172_new_n7431_; 
wire core__abc_22172_new_n7432_; 
wire core__abc_22172_new_n7433_; 
wire core__abc_22172_new_n7434_; 
wire core__abc_22172_new_n7435_; 
wire core__abc_22172_new_n7436_; 
wire core__abc_22172_new_n7437_; 
wire core__abc_22172_new_n7438_; 
wire core__abc_22172_new_n7439_; 
wire core__abc_22172_new_n7440_; 
wire core__abc_22172_new_n7441_; 
wire core__abc_22172_new_n7443_; 
wire core__abc_22172_new_n7444_; 
wire core__abc_22172_new_n7445_; 
wire core__abc_22172_new_n7446_; 
wire core__abc_22172_new_n7447_; 
wire core__abc_22172_new_n7448_; 
wire core__abc_22172_new_n7449_; 
wire core__abc_22172_new_n7450_; 
wire core__abc_22172_new_n7451_; 
wire core__abc_22172_new_n7452_; 
wire core__abc_22172_new_n7453_; 
wire core__abc_22172_new_n7454_; 
wire core__abc_22172_new_n7455_; 
wire core__abc_22172_new_n7456_; 
wire core__abc_22172_new_n7457_; 
wire core__abc_22172_new_n7458_; 
wire core__abc_22172_new_n7459_; 
wire core__abc_22172_new_n7460_; 
wire core__abc_22172_new_n7461_; 
wire core__abc_22172_new_n7462_; 
wire core__abc_22172_new_n7463_; 
wire core__abc_22172_new_n7464_; 
wire core__abc_22172_new_n7465_; 
wire core__abc_22172_new_n7466_; 
wire core__abc_22172_new_n7467_; 
wire core__abc_22172_new_n7468_; 
wire core__abc_22172_new_n7469_; 
wire core__abc_22172_new_n7470_; 
wire core__abc_22172_new_n7471_; 
wire core__abc_22172_new_n7472_; 
wire core__abc_22172_new_n7473_; 
wire core__abc_22172_new_n7474_; 
wire core__abc_22172_new_n7475_; 
wire core__abc_22172_new_n7476_; 
wire core__abc_22172_new_n7478_; 
wire core__abc_22172_new_n7479_; 
wire core__abc_22172_new_n7480_; 
wire core__abc_22172_new_n7481_; 
wire core__abc_22172_new_n7482_; 
wire core__abc_22172_new_n7483_; 
wire core__abc_22172_new_n7484_; 
wire core__abc_22172_new_n7485_; 
wire core__abc_22172_new_n7486_; 
wire core__abc_22172_new_n7487_; 
wire core__abc_22172_new_n7488_; 
wire core__abc_22172_new_n7489_; 
wire core__abc_22172_new_n7490_; 
wire core__abc_22172_new_n7491_; 
wire core__abc_22172_new_n7492_; 
wire core__abc_22172_new_n7493_; 
wire core__abc_22172_new_n7494_; 
wire core__abc_22172_new_n7495_; 
wire core__abc_22172_new_n7496_; 
wire core__abc_22172_new_n7497_; 
wire core__abc_22172_new_n7498_; 
wire core__abc_22172_new_n7499_; 
wire core__abc_22172_new_n7500_; 
wire core__abc_22172_new_n7501_; 
wire core__abc_22172_new_n7502_; 
wire core__abc_22172_new_n7503_; 
wire core__abc_22172_new_n7504_; 
wire core__abc_22172_new_n7506_; 
wire core__abc_22172_new_n7507_; 
wire core__abc_22172_new_n7508_; 
wire core__abc_22172_new_n7509_; 
wire core__abc_22172_new_n7510_; 
wire core__abc_22172_new_n7511_; 
wire core__abc_22172_new_n7512_; 
wire core__abc_22172_new_n7513_; 
wire core__abc_22172_new_n7514_; 
wire core__abc_22172_new_n7515_; 
wire core__abc_22172_new_n7516_; 
wire core__abc_22172_new_n7517_; 
wire core__abc_22172_new_n7518_; 
wire core__abc_22172_new_n7519_; 
wire core__abc_22172_new_n7520_; 
wire core__abc_22172_new_n7521_; 
wire core__abc_22172_new_n7522_; 
wire core__abc_22172_new_n7523_; 
wire core__abc_22172_new_n7524_; 
wire core__abc_22172_new_n7525_; 
wire core__abc_22172_new_n7526_; 
wire core__abc_22172_new_n7527_; 
wire core__abc_22172_new_n7528_; 
wire core__abc_22172_new_n7529_; 
wire core__abc_22172_new_n7530_; 
wire core__abc_22172_new_n7531_; 
wire core__abc_22172_new_n7532_; 
wire core__abc_22172_new_n7533_; 
wire core__abc_22172_new_n7535_; 
wire core__abc_22172_new_n7536_; 
wire core__abc_22172_new_n7537_; 
wire core__abc_22172_new_n7538_; 
wire core__abc_22172_new_n7539_; 
wire core__abc_22172_new_n7540_; 
wire core__abc_22172_new_n7541_; 
wire core__abc_22172_new_n7542_; 
wire core__abc_22172_new_n7543_; 
wire core__abc_22172_new_n7544_; 
wire core__abc_22172_new_n7545_; 
wire core__abc_22172_new_n7546_; 
wire core__abc_22172_new_n7547_; 
wire core__abc_22172_new_n7548_; 
wire core__abc_22172_new_n7549_; 
wire core__abc_22172_new_n7550_; 
wire core__abc_22172_new_n7551_; 
wire core__abc_22172_new_n7552_; 
wire core__abc_22172_new_n7553_; 
wire core__abc_22172_new_n7554_; 
wire core__abc_22172_new_n7555_; 
wire core__abc_22172_new_n7556_; 
wire core__abc_22172_new_n7557_; 
wire core__abc_22172_new_n7558_; 
wire core__abc_22172_new_n7559_; 
wire core__abc_22172_new_n7560_; 
wire core__abc_22172_new_n7561_; 
wire core__abc_22172_new_n7563_; 
wire core__abc_22172_new_n7564_; 
wire core__abc_22172_new_n7565_; 
wire core__abc_22172_new_n7566_; 
wire core__abc_22172_new_n7567_; 
wire core__abc_22172_new_n7568_; 
wire core__abc_22172_new_n7569_; 
wire core__abc_22172_new_n7570_; 
wire core__abc_22172_new_n7571_; 
wire core__abc_22172_new_n7572_; 
wire core__abc_22172_new_n7573_; 
wire core__abc_22172_new_n7574_; 
wire core__abc_22172_new_n7575_; 
wire core__abc_22172_new_n7576_; 
wire core__abc_22172_new_n7577_; 
wire core__abc_22172_new_n7578_; 
wire core__abc_22172_new_n7579_; 
wire core__abc_22172_new_n7580_; 
wire core__abc_22172_new_n7581_; 
wire core__abc_22172_new_n7582_; 
wire core__abc_22172_new_n7583_; 
wire core__abc_22172_new_n7584_; 
wire core__abc_22172_new_n7585_; 
wire core__abc_22172_new_n7586_; 
wire core__abc_22172_new_n7587_; 
wire core__abc_22172_new_n7588_; 
wire core__abc_22172_new_n7589_; 
wire core__abc_22172_new_n7590_; 
wire core__abc_22172_new_n7591_; 
wire core__abc_22172_new_n7592_; 
wire core__abc_22172_new_n7593_; 
wire core__abc_22172_new_n7594_; 
wire core__abc_22172_new_n7595_; 
wire core__abc_22172_new_n7596_; 
wire core__abc_22172_new_n7597_; 
wire core__abc_22172_new_n7598_; 
wire core__abc_22172_new_n7599_; 
wire core__abc_22172_new_n7601_; 
wire core__abc_22172_new_n7602_; 
wire core__abc_22172_new_n7603_; 
wire core__abc_22172_new_n7604_; 
wire core__abc_22172_new_n7605_; 
wire core__abc_22172_new_n7606_; 
wire core__abc_22172_new_n7607_; 
wire core__abc_22172_new_n7608_; 
wire core__abc_22172_new_n7609_; 
wire core__abc_22172_new_n7610_; 
wire core__abc_22172_new_n7611_; 
wire core__abc_22172_new_n7612_; 
wire core__abc_22172_new_n7613_; 
wire core__abc_22172_new_n7614_; 
wire core__abc_22172_new_n7615_; 
wire core__abc_22172_new_n7616_; 
wire core__abc_22172_new_n7617_; 
wire core__abc_22172_new_n7618_; 
wire core__abc_22172_new_n7619_; 
wire core__abc_22172_new_n7620_; 
wire core__abc_22172_new_n7621_; 
wire core__abc_22172_new_n7622_; 
wire core__abc_22172_new_n7623_; 
wire core__abc_22172_new_n7624_; 
wire core__abc_22172_new_n7625_; 
wire core__abc_22172_new_n7627_; 
wire core__abc_22172_new_n7628_; 
wire core__abc_22172_new_n7629_; 
wire core__abc_22172_new_n7630_; 
wire core__abc_22172_new_n7631_; 
wire core__abc_22172_new_n7632_; 
wire core__abc_22172_new_n7633_; 
wire core__abc_22172_new_n7634_; 
wire core__abc_22172_new_n7635_; 
wire core__abc_22172_new_n7636_; 
wire core__abc_22172_new_n7637_; 
wire core__abc_22172_new_n7638_; 
wire core__abc_22172_new_n7639_; 
wire core__abc_22172_new_n7640_; 
wire core__abc_22172_new_n7641_; 
wire core__abc_22172_new_n7642_; 
wire core__abc_22172_new_n7643_; 
wire core__abc_22172_new_n7644_; 
wire core__abc_22172_new_n7645_; 
wire core__abc_22172_new_n7646_; 
wire core__abc_22172_new_n7647_; 
wire core__abc_22172_new_n7648_; 
wire core__abc_22172_new_n7649_; 
wire core__abc_22172_new_n7650_; 
wire core__abc_22172_new_n7651_; 
wire core__abc_22172_new_n7652_; 
wire core__abc_22172_new_n7653_; 
wire core__abc_22172_new_n7654_; 
wire core__abc_22172_new_n7655_; 
wire core__abc_22172_new_n7657_; 
wire core__abc_22172_new_n7658_; 
wire core__abc_22172_new_n7659_; 
wire core__abc_22172_new_n7660_; 
wire core__abc_22172_new_n7661_; 
wire core__abc_22172_new_n7662_; 
wire core__abc_22172_new_n7663_; 
wire core__abc_22172_new_n7664_; 
wire core__abc_22172_new_n7665_; 
wire core__abc_22172_new_n7666_; 
wire core__abc_22172_new_n7667_; 
wire core__abc_22172_new_n7668_; 
wire core__abc_22172_new_n7669_; 
wire core__abc_22172_new_n7670_; 
wire core__abc_22172_new_n7671_; 
wire core__abc_22172_new_n7672_; 
wire core__abc_22172_new_n7673_; 
wire core__abc_22172_new_n7674_; 
wire core__abc_22172_new_n7675_; 
wire core__abc_22172_new_n7676_; 
wire core__abc_22172_new_n7677_; 
wire core__abc_22172_new_n7678_; 
wire core__abc_22172_new_n7679_; 
wire core__abc_22172_new_n7680_; 
wire core__abc_22172_new_n7682_; 
wire core__abc_22172_new_n7683_; 
wire core__abc_22172_new_n7684_; 
wire core__abc_22172_new_n7685_; 
wire core__abc_22172_new_n7686_; 
wire core__abc_22172_new_n7687_; 
wire core__abc_22172_new_n7688_; 
wire core__abc_22172_new_n7689_; 
wire core__abc_22172_new_n7690_; 
wire core__abc_22172_new_n7691_; 
wire core__abc_22172_new_n7692_; 
wire core__abc_22172_new_n7693_; 
wire core__abc_22172_new_n7694_; 
wire core__abc_22172_new_n7695_; 
wire core__abc_22172_new_n7696_; 
wire core__abc_22172_new_n7697_; 
wire core__abc_22172_new_n7698_; 
wire core__abc_22172_new_n7699_; 
wire core__abc_22172_new_n7700_; 
wire core__abc_22172_new_n7701_; 
wire core__abc_22172_new_n7702_; 
wire core__abc_22172_new_n7703_; 
wire core__abc_22172_new_n7704_; 
wire core__abc_22172_new_n7705_; 
wire core__abc_22172_new_n7706_; 
wire core__abc_22172_new_n7707_; 
wire core__abc_22172_new_n7708_; 
wire core__abc_22172_new_n7709_; 
wire core__abc_22172_new_n7710_; 
wire core__abc_22172_new_n7711_; 
wire core__abc_22172_new_n7713_; 
wire core__abc_22172_new_n7714_; 
wire core__abc_22172_new_n7715_; 
wire core__abc_22172_new_n7716_; 
wire core__abc_22172_new_n7717_; 
wire core__abc_22172_new_n7718_; 
wire core__abc_22172_new_n7719_; 
wire core__abc_22172_new_n7720_; 
wire core__abc_22172_new_n7721_; 
wire core__abc_22172_new_n7722_; 
wire core__abc_22172_new_n7723_; 
wire core__abc_22172_new_n7724_; 
wire core__abc_22172_new_n7725_; 
wire core__abc_22172_new_n7726_; 
wire core__abc_22172_new_n7727_; 
wire core__abc_22172_new_n7728_; 
wire core__abc_22172_new_n7729_; 
wire core__abc_22172_new_n7730_; 
wire core__abc_22172_new_n7731_; 
wire core__abc_22172_new_n7732_; 
wire core__abc_22172_new_n7733_; 
wire core__abc_22172_new_n7734_; 
wire core__abc_22172_new_n7735_; 
wire core__abc_22172_new_n7736_; 
wire core__abc_22172_new_n7738_; 
wire core__abc_22172_new_n7739_; 
wire core__abc_22172_new_n7740_; 
wire core__abc_22172_new_n7741_; 
wire core__abc_22172_new_n7742_; 
wire core__abc_22172_new_n7743_; 
wire core__abc_22172_new_n7744_; 
wire core__abc_22172_new_n7745_; 
wire core__abc_22172_new_n7746_; 
wire core__abc_22172_new_n7747_; 
wire core__abc_22172_new_n7748_; 
wire core__abc_22172_new_n7749_; 
wire core__abc_22172_new_n7750_; 
wire core__abc_22172_new_n7751_; 
wire core__abc_22172_new_n7752_; 
wire core__abc_22172_new_n7753_; 
wire core__abc_22172_new_n7754_; 
wire core__abc_22172_new_n7755_; 
wire core__abc_22172_new_n7756_; 
wire core__abc_22172_new_n7757_; 
wire core__abc_22172_new_n7758_; 
wire core__abc_22172_new_n7759_; 
wire core__abc_22172_new_n7760_; 
wire core__abc_22172_new_n7761_; 
wire core__abc_22172_new_n7762_; 
wire core__abc_22172_new_n7763_; 
wire core__abc_22172_new_n7764_; 
wire core__abc_22172_new_n7765_; 
wire core__abc_22172_new_n7767_; 
wire core__abc_22172_new_n7768_; 
wire core__abc_22172_new_n7769_; 
wire core__abc_22172_new_n7770_; 
wire core__abc_22172_new_n7771_; 
wire core__abc_22172_new_n7772_; 
wire core__abc_22172_new_n7773_; 
wire core__abc_22172_new_n7774_; 
wire core__abc_22172_new_n7775_; 
wire core__abc_22172_new_n7776_; 
wire core__abc_22172_new_n7777_; 
wire core__abc_22172_new_n7778_; 
wire core__abc_22172_new_n7779_; 
wire core__abc_22172_new_n7780_; 
wire core__abc_22172_new_n7781_; 
wire core__abc_22172_new_n7782_; 
wire core__abc_22172_new_n7783_; 
wire core__abc_22172_new_n7784_; 
wire core__abc_22172_new_n7785_; 
wire core__abc_22172_new_n7786_; 
wire core__abc_22172_new_n7787_; 
wire core__abc_22172_new_n7788_; 
wire core__abc_22172_new_n7790_; 
wire core__abc_22172_new_n7791_; 
wire core__abc_22172_new_n7792_; 
wire core__abc_22172_new_n7793_; 
wire core__abc_22172_new_n7794_; 
wire core__abc_22172_new_n7795_; 
wire core__abc_22172_new_n7796_; 
wire core__abc_22172_new_n7797_; 
wire core__abc_22172_new_n7798_; 
wire core__abc_22172_new_n7799_; 
wire core__abc_22172_new_n7800_; 
wire core__abc_22172_new_n7802_; 
wire core__abc_22172_new_n7803_; 
wire core__abc_22172_new_n7804_; 
wire core__abc_22172_new_n7805_; 
wire core__abc_22172_new_n7806_; 
wire core__abc_22172_new_n7807_; 
wire core__abc_22172_new_n7808_; 
wire core__abc_22172_new_n7809_; 
wire core__abc_22172_new_n7810_; 
wire core__abc_22172_new_n7812_; 
wire core__abc_22172_new_n7813_; 
wire core__abc_22172_new_n7814_; 
wire core__abc_22172_new_n7815_; 
wire core__abc_22172_new_n7816_; 
wire core__abc_22172_new_n7817_; 
wire core__abc_22172_new_n7818_; 
wire core__abc_22172_new_n7819_; 
wire core__abc_22172_new_n7820_; 
wire core__abc_22172_new_n7821_; 
wire core__abc_22172_new_n7822_; 
wire core__abc_22172_new_n7823_; 
wire core__abc_22172_new_n7825_; 
wire core__abc_22172_new_n7826_; 
wire core__abc_22172_new_n7827_; 
wire core__abc_22172_new_n7828_; 
wire core__abc_22172_new_n7829_; 
wire core__abc_22172_new_n7830_; 
wire core__abc_22172_new_n7831_; 
wire core__abc_22172_new_n7832_; 
wire core__abc_22172_new_n7833_; 
wire core__abc_22172_new_n7834_; 
wire core__abc_22172_new_n7835_; 
wire core__abc_22172_new_n7836_; 
wire core__abc_22172_new_n7837_; 
wire core__abc_22172_new_n7838_; 
wire core__abc_22172_new_n7839_; 
wire core__abc_22172_new_n7840_; 
wire core__abc_22172_new_n7842_; 
wire core__abc_22172_new_n7843_; 
wire core__abc_22172_new_n7844_; 
wire core__abc_22172_new_n7845_; 
wire core__abc_22172_new_n7846_; 
wire core__abc_22172_new_n7847_; 
wire core__abc_22172_new_n7848_; 
wire core__abc_22172_new_n7849_; 
wire core__abc_22172_new_n7850_; 
wire core__abc_22172_new_n7851_; 
wire core__abc_22172_new_n7852_; 
wire core__abc_22172_new_n7854_; 
wire core__abc_22172_new_n7855_; 
wire core__abc_22172_new_n7856_; 
wire core__abc_22172_new_n7857_; 
wire core__abc_22172_new_n7858_; 
wire core__abc_22172_new_n7859_; 
wire core__abc_22172_new_n7860_; 
wire core__abc_22172_new_n7861_; 
wire core__abc_22172_new_n7862_; 
wire core__abc_22172_new_n7863_; 
wire core__abc_22172_new_n7864_; 
wire core__abc_22172_new_n7865_; 
wire core__abc_22172_new_n7866_; 
wire core__abc_22172_new_n7867_; 
wire core__abc_22172_new_n7868_; 
wire core__abc_22172_new_n7869_; 
wire core__abc_22172_new_n7870_; 
wire core__abc_22172_new_n7872_; 
wire core__abc_22172_new_n7873_; 
wire core__abc_22172_new_n7874_; 
wire core__abc_22172_new_n7875_; 
wire core__abc_22172_new_n7876_; 
wire core__abc_22172_new_n7877_; 
wire core__abc_22172_new_n7878_; 
wire core__abc_22172_new_n7879_; 
wire core__abc_22172_new_n7880_; 
wire core__abc_22172_new_n7881_; 
wire core__abc_22172_new_n7882_; 
wire core__abc_22172_new_n7883_; 
wire core__abc_22172_new_n7884_; 
wire core__abc_22172_new_n7886_; 
wire core__abc_22172_new_n7887_; 
wire core__abc_22172_new_n7888_; 
wire core__abc_22172_new_n7889_; 
wire core__abc_22172_new_n7890_; 
wire core__abc_22172_new_n7891_; 
wire core__abc_22172_new_n7892_; 
wire core__abc_22172_new_n7893_; 
wire core__abc_22172_new_n7894_; 
wire core__abc_22172_new_n7895_; 
wire core__abc_22172_new_n7896_; 
wire core__abc_22172_new_n7897_; 
wire core__abc_22172_new_n7898_; 
wire core__abc_22172_new_n7899_; 
wire core__abc_22172_new_n7901_; 
wire core__abc_22172_new_n7902_; 
wire core__abc_22172_new_n7903_; 
wire core__abc_22172_new_n7904_; 
wire core__abc_22172_new_n7905_; 
wire core__abc_22172_new_n7906_; 
wire core__abc_22172_new_n7907_; 
wire core__abc_22172_new_n7908_; 
wire core__abc_22172_new_n7909_; 
wire core__abc_22172_new_n7910_; 
wire core__abc_22172_new_n7911_; 
wire core__abc_22172_new_n7912_; 
wire core__abc_22172_new_n7913_; 
wire core__abc_22172_new_n7915_; 
wire core__abc_22172_new_n7916_; 
wire core__abc_22172_new_n7917_; 
wire core__abc_22172_new_n7918_; 
wire core__abc_22172_new_n7919_; 
wire core__abc_22172_new_n7920_; 
wire core__abc_22172_new_n7921_; 
wire core__abc_22172_new_n7922_; 
wire core__abc_22172_new_n7923_; 
wire core__abc_22172_new_n7924_; 
wire core__abc_22172_new_n7925_; 
wire core__abc_22172_new_n7926_; 
wire core__abc_22172_new_n7927_; 
wire core__abc_22172_new_n7928_; 
wire core__abc_22172_new_n7929_; 
wire core__abc_22172_new_n7930_; 
wire core__abc_22172_new_n7932_; 
wire core__abc_22172_new_n7933_; 
wire core__abc_22172_new_n7934_; 
wire core__abc_22172_new_n7935_; 
wire core__abc_22172_new_n7936_; 
wire core__abc_22172_new_n7937_; 
wire core__abc_22172_new_n7938_; 
wire core__abc_22172_new_n7939_; 
wire core__abc_22172_new_n7940_; 
wire core__abc_22172_new_n7941_; 
wire core__abc_22172_new_n7942_; 
wire core__abc_22172_new_n7943_; 
wire core__abc_22172_new_n7944_; 
wire core__abc_22172_new_n7945_; 
wire core__abc_22172_new_n7946_; 
wire core__abc_22172_new_n7948_; 
wire core__abc_22172_new_n7949_; 
wire core__abc_22172_new_n7950_; 
wire core__abc_22172_new_n7951_; 
wire core__abc_22172_new_n7952_; 
wire core__abc_22172_new_n7953_; 
wire core__abc_22172_new_n7954_; 
wire core__abc_22172_new_n7955_; 
wire core__abc_22172_new_n7956_; 
wire core__abc_22172_new_n7957_; 
wire core__abc_22172_new_n7958_; 
wire core__abc_22172_new_n7959_; 
wire core__abc_22172_new_n7960_; 
wire core__abc_22172_new_n7961_; 
wire core__abc_22172_new_n7962_; 
wire core__abc_22172_new_n7964_; 
wire core__abc_22172_new_n7965_; 
wire core__abc_22172_new_n7966_; 
wire core__abc_22172_new_n7967_; 
wire core__abc_22172_new_n7968_; 
wire core__abc_22172_new_n7969_; 
wire core__abc_22172_new_n7970_; 
wire core__abc_22172_new_n7971_; 
wire core__abc_22172_new_n7972_; 
wire core__abc_22172_new_n7973_; 
wire core__abc_22172_new_n7974_; 
wire core__abc_22172_new_n7975_; 
wire core__abc_22172_new_n7977_; 
wire core__abc_22172_new_n7978_; 
wire core__abc_22172_new_n7979_; 
wire core__abc_22172_new_n7980_; 
wire core__abc_22172_new_n7981_; 
wire core__abc_22172_new_n7982_; 
wire core__abc_22172_new_n7983_; 
wire core__abc_22172_new_n7984_; 
wire core__abc_22172_new_n7985_; 
wire core__abc_22172_new_n7986_; 
wire core__abc_22172_new_n7987_; 
wire core__abc_22172_new_n7988_; 
wire core__abc_22172_new_n7989_; 
wire core__abc_22172_new_n7990_; 
wire core__abc_22172_new_n7991_; 
wire core__abc_22172_new_n7993_; 
wire core__abc_22172_new_n7994_; 
wire core__abc_22172_new_n7995_; 
wire core__abc_22172_new_n7996_; 
wire core__abc_22172_new_n7997_; 
wire core__abc_22172_new_n7998_; 
wire core__abc_22172_new_n7999_; 
wire core__abc_22172_new_n8000_; 
wire core__abc_22172_new_n8001_; 
wire core__abc_22172_new_n8002_; 
wire core__abc_22172_new_n8003_; 
wire core__abc_22172_new_n8004_; 
wire core__abc_22172_new_n8005_; 
wire core__abc_22172_new_n8006_; 
wire core__abc_22172_new_n8007_; 
wire core__abc_22172_new_n8008_; 
wire core__abc_22172_new_n8010_; 
wire core__abc_22172_new_n8011_; 
wire core__abc_22172_new_n8012_; 
wire core__abc_22172_new_n8013_; 
wire core__abc_22172_new_n8014_; 
wire core__abc_22172_new_n8015_; 
wire core__abc_22172_new_n8016_; 
wire core__abc_22172_new_n8017_; 
wire core__abc_22172_new_n8018_; 
wire core__abc_22172_new_n8019_; 
wire core__abc_22172_new_n8020_; 
wire core__abc_22172_new_n8021_; 
wire core__abc_22172_new_n8022_; 
wire core__abc_22172_new_n8023_; 
wire core__abc_22172_new_n8024_; 
wire core__abc_22172_new_n8026_; 
wire core__abc_22172_new_n8027_; 
wire core__abc_22172_new_n8028_; 
wire core__abc_22172_new_n8029_; 
wire core__abc_22172_new_n8030_; 
wire core__abc_22172_new_n8031_; 
wire core__abc_22172_new_n8032_; 
wire core__abc_22172_new_n8033_; 
wire core__abc_22172_new_n8034_; 
wire core__abc_22172_new_n8035_; 
wire core__abc_22172_new_n8036_; 
wire core__abc_22172_new_n8037_; 
wire core__abc_22172_new_n8038_; 
wire core__abc_22172_new_n8039_; 
wire core__abc_22172_new_n8041_; 
wire core__abc_22172_new_n8042_; 
wire core__abc_22172_new_n8043_; 
wire core__abc_22172_new_n8044_; 
wire core__abc_22172_new_n8045_; 
wire core__abc_22172_new_n8046_; 
wire core__abc_22172_new_n8047_; 
wire core__abc_22172_new_n8048_; 
wire core__abc_22172_new_n8049_; 
wire core__abc_22172_new_n8050_; 
wire core__abc_22172_new_n8051_; 
wire core__abc_22172_new_n8052_; 
wire core__abc_22172_new_n8053_; 
wire core__abc_22172_new_n8054_; 
wire core__abc_22172_new_n8056_; 
wire core__abc_22172_new_n8057_; 
wire core__abc_22172_new_n8058_; 
wire core__abc_22172_new_n8059_; 
wire core__abc_22172_new_n8060_; 
wire core__abc_22172_new_n8061_; 
wire core__abc_22172_new_n8062_; 
wire core__abc_22172_new_n8063_; 
wire core__abc_22172_new_n8064_; 
wire core__abc_22172_new_n8065_; 
wire core__abc_22172_new_n8066_; 
wire core__abc_22172_new_n8067_; 
wire core__abc_22172_new_n8068_; 
wire core__abc_22172_new_n8069_; 
wire core__abc_22172_new_n8071_; 
wire core__abc_22172_new_n8072_; 
wire core__abc_22172_new_n8073_; 
wire core__abc_22172_new_n8074_; 
wire core__abc_22172_new_n8075_; 
wire core__abc_22172_new_n8076_; 
wire core__abc_22172_new_n8077_; 
wire core__abc_22172_new_n8078_; 
wire core__abc_22172_new_n8079_; 
wire core__abc_22172_new_n8080_; 
wire core__abc_22172_new_n8081_; 
wire core__abc_22172_new_n8082_; 
wire core__abc_22172_new_n8083_; 
wire core__abc_22172_new_n8084_; 
wire core__abc_22172_new_n8085_; 
wire core__abc_22172_new_n8087_; 
wire core__abc_22172_new_n8088_; 
wire core__abc_22172_new_n8089_; 
wire core__abc_22172_new_n8090_; 
wire core__abc_22172_new_n8091_; 
wire core__abc_22172_new_n8092_; 
wire core__abc_22172_new_n8093_; 
wire core__abc_22172_new_n8094_; 
wire core__abc_22172_new_n8095_; 
wire core__abc_22172_new_n8096_; 
wire core__abc_22172_new_n8097_; 
wire core__abc_22172_new_n8098_; 
wire core__abc_22172_new_n8099_; 
wire core__abc_22172_new_n8100_; 
wire core__abc_22172_new_n8101_; 
wire core__abc_22172_new_n8102_; 
wire core__abc_22172_new_n8103_; 
wire core__abc_22172_new_n8105_; 
wire core__abc_22172_new_n8106_; 
wire core__abc_22172_new_n8107_; 
wire core__abc_22172_new_n8108_; 
wire core__abc_22172_new_n8109_; 
wire core__abc_22172_new_n8110_; 
wire core__abc_22172_new_n8111_; 
wire core__abc_22172_new_n8112_; 
wire core__abc_22172_new_n8113_; 
wire core__abc_22172_new_n8114_; 
wire core__abc_22172_new_n8115_; 
wire core__abc_22172_new_n8116_; 
wire core__abc_22172_new_n8117_; 
wire core__abc_22172_new_n8118_; 
wire core__abc_22172_new_n8119_; 
wire core__abc_22172_new_n8120_; 
wire core__abc_22172_new_n8122_; 
wire core__abc_22172_new_n8123_; 
wire core__abc_22172_new_n8124_; 
wire core__abc_22172_new_n8125_; 
wire core__abc_22172_new_n8126_; 
wire core__abc_22172_new_n8127_; 
wire core__abc_22172_new_n8128_; 
wire core__abc_22172_new_n8129_; 
wire core__abc_22172_new_n8130_; 
wire core__abc_22172_new_n8131_; 
wire core__abc_22172_new_n8132_; 
wire core__abc_22172_new_n8133_; 
wire core__abc_22172_new_n8134_; 
wire core__abc_22172_new_n8135_; 
wire core__abc_22172_new_n8136_; 
wire core__abc_22172_new_n8138_; 
wire core__abc_22172_new_n8139_; 
wire core__abc_22172_new_n8140_; 
wire core__abc_22172_new_n8141_; 
wire core__abc_22172_new_n8142_; 
wire core__abc_22172_new_n8143_; 
wire core__abc_22172_new_n8144_; 
wire core__abc_22172_new_n8145_; 
wire core__abc_22172_new_n8146_; 
wire core__abc_22172_new_n8147_; 
wire core__abc_22172_new_n8148_; 
wire core__abc_22172_new_n8149_; 
wire core__abc_22172_new_n8150_; 
wire core__abc_22172_new_n8151_; 
wire core__abc_22172_new_n8152_; 
wire core__abc_22172_new_n8154_; 
wire core__abc_22172_new_n8155_; 
wire core__abc_22172_new_n8156_; 
wire core__abc_22172_new_n8157_; 
wire core__abc_22172_new_n8158_; 
wire core__abc_22172_new_n8159_; 
wire core__abc_22172_new_n8160_; 
wire core__abc_22172_new_n8161_; 
wire core__abc_22172_new_n8162_; 
wire core__abc_22172_new_n8163_; 
wire core__abc_22172_new_n8164_; 
wire core__abc_22172_new_n8165_; 
wire core__abc_22172_new_n8166_; 
wire core__abc_22172_new_n8168_; 
wire core__abc_22172_new_n8169_; 
wire core__abc_22172_new_n8170_; 
wire core__abc_22172_new_n8171_; 
wire core__abc_22172_new_n8172_; 
wire core__abc_22172_new_n8173_; 
wire core__abc_22172_new_n8174_; 
wire core__abc_22172_new_n8175_; 
wire core__abc_22172_new_n8176_; 
wire core__abc_22172_new_n8177_; 
wire core__abc_22172_new_n8178_; 
wire core__abc_22172_new_n8179_; 
wire core__abc_22172_new_n8180_; 
wire core__abc_22172_new_n8181_; 
wire core__abc_22172_new_n8182_; 
wire core__abc_22172_new_n8184_; 
wire core__abc_22172_new_n8185_; 
wire core__abc_22172_new_n8186_; 
wire core__abc_22172_new_n8187_; 
wire core__abc_22172_new_n8188_; 
wire core__abc_22172_new_n8189_; 
wire core__abc_22172_new_n8190_; 
wire core__abc_22172_new_n8191_; 
wire core__abc_22172_new_n8192_; 
wire core__abc_22172_new_n8193_; 
wire core__abc_22172_new_n8194_; 
wire core__abc_22172_new_n8195_; 
wire core__abc_22172_new_n8196_; 
wire core__abc_22172_new_n8197_; 
wire core__abc_22172_new_n8198_; 
wire core__abc_22172_new_n8200_; 
wire core__abc_22172_new_n8201_; 
wire core__abc_22172_new_n8202_; 
wire core__abc_22172_new_n8203_; 
wire core__abc_22172_new_n8204_; 
wire core__abc_22172_new_n8205_; 
wire core__abc_22172_new_n8206_; 
wire core__abc_22172_new_n8207_; 
wire core__abc_22172_new_n8208_; 
wire core__abc_22172_new_n8209_; 
wire core__abc_22172_new_n8210_; 
wire core__abc_22172_new_n8211_; 
wire core__abc_22172_new_n8212_; 
wire core__abc_22172_new_n8213_; 
wire core__abc_22172_new_n8214_; 
wire core__abc_22172_new_n8216_; 
wire core__abc_22172_new_n8217_; 
wire core__abc_22172_new_n8218_; 
wire core__abc_22172_new_n8219_; 
wire core__abc_22172_new_n8220_; 
wire core__abc_22172_new_n8221_; 
wire core__abc_22172_new_n8222_; 
wire core__abc_22172_new_n8223_; 
wire core__abc_22172_new_n8224_; 
wire core__abc_22172_new_n8225_; 
wire core__abc_22172_new_n8226_; 
wire core__abc_22172_new_n8227_; 
wire core__abc_22172_new_n8228_; 
wire core__abc_22172_new_n8229_; 
wire core__abc_22172_new_n8230_; 
wire core__abc_22172_new_n8231_; 
wire core__abc_22172_new_n8233_; 
wire core__abc_22172_new_n8234_; 
wire core__abc_22172_new_n8235_; 
wire core__abc_22172_new_n8236_; 
wire core__abc_22172_new_n8237_; 
wire core__abc_22172_new_n8238_; 
wire core__abc_22172_new_n8239_; 
wire core__abc_22172_new_n8240_; 
wire core__abc_22172_new_n8241_; 
wire core__abc_22172_new_n8242_; 
wire core__abc_22172_new_n8243_; 
wire core__abc_22172_new_n8244_; 
wire core__abc_22172_new_n8245_; 
wire core__abc_22172_new_n8246_; 
wire core__abc_22172_new_n8247_; 
wire core__abc_22172_new_n8248_; 
wire core__abc_22172_new_n8250_; 
wire core__abc_22172_new_n8251_; 
wire core__abc_22172_new_n8252_; 
wire core__abc_22172_new_n8253_; 
wire core__abc_22172_new_n8254_; 
wire core__abc_22172_new_n8255_; 
wire core__abc_22172_new_n8256_; 
wire core__abc_22172_new_n8257_; 
wire core__abc_22172_new_n8258_; 
wire core__abc_22172_new_n8259_; 
wire core__abc_22172_new_n8260_; 
wire core__abc_22172_new_n8261_; 
wire core__abc_22172_new_n8262_; 
wire core__abc_22172_new_n8263_; 
wire core__abc_22172_new_n8264_; 
wire core__abc_22172_new_n8266_; 
wire core__abc_22172_new_n8267_; 
wire core__abc_22172_new_n8268_; 
wire core__abc_22172_new_n8269_; 
wire core__abc_22172_new_n8270_; 
wire core__abc_22172_new_n8271_; 
wire core__abc_22172_new_n8272_; 
wire core__abc_22172_new_n8273_; 
wire core__abc_22172_new_n8274_; 
wire core__abc_22172_new_n8275_; 
wire core__abc_22172_new_n8276_; 
wire core__abc_22172_new_n8277_; 
wire core__abc_22172_new_n8278_; 
wire core__abc_22172_new_n8279_; 
wire core__abc_22172_new_n8280_; 
wire core__abc_22172_new_n8282_; 
wire core__abc_22172_new_n8283_; 
wire core__abc_22172_new_n8284_; 
wire core__abc_22172_new_n8285_; 
wire core__abc_22172_new_n8286_; 
wire core__abc_22172_new_n8287_; 
wire core__abc_22172_new_n8288_; 
wire core__abc_22172_new_n8289_; 
wire core__abc_22172_new_n8290_; 
wire core__abc_22172_new_n8291_; 
wire core__abc_22172_new_n8292_; 
wire core__abc_22172_new_n8293_; 
wire core__abc_22172_new_n8294_; 
wire core__abc_22172_new_n8295_; 
wire core__abc_22172_new_n8297_; 
wire core__abc_22172_new_n8298_; 
wire core__abc_22172_new_n8299_; 
wire core__abc_22172_new_n8300_; 
wire core__abc_22172_new_n8301_; 
wire core__abc_22172_new_n8302_; 
wire core__abc_22172_new_n8303_; 
wire core__abc_22172_new_n8304_; 
wire core__abc_22172_new_n8305_; 
wire core__abc_22172_new_n8306_; 
wire core__abc_22172_new_n8307_; 
wire core__abc_22172_new_n8308_; 
wire core__abc_22172_new_n8309_; 
wire core__abc_22172_new_n8310_; 
wire core__abc_22172_new_n8311_; 
wire core__abc_22172_new_n8312_; 
wire core__abc_22172_new_n8314_; 
wire core__abc_22172_new_n8315_; 
wire core__abc_22172_new_n8316_; 
wire core__abc_22172_new_n8317_; 
wire core__abc_22172_new_n8318_; 
wire core__abc_22172_new_n8319_; 
wire core__abc_22172_new_n8320_; 
wire core__abc_22172_new_n8321_; 
wire core__abc_22172_new_n8322_; 
wire core__abc_22172_new_n8323_; 
wire core__abc_22172_new_n8324_; 
wire core__abc_22172_new_n8325_; 
wire core__abc_22172_new_n8326_; 
wire core__abc_22172_new_n8327_; 
wire core__abc_22172_new_n8328_; 
wire core__abc_22172_new_n8329_; 
wire core__abc_22172_new_n8331_; 
wire core__abc_22172_new_n8332_; 
wire core__abc_22172_new_n8333_; 
wire core__abc_22172_new_n8334_; 
wire core__abc_22172_new_n8335_; 
wire core__abc_22172_new_n8336_; 
wire core__abc_22172_new_n8337_; 
wire core__abc_22172_new_n8338_; 
wire core__abc_22172_new_n8339_; 
wire core__abc_22172_new_n8340_; 
wire core__abc_22172_new_n8341_; 
wire core__abc_22172_new_n8342_; 
wire core__abc_22172_new_n8343_; 
wire core__abc_22172_new_n8344_; 
wire core__abc_22172_new_n8345_; 
wire core__abc_22172_new_n8347_; 
wire core__abc_22172_new_n8348_; 
wire core__abc_22172_new_n8349_; 
wire core__abc_22172_new_n8350_; 
wire core__abc_22172_new_n8351_; 
wire core__abc_22172_new_n8352_; 
wire core__abc_22172_new_n8353_; 
wire core__abc_22172_new_n8354_; 
wire core__abc_22172_new_n8355_; 
wire core__abc_22172_new_n8356_; 
wire core__abc_22172_new_n8357_; 
wire core__abc_22172_new_n8358_; 
wire core__abc_22172_new_n8360_; 
wire core__abc_22172_new_n8361_; 
wire core__abc_22172_new_n8362_; 
wire core__abc_22172_new_n8363_; 
wire core__abc_22172_new_n8364_; 
wire core__abc_22172_new_n8365_; 
wire core__abc_22172_new_n8366_; 
wire core__abc_22172_new_n8367_; 
wire core__abc_22172_new_n8368_; 
wire core__abc_22172_new_n8369_; 
wire core__abc_22172_new_n8370_; 
wire core__abc_22172_new_n8371_; 
wire core__abc_22172_new_n8372_; 
wire core__abc_22172_new_n8373_; 
wire core__abc_22172_new_n8375_; 
wire core__abc_22172_new_n8376_; 
wire core__abc_22172_new_n8377_; 
wire core__abc_22172_new_n8378_; 
wire core__abc_22172_new_n8379_; 
wire core__abc_22172_new_n8380_; 
wire core__abc_22172_new_n8381_; 
wire core__abc_22172_new_n8382_; 
wire core__abc_22172_new_n8383_; 
wire core__abc_22172_new_n8384_; 
wire core__abc_22172_new_n8385_; 
wire core__abc_22172_new_n8386_; 
wire core__abc_22172_new_n8387_; 
wire core__abc_22172_new_n8388_; 
wire core__abc_22172_new_n8389_; 
wire core__abc_22172_new_n8391_; 
wire core__abc_22172_new_n8392_; 
wire core__abc_22172_new_n8393_; 
wire core__abc_22172_new_n8394_; 
wire core__abc_22172_new_n8395_; 
wire core__abc_22172_new_n8396_; 
wire core__abc_22172_new_n8397_; 
wire core__abc_22172_new_n8398_; 
wire core__abc_22172_new_n8399_; 
wire core__abc_22172_new_n8400_; 
wire core__abc_22172_new_n8401_; 
wire core__abc_22172_new_n8402_; 
wire core__abc_22172_new_n8403_; 
wire core__abc_22172_new_n8404_; 
wire core__abc_22172_new_n8405_; 
wire core__abc_22172_new_n8406_; 
wire core__abc_22172_new_n8408_; 
wire core__abc_22172_new_n8409_; 
wire core__abc_22172_new_n8410_; 
wire core__abc_22172_new_n8411_; 
wire core__abc_22172_new_n8412_; 
wire core__abc_22172_new_n8413_; 
wire core__abc_22172_new_n8414_; 
wire core__abc_22172_new_n8415_; 
wire core__abc_22172_new_n8416_; 
wire core__abc_22172_new_n8417_; 
wire core__abc_22172_new_n8418_; 
wire core__abc_22172_new_n8420_; 
wire core__abc_22172_new_n8421_; 
wire core__abc_22172_new_n8422_; 
wire core__abc_22172_new_n8423_; 
wire core__abc_22172_new_n8424_; 
wire core__abc_22172_new_n8425_; 
wire core__abc_22172_new_n8426_; 
wire core__abc_22172_new_n8427_; 
wire core__abc_22172_new_n8428_; 
wire core__abc_22172_new_n8429_; 
wire core__abc_22172_new_n8430_; 
wire core__abc_22172_new_n8431_; 
wire core__abc_22172_new_n8433_; 
wire core__abc_22172_new_n8434_; 
wire core__abc_22172_new_n8435_; 
wire core__abc_22172_new_n8436_; 
wire core__abc_22172_new_n8437_; 
wire core__abc_22172_new_n8438_; 
wire core__abc_22172_new_n8439_; 
wire core__abc_22172_new_n8440_; 
wire core__abc_22172_new_n8441_; 
wire core__abc_22172_new_n8442_; 
wire core__abc_22172_new_n8443_; 
wire core__abc_22172_new_n8445_; 
wire core__abc_22172_new_n8446_; 
wire core__abc_22172_new_n8447_; 
wire core__abc_22172_new_n8448_; 
wire core__abc_22172_new_n8449_; 
wire core__abc_22172_new_n8450_; 
wire core__abc_22172_new_n8451_; 
wire core__abc_22172_new_n8452_; 
wire core__abc_22172_new_n8453_; 
wire core__abc_22172_new_n8454_; 
wire core__abc_22172_new_n8455_; 
wire core__abc_22172_new_n8456_; 
wire core__abc_22172_new_n8458_; 
wire core__abc_22172_new_n8459_; 
wire core__abc_22172_new_n8460_; 
wire core__abc_22172_new_n8461_; 
wire core__abc_22172_new_n8462_; 
wire core__abc_22172_new_n8463_; 
wire core__abc_22172_new_n8464_; 
wire core__abc_22172_new_n8465_; 
wire core__abc_22172_new_n8466_; 
wire core__abc_22172_new_n8467_; 
wire core__abc_22172_new_n8468_; 
wire core__abc_22172_new_n8470_; 
wire core__abc_22172_new_n8471_; 
wire core__abc_22172_new_n8472_; 
wire core__abc_22172_new_n8473_; 
wire core__abc_22172_new_n8474_; 
wire core__abc_22172_new_n8475_; 
wire core__abc_22172_new_n8476_; 
wire core__abc_22172_new_n8477_; 
wire core__abc_22172_new_n8478_; 
wire core__abc_22172_new_n8479_; 
wire core__abc_22172_new_n8480_; 
wire core__abc_22172_new_n8482_; 
wire core__abc_22172_new_n8483_; 
wire core__abc_22172_new_n8484_; 
wire core__abc_22172_new_n8485_; 
wire core__abc_22172_new_n8486_; 
wire core__abc_22172_new_n8487_; 
wire core__abc_22172_new_n8488_; 
wire core__abc_22172_new_n8489_; 
wire core__abc_22172_new_n8490_; 
wire core__abc_22172_new_n8491_; 
wire core__abc_22172_new_n8493_; 
wire core__abc_22172_new_n8494_; 
wire core__abc_22172_new_n8495_; 
wire core__abc_22172_new_n8496_; 
wire core__abc_22172_new_n8497_; 
wire core__abc_22172_new_n8498_; 
wire core__abc_22172_new_n8499_; 
wire core__abc_22172_new_n8500_; 
wire core__abc_22172_new_n8501_; 
wire core__abc_22172_new_n8502_; 
wire core__abc_22172_new_n8504_; 
wire core__abc_22172_new_n8505_; 
wire core__abc_22172_new_n8506_; 
wire core__abc_22172_new_n8507_; 
wire core__abc_22172_new_n8508_; 
wire core__abc_22172_new_n8509_; 
wire core__abc_22172_new_n8510_; 
wire core__abc_22172_new_n8511_; 
wire core__abc_22172_new_n8512_; 
wire core__abc_22172_new_n8513_; 
wire core__abc_22172_new_n8515_; 
wire core__abc_22172_new_n8516_; 
wire core__abc_22172_new_n8517_; 
wire core__abc_22172_new_n8518_; 
wire core__abc_22172_new_n8519_; 
wire core__abc_22172_new_n8520_; 
wire core__abc_22172_new_n8521_; 
wire core__abc_22172_new_n8522_; 
wire core__abc_22172_new_n8523_; 
wire core__abc_22172_new_n8524_; 
wire core__abc_22172_new_n8525_; 
wire core__abc_22172_new_n8527_; 
wire core__abc_22172_new_n8528_; 
wire core__abc_22172_new_n8529_; 
wire core__abc_22172_new_n8530_; 
wire core__abc_22172_new_n8531_; 
wire core__abc_22172_new_n8532_; 
wire core__abc_22172_new_n8533_; 
wire core__abc_22172_new_n8534_; 
wire core__abc_22172_new_n8535_; 
wire core__abc_22172_new_n8536_; 
wire core__abc_22172_new_n8537_; 
wire core__abc_22172_new_n8539_; 
wire core__abc_22172_new_n8540_; 
wire core__abc_22172_new_n8541_; 
wire core__abc_22172_new_n8542_; 
wire core__abc_22172_new_n8543_; 
wire core__abc_22172_new_n8544_; 
wire core__abc_22172_new_n8545_; 
wire core__abc_22172_new_n8546_; 
wire core__abc_22172_new_n8547_; 
wire core__abc_22172_new_n8548_; 
wire core__abc_22172_new_n8549_; 
wire core__abc_22172_new_n8551_; 
wire core__abc_22172_new_n8552_; 
wire core__abc_22172_new_n8553_; 
wire core__abc_22172_new_n8554_; 
wire core__abc_22172_new_n8555_; 
wire core__abc_22172_new_n8556_; 
wire core__abc_22172_new_n8557_; 
wire core__abc_22172_new_n8558_; 
wire core__abc_22172_new_n8559_; 
wire core__abc_22172_new_n8560_; 
wire core__abc_22172_new_n8561_; 
wire core__abc_22172_new_n8563_; 
wire core__abc_22172_new_n8564_; 
wire core__abc_22172_new_n8565_; 
wire core__abc_22172_new_n8566_; 
wire core__abc_22172_new_n8567_; 
wire core__abc_22172_new_n8568_; 
wire core__abc_22172_new_n8569_; 
wire core__abc_22172_new_n8570_; 
wire core__abc_22172_new_n8571_; 
wire core__abc_22172_new_n8572_; 
wire core__abc_22172_new_n8574_; 
wire core__abc_22172_new_n8575_; 
wire core__abc_22172_new_n8576_; 
wire core__abc_22172_new_n8577_; 
wire core__abc_22172_new_n8578_; 
wire core__abc_22172_new_n8579_; 
wire core__abc_22172_new_n8580_; 
wire core__abc_22172_new_n8581_; 
wire core__abc_22172_new_n8582_; 
wire core__abc_22172_new_n8583_; 
wire core__abc_22172_new_n8584_; 
wire core__abc_22172_new_n8586_; 
wire core__abc_22172_new_n8587_; 
wire core__abc_22172_new_n8588_; 
wire core__abc_22172_new_n8589_; 
wire core__abc_22172_new_n8590_; 
wire core__abc_22172_new_n8591_; 
wire core__abc_22172_new_n8592_; 
wire core__abc_22172_new_n8593_; 
wire core__abc_22172_new_n8594_; 
wire core__abc_22172_new_n8595_; 
wire core__abc_22172_new_n8597_; 
wire core__abc_22172_new_n8598_; 
wire core__abc_22172_new_n8599_; 
wire core__abc_22172_new_n8600_; 
wire core__abc_22172_new_n8601_; 
wire core__abc_22172_new_n8602_; 
wire core__abc_22172_new_n8603_; 
wire core__abc_22172_new_n8604_; 
wire core__abc_22172_new_n8605_; 
wire core__abc_22172_new_n8606_; 
wire core__abc_22172_new_n8607_; 
wire core__abc_22172_new_n8608_; 
wire core__abc_22172_new_n8610_; 
wire core__abc_22172_new_n8611_; 
wire core__abc_22172_new_n8612_; 
wire core__abc_22172_new_n8613_; 
wire core__abc_22172_new_n8614_; 
wire core__abc_22172_new_n8615_; 
wire core__abc_22172_new_n8616_; 
wire core__abc_22172_new_n8617_; 
wire core__abc_22172_new_n8618_; 
wire core__abc_22172_new_n8619_; 
wire core__abc_22172_new_n8620_; 
wire core__abc_22172_new_n8621_; 
wire core__abc_22172_new_n8622_; 
wire core__abc_22172_new_n8624_; 
wire core__abc_22172_new_n8625_; 
wire core__abc_22172_new_n8626_; 
wire core__abc_22172_new_n8627_; 
wire core__abc_22172_new_n8628_; 
wire core__abc_22172_new_n8629_; 
wire core__abc_22172_new_n8630_; 
wire core__abc_22172_new_n8631_; 
wire core__abc_22172_new_n8632_; 
wire core__abc_22172_new_n8633_; 
wire core__abc_22172_new_n8634_; 
wire core__abc_22172_new_n8635_; 
wire core__abc_22172_new_n8636_; 
wire core__abc_22172_new_n8637_; 
wire core__abc_22172_new_n8639_; 
wire core__abc_22172_new_n8640_; 
wire core__abc_22172_new_n8641_; 
wire core__abc_22172_new_n8642_; 
wire core__abc_22172_new_n8643_; 
wire core__abc_22172_new_n8644_; 
wire core__abc_22172_new_n8645_; 
wire core__abc_22172_new_n8646_; 
wire core__abc_22172_new_n8647_; 
wire core__abc_22172_new_n8648_; 
wire core__abc_22172_new_n8649_; 
wire core__abc_22172_new_n8651_; 
wire core__abc_22172_new_n8652_; 
wire core__abc_22172_new_n8653_; 
wire core__abc_22172_new_n8654_; 
wire core__abc_22172_new_n8655_; 
wire core__abc_22172_new_n8656_; 
wire core__abc_22172_new_n8657_; 
wire core__abc_22172_new_n8658_; 
wire core__abc_22172_new_n8659_; 
wire core__abc_22172_new_n8660_; 
wire core__abc_22172_new_n8661_; 
wire core__abc_22172_new_n8663_; 
wire core__abc_22172_new_n8664_; 
wire core__abc_22172_new_n8665_; 
wire core__abc_22172_new_n8666_; 
wire core__abc_22172_new_n8667_; 
wire core__abc_22172_new_n8668_; 
wire core__abc_22172_new_n8669_; 
wire core__abc_22172_new_n8670_; 
wire core__abc_22172_new_n8671_; 
wire core__abc_22172_new_n8672_; 
wire core__abc_22172_new_n8674_; 
wire core__abc_22172_new_n8675_; 
wire core__abc_22172_new_n8676_; 
wire core__abc_22172_new_n8677_; 
wire core__abc_22172_new_n8678_; 
wire core__abc_22172_new_n8679_; 
wire core__abc_22172_new_n8680_; 
wire core__abc_22172_new_n8681_; 
wire core__abc_22172_new_n8682_; 
wire core__abc_22172_new_n8683_; 
wire core__abc_22172_new_n8684_; 
wire core__abc_22172_new_n8686_; 
wire core__abc_22172_new_n8687_; 
wire core__abc_22172_new_n8688_; 
wire core__abc_22172_new_n8689_; 
wire core__abc_22172_new_n8690_; 
wire core__abc_22172_new_n8691_; 
wire core__abc_22172_new_n8692_; 
wire core__abc_22172_new_n8693_; 
wire core__abc_22172_new_n8694_; 
wire core__abc_22172_new_n8695_; 
wire core__abc_22172_new_n8697_; 
wire core__abc_22172_new_n8698_; 
wire core__abc_22172_new_n8699_; 
wire core__abc_22172_new_n8700_; 
wire core__abc_22172_new_n8701_; 
wire core__abc_22172_new_n8702_; 
wire core__abc_22172_new_n8703_; 
wire core__abc_22172_new_n8704_; 
wire core__abc_22172_new_n8705_; 
wire core__abc_22172_new_n8706_; 
wire core__abc_22172_new_n8707_; 
wire core__abc_22172_new_n8708_; 
wire core__abc_22172_new_n8710_; 
wire core__abc_22172_new_n8711_; 
wire core__abc_22172_new_n8712_; 
wire core__abc_22172_new_n8713_; 
wire core__abc_22172_new_n8714_; 
wire core__abc_22172_new_n8715_; 
wire core__abc_22172_new_n8716_; 
wire core__abc_22172_new_n8717_; 
wire core__abc_22172_new_n8718_; 
wire core__abc_22172_new_n8719_; 
wire core__abc_22172_new_n8720_; 
wire core__abc_22172_new_n8722_; 
wire core__abc_22172_new_n8723_; 
wire core__abc_22172_new_n8724_; 
wire core__abc_22172_new_n8725_; 
wire core__abc_22172_new_n8726_; 
wire core__abc_22172_new_n8727_; 
wire core__abc_22172_new_n8728_; 
wire core__abc_22172_new_n8729_; 
wire core__abc_22172_new_n8730_; 
wire core__abc_22172_new_n8731_; 
wire core__abc_22172_new_n8732_; 
wire core__abc_22172_new_n8734_; 
wire core__abc_22172_new_n8735_; 
wire core__abc_22172_new_n8736_; 
wire core__abc_22172_new_n8737_; 
wire core__abc_22172_new_n8738_; 
wire core__abc_22172_new_n8739_; 
wire core__abc_22172_new_n8740_; 
wire core__abc_22172_new_n8741_; 
wire core__abc_22172_new_n8742_; 
wire core__abc_22172_new_n8743_; 
wire core__abc_22172_new_n8744_; 
wire core__abc_22172_new_n8746_; 
wire core__abc_22172_new_n8747_; 
wire core__abc_22172_new_n8748_; 
wire core__abc_22172_new_n8749_; 
wire core__abc_22172_new_n8750_; 
wire core__abc_22172_new_n8751_; 
wire core__abc_22172_new_n8752_; 
wire core__abc_22172_new_n8753_; 
wire core__abc_22172_new_n8754_; 
wire core__abc_22172_new_n8755_; 
wire core__abc_22172_new_n8757_; 
wire core__abc_22172_new_n8758_; 
wire core__abc_22172_new_n8759_; 
wire core__abc_22172_new_n8760_; 
wire core__abc_22172_new_n8761_; 
wire core__abc_22172_new_n8762_; 
wire core__abc_22172_new_n8763_; 
wire core__abc_22172_new_n8764_; 
wire core__abc_22172_new_n8765_; 
wire core__abc_22172_new_n8766_; 
wire core__abc_22172_new_n8768_; 
wire core__abc_22172_new_n8769_; 
wire core__abc_22172_new_n8770_; 
wire core__abc_22172_new_n8771_; 
wire core__abc_22172_new_n8772_; 
wire core__abc_22172_new_n8773_; 
wire core__abc_22172_new_n8774_; 
wire core__abc_22172_new_n8775_; 
wire core__abc_22172_new_n8776_; 
wire core__abc_22172_new_n8777_; 
wire core__abc_22172_new_n8778_; 
wire core__abc_22172_new_n8780_; 
wire core__abc_22172_new_n8781_; 
wire core__abc_22172_new_n8782_; 
wire core__abc_22172_new_n8783_; 
wire core__abc_22172_new_n8784_; 
wire core__abc_22172_new_n8785_; 
wire core__abc_22172_new_n8786_; 
wire core__abc_22172_new_n8787_; 
wire core__abc_22172_new_n8788_; 
wire core__abc_22172_new_n8789_; 
wire core__abc_22172_new_n8790_; 
wire core__abc_22172_new_n8792_; 
wire core__abc_22172_new_n8793_; 
wire core__abc_22172_new_n8794_; 
wire core__abc_22172_new_n8795_; 
wire core__abc_22172_new_n8796_; 
wire core__abc_22172_new_n8797_; 
wire core__abc_22172_new_n8798_; 
wire core__abc_22172_new_n8799_; 
wire core__abc_22172_new_n8800_; 
wire core__abc_22172_new_n8801_; 
wire core__abc_22172_new_n8803_; 
wire core__abc_22172_new_n8804_; 
wire core__abc_22172_new_n8805_; 
wire core__abc_22172_new_n8806_; 
wire core__abc_22172_new_n8807_; 
wire core__abc_22172_new_n8808_; 
wire core__abc_22172_new_n8809_; 
wire core__abc_22172_new_n8810_; 
wire core__abc_22172_new_n8811_; 
wire core__abc_22172_new_n8812_; 
wire core__abc_22172_new_n8813_; 
wire core__abc_22172_new_n8814_; 
wire core__abc_22172_new_n8816_; 
wire core__abc_22172_new_n8817_; 
wire core__abc_22172_new_n8818_; 
wire core__abc_22172_new_n8819_; 
wire core__abc_22172_new_n8820_; 
wire core__abc_22172_new_n8821_; 
wire core__abc_22172_new_n8822_; 
wire core__abc_22172_new_n8823_; 
wire core__abc_22172_new_n8824_; 
wire core__abc_22172_new_n8825_; 
wire core__abc_22172_new_n8826_; 
wire core__abc_22172_new_n8827_; 
wire core__abc_22172_new_n8829_; 
wire core__abc_22172_new_n8830_; 
wire core__abc_22172_new_n8831_; 
wire core__abc_22172_new_n8832_; 
wire core__abc_22172_new_n8833_; 
wire core__abc_22172_new_n8834_; 
wire core__abc_22172_new_n8835_; 
wire core__abc_22172_new_n8836_; 
wire core__abc_22172_new_n8837_; 
wire core__abc_22172_new_n8838_; 
wire core__abc_22172_new_n8839_; 
wire core__abc_22172_new_n8841_; 
wire core__abc_22172_new_n8842_; 
wire core__abc_22172_new_n8843_; 
wire core__abc_22172_new_n8844_; 
wire core__abc_22172_new_n8845_; 
wire core__abc_22172_new_n8846_; 
wire core__abc_22172_new_n8847_; 
wire core__abc_22172_new_n8848_; 
wire core__abc_22172_new_n8849_; 
wire core__abc_22172_new_n8850_; 
wire core__abc_22172_new_n8851_; 
wire core__abc_22172_new_n8852_; 
wire core__abc_22172_new_n8854_; 
wire core__abc_22172_new_n8855_; 
wire core__abc_22172_new_n8856_; 
wire core__abc_22172_new_n8857_; 
wire core__abc_22172_new_n8858_; 
wire core__abc_22172_new_n8859_; 
wire core__abc_22172_new_n8860_; 
wire core__abc_22172_new_n8861_; 
wire core__abc_22172_new_n8862_; 
wire core__abc_22172_new_n8863_; 
wire core__abc_22172_new_n8864_; 
wire core__abc_22172_new_n8866_; 
wire core__abc_22172_new_n8867_; 
wire core__abc_22172_new_n8868_; 
wire core__abc_22172_new_n8869_; 
wire core__abc_22172_new_n8870_; 
wire core__abc_22172_new_n8871_; 
wire core__abc_22172_new_n8872_; 
wire core__abc_22172_new_n8873_; 
wire core__abc_22172_new_n8874_; 
wire core__abc_22172_new_n8875_; 
wire core__abc_22172_new_n8877_; 
wire core__abc_22172_new_n8878_; 
wire core__abc_22172_new_n8879_; 
wire core__abc_22172_new_n8880_; 
wire core__abc_22172_new_n8881_; 
wire core__abc_22172_new_n8882_; 
wire core__abc_22172_new_n8883_; 
wire core__abc_22172_new_n8884_; 
wire core__abc_22172_new_n8885_; 
wire core__abc_22172_new_n8886_; 
wire core__abc_22172_new_n8888_; 
wire core__abc_22172_new_n8889_; 
wire core__abc_22172_new_n8890_; 
wire core__abc_22172_new_n8891_; 
wire core__abc_22172_new_n8892_; 
wire core__abc_22172_new_n8893_; 
wire core__abc_22172_new_n8894_; 
wire core__abc_22172_new_n8895_; 
wire core__abc_22172_new_n8896_; 
wire core__abc_22172_new_n8897_; 
wire core__abc_22172_new_n8898_; 
wire core__abc_22172_new_n8900_; 
wire core__abc_22172_new_n8901_; 
wire core__abc_22172_new_n8902_; 
wire core__abc_22172_new_n8903_; 
wire core__abc_22172_new_n8904_; 
wire core__abc_22172_new_n8905_; 
wire core__abc_22172_new_n8906_; 
wire core__abc_22172_new_n8907_; 
wire core__abc_22172_new_n8908_; 
wire core__abc_22172_new_n8909_; 
wire core__abc_22172_new_n8910_; 
wire core__abc_22172_new_n8911_; 
wire core__abc_22172_new_n8913_; 
wire core__abc_22172_new_n8914_; 
wire core__abc_22172_new_n8915_; 
wire core__abc_22172_new_n8916_; 
wire core__abc_22172_new_n8917_; 
wire core__abc_22172_new_n8918_; 
wire core__abc_22172_new_n8919_; 
wire core__abc_22172_new_n8920_; 
wire core__abc_22172_new_n8921_; 
wire core__abc_22172_new_n8922_; 
wire core__abc_22172_new_n8924_; 
wire core__abc_22172_new_n8925_; 
wire core__abc_22172_new_n8926_; 
wire core__abc_22172_new_n8927_; 
wire core__abc_22172_new_n8928_; 
wire core__abc_22172_new_n8929_; 
wire core__abc_22172_new_n8930_; 
wire core__abc_22172_new_n8931_; 
wire core__abc_22172_new_n8932_; 
wire core__abc_22172_new_n8933_; 
wire core__abc_22172_new_n8934_; 
wire core__abc_22172_new_n8935_; 
wire core__abc_22172_new_n8936_; 
wire core__abc_22172_new_n8938_; 
wire core__abc_22172_new_n8939_; 
wire core__abc_22172_new_n8940_; 
wire core__abc_22172_new_n8941_; 
wire core__abc_22172_new_n8942_; 
wire core__abc_22172_new_n8943_; 
wire core__abc_22172_new_n8944_; 
wire core__abc_22172_new_n8945_; 
wire core__abc_22172_new_n8946_; 
wire core__abc_22172_new_n8947_; 
wire core__abc_22172_new_n8949_; 
wire core__abc_22172_new_n8950_; 
wire core__abc_22172_new_n8951_; 
wire core__abc_22172_new_n8952_; 
wire core__abc_22172_new_n8953_; 
wire core__abc_22172_new_n8954_; 
wire core__abc_22172_new_n8955_; 
wire core__abc_22172_new_n8956_; 
wire core__abc_22172_new_n8957_; 
wire core__abc_22172_new_n8958_; 
wire core__abc_22172_new_n8959_; 
wire core__abc_22172_new_n8961_; 
wire core__abc_22172_new_n8962_; 
wire core__abc_22172_new_n8963_; 
wire core__abc_22172_new_n8964_; 
wire core__abc_22172_new_n8965_; 
wire core__abc_22172_new_n8966_; 
wire core__abc_22172_new_n8967_; 
wire core__abc_22172_new_n8968_; 
wire core__abc_22172_new_n8969_; 
wire core__abc_22172_new_n8970_; 
wire core__abc_22172_new_n8971_; 
wire core__abc_22172_new_n8973_; 
wire core__abc_22172_new_n8974_; 
wire core__abc_22172_new_n8975_; 
wire core__abc_22172_new_n8976_; 
wire core__abc_22172_new_n8977_; 
wire core__abc_22172_new_n8978_; 
wire core__abc_22172_new_n8979_; 
wire core__abc_22172_new_n8980_; 
wire core__abc_22172_new_n8981_; 
wire core__abc_22172_new_n8982_; 
wire core__abc_22172_new_n8984_; 
wire core__abc_22172_new_n8985_; 
wire core__abc_22172_new_n8986_; 
wire core__abc_22172_new_n8987_; 
wire core__abc_22172_new_n8988_; 
wire core__abc_22172_new_n8989_; 
wire core__abc_22172_new_n8990_; 
wire core__abc_22172_new_n8991_; 
wire core__abc_22172_new_n8992_; 
wire core__abc_22172_new_n8993_; 
wire core__abc_22172_new_n8995_; 
wire core__abc_22172_new_n8996_; 
wire core__abc_22172_new_n8997_; 
wire core__abc_22172_new_n8998_; 
wire core__abc_22172_new_n8999_; 
wire core__abc_22172_new_n9000_; 
wire core__abc_22172_new_n9001_; 
wire core__abc_22172_new_n9002_; 
wire core__abc_22172_new_n9003_; 
wire core__abc_22172_new_n9004_; 
wire core__abc_22172_new_n9005_; 
wire core__abc_22172_new_n9007_; 
wire core__abc_22172_new_n9008_; 
wire core__abc_22172_new_n9009_; 
wire core__abc_22172_new_n9010_; 
wire core__abc_22172_new_n9011_; 
wire core__abc_22172_new_n9012_; 
wire core__abc_22172_new_n9013_; 
wire core__abc_22172_new_n9014_; 
wire core__abc_22172_new_n9015_; 
wire core__abc_22172_new_n9016_; 
wire core__abc_22172_new_n9017_; 
wire core__abc_22172_new_n9018_; 
wire core__abc_22172_new_n9020_; 
wire core__abc_22172_new_n9021_; 
wire core__abc_22172_new_n9022_; 
wire core__abc_22172_new_n9023_; 
wire core__abc_22172_new_n9024_; 
wire core__abc_22172_new_n9025_; 
wire core__abc_22172_new_n9026_; 
wire core__abc_22172_new_n9027_; 
wire core__abc_22172_new_n9028_; 
wire core__abc_22172_new_n9029_; 
wire core__abc_22172_new_n9030_; 
wire core__abc_22172_new_n9032_; 
wire core__abc_22172_new_n9033_; 
wire core__abc_22172_new_n9034_; 
wire core__abc_22172_new_n9035_; 
wire core__abc_22172_new_n9036_; 
wire core__abc_22172_new_n9037_; 
wire core__abc_22172_new_n9038_; 
wire core__abc_22172_new_n9039_; 
wire core__abc_22172_new_n9040_; 
wire core__abc_22172_new_n9041_; 
wire core__abc_22172_new_n9042_; 
wire core__abc_22172_new_n9043_; 
wire core__abc_22172_new_n9045_; 
wire core__abc_22172_new_n9046_; 
wire core__abc_22172_new_n9047_; 
wire core__abc_22172_new_n9048_; 
wire core__abc_22172_new_n9049_; 
wire core__abc_22172_new_n9050_; 
wire core__abc_22172_new_n9051_; 
wire core__abc_22172_new_n9052_; 
wire core__abc_22172_new_n9053_; 
wire core__abc_22172_new_n9054_; 
wire core__abc_22172_new_n9056_; 
wire core__abc_22172_new_n9057_; 
wire core__abc_22172_new_n9058_; 
wire core__abc_22172_new_n9059_; 
wire core__abc_22172_new_n9060_; 
wire core__abc_22172_new_n9061_; 
wire core__abc_22172_new_n9062_; 
wire core__abc_22172_new_n9063_; 
wire core__abc_22172_new_n9064_; 
wire core__abc_22172_new_n9065_; 
wire core__abc_22172_new_n9067_; 
wire core__abc_22172_new_n9068_; 
wire core__abc_22172_new_n9069_; 
wire core__abc_22172_new_n9070_; 
wire core__abc_22172_new_n9071_; 
wire core__abc_22172_new_n9072_; 
wire core__abc_22172_new_n9073_; 
wire core__abc_22172_new_n9074_; 
wire core__abc_22172_new_n9075_; 
wire core__abc_22172_new_n9076_; 
wire core__abc_22172_new_n9077_; 
wire core__abc_22172_new_n9079_; 
wire core__abc_22172_new_n9080_; 
wire core__abc_22172_new_n9081_; 
wire core__abc_22172_new_n9082_; 
wire core__abc_22172_new_n9083_; 
wire core__abc_22172_new_n9084_; 
wire core__abc_22172_new_n9085_; 
wire core__abc_22172_new_n9086_; 
wire core__abc_22172_new_n9087_; 
wire core__abc_22172_new_n9088_; 
wire core__abc_22172_new_n9089_; 
wire core__abc_22172_new_n9090_; 
wire core__abc_22172_new_n9091_; 
wire core__abc_22172_new_n9092_; 
wire core__abc_22172_new_n9093_; 
wire core__abc_22172_new_n9094_; 
wire core__abc_22172_new_n9096_; 
wire core__abc_22172_new_n9097_; 
wire core__abc_22172_new_n9098_; 
wire core__abc_22172_new_n9099_; 
wire core__abc_22172_new_n9100_; 
wire core__abc_22172_new_n9101_; 
wire core__abc_22172_new_n9102_; 
wire core__abc_22172_new_n9103_; 
wire core__abc_22172_new_n9104_; 
wire core__abc_22172_new_n9105_; 
wire core__abc_22172_new_n9106_; 
wire core__abc_22172_new_n9108_; 
wire core__abc_22172_new_n9109_; 
wire core__abc_22172_new_n9110_; 
wire core__abc_22172_new_n9111_; 
wire core__abc_22172_new_n9112_; 
wire core__abc_22172_new_n9113_; 
wire core__abc_22172_new_n9114_; 
wire core__abc_22172_new_n9115_; 
wire core__abc_22172_new_n9116_; 
wire core__abc_22172_new_n9117_; 
wire core__abc_22172_new_n9118_; 
wire core__abc_22172_new_n9119_; 
wire core__abc_22172_new_n9120_; 
wire core__abc_22172_new_n9122_; 
wire core__abc_22172_new_n9123_; 
wire core__abc_22172_new_n9124_; 
wire core__abc_22172_new_n9125_; 
wire core__abc_22172_new_n9126_; 
wire core__abc_22172_new_n9127_; 
wire core__abc_22172_new_n9128_; 
wire core__abc_22172_new_n9129_; 
wire core__abc_22172_new_n9130_; 
wire core__abc_22172_new_n9131_; 
wire core__abc_22172_new_n9132_; 
wire core__abc_22172_new_n9134_; 
wire core__abc_22172_new_n9135_; 
wire core__abc_22172_new_n9136_; 
wire core__abc_22172_new_n9137_; 
wire core__abc_22172_new_n9138_; 
wire core__abc_22172_new_n9139_; 
wire core__abc_22172_new_n9140_; 
wire core__abc_22172_new_n9141_; 
wire core__abc_22172_new_n9142_; 
wire core__abc_22172_new_n9143_; 
wire core__abc_22172_new_n9144_; 
wire core__abc_22172_new_n9145_; 
wire core__abc_22172_new_n9146_; 
wire core__abc_22172_new_n9148_; 
wire core__abc_22172_new_n9149_; 
wire core__abc_22172_new_n9150_; 
wire core__abc_22172_new_n9151_; 
wire core__abc_22172_new_n9152_; 
wire core__abc_22172_new_n9153_; 
wire core__abc_22172_new_n9154_; 
wire core__abc_22172_new_n9155_; 
wire core__abc_22172_new_n9156_; 
wire core__abc_22172_new_n9157_; 
wire core__abc_22172_new_n9158_; 
wire core__abc_22172_new_n9160_; 
wire core__abc_22172_new_n9161_; 
wire core__abc_22172_new_n9162_; 
wire core__abc_22172_new_n9163_; 
wire core__abc_22172_new_n9164_; 
wire core__abc_22172_new_n9165_; 
wire core__abc_22172_new_n9166_; 
wire core__abc_22172_new_n9167_; 
wire core__abc_22172_new_n9168_; 
wire core__abc_22172_new_n9169_; 
wire core__abc_22172_new_n9170_; 
wire core__abc_22172_new_n9172_; 
wire core__abc_22172_new_n9173_; 
wire core__abc_22172_new_n9174_; 
wire core__abc_22172_new_n9175_; 
wire core__abc_22172_new_n9176_; 
wire core__abc_22172_new_n9177_; 
wire core__abc_22172_new_n9178_; 
wire core__abc_22172_new_n9179_; 
wire core__abc_22172_new_n9180_; 
wire core__abc_22172_new_n9181_; 
wire core__abc_22172_new_n9182_; 
wire core__abc_22172_new_n9184_; 
wire core__abc_22172_new_n9185_; 
wire core__abc_22172_new_n9186_; 
wire core__abc_22172_new_n9187_; 
wire core__abc_22172_new_n9188_; 
wire core__abc_22172_new_n9189_; 
wire core__abc_22172_new_n9190_; 
wire core__abc_22172_new_n9191_; 
wire core__abc_22172_new_n9192_; 
wire core__abc_22172_new_n9193_; 
wire core__abc_22172_new_n9194_; 
wire core__abc_22172_new_n9195_; 
wire core__abc_22172_new_n9196_; 
wire core__abc_22172_new_n9198_; 
wire core__abc_22172_new_n9199_; 
wire core__abc_22172_new_n9200_; 
wire core__abc_22172_new_n9201_; 
wire core__abc_22172_new_n9202_; 
wire core__abc_22172_new_n9203_; 
wire core__abc_22172_new_n9204_; 
wire core__abc_22172_new_n9205_; 
wire core__abc_22172_new_n9206_; 
wire core__abc_22172_new_n9207_; 
wire core__abc_22172_new_n9208_; 
wire core__abc_22172_new_n9209_; 
wire core__abc_22172_new_n9211_; 
wire core__abc_22172_new_n9212_; 
wire core__abc_22172_new_n9213_; 
wire core__abc_22172_new_n9214_; 
wire core__abc_22172_new_n9215_; 
wire core__abc_22172_new_n9216_; 
wire core__abc_22172_new_n9217_; 
wire core__abc_22172_new_n9218_; 
wire core__abc_22172_new_n9219_; 
wire core__abc_22172_new_n9220_; 
wire core__abc_22172_new_n9221_; 
wire core__abc_22172_new_n9222_; 
wire core__abc_22172_new_n9223_; 
wire core__abc_22172_new_n9225_; 
wire core__abc_22172_new_n9226_; 
wire core__abc_22172_new_n9227_; 
wire core__abc_22172_new_n9228_; 
wire core__abc_22172_new_n9229_; 
wire core__abc_22172_new_n9230_; 
wire core__abc_22172_new_n9231_; 
wire core__abc_22172_new_n9232_; 
wire core__abc_22172_new_n9233_; 
wire core__abc_22172_new_n9234_; 
wire core__abc_22172_new_n9235_; 
wire core__abc_22172_new_n9237_; 
wire core__abc_22172_new_n9238_; 
wire core__abc_22172_new_n9239_; 
wire core__abc_22172_new_n9240_; 
wire core__abc_22172_new_n9241_; 
wire core__abc_22172_new_n9242_; 
wire core__abc_22172_new_n9243_; 
wire core__abc_22172_new_n9244_; 
wire core__abc_22172_new_n9245_; 
wire core__abc_22172_new_n9246_; 
wire core__abc_22172_new_n9247_; 
wire core__abc_22172_new_n9248_; 
wire core__abc_22172_new_n9250_; 
wire core__abc_22172_new_n9251_; 
wire core__abc_22172_new_n9252_; 
wire core__abc_22172_new_n9253_; 
wire core__abc_22172_new_n9254_; 
wire core__abc_22172_new_n9255_; 
wire core__abc_22172_new_n9256_; 
wire core__abc_22172_new_n9257_; 
wire core__abc_22172_new_n9258_; 
wire core__abc_22172_new_n9259_; 
wire core__abc_22172_new_n9260_; 
wire core__abc_22172_new_n9262_; 
wire core__abc_22172_new_n9263_; 
wire core__abc_22172_new_n9264_; 
wire core__abc_22172_new_n9265_; 
wire core__abc_22172_new_n9266_; 
wire core__abc_22172_new_n9267_; 
wire core__abc_22172_new_n9268_; 
wire core__abc_22172_new_n9269_; 
wire core__abc_22172_new_n9270_; 
wire core__abc_22172_new_n9271_; 
wire core__abc_22172_new_n9272_; 
wire core__abc_22172_new_n9274_; 
wire core__abc_22172_new_n9275_; 
wire core__abc_22172_new_n9276_; 
wire core__abc_22172_new_n9277_; 
wire core__abc_22172_new_n9278_; 
wire core__abc_22172_new_n9279_; 
wire core__abc_22172_new_n9280_; 
wire core__abc_22172_new_n9281_; 
wire core__abc_22172_new_n9282_; 
wire core__abc_22172_new_n9283_; 
wire core__abc_22172_new_n9284_; 
wire core__abc_22172_new_n9286_; 
wire core__abc_22172_new_n9287_; 
wire core__abc_22172_new_n9288_; 
wire core__abc_22172_new_n9289_; 
wire core__abc_22172_new_n9290_; 
wire core__abc_22172_new_n9291_; 
wire core__abc_22172_new_n9292_; 
wire core__abc_22172_new_n9293_; 
wire core__abc_22172_new_n9294_; 
wire core__abc_22172_new_n9295_; 
wire core__abc_22172_new_n9296_; 
wire core__abc_22172_new_n9298_; 
wire core__abc_22172_new_n9299_; 
wire core__abc_22172_new_n9300_; 
wire core__abc_22172_new_n9301_; 
wire core__abc_22172_new_n9302_; 
wire core__abc_22172_new_n9303_; 
wire core__abc_22172_new_n9304_; 
wire core__abc_22172_new_n9305_; 
wire core__abc_22172_new_n9306_; 
wire core__abc_22172_new_n9307_; 
wire core__abc_22172_new_n9308_; 
wire core__abc_22172_new_n9309_; 
wire core__abc_22172_new_n9310_; 
wire core__abc_22172_new_n9312_; 
wire core__abc_22172_new_n9313_; 
wire core__abc_22172_new_n9314_; 
wire core__abc_22172_new_n9315_; 
wire core__abc_22172_new_n9316_; 
wire core__abc_22172_new_n9317_; 
wire core__abc_22172_new_n9318_; 
wire core__abc_22172_new_n9319_; 
wire core__abc_22172_new_n9320_; 
wire core__abc_22172_new_n9321_; 
wire core__abc_22172_new_n9322_; 
wire core__abc_22172_new_n9323_; 
wire core__abc_22172_new_n9325_; 
wire core__abc_22172_new_n9326_; 
wire core__abc_22172_new_n9327_; 
wire core__abc_22172_new_n9328_; 
wire core__abc_22172_new_n9329_; 
wire core__abc_22172_new_n9330_; 
wire core__abc_22172_new_n9331_; 
wire core__abc_22172_new_n9332_; 
wire core__abc_22172_new_n9333_; 
wire core__abc_22172_new_n9334_; 
wire core__abc_22172_new_n9335_; 
wire core__abc_22172_new_n9337_; 
wire core__abc_22172_new_n9338_; 
wire core__abc_22172_new_n9339_; 
wire core__abc_22172_new_n9340_; 
wire core__abc_22172_new_n9341_; 
wire core__abc_22172_new_n9342_; 
wire core__abc_22172_new_n9343_; 
wire core__abc_22172_new_n9344_; 
wire core__abc_22172_new_n9345_; 
wire core__abc_22172_new_n9346_; 
wire core__abc_22172_new_n9347_; 
wire core__abc_22172_new_n9348_; 
wire core__abc_22172_new_n9349_; 
wire core__abc_22172_new_n9351_; 
wire core__abc_22172_new_n9352_; 
wire core__abc_22172_new_n9353_; 
wire core__abc_22172_new_n9354_; 
wire core__abc_22172_new_n9355_; 
wire core__abc_22172_new_n9356_; 
wire core__abc_22172_new_n9357_; 
wire core__abc_22172_new_n9358_; 
wire core__abc_22172_new_n9359_; 
wire core__abc_22172_new_n9360_; 
wire core__abc_22172_new_n9361_; 
wire core__abc_22172_new_n9363_; 
wire core__abc_22172_new_n9364_; 
wire core__abc_22172_new_n9365_; 
wire core__abc_22172_new_n9366_; 
wire core__abc_22172_new_n9367_; 
wire core__abc_22172_new_n9368_; 
wire core__abc_22172_new_n9369_; 
wire core__abc_22172_new_n9370_; 
wire core__abc_22172_new_n9371_; 
wire core__abc_22172_new_n9372_; 
wire core__abc_22172_new_n9373_; 
wire core__abc_22172_new_n9375_; 
wire core__abc_22172_new_n9376_; 
wire core__abc_22172_new_n9377_; 
wire core__abc_22172_new_n9378_; 
wire core__abc_22172_new_n9379_; 
wire core__abc_22172_new_n9380_; 
wire core__abc_22172_new_n9381_; 
wire core__abc_22172_new_n9382_; 
wire core__abc_22172_new_n9383_; 
wire core__abc_22172_new_n9384_; 
wire core__abc_22172_new_n9385_; 
wire core__abc_22172_new_n9387_; 
wire core__abc_22172_new_n9388_; 
wire core__abc_22172_new_n9389_; 
wire core__abc_22172_new_n9390_; 
wire core__abc_22172_new_n9391_; 
wire core__abc_22172_new_n9392_; 
wire core__abc_22172_new_n9393_; 
wire core__abc_22172_new_n9394_; 
wire core__abc_22172_new_n9395_; 
wire core__abc_22172_new_n9396_; 
wire core__abc_22172_new_n9397_; 
wire core__abc_22172_new_n9399_; 
wire core__abc_22172_new_n9400_; 
wire core__abc_22172_new_n9401_; 
wire core__abc_22172_new_n9402_; 
wire core__abc_22172_new_n9403_; 
wire core__abc_22172_new_n9404_; 
wire core__abc_22172_new_n9405_; 
wire core__abc_22172_new_n9406_; 
wire core__abc_22172_new_n9407_; 
wire core__abc_22172_new_n9408_; 
wire core__abc_22172_new_n9409_; 
wire core__abc_22172_new_n9410_; 
wire core__abc_22172_new_n9412_; 
wire core__abc_22172_new_n9413_; 
wire core__abc_22172_new_n9414_; 
wire core__abc_22172_new_n9415_; 
wire core__abc_22172_new_n9416_; 
wire core__abc_22172_new_n9417_; 
wire core__abc_22172_new_n9418_; 
wire core__abc_22172_new_n9419_; 
wire core__abc_22172_new_n9420_; 
wire core__abc_22172_new_n9421_; 
wire core__abc_22172_new_n9422_; 
wire core__abc_22172_new_n9423_; 
wire core__abc_22172_new_n9425_; 
wire core__abc_22172_new_n9426_; 
wire core__abc_22172_new_n9427_; 
wire core__abc_22172_new_n9428_; 
wire core__abc_22172_new_n9429_; 
wire core__abc_22172_new_n9430_; 
wire core__abc_22172_new_n9431_; 
wire core__abc_22172_new_n9432_; 
wire core__abc_22172_new_n9433_; 
wire core__abc_22172_new_n9434_; 
wire core__abc_22172_new_n9435_; 
wire core__abc_22172_new_n9436_; 
wire core__abc_22172_new_n9438_; 
wire core__abc_22172_new_n9439_; 
wire core__abc_22172_new_n9440_; 
wire core__abc_22172_new_n9441_; 
wire core__abc_22172_new_n9442_; 
wire core__abc_22172_new_n9443_; 
wire core__abc_22172_new_n9444_; 
wire core__abc_22172_new_n9445_; 
wire core__abc_22172_new_n9446_; 
wire core__abc_22172_new_n9447_; 
wire core__abc_22172_new_n9448_; 
wire core__abc_22172_new_n9449_; 
wire core__abc_22172_new_n9450_; 
wire core__abc_22172_new_n9452_; 
wire core__abc_22172_new_n9453_; 
wire core__abc_22172_new_n9454_; 
wire core__abc_22172_new_n9455_; 
wire core__abc_22172_new_n9456_; 
wire core__abc_22172_new_n9457_; 
wire core__abc_22172_new_n9458_; 
wire core__abc_22172_new_n9459_; 
wire core__abc_22172_new_n9460_; 
wire core__abc_22172_new_n9461_; 
wire core__abc_22172_new_n9462_; 
wire core__abc_22172_new_n9464_; 
wire core__abc_22172_new_n9465_; 
wire core__abc_22172_new_n9466_; 
wire core__abc_22172_new_n9467_; 
wire core__abc_22172_new_n9468_; 
wire core__abc_22172_new_n9469_; 
wire core__abc_22172_new_n9470_; 
wire core__abc_22172_new_n9471_; 
wire core__abc_22172_new_n9472_; 
wire core__abc_22172_new_n9473_; 
wire core__abc_22172_new_n9474_; 
wire core__abc_22172_new_n9476_; 
wire core__abc_22172_new_n9477_; 
wire core__abc_22172_new_n9478_; 
wire core__abc_22172_new_n9479_; 
wire core__abc_22172_new_n9480_; 
wire core__abc_22172_new_n9481_; 
wire core__abc_22172_new_n9482_; 
wire core__abc_22172_new_n9483_; 
wire core__abc_22172_new_n9484_; 
wire core__abc_22172_new_n9485_; 
wire core__abc_22172_new_n9486_; 
wire core__abc_22172_new_n9488_; 
wire core__abc_22172_new_n9489_; 
wire core__abc_22172_new_n9490_; 
wire core__abc_22172_new_n9491_; 
wire core__abc_22172_new_n9492_; 
wire core__abc_22172_new_n9493_; 
wire core__abc_22172_new_n9494_; 
wire core__abc_22172_new_n9495_; 
wire core__abc_22172_new_n9496_; 
wire core__abc_22172_new_n9497_; 
wire core__abc_22172_new_n9498_; 
wire core__abc_22172_new_n9500_; 
wire core__abc_22172_new_n9501_; 
wire core__abc_22172_new_n9502_; 
wire core__abc_22172_new_n9503_; 
wire core__abc_22172_new_n9504_; 
wire core__abc_22172_new_n9505_; 
wire core__abc_22172_new_n9506_; 
wire core__abc_22172_new_n9507_; 
wire core__abc_22172_new_n9508_; 
wire core__abc_22172_new_n9509_; 
wire core__abc_22172_new_n9510_; 
wire core__abc_22172_new_n9512_; 
wire core__abc_22172_new_n9513_; 
wire core__abc_22172_new_n9514_; 
wire core__abc_22172_new_n9515_; 
wire core__abc_22172_new_n9516_; 
wire core__abc_22172_new_n9517_; 
wire core__abc_22172_new_n9518_; 
wire core__abc_22172_new_n9519_; 
wire core__abc_22172_new_n9520_; 
wire core__abc_22172_new_n9521_; 
wire core__abc_22172_new_n9522_; 
wire core__abc_22172_new_n9524_; 
wire core__abc_22172_new_n9525_; 
wire core__abc_22172_new_n9526_; 
wire core__abc_22172_new_n9527_; 
wire core__abc_22172_new_n9528_; 
wire core__abc_22172_new_n9529_; 
wire core__abc_22172_new_n9530_; 
wire core__abc_22172_new_n9531_; 
wire core__abc_22172_new_n9532_; 
wire core__abc_22172_new_n9533_; 
wire core__abc_22172_new_n9534_; 
wire core__abc_22172_new_n9536_; 
wire core__abc_22172_new_n9537_; 
wire core__abc_22172_new_n9538_; 
wire core__abc_22172_new_n9539_; 
wire core__abc_22172_new_n9540_; 
wire core__abc_22172_new_n9541_; 
wire core__abc_22172_new_n9542_; 
wire core__abc_22172_new_n9543_; 
wire core__abc_22172_new_n9544_; 
wire core__abc_22172_new_n9545_; 
wire core__abc_22172_new_n9546_; 
wire core__abc_22172_new_n9548_; 
wire core__abc_22172_new_n9549_; 
wire core__abc_22172_new_n9550_; 
wire core__abc_22172_new_n9551_; 
wire core__abc_22172_new_n9552_; 
wire core__abc_22172_new_n9553_; 
wire core__abc_22172_new_n9554_; 
wire core__abc_22172_new_n9555_; 
wire core__abc_22172_new_n9556_; 
wire core__abc_22172_new_n9557_; 
wire core__abc_22172_new_n9558_; 
wire core__abc_22172_new_n9560_; 
wire core__abc_22172_new_n9561_; 
wire core__abc_22172_new_n9562_; 
wire core__abc_22172_new_n9563_; 
wire core__abc_22172_new_n9564_; 
wire core__abc_22172_new_n9565_; 
wire core__abc_22172_new_n9566_; 
wire core__abc_22172_new_n9567_; 
wire core__abc_22172_new_n9568_; 
wire core__abc_22172_new_n9569_; 
wire core__abc_22172_new_n9570_; 
wire core__abc_22172_new_n9572_; 
wire core__abc_22172_new_n9573_; 
wire core__abc_22172_new_n9574_; 
wire core__abc_22172_new_n9575_; 
wire core__abc_22172_new_n9576_; 
wire core__abc_22172_new_n9577_; 
wire core__abc_22172_new_n9578_; 
wire core__abc_22172_new_n9579_; 
wire core__abc_22172_new_n9580_; 
wire core__abc_22172_new_n9581_; 
wire core__abc_22172_new_n9582_; 
wire core__abc_22172_new_n9584_; 
wire core__abc_22172_new_n9585_; 
wire core__abc_22172_new_n9586_; 
wire core__abc_22172_new_n9587_; 
wire core__abc_22172_new_n9588_; 
wire core__abc_22172_new_n9589_; 
wire core__abc_22172_new_n9590_; 
wire core__abc_22172_new_n9591_; 
wire core__abc_22172_new_n9592_; 
wire core__abc_22172_new_n9593_; 
wire core__abc_22172_new_n9594_; 
wire core__abc_22172_new_n9596_; 
wire core__abc_22172_new_n9597_; 
wire core__abc_22172_new_n9598_; 
wire core__abc_22172_new_n9599_; 
wire core__abc_22172_new_n9600_; 
wire core__abc_22172_new_n9601_; 
wire core__abc_22172_new_n9602_; 
wire core__abc_22172_new_n9603_; 
wire core__abc_22172_new_n9604_; 
wire core__abc_22172_new_n9605_; 
wire core__abc_22172_new_n9606_; 
wire core__abc_22172_new_n9607_; 
wire core__abc_22172_new_n9609_; 
wire core__abc_22172_new_n9610_; 
wire core__abc_22172_new_n9611_; 
wire core__abc_22172_new_n9612_; 
wire core__abc_22172_new_n9613_; 
wire core__abc_22172_new_n9614_; 
wire core__abc_22172_new_n9615_; 
wire core__abc_22172_new_n9616_; 
wire core__abc_22172_new_n9617_; 
wire core__abc_22172_new_n9618_; 
wire core__abc_22172_new_n9619_; 
wire core__abc_22172_new_n9621_; 
wire core__abc_22172_new_n9622_; 
wire core__abc_22172_new_n9623_; 
wire core__abc_22172_new_n9624_; 
wire core__abc_22172_new_n9625_; 
wire core__abc_22172_new_n9626_; 
wire core__abc_22172_new_n9627_; 
wire core__abc_22172_new_n9628_; 
wire core__abc_22172_new_n9629_; 
wire core__abc_22172_new_n9630_; 
wire core__abc_22172_new_n9631_; 
wire core__abc_22172_new_n9632_; 
wire core__abc_22172_new_n9633_; 
wire core__abc_22172_new_n9635_; 
wire core__abc_22172_new_n9636_; 
wire core__abc_22172_new_n9637_; 
wire core__abc_22172_new_n9638_; 
wire core__abc_22172_new_n9639_; 
wire core__abc_22172_new_n9640_; 
wire core__abc_22172_new_n9641_; 
wire core__abc_22172_new_n9642_; 
wire core__abc_22172_new_n9643_; 
wire core__abc_22172_new_n9644_; 
wire core__abc_22172_new_n9645_; 
wire core__abc_22172_new_n9647_; 
wire core__abc_22172_new_n9648_; 
wire core__abc_22172_new_n9649_; 
wire core__abc_22172_new_n9650_; 
wire core__abc_22172_new_n9651_; 
wire core__abc_22172_new_n9652_; 
wire core__abc_22172_new_n9653_; 
wire core__abc_22172_new_n9654_; 
wire core__abc_22172_new_n9655_; 
wire core__abc_22172_new_n9656_; 
wire core__abc_22172_new_n9657_; 
wire core__abc_22172_new_n9659_; 
wire core__abc_22172_new_n9660_; 
wire core__abc_22172_new_n9661_; 
wire core__abc_22172_new_n9662_; 
wire core__abc_22172_new_n9663_; 
wire core__abc_22172_new_n9664_; 
wire core__abc_22172_new_n9665_; 
wire core__abc_22172_new_n9666_; 
wire core__abc_22172_new_n9667_; 
wire core__abc_22172_new_n9668_; 
wire core__abc_22172_new_n9669_; 
wire core__abc_22172_new_n9671_; 
wire core__abc_22172_new_n9672_; 
wire core__abc_22172_new_n9673_; 
wire core__abc_22172_new_n9674_; 
wire core__abc_22172_new_n9675_; 
wire core__abc_22172_new_n9676_; 
wire core__abc_22172_new_n9677_; 
wire core__abc_22172_new_n9678_; 
wire core__abc_22172_new_n9679_; 
wire core__abc_22172_new_n9680_; 
wire core__abc_22172_new_n9681_; 
wire core__abc_22172_new_n9683_; 
wire core__abc_22172_new_n9684_; 
wire core__abc_22172_new_n9685_; 
wire core__abc_22172_new_n9686_; 
wire core__abc_22172_new_n9687_; 
wire core__abc_22172_new_n9688_; 
wire core__abc_22172_new_n9689_; 
wire core__abc_22172_new_n9690_; 
wire core__abc_22172_new_n9691_; 
wire core__abc_22172_new_n9692_; 
wire core__abc_22172_new_n9693_; 
wire core__abc_22172_new_n9695_; 
wire core__abc_22172_new_n9696_; 
wire core__abc_22172_new_n9697_; 
wire core__abc_22172_new_n9698_; 
wire core__abc_22172_new_n9699_; 
wire core__abc_22172_new_n9700_; 
wire core__abc_22172_new_n9701_; 
wire core__abc_22172_new_n9702_; 
wire core__abc_22172_new_n9703_; 
wire core__abc_22172_new_n9704_; 
wire core__abc_22172_new_n9705_; 
wire core__abc_22172_new_n9706_; 
wire core__abc_22172_new_n9707_; 
wire core__abc_22172_new_n9709_; 
wire core__abc_22172_new_n9710_; 
wire core__abc_22172_new_n9711_; 
wire core__abc_22172_new_n9712_; 
wire core__abc_22172_new_n9713_; 
wire core__abc_22172_new_n9714_; 
wire core__abc_22172_new_n9715_; 
wire core__abc_22172_new_n9716_; 
wire core__abc_22172_new_n9717_; 
wire core__abc_22172_new_n9718_; 
wire core__abc_22172_new_n9719_; 
wire core__abc_22172_new_n9720_; 
wire core__abc_22172_new_n9721_; 
wire core__abc_22172_new_n9723_; 
wire core__abc_22172_new_n9724_; 
wire core__abc_22172_new_n9725_; 
wire core__abc_22172_new_n9726_; 
wire core__abc_22172_new_n9727_; 
wire core__abc_22172_new_n9728_; 
wire core__abc_22172_new_n9729_; 
wire core__abc_22172_new_n9730_; 
wire core__abc_22172_new_n9731_; 
wire core__abc_22172_new_n9732_; 
wire core__abc_22172_new_n9733_; 
wire core__abc_22172_new_n9735_; 
wire core__abc_22172_new_n9736_; 
wire core__abc_22172_new_n9737_; 
wire core__abc_22172_new_n9738_; 
wire core__abc_22172_new_n9739_; 
wire core__abc_22172_new_n9740_; 
wire core__abc_22172_new_n9741_; 
wire core__abc_22172_new_n9742_; 
wire core__abc_22172_new_n9743_; 
wire core__abc_22172_new_n9744_; 
wire core__abc_22172_new_n9745_; 
wire core__abc_22172_new_n9746_; 
wire core__abc_22172_new_n9748_; 
wire core__abc_22172_new_n9749_; 
wire core__abc_22172_new_n9750_; 
wire core__abc_22172_new_n9751_; 
wire core__abc_22172_new_n9752_; 
wire core__abc_22172_new_n9753_; 
wire core__abc_22172_new_n9754_; 
wire core__abc_22172_new_n9755_; 
wire core__abc_22172_new_n9756_; 
wire core__abc_22172_new_n9757_; 
wire core__abc_22172_new_n9758_; 
wire core__abc_22172_new_n9760_; 
wire core__abc_22172_new_n9761_; 
wire core__abc_22172_new_n9762_; 
wire core__abc_22172_new_n9763_; 
wire core__abc_22172_new_n9764_; 
wire core__abc_22172_new_n9765_; 
wire core__abc_22172_new_n9766_; 
wire core__abc_22172_new_n9767_; 
wire core__abc_22172_new_n9768_; 
wire core__abc_22172_new_n9769_; 
wire core__abc_22172_new_n9770_; 
wire core__abc_22172_new_n9772_; 
wire core__abc_22172_new_n9773_; 
wire core__abc_22172_new_n9774_; 
wire core__abc_22172_new_n9775_; 
wire core__abc_22172_new_n9776_; 
wire core__abc_22172_new_n9777_; 
wire core__abc_22172_new_n9778_; 
wire core__abc_22172_new_n9779_; 
wire core__abc_22172_new_n9780_; 
wire core__abc_22172_new_n9781_; 
wire core__abc_22172_new_n9782_; 
wire core__abc_22172_new_n9784_; 
wire core__abc_22172_new_n9785_; 
wire core__abc_22172_new_n9786_; 
wire core__abc_22172_new_n9787_; 
wire core__abc_22172_new_n9788_; 
wire core__abc_22172_new_n9789_; 
wire core__abc_22172_new_n9790_; 
wire core__abc_22172_new_n9791_; 
wire core__abc_22172_new_n9792_; 
wire core__abc_22172_new_n9793_; 
wire core__abc_22172_new_n9794_; 
wire core__abc_22172_new_n9795_; 
wire core__abc_22172_new_n9796_; 
wire core__abc_22172_new_n9798_; 
wire core__abc_22172_new_n9799_; 
wire core__abc_22172_new_n9800_; 
wire core__abc_22172_new_n9801_; 
wire core__abc_22172_new_n9802_; 
wire core__abc_22172_new_n9803_; 
wire core__abc_22172_new_n9804_; 
wire core__abc_22172_new_n9805_; 
wire core__abc_22172_new_n9806_; 
wire core__abc_22172_new_n9807_; 
wire core__abc_22172_new_n9808_; 
wire core__abc_22172_new_n9809_; 
wire core__abc_22172_new_n9810_; 
wire core__abc_22172_new_n9812_; 
wire core__abc_22172_new_n9813_; 
wire core__abc_22172_new_n9814_; 
wire core__abc_22172_new_n9815_; 
wire core__abc_22172_new_n9816_; 
wire core__abc_22172_new_n9817_; 
wire core__abc_22172_new_n9818_; 
wire core__abc_22172_new_n9819_; 
wire core__abc_22172_new_n9820_; 
wire core__abc_22172_new_n9821_; 
wire core__abc_22172_new_n9822_; 
wire core__abc_22172_new_n9823_; 
wire core__abc_22172_new_n9825_; 
wire core__abc_22172_new_n9826_; 
wire core__abc_22172_new_n9827_; 
wire core__abc_22172_new_n9828_; 
wire core__abc_22172_new_n9829_; 
wire core__abc_22172_new_n9830_; 
wire core__abc_22172_new_n9831_; 
wire core__abc_22172_new_n9832_; 
wire core__abc_22172_new_n9833_; 
wire core__abc_22172_new_n9834_; 
wire core__abc_22172_new_n9835_; 
wire core__abc_22172_new_n9836_; 
wire core__abc_22172_new_n9838_; 
wire core__abc_22172_new_n9839_; 
wire core__abc_22172_new_n9840_; 
wire core__abc_22172_new_n9841_; 
wire core__abc_22172_new_n9842_; 
wire core__abc_22172_new_n9843_; 
wire core__abc_22172_new_n9844_; 
wire core__abc_22172_new_n9845_; 
wire core__abc_22172_new_n9846_; 
wire core__abc_22172_new_n9847_; 
wire core__abc_22172_new_n9848_; 
wire core__abc_22172_new_n9849_; 
wire core__abc_22172_new_n9850_; 
wire core__abc_22172_new_n9852_; 
wire core__abc_22172_new_n9853_; 
wire core__abc_22172_new_n9854_; 
wire core__abc_22172_new_n9855_; 
wire core__abc_22172_new_n9856_; 
wire core__abc_22172_new_n9857_; 
wire core__abc_22172_new_n9858_; 
wire core__abc_22172_new_n9859_; 
wire core__abc_22172_new_n9860_; 
wire core__abc_22172_new_n9861_; 
wire core__abc_22172_new_n9862_; 
wire core__abc_22172_new_n9864_; 
wire core__abc_22172_new_n9865_; 
wire core__abc_22172_new_n9866_; 
wire core__abc_22172_new_n9867_; 
wire core__abc_22172_new_n9868_; 
wire core__abc_22172_new_n9869_; 
wire core__abc_22172_new_n9870_; 
wire core__abc_22172_new_n9871_; 
wire core__abc_22172_new_n9872_; 
wire core__abc_22172_new_n9873_; 
wire core__abc_22172_new_n9874_; 
wire core__abc_22172_new_n9876_; 
wire core__abc_22172_new_n9877_; 
wire core__abc_22172_new_n9878_; 
wire core__abc_22172_new_n9879_; 
wire core__abc_22172_new_n9880_; 
wire core__abc_22172_new_n9881_; 
wire core__abc_22172_new_n9882_; 
wire core__abc_22172_new_n9883_; 
wire core__abc_22172_new_n9884_; 
wire core__abc_22172_new_n9885_; 
wire core__abc_22172_new_n9886_; 
wire core__abc_22172_new_n9888_; 
wire core__abc_22172_new_n9890_; 
wire core__abc_22172_new_n9891_; 
wire core__abc_22172_new_n9895_; 
wire core__abc_22172_new_n9896_; 
wire core__abc_22172_new_n9897_; 
wire core__abc_22172_new_n9898_; 
wire core_compress; 
wire core_compression_rounds_0_; 
wire core_compression_rounds_1_; 
wire core_compression_rounds_2_; 
wire core_compression_rounds_3_; 
wire core_final_rounds_0_; 
wire core_final_rounds_1_; 
wire core_final_rounds_2_; 
wire core_final_rounds_3_; 
wire core_finalize; 
wire core_initalize; 
wire core_key_0_; 
wire core_key_100_; 
wire core_key_101_; 
wire core_key_102_; 
wire core_key_103_; 
wire core_key_104_; 
wire core_key_105_; 
wire core_key_106_; 
wire core_key_107_; 
wire core_key_108_; 
wire core_key_109_; 
wire core_key_10_; 
wire core_key_110_; 
wire core_key_111_; 
wire core_key_112_; 
wire core_key_113_; 
wire core_key_114_; 
wire core_key_115_; 
wire core_key_116_; 
wire core_key_117_; 
wire core_key_118_; 
wire core_key_119_; 
wire core_key_11_; 
wire core_key_120_; 
wire core_key_121_; 
wire core_key_122_; 
wire core_key_123_; 
wire core_key_124_; 
wire core_key_125_; 
wire core_key_126_; 
wire core_key_127_; 
wire core_key_12_; 
wire core_key_13_; 
wire core_key_14_; 
wire core_key_15_; 
wire core_key_16_; 
wire core_key_17_; 
wire core_key_18_; 
wire core_key_19_; 
wire core_key_1_; 
wire core_key_20_; 
wire core_key_21_; 
wire core_key_22_; 
wire core_key_23_; 
wire core_key_24_; 
wire core_key_25_; 
wire core_key_26_; 
wire core_key_27_; 
wire core_key_28_; 
wire core_key_29_; 
wire core_key_2_; 
wire core_key_30_; 
wire core_key_31_; 
wire core_key_32_; 
wire core_key_33_; 
wire core_key_34_; 
wire core_key_35_; 
wire core_key_36_; 
wire core_key_37_; 
wire core_key_38_; 
wire core_key_39_; 
wire core_key_3_; 
wire core_key_40_; 
wire core_key_41_; 
wire core_key_42_; 
wire core_key_43_; 
wire core_key_44_; 
wire core_key_45_; 
wire core_key_46_; 
wire core_key_47_; 
wire core_key_48_; 
wire core_key_49_; 
wire core_key_4_; 
wire core_key_50_; 
wire core_key_51_; 
wire core_key_52_; 
wire core_key_53_; 
wire core_key_54_; 
wire core_key_55_; 
wire core_key_56_; 
wire core_key_57_; 
wire core_key_58_; 
wire core_key_59_; 
wire core_key_5_; 
wire core_key_60_; 
wire core_key_61_; 
wire core_key_62_; 
wire core_key_63_; 
wire core_key_64_; 
wire core_key_65_; 
wire core_key_66_; 
wire core_key_67_; 
wire core_key_68_; 
wire core_key_69_; 
wire core_key_6_; 
wire core_key_70_; 
wire core_key_71_; 
wire core_key_72_; 
wire core_key_73_; 
wire core_key_74_; 
wire core_key_75_; 
wire core_key_76_; 
wire core_key_77_; 
wire core_key_78_; 
wire core_key_79_; 
wire core_key_7_; 
wire core_key_80_; 
wire core_key_81_; 
wire core_key_82_; 
wire core_key_83_; 
wire core_key_84_; 
wire core_key_85_; 
wire core_key_86_; 
wire core_key_87_; 
wire core_key_88_; 
wire core_key_89_; 
wire core_key_8_; 
wire core_key_90_; 
wire core_key_91_; 
wire core_key_92_; 
wire core_key_93_; 
wire core_key_94_; 
wire core_key_95_; 
wire core_key_96_; 
wire core_key_97_; 
wire core_key_98_; 
wire core_key_99_; 
wire core_key_9_; 
wire core_long; 
wire core_loop_ctr_reg_0_; 
wire core_loop_ctr_reg_1_; 
wire core_loop_ctr_reg_2_; 
wire core_loop_ctr_reg_3_; 
wire core_mi_0_; 
wire core_mi_10_; 
wire core_mi_11_; 
wire core_mi_12_; 
wire core_mi_13_; 
wire core_mi_14_; 
wire core_mi_15_; 
wire core_mi_16_; 
wire core_mi_17_; 
wire core_mi_18_; 
wire core_mi_19_; 
wire core_mi_1_; 
wire core_mi_20_; 
wire core_mi_21_; 
wire core_mi_22_; 
wire core_mi_23_; 
wire core_mi_24_; 
wire core_mi_25_; 
wire core_mi_26_; 
wire core_mi_27_; 
wire core_mi_28_; 
wire core_mi_29_; 
wire core_mi_2_; 
wire core_mi_30_; 
wire core_mi_31_; 
wire core_mi_32_; 
wire core_mi_33_; 
wire core_mi_34_; 
wire core_mi_35_; 
wire core_mi_36_; 
wire core_mi_37_; 
wire core_mi_38_; 
wire core_mi_39_; 
wire core_mi_3_; 
wire core_mi_40_; 
wire core_mi_41_; 
wire core_mi_42_; 
wire core_mi_43_; 
wire core_mi_44_; 
wire core_mi_45_; 
wire core_mi_46_; 
wire core_mi_47_; 
wire core_mi_48_; 
wire core_mi_49_; 
wire core_mi_4_; 
wire core_mi_50_; 
wire core_mi_51_; 
wire core_mi_52_; 
wire core_mi_53_; 
wire core_mi_54_; 
wire core_mi_55_; 
wire core_mi_56_; 
wire core_mi_57_; 
wire core_mi_58_; 
wire core_mi_59_; 
wire core_mi_5_; 
wire core_mi_60_; 
wire core_mi_61_; 
wire core_mi_62_; 
wire core_mi_63_; 
wire core_mi_6_; 
wire core_mi_7_; 
wire core_mi_8_; 
wire core_mi_9_; 
wire core_mi_reg_0_; 
wire core_mi_reg_10_; 
wire core_mi_reg_11_; 
wire core_mi_reg_12_; 
wire core_mi_reg_13_; 
wire core_mi_reg_14_; 
wire core_mi_reg_15_; 
wire core_mi_reg_16_; 
wire core_mi_reg_17_; 
wire core_mi_reg_18_; 
wire core_mi_reg_19_; 
wire core_mi_reg_1_; 
wire core_mi_reg_20_; 
wire core_mi_reg_21_; 
wire core_mi_reg_22_; 
wire core_mi_reg_23_; 
wire core_mi_reg_24_; 
wire core_mi_reg_25_; 
wire core_mi_reg_26_; 
wire core_mi_reg_27_; 
wire core_mi_reg_28_; 
wire core_mi_reg_29_; 
wire core_mi_reg_2_; 
wire core_mi_reg_30_; 
wire core_mi_reg_31_; 
wire core_mi_reg_32_; 
wire core_mi_reg_33_; 
wire core_mi_reg_34_; 
wire core_mi_reg_35_; 
wire core_mi_reg_36_; 
wire core_mi_reg_37_; 
wire core_mi_reg_38_; 
wire core_mi_reg_39_; 
wire core_mi_reg_3_; 
wire core_mi_reg_40_; 
wire core_mi_reg_41_; 
wire core_mi_reg_42_; 
wire core_mi_reg_43_; 
wire core_mi_reg_44_; 
wire core_mi_reg_45_; 
wire core_mi_reg_46_; 
wire core_mi_reg_47_; 
wire core_mi_reg_48_; 
wire core_mi_reg_49_; 
wire core_mi_reg_4_; 
wire core_mi_reg_50_; 
wire core_mi_reg_51_; 
wire core_mi_reg_52_; 
wire core_mi_reg_53_; 
wire core_mi_reg_54_; 
wire core_mi_reg_55_; 
wire core_mi_reg_56_; 
wire core_mi_reg_57_; 
wire core_mi_reg_58_; 
wire core_mi_reg_59_; 
wire core_mi_reg_5_; 
wire core_mi_reg_60_; 
wire core_mi_reg_61_; 
wire core_mi_reg_62_; 
wire core_mi_reg_63_; 
wire core_mi_reg_6_; 
wire core_mi_reg_7_; 
wire core_mi_reg_8_; 
wire core_mi_reg_9_; 
wire core_ready; 
wire core_siphash_ctrl_reg_0_; 
wire core_siphash_ctrl_reg_1_; 
wire core_siphash_ctrl_reg_2_; 
wire core_siphash_ctrl_reg_3_; 
wire core_siphash_ctrl_reg_4_; 
wire core_siphash_ctrl_reg_5_; 
wire core_siphash_ctrl_reg_6_; 
wire core_siphash_valid_reg; 
wire core_siphash_word1_we; 
wire core_siphash_word_0_; 
wire core_siphash_word_100_; 
wire core_siphash_word_101_; 
wire core_siphash_word_102_; 
wire core_siphash_word_103_; 
wire core_siphash_word_104_; 
wire core_siphash_word_105_; 
wire core_siphash_word_106_; 
wire core_siphash_word_107_; 
wire core_siphash_word_108_; 
wire core_siphash_word_109_; 
wire core_siphash_word_10_; 
wire core_siphash_word_110_; 
wire core_siphash_word_111_; 
wire core_siphash_word_112_; 
wire core_siphash_word_113_; 
wire core_siphash_word_114_; 
wire core_siphash_word_115_; 
wire core_siphash_word_116_; 
wire core_siphash_word_117_; 
wire core_siphash_word_118_; 
wire core_siphash_word_119_; 
wire core_siphash_word_11_; 
wire core_siphash_word_120_; 
wire core_siphash_word_121_; 
wire core_siphash_word_122_; 
wire core_siphash_word_123_; 
wire core_siphash_word_124_; 
wire core_siphash_word_125_; 
wire core_siphash_word_126_; 
wire core_siphash_word_127_; 
wire core_siphash_word_12_; 
wire core_siphash_word_13_; 
wire core_siphash_word_14_; 
wire core_siphash_word_15_; 
wire core_siphash_word_16_; 
wire core_siphash_word_17_; 
wire core_siphash_word_18_; 
wire core_siphash_word_19_; 
wire core_siphash_word_1_; 
wire core_siphash_word_20_; 
wire core_siphash_word_21_; 
wire core_siphash_word_22_; 
wire core_siphash_word_23_; 
wire core_siphash_word_24_; 
wire core_siphash_word_25_; 
wire core_siphash_word_26_; 
wire core_siphash_word_27_; 
wire core_siphash_word_28_; 
wire core_siphash_word_29_; 
wire core_siphash_word_2_; 
wire core_siphash_word_30_; 
wire core_siphash_word_31_; 
wire core_siphash_word_32_; 
wire core_siphash_word_33_; 
wire core_siphash_word_34_; 
wire core_siphash_word_35_; 
wire core_siphash_word_36_; 
wire core_siphash_word_37_; 
wire core_siphash_word_38_; 
wire core_siphash_word_39_; 
wire core_siphash_word_3_; 
wire core_siphash_word_40_; 
wire core_siphash_word_41_; 
wire core_siphash_word_42_; 
wire core_siphash_word_43_; 
wire core_siphash_word_44_; 
wire core_siphash_word_45_; 
wire core_siphash_word_46_; 
wire core_siphash_word_47_; 
wire core_siphash_word_48_; 
wire core_siphash_word_49_; 
wire core_siphash_word_4_; 
wire core_siphash_word_50_; 
wire core_siphash_word_51_; 
wire core_siphash_word_52_; 
wire core_siphash_word_53_; 
wire core_siphash_word_54_; 
wire core_siphash_word_55_; 
wire core_siphash_word_56_; 
wire core_siphash_word_57_; 
wire core_siphash_word_58_; 
wire core_siphash_word_59_; 
wire core_siphash_word_5_; 
wire core_siphash_word_60_; 
wire core_siphash_word_61_; 
wire core_siphash_word_62_; 
wire core_siphash_word_63_; 
wire core_siphash_word_64_; 
wire core_siphash_word_65_; 
wire core_siphash_word_66_; 
wire core_siphash_word_67_; 
wire core_siphash_word_68_; 
wire core_siphash_word_69_; 
wire core_siphash_word_6_; 
wire core_siphash_word_70_; 
wire core_siphash_word_71_; 
wire core_siphash_word_72_; 
wire core_siphash_word_73_; 
wire core_siphash_word_74_; 
wire core_siphash_word_75_; 
wire core_siphash_word_76_; 
wire core_siphash_word_77_; 
wire core_siphash_word_78_; 
wire core_siphash_word_79_; 
wire core_siphash_word_7_; 
wire core_siphash_word_80_; 
wire core_siphash_word_81_; 
wire core_siphash_word_82_; 
wire core_siphash_word_83_; 
wire core_siphash_word_84_; 
wire core_siphash_word_85_; 
wire core_siphash_word_86_; 
wire core_siphash_word_87_; 
wire core_siphash_word_88_; 
wire core_siphash_word_89_; 
wire core_siphash_word_8_; 
wire core_siphash_word_90_; 
wire core_siphash_word_91_; 
wire core_siphash_word_92_; 
wire core_siphash_word_93_; 
wire core_siphash_word_94_; 
wire core_siphash_word_95_; 
wire core_siphash_word_96_; 
wire core_siphash_word_97_; 
wire core_siphash_word_98_; 
wire core_siphash_word_99_; 
wire core_siphash_word_9_; 
wire core_v0_reg_0_; 
wire core_v0_reg_10_; 
wire core_v0_reg_11_; 
wire core_v0_reg_12_; 
wire core_v0_reg_13_; 
wire core_v0_reg_14_; 
wire core_v0_reg_15_; 
wire core_v0_reg_16_; 
wire core_v0_reg_17_; 
wire core_v0_reg_18_; 
wire core_v0_reg_19_; 
wire core_v0_reg_1_; 
wire core_v0_reg_20_; 
wire core_v0_reg_21_; 
wire core_v0_reg_22_; 
wire core_v0_reg_23_; 
wire core_v0_reg_24_; 
wire core_v0_reg_25_; 
wire core_v0_reg_26_; 
wire core_v0_reg_27_; 
wire core_v0_reg_28_; 
wire core_v0_reg_29_; 
wire core_v0_reg_2_; 
wire core_v0_reg_30_; 
wire core_v0_reg_31_; 
wire core_v0_reg_32_; 
wire core_v0_reg_33_; 
wire core_v0_reg_34_; 
wire core_v0_reg_35_; 
wire core_v0_reg_36_; 
wire core_v0_reg_37_; 
wire core_v0_reg_38_; 
wire core_v0_reg_39_; 
wire core_v0_reg_3_; 
wire core_v0_reg_40_; 
wire core_v0_reg_41_; 
wire core_v0_reg_42_; 
wire core_v0_reg_43_; 
wire core_v0_reg_44_; 
wire core_v0_reg_45_; 
wire core_v0_reg_46_; 
wire core_v0_reg_47_; 
wire core_v0_reg_48_; 
wire core_v0_reg_49_; 
wire core_v0_reg_4_; 
wire core_v0_reg_50_; 
wire core_v0_reg_51_; 
wire core_v0_reg_52_; 
wire core_v0_reg_53_; 
wire core_v0_reg_54_; 
wire core_v0_reg_55_; 
wire core_v0_reg_56_; 
wire core_v0_reg_57_; 
wire core_v0_reg_58_; 
wire core_v0_reg_59_; 
wire core_v0_reg_5_; 
wire core_v0_reg_60_; 
wire core_v0_reg_61_; 
wire core_v0_reg_62_; 
wire core_v0_reg_63_; 
wire core_v0_reg_6_; 
wire core_v0_reg_7_; 
wire core_v0_reg_8_; 
wire core_v0_reg_9_; 
wire core_v1_reg_0_; 
wire core_v1_reg_10_; 
wire core_v1_reg_11_; 
wire core_v1_reg_12_; 
wire core_v1_reg_13_; 
wire core_v1_reg_14_; 
wire core_v1_reg_15_; 
wire core_v1_reg_16_; 
wire core_v1_reg_17_; 
wire core_v1_reg_18_; 
wire core_v1_reg_19_; 
wire core_v1_reg_1_; 
wire core_v1_reg_20_; 
wire core_v1_reg_21_; 
wire core_v1_reg_22_; 
wire core_v1_reg_23_; 
wire core_v1_reg_24_; 
wire core_v1_reg_25_; 
wire core_v1_reg_26_; 
wire core_v1_reg_27_; 
wire core_v1_reg_28_; 
wire core_v1_reg_29_; 
wire core_v1_reg_2_; 
wire core_v1_reg_30_; 
wire core_v1_reg_31_; 
wire core_v1_reg_32_; 
wire core_v1_reg_33_; 
wire core_v1_reg_34_; 
wire core_v1_reg_35_; 
wire core_v1_reg_36_; 
wire core_v1_reg_37_; 
wire core_v1_reg_38_; 
wire core_v1_reg_39_; 
wire core_v1_reg_3_; 
wire core_v1_reg_40_; 
wire core_v1_reg_41_; 
wire core_v1_reg_42_; 
wire core_v1_reg_43_; 
wire core_v1_reg_44_; 
wire core_v1_reg_45_; 
wire core_v1_reg_46_; 
wire core_v1_reg_47_; 
wire core_v1_reg_48_; 
wire core_v1_reg_49_; 
wire core_v1_reg_4_; 
wire core_v1_reg_50_; 
wire core_v1_reg_51_; 
wire core_v1_reg_52_; 
wire core_v1_reg_53_; 
wire core_v1_reg_54_; 
wire core_v1_reg_55_; 
wire core_v1_reg_56_; 
wire core_v1_reg_57_; 
wire core_v1_reg_58_; 
wire core_v1_reg_59_; 
wire core_v1_reg_5_; 
wire core_v1_reg_60_; 
wire core_v1_reg_61_; 
wire core_v1_reg_62_; 
wire core_v1_reg_63_; 
wire core_v1_reg_6_; 
wire core_v1_reg_7_; 
wire core_v1_reg_8_; 
wire core_v1_reg_9_; 
wire core_v2_reg_0_; 
wire core_v2_reg_10_; 
wire core_v2_reg_11_; 
wire core_v2_reg_12_; 
wire core_v2_reg_13_; 
wire core_v2_reg_14_; 
wire core_v2_reg_15_; 
wire core_v2_reg_16_; 
wire core_v2_reg_17_; 
wire core_v2_reg_18_; 
wire core_v2_reg_19_; 
wire core_v2_reg_1_; 
wire core_v2_reg_20_; 
wire core_v2_reg_21_; 
wire core_v2_reg_22_; 
wire core_v2_reg_23_; 
wire core_v2_reg_24_; 
wire core_v2_reg_25_; 
wire core_v2_reg_26_; 
wire core_v2_reg_27_; 
wire core_v2_reg_28_; 
wire core_v2_reg_29_; 
wire core_v2_reg_2_; 
wire core_v2_reg_30_; 
wire core_v2_reg_31_; 
wire core_v2_reg_32_; 
wire core_v2_reg_33_; 
wire core_v2_reg_34_; 
wire core_v2_reg_35_; 
wire core_v2_reg_36_; 
wire core_v2_reg_37_; 
wire core_v2_reg_38_; 
wire core_v2_reg_39_; 
wire core_v2_reg_3_; 
wire core_v2_reg_40_; 
wire core_v2_reg_41_; 
wire core_v2_reg_42_; 
wire core_v2_reg_43_; 
wire core_v2_reg_44_; 
wire core_v2_reg_45_; 
wire core_v2_reg_46_; 
wire core_v2_reg_47_; 
wire core_v2_reg_48_; 
wire core_v2_reg_49_; 
wire core_v2_reg_4_; 
wire core_v2_reg_50_; 
wire core_v2_reg_51_; 
wire core_v2_reg_52_; 
wire core_v2_reg_53_; 
wire core_v2_reg_54_; 
wire core_v2_reg_55_; 
wire core_v2_reg_56_; 
wire core_v2_reg_57_; 
wire core_v2_reg_58_; 
wire core_v2_reg_59_; 
wire core_v2_reg_5_; 
wire core_v2_reg_60_; 
wire core_v2_reg_61_; 
wire core_v2_reg_62_; 
wire core_v2_reg_63_; 
wire core_v2_reg_6_; 
wire core_v2_reg_7_; 
wire core_v2_reg_8_; 
wire core_v2_reg_9_; 
wire core_v3_reg_0_; 
wire core_v3_reg_10_; 
wire core_v3_reg_11_; 
wire core_v3_reg_12_; 
wire core_v3_reg_13_; 
wire core_v3_reg_14_; 
wire core_v3_reg_15_; 
wire core_v3_reg_16_; 
wire core_v3_reg_17_; 
wire core_v3_reg_18_; 
wire core_v3_reg_19_; 
wire core_v3_reg_1_; 
wire core_v3_reg_20_; 
wire core_v3_reg_21_; 
wire core_v3_reg_22_; 
wire core_v3_reg_23_; 
wire core_v3_reg_24_; 
wire core_v3_reg_25_; 
wire core_v3_reg_26_; 
wire core_v3_reg_27_; 
wire core_v3_reg_28_; 
wire core_v3_reg_29_; 
wire core_v3_reg_2_; 
wire core_v3_reg_30_; 
wire core_v3_reg_31_; 
wire core_v3_reg_32_; 
wire core_v3_reg_33_; 
wire core_v3_reg_34_; 
wire core_v3_reg_35_; 
wire core_v3_reg_36_; 
wire core_v3_reg_37_; 
wire core_v3_reg_38_; 
wire core_v3_reg_39_; 
wire core_v3_reg_3_; 
wire core_v3_reg_40_; 
wire core_v3_reg_41_; 
wire core_v3_reg_42_; 
wire core_v3_reg_43_; 
wire core_v3_reg_44_; 
wire core_v3_reg_45_; 
wire core_v3_reg_46_; 
wire core_v3_reg_47_; 
wire core_v3_reg_48_; 
wire core_v3_reg_49_; 
wire core_v3_reg_4_; 
wire core_v3_reg_50_; 
wire core_v3_reg_51_; 
wire core_v3_reg_52_; 
wire core_v3_reg_53_; 
wire core_v3_reg_54_; 
wire core_v3_reg_55_; 
wire core_v3_reg_56_; 
wire core_v3_reg_57_; 
wire core_v3_reg_58_; 
wire core_v3_reg_59_; 
wire core_v3_reg_5_; 
wire core_v3_reg_60_; 
wire core_v3_reg_61_; 
wire core_v3_reg_62_; 
wire core_v3_reg_63_; 
wire core_v3_reg_6_; 
wire core_v3_reg_7_; 
wire core_v3_reg_8_; 
wire core_v3_reg_9_; 
input cs;
output \read_data[0] ;
output \read_data[10] ;
output \read_data[11] ;
output \read_data[12] ;
output \read_data[13] ;
output \read_data[14] ;
output \read_data[15] ;
output \read_data[16] ;
output \read_data[17] ;
output \read_data[18] ;
output \read_data[19] ;
output \read_data[1] ;
output \read_data[20] ;
output \read_data[21] ;
output \read_data[22] ;
output \read_data[23] ;
output \read_data[24] ;
output \read_data[25] ;
output \read_data[26] ;
output \read_data[27] ;
output \read_data[28] ;
output \read_data[29] ;
output \read_data[2] ;
output \read_data[30] ;
output \read_data[31] ;
output \read_data[3] ;
output \read_data[4] ;
output \read_data[5] ;
output \read_data[6] ;
output \read_data[7] ;
output \read_data[8] ;
output \read_data[9] ;
input reset_n;
input we;
wire word0_reg_0_; 
wire word0_reg_10_; 
wire word0_reg_11_; 
wire word0_reg_12_; 
wire word0_reg_13_; 
wire word0_reg_14_; 
wire word0_reg_15_; 
wire word0_reg_16_; 
wire word0_reg_17_; 
wire word0_reg_18_; 
wire word0_reg_19_; 
wire word0_reg_1_; 
wire word0_reg_20_; 
wire word0_reg_21_; 
wire word0_reg_22_; 
wire word0_reg_23_; 
wire word0_reg_24_; 
wire word0_reg_25_; 
wire word0_reg_26_; 
wire word0_reg_27_; 
wire word0_reg_28_; 
wire word0_reg_29_; 
wire word0_reg_2_; 
wire word0_reg_30_; 
wire word0_reg_31_; 
wire word0_reg_3_; 
wire word0_reg_4_; 
wire word0_reg_5_; 
wire word0_reg_6_; 
wire word0_reg_7_; 
wire word0_reg_8_; 
wire word0_reg_9_; 
wire word1_reg_0_; 
wire word1_reg_10_; 
wire word1_reg_11_; 
wire word1_reg_12_; 
wire word1_reg_13_; 
wire word1_reg_14_; 
wire word1_reg_15_; 
wire word1_reg_16_; 
wire word1_reg_17_; 
wire word1_reg_18_; 
wire word1_reg_19_; 
wire word1_reg_1_; 
wire word1_reg_20_; 
wire word1_reg_21_; 
wire word1_reg_22_; 
wire word1_reg_23_; 
wire word1_reg_24_; 
wire word1_reg_25_; 
wire word1_reg_26_; 
wire word1_reg_27_; 
wire word1_reg_28_; 
wire word1_reg_29_; 
wire word1_reg_2_; 
wire word1_reg_30_; 
wire word1_reg_31_; 
wire word1_reg_3_; 
wire word1_reg_4_; 
wire word1_reg_5_; 
wire word1_reg_6_; 
wire word1_reg_7_; 
wire word1_reg_8_; 
wire word1_reg_9_; 
wire word2_reg_0_; 
wire word2_reg_10_; 
wire word2_reg_11_; 
wire word2_reg_12_; 
wire word2_reg_13_; 
wire word2_reg_14_; 
wire word2_reg_15_; 
wire word2_reg_16_; 
wire word2_reg_17_; 
wire word2_reg_18_; 
wire word2_reg_19_; 
wire word2_reg_1_; 
wire word2_reg_20_; 
wire word2_reg_21_; 
wire word2_reg_22_; 
wire word2_reg_23_; 
wire word2_reg_24_; 
wire word2_reg_25_; 
wire word2_reg_26_; 
wire word2_reg_27_; 
wire word2_reg_28_; 
wire word2_reg_29_; 
wire word2_reg_2_; 
wire word2_reg_30_; 
wire word2_reg_31_; 
wire word2_reg_3_; 
wire word2_reg_4_; 
wire word2_reg_5_; 
wire word2_reg_6_; 
wire word2_reg_7_; 
wire word2_reg_8_; 
wire word2_reg_9_; 
wire word3_reg_0_; 
wire word3_reg_10_; 
wire word3_reg_11_; 
wire word3_reg_12_; 
wire word3_reg_13_; 
wire word3_reg_14_; 
wire word3_reg_15_; 
wire word3_reg_16_; 
wire word3_reg_17_; 
wire word3_reg_18_; 
wire word3_reg_19_; 
wire word3_reg_1_; 
wire word3_reg_20_; 
wire word3_reg_21_; 
wire word3_reg_22_; 
wire word3_reg_23_; 
wire word3_reg_24_; 
wire word3_reg_25_; 
wire word3_reg_26_; 
wire word3_reg_27_; 
wire word3_reg_28_; 
wire word3_reg_29_; 
wire word3_reg_2_; 
wire word3_reg_30_; 
wire word3_reg_31_; 
wire word3_reg_3_; 
wire word3_reg_4_; 
wire word3_reg_5_; 
wire word3_reg_6_; 
wire word3_reg_7_; 
wire word3_reg_8_; 
wire word3_reg_9_; 
input \write_data[0] ;
input \write_data[10] ;
input \write_data[11] ;
input \write_data[12] ;
input \write_data[13] ;
input \write_data[14] ;
input \write_data[15] ;
input \write_data[16] ;
input \write_data[17] ;
input \write_data[18] ;
input \write_data[19] ;
input \write_data[1] ;
input \write_data[20] ;
input \write_data[21] ;
input \write_data[22] ;
input \write_data[23] ;
input \write_data[24] ;
input \write_data[25] ;
input \write_data[26] ;
input \write_data[27] ;
input \write_data[28] ;
input \write_data[29] ;
input \write_data[2] ;
input \write_data[30] ;
input \write_data[31] ;
input \write_data[3] ;
input \write_data[4] ;
input \write_data[5] ;
input \write_data[6] ;
input \write_data[7] ;
input \write_data[8] ;
input \write_data[9] ;
AND2X2 AND2X2_1 ( .A(_abc_19873_new_n870_), .B(_abc_19873_new_n871_), .Y(_abc_19873_new_n872_));
AND2X2 AND2X2_10 ( .A(_abc_19873_new_n878_), .B(\addr[3] ), .Y(_abc_19873_new_n886_));
AND2X2 AND2X2_100 ( .A(_abc_19873_new_n916_), .B(core_key_68_), .Y(_abc_19873_new_n1031_));
AND2X2 AND2X2_1000 ( .A(_abc_19873_new_n2503_), .B(_abc_19873_new_n2500_), .Y(_0key3_reg_31_0__5_));
AND2X2 AND2X2_1001 ( .A(_abc_19873_new_n2474_), .B(_abc_19873_new_n2158_), .Y(_abc_19873_new_n2506_));
AND2X2 AND2X2_1002 ( .A(_abc_19873_new_n2507_), .B(reset_n), .Y(_abc_19873_new_n2508_));
AND2X2 AND2X2_1003 ( .A(_abc_19873_new_n2508_), .B(_abc_19873_new_n2505_), .Y(_0key3_reg_31_0__6_));
AND2X2 AND2X2_1004 ( .A(_abc_19873_new_n2474_), .B(_abc_19873_new_n2164_), .Y(_abc_19873_new_n2511_));
AND2X2 AND2X2_1005 ( .A(_abc_19873_new_n2512_), .B(reset_n), .Y(_abc_19873_new_n2513_));
AND2X2 AND2X2_1006 ( .A(_abc_19873_new_n2513_), .B(_abc_19873_new_n2510_), .Y(_0key3_reg_31_0__7_));
AND2X2 AND2X2_1007 ( .A(_abc_19873_new_n2474_), .B(_abc_19873_new_n2170_), .Y(_abc_19873_new_n2516_));
AND2X2 AND2X2_1008 ( .A(_abc_19873_new_n2517_), .B(reset_n), .Y(_abc_19873_new_n2518_));
AND2X2 AND2X2_1009 ( .A(_abc_19873_new_n2518_), .B(_abc_19873_new_n2515_), .Y(_0key3_reg_31_0__8_));
AND2X2 AND2X2_101 ( .A(_abc_19873_new_n1035_), .B(_abc_19873_new_n937_), .Y(\read_data[4] ));
AND2X2 AND2X2_1010 ( .A(_abc_19873_new_n2474_), .B(_abc_19873_new_n2176_), .Y(_abc_19873_new_n2521_));
AND2X2 AND2X2_1011 ( .A(_abc_19873_new_n2522_), .B(reset_n), .Y(_abc_19873_new_n2523_));
AND2X2 AND2X2_1012 ( .A(_abc_19873_new_n2523_), .B(_abc_19873_new_n2520_), .Y(_0key3_reg_31_0__9_));
AND2X2 AND2X2_1013 ( .A(_abc_19873_new_n2474_), .B(_abc_19873_new_n2182_), .Y(_abc_19873_new_n2526_));
AND2X2 AND2X2_1014 ( .A(_abc_19873_new_n2527_), .B(reset_n), .Y(_abc_19873_new_n2528_));
AND2X2 AND2X2_1015 ( .A(_abc_19873_new_n2528_), .B(_abc_19873_new_n2525_), .Y(_0key3_reg_31_0__10_));
AND2X2 AND2X2_1016 ( .A(_abc_19873_new_n2474_), .B(_abc_19873_new_n2188_), .Y(_abc_19873_new_n2531_));
AND2X2 AND2X2_1017 ( .A(_abc_19873_new_n2532_), .B(reset_n), .Y(_abc_19873_new_n2533_));
AND2X2 AND2X2_1018 ( .A(_abc_19873_new_n2533_), .B(_abc_19873_new_n2530_), .Y(_0key3_reg_31_0__11_));
AND2X2 AND2X2_1019 ( .A(_abc_19873_new_n2474_), .B(_abc_19873_new_n2194_), .Y(_abc_19873_new_n2536_));
AND2X2 AND2X2_102 ( .A(_abc_19873_new_n893_), .B(_abc_19873_new_n904_), .Y(_abc_19873_new_n1037_));
AND2X2 AND2X2_1020 ( .A(_abc_19873_new_n2537_), .B(reset_n), .Y(_abc_19873_new_n2538_));
AND2X2 AND2X2_1021 ( .A(_abc_19873_new_n2538_), .B(_abc_19873_new_n2535_), .Y(_0key3_reg_31_0__12_));
AND2X2 AND2X2_1022 ( .A(_abc_19873_new_n2474_), .B(_abc_19873_new_n2200_), .Y(_abc_19873_new_n2541_));
AND2X2 AND2X2_1023 ( .A(_abc_19873_new_n2542_), .B(reset_n), .Y(_abc_19873_new_n2543_));
AND2X2 AND2X2_1024 ( .A(_abc_19873_new_n2543_), .B(_abc_19873_new_n2540_), .Y(_0key3_reg_31_0__13_));
AND2X2 AND2X2_1025 ( .A(_abc_19873_new_n2474_), .B(_abc_19873_new_n2206_), .Y(_abc_19873_new_n2546_));
AND2X2 AND2X2_1026 ( .A(_abc_19873_new_n2547_), .B(reset_n), .Y(_abc_19873_new_n2548_));
AND2X2 AND2X2_1027 ( .A(_abc_19873_new_n2548_), .B(_abc_19873_new_n2545_), .Y(_0key3_reg_31_0__14_));
AND2X2 AND2X2_1028 ( .A(_abc_19873_new_n2474_), .B(_abc_19873_new_n2212_), .Y(_abc_19873_new_n2551_));
AND2X2 AND2X2_1029 ( .A(_abc_19873_new_n2552_), .B(reset_n), .Y(_abc_19873_new_n2553_));
AND2X2 AND2X2_103 ( .A(_abc_19873_new_n897_), .B(core_final_rounds_1_), .Y(_abc_19873_new_n1040_));
AND2X2 AND2X2_1030 ( .A(_abc_19873_new_n2553_), .B(_abc_19873_new_n2550_), .Y(_0key3_reg_31_0__15_));
AND2X2 AND2X2_1031 ( .A(_abc_19873_new_n2474_), .B(_abc_19873_new_n2218_), .Y(_abc_19873_new_n2556_));
AND2X2 AND2X2_1032 ( .A(_abc_19873_new_n2557_), .B(reset_n), .Y(_abc_19873_new_n2558_));
AND2X2 AND2X2_1033 ( .A(_abc_19873_new_n2558_), .B(_abc_19873_new_n2555_), .Y(_0key3_reg_31_0__16_));
AND2X2 AND2X2_1034 ( .A(_abc_19873_new_n2474_), .B(_abc_19873_new_n2224_), .Y(_abc_19873_new_n2561_));
AND2X2 AND2X2_1035 ( .A(_abc_19873_new_n2562_), .B(reset_n), .Y(_abc_19873_new_n2563_));
AND2X2 AND2X2_1036 ( .A(_abc_19873_new_n2563_), .B(_abc_19873_new_n2560_), .Y(_0key3_reg_31_0__17_));
AND2X2 AND2X2_1037 ( .A(_abc_19873_new_n2474_), .B(_abc_19873_new_n2230_), .Y(_abc_19873_new_n2566_));
AND2X2 AND2X2_1038 ( .A(_abc_19873_new_n2567_), .B(reset_n), .Y(_abc_19873_new_n2568_));
AND2X2 AND2X2_1039 ( .A(_abc_19873_new_n2568_), .B(_abc_19873_new_n2565_), .Y(_0key3_reg_31_0__18_));
AND2X2 AND2X2_104 ( .A(_abc_19873_new_n916_), .B(core_key_69_), .Y(_abc_19873_new_n1041_));
AND2X2 AND2X2_1040 ( .A(_abc_19873_new_n2474_), .B(_abc_19873_new_n2236_), .Y(_abc_19873_new_n2571_));
AND2X2 AND2X2_1041 ( .A(_abc_19873_new_n2572_), .B(reset_n), .Y(_abc_19873_new_n2573_));
AND2X2 AND2X2_1042 ( .A(_abc_19873_new_n2573_), .B(_abc_19873_new_n2570_), .Y(_0key3_reg_31_0__19_));
AND2X2 AND2X2_1043 ( .A(_abc_19873_new_n2474_), .B(_abc_19873_new_n2242_), .Y(_abc_19873_new_n2576_));
AND2X2 AND2X2_1044 ( .A(_abc_19873_new_n2577_), .B(reset_n), .Y(_abc_19873_new_n2578_));
AND2X2 AND2X2_1045 ( .A(_abc_19873_new_n2578_), .B(_abc_19873_new_n2575_), .Y(_0key3_reg_31_0__20_));
AND2X2 AND2X2_1046 ( .A(_abc_19873_new_n2474_), .B(_abc_19873_new_n2248_), .Y(_abc_19873_new_n2581_));
AND2X2 AND2X2_1047 ( .A(_abc_19873_new_n2582_), .B(reset_n), .Y(_abc_19873_new_n2583_));
AND2X2 AND2X2_1048 ( .A(_abc_19873_new_n2583_), .B(_abc_19873_new_n2580_), .Y(_0key3_reg_31_0__21_));
AND2X2 AND2X2_1049 ( .A(_abc_19873_new_n2474_), .B(_abc_19873_new_n2254_), .Y(_abc_19873_new_n2586_));
AND2X2 AND2X2_105 ( .A(_abc_19873_new_n925_), .B(word2_reg_5_), .Y(_abc_19873_new_n1044_));
AND2X2 AND2X2_1050 ( .A(_abc_19873_new_n2587_), .B(reset_n), .Y(_abc_19873_new_n2588_));
AND2X2 AND2X2_1051 ( .A(_abc_19873_new_n2588_), .B(_abc_19873_new_n2585_), .Y(_0key3_reg_31_0__22_));
AND2X2 AND2X2_1052 ( .A(_abc_19873_new_n2474_), .B(_abc_19873_new_n2260_), .Y(_abc_19873_new_n2591_));
AND2X2 AND2X2_1053 ( .A(_abc_19873_new_n2592_), .B(reset_n), .Y(_abc_19873_new_n2593_));
AND2X2 AND2X2_1054 ( .A(_abc_19873_new_n2593_), .B(_abc_19873_new_n2590_), .Y(_0key3_reg_31_0__23_));
AND2X2 AND2X2_1055 ( .A(_abc_19873_new_n2474_), .B(_abc_19873_new_n2266_), .Y(_abc_19873_new_n2596_));
AND2X2 AND2X2_1056 ( .A(_abc_19873_new_n2597_), .B(reset_n), .Y(_abc_19873_new_n2598_));
AND2X2 AND2X2_1057 ( .A(_abc_19873_new_n2598_), .B(_abc_19873_new_n2595_), .Y(_0key3_reg_31_0__24_));
AND2X2 AND2X2_1058 ( .A(_abc_19873_new_n2474_), .B(_abc_19873_new_n2272_), .Y(_abc_19873_new_n2601_));
AND2X2 AND2X2_1059 ( .A(_abc_19873_new_n2602_), .B(reset_n), .Y(_abc_19873_new_n2603_));
AND2X2 AND2X2_106 ( .A(_abc_19873_new_n919_), .B(core_mi_37_), .Y(_abc_19873_new_n1045_));
AND2X2 AND2X2_1060 ( .A(_abc_19873_new_n2603_), .B(_abc_19873_new_n2600_), .Y(_0key3_reg_31_0__25_));
AND2X2 AND2X2_1061 ( .A(_abc_19873_new_n2474_), .B(_abc_19873_new_n2278_), .Y(_abc_19873_new_n2606_));
AND2X2 AND2X2_1062 ( .A(_abc_19873_new_n2607_), .B(reset_n), .Y(_abc_19873_new_n2608_));
AND2X2 AND2X2_1063 ( .A(_abc_19873_new_n2608_), .B(_abc_19873_new_n2605_), .Y(_0key3_reg_31_0__26_));
AND2X2 AND2X2_1064 ( .A(_abc_19873_new_n2474_), .B(_abc_19873_new_n2284_), .Y(_abc_19873_new_n2611_));
AND2X2 AND2X2_1065 ( .A(_abc_19873_new_n2612_), .B(reset_n), .Y(_abc_19873_new_n2613_));
AND2X2 AND2X2_1066 ( .A(_abc_19873_new_n2613_), .B(_abc_19873_new_n2610_), .Y(_0key3_reg_31_0__27_));
AND2X2 AND2X2_1067 ( .A(_abc_19873_new_n2474_), .B(_abc_19873_new_n2290_), .Y(_abc_19873_new_n2616_));
AND2X2 AND2X2_1068 ( .A(_abc_19873_new_n2617_), .B(reset_n), .Y(_abc_19873_new_n2618_));
AND2X2 AND2X2_1069 ( .A(_abc_19873_new_n2618_), .B(_abc_19873_new_n2615_), .Y(_0key3_reg_31_0__28_));
AND2X2 AND2X2_107 ( .A(_abc_19873_new_n930_), .B(word0_reg_5_), .Y(_abc_19873_new_n1046_));
AND2X2 AND2X2_1070 ( .A(_abc_19873_new_n2474_), .B(_abc_19873_new_n2296_), .Y(_abc_19873_new_n2621_));
AND2X2 AND2X2_1071 ( .A(_abc_19873_new_n2622_), .B(reset_n), .Y(_abc_19873_new_n2623_));
AND2X2 AND2X2_1072 ( .A(_abc_19873_new_n2623_), .B(_abc_19873_new_n2620_), .Y(_0key3_reg_31_0__29_));
AND2X2 AND2X2_1073 ( .A(_abc_19873_new_n2474_), .B(_abc_19873_new_n2302_), .Y(_abc_19873_new_n2626_));
AND2X2 AND2X2_1074 ( .A(_abc_19873_new_n2627_), .B(reset_n), .Y(_abc_19873_new_n2628_));
AND2X2 AND2X2_1075 ( .A(_abc_19873_new_n2628_), .B(_abc_19873_new_n2625_), .Y(_0key3_reg_31_0__30_));
AND2X2 AND2X2_1076 ( .A(_abc_19873_new_n2474_), .B(_abc_19873_new_n2308_), .Y(_abc_19873_new_n2631_));
AND2X2 AND2X2_1077 ( .A(_abc_19873_new_n2632_), .B(reset_n), .Y(_abc_19873_new_n2633_));
AND2X2 AND2X2_1078 ( .A(_abc_19873_new_n2633_), .B(_abc_19873_new_n2630_), .Y(_0key3_reg_31_0__31_));
AND2X2 AND2X2_1079 ( .A(_abc_19873_new_n916_), .B(_abc_19873_new_n2119_), .Y(_abc_19873_new_n2635_));
AND2X2 AND2X2_108 ( .A(_abc_19873_new_n928_), .B(core_key_37_), .Y(_abc_19873_new_n1050_));
AND2X2 AND2X2_1080 ( .A(_abc_19873_new_n2635_), .B(_abc_19873_new_n2122_), .Y(_abc_19873_new_n2637_));
AND2X2 AND2X2_1081 ( .A(_abc_19873_new_n2638_), .B(_abc_19873_new_n2636_), .Y(_abc_19873_new_n2639_));
AND2X2 AND2X2_1082 ( .A(_abc_19873_new_n2639_), .B(reset_n), .Y(_0key2_reg_31_0__0_));
AND2X2 AND2X2_1083 ( .A(_abc_19873_new_n2635_), .B(_abc_19873_new_n2128_), .Y(_abc_19873_new_n2642_));
AND2X2 AND2X2_1084 ( .A(_abc_19873_new_n2643_), .B(_abc_19873_new_n2641_), .Y(_abc_19873_new_n2644_));
AND2X2 AND2X2_1085 ( .A(_abc_19873_new_n2644_), .B(reset_n), .Y(_0key2_reg_31_0__1_));
AND2X2 AND2X2_1086 ( .A(_abc_19873_new_n2635_), .B(_abc_19873_new_n2134_), .Y(_abc_19873_new_n2647_));
AND2X2 AND2X2_1087 ( .A(_abc_19873_new_n2648_), .B(_abc_19873_new_n2646_), .Y(_abc_19873_new_n2649_));
AND2X2 AND2X2_1088 ( .A(_abc_19873_new_n2649_), .B(reset_n), .Y(_0key2_reg_31_0__2_));
AND2X2 AND2X2_1089 ( .A(_abc_19873_new_n2635_), .B(_abc_19873_new_n2140_), .Y(_abc_19873_new_n2652_));
AND2X2 AND2X2_109 ( .A(_abc_19873_new_n901_), .B(core_key_5_), .Y(_abc_19873_new_n1051_));
AND2X2 AND2X2_1090 ( .A(_abc_19873_new_n2653_), .B(_abc_19873_new_n2651_), .Y(_abc_19873_new_n2654_));
AND2X2 AND2X2_1091 ( .A(_abc_19873_new_n2654_), .B(reset_n), .Y(_0key2_reg_31_0__3_));
AND2X2 AND2X2_1092 ( .A(_abc_19873_new_n2635_), .B(_abc_19873_new_n2146_), .Y(_abc_19873_new_n2657_));
AND2X2 AND2X2_1093 ( .A(_abc_19873_new_n2658_), .B(_abc_19873_new_n2656_), .Y(_abc_19873_new_n2659_));
AND2X2 AND2X2_1094 ( .A(_abc_19873_new_n2659_), .B(reset_n), .Y(_0key2_reg_31_0__4_));
AND2X2 AND2X2_1095 ( .A(_abc_19873_new_n2635_), .B(_abc_19873_new_n2152_), .Y(_abc_19873_new_n2662_));
AND2X2 AND2X2_1096 ( .A(_abc_19873_new_n2663_), .B(_abc_19873_new_n2661_), .Y(_abc_19873_new_n2664_));
AND2X2 AND2X2_1097 ( .A(_abc_19873_new_n2664_), .B(reset_n), .Y(_0key2_reg_31_0__5_));
AND2X2 AND2X2_1098 ( .A(_abc_19873_new_n2635_), .B(_abc_19873_new_n2158_), .Y(_abc_19873_new_n2667_));
AND2X2 AND2X2_1099 ( .A(_abc_19873_new_n2668_), .B(_abc_19873_new_n2666_), .Y(_abc_19873_new_n2669_));
AND2X2 AND2X2_11 ( .A(_abc_19873_new_n885_), .B(_abc_19873_new_n886_), .Y(_abc_19873_new_n887_));
AND2X2 AND2X2_110 ( .A(_abc_19873_new_n881_), .B(core_key_101_), .Y(_abc_19873_new_n1053_));
AND2X2 AND2X2_1100 ( .A(_abc_19873_new_n2669_), .B(reset_n), .Y(_0key2_reg_31_0__6_));
AND2X2 AND2X2_1101 ( .A(_abc_19873_new_n2635_), .B(_abc_19873_new_n2164_), .Y(_abc_19873_new_n2672_));
AND2X2 AND2X2_1102 ( .A(_abc_19873_new_n2673_), .B(_abc_19873_new_n2671_), .Y(_abc_19873_new_n2674_));
AND2X2 AND2X2_1103 ( .A(_abc_19873_new_n2674_), .B(reset_n), .Y(_0key2_reg_31_0__7_));
AND2X2 AND2X2_1104 ( .A(_abc_19873_new_n2635_), .B(_abc_19873_new_n2170_), .Y(_abc_19873_new_n2677_));
AND2X2 AND2X2_1105 ( .A(_abc_19873_new_n2678_), .B(_abc_19873_new_n2676_), .Y(_abc_19873_new_n2679_));
AND2X2 AND2X2_1106 ( .A(_abc_19873_new_n2679_), .B(reset_n), .Y(_0key2_reg_31_0__8_));
AND2X2 AND2X2_1107 ( .A(_abc_19873_new_n2635_), .B(_abc_19873_new_n2176_), .Y(_abc_19873_new_n2682_));
AND2X2 AND2X2_1108 ( .A(_abc_19873_new_n2683_), .B(_abc_19873_new_n2681_), .Y(_abc_19873_new_n2684_));
AND2X2 AND2X2_1109 ( .A(_abc_19873_new_n2684_), .B(reset_n), .Y(_0key2_reg_31_0__9_));
AND2X2 AND2X2_111 ( .A(_abc_19873_new_n888_), .B(core_mi_5_), .Y(_abc_19873_new_n1054_));
AND2X2 AND2X2_1110 ( .A(_abc_19873_new_n2635_), .B(_abc_19873_new_n2182_), .Y(_abc_19873_new_n2687_));
AND2X2 AND2X2_1111 ( .A(_abc_19873_new_n2688_), .B(_abc_19873_new_n2686_), .Y(_abc_19873_new_n2689_));
AND2X2 AND2X2_1112 ( .A(_abc_19873_new_n2689_), .B(reset_n), .Y(_0key2_reg_31_0__10_));
AND2X2 AND2X2_1113 ( .A(_abc_19873_new_n2635_), .B(_abc_19873_new_n2188_), .Y(_abc_19873_new_n2692_));
AND2X2 AND2X2_1114 ( .A(_abc_19873_new_n2693_), .B(_abc_19873_new_n2691_), .Y(_abc_19873_new_n2694_));
AND2X2 AND2X2_1115 ( .A(_abc_19873_new_n2694_), .B(reset_n), .Y(_0key2_reg_31_0__11_));
AND2X2 AND2X2_1116 ( .A(_abc_19873_new_n2635_), .B(_abc_19873_new_n2194_), .Y(_abc_19873_new_n2697_));
AND2X2 AND2X2_1117 ( .A(_abc_19873_new_n2698_), .B(_abc_19873_new_n2696_), .Y(_abc_19873_new_n2699_));
AND2X2 AND2X2_1118 ( .A(_abc_19873_new_n2699_), .B(reset_n), .Y(_0key2_reg_31_0__12_));
AND2X2 AND2X2_1119 ( .A(_abc_19873_new_n2635_), .B(_abc_19873_new_n2200_), .Y(_abc_19873_new_n2702_));
AND2X2 AND2X2_112 ( .A(_abc_19873_new_n907_), .B(word1_reg_5_), .Y(_abc_19873_new_n1056_));
AND2X2 AND2X2_1120 ( .A(_abc_19873_new_n2703_), .B(_abc_19873_new_n2701_), .Y(_abc_19873_new_n2704_));
AND2X2 AND2X2_1121 ( .A(_abc_19873_new_n2704_), .B(reset_n), .Y(_0key2_reg_31_0__13_));
AND2X2 AND2X2_1122 ( .A(_abc_19873_new_n2635_), .B(_abc_19873_new_n2206_), .Y(_abc_19873_new_n2707_));
AND2X2 AND2X2_1123 ( .A(_abc_19873_new_n2708_), .B(_abc_19873_new_n2706_), .Y(_abc_19873_new_n2709_));
AND2X2 AND2X2_1124 ( .A(_abc_19873_new_n2709_), .B(reset_n), .Y(_0key2_reg_31_0__14_));
AND2X2 AND2X2_1125 ( .A(_abc_19873_new_n2635_), .B(_abc_19873_new_n2212_), .Y(_abc_19873_new_n2712_));
AND2X2 AND2X2_1126 ( .A(_abc_19873_new_n2713_), .B(_abc_19873_new_n2711_), .Y(_abc_19873_new_n2714_));
AND2X2 AND2X2_1127 ( .A(_abc_19873_new_n2714_), .B(reset_n), .Y(_0key2_reg_31_0__15_));
AND2X2 AND2X2_1128 ( .A(_abc_19873_new_n2635_), .B(_abc_19873_new_n2218_), .Y(_abc_19873_new_n2717_));
AND2X2 AND2X2_1129 ( .A(_abc_19873_new_n2718_), .B(_abc_19873_new_n2716_), .Y(_abc_19873_new_n2719_));
AND2X2 AND2X2_113 ( .A(_abc_19873_new_n912_), .B(word3_reg_5_), .Y(_abc_19873_new_n1057_));
AND2X2 AND2X2_1130 ( .A(_abc_19873_new_n2719_), .B(reset_n), .Y(_0key2_reg_31_0__16_));
AND2X2 AND2X2_1131 ( .A(_abc_19873_new_n2635_), .B(_abc_19873_new_n2224_), .Y(_abc_19873_new_n2722_));
AND2X2 AND2X2_1132 ( .A(_abc_19873_new_n2723_), .B(_abc_19873_new_n2721_), .Y(_abc_19873_new_n2724_));
AND2X2 AND2X2_1133 ( .A(_abc_19873_new_n2724_), .B(reset_n), .Y(_0key2_reg_31_0__17_));
AND2X2 AND2X2_1134 ( .A(_abc_19873_new_n2635_), .B(_abc_19873_new_n2230_), .Y(_abc_19873_new_n2727_));
AND2X2 AND2X2_1135 ( .A(_abc_19873_new_n2728_), .B(_abc_19873_new_n2726_), .Y(_abc_19873_new_n2729_));
AND2X2 AND2X2_1136 ( .A(_abc_19873_new_n2729_), .B(reset_n), .Y(_0key2_reg_31_0__18_));
AND2X2 AND2X2_1137 ( .A(_abc_19873_new_n2635_), .B(_abc_19873_new_n2236_), .Y(_abc_19873_new_n2732_));
AND2X2 AND2X2_1138 ( .A(_abc_19873_new_n2733_), .B(_abc_19873_new_n2731_), .Y(_abc_19873_new_n2734_));
AND2X2 AND2X2_1139 ( .A(_abc_19873_new_n2734_), .B(reset_n), .Y(_0key2_reg_31_0__19_));
AND2X2 AND2X2_114 ( .A(_abc_19873_new_n1061_), .B(_abc_19873_new_n937_), .Y(\read_data[5] ));
AND2X2 AND2X2_1140 ( .A(_abc_19873_new_n2635_), .B(_abc_19873_new_n2242_), .Y(_abc_19873_new_n2737_));
AND2X2 AND2X2_1141 ( .A(_abc_19873_new_n2738_), .B(_abc_19873_new_n2736_), .Y(_abc_19873_new_n2739_));
AND2X2 AND2X2_1142 ( .A(_abc_19873_new_n2739_), .B(reset_n), .Y(_0key2_reg_31_0__20_));
AND2X2 AND2X2_1143 ( .A(_abc_19873_new_n2635_), .B(_abc_19873_new_n2248_), .Y(_abc_19873_new_n2742_));
AND2X2 AND2X2_1144 ( .A(_abc_19873_new_n2743_), .B(_abc_19873_new_n2741_), .Y(_abc_19873_new_n2744_));
AND2X2 AND2X2_1145 ( .A(_abc_19873_new_n2744_), .B(reset_n), .Y(_0key2_reg_31_0__21_));
AND2X2 AND2X2_1146 ( .A(_abc_19873_new_n2635_), .B(_abc_19873_new_n2254_), .Y(_abc_19873_new_n2747_));
AND2X2 AND2X2_1147 ( .A(_abc_19873_new_n2748_), .B(_abc_19873_new_n2746_), .Y(_abc_19873_new_n2749_));
AND2X2 AND2X2_1148 ( .A(_abc_19873_new_n2749_), .B(reset_n), .Y(_0key2_reg_31_0__22_));
AND2X2 AND2X2_1149 ( .A(_abc_19873_new_n2635_), .B(_abc_19873_new_n2260_), .Y(_abc_19873_new_n2752_));
AND2X2 AND2X2_115 ( .A(_abc_19873_new_n897_), .B(core_final_rounds_2_), .Y(_abc_19873_new_n1063_));
AND2X2 AND2X2_1150 ( .A(_abc_19873_new_n2753_), .B(_abc_19873_new_n2751_), .Y(_abc_19873_new_n2754_));
AND2X2 AND2X2_1151 ( .A(_abc_19873_new_n2754_), .B(reset_n), .Y(_0key2_reg_31_0__23_));
AND2X2 AND2X2_1152 ( .A(_abc_19873_new_n2635_), .B(_abc_19873_new_n2266_), .Y(_abc_19873_new_n2757_));
AND2X2 AND2X2_1153 ( .A(_abc_19873_new_n2758_), .B(_abc_19873_new_n2756_), .Y(_abc_19873_new_n2759_));
AND2X2 AND2X2_1154 ( .A(_abc_19873_new_n2759_), .B(reset_n), .Y(_0key2_reg_31_0__24_));
AND2X2 AND2X2_1155 ( .A(_abc_19873_new_n2635_), .B(_abc_19873_new_n2272_), .Y(_abc_19873_new_n2762_));
AND2X2 AND2X2_1156 ( .A(_abc_19873_new_n2763_), .B(_abc_19873_new_n2761_), .Y(_abc_19873_new_n2764_));
AND2X2 AND2X2_1157 ( .A(_abc_19873_new_n2764_), .B(reset_n), .Y(_0key2_reg_31_0__25_));
AND2X2 AND2X2_1158 ( .A(_abc_19873_new_n2635_), .B(_abc_19873_new_n2278_), .Y(_abc_19873_new_n2767_));
AND2X2 AND2X2_1159 ( .A(_abc_19873_new_n2768_), .B(_abc_19873_new_n2766_), .Y(_abc_19873_new_n2769_));
AND2X2 AND2X2_116 ( .A(_abc_19873_new_n919_), .B(core_mi_38_), .Y(_abc_19873_new_n1064_));
AND2X2 AND2X2_1160 ( .A(_abc_19873_new_n2769_), .B(reset_n), .Y(_0key2_reg_31_0__26_));
AND2X2 AND2X2_1161 ( .A(_abc_19873_new_n2635_), .B(_abc_19873_new_n2284_), .Y(_abc_19873_new_n2772_));
AND2X2 AND2X2_1162 ( .A(_abc_19873_new_n2773_), .B(_abc_19873_new_n2771_), .Y(_abc_19873_new_n2774_));
AND2X2 AND2X2_1163 ( .A(_abc_19873_new_n2774_), .B(reset_n), .Y(_0key2_reg_31_0__27_));
AND2X2 AND2X2_1164 ( .A(_abc_19873_new_n2635_), .B(_abc_19873_new_n2290_), .Y(_abc_19873_new_n2777_));
AND2X2 AND2X2_1165 ( .A(_abc_19873_new_n2778_), .B(_abc_19873_new_n2776_), .Y(_abc_19873_new_n2779_));
AND2X2 AND2X2_1166 ( .A(_abc_19873_new_n2779_), .B(reset_n), .Y(_0key2_reg_31_0__28_));
AND2X2 AND2X2_1167 ( .A(_abc_19873_new_n2635_), .B(_abc_19873_new_n2296_), .Y(_abc_19873_new_n2782_));
AND2X2 AND2X2_1168 ( .A(_abc_19873_new_n2783_), .B(_abc_19873_new_n2781_), .Y(_abc_19873_new_n2784_));
AND2X2 AND2X2_1169 ( .A(_abc_19873_new_n2784_), .B(reset_n), .Y(_0key2_reg_31_0__29_));
AND2X2 AND2X2_117 ( .A(_abc_19873_new_n928_), .B(core_key_38_), .Y(_abc_19873_new_n1066_));
AND2X2 AND2X2_1170 ( .A(_abc_19873_new_n2635_), .B(_abc_19873_new_n2302_), .Y(_abc_19873_new_n2787_));
AND2X2 AND2X2_1171 ( .A(_abc_19873_new_n2788_), .B(_abc_19873_new_n2786_), .Y(_abc_19873_new_n2789_));
AND2X2 AND2X2_1172 ( .A(_abc_19873_new_n2789_), .B(reset_n), .Y(_0key2_reg_31_0__30_));
AND2X2 AND2X2_1173 ( .A(_abc_19873_new_n2635_), .B(_abc_19873_new_n2308_), .Y(_abc_19873_new_n2792_));
AND2X2 AND2X2_1174 ( .A(_abc_19873_new_n2793_), .B(_abc_19873_new_n2791_), .Y(_abc_19873_new_n2794_));
AND2X2 AND2X2_1175 ( .A(_abc_19873_new_n2794_), .B(reset_n), .Y(_0key2_reg_31_0__31_));
AND2X2 AND2X2_1176 ( .A(_abc_19873_new_n928_), .B(_abc_19873_new_n2119_), .Y(_abc_19873_new_n2796_));
AND2X2 AND2X2_1177 ( .A(_abc_19873_new_n2796_), .B(_abc_19873_new_n2122_), .Y(_abc_19873_new_n2798_));
AND2X2 AND2X2_1178 ( .A(_abc_19873_new_n2799_), .B(reset_n), .Y(_abc_19873_new_n2800_));
AND2X2 AND2X2_1179 ( .A(_abc_19873_new_n2800_), .B(_abc_19873_new_n2797_), .Y(_0key1_reg_31_0__0_));
AND2X2 AND2X2_118 ( .A(_abc_19873_new_n916_), .B(core_key_70_), .Y(_abc_19873_new_n1067_));
AND2X2 AND2X2_1180 ( .A(_abc_19873_new_n2796_), .B(_abc_19873_new_n2128_), .Y(_abc_19873_new_n2803_));
AND2X2 AND2X2_1181 ( .A(_abc_19873_new_n2804_), .B(reset_n), .Y(_abc_19873_new_n2805_));
AND2X2 AND2X2_1182 ( .A(_abc_19873_new_n2805_), .B(_abc_19873_new_n2802_), .Y(_0key1_reg_31_0__1_));
AND2X2 AND2X2_1183 ( .A(_abc_19873_new_n2796_), .B(_abc_19873_new_n2134_), .Y(_abc_19873_new_n2808_));
AND2X2 AND2X2_1184 ( .A(_abc_19873_new_n2809_), .B(_abc_19873_new_n2807_), .Y(_abc_19873_new_n2810_));
AND2X2 AND2X2_1185 ( .A(_abc_19873_new_n2810_), .B(reset_n), .Y(_0key1_reg_31_0__2_));
AND2X2 AND2X2_1186 ( .A(_abc_19873_new_n2796_), .B(_abc_19873_new_n2140_), .Y(_abc_19873_new_n2813_));
AND2X2 AND2X2_1187 ( .A(_abc_19873_new_n2814_), .B(reset_n), .Y(_abc_19873_new_n2815_));
AND2X2 AND2X2_1188 ( .A(_abc_19873_new_n2815_), .B(_abc_19873_new_n2812_), .Y(_0key1_reg_31_0__3_));
AND2X2 AND2X2_1189 ( .A(_abc_19873_new_n2796_), .B(_abc_19873_new_n2146_), .Y(_abc_19873_new_n2818_));
AND2X2 AND2X2_119 ( .A(_abc_19873_new_n888_), .B(core_mi_6_), .Y(_abc_19873_new_n1070_));
AND2X2 AND2X2_1190 ( .A(_abc_19873_new_n2819_), .B(reset_n), .Y(_abc_19873_new_n2820_));
AND2X2 AND2X2_1191 ( .A(_abc_19873_new_n2820_), .B(_abc_19873_new_n2817_), .Y(_0key1_reg_31_0__4_));
AND2X2 AND2X2_1192 ( .A(_abc_19873_new_n2796_), .B(_abc_19873_new_n2152_), .Y(_abc_19873_new_n2823_));
AND2X2 AND2X2_1193 ( .A(_abc_19873_new_n2824_), .B(reset_n), .Y(_abc_19873_new_n2825_));
AND2X2 AND2X2_1194 ( .A(_abc_19873_new_n2825_), .B(_abc_19873_new_n2822_), .Y(_0key1_reg_31_0__5_));
AND2X2 AND2X2_1195 ( .A(_abc_19873_new_n2796_), .B(_abc_19873_new_n2158_), .Y(_abc_19873_new_n2828_));
AND2X2 AND2X2_1196 ( .A(_abc_19873_new_n2829_), .B(_abc_19873_new_n2827_), .Y(_abc_19873_new_n2830_));
AND2X2 AND2X2_1197 ( .A(_abc_19873_new_n2830_), .B(reset_n), .Y(_0key1_reg_31_0__6_));
AND2X2 AND2X2_1198 ( .A(_abc_19873_new_n2796_), .B(_abc_19873_new_n2164_), .Y(_abc_19873_new_n2833_));
AND2X2 AND2X2_1199 ( .A(_abc_19873_new_n2834_), .B(reset_n), .Y(_abc_19873_new_n2835_));
AND2X2 AND2X2_12 ( .A(_abc_19873_new_n875_), .B(_abc_19873_new_n887_), .Y(_abc_19873_new_n888_));
AND2X2 AND2X2_120 ( .A(_abc_19873_new_n881_), .B(core_key_102_), .Y(_abc_19873_new_n1071_));
AND2X2 AND2X2_1200 ( .A(_abc_19873_new_n2835_), .B(_abc_19873_new_n2832_), .Y(_0key1_reg_31_0__7_));
AND2X2 AND2X2_1201 ( .A(_abc_19873_new_n2796_), .B(_abc_19873_new_n2170_), .Y(_abc_19873_new_n2838_));
AND2X2 AND2X2_1202 ( .A(_abc_19873_new_n2839_), .B(_abc_19873_new_n2837_), .Y(_abc_19873_new_n2840_));
AND2X2 AND2X2_1203 ( .A(_abc_19873_new_n2840_), .B(reset_n), .Y(_0key1_reg_31_0__8_));
AND2X2 AND2X2_1204 ( .A(_abc_19873_new_n2796_), .B(_abc_19873_new_n2176_), .Y(_abc_19873_new_n2843_));
AND2X2 AND2X2_1205 ( .A(_abc_19873_new_n2844_), .B(_abc_19873_new_n2842_), .Y(_abc_19873_new_n2845_));
AND2X2 AND2X2_1206 ( .A(_abc_19873_new_n2845_), .B(reset_n), .Y(_0key1_reg_31_0__9_));
AND2X2 AND2X2_1207 ( .A(_abc_19873_new_n2796_), .B(_abc_19873_new_n2182_), .Y(_abc_19873_new_n2848_));
AND2X2 AND2X2_1208 ( .A(_abc_19873_new_n2849_), .B(_abc_19873_new_n2847_), .Y(_abc_19873_new_n2850_));
AND2X2 AND2X2_1209 ( .A(_abc_19873_new_n2850_), .B(reset_n), .Y(_0key1_reg_31_0__10_));
AND2X2 AND2X2_121 ( .A(_abc_19873_new_n907_), .B(word1_reg_6_), .Y(_abc_19873_new_n1073_));
AND2X2 AND2X2_1210 ( .A(_abc_19873_new_n2796_), .B(_abc_19873_new_n2188_), .Y(_abc_19873_new_n2853_));
AND2X2 AND2X2_1211 ( .A(_abc_19873_new_n2854_), .B(_abc_19873_new_n2852_), .Y(_abc_19873_new_n2855_));
AND2X2 AND2X2_1212 ( .A(_abc_19873_new_n2855_), .B(reset_n), .Y(_0key1_reg_31_0__11_));
AND2X2 AND2X2_1213 ( .A(_abc_19873_new_n2796_), .B(_abc_19873_new_n2194_), .Y(_abc_19873_new_n2858_));
AND2X2 AND2X2_1214 ( .A(_abc_19873_new_n2859_), .B(_abc_19873_new_n2857_), .Y(_abc_19873_new_n2860_));
AND2X2 AND2X2_1215 ( .A(_abc_19873_new_n2860_), .B(reset_n), .Y(_0key1_reg_31_0__12_));
AND2X2 AND2X2_1216 ( .A(_abc_19873_new_n2796_), .B(_abc_19873_new_n2200_), .Y(_abc_19873_new_n2863_));
AND2X2 AND2X2_1217 ( .A(_abc_19873_new_n2864_), .B(_abc_19873_new_n2862_), .Y(_abc_19873_new_n2865_));
AND2X2 AND2X2_1218 ( .A(_abc_19873_new_n2865_), .B(reset_n), .Y(_0key1_reg_31_0__13_));
AND2X2 AND2X2_1219 ( .A(_abc_19873_new_n2796_), .B(_abc_19873_new_n2206_), .Y(_abc_19873_new_n2868_));
AND2X2 AND2X2_122 ( .A(_abc_19873_new_n925_), .B(word2_reg_6_), .Y(_abc_19873_new_n1074_));
AND2X2 AND2X2_1220 ( .A(_abc_19873_new_n2869_), .B(_abc_19873_new_n2867_), .Y(_abc_19873_new_n2870_));
AND2X2 AND2X2_1221 ( .A(_abc_19873_new_n2870_), .B(reset_n), .Y(_0key1_reg_31_0__14_));
AND2X2 AND2X2_1222 ( .A(_abc_19873_new_n2796_), .B(_abc_19873_new_n2212_), .Y(_abc_19873_new_n2873_));
AND2X2 AND2X2_1223 ( .A(_abc_19873_new_n2874_), .B(_abc_19873_new_n2872_), .Y(_abc_19873_new_n2875_));
AND2X2 AND2X2_1224 ( .A(_abc_19873_new_n2875_), .B(reset_n), .Y(_0key1_reg_31_0__15_));
AND2X2 AND2X2_1225 ( .A(_abc_19873_new_n2796_), .B(_abc_19873_new_n2218_), .Y(_abc_19873_new_n2878_));
AND2X2 AND2X2_1226 ( .A(_abc_19873_new_n2879_), .B(_abc_19873_new_n2877_), .Y(_abc_19873_new_n2880_));
AND2X2 AND2X2_1227 ( .A(_abc_19873_new_n2880_), .B(reset_n), .Y(_0key1_reg_31_0__16_));
AND2X2 AND2X2_1228 ( .A(_abc_19873_new_n2796_), .B(_abc_19873_new_n2224_), .Y(_abc_19873_new_n2883_));
AND2X2 AND2X2_1229 ( .A(_abc_19873_new_n2884_), .B(_abc_19873_new_n2882_), .Y(_abc_19873_new_n2885_));
AND2X2 AND2X2_123 ( .A(_abc_19873_new_n930_), .B(word0_reg_6_), .Y(_abc_19873_new_n1077_));
AND2X2 AND2X2_1230 ( .A(_abc_19873_new_n2885_), .B(reset_n), .Y(_0key1_reg_31_0__17_));
AND2X2 AND2X2_1231 ( .A(_abc_19873_new_n2796_), .B(_abc_19873_new_n2230_), .Y(_abc_19873_new_n2888_));
AND2X2 AND2X2_1232 ( .A(_abc_19873_new_n2889_), .B(_abc_19873_new_n2887_), .Y(_abc_19873_new_n2890_));
AND2X2 AND2X2_1233 ( .A(_abc_19873_new_n2890_), .B(reset_n), .Y(_0key1_reg_31_0__18_));
AND2X2 AND2X2_1234 ( .A(_abc_19873_new_n2796_), .B(_abc_19873_new_n2236_), .Y(_abc_19873_new_n2893_));
AND2X2 AND2X2_1235 ( .A(_abc_19873_new_n2894_), .B(_abc_19873_new_n2892_), .Y(_abc_19873_new_n2895_));
AND2X2 AND2X2_1236 ( .A(_abc_19873_new_n2895_), .B(reset_n), .Y(_0key1_reg_31_0__19_));
AND2X2 AND2X2_1237 ( .A(_abc_19873_new_n2796_), .B(_abc_19873_new_n2242_), .Y(_abc_19873_new_n2898_));
AND2X2 AND2X2_1238 ( .A(_abc_19873_new_n2899_), .B(_abc_19873_new_n2897_), .Y(_abc_19873_new_n2900_));
AND2X2 AND2X2_1239 ( .A(_abc_19873_new_n2900_), .B(reset_n), .Y(_0key1_reg_31_0__20_));
AND2X2 AND2X2_124 ( .A(_abc_19873_new_n901_), .B(core_key_6_), .Y(_abc_19873_new_n1079_));
AND2X2 AND2X2_1240 ( .A(_abc_19873_new_n2796_), .B(_abc_19873_new_n2248_), .Y(_abc_19873_new_n2903_));
AND2X2 AND2X2_1241 ( .A(_abc_19873_new_n2904_), .B(_abc_19873_new_n2902_), .Y(_abc_19873_new_n2905_));
AND2X2 AND2X2_1242 ( .A(_abc_19873_new_n2905_), .B(reset_n), .Y(_0key1_reg_31_0__21_));
AND2X2 AND2X2_1243 ( .A(_abc_19873_new_n2796_), .B(_abc_19873_new_n2254_), .Y(_abc_19873_new_n2908_));
AND2X2 AND2X2_1244 ( .A(_abc_19873_new_n2909_), .B(_abc_19873_new_n2907_), .Y(_abc_19873_new_n2910_));
AND2X2 AND2X2_1245 ( .A(_abc_19873_new_n2910_), .B(reset_n), .Y(_0key1_reg_31_0__22_));
AND2X2 AND2X2_1246 ( .A(_abc_19873_new_n2796_), .B(_abc_19873_new_n2260_), .Y(_abc_19873_new_n2913_));
AND2X2 AND2X2_1247 ( .A(_abc_19873_new_n2914_), .B(_abc_19873_new_n2912_), .Y(_abc_19873_new_n2915_));
AND2X2 AND2X2_1248 ( .A(_abc_19873_new_n2915_), .B(reset_n), .Y(_0key1_reg_31_0__23_));
AND2X2 AND2X2_1249 ( .A(_abc_19873_new_n2796_), .B(_abc_19873_new_n2266_), .Y(_abc_19873_new_n2918_));
AND2X2 AND2X2_125 ( .A(_abc_19873_new_n912_), .B(word3_reg_6_), .Y(_abc_19873_new_n1080_));
AND2X2 AND2X2_1250 ( .A(_abc_19873_new_n2919_), .B(_abc_19873_new_n2917_), .Y(_abc_19873_new_n2920_));
AND2X2 AND2X2_1251 ( .A(_abc_19873_new_n2920_), .B(reset_n), .Y(_0key1_reg_31_0__24_));
AND2X2 AND2X2_1252 ( .A(_abc_19873_new_n2796_), .B(_abc_19873_new_n2272_), .Y(_abc_19873_new_n2923_));
AND2X2 AND2X2_1253 ( .A(_abc_19873_new_n2924_), .B(_abc_19873_new_n2922_), .Y(_abc_19873_new_n2925_));
AND2X2 AND2X2_1254 ( .A(_abc_19873_new_n2925_), .B(reset_n), .Y(_0key1_reg_31_0__25_));
AND2X2 AND2X2_1255 ( .A(_abc_19873_new_n2796_), .B(_abc_19873_new_n2278_), .Y(_abc_19873_new_n2928_));
AND2X2 AND2X2_1256 ( .A(_abc_19873_new_n2929_), .B(_abc_19873_new_n2927_), .Y(_abc_19873_new_n2930_));
AND2X2 AND2X2_1257 ( .A(_abc_19873_new_n2930_), .B(reset_n), .Y(_0key1_reg_31_0__26_));
AND2X2 AND2X2_1258 ( .A(_abc_19873_new_n2796_), .B(_abc_19873_new_n2284_), .Y(_abc_19873_new_n2933_));
AND2X2 AND2X2_1259 ( .A(_abc_19873_new_n2934_), .B(_abc_19873_new_n2932_), .Y(_abc_19873_new_n2935_));
AND2X2 AND2X2_126 ( .A(_abc_19873_new_n1084_), .B(_abc_19873_new_n937_), .Y(\read_data[6] ));
AND2X2 AND2X2_1260 ( .A(_abc_19873_new_n2935_), .B(reset_n), .Y(_0key1_reg_31_0__27_));
AND2X2 AND2X2_1261 ( .A(_abc_19873_new_n2796_), .B(_abc_19873_new_n2290_), .Y(_abc_19873_new_n2938_));
AND2X2 AND2X2_1262 ( .A(_abc_19873_new_n2939_), .B(_abc_19873_new_n2937_), .Y(_abc_19873_new_n2940_));
AND2X2 AND2X2_1263 ( .A(_abc_19873_new_n2940_), .B(reset_n), .Y(_0key1_reg_31_0__28_));
AND2X2 AND2X2_1264 ( .A(_abc_19873_new_n2796_), .B(_abc_19873_new_n2296_), .Y(_abc_19873_new_n2943_));
AND2X2 AND2X2_1265 ( .A(_abc_19873_new_n2944_), .B(_abc_19873_new_n2942_), .Y(_abc_19873_new_n2945_));
AND2X2 AND2X2_1266 ( .A(_abc_19873_new_n2945_), .B(reset_n), .Y(_0key1_reg_31_0__29_));
AND2X2 AND2X2_1267 ( .A(_abc_19873_new_n2796_), .B(_abc_19873_new_n2302_), .Y(_abc_19873_new_n2948_));
AND2X2 AND2X2_1268 ( .A(_abc_19873_new_n2949_), .B(_abc_19873_new_n2947_), .Y(_abc_19873_new_n2950_));
AND2X2 AND2X2_1269 ( .A(_abc_19873_new_n2950_), .B(reset_n), .Y(_0key1_reg_31_0__30_));
AND2X2 AND2X2_127 ( .A(_abc_19873_new_n901_), .B(core_key_7_), .Y(_abc_19873_new_n1086_));
AND2X2 AND2X2_1270 ( .A(_abc_19873_new_n2796_), .B(_abc_19873_new_n2308_), .Y(_abc_19873_new_n2953_));
AND2X2 AND2X2_1271 ( .A(_abc_19873_new_n2954_), .B(_abc_19873_new_n2952_), .Y(_abc_19873_new_n2955_));
AND2X2 AND2X2_1272 ( .A(_abc_19873_new_n2955_), .B(reset_n), .Y(_0key1_reg_31_0__31_));
AND2X2 AND2X2_1273 ( .A(_abc_19873_new_n901_), .B(_abc_19873_new_n2119_), .Y(_abc_19873_new_n2957_));
AND2X2 AND2X2_1274 ( .A(_abc_19873_new_n2957_), .B(_abc_19873_new_n2122_), .Y(_abc_19873_new_n2959_));
AND2X2 AND2X2_1275 ( .A(_abc_19873_new_n2960_), .B(reset_n), .Y(_abc_19873_new_n2961_));
AND2X2 AND2X2_1276 ( .A(_abc_19873_new_n2961_), .B(_abc_19873_new_n2958_), .Y(_0key0_reg_31_0__0_));
AND2X2 AND2X2_1277 ( .A(_abc_19873_new_n2957_), .B(_abc_19873_new_n2128_), .Y(_abc_19873_new_n2964_));
AND2X2 AND2X2_1278 ( .A(_abc_19873_new_n2965_), .B(reset_n), .Y(_abc_19873_new_n2966_));
AND2X2 AND2X2_1279 ( .A(_abc_19873_new_n2966_), .B(_abc_19873_new_n2963_), .Y(_0key0_reg_31_0__1_));
AND2X2 AND2X2_128 ( .A(_abc_19873_new_n928_), .B(core_key_39_), .Y(_abc_19873_new_n1087_));
AND2X2 AND2X2_1280 ( .A(_abc_19873_new_n2957_), .B(_abc_19873_new_n2134_), .Y(_abc_19873_new_n2969_));
AND2X2 AND2X2_1281 ( .A(_abc_19873_new_n2970_), .B(reset_n), .Y(_abc_19873_new_n2971_));
AND2X2 AND2X2_1282 ( .A(_abc_19873_new_n2971_), .B(_abc_19873_new_n2968_), .Y(_0key0_reg_31_0__2_));
AND2X2 AND2X2_1283 ( .A(_abc_19873_new_n2957_), .B(_abc_19873_new_n2140_), .Y(_abc_19873_new_n2974_));
AND2X2 AND2X2_1284 ( .A(_abc_19873_new_n2975_), .B(reset_n), .Y(_abc_19873_new_n2976_));
AND2X2 AND2X2_1285 ( .A(_abc_19873_new_n2976_), .B(_abc_19873_new_n2973_), .Y(_0key0_reg_31_0__3_));
AND2X2 AND2X2_1286 ( .A(_abc_19873_new_n2957_), .B(_abc_19873_new_n2146_), .Y(_abc_19873_new_n2979_));
AND2X2 AND2X2_1287 ( .A(_abc_19873_new_n2980_), .B(reset_n), .Y(_abc_19873_new_n2981_));
AND2X2 AND2X2_1288 ( .A(_abc_19873_new_n2981_), .B(_abc_19873_new_n2978_), .Y(_0key0_reg_31_0__4_));
AND2X2 AND2X2_1289 ( .A(_abc_19873_new_n2957_), .B(_abc_19873_new_n2152_), .Y(_abc_19873_new_n2984_));
AND2X2 AND2X2_129 ( .A(_abc_19873_new_n919_), .B(core_mi_39_), .Y(_abc_19873_new_n1089_));
AND2X2 AND2X2_1290 ( .A(_abc_19873_new_n2985_), .B(reset_n), .Y(_abc_19873_new_n2986_));
AND2X2 AND2X2_1291 ( .A(_abc_19873_new_n2986_), .B(_abc_19873_new_n2983_), .Y(_0key0_reg_31_0__5_));
AND2X2 AND2X2_1292 ( .A(_abc_19873_new_n2957_), .B(_abc_19873_new_n2158_), .Y(_abc_19873_new_n2989_));
AND2X2 AND2X2_1293 ( .A(_abc_19873_new_n2990_), .B(reset_n), .Y(_abc_19873_new_n2991_));
AND2X2 AND2X2_1294 ( .A(_abc_19873_new_n2991_), .B(_abc_19873_new_n2988_), .Y(_0key0_reg_31_0__6_));
AND2X2 AND2X2_1295 ( .A(_abc_19873_new_n2957_), .B(_abc_19873_new_n2164_), .Y(_abc_19873_new_n2994_));
AND2X2 AND2X2_1296 ( .A(_abc_19873_new_n2995_), .B(reset_n), .Y(_abc_19873_new_n2996_));
AND2X2 AND2X2_1297 ( .A(_abc_19873_new_n2996_), .B(_abc_19873_new_n2993_), .Y(_0key0_reg_31_0__7_));
AND2X2 AND2X2_1298 ( .A(_abc_19873_new_n2957_), .B(_abc_19873_new_n2170_), .Y(_abc_19873_new_n2999_));
AND2X2 AND2X2_1299 ( .A(_abc_19873_new_n3000_), .B(reset_n), .Y(_abc_19873_new_n3001_));
AND2X2 AND2X2_13 ( .A(_abc_19873_new_n888_), .B(core_mi_0_), .Y(_abc_19873_new_n889_));
AND2X2 AND2X2_130 ( .A(_abc_19873_new_n930_), .B(word0_reg_7_), .Y(_abc_19873_new_n1090_));
AND2X2 AND2X2_1300 ( .A(_abc_19873_new_n3001_), .B(_abc_19873_new_n2998_), .Y(_0key0_reg_31_0__8_));
AND2X2 AND2X2_1301 ( .A(_abc_19873_new_n2957_), .B(_abc_19873_new_n2176_), .Y(_abc_19873_new_n3004_));
AND2X2 AND2X2_1302 ( .A(_abc_19873_new_n3005_), .B(reset_n), .Y(_abc_19873_new_n3006_));
AND2X2 AND2X2_1303 ( .A(_abc_19873_new_n3006_), .B(_abc_19873_new_n3003_), .Y(_0key0_reg_31_0__9_));
AND2X2 AND2X2_1304 ( .A(_abc_19873_new_n2957_), .B(_abc_19873_new_n2182_), .Y(_abc_19873_new_n3009_));
AND2X2 AND2X2_1305 ( .A(_abc_19873_new_n3010_), .B(reset_n), .Y(_abc_19873_new_n3011_));
AND2X2 AND2X2_1306 ( .A(_abc_19873_new_n3011_), .B(_abc_19873_new_n3008_), .Y(_0key0_reg_31_0__10_));
AND2X2 AND2X2_1307 ( .A(_abc_19873_new_n2957_), .B(_abc_19873_new_n2188_), .Y(_abc_19873_new_n3014_));
AND2X2 AND2X2_1308 ( .A(_abc_19873_new_n3015_), .B(reset_n), .Y(_abc_19873_new_n3016_));
AND2X2 AND2X2_1309 ( .A(_abc_19873_new_n3016_), .B(_abc_19873_new_n3013_), .Y(_0key0_reg_31_0__11_));
AND2X2 AND2X2_131 ( .A(_abc_19873_new_n925_), .B(word2_reg_7_), .Y(_abc_19873_new_n1093_));
AND2X2 AND2X2_1310 ( .A(_abc_19873_new_n2957_), .B(_abc_19873_new_n2194_), .Y(_abc_19873_new_n3019_));
AND2X2 AND2X2_1311 ( .A(_abc_19873_new_n3020_), .B(reset_n), .Y(_abc_19873_new_n3021_));
AND2X2 AND2X2_1312 ( .A(_abc_19873_new_n3021_), .B(_abc_19873_new_n3018_), .Y(_0key0_reg_31_0__12_));
AND2X2 AND2X2_1313 ( .A(_abc_19873_new_n2957_), .B(_abc_19873_new_n2200_), .Y(_abc_19873_new_n3024_));
AND2X2 AND2X2_1314 ( .A(_abc_19873_new_n3025_), .B(reset_n), .Y(_abc_19873_new_n3026_));
AND2X2 AND2X2_1315 ( .A(_abc_19873_new_n3026_), .B(_abc_19873_new_n3023_), .Y(_0key0_reg_31_0__13_));
AND2X2 AND2X2_1316 ( .A(_abc_19873_new_n2957_), .B(_abc_19873_new_n2206_), .Y(_abc_19873_new_n3029_));
AND2X2 AND2X2_1317 ( .A(_abc_19873_new_n3030_), .B(reset_n), .Y(_abc_19873_new_n3031_));
AND2X2 AND2X2_1318 ( .A(_abc_19873_new_n3031_), .B(_abc_19873_new_n3028_), .Y(_0key0_reg_31_0__14_));
AND2X2 AND2X2_1319 ( .A(_abc_19873_new_n2957_), .B(_abc_19873_new_n2212_), .Y(_abc_19873_new_n3034_));
AND2X2 AND2X2_132 ( .A(_abc_19873_new_n907_), .B(word1_reg_7_), .Y(_abc_19873_new_n1094_));
AND2X2 AND2X2_1320 ( .A(_abc_19873_new_n3035_), .B(reset_n), .Y(_abc_19873_new_n3036_));
AND2X2 AND2X2_1321 ( .A(_abc_19873_new_n3036_), .B(_abc_19873_new_n3033_), .Y(_0key0_reg_31_0__15_));
AND2X2 AND2X2_1322 ( .A(_abc_19873_new_n2957_), .B(_abc_19873_new_n2218_), .Y(_abc_19873_new_n3039_));
AND2X2 AND2X2_1323 ( .A(_abc_19873_new_n3040_), .B(reset_n), .Y(_abc_19873_new_n3041_));
AND2X2 AND2X2_1324 ( .A(_abc_19873_new_n3041_), .B(_abc_19873_new_n3038_), .Y(_0key0_reg_31_0__16_));
AND2X2 AND2X2_1325 ( .A(_abc_19873_new_n2957_), .B(_abc_19873_new_n2224_), .Y(_abc_19873_new_n3044_));
AND2X2 AND2X2_1326 ( .A(_abc_19873_new_n3045_), .B(reset_n), .Y(_abc_19873_new_n3046_));
AND2X2 AND2X2_1327 ( .A(_abc_19873_new_n3046_), .B(_abc_19873_new_n3043_), .Y(_0key0_reg_31_0__17_));
AND2X2 AND2X2_1328 ( .A(_abc_19873_new_n2957_), .B(_abc_19873_new_n2230_), .Y(_abc_19873_new_n3049_));
AND2X2 AND2X2_1329 ( .A(_abc_19873_new_n3050_), .B(reset_n), .Y(_abc_19873_new_n3051_));
AND2X2 AND2X2_133 ( .A(_abc_19873_new_n912_), .B(word3_reg_7_), .Y(_abc_19873_new_n1095_));
AND2X2 AND2X2_1330 ( .A(_abc_19873_new_n3051_), .B(_abc_19873_new_n3048_), .Y(_0key0_reg_31_0__18_));
AND2X2 AND2X2_1331 ( .A(_abc_19873_new_n2957_), .B(_abc_19873_new_n2236_), .Y(_abc_19873_new_n3054_));
AND2X2 AND2X2_1332 ( .A(_abc_19873_new_n3055_), .B(reset_n), .Y(_abc_19873_new_n3056_));
AND2X2 AND2X2_1333 ( .A(_abc_19873_new_n3056_), .B(_abc_19873_new_n3053_), .Y(_0key0_reg_31_0__19_));
AND2X2 AND2X2_1334 ( .A(_abc_19873_new_n2957_), .B(_abc_19873_new_n2242_), .Y(_abc_19873_new_n3059_));
AND2X2 AND2X2_1335 ( .A(_abc_19873_new_n3060_), .B(reset_n), .Y(_abc_19873_new_n3061_));
AND2X2 AND2X2_1336 ( .A(_abc_19873_new_n3061_), .B(_abc_19873_new_n3058_), .Y(_0key0_reg_31_0__20_));
AND2X2 AND2X2_1337 ( .A(_abc_19873_new_n2957_), .B(_abc_19873_new_n2248_), .Y(_abc_19873_new_n3064_));
AND2X2 AND2X2_1338 ( .A(_abc_19873_new_n3065_), .B(reset_n), .Y(_abc_19873_new_n3066_));
AND2X2 AND2X2_1339 ( .A(_abc_19873_new_n3066_), .B(_abc_19873_new_n3063_), .Y(_0key0_reg_31_0__21_));
AND2X2 AND2X2_134 ( .A(_abc_19873_new_n897_), .B(core_final_rounds_3_), .Y(_abc_19873_new_n1098_));
AND2X2 AND2X2_1340 ( .A(_abc_19873_new_n2957_), .B(_abc_19873_new_n2254_), .Y(_abc_19873_new_n3069_));
AND2X2 AND2X2_1341 ( .A(_abc_19873_new_n3070_), .B(reset_n), .Y(_abc_19873_new_n3071_));
AND2X2 AND2X2_1342 ( .A(_abc_19873_new_n3071_), .B(_abc_19873_new_n3068_), .Y(_0key0_reg_31_0__22_));
AND2X2 AND2X2_1343 ( .A(_abc_19873_new_n2957_), .B(_abc_19873_new_n2260_), .Y(_abc_19873_new_n3074_));
AND2X2 AND2X2_1344 ( .A(_abc_19873_new_n3075_), .B(reset_n), .Y(_abc_19873_new_n3076_));
AND2X2 AND2X2_1345 ( .A(_abc_19873_new_n3076_), .B(_abc_19873_new_n3073_), .Y(_0key0_reg_31_0__23_));
AND2X2 AND2X2_1346 ( .A(_abc_19873_new_n2957_), .B(_abc_19873_new_n2266_), .Y(_abc_19873_new_n3079_));
AND2X2 AND2X2_1347 ( .A(_abc_19873_new_n3080_), .B(reset_n), .Y(_abc_19873_new_n3081_));
AND2X2 AND2X2_1348 ( .A(_abc_19873_new_n3081_), .B(_abc_19873_new_n3078_), .Y(_0key0_reg_31_0__24_));
AND2X2 AND2X2_1349 ( .A(_abc_19873_new_n2957_), .B(_abc_19873_new_n2272_), .Y(_abc_19873_new_n3084_));
AND2X2 AND2X2_135 ( .A(_abc_19873_new_n916_), .B(core_key_71_), .Y(_abc_19873_new_n1099_));
AND2X2 AND2X2_1350 ( .A(_abc_19873_new_n3085_), .B(reset_n), .Y(_abc_19873_new_n3086_));
AND2X2 AND2X2_1351 ( .A(_abc_19873_new_n3086_), .B(_abc_19873_new_n3083_), .Y(_0key0_reg_31_0__25_));
AND2X2 AND2X2_1352 ( .A(_abc_19873_new_n2957_), .B(_abc_19873_new_n2278_), .Y(_abc_19873_new_n3089_));
AND2X2 AND2X2_1353 ( .A(_abc_19873_new_n3090_), .B(reset_n), .Y(_abc_19873_new_n3091_));
AND2X2 AND2X2_1354 ( .A(_abc_19873_new_n3091_), .B(_abc_19873_new_n3088_), .Y(_0key0_reg_31_0__26_));
AND2X2 AND2X2_1355 ( .A(_abc_19873_new_n2957_), .B(_abc_19873_new_n2284_), .Y(_abc_19873_new_n3094_));
AND2X2 AND2X2_1356 ( .A(_abc_19873_new_n3095_), .B(reset_n), .Y(_abc_19873_new_n3096_));
AND2X2 AND2X2_1357 ( .A(_abc_19873_new_n3096_), .B(_abc_19873_new_n3093_), .Y(_0key0_reg_31_0__27_));
AND2X2 AND2X2_1358 ( .A(_abc_19873_new_n2957_), .B(_abc_19873_new_n2290_), .Y(_abc_19873_new_n3099_));
AND2X2 AND2X2_1359 ( .A(_abc_19873_new_n3100_), .B(reset_n), .Y(_abc_19873_new_n3101_));
AND2X2 AND2X2_136 ( .A(_abc_19873_new_n881_), .B(core_key_103_), .Y(_abc_19873_new_n1101_));
AND2X2 AND2X2_1360 ( .A(_abc_19873_new_n3101_), .B(_abc_19873_new_n3098_), .Y(_0key0_reg_31_0__28_));
AND2X2 AND2X2_1361 ( .A(_abc_19873_new_n2957_), .B(_abc_19873_new_n2296_), .Y(_abc_19873_new_n3104_));
AND2X2 AND2X2_1362 ( .A(_abc_19873_new_n3105_), .B(reset_n), .Y(_abc_19873_new_n3106_));
AND2X2 AND2X2_1363 ( .A(_abc_19873_new_n3106_), .B(_abc_19873_new_n3103_), .Y(_0key0_reg_31_0__29_));
AND2X2 AND2X2_1364 ( .A(_abc_19873_new_n2957_), .B(_abc_19873_new_n2302_), .Y(_abc_19873_new_n3109_));
AND2X2 AND2X2_1365 ( .A(_abc_19873_new_n3110_), .B(reset_n), .Y(_abc_19873_new_n3111_));
AND2X2 AND2X2_1366 ( .A(_abc_19873_new_n3111_), .B(_abc_19873_new_n3108_), .Y(_0key0_reg_31_0__30_));
AND2X2 AND2X2_1367 ( .A(_abc_19873_new_n2957_), .B(_abc_19873_new_n2308_), .Y(_abc_19873_new_n3114_));
AND2X2 AND2X2_1368 ( .A(_abc_19873_new_n3115_), .B(reset_n), .Y(_abc_19873_new_n3116_));
AND2X2 AND2X2_1369 ( .A(_abc_19873_new_n3116_), .B(_abc_19873_new_n3113_), .Y(_0key0_reg_31_0__31_));
AND2X2 AND2X2_137 ( .A(_abc_19873_new_n888_), .B(core_mi_7_), .Y(_abc_19873_new_n1102_));
AND2X2 AND2X2_1370 ( .A(_abc_19873_new_n897_), .B(_abc_19873_new_n2119_), .Y(_abc_19873_new_n3118_));
AND2X2 AND2X2_1371 ( .A(_abc_19873_new_n3118_), .B(\write_data[0] ), .Y(_abc_19873_new_n3119_));
AND2X2 AND2X2_1372 ( .A(_abc_19873_new_n3120_), .B(core_compression_rounds_0_), .Y(_abc_19873_new_n3121_));
AND2X2 AND2X2_1373 ( .A(_abc_19873_new_n3122_), .B(reset_n), .Y(_0param_reg_7_0__0_));
AND2X2 AND2X2_1374 ( .A(_abc_19873_new_n3120_), .B(core_compression_rounds_1_), .Y(_abc_19873_new_n3124_));
AND2X2 AND2X2_1375 ( .A(_abc_19873_new_n3118_), .B(\write_data[1] ), .Y(_abc_19873_new_n3126_));
AND2X2 AND2X2_1376 ( .A(_abc_19873_new_n3120_), .B(core_compression_rounds_2_), .Y(_abc_19873_new_n3129_));
AND2X2 AND2X2_1377 ( .A(_abc_19873_new_n3118_), .B(\write_data[2] ), .Y(_abc_19873_new_n3130_));
AND2X2 AND2X2_1378 ( .A(_abc_19873_new_n3131_), .B(reset_n), .Y(_0param_reg_7_0__2_));
AND2X2 AND2X2_1379 ( .A(_abc_19873_new_n3118_), .B(\write_data[3] ), .Y(_abc_19873_new_n3133_));
AND2X2 AND2X2_138 ( .A(_abc_19873_new_n1106_), .B(_abc_19873_new_n937_), .Y(\read_data[7] ));
AND2X2 AND2X2_1380 ( .A(_abc_19873_new_n3120_), .B(core_compression_rounds_3_), .Y(_abc_19873_new_n3134_));
AND2X2 AND2X2_1381 ( .A(_abc_19873_new_n3135_), .B(reset_n), .Y(_0param_reg_7_0__3_));
AND2X2 AND2X2_1382 ( .A(_abc_19873_new_n3118_), .B(\write_data[4] ), .Y(_abc_19873_new_n3137_));
AND2X2 AND2X2_1383 ( .A(_abc_19873_new_n3120_), .B(core_final_rounds_0_), .Y(_abc_19873_new_n3138_));
AND2X2 AND2X2_1384 ( .A(_abc_19873_new_n3139_), .B(reset_n), .Y(_0param_reg_7_0__4_));
AND2X2 AND2X2_1385 ( .A(_abc_19873_new_n3118_), .B(\write_data[5] ), .Y(_abc_19873_new_n3141_));
AND2X2 AND2X2_1386 ( .A(_abc_19873_new_n3120_), .B(core_final_rounds_1_), .Y(_abc_19873_new_n3142_));
AND2X2 AND2X2_1387 ( .A(_abc_19873_new_n3143_), .B(reset_n), .Y(_0param_reg_7_0__5_));
AND2X2 AND2X2_1388 ( .A(_abc_19873_new_n3120_), .B(core_final_rounds_2_), .Y(_abc_19873_new_n3145_));
AND2X2 AND2X2_1389 ( .A(_abc_19873_new_n3118_), .B(\write_data[6] ), .Y(_abc_19873_new_n3146_));
AND2X2 AND2X2_139 ( .A(_abc_19873_new_n881_), .B(core_key_104_), .Y(_abc_19873_new_n1108_));
AND2X2 AND2X2_1390 ( .A(_abc_19873_new_n3118_), .B(\write_data[7] ), .Y(_abc_19873_new_n3149_));
AND2X2 AND2X2_1391 ( .A(_abc_19873_new_n3120_), .B(core_final_rounds_3_), .Y(_abc_19873_new_n3150_));
AND2X2 AND2X2_1392 ( .A(_abc_19873_new_n3151_), .B(reset_n), .Y(_0param_reg_7_0__7_));
AND2X2 AND2X2_1393 ( .A(_abc_19873_new_n2119_), .B(reset_n), .Y(_abc_19873_new_n3153_));
AND2X2 AND2X2_1394 ( .A(_abc_19873_new_n3153_), .B(\write_data[0] ), .Y(_abc_19873_new_n3154_));
AND2X2 AND2X2_1395 ( .A(_abc_19873_new_n894_), .B(_abc_19873_new_n3154_), .Y(_0ctrl_reg_2_0__0_));
AND2X2 AND2X2_1396 ( .A(_abc_19873_new_n3153_), .B(\write_data[1] ), .Y(_abc_19873_new_n3156_));
AND2X2 AND2X2_1397 ( .A(_abc_19873_new_n894_), .B(_abc_19873_new_n3156_), .Y(_0ctrl_reg_2_0__1_));
AND2X2 AND2X2_1398 ( .A(_abc_19873_new_n3153_), .B(\write_data[2] ), .Y(_abc_19873_new_n3158_));
AND2X2 AND2X2_1399 ( .A(_abc_19873_new_n894_), .B(_abc_19873_new_n3158_), .Y(_0ctrl_reg_2_0__2_));
AND2X2 AND2X2_14 ( .A(_abc_19873_new_n891_), .B(_abc_19873_new_n873_), .Y(_abc_19873_new_n892_));
AND2X2 AND2X2_140 ( .A(_abc_19873_new_n916_), .B(core_key_72_), .Y(_abc_19873_new_n1109_));
AND2X2 AND2X2_1400 ( .A(_abc_19873_new_n886_), .B(_abc_19873_new_n914_), .Y(_abc_19873_new_n3160_));
AND2X2 AND2X2_1401 ( .A(_abc_19873_new_n3160_), .B(_abc_19873_new_n2119_), .Y(_abc_19873_new_n3161_));
AND2X2 AND2X2_1402 ( .A(_abc_19873_new_n3161_), .B(_abc_19873_new_n893_), .Y(_abc_19873_new_n3162_));
AND2X2 AND2X2_1403 ( .A(_abc_19873_new_n3162_), .B(_abc_19873_new_n2122_), .Y(_abc_19873_new_n3163_));
AND2X2 AND2X2_1404 ( .A(_abc_19873_new_n3165_), .B(reset_n), .Y(_abc_19873_new_n3166_));
AND2X2 AND2X2_1405 ( .A(_abc_19873_new_n3166_), .B(_abc_19873_new_n3164_), .Y(_0long_reg_0_0_));
AND2X2 AND2X2_1406 ( .A(core__abc_22172_new_n1132_), .B(core__abc_22172_new_n1133_), .Y(core__abc_22172_new_n1134_));
AND2X2 AND2X2_1407 ( .A(core__abc_22172_new_n1134_), .B(core__abc_22172_new_n1131_), .Y(core__abc_22172_new_n1135_));
AND2X2 AND2X2_1408 ( .A(core__abc_22172_new_n1135_), .B(core__abc_22172_new_n1130_), .Y(core__abc_22172_new_n1136_));
AND2X2 AND2X2_1409 ( .A(core__abc_22172_new_n1137_), .B(core_final_rounds_3_), .Y(core__abc_22172_new_n1138_));
AND2X2 AND2X2_141 ( .A(_abc_19873_new_n925_), .B(word2_reg_8_), .Y(_abc_19873_new_n1111_));
AND2X2 AND2X2_1410 ( .A(core__abc_22172_new_n1140_), .B(core_loop_ctr_reg_3_), .Y(core__abc_22172_new_n1141_));
AND2X2 AND2X2_1411 ( .A(core__abc_22172_new_n1139_), .B(core__abc_22172_new_n1142_), .Y(core__abc_22172_new_n1143_));
AND2X2 AND2X2_1412 ( .A(core__abc_22172_new_n1137_), .B(core__abc_22172_new_n1146_), .Y(core__abc_22172_new_n1147_));
AND2X2 AND2X2_1413 ( .A(core__abc_22172_new_n1147_), .B(core_loop_ctr_reg_2_), .Y(core__abc_22172_new_n1148_));
AND2X2 AND2X2_1414 ( .A(core__abc_22172_new_n1149_), .B(core__abc_22172_new_n1150_), .Y(core__abc_22172_new_n1151_));
AND2X2 AND2X2_1415 ( .A(core_final_rounds_0_), .B(core_loop_ctr_reg_0_), .Y(core__abc_22172_new_n1152_));
AND2X2 AND2X2_1416 ( .A(core__abc_22172_new_n1132_), .B(core__abc_22172_new_n1155_), .Y(core__abc_22172_new_n1156_));
AND2X2 AND2X2_1417 ( .A(core_final_rounds_1_), .B(core_loop_ctr_reg_1_), .Y(core__abc_22172_new_n1157_));
AND2X2 AND2X2_1418 ( .A(core__abc_22172_new_n1158_), .B(core__abc_22172_new_n1133_), .Y(core__abc_22172_new_n1159_));
AND2X2 AND2X2_1419 ( .A(core__abc_22172_new_n1160_), .B(core__abc_22172_new_n1161_), .Y(core__abc_22172_new_n1162_));
AND2X2 AND2X2_142 ( .A(_abc_19873_new_n907_), .B(word1_reg_8_), .Y(_abc_19873_new_n1112_));
AND2X2 AND2X2_1420 ( .A(core__abc_22172_new_n1162_), .B(core__abc_22172_new_n1154_), .Y(core__abc_22172_new_n1163_));
AND2X2 AND2X2_1421 ( .A(core__abc_22172_new_n1151_), .B(core__abc_22172_new_n1163_), .Y(core__abc_22172_new_n1164_));
AND2X2 AND2X2_1422 ( .A(core__abc_22172_new_n1145_), .B(core__abc_22172_new_n1164_), .Y(core__abc_22172_new_n1165_));
AND2X2 AND2X2_1423 ( .A(core__abc_22172_new_n1165_), .B(core__abc_22172_new_n1166_), .Y(core__abc_22172_new_n1167_));
AND2X2 AND2X2_1424 ( .A(core__abc_22172_new_n1171_), .B(core__abc_22172_new_n1169_), .Y(core__abc_22172_new_n1172_));
AND2X2 AND2X2_1425 ( .A(core__abc_22172_new_n1172_), .B(core__abc_22172_new_n1168_), .Y(core__abc_22172_new_n1173_));
AND2X2 AND2X2_1426 ( .A(core__abc_22172_new_n1178_), .B(core__abc_22172_new_n1179_), .Y(core__abc_22172_new_n1180_));
AND2X2 AND2X2_1427 ( .A(core__abc_22172_new_n1180_), .B(core__abc_22172_new_n1177_), .Y(core__abc_22172_new_n1181_));
AND2X2 AND2X2_1428 ( .A(core__abc_22172_new_n1181_), .B(core__abc_22172_new_n1176_), .Y(core__abc_22172_new_n1182_));
AND2X2 AND2X2_1429 ( .A(core__abc_22172_new_n1183_), .B(core_compression_rounds_3_), .Y(core__abc_22172_new_n1184_));
AND2X2 AND2X2_143 ( .A(_abc_19873_new_n930_), .B(word0_reg_8_), .Y(_abc_19873_new_n1113_));
AND2X2 AND2X2_1430 ( .A(core__abc_22172_new_n1186_), .B(core_loop_ctr_reg_3_), .Y(core__abc_22172_new_n1187_));
AND2X2 AND2X2_1431 ( .A(core_loop_ctr_reg_0_), .B(core_compression_rounds_0_), .Y(core__abc_22172_new_n1189_));
AND2X2 AND2X2_1432 ( .A(core__abc_22172_new_n1155_), .B(core__abc_22172_new_n1178_), .Y(core__abc_22172_new_n1192_));
AND2X2 AND2X2_1433 ( .A(core_loop_ctr_reg_1_), .B(core_compression_rounds_1_), .Y(core__abc_22172_new_n1193_));
AND2X2 AND2X2_1434 ( .A(core__abc_22172_new_n1194_), .B(core__abc_22172_new_n1179_), .Y(core__abc_22172_new_n1195_));
AND2X2 AND2X2_1435 ( .A(core__abc_22172_new_n1196_), .B(core__abc_22172_new_n1197_), .Y(core__abc_22172_new_n1198_));
AND2X2 AND2X2_1436 ( .A(core__abc_22172_new_n1198_), .B(core__abc_22172_new_n1191_), .Y(core__abc_22172_new_n1199_));
AND2X2 AND2X2_1437 ( .A(core__abc_22172_new_n1188_), .B(core__abc_22172_new_n1199_), .Y(core__abc_22172_new_n1200_));
AND2X2 AND2X2_1438 ( .A(core__abc_22172_new_n1183_), .B(core__abc_22172_new_n1201_), .Y(core__abc_22172_new_n1202_));
AND2X2 AND2X2_1439 ( .A(core__abc_22172_new_n1204_), .B(core__abc_22172_new_n1206_), .Y(core__abc_22172_new_n1207_));
AND2X2 AND2X2_144 ( .A(_abc_19873_new_n912_), .B(word3_reg_8_), .Y(_abc_19873_new_n1117_));
AND2X2 AND2X2_1440 ( .A(core__abc_22172_new_n1185_), .B(core__abc_22172_new_n1142_), .Y(core__abc_22172_new_n1208_));
AND2X2 AND2X2_1441 ( .A(core__abc_22172_new_n1210_), .B(core__abc_22172_new_n1200_), .Y(core__abc_22172_new_n1211_));
AND2X2 AND2X2_1442 ( .A(core__abc_22172_new_n1211_), .B(core_siphash_ctrl_reg_4_), .Y(core__abc_22172_new_n1212_));
AND2X2 AND2X2_1443 ( .A(core__abc_22172_new_n1213_), .B(core_compress), .Y(core__abc_22172_new_n1214_));
AND2X2 AND2X2_1444 ( .A(core__abc_22172_new_n1213_), .B(core_finalize), .Y(core__abc_22172_new_n1215_));
AND2X2 AND2X2_1445 ( .A(core__abc_22172_new_n1218_), .B(core__abc_22172_new_n1172_), .Y(core__abc_22172_new_n1219_));
AND2X2 AND2X2_1446 ( .A(core__abc_22172_new_n1219_), .B(core__abc_22172_new_n1216_), .Y(core__abc_22172_new_n1220_));
AND2X2 AND2X2_1447 ( .A(core_siphash_ctrl_reg_0_), .B(reset_n), .Y(core__abc_22172_new_n1228_));
AND2X2 AND2X2_1448 ( .A(core__abc_22172_new_n1227_), .B(core__abc_22172_new_n1228_), .Y(core__abc_22172_new_n1229_));
AND2X2 AND2X2_1449 ( .A(core__abc_22172_new_n1230_), .B(core_siphash_ctrl_reg_4_), .Y(core__abc_22172_new_n1231_));
AND2X2 AND2X2_145 ( .A(_abc_19873_new_n928_), .B(core_key_40_), .Y(_abc_19873_new_n1118_));
AND2X2 AND2X2_1450 ( .A(core__abc_22172_new_n1232_), .B(core__abc_22172_new_n1166_), .Y(core__abc_22172_new_n1233_));
AND2X2 AND2X2_1451 ( .A(core_siphash_ctrl_reg_0_), .B(core_initalize), .Y(core__abc_22172_new_n1234_));
AND2X2 AND2X2_1452 ( .A(core__abc_22172_new_n1236_), .B(core__abc_22172_new_n1222_), .Y(core__abc_22172_new_n1237_));
AND2X2 AND2X2_1453 ( .A(core_siphash_ctrl_reg_5_), .B(reset_n), .Y(core__abc_22172_new_n1243_));
AND2X2 AND2X2_1454 ( .A(core__abc_22172_new_n1223_), .B(reset_n), .Y(core__abc_22172_new_n1244_));
AND2X2 AND2X2_1455 ( .A(core__abc_22172_new_n1244_), .B(core_siphash_ctrl_reg_3_), .Y(core__abc_22172_new_n1245_));
AND2X2 AND2X2_1456 ( .A(core__abc_22172_new_n1244_), .B(core_siphash_ctrl_reg_4_), .Y(core__abc_22172_new_n1247_));
AND2X2 AND2X2_1457 ( .A(core__abc_22172_new_n1222_), .B(core__abc_22172_new_n1228_), .Y(core__abc_22172_new_n1248_));
AND2X2 AND2X2_1458 ( .A(core__abc_22172_new_n1248_), .B(core__abc_22172_new_n1214_), .Y(core__abc_22172_new_n1249_));
AND2X2 AND2X2_1459 ( .A(core__abc_22172_new_n1244_), .B(core_siphash_ctrl_reg_6_), .Y(core__abc_22172_new_n1251_));
AND2X2 AND2X2_146 ( .A(_abc_19873_new_n901_), .B(core_key_8_), .Y(_abc_19873_new_n1119_));
AND2X2 AND2X2_1460 ( .A(core__abc_22172_new_n1215_), .B(core__abc_22172_new_n1252_), .Y(core__abc_22172_new_n1253_));
AND2X2 AND2X2_1461 ( .A(core__abc_22172_new_n1248_), .B(core__abc_22172_new_n1253_), .Y(core__abc_22172_new_n1254_));
AND2X2 AND2X2_1462 ( .A(core_v1_reg_0_), .B(core_v0_reg_0_), .Y(core__abc_22172_new_n1258_));
AND2X2 AND2X2_1463 ( .A(core__abc_22172_new_n1259_), .B(core__abc_22172_new_n1257_), .Y(core__abc_22172_new_n1260_));
AND2X2 AND2X2_1464 ( .A(core__abc_22172_new_n1261_), .B(core__abc_22172_new_n1262_), .Y(core__abc_22172_new_n1263_));
AND2X2 AND2X2_1465 ( .A(core_v2_reg_0_), .B(core_v3_reg_0_), .Y(core__abc_22172_new_n1264_));
AND2X2 AND2X2_1466 ( .A(core__abc_22172_new_n1267_), .B(core__abc_22172_new_n1269_), .Y(core__abc_22172_new_n1270_));
AND2X2 AND2X2_1467 ( .A(core__abc_22172_new_n1272_), .B(reset_n), .Y(core__abc_22172_new_n1273_));
AND2X2 AND2X2_1468 ( .A(core__abc_22172_new_n1271_), .B(core__abc_22172_new_n1273_), .Y(core__0siphash_word1_reg_63_0__0_));
AND2X2 AND2X2_1469 ( .A(core_v1_reg_1_), .B(core_v0_reg_1_), .Y(core__abc_22172_new_n1276_));
AND2X2 AND2X2_147 ( .A(_abc_19873_new_n919_), .B(core_mi_40_), .Y(_abc_19873_new_n1121_));
AND2X2 AND2X2_1470 ( .A(core__abc_22172_new_n1277_), .B(core__abc_22172_new_n1275_), .Y(core__abc_22172_new_n1278_));
AND2X2 AND2X2_1471 ( .A(core_v2_reg_1_), .B(core_v3_reg_1_), .Y(core__abc_22172_new_n1279_));
AND2X2 AND2X2_1472 ( .A(core__abc_22172_new_n1280_), .B(core__abc_22172_new_n1281_), .Y(core__abc_22172_new_n1282_));
AND2X2 AND2X2_1473 ( .A(core__abc_22172_new_n1286_), .B(core__abc_22172_new_n1287_), .Y(core__abc_22172_new_n1288_));
AND2X2 AND2X2_1474 ( .A(core__abc_22172_new_n1285_), .B(core__abc_22172_new_n1290_), .Y(core__abc_22172_new_n1291_));
AND2X2 AND2X2_1475 ( .A(core__abc_22172_new_n1293_), .B(reset_n), .Y(core__abc_22172_new_n1294_));
AND2X2 AND2X2_1476 ( .A(core__abc_22172_new_n1292_), .B(core__abc_22172_new_n1294_), .Y(core__0siphash_word1_reg_63_0__1_));
AND2X2 AND2X2_1477 ( .A(core_v1_reg_2_), .B(core_v0_reg_2_), .Y(core__abc_22172_new_n1296_));
AND2X2 AND2X2_1478 ( .A(core__abc_22172_new_n1297_), .B(core__abc_22172_new_n1298_), .Y(core__abc_22172_new_n1299_));
AND2X2 AND2X2_1479 ( .A(core_v2_reg_2_), .B(core_v3_reg_2_), .Y(core__abc_22172_new_n1301_));
AND2X2 AND2X2_148 ( .A(_abc_19873_new_n888_), .B(core_mi_8_), .Y(_abc_19873_new_n1122_));
AND2X2 AND2X2_1480 ( .A(core__abc_22172_new_n1302_), .B(core__abc_22172_new_n1303_), .Y(core__abc_22172_new_n1304_));
AND2X2 AND2X2_1481 ( .A(core__abc_22172_new_n1306_), .B(core__abc_22172_new_n1300_), .Y(core__abc_22172_new_n1307_));
AND2X2 AND2X2_1482 ( .A(core__abc_22172_new_n1305_), .B(core__abc_22172_new_n1299_), .Y(core__abc_22172_new_n1308_));
AND2X2 AND2X2_1483 ( .A(core__abc_22172_new_n1311_), .B(reset_n), .Y(core__abc_22172_new_n1312_));
AND2X2 AND2X2_1484 ( .A(core__abc_22172_new_n1310_), .B(core__abc_22172_new_n1312_), .Y(core__0siphash_word1_reg_63_0__2_));
AND2X2 AND2X2_1485 ( .A(core_v1_reg_3_), .B(core_v0_reg_3_), .Y(core__abc_22172_new_n1315_));
AND2X2 AND2X2_1486 ( .A(core__abc_22172_new_n1316_), .B(core__abc_22172_new_n1314_), .Y(core__abc_22172_new_n1317_));
AND2X2 AND2X2_1487 ( .A(core_v2_reg_3_), .B(core_v3_reg_3_), .Y(core__abc_22172_new_n1318_));
AND2X2 AND2X2_1488 ( .A(core__abc_22172_new_n1319_), .B(core__abc_22172_new_n1320_), .Y(core__abc_22172_new_n1321_));
AND2X2 AND2X2_1489 ( .A(core__abc_22172_new_n1324_), .B(core__abc_22172_new_n1326_), .Y(core__abc_22172_new_n1327_));
AND2X2 AND2X2_149 ( .A(_abc_19873_new_n1126_), .B(_abc_19873_new_n937_), .Y(\read_data[8] ));
AND2X2 AND2X2_1490 ( .A(core__abc_22172_new_n1329_), .B(reset_n), .Y(core__abc_22172_new_n1330_));
AND2X2 AND2X2_1491 ( .A(core__abc_22172_new_n1328_), .B(core__abc_22172_new_n1330_), .Y(core__0siphash_word1_reg_63_0__3_));
AND2X2 AND2X2_1492 ( .A(core_v1_reg_4_), .B(core_v0_reg_4_), .Y(core__abc_22172_new_n1333_));
AND2X2 AND2X2_1493 ( .A(core__abc_22172_new_n1334_), .B(core__abc_22172_new_n1332_), .Y(core__abc_22172_new_n1335_));
AND2X2 AND2X2_1494 ( .A(core_v2_reg_4_), .B(core_v3_reg_4_), .Y(core__abc_22172_new_n1336_));
AND2X2 AND2X2_1495 ( .A(core__abc_22172_new_n1337_), .B(core__abc_22172_new_n1338_), .Y(core__abc_22172_new_n1339_));
AND2X2 AND2X2_1496 ( .A(core__abc_22172_new_n1342_), .B(core__abc_22172_new_n1344_), .Y(core__abc_22172_new_n1345_));
AND2X2 AND2X2_1497 ( .A(core__abc_22172_new_n1347_), .B(reset_n), .Y(core__abc_22172_new_n1348_));
AND2X2 AND2X2_1498 ( .A(core__abc_22172_new_n1346_), .B(core__abc_22172_new_n1348_), .Y(core__0siphash_word1_reg_63_0__4_));
AND2X2 AND2X2_1499 ( .A(core_v1_reg_5_), .B(core_v0_reg_5_), .Y(core__abc_22172_new_n1351_));
AND2X2 AND2X2_15 ( .A(_abc_19873_new_n872_), .B(_abc_19873_new_n892_), .Y(_abc_19873_new_n893_));
AND2X2 AND2X2_150 ( .A(_abc_19873_new_n881_), .B(core_key_105_), .Y(_abc_19873_new_n1128_));
AND2X2 AND2X2_1500 ( .A(core__abc_22172_new_n1352_), .B(core__abc_22172_new_n1350_), .Y(core__abc_22172_new_n1353_));
AND2X2 AND2X2_1501 ( .A(core_v2_reg_5_), .B(core_v3_reg_5_), .Y(core__abc_22172_new_n1354_));
AND2X2 AND2X2_1502 ( .A(core__abc_22172_new_n1356_), .B(core__abc_22172_new_n1357_), .Y(core__abc_22172_new_n1358_));
AND2X2 AND2X2_1503 ( .A(core__abc_22172_new_n1359_), .B(core__abc_22172_new_n1355_), .Y(core__abc_22172_new_n1360_));
AND2X2 AND2X2_1504 ( .A(core__abc_22172_new_n1364_), .B(core__abc_22172_new_n1361_), .Y(core__abc_22172_new_n1365_));
AND2X2 AND2X2_1505 ( .A(core__abc_22172_new_n1367_), .B(reset_n), .Y(core__abc_22172_new_n1368_));
AND2X2 AND2X2_1506 ( .A(core__abc_22172_new_n1366_), .B(core__abc_22172_new_n1368_), .Y(core__0siphash_word1_reg_63_0__5_));
AND2X2 AND2X2_1507 ( .A(core_v1_reg_6_), .B(core_v0_reg_6_), .Y(core__abc_22172_new_n1371_));
AND2X2 AND2X2_1508 ( .A(core__abc_22172_new_n1372_), .B(core__abc_22172_new_n1370_), .Y(core__abc_22172_new_n1373_));
AND2X2 AND2X2_1509 ( .A(core_v2_reg_6_), .B(core_v3_reg_6_), .Y(core__abc_22172_new_n1374_));
AND2X2 AND2X2_151 ( .A(_abc_19873_new_n916_), .B(core_key_73_), .Y(_abc_19873_new_n1129_));
AND2X2 AND2X2_1510 ( .A(core__abc_22172_new_n1375_), .B(core__abc_22172_new_n1376_), .Y(core__abc_22172_new_n1377_));
AND2X2 AND2X2_1511 ( .A(core__abc_22172_new_n1380_), .B(core__abc_22172_new_n1382_), .Y(core__abc_22172_new_n1383_));
AND2X2 AND2X2_1512 ( .A(core__abc_22172_new_n1385_), .B(reset_n), .Y(core__abc_22172_new_n1386_));
AND2X2 AND2X2_1513 ( .A(core__abc_22172_new_n1384_), .B(core__abc_22172_new_n1386_), .Y(core__0siphash_word1_reg_63_0__6_));
AND2X2 AND2X2_1514 ( .A(core_v1_reg_7_), .B(core_v0_reg_7_), .Y(core__abc_22172_new_n1389_));
AND2X2 AND2X2_1515 ( .A(core__abc_22172_new_n1390_), .B(core__abc_22172_new_n1388_), .Y(core__abc_22172_new_n1391_));
AND2X2 AND2X2_1516 ( .A(core_v2_reg_7_), .B(core_v3_reg_7_), .Y(core__abc_22172_new_n1392_));
AND2X2 AND2X2_1517 ( .A(core__abc_22172_new_n1394_), .B(core__abc_22172_new_n1395_), .Y(core__abc_22172_new_n1396_));
AND2X2 AND2X2_1518 ( .A(core__abc_22172_new_n1397_), .B(core__abc_22172_new_n1393_), .Y(core__abc_22172_new_n1398_));
AND2X2 AND2X2_1519 ( .A(core__abc_22172_new_n1402_), .B(core__abc_22172_new_n1399_), .Y(core__abc_22172_new_n1403_));
AND2X2 AND2X2_152 ( .A(_abc_19873_new_n912_), .B(word3_reg_9_), .Y(_abc_19873_new_n1131_));
AND2X2 AND2X2_1520 ( .A(core__abc_22172_new_n1405_), .B(reset_n), .Y(core__abc_22172_new_n1406_));
AND2X2 AND2X2_1521 ( .A(core__abc_22172_new_n1404_), .B(core__abc_22172_new_n1406_), .Y(core__0siphash_word1_reg_63_0__7_));
AND2X2 AND2X2_1522 ( .A(core_v1_reg_8_), .B(core_v0_reg_8_), .Y(core__abc_22172_new_n1409_));
AND2X2 AND2X2_1523 ( .A(core__abc_22172_new_n1410_), .B(core__abc_22172_new_n1408_), .Y(core__abc_22172_new_n1411_));
AND2X2 AND2X2_1524 ( .A(core_v2_reg_8_), .B(core_v3_reg_8_), .Y(core__abc_22172_new_n1412_));
AND2X2 AND2X2_1525 ( .A(core__abc_22172_new_n1413_), .B(core__abc_22172_new_n1414_), .Y(core__abc_22172_new_n1415_));
AND2X2 AND2X2_1526 ( .A(core__abc_22172_new_n1419_), .B(core__abc_22172_new_n1416_), .Y(core__abc_22172_new_n1420_));
AND2X2 AND2X2_1527 ( .A(core__abc_22172_new_n1422_), .B(reset_n), .Y(core__abc_22172_new_n1423_));
AND2X2 AND2X2_1528 ( .A(core__abc_22172_new_n1421_), .B(core__abc_22172_new_n1423_), .Y(core__0siphash_word1_reg_63_0__8_));
AND2X2 AND2X2_1529 ( .A(core_v1_reg_9_), .B(core_v0_reg_9_), .Y(core__abc_22172_new_n1426_));
AND2X2 AND2X2_153 ( .A(_abc_19873_new_n907_), .B(word1_reg_9_), .Y(_abc_19873_new_n1132_));
AND2X2 AND2X2_1530 ( .A(core__abc_22172_new_n1427_), .B(core__abc_22172_new_n1425_), .Y(core__abc_22172_new_n1428_));
AND2X2 AND2X2_1531 ( .A(core_v2_reg_9_), .B(core_v3_reg_9_), .Y(core__abc_22172_new_n1429_));
AND2X2 AND2X2_1532 ( .A(core__abc_22172_new_n1430_), .B(core__abc_22172_new_n1431_), .Y(core__abc_22172_new_n1432_));
AND2X2 AND2X2_1533 ( .A(core__abc_22172_new_n1436_), .B(core__abc_22172_new_n1433_), .Y(core__abc_22172_new_n1437_));
AND2X2 AND2X2_1534 ( .A(core__abc_22172_new_n1439_), .B(reset_n), .Y(core__abc_22172_new_n1440_));
AND2X2 AND2X2_1535 ( .A(core__abc_22172_new_n1438_), .B(core__abc_22172_new_n1440_), .Y(core__0siphash_word1_reg_63_0__9_));
AND2X2 AND2X2_1536 ( .A(core_v1_reg_10_), .B(core_v0_reg_10_), .Y(core__abc_22172_new_n1443_));
AND2X2 AND2X2_1537 ( .A(core__abc_22172_new_n1444_), .B(core__abc_22172_new_n1442_), .Y(core__abc_22172_new_n1445_));
AND2X2 AND2X2_1538 ( .A(core_v2_reg_10_), .B(core_v3_reg_10_), .Y(core__abc_22172_new_n1446_));
AND2X2 AND2X2_1539 ( .A(core__abc_22172_new_n1447_), .B(core__abc_22172_new_n1448_), .Y(core__abc_22172_new_n1449_));
AND2X2 AND2X2_154 ( .A(_abc_19873_new_n930_), .B(word0_reg_9_), .Y(_abc_19873_new_n1133_));
AND2X2 AND2X2_1540 ( .A(core__abc_22172_new_n1453_), .B(core__abc_22172_new_n1450_), .Y(core__abc_22172_new_n1454_));
AND2X2 AND2X2_1541 ( .A(core__abc_22172_new_n1456_), .B(reset_n), .Y(core__abc_22172_new_n1457_));
AND2X2 AND2X2_1542 ( .A(core__abc_22172_new_n1455_), .B(core__abc_22172_new_n1457_), .Y(core__0siphash_word1_reg_63_0__10_));
AND2X2 AND2X2_1543 ( .A(core_v1_reg_11_), .B(core_v0_reg_11_), .Y(core__abc_22172_new_n1460_));
AND2X2 AND2X2_1544 ( .A(core__abc_22172_new_n1461_), .B(core__abc_22172_new_n1459_), .Y(core__abc_22172_new_n1462_));
AND2X2 AND2X2_1545 ( .A(core_v2_reg_11_), .B(core_v3_reg_11_), .Y(core__abc_22172_new_n1463_));
AND2X2 AND2X2_1546 ( .A(core__abc_22172_new_n1464_), .B(core__abc_22172_new_n1465_), .Y(core__abc_22172_new_n1466_));
AND2X2 AND2X2_1547 ( .A(core__abc_22172_new_n1470_), .B(core__abc_22172_new_n1467_), .Y(core__abc_22172_new_n1471_));
AND2X2 AND2X2_1548 ( .A(core__abc_22172_new_n1473_), .B(reset_n), .Y(core__abc_22172_new_n1474_));
AND2X2 AND2X2_1549 ( .A(core__abc_22172_new_n1472_), .B(core__abc_22172_new_n1474_), .Y(core__0siphash_word1_reg_63_0__11_));
AND2X2 AND2X2_155 ( .A(_abc_19873_new_n925_), .B(word2_reg_9_), .Y(_abc_19873_new_n1137_));
AND2X2 AND2X2_1550 ( .A(core_v1_reg_12_), .B(core_v0_reg_12_), .Y(core__abc_22172_new_n1477_));
AND2X2 AND2X2_1551 ( .A(core__abc_22172_new_n1478_), .B(core__abc_22172_new_n1476_), .Y(core__abc_22172_new_n1479_));
AND2X2 AND2X2_1552 ( .A(core_v2_reg_12_), .B(core_v3_reg_12_), .Y(core__abc_22172_new_n1480_));
AND2X2 AND2X2_1553 ( .A(core__abc_22172_new_n1481_), .B(core__abc_22172_new_n1482_), .Y(core__abc_22172_new_n1483_));
AND2X2 AND2X2_1554 ( .A(core__abc_22172_new_n1487_), .B(core__abc_22172_new_n1484_), .Y(core__abc_22172_new_n1488_));
AND2X2 AND2X2_1555 ( .A(core__abc_22172_new_n1490_), .B(reset_n), .Y(core__abc_22172_new_n1491_));
AND2X2 AND2X2_1556 ( .A(core__abc_22172_new_n1489_), .B(core__abc_22172_new_n1491_), .Y(core__0siphash_word1_reg_63_0__12_));
AND2X2 AND2X2_1557 ( .A(core_v1_reg_13_), .B(core_v0_reg_13_), .Y(core__abc_22172_new_n1494_));
AND2X2 AND2X2_1558 ( .A(core__abc_22172_new_n1495_), .B(core__abc_22172_new_n1493_), .Y(core__abc_22172_new_n1496_));
AND2X2 AND2X2_1559 ( .A(core_v2_reg_13_), .B(core_v3_reg_13_), .Y(core__abc_22172_new_n1497_));
AND2X2 AND2X2_156 ( .A(_abc_19873_new_n928_), .B(core_key_41_), .Y(_abc_19873_new_n1138_));
AND2X2 AND2X2_1560 ( .A(core__abc_22172_new_n1498_), .B(core__abc_22172_new_n1499_), .Y(core__abc_22172_new_n1500_));
AND2X2 AND2X2_1561 ( .A(core__abc_22172_new_n1504_), .B(core__abc_22172_new_n1501_), .Y(core__abc_22172_new_n1505_));
AND2X2 AND2X2_1562 ( .A(core__abc_22172_new_n1507_), .B(reset_n), .Y(core__abc_22172_new_n1508_));
AND2X2 AND2X2_1563 ( .A(core__abc_22172_new_n1506_), .B(core__abc_22172_new_n1508_), .Y(core__0siphash_word1_reg_63_0__13_));
AND2X2 AND2X2_1564 ( .A(core_v1_reg_14_), .B(core_v0_reg_14_), .Y(core__abc_22172_new_n1511_));
AND2X2 AND2X2_1565 ( .A(core__abc_22172_new_n1512_), .B(core__abc_22172_new_n1510_), .Y(core__abc_22172_new_n1513_));
AND2X2 AND2X2_1566 ( .A(core_v2_reg_14_), .B(core_v3_reg_14_), .Y(core__abc_22172_new_n1514_));
AND2X2 AND2X2_1567 ( .A(core__abc_22172_new_n1515_), .B(core__abc_22172_new_n1516_), .Y(core__abc_22172_new_n1517_));
AND2X2 AND2X2_1568 ( .A(core__abc_22172_new_n1521_), .B(core__abc_22172_new_n1518_), .Y(core__abc_22172_new_n1522_));
AND2X2 AND2X2_1569 ( .A(core__abc_22172_new_n1524_), .B(reset_n), .Y(core__abc_22172_new_n1525_));
AND2X2 AND2X2_157 ( .A(_abc_19873_new_n901_), .B(core_key_9_), .Y(_abc_19873_new_n1139_));
AND2X2 AND2X2_1570 ( .A(core__abc_22172_new_n1523_), .B(core__abc_22172_new_n1525_), .Y(core__0siphash_word1_reg_63_0__14_));
AND2X2 AND2X2_1571 ( .A(core_v1_reg_15_), .B(core_v0_reg_15_), .Y(core__abc_22172_new_n1528_));
AND2X2 AND2X2_1572 ( .A(core__abc_22172_new_n1529_), .B(core__abc_22172_new_n1527_), .Y(core__abc_22172_new_n1530_));
AND2X2 AND2X2_1573 ( .A(core_v2_reg_15_), .B(core_v3_reg_15_), .Y(core__abc_22172_new_n1531_));
AND2X2 AND2X2_1574 ( .A(core__abc_22172_new_n1532_), .B(core__abc_22172_new_n1533_), .Y(core__abc_22172_new_n1534_));
AND2X2 AND2X2_1575 ( .A(core__abc_22172_new_n1538_), .B(core__abc_22172_new_n1535_), .Y(core__abc_22172_new_n1539_));
AND2X2 AND2X2_1576 ( .A(core__abc_22172_new_n1541_), .B(reset_n), .Y(core__abc_22172_new_n1542_));
AND2X2 AND2X2_1577 ( .A(core__abc_22172_new_n1540_), .B(core__abc_22172_new_n1542_), .Y(core__0siphash_word1_reg_63_0__15_));
AND2X2 AND2X2_1578 ( .A(core_v1_reg_16_), .B(core_v0_reg_16_), .Y(core__abc_22172_new_n1545_));
AND2X2 AND2X2_1579 ( .A(core__abc_22172_new_n1546_), .B(core__abc_22172_new_n1544_), .Y(core__abc_22172_new_n1547_));
AND2X2 AND2X2_158 ( .A(_abc_19873_new_n888_), .B(core_mi_9_), .Y(_abc_19873_new_n1141_));
AND2X2 AND2X2_1580 ( .A(core_v2_reg_16_), .B(core_v3_reg_16_), .Y(core__abc_22172_new_n1548_));
AND2X2 AND2X2_1581 ( .A(core__abc_22172_new_n1549_), .B(core__abc_22172_new_n1550_), .Y(core__abc_22172_new_n1551_));
AND2X2 AND2X2_1582 ( .A(core__abc_22172_new_n1555_), .B(core__abc_22172_new_n1552_), .Y(core__abc_22172_new_n1556_));
AND2X2 AND2X2_1583 ( .A(core__abc_22172_new_n1558_), .B(reset_n), .Y(core__abc_22172_new_n1559_));
AND2X2 AND2X2_1584 ( .A(core__abc_22172_new_n1557_), .B(core__abc_22172_new_n1559_), .Y(core__0siphash_word1_reg_63_0__16_));
AND2X2 AND2X2_1585 ( .A(core_v1_reg_17_), .B(core_v0_reg_17_), .Y(core__abc_22172_new_n1562_));
AND2X2 AND2X2_1586 ( .A(core__abc_22172_new_n1563_), .B(core__abc_22172_new_n1561_), .Y(core__abc_22172_new_n1564_));
AND2X2 AND2X2_1587 ( .A(core_v2_reg_17_), .B(core_v3_reg_17_), .Y(core__abc_22172_new_n1565_));
AND2X2 AND2X2_1588 ( .A(core__abc_22172_new_n1566_), .B(core__abc_22172_new_n1567_), .Y(core__abc_22172_new_n1568_));
AND2X2 AND2X2_1589 ( .A(core__abc_22172_new_n1572_), .B(core__abc_22172_new_n1569_), .Y(core__abc_22172_new_n1573_));
AND2X2 AND2X2_159 ( .A(_abc_19873_new_n919_), .B(core_mi_41_), .Y(_abc_19873_new_n1142_));
AND2X2 AND2X2_1590 ( .A(core__abc_22172_new_n1575_), .B(reset_n), .Y(core__abc_22172_new_n1576_));
AND2X2 AND2X2_1591 ( .A(core__abc_22172_new_n1574_), .B(core__abc_22172_new_n1576_), .Y(core__0siphash_word1_reg_63_0__17_));
AND2X2 AND2X2_1592 ( .A(core_v1_reg_18_), .B(core_v0_reg_18_), .Y(core__abc_22172_new_n1579_));
AND2X2 AND2X2_1593 ( .A(core__abc_22172_new_n1580_), .B(core__abc_22172_new_n1578_), .Y(core__abc_22172_new_n1581_));
AND2X2 AND2X2_1594 ( .A(core_v2_reg_18_), .B(core_v3_reg_18_), .Y(core__abc_22172_new_n1582_));
AND2X2 AND2X2_1595 ( .A(core__abc_22172_new_n1583_), .B(core__abc_22172_new_n1584_), .Y(core__abc_22172_new_n1585_));
AND2X2 AND2X2_1596 ( .A(core__abc_22172_new_n1589_), .B(core__abc_22172_new_n1586_), .Y(core__abc_22172_new_n1590_));
AND2X2 AND2X2_1597 ( .A(core__abc_22172_new_n1592_), .B(reset_n), .Y(core__abc_22172_new_n1593_));
AND2X2 AND2X2_1598 ( .A(core__abc_22172_new_n1591_), .B(core__abc_22172_new_n1593_), .Y(core__0siphash_word1_reg_63_0__18_));
AND2X2 AND2X2_1599 ( .A(core_v1_reg_19_), .B(core_v0_reg_19_), .Y(core__abc_22172_new_n1596_));
AND2X2 AND2X2_16 ( .A(_abc_19873_new_n893_), .B(_abc_19873_new_n887_), .Y(_abc_19873_new_n894_));
AND2X2 AND2X2_160 ( .A(_abc_19873_new_n1146_), .B(_abc_19873_new_n937_), .Y(\read_data[9] ));
AND2X2 AND2X2_1600 ( .A(core__abc_22172_new_n1597_), .B(core__abc_22172_new_n1595_), .Y(core__abc_22172_new_n1598_));
AND2X2 AND2X2_1601 ( .A(core_v2_reg_19_), .B(core_v3_reg_19_), .Y(core__abc_22172_new_n1599_));
AND2X2 AND2X2_1602 ( .A(core__abc_22172_new_n1600_), .B(core__abc_22172_new_n1601_), .Y(core__abc_22172_new_n1602_));
AND2X2 AND2X2_1603 ( .A(core__abc_22172_new_n1606_), .B(core__abc_22172_new_n1603_), .Y(core__abc_22172_new_n1607_));
AND2X2 AND2X2_1604 ( .A(core__abc_22172_new_n1609_), .B(reset_n), .Y(core__abc_22172_new_n1610_));
AND2X2 AND2X2_1605 ( .A(core__abc_22172_new_n1608_), .B(core__abc_22172_new_n1610_), .Y(core__0siphash_word1_reg_63_0__19_));
AND2X2 AND2X2_1606 ( .A(core_v1_reg_20_), .B(core_v0_reg_20_), .Y(core__abc_22172_new_n1613_));
AND2X2 AND2X2_1607 ( .A(core__abc_22172_new_n1614_), .B(core__abc_22172_new_n1612_), .Y(core__abc_22172_new_n1615_));
AND2X2 AND2X2_1608 ( .A(core_v2_reg_20_), .B(core_v3_reg_20_), .Y(core__abc_22172_new_n1616_));
AND2X2 AND2X2_1609 ( .A(core__abc_22172_new_n1617_), .B(core__abc_22172_new_n1618_), .Y(core__abc_22172_new_n1619_));
AND2X2 AND2X2_161 ( .A(_abc_19873_new_n881_), .B(core_key_106_), .Y(_abc_19873_new_n1148_));
AND2X2 AND2X2_1610 ( .A(core__abc_22172_new_n1623_), .B(core__abc_22172_new_n1620_), .Y(core__abc_22172_new_n1624_));
AND2X2 AND2X2_1611 ( .A(core__abc_22172_new_n1626_), .B(reset_n), .Y(core__abc_22172_new_n1627_));
AND2X2 AND2X2_1612 ( .A(core__abc_22172_new_n1625_), .B(core__abc_22172_new_n1627_), .Y(core__0siphash_word1_reg_63_0__20_));
AND2X2 AND2X2_1613 ( .A(core_v1_reg_21_), .B(core_v0_reg_21_), .Y(core__abc_22172_new_n1630_));
AND2X2 AND2X2_1614 ( .A(core__abc_22172_new_n1631_), .B(core__abc_22172_new_n1629_), .Y(core__abc_22172_new_n1632_));
AND2X2 AND2X2_1615 ( .A(core_v2_reg_21_), .B(core_v3_reg_21_), .Y(core__abc_22172_new_n1633_));
AND2X2 AND2X2_1616 ( .A(core__abc_22172_new_n1634_), .B(core__abc_22172_new_n1635_), .Y(core__abc_22172_new_n1636_));
AND2X2 AND2X2_1617 ( .A(core__abc_22172_new_n1640_), .B(core__abc_22172_new_n1637_), .Y(core__abc_22172_new_n1641_));
AND2X2 AND2X2_1618 ( .A(core__abc_22172_new_n1643_), .B(reset_n), .Y(core__abc_22172_new_n1644_));
AND2X2 AND2X2_1619 ( .A(core__abc_22172_new_n1642_), .B(core__abc_22172_new_n1644_), .Y(core__0siphash_word1_reg_63_0__21_));
AND2X2 AND2X2_162 ( .A(_abc_19873_new_n916_), .B(core_key_74_), .Y(_abc_19873_new_n1149_));
AND2X2 AND2X2_1620 ( .A(core_v1_reg_22_), .B(core_v0_reg_22_), .Y(core__abc_22172_new_n1647_));
AND2X2 AND2X2_1621 ( .A(core__abc_22172_new_n1648_), .B(core__abc_22172_new_n1646_), .Y(core__abc_22172_new_n1649_));
AND2X2 AND2X2_1622 ( .A(core_v2_reg_22_), .B(core_v3_reg_22_), .Y(core__abc_22172_new_n1650_));
AND2X2 AND2X2_1623 ( .A(core__abc_22172_new_n1651_), .B(core__abc_22172_new_n1652_), .Y(core__abc_22172_new_n1653_));
AND2X2 AND2X2_1624 ( .A(core__abc_22172_new_n1657_), .B(core__abc_22172_new_n1654_), .Y(core__abc_22172_new_n1658_));
AND2X2 AND2X2_1625 ( .A(core__abc_22172_new_n1660_), .B(reset_n), .Y(core__abc_22172_new_n1661_));
AND2X2 AND2X2_1626 ( .A(core__abc_22172_new_n1659_), .B(core__abc_22172_new_n1661_), .Y(core__0siphash_word1_reg_63_0__22_));
AND2X2 AND2X2_1627 ( .A(core_v1_reg_23_), .B(core_v0_reg_23_), .Y(core__abc_22172_new_n1664_));
AND2X2 AND2X2_1628 ( .A(core__abc_22172_new_n1665_), .B(core__abc_22172_new_n1663_), .Y(core__abc_22172_new_n1666_));
AND2X2 AND2X2_1629 ( .A(core_v2_reg_23_), .B(core_v3_reg_23_), .Y(core__abc_22172_new_n1667_));
AND2X2 AND2X2_163 ( .A(_abc_19873_new_n925_), .B(word2_reg_10_), .Y(_abc_19873_new_n1151_));
AND2X2 AND2X2_1630 ( .A(core__abc_22172_new_n1668_), .B(core__abc_22172_new_n1669_), .Y(core__abc_22172_new_n1670_));
AND2X2 AND2X2_1631 ( .A(core__abc_22172_new_n1674_), .B(core__abc_22172_new_n1671_), .Y(core__abc_22172_new_n1675_));
AND2X2 AND2X2_1632 ( .A(core__abc_22172_new_n1677_), .B(reset_n), .Y(core__abc_22172_new_n1678_));
AND2X2 AND2X2_1633 ( .A(core__abc_22172_new_n1676_), .B(core__abc_22172_new_n1678_), .Y(core__0siphash_word1_reg_63_0__23_));
AND2X2 AND2X2_1634 ( .A(core_v1_reg_24_), .B(core_v0_reg_24_), .Y(core__abc_22172_new_n1681_));
AND2X2 AND2X2_1635 ( .A(core__abc_22172_new_n1682_), .B(core__abc_22172_new_n1680_), .Y(core__abc_22172_new_n1683_));
AND2X2 AND2X2_1636 ( .A(core_v2_reg_24_), .B(core_v3_reg_24_), .Y(core__abc_22172_new_n1684_));
AND2X2 AND2X2_1637 ( .A(core__abc_22172_new_n1685_), .B(core__abc_22172_new_n1686_), .Y(core__abc_22172_new_n1687_));
AND2X2 AND2X2_1638 ( .A(core__abc_22172_new_n1691_), .B(core__abc_22172_new_n1688_), .Y(core__abc_22172_new_n1692_));
AND2X2 AND2X2_1639 ( .A(core__abc_22172_new_n1694_), .B(reset_n), .Y(core__abc_22172_new_n1695_));
AND2X2 AND2X2_164 ( .A(_abc_19873_new_n907_), .B(word1_reg_10_), .Y(_abc_19873_new_n1152_));
AND2X2 AND2X2_1640 ( .A(core__abc_22172_new_n1693_), .B(core__abc_22172_new_n1695_), .Y(core__0siphash_word1_reg_63_0__24_));
AND2X2 AND2X2_1641 ( .A(core_v1_reg_25_), .B(core_v0_reg_25_), .Y(core__abc_22172_new_n1698_));
AND2X2 AND2X2_1642 ( .A(core__abc_22172_new_n1699_), .B(core__abc_22172_new_n1697_), .Y(core__abc_22172_new_n1700_));
AND2X2 AND2X2_1643 ( .A(core_v2_reg_25_), .B(core_v3_reg_25_), .Y(core__abc_22172_new_n1701_));
AND2X2 AND2X2_1644 ( .A(core__abc_22172_new_n1702_), .B(core__abc_22172_new_n1703_), .Y(core__abc_22172_new_n1704_));
AND2X2 AND2X2_1645 ( .A(core__abc_22172_new_n1708_), .B(core__abc_22172_new_n1705_), .Y(core__abc_22172_new_n1709_));
AND2X2 AND2X2_1646 ( .A(core__abc_22172_new_n1711_), .B(reset_n), .Y(core__abc_22172_new_n1712_));
AND2X2 AND2X2_1647 ( .A(core__abc_22172_new_n1710_), .B(core__abc_22172_new_n1712_), .Y(core__0siphash_word1_reg_63_0__25_));
AND2X2 AND2X2_1648 ( .A(core_v1_reg_26_), .B(core_v0_reg_26_), .Y(core__abc_22172_new_n1715_));
AND2X2 AND2X2_1649 ( .A(core__abc_22172_new_n1716_), .B(core__abc_22172_new_n1714_), .Y(core__abc_22172_new_n1717_));
AND2X2 AND2X2_165 ( .A(_abc_19873_new_n930_), .B(word0_reg_10_), .Y(_abc_19873_new_n1153_));
AND2X2 AND2X2_1650 ( .A(core_v2_reg_26_), .B(core_v3_reg_26_), .Y(core__abc_22172_new_n1718_));
AND2X2 AND2X2_1651 ( .A(core__abc_22172_new_n1719_), .B(core__abc_22172_new_n1720_), .Y(core__abc_22172_new_n1721_));
AND2X2 AND2X2_1652 ( .A(core__abc_22172_new_n1725_), .B(core__abc_22172_new_n1722_), .Y(core__abc_22172_new_n1726_));
AND2X2 AND2X2_1653 ( .A(core__abc_22172_new_n1728_), .B(reset_n), .Y(core__abc_22172_new_n1729_));
AND2X2 AND2X2_1654 ( .A(core__abc_22172_new_n1727_), .B(core__abc_22172_new_n1729_), .Y(core__0siphash_word1_reg_63_0__26_));
AND2X2 AND2X2_1655 ( .A(core_v1_reg_27_), .B(core_v0_reg_27_), .Y(core__abc_22172_new_n1732_));
AND2X2 AND2X2_1656 ( .A(core__abc_22172_new_n1733_), .B(core__abc_22172_new_n1731_), .Y(core__abc_22172_new_n1734_));
AND2X2 AND2X2_1657 ( .A(core_v2_reg_27_), .B(core_v3_reg_27_), .Y(core__abc_22172_new_n1735_));
AND2X2 AND2X2_1658 ( .A(core__abc_22172_new_n1736_), .B(core__abc_22172_new_n1737_), .Y(core__abc_22172_new_n1738_));
AND2X2 AND2X2_1659 ( .A(core__abc_22172_new_n1742_), .B(core__abc_22172_new_n1739_), .Y(core__abc_22172_new_n1743_));
AND2X2 AND2X2_166 ( .A(_abc_19873_new_n912_), .B(word3_reg_10_), .Y(_abc_19873_new_n1157_));
AND2X2 AND2X2_1660 ( .A(core__abc_22172_new_n1745_), .B(reset_n), .Y(core__abc_22172_new_n1746_));
AND2X2 AND2X2_1661 ( .A(core__abc_22172_new_n1744_), .B(core__abc_22172_new_n1746_), .Y(core__0siphash_word1_reg_63_0__27_));
AND2X2 AND2X2_1662 ( .A(core_v1_reg_28_), .B(core_v0_reg_28_), .Y(core__abc_22172_new_n1749_));
AND2X2 AND2X2_1663 ( .A(core__abc_22172_new_n1750_), .B(core__abc_22172_new_n1748_), .Y(core__abc_22172_new_n1751_));
AND2X2 AND2X2_1664 ( .A(core_v2_reg_28_), .B(core_v3_reg_28_), .Y(core__abc_22172_new_n1752_));
AND2X2 AND2X2_1665 ( .A(core__abc_22172_new_n1753_), .B(core__abc_22172_new_n1754_), .Y(core__abc_22172_new_n1755_));
AND2X2 AND2X2_1666 ( .A(core__abc_22172_new_n1759_), .B(core__abc_22172_new_n1756_), .Y(core__abc_22172_new_n1760_));
AND2X2 AND2X2_1667 ( .A(core__abc_22172_new_n1762_), .B(reset_n), .Y(core__abc_22172_new_n1763_));
AND2X2 AND2X2_1668 ( .A(core__abc_22172_new_n1761_), .B(core__abc_22172_new_n1763_), .Y(core__0siphash_word1_reg_63_0__28_));
AND2X2 AND2X2_1669 ( .A(core_v1_reg_29_), .B(core_v0_reg_29_), .Y(core__abc_22172_new_n1766_));
AND2X2 AND2X2_167 ( .A(_abc_19873_new_n928_), .B(core_key_42_), .Y(_abc_19873_new_n1158_));
AND2X2 AND2X2_1670 ( .A(core__abc_22172_new_n1767_), .B(core__abc_22172_new_n1765_), .Y(core__abc_22172_new_n1768_));
AND2X2 AND2X2_1671 ( .A(core_v2_reg_29_), .B(core_v3_reg_29_), .Y(core__abc_22172_new_n1769_));
AND2X2 AND2X2_1672 ( .A(core__abc_22172_new_n1770_), .B(core__abc_22172_new_n1771_), .Y(core__abc_22172_new_n1772_));
AND2X2 AND2X2_1673 ( .A(core__abc_22172_new_n1776_), .B(core__abc_22172_new_n1773_), .Y(core__abc_22172_new_n1777_));
AND2X2 AND2X2_1674 ( .A(core__abc_22172_new_n1779_), .B(reset_n), .Y(core__abc_22172_new_n1780_));
AND2X2 AND2X2_1675 ( .A(core__abc_22172_new_n1778_), .B(core__abc_22172_new_n1780_), .Y(core__0siphash_word1_reg_63_0__29_));
AND2X2 AND2X2_1676 ( .A(core_v1_reg_30_), .B(core_v0_reg_30_), .Y(core__abc_22172_new_n1783_));
AND2X2 AND2X2_1677 ( .A(core__abc_22172_new_n1784_), .B(core__abc_22172_new_n1782_), .Y(core__abc_22172_new_n1785_));
AND2X2 AND2X2_1678 ( .A(core_v2_reg_30_), .B(core_v3_reg_30_), .Y(core__abc_22172_new_n1786_));
AND2X2 AND2X2_1679 ( .A(core__abc_22172_new_n1787_), .B(core__abc_22172_new_n1788_), .Y(core__abc_22172_new_n1789_));
AND2X2 AND2X2_168 ( .A(_abc_19873_new_n901_), .B(core_key_10_), .Y(_abc_19873_new_n1159_));
AND2X2 AND2X2_1680 ( .A(core__abc_22172_new_n1793_), .B(core__abc_22172_new_n1790_), .Y(core__abc_22172_new_n1794_));
AND2X2 AND2X2_1681 ( .A(core__abc_22172_new_n1796_), .B(reset_n), .Y(core__abc_22172_new_n1797_));
AND2X2 AND2X2_1682 ( .A(core__abc_22172_new_n1795_), .B(core__abc_22172_new_n1797_), .Y(core__0siphash_word1_reg_63_0__30_));
AND2X2 AND2X2_1683 ( .A(core_v1_reg_31_), .B(core_v0_reg_31_), .Y(core__abc_22172_new_n1800_));
AND2X2 AND2X2_1684 ( .A(core__abc_22172_new_n1801_), .B(core__abc_22172_new_n1799_), .Y(core__abc_22172_new_n1802_));
AND2X2 AND2X2_1685 ( .A(core_v2_reg_31_), .B(core_v3_reg_31_), .Y(core__abc_22172_new_n1803_));
AND2X2 AND2X2_1686 ( .A(core__abc_22172_new_n1804_), .B(core__abc_22172_new_n1805_), .Y(core__abc_22172_new_n1806_));
AND2X2 AND2X2_1687 ( .A(core__abc_22172_new_n1810_), .B(core__abc_22172_new_n1807_), .Y(core__abc_22172_new_n1811_));
AND2X2 AND2X2_1688 ( .A(core__abc_22172_new_n1813_), .B(reset_n), .Y(core__abc_22172_new_n1814_));
AND2X2 AND2X2_1689 ( .A(core__abc_22172_new_n1812_), .B(core__abc_22172_new_n1814_), .Y(core__0siphash_word1_reg_63_0__31_));
AND2X2 AND2X2_169 ( .A(_abc_19873_new_n919_), .B(core_mi_42_), .Y(_abc_19873_new_n1161_));
AND2X2 AND2X2_1690 ( .A(core_v1_reg_32_), .B(core_v0_reg_32_), .Y(core__abc_22172_new_n1817_));
AND2X2 AND2X2_1691 ( .A(core__abc_22172_new_n1818_), .B(core__abc_22172_new_n1816_), .Y(core__abc_22172_new_n1819_));
AND2X2 AND2X2_1692 ( .A(core_v2_reg_32_), .B(core_v3_reg_32_), .Y(core__abc_22172_new_n1820_));
AND2X2 AND2X2_1693 ( .A(core__abc_22172_new_n1821_), .B(core__abc_22172_new_n1822_), .Y(core__abc_22172_new_n1823_));
AND2X2 AND2X2_1694 ( .A(core__abc_22172_new_n1827_), .B(core__abc_22172_new_n1824_), .Y(core__abc_22172_new_n1828_));
AND2X2 AND2X2_1695 ( .A(core__abc_22172_new_n1830_), .B(reset_n), .Y(core__abc_22172_new_n1831_));
AND2X2 AND2X2_1696 ( .A(core__abc_22172_new_n1829_), .B(core__abc_22172_new_n1831_), .Y(core__0siphash_word1_reg_63_0__32_));
AND2X2 AND2X2_1697 ( .A(core_v1_reg_33_), .B(core_v0_reg_33_), .Y(core__abc_22172_new_n1834_));
AND2X2 AND2X2_1698 ( .A(core__abc_22172_new_n1835_), .B(core__abc_22172_new_n1833_), .Y(core__abc_22172_new_n1836_));
AND2X2 AND2X2_1699 ( .A(core_v2_reg_33_), .B(core_v3_reg_33_), .Y(core__abc_22172_new_n1837_));
AND2X2 AND2X2_17 ( .A(_abc_19873_new_n894_), .B(core_initalize), .Y(_abc_19873_new_n895_));
AND2X2 AND2X2_170 ( .A(_abc_19873_new_n888_), .B(core_mi_10_), .Y(_abc_19873_new_n1162_));
AND2X2 AND2X2_1700 ( .A(core__abc_22172_new_n1838_), .B(core__abc_22172_new_n1839_), .Y(core__abc_22172_new_n1840_));
AND2X2 AND2X2_1701 ( .A(core__abc_22172_new_n1844_), .B(core__abc_22172_new_n1841_), .Y(core__abc_22172_new_n1845_));
AND2X2 AND2X2_1702 ( .A(core__abc_22172_new_n1847_), .B(reset_n), .Y(core__abc_22172_new_n1848_));
AND2X2 AND2X2_1703 ( .A(core__abc_22172_new_n1846_), .B(core__abc_22172_new_n1848_), .Y(core__0siphash_word1_reg_63_0__33_));
AND2X2 AND2X2_1704 ( .A(core_v1_reg_34_), .B(core_v0_reg_34_), .Y(core__abc_22172_new_n1851_));
AND2X2 AND2X2_1705 ( .A(core__abc_22172_new_n1852_), .B(core__abc_22172_new_n1850_), .Y(core__abc_22172_new_n1853_));
AND2X2 AND2X2_1706 ( .A(core_v2_reg_34_), .B(core_v3_reg_34_), .Y(core__abc_22172_new_n1855_));
AND2X2 AND2X2_1707 ( .A(core__abc_22172_new_n1856_), .B(core__abc_22172_new_n1854_), .Y(core__abc_22172_new_n1857_));
AND2X2 AND2X2_1708 ( .A(core__abc_22172_new_n1861_), .B(core__abc_22172_new_n1858_), .Y(core__abc_22172_new_n1862_));
AND2X2 AND2X2_1709 ( .A(core__abc_22172_new_n1864_), .B(reset_n), .Y(core__abc_22172_new_n1865_));
AND2X2 AND2X2_171 ( .A(_abc_19873_new_n1166_), .B(_abc_19873_new_n937_), .Y(\read_data[10] ));
AND2X2 AND2X2_1710 ( .A(core__abc_22172_new_n1863_), .B(core__abc_22172_new_n1865_), .Y(core__0siphash_word1_reg_63_0__34_));
AND2X2 AND2X2_1711 ( .A(core_v1_reg_35_), .B(core_v0_reg_35_), .Y(core__abc_22172_new_n1868_));
AND2X2 AND2X2_1712 ( .A(core__abc_22172_new_n1869_), .B(core__abc_22172_new_n1867_), .Y(core__abc_22172_new_n1870_));
AND2X2 AND2X2_1713 ( .A(core_v2_reg_35_), .B(core_v3_reg_35_), .Y(core__abc_22172_new_n1871_));
AND2X2 AND2X2_1714 ( .A(core__abc_22172_new_n1872_), .B(core__abc_22172_new_n1873_), .Y(core__abc_22172_new_n1874_));
AND2X2 AND2X2_1715 ( .A(core__abc_22172_new_n1878_), .B(core__abc_22172_new_n1875_), .Y(core__abc_22172_new_n1879_));
AND2X2 AND2X2_1716 ( .A(core__abc_22172_new_n1881_), .B(reset_n), .Y(core__abc_22172_new_n1882_));
AND2X2 AND2X2_1717 ( .A(core__abc_22172_new_n1880_), .B(core__abc_22172_new_n1882_), .Y(core__0siphash_word1_reg_63_0__35_));
AND2X2 AND2X2_1718 ( .A(core_v1_reg_36_), .B(core_v0_reg_36_), .Y(core__abc_22172_new_n1885_));
AND2X2 AND2X2_1719 ( .A(core__abc_22172_new_n1886_), .B(core__abc_22172_new_n1884_), .Y(core__abc_22172_new_n1887_));
AND2X2 AND2X2_172 ( .A(_abc_19873_new_n912_), .B(word3_reg_11_), .Y(_abc_19873_new_n1168_));
AND2X2 AND2X2_1720 ( .A(core_v2_reg_36_), .B(core_v3_reg_36_), .Y(core__abc_22172_new_n1889_));
AND2X2 AND2X2_1721 ( .A(core__abc_22172_new_n1890_), .B(core__abc_22172_new_n1888_), .Y(core__abc_22172_new_n1891_));
AND2X2 AND2X2_1722 ( .A(core__abc_22172_new_n1895_), .B(core__abc_22172_new_n1892_), .Y(core__abc_22172_new_n1896_));
AND2X2 AND2X2_1723 ( .A(core__abc_22172_new_n1898_), .B(reset_n), .Y(core__abc_22172_new_n1899_));
AND2X2 AND2X2_1724 ( .A(core__abc_22172_new_n1897_), .B(core__abc_22172_new_n1899_), .Y(core__0siphash_word1_reg_63_0__36_));
AND2X2 AND2X2_1725 ( .A(core_v1_reg_37_), .B(core_v0_reg_37_), .Y(core__abc_22172_new_n1902_));
AND2X2 AND2X2_1726 ( .A(core__abc_22172_new_n1903_), .B(core__abc_22172_new_n1901_), .Y(core__abc_22172_new_n1904_));
AND2X2 AND2X2_1727 ( .A(core_v2_reg_37_), .B(core_v3_reg_37_), .Y(core__abc_22172_new_n1905_));
AND2X2 AND2X2_1728 ( .A(core__abc_22172_new_n1906_), .B(core__abc_22172_new_n1907_), .Y(core__abc_22172_new_n1908_));
AND2X2 AND2X2_1729 ( .A(core__abc_22172_new_n1912_), .B(core__abc_22172_new_n1909_), .Y(core__abc_22172_new_n1913_));
AND2X2 AND2X2_173 ( .A(_abc_19873_new_n901_), .B(core_key_11_), .Y(_abc_19873_new_n1169_));
AND2X2 AND2X2_1730 ( .A(core__abc_22172_new_n1915_), .B(reset_n), .Y(core__abc_22172_new_n1916_));
AND2X2 AND2X2_1731 ( .A(core__abc_22172_new_n1914_), .B(core__abc_22172_new_n1916_), .Y(core__0siphash_word1_reg_63_0__37_));
AND2X2 AND2X2_1732 ( .A(core_v1_reg_38_), .B(core_v0_reg_38_), .Y(core__abc_22172_new_n1919_));
AND2X2 AND2X2_1733 ( .A(core__abc_22172_new_n1920_), .B(core__abc_22172_new_n1918_), .Y(core__abc_22172_new_n1921_));
AND2X2 AND2X2_1734 ( .A(core_v2_reg_38_), .B(core_v3_reg_38_), .Y(core__abc_22172_new_n1923_));
AND2X2 AND2X2_1735 ( .A(core__abc_22172_new_n1924_), .B(core__abc_22172_new_n1922_), .Y(core__abc_22172_new_n1925_));
AND2X2 AND2X2_1736 ( .A(core__abc_22172_new_n1929_), .B(core__abc_22172_new_n1926_), .Y(core__abc_22172_new_n1930_));
AND2X2 AND2X2_1737 ( .A(core__abc_22172_new_n1932_), .B(reset_n), .Y(core__abc_22172_new_n1933_));
AND2X2 AND2X2_1738 ( .A(core__abc_22172_new_n1931_), .B(core__abc_22172_new_n1933_), .Y(core__0siphash_word1_reg_63_0__38_));
AND2X2 AND2X2_1739 ( .A(core_v1_reg_39_), .B(core_v0_reg_39_), .Y(core__abc_22172_new_n1936_));
AND2X2 AND2X2_174 ( .A(_abc_19873_new_n925_), .B(word2_reg_11_), .Y(_abc_19873_new_n1170_));
AND2X2 AND2X2_1740 ( .A(core__abc_22172_new_n1937_), .B(core__abc_22172_new_n1935_), .Y(core__abc_22172_new_n1938_));
AND2X2 AND2X2_1741 ( .A(core_v2_reg_39_), .B(core_v3_reg_39_), .Y(core__abc_22172_new_n1939_));
AND2X2 AND2X2_1742 ( .A(core__abc_22172_new_n1940_), .B(core__abc_22172_new_n1941_), .Y(core__abc_22172_new_n1942_));
AND2X2 AND2X2_1743 ( .A(core__abc_22172_new_n1946_), .B(core__abc_22172_new_n1943_), .Y(core__abc_22172_new_n1947_));
AND2X2 AND2X2_1744 ( .A(core__abc_22172_new_n1949_), .B(reset_n), .Y(core__abc_22172_new_n1950_));
AND2X2 AND2X2_1745 ( .A(core__abc_22172_new_n1948_), .B(core__abc_22172_new_n1950_), .Y(core__0siphash_word1_reg_63_0__39_));
AND2X2 AND2X2_1746 ( .A(core_v1_reg_40_), .B(core_v0_reg_40_), .Y(core__abc_22172_new_n1953_));
AND2X2 AND2X2_1747 ( .A(core__abc_22172_new_n1954_), .B(core__abc_22172_new_n1952_), .Y(core__abc_22172_new_n1955_));
AND2X2 AND2X2_1748 ( .A(core_v2_reg_40_), .B(core_v3_reg_40_), .Y(core__abc_22172_new_n1956_));
AND2X2 AND2X2_1749 ( .A(core__abc_22172_new_n1957_), .B(core__abc_22172_new_n1958_), .Y(core__abc_22172_new_n1959_));
AND2X2 AND2X2_175 ( .A(_abc_19873_new_n881_), .B(core_key_107_), .Y(_abc_19873_new_n1173_));
AND2X2 AND2X2_1750 ( .A(core__abc_22172_new_n1963_), .B(core__abc_22172_new_n1960_), .Y(core__abc_22172_new_n1964_));
AND2X2 AND2X2_1751 ( .A(core__abc_22172_new_n1966_), .B(reset_n), .Y(core__abc_22172_new_n1967_));
AND2X2 AND2X2_1752 ( .A(core__abc_22172_new_n1965_), .B(core__abc_22172_new_n1967_), .Y(core__0siphash_word1_reg_63_0__40_));
AND2X2 AND2X2_1753 ( .A(core_v1_reg_41_), .B(core_v0_reg_41_), .Y(core__abc_22172_new_n1970_));
AND2X2 AND2X2_1754 ( .A(core__abc_22172_new_n1971_), .B(core__abc_22172_new_n1969_), .Y(core__abc_22172_new_n1972_));
AND2X2 AND2X2_1755 ( .A(core_v2_reg_41_), .B(core_v3_reg_41_), .Y(core__abc_22172_new_n1973_));
AND2X2 AND2X2_1756 ( .A(core__abc_22172_new_n1974_), .B(core__abc_22172_new_n1975_), .Y(core__abc_22172_new_n1976_));
AND2X2 AND2X2_1757 ( .A(core__abc_22172_new_n1980_), .B(core__abc_22172_new_n1977_), .Y(core__abc_22172_new_n1981_));
AND2X2 AND2X2_1758 ( .A(core__abc_22172_new_n1983_), .B(reset_n), .Y(core__abc_22172_new_n1984_));
AND2X2 AND2X2_1759 ( .A(core__abc_22172_new_n1982_), .B(core__abc_22172_new_n1984_), .Y(core__0siphash_word1_reg_63_0__41_));
AND2X2 AND2X2_176 ( .A(_abc_19873_new_n888_), .B(core_mi_11_), .Y(_abc_19873_new_n1174_));
AND2X2 AND2X2_1760 ( .A(core_v1_reg_42_), .B(core_v0_reg_42_), .Y(core__abc_22172_new_n1987_));
AND2X2 AND2X2_1761 ( .A(core__abc_22172_new_n1988_), .B(core__abc_22172_new_n1986_), .Y(core__abc_22172_new_n1989_));
AND2X2 AND2X2_1762 ( .A(core_v2_reg_42_), .B(core_v3_reg_42_), .Y(core__abc_22172_new_n1990_));
AND2X2 AND2X2_1763 ( .A(core__abc_22172_new_n1991_), .B(core__abc_22172_new_n1992_), .Y(core__abc_22172_new_n1993_));
AND2X2 AND2X2_1764 ( .A(core__abc_22172_new_n1997_), .B(core__abc_22172_new_n1994_), .Y(core__abc_22172_new_n1998_));
AND2X2 AND2X2_1765 ( .A(core__abc_22172_new_n2000_), .B(reset_n), .Y(core__abc_22172_new_n2001_));
AND2X2 AND2X2_1766 ( .A(core__abc_22172_new_n1999_), .B(core__abc_22172_new_n2001_), .Y(core__0siphash_word1_reg_63_0__42_));
AND2X2 AND2X2_1767 ( .A(core_v1_reg_43_), .B(core_v0_reg_43_), .Y(core__abc_22172_new_n2004_));
AND2X2 AND2X2_1768 ( .A(core__abc_22172_new_n2005_), .B(core__abc_22172_new_n2003_), .Y(core__abc_22172_new_n2006_));
AND2X2 AND2X2_1769 ( .A(core_v2_reg_43_), .B(core_v3_reg_43_), .Y(core__abc_22172_new_n2008_));
AND2X2 AND2X2_177 ( .A(_abc_19873_new_n928_), .B(core_key_43_), .Y(_abc_19873_new_n1176_));
AND2X2 AND2X2_1770 ( .A(core__abc_22172_new_n2009_), .B(core__abc_22172_new_n2007_), .Y(core__abc_22172_new_n2010_));
AND2X2 AND2X2_1771 ( .A(core__abc_22172_new_n2014_), .B(core__abc_22172_new_n2011_), .Y(core__abc_22172_new_n2015_));
AND2X2 AND2X2_1772 ( .A(core__abc_22172_new_n2017_), .B(reset_n), .Y(core__abc_22172_new_n2018_));
AND2X2 AND2X2_1773 ( .A(core__abc_22172_new_n2016_), .B(core__abc_22172_new_n2018_), .Y(core__0siphash_word1_reg_63_0__43_));
AND2X2 AND2X2_1774 ( .A(core_v1_reg_44_), .B(core_v0_reg_44_), .Y(core__abc_22172_new_n2021_));
AND2X2 AND2X2_1775 ( .A(core__abc_22172_new_n2022_), .B(core__abc_22172_new_n2020_), .Y(core__abc_22172_new_n2023_));
AND2X2 AND2X2_1776 ( .A(core_v2_reg_44_), .B(core_v3_reg_44_), .Y(core__abc_22172_new_n2025_));
AND2X2 AND2X2_1777 ( .A(core__abc_22172_new_n2026_), .B(core__abc_22172_new_n2024_), .Y(core__abc_22172_new_n2027_));
AND2X2 AND2X2_1778 ( .A(core__abc_22172_new_n2031_), .B(core__abc_22172_new_n2028_), .Y(core__abc_22172_new_n2032_));
AND2X2 AND2X2_1779 ( .A(core__abc_22172_new_n2034_), .B(reset_n), .Y(core__abc_22172_new_n2035_));
AND2X2 AND2X2_178 ( .A(_abc_19873_new_n916_), .B(core_key_75_), .Y(_abc_19873_new_n1177_));
AND2X2 AND2X2_1780 ( .A(core__abc_22172_new_n2033_), .B(core__abc_22172_new_n2035_), .Y(core__0siphash_word1_reg_63_0__44_));
AND2X2 AND2X2_1781 ( .A(core_v1_reg_45_), .B(core_v0_reg_45_), .Y(core__abc_22172_new_n2038_));
AND2X2 AND2X2_1782 ( .A(core__abc_22172_new_n2039_), .B(core__abc_22172_new_n2037_), .Y(core__abc_22172_new_n2040_));
AND2X2 AND2X2_1783 ( .A(core_v2_reg_45_), .B(core_v3_reg_45_), .Y(core__abc_22172_new_n2042_));
AND2X2 AND2X2_1784 ( .A(core__abc_22172_new_n2043_), .B(core__abc_22172_new_n2041_), .Y(core__abc_22172_new_n2044_));
AND2X2 AND2X2_1785 ( .A(core__abc_22172_new_n2048_), .B(core__abc_22172_new_n2045_), .Y(core__abc_22172_new_n2049_));
AND2X2 AND2X2_1786 ( .A(core__abc_22172_new_n2051_), .B(reset_n), .Y(core__abc_22172_new_n2052_));
AND2X2 AND2X2_1787 ( .A(core__abc_22172_new_n2050_), .B(core__abc_22172_new_n2052_), .Y(core__0siphash_word1_reg_63_0__45_));
AND2X2 AND2X2_1788 ( .A(core_v1_reg_46_), .B(core_v0_reg_46_), .Y(core__abc_22172_new_n2055_));
AND2X2 AND2X2_1789 ( .A(core__abc_22172_new_n2056_), .B(core__abc_22172_new_n2054_), .Y(core__abc_22172_new_n2057_));
AND2X2 AND2X2_179 ( .A(_abc_19873_new_n930_), .B(word0_reg_11_), .Y(_abc_19873_new_n1180_));
AND2X2 AND2X2_1790 ( .A(core_v2_reg_46_), .B(core_v3_reg_46_), .Y(core__abc_22172_new_n2059_));
AND2X2 AND2X2_1791 ( .A(core__abc_22172_new_n2060_), .B(core__abc_22172_new_n2058_), .Y(core__abc_22172_new_n2061_));
AND2X2 AND2X2_1792 ( .A(core__abc_22172_new_n2065_), .B(core__abc_22172_new_n2062_), .Y(core__abc_22172_new_n2066_));
AND2X2 AND2X2_1793 ( .A(core__abc_22172_new_n2068_), .B(reset_n), .Y(core__abc_22172_new_n2069_));
AND2X2 AND2X2_1794 ( .A(core__abc_22172_new_n2067_), .B(core__abc_22172_new_n2069_), .Y(core__0siphash_word1_reg_63_0__46_));
AND2X2 AND2X2_1795 ( .A(core_v1_reg_47_), .B(core_v0_reg_47_), .Y(core__abc_22172_new_n2072_));
AND2X2 AND2X2_1796 ( .A(core__abc_22172_new_n2073_), .B(core__abc_22172_new_n2071_), .Y(core__abc_22172_new_n2074_));
AND2X2 AND2X2_1797 ( .A(core_v2_reg_47_), .B(core_v3_reg_47_), .Y(core__abc_22172_new_n2076_));
AND2X2 AND2X2_1798 ( .A(core__abc_22172_new_n2077_), .B(core__abc_22172_new_n2075_), .Y(core__abc_22172_new_n2078_));
AND2X2 AND2X2_1799 ( .A(core__abc_22172_new_n2082_), .B(core__abc_22172_new_n2079_), .Y(core__abc_22172_new_n2083_));
AND2X2 AND2X2_18 ( .A(_abc_19873_new_n886_), .B(_abc_19873_new_n876_), .Y(_abc_19873_new_n896_));
AND2X2 AND2X2_180 ( .A(_abc_19873_new_n907_), .B(word1_reg_11_), .Y(_abc_19873_new_n1181_));
AND2X2 AND2X2_1800 ( .A(core__abc_22172_new_n2085_), .B(reset_n), .Y(core__abc_22172_new_n2086_));
AND2X2 AND2X2_1801 ( .A(core__abc_22172_new_n2084_), .B(core__abc_22172_new_n2086_), .Y(core__0siphash_word1_reg_63_0__47_));
AND2X2 AND2X2_1802 ( .A(core_v1_reg_48_), .B(core_v0_reg_48_), .Y(core__abc_22172_new_n2089_));
AND2X2 AND2X2_1803 ( .A(core__abc_22172_new_n2090_), .B(core__abc_22172_new_n2088_), .Y(core__abc_22172_new_n2091_));
AND2X2 AND2X2_1804 ( .A(core_v2_reg_48_), .B(core_v3_reg_48_), .Y(core__abc_22172_new_n2093_));
AND2X2 AND2X2_1805 ( .A(core__abc_22172_new_n2094_), .B(core__abc_22172_new_n2092_), .Y(core__abc_22172_new_n2095_));
AND2X2 AND2X2_1806 ( .A(core__abc_22172_new_n2099_), .B(core__abc_22172_new_n2096_), .Y(core__abc_22172_new_n2100_));
AND2X2 AND2X2_1807 ( .A(core__abc_22172_new_n2102_), .B(reset_n), .Y(core__abc_22172_new_n2103_));
AND2X2 AND2X2_1808 ( .A(core__abc_22172_new_n2101_), .B(core__abc_22172_new_n2103_), .Y(core__0siphash_word1_reg_63_0__48_));
AND2X2 AND2X2_1809 ( .A(core_v1_reg_49_), .B(core_v0_reg_49_), .Y(core__abc_22172_new_n2105_));
AND2X2 AND2X2_181 ( .A(_abc_19873_new_n919_), .B(core_mi_43_), .Y(_abc_19873_new_n1183_));
AND2X2 AND2X2_1810 ( .A(core__abc_22172_new_n2106_), .B(core__abc_22172_new_n2107_), .Y(core__abc_22172_new_n2108_));
AND2X2 AND2X2_1811 ( .A(core_v2_reg_49_), .B(core_v3_reg_49_), .Y(core__abc_22172_new_n2111_));
AND2X2 AND2X2_1812 ( .A(core__abc_22172_new_n2112_), .B(core__abc_22172_new_n2110_), .Y(core__abc_22172_new_n2113_));
AND2X2 AND2X2_1813 ( .A(core__abc_22172_new_n2109_), .B(core__abc_22172_new_n2113_), .Y(core__abc_22172_new_n2114_));
AND2X2 AND2X2_1814 ( .A(core__abc_22172_new_n2115_), .B(core__abc_22172_new_n2108_), .Y(core__abc_22172_new_n2116_));
AND2X2 AND2X2_1815 ( .A(core__abc_22172_new_n2119_), .B(reset_n), .Y(core__abc_22172_new_n2120_));
AND2X2 AND2X2_1816 ( .A(core__abc_22172_new_n2118_), .B(core__abc_22172_new_n2120_), .Y(core__0siphash_word1_reg_63_0__49_));
AND2X2 AND2X2_1817 ( .A(core_v1_reg_50_), .B(core_v0_reg_50_), .Y(core__abc_22172_new_n2123_));
AND2X2 AND2X2_1818 ( .A(core__abc_22172_new_n2124_), .B(core__abc_22172_new_n2122_), .Y(core__abc_22172_new_n2125_));
AND2X2 AND2X2_1819 ( .A(core_v2_reg_50_), .B(core_v3_reg_50_), .Y(core__abc_22172_new_n2127_));
AND2X2 AND2X2_182 ( .A(_abc_19873_new_n1187_), .B(_abc_19873_new_n937_), .Y(\read_data[11] ));
AND2X2 AND2X2_1820 ( .A(core__abc_22172_new_n2128_), .B(core__abc_22172_new_n2126_), .Y(core__abc_22172_new_n2129_));
AND2X2 AND2X2_1821 ( .A(core__abc_22172_new_n2133_), .B(core__abc_22172_new_n2130_), .Y(core__abc_22172_new_n2134_));
AND2X2 AND2X2_1822 ( .A(core__abc_22172_new_n2136_), .B(reset_n), .Y(core__abc_22172_new_n2137_));
AND2X2 AND2X2_1823 ( .A(core__abc_22172_new_n2135_), .B(core__abc_22172_new_n2137_), .Y(core__0siphash_word1_reg_63_0__50_));
AND2X2 AND2X2_1824 ( .A(core_v1_reg_51_), .B(core_v0_reg_51_), .Y(core__abc_22172_new_n2140_));
AND2X2 AND2X2_1825 ( .A(core__abc_22172_new_n2141_), .B(core__abc_22172_new_n2139_), .Y(core__abc_22172_new_n2142_));
AND2X2 AND2X2_1826 ( .A(core_v2_reg_51_), .B(core_v3_reg_51_), .Y(core__abc_22172_new_n2144_));
AND2X2 AND2X2_1827 ( .A(core__abc_22172_new_n2145_), .B(core__abc_22172_new_n2143_), .Y(core__abc_22172_new_n2146_));
AND2X2 AND2X2_1828 ( .A(core__abc_22172_new_n2150_), .B(core__abc_22172_new_n2147_), .Y(core__abc_22172_new_n2151_));
AND2X2 AND2X2_1829 ( .A(core__abc_22172_new_n2153_), .B(reset_n), .Y(core__abc_22172_new_n2154_));
AND2X2 AND2X2_183 ( .A(_abc_19873_new_n881_), .B(core_key_108_), .Y(_abc_19873_new_n1189_));
AND2X2 AND2X2_1830 ( .A(core__abc_22172_new_n2152_), .B(core__abc_22172_new_n2154_), .Y(core__0siphash_word1_reg_63_0__51_));
AND2X2 AND2X2_1831 ( .A(core_v1_reg_52_), .B(core_v0_reg_52_), .Y(core__abc_22172_new_n2157_));
AND2X2 AND2X2_1832 ( .A(core__abc_22172_new_n2158_), .B(core__abc_22172_new_n2156_), .Y(core__abc_22172_new_n2159_));
AND2X2 AND2X2_1833 ( .A(core_v2_reg_52_), .B(core_v3_reg_52_), .Y(core__abc_22172_new_n2161_));
AND2X2 AND2X2_1834 ( .A(core__abc_22172_new_n2162_), .B(core__abc_22172_new_n2160_), .Y(core__abc_22172_new_n2163_));
AND2X2 AND2X2_1835 ( .A(core__abc_22172_new_n2167_), .B(core__abc_22172_new_n2164_), .Y(core__abc_22172_new_n2168_));
AND2X2 AND2X2_1836 ( .A(core__abc_22172_new_n2170_), .B(reset_n), .Y(core__abc_22172_new_n2171_));
AND2X2 AND2X2_1837 ( .A(core__abc_22172_new_n2169_), .B(core__abc_22172_new_n2171_), .Y(core__0siphash_word1_reg_63_0__52_));
AND2X2 AND2X2_1838 ( .A(core_v1_reg_53_), .B(core_v0_reg_53_), .Y(core__abc_22172_new_n2173_));
AND2X2 AND2X2_1839 ( .A(core__abc_22172_new_n2174_), .B(core__abc_22172_new_n2175_), .Y(core__abc_22172_new_n2176_));
AND2X2 AND2X2_184 ( .A(_abc_19873_new_n888_), .B(core_mi_12_), .Y(_abc_19873_new_n1190_));
AND2X2 AND2X2_1840 ( .A(core_v2_reg_53_), .B(core_v3_reg_53_), .Y(core__abc_22172_new_n2179_));
AND2X2 AND2X2_1841 ( .A(core__abc_22172_new_n2180_), .B(core__abc_22172_new_n2178_), .Y(core__abc_22172_new_n2181_));
AND2X2 AND2X2_1842 ( .A(core__abc_22172_new_n2177_), .B(core__abc_22172_new_n2181_), .Y(core__abc_22172_new_n2182_));
AND2X2 AND2X2_1843 ( .A(core__abc_22172_new_n2183_), .B(core__abc_22172_new_n2176_), .Y(core__abc_22172_new_n2184_));
AND2X2 AND2X2_1844 ( .A(core__abc_22172_new_n2187_), .B(reset_n), .Y(core__abc_22172_new_n2188_));
AND2X2 AND2X2_1845 ( .A(core__abc_22172_new_n2186_), .B(core__abc_22172_new_n2188_), .Y(core__0siphash_word1_reg_63_0__53_));
AND2X2 AND2X2_1846 ( .A(core_v1_reg_54_), .B(core_v0_reg_54_), .Y(core__abc_22172_new_n2191_));
AND2X2 AND2X2_1847 ( .A(core__abc_22172_new_n2192_), .B(core__abc_22172_new_n2190_), .Y(core__abc_22172_new_n2193_));
AND2X2 AND2X2_1848 ( .A(core_v2_reg_54_), .B(core_v3_reg_54_), .Y(core__abc_22172_new_n2195_));
AND2X2 AND2X2_1849 ( .A(core__abc_22172_new_n2196_), .B(core__abc_22172_new_n2194_), .Y(core__abc_22172_new_n2197_));
AND2X2 AND2X2_185 ( .A(_abc_19873_new_n916_), .B(core_key_76_), .Y(_abc_19873_new_n1193_));
AND2X2 AND2X2_1850 ( .A(core__abc_22172_new_n2201_), .B(core__abc_22172_new_n2198_), .Y(core__abc_22172_new_n2202_));
AND2X2 AND2X2_1851 ( .A(core__abc_22172_new_n2204_), .B(reset_n), .Y(core__abc_22172_new_n2205_));
AND2X2 AND2X2_1852 ( .A(core__abc_22172_new_n2203_), .B(core__abc_22172_new_n2205_), .Y(core__0siphash_word1_reg_63_0__54_));
AND2X2 AND2X2_1853 ( .A(core_v1_reg_55_), .B(core_v0_reg_55_), .Y(core__abc_22172_new_n2208_));
AND2X2 AND2X2_1854 ( .A(core__abc_22172_new_n2209_), .B(core__abc_22172_new_n2207_), .Y(core__abc_22172_new_n2210_));
AND2X2 AND2X2_1855 ( .A(core_v2_reg_55_), .B(core_v3_reg_55_), .Y(core__abc_22172_new_n2212_));
AND2X2 AND2X2_1856 ( .A(core__abc_22172_new_n2213_), .B(core__abc_22172_new_n2211_), .Y(core__abc_22172_new_n2214_));
AND2X2 AND2X2_1857 ( .A(core__abc_22172_new_n2218_), .B(core__abc_22172_new_n2215_), .Y(core__abc_22172_new_n2219_));
AND2X2 AND2X2_1858 ( .A(core__abc_22172_new_n2221_), .B(reset_n), .Y(core__abc_22172_new_n2222_));
AND2X2 AND2X2_1859 ( .A(core__abc_22172_new_n2220_), .B(core__abc_22172_new_n2222_), .Y(core__0siphash_word1_reg_63_0__55_));
AND2X2 AND2X2_186 ( .A(_abc_19873_new_n925_), .B(word2_reg_12_), .Y(_abc_19873_new_n1196_));
AND2X2 AND2X2_1860 ( .A(core_v1_reg_56_), .B(core_v0_reg_56_), .Y(core__abc_22172_new_n2225_));
AND2X2 AND2X2_1861 ( .A(core__abc_22172_new_n2226_), .B(core__abc_22172_new_n2224_), .Y(core__abc_22172_new_n2227_));
AND2X2 AND2X2_1862 ( .A(core_v2_reg_56_), .B(core_v3_reg_56_), .Y(core__abc_22172_new_n2229_));
AND2X2 AND2X2_1863 ( .A(core__abc_22172_new_n2230_), .B(core__abc_22172_new_n2228_), .Y(core__abc_22172_new_n2231_));
AND2X2 AND2X2_1864 ( .A(core__abc_22172_new_n2235_), .B(core__abc_22172_new_n2232_), .Y(core__abc_22172_new_n2236_));
AND2X2 AND2X2_1865 ( .A(core__abc_22172_new_n2238_), .B(reset_n), .Y(core__abc_22172_new_n2239_));
AND2X2 AND2X2_1866 ( .A(core__abc_22172_new_n2237_), .B(core__abc_22172_new_n2239_), .Y(core__0siphash_word1_reg_63_0__56_));
AND2X2 AND2X2_1867 ( .A(core_v1_reg_57_), .B(core_v0_reg_57_), .Y(core__abc_22172_new_n2242_));
AND2X2 AND2X2_1868 ( .A(core__abc_22172_new_n2243_), .B(core__abc_22172_new_n2241_), .Y(core__abc_22172_new_n2244_));
AND2X2 AND2X2_1869 ( .A(core_v2_reg_57_), .B(core_v3_reg_57_), .Y(core__abc_22172_new_n2246_));
AND2X2 AND2X2_187 ( .A(_abc_19873_new_n907_), .B(word1_reg_12_), .Y(_abc_19873_new_n1197_));
AND2X2 AND2X2_1870 ( .A(core__abc_22172_new_n2247_), .B(core__abc_22172_new_n2245_), .Y(core__abc_22172_new_n2248_));
AND2X2 AND2X2_1871 ( .A(core__abc_22172_new_n2252_), .B(core__abc_22172_new_n2249_), .Y(core__abc_22172_new_n2253_));
AND2X2 AND2X2_1872 ( .A(core__abc_22172_new_n2255_), .B(reset_n), .Y(core__abc_22172_new_n2256_));
AND2X2 AND2X2_1873 ( .A(core__abc_22172_new_n2254_), .B(core__abc_22172_new_n2256_), .Y(core__0siphash_word1_reg_63_0__57_));
AND2X2 AND2X2_1874 ( .A(core_v1_reg_58_), .B(core_v0_reg_58_), .Y(core__abc_22172_new_n2259_));
AND2X2 AND2X2_1875 ( .A(core__abc_22172_new_n2260_), .B(core__abc_22172_new_n2258_), .Y(core__abc_22172_new_n2261_));
AND2X2 AND2X2_1876 ( .A(core_v2_reg_58_), .B(core_v3_reg_58_), .Y(core__abc_22172_new_n2263_));
AND2X2 AND2X2_1877 ( .A(core__abc_22172_new_n2264_), .B(core__abc_22172_new_n2262_), .Y(core__abc_22172_new_n2265_));
AND2X2 AND2X2_1878 ( .A(core__abc_22172_new_n2269_), .B(core__abc_22172_new_n2266_), .Y(core__abc_22172_new_n2270_));
AND2X2 AND2X2_1879 ( .A(core__abc_22172_new_n2272_), .B(reset_n), .Y(core__abc_22172_new_n2273_));
AND2X2 AND2X2_188 ( .A(_abc_19873_new_n912_), .B(word3_reg_12_), .Y(_abc_19873_new_n1198_));
AND2X2 AND2X2_1880 ( .A(core__abc_22172_new_n2271_), .B(core__abc_22172_new_n2273_), .Y(core__0siphash_word1_reg_63_0__58_));
AND2X2 AND2X2_1881 ( .A(core_v1_reg_59_), .B(core_v0_reg_59_), .Y(core__abc_22172_new_n2276_));
AND2X2 AND2X2_1882 ( .A(core__abc_22172_new_n2277_), .B(core__abc_22172_new_n2275_), .Y(core__abc_22172_new_n2278_));
AND2X2 AND2X2_1883 ( .A(core_v2_reg_59_), .B(core_v3_reg_59_), .Y(core__abc_22172_new_n2280_));
AND2X2 AND2X2_1884 ( .A(core__abc_22172_new_n2281_), .B(core__abc_22172_new_n2279_), .Y(core__abc_22172_new_n2282_));
AND2X2 AND2X2_1885 ( .A(core__abc_22172_new_n2286_), .B(core__abc_22172_new_n2283_), .Y(core__abc_22172_new_n2287_));
AND2X2 AND2X2_1886 ( .A(core__abc_22172_new_n2289_), .B(reset_n), .Y(core__abc_22172_new_n2290_));
AND2X2 AND2X2_1887 ( .A(core__abc_22172_new_n2288_), .B(core__abc_22172_new_n2290_), .Y(core__0siphash_word1_reg_63_0__59_));
AND2X2 AND2X2_1888 ( .A(core_v1_reg_60_), .B(core_v0_reg_60_), .Y(core__abc_22172_new_n2293_));
AND2X2 AND2X2_1889 ( .A(core__abc_22172_new_n2294_), .B(core__abc_22172_new_n2292_), .Y(core__abc_22172_new_n2295_));
AND2X2 AND2X2_189 ( .A(_abc_19873_new_n928_), .B(core_key_44_), .Y(_abc_19873_new_n1201_));
AND2X2 AND2X2_1890 ( .A(core_v2_reg_60_), .B(core_v3_reg_60_), .Y(core__abc_22172_new_n2297_));
AND2X2 AND2X2_1891 ( .A(core__abc_22172_new_n2298_), .B(core__abc_22172_new_n2296_), .Y(core__abc_22172_new_n2299_));
AND2X2 AND2X2_1892 ( .A(core__abc_22172_new_n2303_), .B(core__abc_22172_new_n2300_), .Y(core__abc_22172_new_n2304_));
AND2X2 AND2X2_1893 ( .A(core__abc_22172_new_n2306_), .B(reset_n), .Y(core__abc_22172_new_n2307_));
AND2X2 AND2X2_1894 ( .A(core__abc_22172_new_n2305_), .B(core__abc_22172_new_n2307_), .Y(core__0siphash_word1_reg_63_0__60_));
AND2X2 AND2X2_1895 ( .A(core_v1_reg_61_), .B(core_v0_reg_61_), .Y(core__abc_22172_new_n2310_));
AND2X2 AND2X2_1896 ( .A(core__abc_22172_new_n2311_), .B(core__abc_22172_new_n2309_), .Y(core__abc_22172_new_n2312_));
AND2X2 AND2X2_1897 ( .A(core_v2_reg_61_), .B(core_v3_reg_61_), .Y(core__abc_22172_new_n2314_));
AND2X2 AND2X2_1898 ( .A(core__abc_22172_new_n2315_), .B(core__abc_22172_new_n2313_), .Y(core__abc_22172_new_n2316_));
AND2X2 AND2X2_1899 ( .A(core__abc_22172_new_n2320_), .B(core__abc_22172_new_n2317_), .Y(core__abc_22172_new_n2321_));
AND2X2 AND2X2_19 ( .A(_abc_19873_new_n893_), .B(_abc_19873_new_n896_), .Y(_abc_19873_new_n897_));
AND2X2 AND2X2_190 ( .A(_abc_19873_new_n901_), .B(core_key_12_), .Y(_abc_19873_new_n1202_));
AND2X2 AND2X2_1900 ( .A(core__abc_22172_new_n2323_), .B(reset_n), .Y(core__abc_22172_new_n2324_));
AND2X2 AND2X2_1901 ( .A(core__abc_22172_new_n2322_), .B(core__abc_22172_new_n2324_), .Y(core__0siphash_word1_reg_63_0__61_));
AND2X2 AND2X2_1902 ( .A(core_v1_reg_62_), .B(core_v0_reg_62_), .Y(core__abc_22172_new_n2327_));
AND2X2 AND2X2_1903 ( .A(core__abc_22172_new_n2328_), .B(core__abc_22172_new_n2326_), .Y(core__abc_22172_new_n2329_));
AND2X2 AND2X2_1904 ( .A(core_v2_reg_62_), .B(core_v3_reg_62_), .Y(core__abc_22172_new_n2331_));
AND2X2 AND2X2_1905 ( .A(core__abc_22172_new_n2332_), .B(core__abc_22172_new_n2330_), .Y(core__abc_22172_new_n2333_));
AND2X2 AND2X2_1906 ( .A(core__abc_22172_new_n2337_), .B(core__abc_22172_new_n2334_), .Y(core__abc_22172_new_n2338_));
AND2X2 AND2X2_1907 ( .A(core__abc_22172_new_n2340_), .B(reset_n), .Y(core__abc_22172_new_n2341_));
AND2X2 AND2X2_1908 ( .A(core__abc_22172_new_n2339_), .B(core__abc_22172_new_n2341_), .Y(core__0siphash_word1_reg_63_0__62_));
AND2X2 AND2X2_1909 ( .A(core__abc_22172_new_n2344_), .B(core__abc_22172_new_n2346_), .Y(core__abc_22172_new_n2347_));
AND2X2 AND2X2_191 ( .A(_abc_19873_new_n919_), .B(core_mi_44_), .Y(_abc_19873_new_n1204_));
AND2X2 AND2X2_1910 ( .A(core_v2_reg_63_), .B(core_v3_reg_63_), .Y(core__abc_22172_new_n2350_));
AND2X2 AND2X2_1911 ( .A(core__abc_22172_new_n2351_), .B(core__abc_22172_new_n2349_), .Y(core__abc_22172_new_n2352_));
AND2X2 AND2X2_1912 ( .A(core__abc_22172_new_n2353_), .B(core__abc_22172_new_n2355_), .Y(core__abc_22172_new_n2356_));
AND2X2 AND2X2_1913 ( .A(core__abc_22172_new_n2358_), .B(reset_n), .Y(core__abc_22172_new_n2359_));
AND2X2 AND2X2_1914 ( .A(core__abc_22172_new_n2357_), .B(core__abc_22172_new_n2359_), .Y(core__0siphash_word1_reg_63_0__63_));
AND2X2 AND2X2_1915 ( .A(core__abc_22172_new_n1256_), .B(core__abc_22172_new_n1169_), .Y(core__abc_22172_new_n2362_));
AND2X2 AND2X2_1916 ( .A(core__abc_22172_new_n2362_), .B(core__abc_22172_new_n2361_), .Y(core__abc_22172_new_n2363_));
AND2X2 AND2X2_1917 ( .A(core__abc_22172_new_n1218_), .B(core__abc_22172_new_n2363_), .Y(core__abc_22172_new_n2364_));
AND2X2 AND2X2_1918 ( .A(core__abc_22172_new_n2367_), .B(core__abc_22172_new_n2365_), .Y(core__abc_22172_new_n2368_));
AND2X2 AND2X2_1919 ( .A(core__abc_22172_new_n2368_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__0_));
AND2X2 AND2X2_192 ( .A(_abc_19873_new_n930_), .B(word0_reg_12_), .Y(_abc_19873_new_n1205_));
AND2X2 AND2X2_1920 ( .A(core__abc_22172_new_n2371_), .B(core__abc_22172_new_n2370_), .Y(core__abc_22172_new_n2372_));
AND2X2 AND2X2_1921 ( .A(core__abc_22172_new_n2372_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__1_));
AND2X2 AND2X2_1922 ( .A(core__abc_22172_new_n2375_), .B(core__abc_22172_new_n2374_), .Y(core__abc_22172_new_n2376_));
AND2X2 AND2X2_1923 ( .A(core__abc_22172_new_n2376_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__2_));
AND2X2 AND2X2_1924 ( .A(core__abc_22172_new_n2379_), .B(core__abc_22172_new_n2378_), .Y(core__abc_22172_new_n2380_));
AND2X2 AND2X2_1925 ( .A(core__abc_22172_new_n2380_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__3_));
AND2X2 AND2X2_1926 ( .A(core__abc_22172_new_n2383_), .B(core__abc_22172_new_n2382_), .Y(core__abc_22172_new_n2384_));
AND2X2 AND2X2_1927 ( .A(core__abc_22172_new_n2384_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__4_));
AND2X2 AND2X2_1928 ( .A(core__abc_22172_new_n2387_), .B(core__abc_22172_new_n2386_), .Y(core__abc_22172_new_n2388_));
AND2X2 AND2X2_1929 ( .A(core__abc_22172_new_n2388_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__5_));
AND2X2 AND2X2_193 ( .A(_abc_19873_new_n1209_), .B(_abc_19873_new_n937_), .Y(\read_data[12] ));
AND2X2 AND2X2_1930 ( .A(core__abc_22172_new_n2391_), .B(core__abc_22172_new_n2390_), .Y(core__abc_22172_new_n2392_));
AND2X2 AND2X2_1931 ( .A(core__abc_22172_new_n2392_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__6_));
AND2X2 AND2X2_1932 ( .A(core__abc_22172_new_n2395_), .B(core__abc_22172_new_n2394_), .Y(core__abc_22172_new_n2396_));
AND2X2 AND2X2_1933 ( .A(core__abc_22172_new_n2396_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__7_));
AND2X2 AND2X2_1934 ( .A(core__abc_22172_new_n2399_), .B(core__abc_22172_new_n2398_), .Y(core__abc_22172_new_n2400_));
AND2X2 AND2X2_1935 ( .A(core__abc_22172_new_n2400_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__8_));
AND2X2 AND2X2_1936 ( .A(core__abc_22172_new_n2403_), .B(core__abc_22172_new_n2402_), .Y(core__abc_22172_new_n2404_));
AND2X2 AND2X2_1937 ( .A(core__abc_22172_new_n2404_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__9_));
AND2X2 AND2X2_1938 ( .A(core__abc_22172_new_n2407_), .B(core__abc_22172_new_n2406_), .Y(core__abc_22172_new_n2408_));
AND2X2 AND2X2_1939 ( .A(core__abc_22172_new_n2408_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__10_));
AND2X2 AND2X2_194 ( .A(_abc_19873_new_n925_), .B(word2_reg_13_), .Y(_abc_19873_new_n1211_));
AND2X2 AND2X2_1940 ( .A(core__abc_22172_new_n2411_), .B(core__abc_22172_new_n2410_), .Y(core__abc_22172_new_n2412_));
AND2X2 AND2X2_1941 ( .A(core__abc_22172_new_n2412_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__11_));
AND2X2 AND2X2_1942 ( .A(core__abc_22172_new_n2415_), .B(core__abc_22172_new_n2414_), .Y(core__abc_22172_new_n2416_));
AND2X2 AND2X2_1943 ( .A(core__abc_22172_new_n2416_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__12_));
AND2X2 AND2X2_1944 ( .A(core__abc_22172_new_n2419_), .B(core__abc_22172_new_n2418_), .Y(core__abc_22172_new_n2420_));
AND2X2 AND2X2_1945 ( .A(core__abc_22172_new_n2420_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__13_));
AND2X2 AND2X2_1946 ( .A(core__abc_22172_new_n2423_), .B(core__abc_22172_new_n2422_), .Y(core__abc_22172_new_n2424_));
AND2X2 AND2X2_1947 ( .A(core__abc_22172_new_n2424_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__14_));
AND2X2 AND2X2_1948 ( .A(core__abc_22172_new_n2427_), .B(core__abc_22172_new_n2426_), .Y(core__abc_22172_new_n2428_));
AND2X2 AND2X2_1949 ( .A(core__abc_22172_new_n2428_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__15_));
AND2X2 AND2X2_195 ( .A(_abc_19873_new_n928_), .B(core_key_45_), .Y(_abc_19873_new_n1212_));
AND2X2 AND2X2_1950 ( .A(core__abc_22172_new_n2431_), .B(core__abc_22172_new_n2430_), .Y(core__abc_22172_new_n2432_));
AND2X2 AND2X2_1951 ( .A(core__abc_22172_new_n2432_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__16_));
AND2X2 AND2X2_1952 ( .A(core__abc_22172_new_n2435_), .B(core__abc_22172_new_n2434_), .Y(core__abc_22172_new_n2436_));
AND2X2 AND2X2_1953 ( .A(core__abc_22172_new_n2436_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__17_));
AND2X2 AND2X2_1954 ( .A(core__abc_22172_new_n2439_), .B(core__abc_22172_new_n2438_), .Y(core__abc_22172_new_n2440_));
AND2X2 AND2X2_1955 ( .A(core__abc_22172_new_n2440_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__18_));
AND2X2 AND2X2_1956 ( .A(core__abc_22172_new_n2443_), .B(core__abc_22172_new_n2442_), .Y(core__abc_22172_new_n2444_));
AND2X2 AND2X2_1957 ( .A(core__abc_22172_new_n2444_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__19_));
AND2X2 AND2X2_1958 ( .A(core__abc_22172_new_n2447_), .B(core__abc_22172_new_n2446_), .Y(core__abc_22172_new_n2448_));
AND2X2 AND2X2_1959 ( .A(core__abc_22172_new_n2448_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__20_));
AND2X2 AND2X2_196 ( .A(_abc_19873_new_n901_), .B(core_key_13_), .Y(_abc_19873_new_n1213_));
AND2X2 AND2X2_1960 ( .A(core__abc_22172_new_n2451_), .B(core__abc_22172_new_n2450_), .Y(core__abc_22172_new_n2452_));
AND2X2 AND2X2_1961 ( .A(core__abc_22172_new_n2452_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__21_));
AND2X2 AND2X2_1962 ( .A(core__abc_22172_new_n2455_), .B(core__abc_22172_new_n2454_), .Y(core__abc_22172_new_n2456_));
AND2X2 AND2X2_1963 ( .A(core__abc_22172_new_n2456_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__22_));
AND2X2 AND2X2_1964 ( .A(core__abc_22172_new_n2459_), .B(core__abc_22172_new_n2458_), .Y(core__abc_22172_new_n2460_));
AND2X2 AND2X2_1965 ( .A(core__abc_22172_new_n2460_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__23_));
AND2X2 AND2X2_1966 ( .A(core__abc_22172_new_n2463_), .B(core__abc_22172_new_n2462_), .Y(core__abc_22172_new_n2464_));
AND2X2 AND2X2_1967 ( .A(core__abc_22172_new_n2464_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__24_));
AND2X2 AND2X2_1968 ( .A(core__abc_22172_new_n2467_), .B(core__abc_22172_new_n2466_), .Y(core__abc_22172_new_n2468_));
AND2X2 AND2X2_1969 ( .A(core__abc_22172_new_n2468_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__25_));
AND2X2 AND2X2_197 ( .A(_abc_19873_new_n881_), .B(core_key_109_), .Y(_abc_19873_new_n1215_));
AND2X2 AND2X2_1970 ( .A(core__abc_22172_new_n2471_), .B(core__abc_22172_new_n2470_), .Y(core__abc_22172_new_n2472_));
AND2X2 AND2X2_1971 ( .A(core__abc_22172_new_n2472_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__26_));
AND2X2 AND2X2_1972 ( .A(core__abc_22172_new_n2475_), .B(core__abc_22172_new_n2474_), .Y(core__abc_22172_new_n2476_));
AND2X2 AND2X2_1973 ( .A(core__abc_22172_new_n2476_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__27_));
AND2X2 AND2X2_1974 ( .A(core__abc_22172_new_n2479_), .B(core__abc_22172_new_n2478_), .Y(core__abc_22172_new_n2480_));
AND2X2 AND2X2_1975 ( .A(core__abc_22172_new_n2480_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__28_));
AND2X2 AND2X2_1976 ( .A(core__abc_22172_new_n2483_), .B(core__abc_22172_new_n2482_), .Y(core__abc_22172_new_n2484_));
AND2X2 AND2X2_1977 ( .A(core__abc_22172_new_n2484_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__29_));
AND2X2 AND2X2_1978 ( .A(core__abc_22172_new_n2487_), .B(core__abc_22172_new_n2486_), .Y(core__abc_22172_new_n2488_));
AND2X2 AND2X2_1979 ( .A(core__abc_22172_new_n2488_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__30_));
AND2X2 AND2X2_198 ( .A(_abc_19873_new_n916_), .B(core_key_77_), .Y(_abc_19873_new_n1216_));
AND2X2 AND2X2_1980 ( .A(core__abc_22172_new_n2491_), .B(core__abc_22172_new_n2490_), .Y(core__abc_22172_new_n2492_));
AND2X2 AND2X2_1981 ( .A(core__abc_22172_new_n2492_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__31_));
AND2X2 AND2X2_1982 ( .A(core__abc_22172_new_n2495_), .B(core__abc_22172_new_n2494_), .Y(core__abc_22172_new_n2496_));
AND2X2 AND2X2_1983 ( .A(core__abc_22172_new_n2496_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__32_));
AND2X2 AND2X2_1984 ( .A(core__abc_22172_new_n2499_), .B(core__abc_22172_new_n2498_), .Y(core__abc_22172_new_n2500_));
AND2X2 AND2X2_1985 ( .A(core__abc_22172_new_n2500_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__33_));
AND2X2 AND2X2_1986 ( .A(core__abc_22172_new_n2503_), .B(core__abc_22172_new_n2502_), .Y(core__abc_22172_new_n2504_));
AND2X2 AND2X2_1987 ( .A(core__abc_22172_new_n2504_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__34_));
AND2X2 AND2X2_1988 ( .A(core__abc_22172_new_n2507_), .B(core__abc_22172_new_n2506_), .Y(core__abc_22172_new_n2508_));
AND2X2 AND2X2_1989 ( .A(core__abc_22172_new_n2508_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__35_));
AND2X2 AND2X2_199 ( .A(_abc_19873_new_n930_), .B(word0_reg_13_), .Y(_abc_19873_new_n1220_));
AND2X2 AND2X2_1990 ( .A(core__abc_22172_new_n2511_), .B(core__abc_22172_new_n2510_), .Y(core__abc_22172_new_n2512_));
AND2X2 AND2X2_1991 ( .A(core__abc_22172_new_n2512_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__36_));
AND2X2 AND2X2_1992 ( .A(core__abc_22172_new_n2515_), .B(core__abc_22172_new_n2514_), .Y(core__abc_22172_new_n2516_));
AND2X2 AND2X2_1993 ( .A(core__abc_22172_new_n2516_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__37_));
AND2X2 AND2X2_1994 ( .A(core__abc_22172_new_n2519_), .B(core__abc_22172_new_n2518_), .Y(core__abc_22172_new_n2520_));
AND2X2 AND2X2_1995 ( .A(core__abc_22172_new_n2520_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__38_));
AND2X2 AND2X2_1996 ( .A(core__abc_22172_new_n2523_), .B(core__abc_22172_new_n2522_), .Y(core__abc_22172_new_n2524_));
AND2X2 AND2X2_1997 ( .A(core__abc_22172_new_n2524_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__39_));
AND2X2 AND2X2_1998 ( .A(core__abc_22172_new_n2527_), .B(core__abc_22172_new_n2526_), .Y(core__abc_22172_new_n2528_));
AND2X2 AND2X2_1999 ( .A(core__abc_22172_new_n2528_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__40_));
AND2X2 AND2X2_2 ( .A(_abc_19873_new_n873_), .B(\addr[4] ), .Y(_abc_19873_new_n874_));
AND2X2 AND2X2_20 ( .A(_abc_19873_new_n897_), .B(core_compression_rounds_0_), .Y(_abc_19873_new_n898_));
AND2X2 AND2X2_200 ( .A(_abc_19873_new_n907_), .B(word1_reg_13_), .Y(_abc_19873_new_n1221_));
AND2X2 AND2X2_2000 ( .A(core__abc_22172_new_n2531_), .B(core__abc_22172_new_n2530_), .Y(core__abc_22172_new_n2532_));
AND2X2 AND2X2_2001 ( .A(core__abc_22172_new_n2532_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__41_));
AND2X2 AND2X2_2002 ( .A(core__abc_22172_new_n2535_), .B(core__abc_22172_new_n2534_), .Y(core__abc_22172_new_n2536_));
AND2X2 AND2X2_2003 ( .A(core__abc_22172_new_n2536_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__42_));
AND2X2 AND2X2_2004 ( .A(core__abc_22172_new_n2539_), .B(core__abc_22172_new_n2538_), .Y(core__abc_22172_new_n2540_));
AND2X2 AND2X2_2005 ( .A(core__abc_22172_new_n2540_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__43_));
AND2X2 AND2X2_2006 ( .A(core__abc_22172_new_n2543_), .B(core__abc_22172_new_n2542_), .Y(core__abc_22172_new_n2544_));
AND2X2 AND2X2_2007 ( .A(core__abc_22172_new_n2544_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__44_));
AND2X2 AND2X2_2008 ( .A(core__abc_22172_new_n2547_), .B(core__abc_22172_new_n2546_), .Y(core__abc_22172_new_n2548_));
AND2X2 AND2X2_2009 ( .A(core__abc_22172_new_n2548_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__45_));
AND2X2 AND2X2_201 ( .A(_abc_19873_new_n912_), .B(word3_reg_13_), .Y(_abc_19873_new_n1223_));
AND2X2 AND2X2_2010 ( .A(core__abc_22172_new_n2551_), .B(core__abc_22172_new_n2550_), .Y(core__abc_22172_new_n2552_));
AND2X2 AND2X2_2011 ( .A(core__abc_22172_new_n2552_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__46_));
AND2X2 AND2X2_2012 ( .A(core__abc_22172_new_n2555_), .B(core__abc_22172_new_n2554_), .Y(core__abc_22172_new_n2556_));
AND2X2 AND2X2_2013 ( .A(core__abc_22172_new_n2556_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__47_));
AND2X2 AND2X2_2014 ( .A(core__abc_22172_new_n2559_), .B(core__abc_22172_new_n2558_), .Y(core__abc_22172_new_n2560_));
AND2X2 AND2X2_2015 ( .A(core__abc_22172_new_n2560_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__48_));
AND2X2 AND2X2_2016 ( .A(core__abc_22172_new_n2563_), .B(core__abc_22172_new_n2562_), .Y(core__abc_22172_new_n2564_));
AND2X2 AND2X2_2017 ( .A(core__abc_22172_new_n2564_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__49_));
AND2X2 AND2X2_2018 ( .A(core__abc_22172_new_n2567_), .B(core__abc_22172_new_n2566_), .Y(core__abc_22172_new_n2568_));
AND2X2 AND2X2_2019 ( .A(core__abc_22172_new_n2568_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__50_));
AND2X2 AND2X2_202 ( .A(_abc_19873_new_n888_), .B(core_mi_13_), .Y(_abc_19873_new_n1225_));
AND2X2 AND2X2_2020 ( .A(core__abc_22172_new_n2571_), .B(core__abc_22172_new_n2570_), .Y(core__abc_22172_new_n2572_));
AND2X2 AND2X2_2021 ( .A(core__abc_22172_new_n2572_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__51_));
AND2X2 AND2X2_2022 ( .A(core__abc_22172_new_n2575_), .B(core__abc_22172_new_n2574_), .Y(core__abc_22172_new_n2576_));
AND2X2 AND2X2_2023 ( .A(core__abc_22172_new_n2576_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__52_));
AND2X2 AND2X2_2024 ( .A(core__abc_22172_new_n2579_), .B(core__abc_22172_new_n2578_), .Y(core__abc_22172_new_n2580_));
AND2X2 AND2X2_2025 ( .A(core__abc_22172_new_n2580_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__53_));
AND2X2 AND2X2_2026 ( .A(core__abc_22172_new_n2583_), .B(core__abc_22172_new_n2582_), .Y(core__abc_22172_new_n2584_));
AND2X2 AND2X2_2027 ( .A(core__abc_22172_new_n2584_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__54_));
AND2X2 AND2X2_2028 ( .A(core__abc_22172_new_n2587_), .B(core__abc_22172_new_n2586_), .Y(core__abc_22172_new_n2588_));
AND2X2 AND2X2_2029 ( .A(core__abc_22172_new_n2588_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__55_));
AND2X2 AND2X2_203 ( .A(_abc_19873_new_n919_), .B(core_mi_45_), .Y(_abc_19873_new_n1226_));
AND2X2 AND2X2_2030 ( .A(core__abc_22172_new_n2591_), .B(core__abc_22172_new_n2590_), .Y(core__abc_22172_new_n2592_));
AND2X2 AND2X2_2031 ( .A(core__abc_22172_new_n2592_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__56_));
AND2X2 AND2X2_2032 ( .A(core__abc_22172_new_n2595_), .B(core__abc_22172_new_n2594_), .Y(core__abc_22172_new_n2596_));
AND2X2 AND2X2_2033 ( .A(core__abc_22172_new_n2596_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__57_));
AND2X2 AND2X2_2034 ( .A(core__abc_22172_new_n2599_), .B(core__abc_22172_new_n2598_), .Y(core__abc_22172_new_n2600_));
AND2X2 AND2X2_2035 ( .A(core__abc_22172_new_n2600_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__58_));
AND2X2 AND2X2_2036 ( .A(core__abc_22172_new_n2603_), .B(core__abc_22172_new_n2602_), .Y(core__abc_22172_new_n2604_));
AND2X2 AND2X2_2037 ( .A(core__abc_22172_new_n2604_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__59_));
AND2X2 AND2X2_2038 ( .A(core__abc_22172_new_n2607_), .B(core__abc_22172_new_n2606_), .Y(core__abc_22172_new_n2608_));
AND2X2 AND2X2_2039 ( .A(core__abc_22172_new_n2608_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__60_));
AND2X2 AND2X2_204 ( .A(_abc_19873_new_n1230_), .B(_abc_19873_new_n937_), .Y(\read_data[13] ));
AND2X2 AND2X2_2040 ( .A(core__abc_22172_new_n2611_), .B(core__abc_22172_new_n2610_), .Y(core__abc_22172_new_n2612_));
AND2X2 AND2X2_2041 ( .A(core__abc_22172_new_n2612_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__61_));
AND2X2 AND2X2_2042 ( .A(core__abc_22172_new_n2615_), .B(core__abc_22172_new_n2614_), .Y(core__abc_22172_new_n2616_));
AND2X2 AND2X2_2043 ( .A(core__abc_22172_new_n2616_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__62_));
AND2X2 AND2X2_2044 ( .A(core__abc_22172_new_n2619_), .B(core__abc_22172_new_n2618_), .Y(core__abc_22172_new_n2620_));
AND2X2 AND2X2_2045 ( .A(core__abc_22172_new_n2620_), .B(reset_n), .Y(core__0siphash_word0_reg_63_0__63_));
AND2X2 AND2X2_2046 ( .A(core__abc_22172_new_n1218_), .B(core__abc_22172_new_n1168_), .Y(core__abc_22172_new_n2623_));
AND2X2 AND2X2_2047 ( .A(core__abc_22172_new_n2625_), .B(core_ready), .Y(core__abc_22172_new_n2626_));
AND2X2 AND2X2_2048 ( .A(core__abc_22172_new_n1173_), .B(core__abc_22172_new_n2361_), .Y(core__abc_22172_new_n2628_));
AND2X2 AND2X2_2049 ( .A(core__abc_22172_new_n2630_), .B(core__abc_22172_new_n1168_), .Y(core__abc_22172_new_n2631_));
AND2X2 AND2X2_205 ( .A(_abc_19873_new_n881_), .B(core_key_110_), .Y(_abc_19873_new_n1232_));
AND2X2 AND2X2_2050 ( .A(core__abc_22172_new_n2631_), .B(core__abc_22172_new_n2629_), .Y(core__abc_22172_new_n2632_));
AND2X2 AND2X2_2051 ( .A(core__abc_22172_new_n2633_), .B(core_loop_ctr_reg_0_), .Y(core__abc_22172_new_n2634_));
AND2X2 AND2X2_2052 ( .A(core__abc_22172_new_n2636_), .B(reset_n), .Y(core__abc_22172_new_n2637_));
AND2X2 AND2X2_2053 ( .A(core__abc_22172_new_n2635_), .B(core__abc_22172_new_n2637_), .Y(core__0loop_ctr_reg_3_0__0_));
AND2X2 AND2X2_2054 ( .A(core_loop_ctr_reg_0_), .B(core_loop_ctr_reg_1_), .Y(core__abc_22172_new_n2640_));
AND2X2 AND2X2_2055 ( .A(core__abc_22172_new_n2628_), .B(core__abc_22172_new_n2641_), .Y(core__abc_22172_new_n2642_));
AND2X2 AND2X2_2056 ( .A(core__abc_22172_new_n2643_), .B(reset_n), .Y(core__abc_22172_new_n2644_));
AND2X2 AND2X2_2057 ( .A(core__abc_22172_new_n2639_), .B(core__abc_22172_new_n2644_), .Y(core__0loop_ctr_reg_3_0__1_));
AND2X2 AND2X2_2058 ( .A(core__abc_22172_new_n2633_), .B(core__abc_22172_new_n2640_), .Y(core__abc_22172_new_n2646_));
AND2X2 AND2X2_2059 ( .A(core__abc_22172_new_n2640_), .B(core_loop_ctr_reg_2_), .Y(core__abc_22172_new_n2648_));
AND2X2 AND2X2_206 ( .A(_abc_19873_new_n888_), .B(core_mi_14_), .Y(_abc_19873_new_n1233_));
AND2X2 AND2X2_2060 ( .A(core__abc_22172_new_n2628_), .B(core__abc_22172_new_n2649_), .Y(core__abc_22172_new_n2650_));
AND2X2 AND2X2_2061 ( .A(core__abc_22172_new_n2651_), .B(reset_n), .Y(core__abc_22172_new_n2652_));
AND2X2 AND2X2_2062 ( .A(core__abc_22172_new_n2647_), .B(core__abc_22172_new_n2652_), .Y(core__0loop_ctr_reg_3_0__2_));
AND2X2 AND2X2_2063 ( .A(core__abc_22172_new_n2628_), .B(core__abc_22172_new_n2648_), .Y(core__abc_22172_new_n2655_));
AND2X2 AND2X2_2064 ( .A(core__abc_22172_new_n2656_), .B(reset_n), .Y(core__abc_22172_new_n2657_));
AND2X2 AND2X2_2065 ( .A(core__abc_22172_new_n2654_), .B(core__abc_22172_new_n2657_), .Y(core__0loop_ctr_reg_3_0__3_));
AND2X2 AND2X2_2066 ( .A(core__abc_22172_new_n1173_), .B(core__abc_22172_new_n1218_), .Y(core__abc_22172_new_n2659_));
AND2X2 AND2X2_2067 ( .A(core__abc_22172_new_n2659_), .B(core__abc_22172_new_n1214_), .Y(core__abc_22172_new_n2660_));
AND2X2 AND2X2_2068 ( .A(core__abc_22172_new_n2663_), .B(reset_n), .Y(core__abc_22172_new_n2664_));
AND2X2 AND2X2_2069 ( .A(core__abc_22172_new_n2664_), .B(core__abc_22172_new_n2661_), .Y(core__0mi_reg_63_0__0_));
AND2X2 AND2X2_207 ( .A(_abc_19873_new_n916_), .B(core_key_78_), .Y(_abc_19873_new_n1235_));
AND2X2 AND2X2_2070 ( .A(core__abc_22172_new_n2667_), .B(reset_n), .Y(core__abc_22172_new_n2668_));
AND2X2 AND2X2_2071 ( .A(core__abc_22172_new_n2668_), .B(core__abc_22172_new_n2666_), .Y(core__0mi_reg_63_0__1_));
AND2X2 AND2X2_2072 ( .A(core__abc_22172_new_n2671_), .B(reset_n), .Y(core__abc_22172_new_n2672_));
AND2X2 AND2X2_2073 ( .A(core__abc_22172_new_n2672_), .B(core__abc_22172_new_n2670_), .Y(core__0mi_reg_63_0__2_));
AND2X2 AND2X2_2074 ( .A(core__abc_22172_new_n2675_), .B(reset_n), .Y(core__abc_22172_new_n2676_));
AND2X2 AND2X2_2075 ( .A(core__abc_22172_new_n2676_), .B(core__abc_22172_new_n2674_), .Y(core__0mi_reg_63_0__3_));
AND2X2 AND2X2_2076 ( .A(core__abc_22172_new_n2679_), .B(reset_n), .Y(core__abc_22172_new_n2680_));
AND2X2 AND2X2_2077 ( .A(core__abc_22172_new_n2680_), .B(core__abc_22172_new_n2678_), .Y(core__0mi_reg_63_0__4_));
AND2X2 AND2X2_2078 ( .A(core__abc_22172_new_n2683_), .B(reset_n), .Y(core__abc_22172_new_n2684_));
AND2X2 AND2X2_2079 ( .A(core__abc_22172_new_n2684_), .B(core__abc_22172_new_n2682_), .Y(core__0mi_reg_63_0__5_));
AND2X2 AND2X2_208 ( .A(_abc_19873_new_n925_), .B(word2_reg_14_), .Y(_abc_19873_new_n1238_));
AND2X2 AND2X2_2080 ( .A(core__abc_22172_new_n2687_), .B(reset_n), .Y(core__abc_22172_new_n2688_));
AND2X2 AND2X2_2081 ( .A(core__abc_22172_new_n2688_), .B(core__abc_22172_new_n2686_), .Y(core__0mi_reg_63_0__6_));
AND2X2 AND2X2_2082 ( .A(core__abc_22172_new_n2691_), .B(reset_n), .Y(core__abc_22172_new_n2692_));
AND2X2 AND2X2_2083 ( .A(core__abc_22172_new_n2692_), .B(core__abc_22172_new_n2690_), .Y(core__0mi_reg_63_0__7_));
AND2X2 AND2X2_2084 ( .A(core__abc_22172_new_n2695_), .B(reset_n), .Y(core__abc_22172_new_n2696_));
AND2X2 AND2X2_2085 ( .A(core__abc_22172_new_n2696_), .B(core__abc_22172_new_n2694_), .Y(core__0mi_reg_63_0__8_));
AND2X2 AND2X2_2086 ( .A(core__abc_22172_new_n2699_), .B(reset_n), .Y(core__abc_22172_new_n2700_));
AND2X2 AND2X2_2087 ( .A(core__abc_22172_new_n2700_), .B(core__abc_22172_new_n2698_), .Y(core__0mi_reg_63_0__9_));
AND2X2 AND2X2_2088 ( .A(core__abc_22172_new_n2703_), .B(reset_n), .Y(core__abc_22172_new_n2704_));
AND2X2 AND2X2_2089 ( .A(core__abc_22172_new_n2704_), .B(core__abc_22172_new_n2702_), .Y(core__0mi_reg_63_0__10_));
AND2X2 AND2X2_209 ( .A(_abc_19873_new_n907_), .B(word1_reg_14_), .Y(_abc_19873_new_n1239_));
AND2X2 AND2X2_2090 ( .A(core__abc_22172_new_n2707_), .B(reset_n), .Y(core__abc_22172_new_n2708_));
AND2X2 AND2X2_2091 ( .A(core__abc_22172_new_n2708_), .B(core__abc_22172_new_n2706_), .Y(core__0mi_reg_63_0__11_));
AND2X2 AND2X2_2092 ( .A(core__abc_22172_new_n2711_), .B(reset_n), .Y(core__abc_22172_new_n2712_));
AND2X2 AND2X2_2093 ( .A(core__abc_22172_new_n2712_), .B(core__abc_22172_new_n2710_), .Y(core__0mi_reg_63_0__12_));
AND2X2 AND2X2_2094 ( .A(core__abc_22172_new_n2715_), .B(reset_n), .Y(core__abc_22172_new_n2716_));
AND2X2 AND2X2_2095 ( .A(core__abc_22172_new_n2716_), .B(core__abc_22172_new_n2714_), .Y(core__0mi_reg_63_0__13_));
AND2X2 AND2X2_2096 ( .A(core__abc_22172_new_n2719_), .B(reset_n), .Y(core__abc_22172_new_n2720_));
AND2X2 AND2X2_2097 ( .A(core__abc_22172_new_n2720_), .B(core__abc_22172_new_n2718_), .Y(core__0mi_reg_63_0__14_));
AND2X2 AND2X2_2098 ( .A(core__abc_22172_new_n2723_), .B(reset_n), .Y(core__abc_22172_new_n2724_));
AND2X2 AND2X2_2099 ( .A(core__abc_22172_new_n2724_), .B(core__abc_22172_new_n2722_), .Y(core__0mi_reg_63_0__15_));
AND2X2 AND2X2_21 ( .A(_abc_19873_new_n879_), .B(_abc_19873_new_n885_), .Y(_abc_19873_new_n900_));
AND2X2 AND2X2_210 ( .A(_abc_19873_new_n912_), .B(word3_reg_14_), .Y(_abc_19873_new_n1240_));
AND2X2 AND2X2_2100 ( .A(core__abc_22172_new_n2727_), .B(reset_n), .Y(core__abc_22172_new_n2728_));
AND2X2 AND2X2_2101 ( .A(core__abc_22172_new_n2728_), .B(core__abc_22172_new_n2726_), .Y(core__0mi_reg_63_0__16_));
AND2X2 AND2X2_2102 ( .A(core__abc_22172_new_n2731_), .B(reset_n), .Y(core__abc_22172_new_n2732_));
AND2X2 AND2X2_2103 ( .A(core__abc_22172_new_n2732_), .B(core__abc_22172_new_n2730_), .Y(core__0mi_reg_63_0__17_));
AND2X2 AND2X2_2104 ( .A(core__abc_22172_new_n2735_), .B(reset_n), .Y(core__abc_22172_new_n2736_));
AND2X2 AND2X2_2105 ( .A(core__abc_22172_new_n2736_), .B(core__abc_22172_new_n2734_), .Y(core__0mi_reg_63_0__18_));
AND2X2 AND2X2_2106 ( .A(core__abc_22172_new_n2739_), .B(reset_n), .Y(core__abc_22172_new_n2740_));
AND2X2 AND2X2_2107 ( .A(core__abc_22172_new_n2740_), .B(core__abc_22172_new_n2738_), .Y(core__0mi_reg_63_0__19_));
AND2X2 AND2X2_2108 ( .A(core__abc_22172_new_n2743_), .B(reset_n), .Y(core__abc_22172_new_n2744_));
AND2X2 AND2X2_2109 ( .A(core__abc_22172_new_n2744_), .B(core__abc_22172_new_n2742_), .Y(core__0mi_reg_63_0__20_));
AND2X2 AND2X2_211 ( .A(_abc_19873_new_n919_), .B(core_mi_46_), .Y(_abc_19873_new_n1243_));
AND2X2 AND2X2_2110 ( .A(core__abc_22172_new_n2747_), .B(reset_n), .Y(core__abc_22172_new_n2748_));
AND2X2 AND2X2_2111 ( .A(core__abc_22172_new_n2748_), .B(core__abc_22172_new_n2746_), .Y(core__0mi_reg_63_0__21_));
AND2X2 AND2X2_2112 ( .A(core__abc_22172_new_n2751_), .B(reset_n), .Y(core__abc_22172_new_n2752_));
AND2X2 AND2X2_2113 ( .A(core__abc_22172_new_n2752_), .B(core__abc_22172_new_n2750_), .Y(core__0mi_reg_63_0__22_));
AND2X2 AND2X2_2114 ( .A(core__abc_22172_new_n2755_), .B(reset_n), .Y(core__abc_22172_new_n2756_));
AND2X2 AND2X2_2115 ( .A(core__abc_22172_new_n2756_), .B(core__abc_22172_new_n2754_), .Y(core__0mi_reg_63_0__23_));
AND2X2 AND2X2_2116 ( .A(core__abc_22172_new_n2759_), .B(reset_n), .Y(core__abc_22172_new_n2760_));
AND2X2 AND2X2_2117 ( .A(core__abc_22172_new_n2760_), .B(core__abc_22172_new_n2758_), .Y(core__0mi_reg_63_0__24_));
AND2X2 AND2X2_2118 ( .A(core__abc_22172_new_n2763_), .B(reset_n), .Y(core__abc_22172_new_n2764_));
AND2X2 AND2X2_2119 ( .A(core__abc_22172_new_n2764_), .B(core__abc_22172_new_n2762_), .Y(core__0mi_reg_63_0__25_));
AND2X2 AND2X2_212 ( .A(_abc_19873_new_n930_), .B(word0_reg_14_), .Y(_abc_19873_new_n1244_));
AND2X2 AND2X2_2120 ( .A(core__abc_22172_new_n2767_), .B(reset_n), .Y(core__abc_22172_new_n2768_));
AND2X2 AND2X2_2121 ( .A(core__abc_22172_new_n2768_), .B(core__abc_22172_new_n2766_), .Y(core__0mi_reg_63_0__26_));
AND2X2 AND2X2_2122 ( .A(core__abc_22172_new_n2771_), .B(reset_n), .Y(core__abc_22172_new_n2772_));
AND2X2 AND2X2_2123 ( .A(core__abc_22172_new_n2772_), .B(core__abc_22172_new_n2770_), .Y(core__0mi_reg_63_0__27_));
AND2X2 AND2X2_2124 ( .A(core__abc_22172_new_n2775_), .B(reset_n), .Y(core__abc_22172_new_n2776_));
AND2X2 AND2X2_2125 ( .A(core__abc_22172_new_n2776_), .B(core__abc_22172_new_n2774_), .Y(core__0mi_reg_63_0__28_));
AND2X2 AND2X2_2126 ( .A(core__abc_22172_new_n2779_), .B(reset_n), .Y(core__abc_22172_new_n2780_));
AND2X2 AND2X2_2127 ( .A(core__abc_22172_new_n2780_), .B(core__abc_22172_new_n2778_), .Y(core__0mi_reg_63_0__29_));
AND2X2 AND2X2_2128 ( .A(core__abc_22172_new_n2783_), .B(reset_n), .Y(core__abc_22172_new_n2784_));
AND2X2 AND2X2_2129 ( .A(core__abc_22172_new_n2784_), .B(core__abc_22172_new_n2782_), .Y(core__0mi_reg_63_0__30_));
AND2X2 AND2X2_213 ( .A(_abc_19873_new_n928_), .B(core_key_46_), .Y(_abc_19873_new_n1246_));
AND2X2 AND2X2_2130 ( .A(core__abc_22172_new_n2787_), .B(reset_n), .Y(core__abc_22172_new_n2788_));
AND2X2 AND2X2_2131 ( .A(core__abc_22172_new_n2788_), .B(core__abc_22172_new_n2786_), .Y(core__0mi_reg_63_0__31_));
AND2X2 AND2X2_2132 ( .A(core__abc_22172_new_n2791_), .B(reset_n), .Y(core__abc_22172_new_n2792_));
AND2X2 AND2X2_2133 ( .A(core__abc_22172_new_n2792_), .B(core__abc_22172_new_n2790_), .Y(core__0mi_reg_63_0__32_));
AND2X2 AND2X2_2134 ( .A(core__abc_22172_new_n2795_), .B(reset_n), .Y(core__abc_22172_new_n2796_));
AND2X2 AND2X2_2135 ( .A(core__abc_22172_new_n2796_), .B(core__abc_22172_new_n2794_), .Y(core__0mi_reg_63_0__33_));
AND2X2 AND2X2_2136 ( .A(core__abc_22172_new_n2799_), .B(reset_n), .Y(core__abc_22172_new_n2800_));
AND2X2 AND2X2_2137 ( .A(core__abc_22172_new_n2800_), .B(core__abc_22172_new_n2798_), .Y(core__0mi_reg_63_0__34_));
AND2X2 AND2X2_2138 ( .A(core__abc_22172_new_n2803_), .B(reset_n), .Y(core__abc_22172_new_n2804_));
AND2X2 AND2X2_2139 ( .A(core__abc_22172_new_n2804_), .B(core__abc_22172_new_n2802_), .Y(core__0mi_reg_63_0__35_));
AND2X2 AND2X2_214 ( .A(_abc_19873_new_n901_), .B(core_key_14_), .Y(_abc_19873_new_n1247_));
AND2X2 AND2X2_2140 ( .A(core__abc_22172_new_n2807_), .B(reset_n), .Y(core__abc_22172_new_n2808_));
AND2X2 AND2X2_2141 ( .A(core__abc_22172_new_n2808_), .B(core__abc_22172_new_n2806_), .Y(core__0mi_reg_63_0__36_));
AND2X2 AND2X2_2142 ( .A(core__abc_22172_new_n2811_), .B(reset_n), .Y(core__abc_22172_new_n2812_));
AND2X2 AND2X2_2143 ( .A(core__abc_22172_new_n2812_), .B(core__abc_22172_new_n2810_), .Y(core__0mi_reg_63_0__37_));
AND2X2 AND2X2_2144 ( .A(core__abc_22172_new_n2815_), .B(reset_n), .Y(core__abc_22172_new_n2816_));
AND2X2 AND2X2_2145 ( .A(core__abc_22172_new_n2816_), .B(core__abc_22172_new_n2814_), .Y(core__0mi_reg_63_0__38_));
AND2X2 AND2X2_2146 ( .A(core__abc_22172_new_n2819_), .B(reset_n), .Y(core__abc_22172_new_n2820_));
AND2X2 AND2X2_2147 ( .A(core__abc_22172_new_n2820_), .B(core__abc_22172_new_n2818_), .Y(core__0mi_reg_63_0__39_));
AND2X2 AND2X2_2148 ( .A(core__abc_22172_new_n2823_), .B(reset_n), .Y(core__abc_22172_new_n2824_));
AND2X2 AND2X2_2149 ( .A(core__abc_22172_new_n2824_), .B(core__abc_22172_new_n2822_), .Y(core__0mi_reg_63_0__40_));
AND2X2 AND2X2_215 ( .A(_abc_19873_new_n1251_), .B(_abc_19873_new_n937_), .Y(\read_data[14] ));
AND2X2 AND2X2_2150 ( .A(core__abc_22172_new_n2827_), .B(reset_n), .Y(core__abc_22172_new_n2828_));
AND2X2 AND2X2_2151 ( .A(core__abc_22172_new_n2828_), .B(core__abc_22172_new_n2826_), .Y(core__0mi_reg_63_0__41_));
AND2X2 AND2X2_2152 ( .A(core__abc_22172_new_n2831_), .B(reset_n), .Y(core__abc_22172_new_n2832_));
AND2X2 AND2X2_2153 ( .A(core__abc_22172_new_n2832_), .B(core__abc_22172_new_n2830_), .Y(core__0mi_reg_63_0__42_));
AND2X2 AND2X2_2154 ( .A(core__abc_22172_new_n2835_), .B(reset_n), .Y(core__abc_22172_new_n2836_));
AND2X2 AND2X2_2155 ( .A(core__abc_22172_new_n2836_), .B(core__abc_22172_new_n2834_), .Y(core__0mi_reg_63_0__43_));
AND2X2 AND2X2_2156 ( .A(core__abc_22172_new_n2839_), .B(reset_n), .Y(core__abc_22172_new_n2840_));
AND2X2 AND2X2_2157 ( .A(core__abc_22172_new_n2840_), .B(core__abc_22172_new_n2838_), .Y(core__0mi_reg_63_0__44_));
AND2X2 AND2X2_2158 ( .A(core__abc_22172_new_n2843_), .B(reset_n), .Y(core__abc_22172_new_n2844_));
AND2X2 AND2X2_2159 ( .A(core__abc_22172_new_n2844_), .B(core__abc_22172_new_n2842_), .Y(core__0mi_reg_63_0__45_));
AND2X2 AND2X2_216 ( .A(_abc_19873_new_n881_), .B(core_key_111_), .Y(_abc_19873_new_n1253_));
AND2X2 AND2X2_2160 ( .A(core__abc_22172_new_n2847_), .B(reset_n), .Y(core__abc_22172_new_n2848_));
AND2X2 AND2X2_2161 ( .A(core__abc_22172_new_n2848_), .B(core__abc_22172_new_n2846_), .Y(core__0mi_reg_63_0__46_));
AND2X2 AND2X2_2162 ( .A(core__abc_22172_new_n2851_), .B(reset_n), .Y(core__abc_22172_new_n2852_));
AND2X2 AND2X2_2163 ( .A(core__abc_22172_new_n2852_), .B(core__abc_22172_new_n2850_), .Y(core__0mi_reg_63_0__47_));
AND2X2 AND2X2_2164 ( .A(core__abc_22172_new_n2855_), .B(reset_n), .Y(core__abc_22172_new_n2856_));
AND2X2 AND2X2_2165 ( .A(core__abc_22172_new_n2856_), .B(core__abc_22172_new_n2854_), .Y(core__0mi_reg_63_0__48_));
AND2X2 AND2X2_2166 ( .A(core__abc_22172_new_n2859_), .B(reset_n), .Y(core__abc_22172_new_n2860_));
AND2X2 AND2X2_2167 ( .A(core__abc_22172_new_n2860_), .B(core__abc_22172_new_n2858_), .Y(core__0mi_reg_63_0__49_));
AND2X2 AND2X2_2168 ( .A(core__abc_22172_new_n2863_), .B(reset_n), .Y(core__abc_22172_new_n2864_));
AND2X2 AND2X2_2169 ( .A(core__abc_22172_new_n2864_), .B(core__abc_22172_new_n2862_), .Y(core__0mi_reg_63_0__50_));
AND2X2 AND2X2_217 ( .A(_abc_19873_new_n916_), .B(core_key_79_), .Y(_abc_19873_new_n1254_));
AND2X2 AND2X2_2170 ( .A(core__abc_22172_new_n2867_), .B(reset_n), .Y(core__abc_22172_new_n2868_));
AND2X2 AND2X2_2171 ( .A(core__abc_22172_new_n2868_), .B(core__abc_22172_new_n2866_), .Y(core__0mi_reg_63_0__51_));
AND2X2 AND2X2_2172 ( .A(core__abc_22172_new_n2871_), .B(reset_n), .Y(core__abc_22172_new_n2872_));
AND2X2 AND2X2_2173 ( .A(core__abc_22172_new_n2872_), .B(core__abc_22172_new_n2870_), .Y(core__0mi_reg_63_0__52_));
AND2X2 AND2X2_2174 ( .A(core__abc_22172_new_n2875_), .B(reset_n), .Y(core__abc_22172_new_n2876_));
AND2X2 AND2X2_2175 ( .A(core__abc_22172_new_n2876_), .B(core__abc_22172_new_n2874_), .Y(core__0mi_reg_63_0__53_));
AND2X2 AND2X2_2176 ( .A(core__abc_22172_new_n2879_), .B(reset_n), .Y(core__abc_22172_new_n2880_));
AND2X2 AND2X2_2177 ( .A(core__abc_22172_new_n2880_), .B(core__abc_22172_new_n2878_), .Y(core__0mi_reg_63_0__54_));
AND2X2 AND2X2_2178 ( .A(core__abc_22172_new_n2883_), .B(reset_n), .Y(core__abc_22172_new_n2884_));
AND2X2 AND2X2_2179 ( .A(core__abc_22172_new_n2884_), .B(core__abc_22172_new_n2882_), .Y(core__0mi_reg_63_0__55_));
AND2X2 AND2X2_218 ( .A(_abc_19873_new_n912_), .B(word3_reg_15_), .Y(_abc_19873_new_n1256_));
AND2X2 AND2X2_2180 ( .A(core__abc_22172_new_n2887_), .B(reset_n), .Y(core__abc_22172_new_n2888_));
AND2X2 AND2X2_2181 ( .A(core__abc_22172_new_n2888_), .B(core__abc_22172_new_n2886_), .Y(core__0mi_reg_63_0__56_));
AND2X2 AND2X2_2182 ( .A(core__abc_22172_new_n2891_), .B(reset_n), .Y(core__abc_22172_new_n2892_));
AND2X2 AND2X2_2183 ( .A(core__abc_22172_new_n2892_), .B(core__abc_22172_new_n2890_), .Y(core__0mi_reg_63_0__57_));
AND2X2 AND2X2_2184 ( .A(core__abc_22172_new_n2895_), .B(reset_n), .Y(core__abc_22172_new_n2896_));
AND2X2 AND2X2_2185 ( .A(core__abc_22172_new_n2896_), .B(core__abc_22172_new_n2894_), .Y(core__0mi_reg_63_0__58_));
AND2X2 AND2X2_2186 ( .A(core__abc_22172_new_n2899_), .B(reset_n), .Y(core__abc_22172_new_n2900_));
AND2X2 AND2X2_2187 ( .A(core__abc_22172_new_n2900_), .B(core__abc_22172_new_n2898_), .Y(core__0mi_reg_63_0__59_));
AND2X2 AND2X2_2188 ( .A(core__abc_22172_new_n2903_), .B(reset_n), .Y(core__abc_22172_new_n2904_));
AND2X2 AND2X2_2189 ( .A(core__abc_22172_new_n2904_), .B(core__abc_22172_new_n2902_), .Y(core__0mi_reg_63_0__60_));
AND2X2 AND2X2_219 ( .A(_abc_19873_new_n907_), .B(word1_reg_15_), .Y(_abc_19873_new_n1257_));
AND2X2 AND2X2_2190 ( .A(core__abc_22172_new_n2907_), .B(reset_n), .Y(core__abc_22172_new_n2908_));
AND2X2 AND2X2_2191 ( .A(core__abc_22172_new_n2908_), .B(core__abc_22172_new_n2906_), .Y(core__0mi_reg_63_0__61_));
AND2X2 AND2X2_2192 ( .A(core__abc_22172_new_n2911_), .B(reset_n), .Y(core__abc_22172_new_n2912_));
AND2X2 AND2X2_2193 ( .A(core__abc_22172_new_n2912_), .B(core__abc_22172_new_n2910_), .Y(core__0mi_reg_63_0__62_));
AND2X2 AND2X2_2194 ( .A(core__abc_22172_new_n2915_), .B(reset_n), .Y(core__abc_22172_new_n2916_));
AND2X2 AND2X2_2195 ( .A(core__abc_22172_new_n2916_), .B(core__abc_22172_new_n2914_), .Y(core__0mi_reg_63_0__63_));
AND2X2 AND2X2_2196 ( .A(core__abc_22172_new_n1278_), .B(core__abc_22172_new_n1258_), .Y(core__abc_22172_new_n2918_));
AND2X2 AND2X2_2197 ( .A(core__abc_22172_new_n1299_), .B(core__abc_22172_new_n1317_), .Y(core__abc_22172_new_n2920_));
AND2X2 AND2X2_2198 ( .A(core__abc_22172_new_n2919_), .B(core__abc_22172_new_n2920_), .Y(core__abc_22172_new_n2921_));
AND2X2 AND2X2_2199 ( .A(core__abc_22172_new_n1314_), .B(core__abc_22172_new_n1296_), .Y(core__abc_22172_new_n2922_));
AND2X2 AND2X2_22 ( .A(_abc_19873_new_n900_), .B(_abc_19873_new_n875_), .Y(_abc_19873_new_n901_));
AND2X2 AND2X2_220 ( .A(_abc_19873_new_n930_), .B(word0_reg_15_), .Y(_abc_19873_new_n1258_));
AND2X2 AND2X2_2200 ( .A(core__abc_22172_new_n1373_), .B(core__abc_22172_new_n1391_), .Y(core__abc_22172_new_n2925_));
AND2X2 AND2X2_2201 ( .A(core__abc_22172_new_n1335_), .B(core__abc_22172_new_n1353_), .Y(core__abc_22172_new_n2926_));
AND2X2 AND2X2_2202 ( .A(core__abc_22172_new_n2925_), .B(core__abc_22172_new_n2926_), .Y(core__abc_22172_new_n2927_));
AND2X2 AND2X2_2203 ( .A(core__abc_22172_new_n2924_), .B(core__abc_22172_new_n2927_), .Y(core__abc_22172_new_n2928_));
AND2X2 AND2X2_2204 ( .A(core__abc_22172_new_n2929_), .B(core__abc_22172_new_n1350_), .Y(core__abc_22172_new_n2930_));
AND2X2 AND2X2_2205 ( .A(core__abc_22172_new_n2925_), .B(core__abc_22172_new_n2930_), .Y(core__abc_22172_new_n2931_));
AND2X2 AND2X2_2206 ( .A(core__abc_22172_new_n1388_), .B(core__abc_22172_new_n1371_), .Y(core__abc_22172_new_n2932_));
AND2X2 AND2X2_2207 ( .A(core__abc_22172_new_n1513_), .B(core__abc_22172_new_n1530_), .Y(core__abc_22172_new_n2936_));
AND2X2 AND2X2_2208 ( .A(core__abc_22172_new_n1479_), .B(core__abc_22172_new_n1496_), .Y(core__abc_22172_new_n2937_));
AND2X2 AND2X2_2209 ( .A(core__abc_22172_new_n2936_), .B(core__abc_22172_new_n2937_), .Y(core__abc_22172_new_n2938_));
AND2X2 AND2X2_221 ( .A(_abc_19873_new_n925_), .B(word2_reg_15_), .Y(_abc_19873_new_n1262_));
AND2X2 AND2X2_2210 ( .A(core__abc_22172_new_n1411_), .B(core__abc_22172_new_n1428_), .Y(core__abc_22172_new_n2939_));
AND2X2 AND2X2_2211 ( .A(core__abc_22172_new_n1445_), .B(core__abc_22172_new_n1462_), .Y(core__abc_22172_new_n2940_));
AND2X2 AND2X2_2212 ( .A(core__abc_22172_new_n2939_), .B(core__abc_22172_new_n2940_), .Y(core__abc_22172_new_n2941_));
AND2X2 AND2X2_2213 ( .A(core__abc_22172_new_n2938_), .B(core__abc_22172_new_n2941_), .Y(core__abc_22172_new_n2942_));
AND2X2 AND2X2_2214 ( .A(core__abc_22172_new_n2935_), .B(core__abc_22172_new_n2942_), .Y(core__abc_22172_new_n2943_));
AND2X2 AND2X2_2215 ( .A(core__abc_22172_new_n2944_), .B(core__abc_22172_new_n1425_), .Y(core__abc_22172_new_n2945_));
AND2X2 AND2X2_2216 ( .A(core__abc_22172_new_n2940_), .B(core__abc_22172_new_n2945_), .Y(core__abc_22172_new_n2946_));
AND2X2 AND2X2_2217 ( .A(core__abc_22172_new_n2947_), .B(core__abc_22172_new_n1461_), .Y(core__abc_22172_new_n2948_));
AND2X2 AND2X2_2218 ( .A(core__abc_22172_new_n2950_), .B(core__abc_22172_new_n2938_), .Y(core__abc_22172_new_n2951_));
AND2X2 AND2X2_2219 ( .A(core__abc_22172_new_n2952_), .B(core__abc_22172_new_n1495_), .Y(core__abc_22172_new_n2953_));
AND2X2 AND2X2_222 ( .A(_abc_19873_new_n928_), .B(core_key_47_), .Y(_abc_19873_new_n1263_));
AND2X2 AND2X2_2220 ( .A(core__abc_22172_new_n2954_), .B(core__abc_22172_new_n2936_), .Y(core__abc_22172_new_n2955_));
AND2X2 AND2X2_2221 ( .A(core__abc_22172_new_n1527_), .B(core__abc_22172_new_n1511_), .Y(core__abc_22172_new_n2956_));
AND2X2 AND2X2_2222 ( .A(core__abc_22172_new_n1785_), .B(core__abc_22172_new_n1802_), .Y(core__abc_22172_new_n2961_));
AND2X2 AND2X2_2223 ( .A(core__abc_22172_new_n1751_), .B(core__abc_22172_new_n1768_), .Y(core__abc_22172_new_n2962_));
AND2X2 AND2X2_2224 ( .A(core__abc_22172_new_n2961_), .B(core__abc_22172_new_n2962_), .Y(core__abc_22172_new_n2963_));
AND2X2 AND2X2_2225 ( .A(core__abc_22172_new_n1683_), .B(core__abc_22172_new_n1700_), .Y(core__abc_22172_new_n2964_));
AND2X2 AND2X2_2226 ( .A(core__abc_22172_new_n1717_), .B(core__abc_22172_new_n1734_), .Y(core__abc_22172_new_n2965_));
AND2X2 AND2X2_2227 ( .A(core__abc_22172_new_n2964_), .B(core__abc_22172_new_n2965_), .Y(core__abc_22172_new_n2966_));
AND2X2 AND2X2_2228 ( .A(core__abc_22172_new_n2963_), .B(core__abc_22172_new_n2966_), .Y(core__abc_22172_new_n2967_));
AND2X2 AND2X2_2229 ( .A(core__abc_22172_new_n1649_), .B(core__abc_22172_new_n1666_), .Y(core__abc_22172_new_n2968_));
AND2X2 AND2X2_223 ( .A(_abc_19873_new_n901_), .B(core_key_15_), .Y(_abc_19873_new_n1264_));
AND2X2 AND2X2_2230 ( .A(core__abc_22172_new_n1615_), .B(core__abc_22172_new_n1632_), .Y(core__abc_22172_new_n2969_));
AND2X2 AND2X2_2231 ( .A(core__abc_22172_new_n2968_), .B(core__abc_22172_new_n2969_), .Y(core__abc_22172_new_n2970_));
AND2X2 AND2X2_2232 ( .A(core__abc_22172_new_n1547_), .B(core__abc_22172_new_n1564_), .Y(core__abc_22172_new_n2971_));
AND2X2 AND2X2_2233 ( .A(core__abc_22172_new_n1581_), .B(core__abc_22172_new_n1598_), .Y(core__abc_22172_new_n2972_));
AND2X2 AND2X2_2234 ( .A(core__abc_22172_new_n2971_), .B(core__abc_22172_new_n2972_), .Y(core__abc_22172_new_n2973_));
AND2X2 AND2X2_2235 ( .A(core__abc_22172_new_n2970_), .B(core__abc_22172_new_n2973_), .Y(core__abc_22172_new_n2974_));
AND2X2 AND2X2_2236 ( .A(core__abc_22172_new_n2967_), .B(core__abc_22172_new_n2974_), .Y(core__abc_22172_new_n2975_));
AND2X2 AND2X2_2237 ( .A(core__abc_22172_new_n2960_), .B(core__abc_22172_new_n2975_), .Y(core__abc_22172_new_n2976_));
AND2X2 AND2X2_2238 ( .A(core__abc_22172_new_n2977_), .B(core__abc_22172_new_n1561_), .Y(core__abc_22172_new_n2978_));
AND2X2 AND2X2_2239 ( .A(core__abc_22172_new_n2972_), .B(core__abc_22172_new_n2978_), .Y(core__abc_22172_new_n2979_));
AND2X2 AND2X2_224 ( .A(_abc_19873_new_n919_), .B(core_mi_47_), .Y(_abc_19873_new_n1266_));
AND2X2 AND2X2_2240 ( .A(core__abc_22172_new_n1595_), .B(core__abc_22172_new_n1579_), .Y(core__abc_22172_new_n2980_));
AND2X2 AND2X2_2241 ( .A(core__abc_22172_new_n2982_), .B(core__abc_22172_new_n2970_), .Y(core__abc_22172_new_n2983_));
AND2X2 AND2X2_2242 ( .A(core__abc_22172_new_n1614_), .B(core__abc_22172_new_n1631_), .Y(core__abc_22172_new_n2985_));
AND2X2 AND2X2_2243 ( .A(core__abc_22172_new_n2987_), .B(core__abc_22172_new_n2968_), .Y(core__abc_22172_new_n2988_));
AND2X2 AND2X2_2244 ( .A(core__abc_22172_new_n1663_), .B(core__abc_22172_new_n1647_), .Y(core__abc_22172_new_n2989_));
AND2X2 AND2X2_2245 ( .A(core__abc_22172_new_n2992_), .B(core__abc_22172_new_n2967_), .Y(core__abc_22172_new_n2993_));
AND2X2 AND2X2_2246 ( .A(core__abc_22172_new_n1682_), .B(core__abc_22172_new_n1699_), .Y(core__abc_22172_new_n2995_));
AND2X2 AND2X2_2247 ( .A(core__abc_22172_new_n2997_), .B(core__abc_22172_new_n2965_), .Y(core__abc_22172_new_n2998_));
AND2X2 AND2X2_2248 ( .A(core__abc_22172_new_n1731_), .B(core__abc_22172_new_n1715_), .Y(core__abc_22172_new_n2999_));
AND2X2 AND2X2_2249 ( .A(core__abc_22172_new_n3001_), .B(core__abc_22172_new_n2963_), .Y(core__abc_22172_new_n3002_));
AND2X2 AND2X2_225 ( .A(_abc_19873_new_n888_), .B(core_mi_15_), .Y(_abc_19873_new_n1267_));
AND2X2 AND2X2_2250 ( .A(core__abc_22172_new_n1799_), .B(core__abc_22172_new_n1783_), .Y(core__abc_22172_new_n3003_));
AND2X2 AND2X2_2251 ( .A(core__abc_22172_new_n1750_), .B(core__abc_22172_new_n1767_), .Y(core__abc_22172_new_n3006_));
AND2X2 AND2X2_2252 ( .A(core__abc_22172_new_n3008_), .B(core__abc_22172_new_n2961_), .Y(core__abc_22172_new_n3009_));
AND2X2 AND2X2_2253 ( .A(core__abc_22172_new_n3013_), .B(core__abc_22172_new_n1819_), .Y(core__abc_22172_new_n3014_));
AND2X2 AND2X2_2254 ( .A(core__abc_22172_new_n3015_), .B(core__abc_22172_new_n1277_), .Y(core__abc_22172_new_n3016_));
AND2X2 AND2X2_2255 ( .A(core__abc_22172_new_n3018_), .B(core__abc_22172_new_n3019_), .Y(core__abc_22172_new_n3020_));
AND2X2 AND2X2_2256 ( .A(core__abc_22172_new_n3022_), .B(core__abc_22172_new_n3023_), .Y(core__abc_22172_new_n3024_));
AND2X2 AND2X2_2257 ( .A(core__abc_22172_new_n3026_), .B(core__abc_22172_new_n3027_), .Y(core__abc_22172_new_n3028_));
AND2X2 AND2X2_2258 ( .A(core__abc_22172_new_n3030_), .B(core__abc_22172_new_n3031_), .Y(core__abc_22172_new_n3032_));
AND2X2 AND2X2_2259 ( .A(core__abc_22172_new_n3032_), .B(core__abc_22172_new_n1825_), .Y(core__abc_22172_new_n3033_));
AND2X2 AND2X2_226 ( .A(_abc_19873_new_n1271_), .B(_abc_19873_new_n937_), .Y(\read_data[15] ));
AND2X2 AND2X2_2260 ( .A(core__abc_22172_new_n1265_), .B(core_v3_reg_48_), .Y(core__abc_22172_new_n3035_));
AND2X2 AND2X2_2261 ( .A(core__abc_22172_new_n3036_), .B(core__abc_22172_new_n3037_), .Y(core__abc_22172_new_n3038_));
AND2X2 AND2X2_2262 ( .A(core__abc_22172_new_n3034_), .B(core__abc_22172_new_n3038_), .Y(core__abc_22172_new_n3039_));
AND2X2 AND2X2_2263 ( .A(core__abc_22172_new_n3040_), .B(core__abc_22172_new_n3041_), .Y(core__abc_22172_new_n3042_));
AND2X2 AND2X2_2264 ( .A(core__abc_22172_new_n1957_), .B(core__abc_22172_new_n1974_), .Y(core__abc_22172_new_n3046_));
AND2X2 AND2X2_2265 ( .A(core__abc_22172_new_n1323_), .B(core__abc_22172_new_n1301_), .Y(core__abc_22172_new_n3049_));
AND2X2 AND2X2_2266 ( .A(core__abc_22172_new_n3054_), .B(core__abc_22172_new_n3052_), .Y(core__abc_22172_new_n3055_));
AND2X2 AND2X2_2267 ( .A(core__abc_22172_new_n1306_), .B(core__abc_22172_new_n1323_), .Y(core__abc_22172_new_n3056_));
AND2X2 AND2X2_2268 ( .A(core__abc_22172_new_n3058_), .B(core__abc_22172_new_n3051_), .Y(core__abc_22172_new_n3059_));
AND2X2 AND2X2_2269 ( .A(core__abc_22172_new_n1379_), .B(core__abc_22172_new_n1398_), .Y(core__abc_22172_new_n3061_));
AND2X2 AND2X2_227 ( .A(_abc_19873_new_n881_), .B(core_key_112_), .Y(_abc_19873_new_n1273_));
AND2X2 AND2X2_2270 ( .A(core__abc_22172_new_n1341_), .B(core__abc_22172_new_n1360_), .Y(core__abc_22172_new_n3062_));
AND2X2 AND2X2_2271 ( .A(core__abc_22172_new_n3061_), .B(core__abc_22172_new_n3062_), .Y(core__abc_22172_new_n3063_));
AND2X2 AND2X2_2272 ( .A(core__abc_22172_new_n3060_), .B(core__abc_22172_new_n3063_), .Y(core__abc_22172_new_n3064_));
AND2X2 AND2X2_2273 ( .A(core__abc_22172_new_n3065_), .B(core__abc_22172_new_n1355_), .Y(core__abc_22172_new_n3066_));
AND2X2 AND2X2_2274 ( .A(core__abc_22172_new_n3068_), .B(core__abc_22172_new_n3061_), .Y(core__abc_22172_new_n3069_));
AND2X2 AND2X2_2275 ( .A(core__abc_22172_new_n1397_), .B(core__abc_22172_new_n1374_), .Y(core__abc_22172_new_n3070_));
AND2X2 AND2X2_2276 ( .A(core__abc_22172_new_n1517_), .B(core__abc_22172_new_n1534_), .Y(core__abc_22172_new_n3074_));
AND2X2 AND2X2_2277 ( .A(core__abc_22172_new_n1483_), .B(core__abc_22172_new_n1500_), .Y(core__abc_22172_new_n3075_));
AND2X2 AND2X2_2278 ( .A(core__abc_22172_new_n3074_), .B(core__abc_22172_new_n3075_), .Y(core__abc_22172_new_n3076_));
AND2X2 AND2X2_2279 ( .A(core__abc_22172_new_n1415_), .B(core__abc_22172_new_n1432_), .Y(core__abc_22172_new_n3077_));
AND2X2 AND2X2_228 ( .A(_abc_19873_new_n888_), .B(core_mi_16_), .Y(_abc_19873_new_n1274_));
AND2X2 AND2X2_2280 ( .A(core__abc_22172_new_n1449_), .B(core__abc_22172_new_n1466_), .Y(core__abc_22172_new_n3078_));
AND2X2 AND2X2_2281 ( .A(core__abc_22172_new_n3077_), .B(core__abc_22172_new_n3078_), .Y(core__abc_22172_new_n3079_));
AND2X2 AND2X2_2282 ( .A(core__abc_22172_new_n3076_), .B(core__abc_22172_new_n3079_), .Y(core__abc_22172_new_n3080_));
AND2X2 AND2X2_2283 ( .A(core__abc_22172_new_n3073_), .B(core__abc_22172_new_n3080_), .Y(core__abc_22172_new_n3081_));
AND2X2 AND2X2_2284 ( .A(core__abc_22172_new_n1413_), .B(core__abc_22172_new_n1430_), .Y(core__abc_22172_new_n3083_));
AND2X2 AND2X2_2285 ( .A(core__abc_22172_new_n3085_), .B(core__abc_22172_new_n3078_), .Y(core__abc_22172_new_n3086_));
AND2X2 AND2X2_2286 ( .A(core__abc_22172_new_n1465_), .B(core__abc_22172_new_n1446_), .Y(core__abc_22172_new_n3087_));
AND2X2 AND2X2_2287 ( .A(core__abc_22172_new_n3089_), .B(core__abc_22172_new_n3076_), .Y(core__abc_22172_new_n3090_));
AND2X2 AND2X2_2288 ( .A(core__abc_22172_new_n3091_), .B(core__abc_22172_new_n1498_), .Y(core__abc_22172_new_n3092_));
AND2X2 AND2X2_2289 ( .A(core__abc_22172_new_n3093_), .B(core__abc_22172_new_n3074_), .Y(core__abc_22172_new_n3094_));
AND2X2 AND2X2_229 ( .A(_abc_19873_new_n916_), .B(core_key_80_), .Y(_abc_19873_new_n1276_));
AND2X2 AND2X2_2290 ( .A(core__abc_22172_new_n1533_), .B(core__abc_22172_new_n1514_), .Y(core__abc_22172_new_n3095_));
AND2X2 AND2X2_2291 ( .A(core__abc_22172_new_n1789_), .B(core__abc_22172_new_n1806_), .Y(core__abc_22172_new_n3100_));
AND2X2 AND2X2_2292 ( .A(core__abc_22172_new_n1755_), .B(core__abc_22172_new_n1772_), .Y(core__abc_22172_new_n3101_));
AND2X2 AND2X2_2293 ( .A(core__abc_22172_new_n3100_), .B(core__abc_22172_new_n3101_), .Y(core__abc_22172_new_n3102_));
AND2X2 AND2X2_2294 ( .A(core__abc_22172_new_n1721_), .B(core__abc_22172_new_n1738_), .Y(core__abc_22172_new_n3103_));
AND2X2 AND2X2_2295 ( .A(core__abc_22172_new_n1687_), .B(core__abc_22172_new_n1704_), .Y(core__abc_22172_new_n3104_));
AND2X2 AND2X2_2296 ( .A(core__abc_22172_new_n3103_), .B(core__abc_22172_new_n3104_), .Y(core__abc_22172_new_n3105_));
AND2X2 AND2X2_2297 ( .A(core__abc_22172_new_n3102_), .B(core__abc_22172_new_n3105_), .Y(core__abc_22172_new_n3106_));
AND2X2 AND2X2_2298 ( .A(core__abc_22172_new_n1653_), .B(core__abc_22172_new_n1670_), .Y(core__abc_22172_new_n3107_));
AND2X2 AND2X2_2299 ( .A(core__abc_22172_new_n1619_), .B(core__abc_22172_new_n1636_), .Y(core__abc_22172_new_n3108_));
AND2X2 AND2X2_23 ( .A(_abc_19873_new_n901_), .B(core_key_0_), .Y(_abc_19873_new_n902_));
AND2X2 AND2X2_230 ( .A(_abc_19873_new_n925_), .B(word2_reg_16_), .Y(_abc_19873_new_n1279_));
AND2X2 AND2X2_2300 ( .A(core__abc_22172_new_n3107_), .B(core__abc_22172_new_n3108_), .Y(core__abc_22172_new_n3109_));
AND2X2 AND2X2_2301 ( .A(core__abc_22172_new_n1585_), .B(core__abc_22172_new_n1602_), .Y(core__abc_22172_new_n3110_));
AND2X2 AND2X2_2302 ( .A(core__abc_22172_new_n1551_), .B(core__abc_22172_new_n1568_), .Y(core__abc_22172_new_n3111_));
AND2X2 AND2X2_2303 ( .A(core__abc_22172_new_n3110_), .B(core__abc_22172_new_n3111_), .Y(core__abc_22172_new_n3112_));
AND2X2 AND2X2_2304 ( .A(core__abc_22172_new_n3109_), .B(core__abc_22172_new_n3112_), .Y(core__abc_22172_new_n3113_));
AND2X2 AND2X2_2305 ( .A(core__abc_22172_new_n3106_), .B(core__abc_22172_new_n3113_), .Y(core__abc_22172_new_n3114_));
AND2X2 AND2X2_2306 ( .A(core__abc_22172_new_n3099_), .B(core__abc_22172_new_n3114_), .Y(core__abc_22172_new_n3115_));
AND2X2 AND2X2_2307 ( .A(core__abc_22172_new_n3116_), .B(core__abc_22172_new_n1566_), .Y(core__abc_22172_new_n3117_));
AND2X2 AND2X2_2308 ( .A(core__abc_22172_new_n3118_), .B(core__abc_22172_new_n3110_), .Y(core__abc_22172_new_n3119_));
AND2X2 AND2X2_2309 ( .A(core__abc_22172_new_n1601_), .B(core__abc_22172_new_n1582_), .Y(core__abc_22172_new_n3120_));
AND2X2 AND2X2_231 ( .A(_abc_19873_new_n907_), .B(word1_reg_16_), .Y(_abc_19873_new_n1280_));
AND2X2 AND2X2_2310 ( .A(core__abc_22172_new_n3122_), .B(core__abc_22172_new_n3109_), .Y(core__abc_22172_new_n3123_));
AND2X2 AND2X2_2311 ( .A(core__abc_22172_new_n1617_), .B(core__abc_22172_new_n1634_), .Y(core__abc_22172_new_n3125_));
AND2X2 AND2X2_2312 ( .A(core__abc_22172_new_n3127_), .B(core__abc_22172_new_n3107_), .Y(core__abc_22172_new_n3128_));
AND2X2 AND2X2_2313 ( .A(core__abc_22172_new_n1669_), .B(core__abc_22172_new_n1650_), .Y(core__abc_22172_new_n3129_));
AND2X2 AND2X2_2314 ( .A(core__abc_22172_new_n3132_), .B(core__abc_22172_new_n3106_), .Y(core__abc_22172_new_n3133_));
AND2X2 AND2X2_2315 ( .A(core__abc_22172_new_n1685_), .B(core__abc_22172_new_n1702_), .Y(core__abc_22172_new_n3135_));
AND2X2 AND2X2_2316 ( .A(core__abc_22172_new_n3137_), .B(core__abc_22172_new_n3103_), .Y(core__abc_22172_new_n3138_));
AND2X2 AND2X2_2317 ( .A(core__abc_22172_new_n1737_), .B(core__abc_22172_new_n1718_), .Y(core__abc_22172_new_n3139_));
AND2X2 AND2X2_2318 ( .A(core__abc_22172_new_n3141_), .B(core__abc_22172_new_n3102_), .Y(core__abc_22172_new_n3142_));
AND2X2 AND2X2_2319 ( .A(core__abc_22172_new_n1805_), .B(core__abc_22172_new_n1786_), .Y(core__abc_22172_new_n3143_));
AND2X2 AND2X2_232 ( .A(_abc_19873_new_n912_), .B(word3_reg_16_), .Y(_abc_19873_new_n1281_));
AND2X2 AND2X2_2320 ( .A(core__abc_22172_new_n1753_), .B(core__abc_22172_new_n1770_), .Y(core__abc_22172_new_n3146_));
AND2X2 AND2X2_2321 ( .A(core__abc_22172_new_n3148_), .B(core__abc_22172_new_n3100_), .Y(core__abc_22172_new_n3149_));
AND2X2 AND2X2_2322 ( .A(core__abc_22172_new_n1925_), .B(core__abc_22172_new_n1942_), .Y(core__abc_22172_new_n3154_));
AND2X2 AND2X2_2323 ( .A(core__abc_22172_new_n1891_), .B(core__abc_22172_new_n1908_), .Y(core__abc_22172_new_n3155_));
AND2X2 AND2X2_2324 ( .A(core__abc_22172_new_n3154_), .B(core__abc_22172_new_n3155_), .Y(core__abc_22172_new_n3156_));
AND2X2 AND2X2_2325 ( .A(core__abc_22172_new_n1823_), .B(core__abc_22172_new_n1840_), .Y(core__abc_22172_new_n3157_));
AND2X2 AND2X2_2326 ( .A(core__abc_22172_new_n1857_), .B(core__abc_22172_new_n1874_), .Y(core__abc_22172_new_n3158_));
AND2X2 AND2X2_2327 ( .A(core__abc_22172_new_n3157_), .B(core__abc_22172_new_n3158_), .Y(core__abc_22172_new_n3159_));
AND2X2 AND2X2_2328 ( .A(core__abc_22172_new_n3156_), .B(core__abc_22172_new_n3159_), .Y(core__abc_22172_new_n3160_));
AND2X2 AND2X2_2329 ( .A(core__abc_22172_new_n3153_), .B(core__abc_22172_new_n3160_), .Y(core__abc_22172_new_n3161_));
AND2X2 AND2X2_233 ( .A(_abc_19873_new_n919_), .B(core_mi_48_), .Y(_abc_19873_new_n1284_));
AND2X2 AND2X2_2330 ( .A(core__abc_22172_new_n1821_), .B(core__abc_22172_new_n1838_), .Y(core__abc_22172_new_n3163_));
AND2X2 AND2X2_2331 ( .A(core__abc_22172_new_n3165_), .B(core__abc_22172_new_n3158_), .Y(core__abc_22172_new_n3166_));
AND2X2 AND2X2_2332 ( .A(core__abc_22172_new_n1873_), .B(core__abc_22172_new_n1855_), .Y(core__abc_22172_new_n3167_));
AND2X2 AND2X2_2333 ( .A(core__abc_22172_new_n3169_), .B(core__abc_22172_new_n3156_), .Y(core__abc_22172_new_n3170_));
AND2X2 AND2X2_2334 ( .A(core__abc_22172_new_n1941_), .B(core__abc_22172_new_n1923_), .Y(core__abc_22172_new_n3171_));
AND2X2 AND2X2_2335 ( .A(core__abc_22172_new_n1890_), .B(core__abc_22172_new_n1906_), .Y(core__abc_22172_new_n3174_));
AND2X2 AND2X2_2336 ( .A(core__abc_22172_new_n3176_), .B(core__abc_22172_new_n3154_), .Y(core__abc_22172_new_n3177_));
AND2X2 AND2X2_2337 ( .A(core__abc_22172_new_n1959_), .B(core__abc_22172_new_n1976_), .Y(core__abc_22172_new_n3181_));
AND2X2 AND2X2_2338 ( .A(core__abc_22172_new_n3180_), .B(core__abc_22172_new_n3181_), .Y(core__abc_22172_new_n3182_));
AND2X2 AND2X2_2339 ( .A(core__abc_22172_new_n3183_), .B(core__abc_22172_new_n1993_), .Y(core__abc_22172_new_n3184_));
AND2X2 AND2X2_234 ( .A(_abc_19873_new_n930_), .B(word0_reg_16_), .Y(_abc_19873_new_n1285_));
AND2X2 AND2X2_2340 ( .A(core__abc_22172_new_n3186_), .B(core__abc_22172_new_n2013_), .Y(core__abc_22172_new_n3187_));
AND2X2 AND2X2_2341 ( .A(core__abc_22172_new_n3185_), .B(core__abc_22172_new_n2010_), .Y(core__abc_22172_new_n3188_));
AND2X2 AND2X2_2342 ( .A(core__abc_22172_new_n3189_), .B(core_v3_reg_27_), .Y(core__abc_22172_new_n3190_));
AND2X2 AND2X2_2343 ( .A(core__abc_22172_new_n3191_), .B(core__abc_22172_new_n3192_), .Y(core__abc_22172_new_n3193_));
AND2X2 AND2X2_2344 ( .A(core__abc_22172_new_n2659_), .B(core__abc_22172_new_n1253_), .Y(core__abc_22172_new_n3196_));
AND2X2 AND2X2_2345 ( .A(core__abc_22172_new_n3197_), .B(core__abc_22172_new_n1169_), .Y(core__abc_22172_new_n3198_));
AND2X2 AND2X2_2346 ( .A(core__abc_22172_new_n2659_), .B(core__abc_22172_new_n1216_), .Y(core__abc_22172_new_n3200_));
AND2X2 AND2X2_2347 ( .A(core__abc_22172_new_n3201_), .B(core__abc_22172_new_n1218_), .Y(core__abc_22172_new_n3202_));
AND2X2 AND2X2_2348 ( .A(core__abc_22172_new_n3204_), .B(core__abc_22172_new_n2624_), .Y(core__abc_22172_new_n3205_));
AND2X2 AND2X2_2349 ( .A(core__abc_22172_new_n3206_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n3207_));
AND2X2 AND2X2_235 ( .A(_abc_19873_new_n928_), .B(core_key_48_), .Y(_abc_19873_new_n1287_));
AND2X2 AND2X2_2350 ( .A(core__abc_22172_new_n3207_), .B(core__abc_22172_new_n3195_), .Y(core__abc_22172_new_n3208_));
AND2X2 AND2X2_2351 ( .A(core__abc_22172_new_n2659_), .B(core__abc_22172_new_n1226_), .Y(core__abc_22172_new_n3209_));
AND2X2 AND2X2_2352 ( .A(core__abc_22172_new_n1170_), .B(core__abc_22172_new_n1169_), .Y(core__abc_22172_new_n3210_));
AND2X2 AND2X2_2353 ( .A(core__abc_22172_new_n2623_), .B(core__abc_22172_new_n3210_), .Y(core__abc_22172_new_n3211_));
AND2X2 AND2X2_2354 ( .A(core__abc_22172_new_n3198_), .B(core__abc_22172_new_n3201_), .Y(core__abc_22172_new_n3213_));
AND2X2 AND2X2_2355 ( .A(core__abc_22172_new_n3213_), .B(core__abc_22172_new_n2623_), .Y(core__abc_22172_new_n3214_));
AND2X2 AND2X2_2356 ( .A(core__abc_22172_new_n3215_), .B(core__abc_22172_new_n3203_), .Y(core__abc_22172_new_n3216_));
AND2X2 AND2X2_2357 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n3218_), .Y(core__abc_22172_new_n3219_));
AND2X2 AND2X2_2358 ( .A(core_v3_reg_0_), .B(core_mi_0_), .Y(core__abc_22172_new_n3220_));
AND2X2 AND2X2_2359 ( .A(core__abc_22172_new_n3221_), .B(core__abc_22172_new_n3222_), .Y(core__abc_22172_new_n3223_));
AND2X2 AND2X2_236 ( .A(_abc_19873_new_n901_), .B(core_key_16_), .Y(_abc_19873_new_n1288_));
AND2X2 AND2X2_2360 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n3223_), .Y(core__abc_22172_new_n3224_));
AND2X2 AND2X2_2361 ( .A(core__abc_22172_new_n3229_), .B(reset_n), .Y(core__abc_22172_new_n3230_));
AND2X2 AND2X2_2362 ( .A(core__abc_22172_new_n3227_), .B(core__abc_22172_new_n3230_), .Y(core__0v3_reg_63_0__0_));
AND2X2 AND2X2_2363 ( .A(core__abc_22172_new_n1842_), .B(core__abc_22172_new_n1818_), .Y(core__abc_22172_new_n3233_));
AND2X2 AND2X2_2364 ( .A(core__abc_22172_new_n3232_), .B(core__abc_22172_new_n3233_), .Y(core__abc_22172_new_n3234_));
AND2X2 AND2X2_2365 ( .A(core__abc_22172_new_n1836_), .B(core__abc_22172_new_n1817_), .Y(core__abc_22172_new_n3235_));
AND2X2 AND2X2_2366 ( .A(core__abc_22172_new_n1819_), .B(core__abc_22172_new_n1836_), .Y(core__abc_22172_new_n3236_));
AND2X2 AND2X2_2367 ( .A(core__abc_22172_new_n3013_), .B(core__abc_22172_new_n3236_), .Y(core__abc_22172_new_n3237_));
AND2X2 AND2X2_2368 ( .A(core__abc_22172_new_n1283_), .B(core__abc_22172_new_n3053_), .Y(core__abc_22172_new_n3242_));
AND2X2 AND2X2_2369 ( .A(core__abc_22172_new_n3245_), .B(core__abc_22172_new_n3246_), .Y(core__abc_22172_new_n3247_));
AND2X2 AND2X2_237 ( .A(_abc_19873_new_n1292_), .B(_abc_19873_new_n937_), .Y(\read_data[16] ));
AND2X2 AND2X2_2370 ( .A(core__abc_22172_new_n3239_), .B(core__abc_22172_new_n3247_), .Y(core__abc_22172_new_n3248_));
AND2X2 AND2X2_2371 ( .A(core__abc_22172_new_n3249_), .B(core__abc_22172_new_n3250_), .Y(core__abc_22172_new_n3251_));
AND2X2 AND2X2_2372 ( .A(core__abc_22172_new_n3251_), .B(core__abc_22172_new_n3042_), .Y(core__abc_22172_new_n3252_));
AND2X2 AND2X2_2373 ( .A(core__abc_22172_new_n3253_), .B(core__abc_22172_new_n3254_), .Y(core__abc_22172_new_n3255_));
AND2X2 AND2X2_2374 ( .A(core__abc_22172_new_n1993_), .B(core__abc_22172_new_n2010_), .Y(core__abc_22172_new_n3257_));
AND2X2 AND2X2_2375 ( .A(core__abc_22172_new_n3048_), .B(core__abc_22172_new_n3257_), .Y(core__abc_22172_new_n3258_));
AND2X2 AND2X2_2376 ( .A(core__abc_22172_new_n2007_), .B(core__abc_22172_new_n1990_), .Y(core__abc_22172_new_n3259_));
AND2X2 AND2X2_2377 ( .A(core__abc_22172_new_n3181_), .B(core__abc_22172_new_n3257_), .Y(core__abc_22172_new_n3262_));
AND2X2 AND2X2_2378 ( .A(core__abc_22172_new_n3180_), .B(core__abc_22172_new_n3262_), .Y(core__abc_22172_new_n3263_));
AND2X2 AND2X2_2379 ( .A(core__abc_22172_new_n3265_), .B(core__abc_22172_new_n2030_), .Y(core__abc_22172_new_n3266_));
AND2X2 AND2X2_238 ( .A(_abc_19873_new_n901_), .B(core_key_17_), .Y(_abc_19873_new_n1294_));
AND2X2 AND2X2_2380 ( .A(core__abc_22172_new_n3264_), .B(core__abc_22172_new_n2027_), .Y(core__abc_22172_new_n3267_));
AND2X2 AND2X2_2381 ( .A(core__abc_22172_new_n3270_), .B(core__abc_22172_new_n3271_), .Y(core__abc_22172_new_n3272_));
AND2X2 AND2X2_2382 ( .A(core__abc_22172_new_n3276_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n3277_));
AND2X2 AND2X2_2383 ( .A(core__abc_22172_new_n3277_), .B(core__abc_22172_new_n3274_), .Y(core__abc_22172_new_n3278_));
AND2X2 AND2X2_2384 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n3279_), .Y(core__abc_22172_new_n3280_));
AND2X2 AND2X2_2385 ( .A(core_v3_reg_1_), .B(core_mi_1_), .Y(core__abc_22172_new_n3281_));
AND2X2 AND2X2_2386 ( .A(core__abc_22172_new_n3282_), .B(core__abc_22172_new_n3283_), .Y(core__abc_22172_new_n3284_));
AND2X2 AND2X2_2387 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n3284_), .Y(core__abc_22172_new_n3285_));
AND2X2 AND2X2_2388 ( .A(core__abc_22172_new_n3289_), .B(reset_n), .Y(core__abc_22172_new_n3290_));
AND2X2 AND2X2_2389 ( .A(core__abc_22172_new_n3288_), .B(core__abc_22172_new_n3290_), .Y(core__0v3_reg_63_0__1_));
AND2X2 AND2X2_239 ( .A(_abc_19873_new_n919_), .B(core_mi_49_), .Y(_abc_19873_new_n1297_));
AND2X2 AND2X2_2390 ( .A(core__abc_22172_new_n3294_), .B(core__abc_22172_new_n1835_), .Y(core__abc_22172_new_n3295_));
AND2X2 AND2X2_2391 ( .A(core__abc_22172_new_n3297_), .B(core__abc_22172_new_n1853_), .Y(core__abc_22172_new_n3298_));
AND2X2 AND2X2_2392 ( .A(core__abc_22172_new_n3299_), .B(core__abc_22172_new_n3300_), .Y(core__abc_22172_new_n3301_));
AND2X2 AND2X2_2393 ( .A(core__abc_22172_new_n3304_), .B(core__abc_22172_new_n1306_), .Y(core__abc_22172_new_n3305_));
AND2X2 AND2X2_2394 ( .A(core__abc_22172_new_n3055_), .B(core__abc_22172_new_n1305_), .Y(core__abc_22172_new_n3306_));
AND2X2 AND2X2_2395 ( .A(core__abc_22172_new_n3309_), .B(core__abc_22172_new_n3310_), .Y(core__abc_22172_new_n3311_));
AND2X2 AND2X2_2396 ( .A(core__abc_22172_new_n3302_), .B(core__abc_22172_new_n3311_), .Y(core__abc_22172_new_n3312_));
AND2X2 AND2X2_2397 ( .A(core__abc_22172_new_n3301_), .B(core__abc_22172_new_n3313_), .Y(core__abc_22172_new_n3314_));
AND2X2 AND2X2_2398 ( .A(core__abc_22172_new_n3293_), .B(core__abc_22172_new_n3316_), .Y(core__abc_22172_new_n3317_));
AND2X2 AND2X2_2399 ( .A(core__abc_22172_new_n3318_), .B(core__abc_22172_new_n3319_), .Y(core__abc_22172_new_n3320_));
AND2X2 AND2X2_24 ( .A(_abc_19873_new_n884_), .B(\addr[0] ), .Y(_abc_19873_new_n903_));
AND2X2 AND2X2_240 ( .A(_abc_19873_new_n930_), .B(word0_reg_17_), .Y(_abc_19873_new_n1298_));
AND2X2 AND2X2_2400 ( .A(core__abc_22172_new_n3322_), .B(core__abc_22172_new_n2047_), .Y(core__abc_22172_new_n3323_));
AND2X2 AND2X2_2401 ( .A(core__abc_22172_new_n3321_), .B(core__abc_22172_new_n2044_), .Y(core__abc_22172_new_n3324_));
AND2X2 AND2X2_2402 ( .A(core__abc_22172_new_n3325_), .B(core_v3_reg_29_), .Y(core__abc_22172_new_n3326_));
AND2X2 AND2X2_2403 ( .A(core__abc_22172_new_n3327_), .B(core__abc_22172_new_n3328_), .Y(core__abc_22172_new_n3329_));
AND2X2 AND2X2_2404 ( .A(core__abc_22172_new_n3333_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n3334_));
AND2X2 AND2X2_2405 ( .A(core__abc_22172_new_n3334_), .B(core__abc_22172_new_n3331_), .Y(core__abc_22172_new_n3335_));
AND2X2 AND2X2_2406 ( .A(core__abc_22172_new_n3214_), .B(core_key_66_), .Y(core__abc_22172_new_n3336_));
AND2X2 AND2X2_2407 ( .A(core_v3_reg_2_), .B(core_mi_2_), .Y(core__abc_22172_new_n3337_));
AND2X2 AND2X2_2408 ( .A(core__abc_22172_new_n3338_), .B(core__abc_22172_new_n3339_), .Y(core__abc_22172_new_n3340_));
AND2X2 AND2X2_2409 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n3340_), .Y(core__abc_22172_new_n3341_));
AND2X2 AND2X2_241 ( .A(_abc_19873_new_n925_), .B(word2_reg_17_), .Y(_abc_19873_new_n1301_));
AND2X2 AND2X2_2410 ( .A(core__abc_22172_new_n3345_), .B(reset_n), .Y(core__abc_22172_new_n3346_));
AND2X2 AND2X2_2411 ( .A(core__abc_22172_new_n3344_), .B(core__abc_22172_new_n3346_), .Y(core__0v3_reg_63_0__2_));
AND2X2 AND2X2_2412 ( .A(core__abc_22172_new_n2027_), .B(core__abc_22172_new_n2044_), .Y(core__abc_22172_new_n3348_));
AND2X2 AND2X2_2413 ( .A(core__abc_22172_new_n3264_), .B(core__abc_22172_new_n3348_), .Y(core__abc_22172_new_n3349_));
AND2X2 AND2X2_2414 ( .A(core__abc_22172_new_n2026_), .B(core__abc_22172_new_n2043_), .Y(core__abc_22172_new_n3351_));
AND2X2 AND2X2_2415 ( .A(core__abc_22172_new_n3354_), .B(core__abc_22172_new_n2061_), .Y(core__abc_22172_new_n3355_));
AND2X2 AND2X2_2416 ( .A(core__abc_22172_new_n3356_), .B(core__abc_22172_new_n2064_), .Y(core__abc_22172_new_n3357_));
AND2X2 AND2X2_2417 ( .A(core__abc_22172_new_n3360_), .B(core__abc_22172_new_n3362_), .Y(core__abc_22172_new_n3363_));
AND2X2 AND2X2_2418 ( .A(core__abc_22172_new_n3299_), .B(core__abc_22172_new_n1852_), .Y(core__abc_22172_new_n3365_));
AND2X2 AND2X2_2419 ( .A(core__abc_22172_new_n3365_), .B(core__abc_22172_new_n1876_), .Y(core__abc_22172_new_n3366_));
AND2X2 AND2X2_242 ( .A(_abc_19873_new_n907_), .B(word1_reg_17_), .Y(_abc_19873_new_n1302_));
AND2X2 AND2X2_2420 ( .A(core__abc_22172_new_n3367_), .B(core__abc_22172_new_n3368_), .Y(core__abc_22172_new_n3369_));
AND2X2 AND2X2_2421 ( .A(core__abc_22172_new_n3371_), .B(core__abc_22172_new_n3370_), .Y(core__abc_22172_new_n3372_));
AND2X2 AND2X2_2422 ( .A(core__abc_22172_new_n3373_), .B(core__abc_22172_new_n1322_), .Y(core__abc_22172_new_n3374_));
AND2X2 AND2X2_2423 ( .A(core__abc_22172_new_n3372_), .B(core__abc_22172_new_n1323_), .Y(core__abc_22172_new_n3375_));
AND2X2 AND2X2_2424 ( .A(core__abc_22172_new_n3376_), .B(core_v3_reg_51_), .Y(core__abc_22172_new_n3377_));
AND2X2 AND2X2_2425 ( .A(core__abc_22172_new_n3378_), .B(core__abc_22172_new_n3379_), .Y(core__abc_22172_new_n3380_));
AND2X2 AND2X2_2426 ( .A(core__abc_22172_new_n3369_), .B(core__abc_22172_new_n3380_), .Y(core__abc_22172_new_n3381_));
AND2X2 AND2X2_2427 ( .A(core__abc_22172_new_n3383_), .B(core__abc_22172_new_n3384_), .Y(core__abc_22172_new_n3385_));
AND2X2 AND2X2_2428 ( .A(core__abc_22172_new_n3386_), .B(core__abc_22172_new_n3382_), .Y(core__abc_22172_new_n3387_));
AND2X2 AND2X2_2429 ( .A(core__abc_22172_new_n3391_), .B(core__abc_22172_new_n3389_), .Y(core__abc_22172_new_n3392_));
AND2X2 AND2X2_243 ( .A(_abc_19873_new_n912_), .B(word3_reg_17_), .Y(_abc_19873_new_n1303_));
AND2X2 AND2X2_2430 ( .A(core__abc_22172_new_n3396_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n3397_));
AND2X2 AND2X2_2431 ( .A(core__abc_22172_new_n3397_), .B(core__abc_22172_new_n3394_), .Y(core__abc_22172_new_n3398_));
AND2X2 AND2X2_2432 ( .A(core__abc_22172_new_n3214_), .B(core_key_67_), .Y(core__abc_22172_new_n3399_));
AND2X2 AND2X2_2433 ( .A(core_v3_reg_3_), .B(core_mi_3_), .Y(core__abc_22172_new_n3400_));
AND2X2 AND2X2_2434 ( .A(core__abc_22172_new_n3401_), .B(core__abc_22172_new_n3402_), .Y(core__abc_22172_new_n3403_));
AND2X2 AND2X2_2435 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n3403_), .Y(core__abc_22172_new_n3404_));
AND2X2 AND2X2_2436 ( .A(core__abc_22172_new_n3408_), .B(reset_n), .Y(core__abc_22172_new_n3409_));
AND2X2 AND2X2_2437 ( .A(core__abc_22172_new_n3407_), .B(core__abc_22172_new_n3409_), .Y(core__0v3_reg_63_0__3_));
AND2X2 AND2X2_2438 ( .A(core__abc_22172_new_n1853_), .B(core__abc_22172_new_n1870_), .Y(core__abc_22172_new_n3411_));
AND2X2 AND2X2_2439 ( .A(core__abc_22172_new_n3296_), .B(core__abc_22172_new_n3411_), .Y(core__abc_22172_new_n3412_));
AND2X2 AND2X2_244 ( .A(_abc_19873_new_n928_), .B(core_key_49_), .Y(_abc_19873_new_n1306_));
AND2X2 AND2X2_2440 ( .A(core__abc_22172_new_n1867_), .B(core__abc_22172_new_n1851_), .Y(core__abc_22172_new_n3413_));
AND2X2 AND2X2_2441 ( .A(core__abc_22172_new_n3236_), .B(core__abc_22172_new_n3411_), .Y(core__abc_22172_new_n3416_));
AND2X2 AND2X2_2442 ( .A(core__abc_22172_new_n3013_), .B(core__abc_22172_new_n3416_), .Y(core__abc_22172_new_n3417_));
AND2X2 AND2X2_2443 ( .A(core__abc_22172_new_n3418_), .B(core__abc_22172_new_n1887_), .Y(core__abc_22172_new_n3419_));
AND2X2 AND2X2_2444 ( .A(core__abc_22172_new_n3420_), .B(core__abc_22172_new_n1893_), .Y(core__abc_22172_new_n3421_));
AND2X2 AND2X2_2445 ( .A(core__abc_22172_new_n3059_), .B(core__abc_22172_new_n1340_), .Y(core__abc_22172_new_n3424_));
AND2X2 AND2X2_2446 ( .A(core__abc_22172_new_n3060_), .B(core__abc_22172_new_n1341_), .Y(core__abc_22172_new_n3425_));
AND2X2 AND2X2_2447 ( .A(core__abc_22172_new_n3426_), .B(core__abc_22172_new_n3423_), .Y(core__abc_22172_new_n3427_));
AND2X2 AND2X2_2448 ( .A(core__abc_22172_new_n3428_), .B(core_v3_reg_52_), .Y(core__abc_22172_new_n3429_));
AND2X2 AND2X2_2449 ( .A(core__abc_22172_new_n3422_), .B(core__abc_22172_new_n3430_), .Y(core__abc_22172_new_n3431_));
AND2X2 AND2X2_245 ( .A(_abc_19873_new_n916_), .B(core_key_81_), .Y(_abc_19873_new_n1307_));
AND2X2 AND2X2_2450 ( .A(core__abc_22172_new_n3432_), .B(core__abc_22172_new_n3433_), .Y(core__abc_22172_new_n3434_));
AND2X2 AND2X2_2451 ( .A(core__abc_22172_new_n3364_), .B(core__abc_22172_new_n3386_), .Y(core__abc_22172_new_n3437_));
AND2X2 AND2X2_2452 ( .A(core__abc_22172_new_n3438_), .B(core__abc_22172_new_n3436_), .Y(core__abc_22172_new_n3439_));
AND2X2 AND2X2_2453 ( .A(core__abc_22172_new_n3440_), .B(core__abc_22172_new_n3441_), .Y(core__abc_22172_new_n3442_));
AND2X2 AND2X2_2454 ( .A(core__abc_22172_new_n3444_), .B(core__abc_22172_new_n2081_), .Y(core__abc_22172_new_n3445_));
AND2X2 AND2X2_2455 ( .A(core__abc_22172_new_n3443_), .B(core__abc_22172_new_n2078_), .Y(core__abc_22172_new_n3446_));
AND2X2 AND2X2_2456 ( .A(core__abc_22172_new_n3447_), .B(core_v3_reg_31_), .Y(core__abc_22172_new_n3448_));
AND2X2 AND2X2_2457 ( .A(core__abc_22172_new_n3450_), .B(core__abc_22172_new_n3449_), .Y(core__abc_22172_new_n3451_));
AND2X2 AND2X2_2458 ( .A(core__abc_22172_new_n3455_), .B(core__abc_22172_new_n3456_), .Y(core__abc_22172_new_n3457_));
AND2X2 AND2X2_2459 ( .A(core__abc_22172_new_n3458_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n3459_));
AND2X2 AND2X2_246 ( .A(_abc_19873_new_n881_), .B(core_key_113_), .Y(_abc_19873_new_n1309_));
AND2X2 AND2X2_2460 ( .A(core__abc_22172_new_n3459_), .B(core__abc_22172_new_n3453_), .Y(core__abc_22172_new_n3460_));
AND2X2 AND2X2_2461 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n3461_), .Y(core__abc_22172_new_n3462_));
AND2X2 AND2X2_2462 ( .A(core_v3_reg_4_), .B(core_mi_4_), .Y(core__abc_22172_new_n3463_));
AND2X2 AND2X2_2463 ( .A(core__abc_22172_new_n3464_), .B(core__abc_22172_new_n3465_), .Y(core__abc_22172_new_n3466_));
AND2X2 AND2X2_2464 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n3466_), .Y(core__abc_22172_new_n3467_));
AND2X2 AND2X2_2465 ( .A(core__abc_22172_new_n3471_), .B(reset_n), .Y(core__abc_22172_new_n3472_));
AND2X2 AND2X2_2466 ( .A(core__abc_22172_new_n3470_), .B(core__abc_22172_new_n3472_), .Y(core__0v3_reg_63_0__4_));
AND2X2 AND2X2_2467 ( .A(core__abc_22172_new_n3476_), .B(core__abc_22172_new_n1904_), .Y(core__abc_22172_new_n3478_));
AND2X2 AND2X2_2468 ( .A(core__abc_22172_new_n3479_), .B(core__abc_22172_new_n3477_), .Y(core__abc_22172_new_n3480_));
AND2X2 AND2X2_2469 ( .A(core__abc_22172_new_n3483_), .B(core__abc_22172_new_n1363_), .Y(core__abc_22172_new_n3484_));
AND2X2 AND2X2_247 ( .A(_abc_19873_new_n888_), .B(core_mi_17_), .Y(_abc_19873_new_n1310_));
AND2X2 AND2X2_2470 ( .A(core__abc_22172_new_n3482_), .B(core__abc_22172_new_n1360_), .Y(core__abc_22172_new_n3485_));
AND2X2 AND2X2_2471 ( .A(core__abc_22172_new_n3486_), .B(core__abc_22172_new_n3481_), .Y(core__abc_22172_new_n3487_));
AND2X2 AND2X2_2472 ( .A(core__abc_22172_new_n3488_), .B(core_v3_reg_53_), .Y(core__abc_22172_new_n3489_));
AND2X2 AND2X2_2473 ( .A(core__abc_22172_new_n3480_), .B(core__abc_22172_new_n3491_), .Y(core__abc_22172_new_n3492_));
AND2X2 AND2X2_2474 ( .A(core__abc_22172_new_n3493_), .B(core__abc_22172_new_n3494_), .Y(core__abc_22172_new_n3495_));
AND2X2 AND2X2_2475 ( .A(core__abc_22172_new_n3496_), .B(core__abc_22172_new_n3498_), .Y(core__abc_22172_new_n3499_));
AND2X2 AND2X2_2476 ( .A(core__abc_22172_new_n2061_), .B(core__abc_22172_new_n2078_), .Y(core__abc_22172_new_n3502_));
AND2X2 AND2X2_2477 ( .A(core__abc_22172_new_n3348_), .B(core__abc_22172_new_n3502_), .Y(core__abc_22172_new_n3503_));
AND2X2 AND2X2_2478 ( .A(core__abc_22172_new_n3261_), .B(core__abc_22172_new_n3503_), .Y(core__abc_22172_new_n3504_));
AND2X2 AND2X2_2479 ( .A(core__abc_22172_new_n3353_), .B(core__abc_22172_new_n3502_), .Y(core__abc_22172_new_n3505_));
AND2X2 AND2X2_248 ( .A(_abc_19873_new_n1314_), .B(_abc_19873_new_n937_), .Y(\read_data[17] ));
AND2X2 AND2X2_2480 ( .A(core__abc_22172_new_n2075_), .B(core__abc_22172_new_n2059_), .Y(core__abc_22172_new_n3506_));
AND2X2 AND2X2_2481 ( .A(core__abc_22172_new_n3263_), .B(core__abc_22172_new_n3503_), .Y(core__abc_22172_new_n3510_));
AND2X2 AND2X2_2482 ( .A(core__abc_22172_new_n3512_), .B(core__abc_22172_new_n2098_), .Y(core__abc_22172_new_n3513_));
AND2X2 AND2X2_2483 ( .A(core__abc_22172_new_n3511_), .B(core__abc_22172_new_n2095_), .Y(core__abc_22172_new_n3514_));
AND2X2 AND2X2_2484 ( .A(core__abc_22172_new_n3517_), .B(core__abc_22172_new_n3518_), .Y(core__abc_22172_new_n3519_));
AND2X2 AND2X2_2485 ( .A(core__abc_22172_new_n3522_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n3523_));
AND2X2 AND2X2_2486 ( .A(core__abc_22172_new_n3523_), .B(core__abc_22172_new_n3521_), .Y(core__abc_22172_new_n3524_));
AND2X2 AND2X2_2487 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n3525_), .Y(core__abc_22172_new_n3526_));
AND2X2 AND2X2_2488 ( .A(core_v3_reg_5_), .B(core_mi_5_), .Y(core__abc_22172_new_n3527_));
AND2X2 AND2X2_2489 ( .A(core__abc_22172_new_n3528_), .B(core__abc_22172_new_n3529_), .Y(core__abc_22172_new_n3530_));
AND2X2 AND2X2_249 ( .A(_abc_19873_new_n912_), .B(word3_reg_18_), .Y(_abc_19873_new_n1316_));
AND2X2 AND2X2_2490 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n3530_), .Y(core__abc_22172_new_n3531_));
AND2X2 AND2X2_2491 ( .A(core__abc_22172_new_n3535_), .B(reset_n), .Y(core__abc_22172_new_n3536_));
AND2X2 AND2X2_2492 ( .A(core__abc_22172_new_n3534_), .B(core__abc_22172_new_n3536_), .Y(core__0v3_reg_63_0__5_));
AND2X2 AND2X2_2493 ( .A(core__abc_22172_new_n1886_), .B(core__abc_22172_new_n1903_), .Y(core__abc_22172_new_n3539_));
AND2X2 AND2X2_2494 ( .A(core__abc_22172_new_n1887_), .B(core__abc_22172_new_n1904_), .Y(core__abc_22172_new_n3542_));
AND2X2 AND2X2_2495 ( .A(core__abc_22172_new_n3418_), .B(core__abc_22172_new_n3542_), .Y(core__abc_22172_new_n3543_));
AND2X2 AND2X2_2496 ( .A(core__abc_22172_new_n3544_), .B(core__abc_22172_new_n1921_), .Y(core__abc_22172_new_n3545_));
AND2X2 AND2X2_2497 ( .A(core__abc_22172_new_n3546_), .B(core__abc_22172_new_n1927_), .Y(core__abc_22172_new_n3547_));
AND2X2 AND2X2_2498 ( .A(core__abc_22172_new_n3551_), .B(core__abc_22172_new_n3067_), .Y(core__abc_22172_new_n3552_));
AND2X2 AND2X2_2499 ( .A(core__abc_22172_new_n3553_), .B(core__abc_22172_new_n1379_), .Y(core__abc_22172_new_n3554_));
AND2X2 AND2X2_25 ( .A(_abc_19873_new_n879_), .B(_abc_19873_new_n903_), .Y(_abc_19873_new_n904_));
AND2X2 AND2X2_250 ( .A(_abc_19873_new_n901_), .B(core_key_18_), .Y(_abc_19873_new_n1317_));
AND2X2 AND2X2_2500 ( .A(core__abc_22172_new_n3552_), .B(core__abc_22172_new_n1378_), .Y(core__abc_22172_new_n3555_));
AND2X2 AND2X2_2501 ( .A(core__abc_22172_new_n3558_), .B(core__abc_22172_new_n3559_), .Y(core__abc_22172_new_n3560_));
AND2X2 AND2X2_2502 ( .A(core__abc_22172_new_n3548_), .B(core__abc_22172_new_n3560_), .Y(core__abc_22172_new_n3561_));
AND2X2 AND2X2_2503 ( .A(core__abc_22172_new_n3562_), .B(core__abc_22172_new_n3563_), .Y(core__abc_22172_new_n3564_));
AND2X2 AND2X2_2504 ( .A(core__abc_22172_new_n3474_), .B(core__abc_22172_new_n3494_), .Y(core__abc_22172_new_n3567_));
AND2X2 AND2X2_2505 ( .A(core__abc_22172_new_n3568_), .B(core__abc_22172_new_n3566_), .Y(core__abc_22172_new_n3569_));
AND2X2 AND2X2_2506 ( .A(core__abc_22172_new_n3570_), .B(core__abc_22172_new_n3565_), .Y(core__abc_22172_new_n3571_));
AND2X2 AND2X2_2507 ( .A(core__abc_22172_new_n2115_), .B(core__abc_22172_new_n2094_), .Y(core__abc_22172_new_n3576_));
AND2X2 AND2X2_2508 ( .A(core__abc_22172_new_n3575_), .B(core__abc_22172_new_n3576_), .Y(core__abc_22172_new_n3577_));
AND2X2 AND2X2_2509 ( .A(core__abc_22172_new_n2113_), .B(core__abc_22172_new_n2093_), .Y(core__abc_22172_new_n3578_));
AND2X2 AND2X2_251 ( .A(_abc_19873_new_n925_), .B(word2_reg_18_), .Y(_abc_19873_new_n1318_));
AND2X2 AND2X2_2510 ( .A(core__abc_22172_new_n2095_), .B(core__abc_22172_new_n2113_), .Y(core__abc_22172_new_n3579_));
AND2X2 AND2X2_2511 ( .A(core__abc_22172_new_n3511_), .B(core__abc_22172_new_n3579_), .Y(core__abc_22172_new_n3580_));
AND2X2 AND2X2_2512 ( .A(core__abc_22172_new_n3582_), .B(core__abc_22172_new_n3574_), .Y(core__abc_22172_new_n3583_));
AND2X2 AND2X2_2513 ( .A(core__abc_22172_new_n3584_), .B(core_v3_reg_33_), .Y(core__abc_22172_new_n3585_));
AND2X2 AND2X2_2514 ( .A(core__abc_22172_new_n3589_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n3590_));
AND2X2 AND2X2_2515 ( .A(core__abc_22172_new_n3590_), .B(core__abc_22172_new_n3588_), .Y(core__abc_22172_new_n3591_));
AND2X2 AND2X2_2516 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n3592_), .Y(core__abc_22172_new_n3593_));
AND2X2 AND2X2_2517 ( .A(core_v3_reg_6_), .B(core_mi_6_), .Y(core__abc_22172_new_n3594_));
AND2X2 AND2X2_2518 ( .A(core__abc_22172_new_n3595_), .B(core__abc_22172_new_n3596_), .Y(core__abc_22172_new_n3597_));
AND2X2 AND2X2_2519 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n3597_), .Y(core__abc_22172_new_n3598_));
AND2X2 AND2X2_252 ( .A(_abc_19873_new_n881_), .B(core_key_114_), .Y(_abc_19873_new_n1321_));
AND2X2 AND2X2_2520 ( .A(core__abc_22172_new_n3602_), .B(reset_n), .Y(core__abc_22172_new_n3603_));
AND2X2 AND2X2_2521 ( .A(core__abc_22172_new_n3601_), .B(core__abc_22172_new_n3603_), .Y(core__0v3_reg_63_0__6_));
AND2X2 AND2X2_2522 ( .A(core__abc_22172_new_n3606_), .B(core__abc_22172_new_n1944_), .Y(core__abc_22172_new_n3607_));
AND2X2 AND2X2_2523 ( .A(core__abc_22172_new_n3605_), .B(core__abc_22172_new_n1938_), .Y(core__abc_22172_new_n3608_));
AND2X2 AND2X2_2524 ( .A(core__abc_22172_new_n3613_), .B(core__abc_22172_new_n1401_), .Y(core__abc_22172_new_n3614_));
AND2X2 AND2X2_2525 ( .A(core__abc_22172_new_n3612_), .B(core__abc_22172_new_n1398_), .Y(core__abc_22172_new_n3615_));
AND2X2 AND2X2_2526 ( .A(core__abc_22172_new_n3616_), .B(core__abc_22172_new_n3611_), .Y(core__abc_22172_new_n3617_));
AND2X2 AND2X2_2527 ( .A(core__abc_22172_new_n3618_), .B(core_v3_reg_55_), .Y(core__abc_22172_new_n3619_));
AND2X2 AND2X2_2528 ( .A(core__abc_22172_new_n3622_), .B(core__abc_22172_new_n3623_), .Y(core__abc_22172_new_n3624_));
AND2X2 AND2X2_2529 ( .A(core__abc_22172_new_n3627_), .B(core__abc_22172_new_n3625_), .Y(core__abc_22172_new_n3628_));
AND2X2 AND2X2_253 ( .A(_abc_19873_new_n888_), .B(core_mi_18_), .Y(_abc_19873_new_n1322_));
AND2X2 AND2X2_2530 ( .A(core__abc_22172_new_n3626_), .B(core__abc_22172_new_n3624_), .Y(core__abc_22172_new_n3629_));
AND2X2 AND2X2_2531 ( .A(core__abc_22172_new_n3635_), .B(core__abc_22172_new_n2132_), .Y(core__abc_22172_new_n3636_));
AND2X2 AND2X2_2532 ( .A(core__abc_22172_new_n3634_), .B(core__abc_22172_new_n2129_), .Y(core__abc_22172_new_n3637_));
AND2X2 AND2X2_2533 ( .A(core__abc_22172_new_n3640_), .B(core__abc_22172_new_n3641_), .Y(core__abc_22172_new_n3642_));
AND2X2 AND2X2_2534 ( .A(core__abc_22172_new_n3645_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n3646_));
AND2X2 AND2X2_2535 ( .A(core__abc_22172_new_n3646_), .B(core__abc_22172_new_n3644_), .Y(core__abc_22172_new_n3647_));
AND2X2 AND2X2_2536 ( .A(core__abc_22172_new_n3214_), .B(core_key_71_), .Y(core__abc_22172_new_n3648_));
AND2X2 AND2X2_2537 ( .A(core_v3_reg_7_), .B(core_mi_7_), .Y(core__abc_22172_new_n3649_));
AND2X2 AND2X2_2538 ( .A(core__abc_22172_new_n3650_), .B(core__abc_22172_new_n3651_), .Y(core__abc_22172_new_n3652_));
AND2X2 AND2X2_2539 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n3652_), .Y(core__abc_22172_new_n3653_));
AND2X2 AND2X2_254 ( .A(_abc_19873_new_n928_), .B(core_key_50_), .Y(_abc_19873_new_n1324_));
AND2X2 AND2X2_2540 ( .A(core__abc_22172_new_n3657_), .B(reset_n), .Y(core__abc_22172_new_n3658_));
AND2X2 AND2X2_2541 ( .A(core__abc_22172_new_n3656_), .B(core__abc_22172_new_n3658_), .Y(core__0v3_reg_63_0__7_));
AND2X2 AND2X2_2542 ( .A(core__abc_22172_new_n3495_), .B(core__abc_22172_new_n3436_), .Y(core__abc_22172_new_n3660_));
AND2X2 AND2X2_2543 ( .A(core__abc_22172_new_n3624_), .B(core__abc_22172_new_n3566_), .Y(core__abc_22172_new_n3661_));
AND2X2 AND2X2_2544 ( .A(core__abc_22172_new_n3661_), .B(core__abc_22172_new_n3660_), .Y(core__abc_22172_new_n3662_));
AND2X2 AND2X2_2545 ( .A(core__abc_22172_new_n3662_), .B(core__abc_22172_new_n3438_), .Y(core__abc_22172_new_n3663_));
AND2X2 AND2X2_2546 ( .A(core__abc_22172_new_n3622_), .B(core__abc_22172_new_n3564_), .Y(core__abc_22172_new_n3665_));
AND2X2 AND2X2_2547 ( .A(core__abc_22172_new_n3495_), .B(core__abc_22172_new_n3434_), .Y(core__abc_22172_new_n3667_));
AND2X2 AND2X2_2548 ( .A(core__abc_22172_new_n3661_), .B(core__abc_22172_new_n3668_), .Y(core__abc_22172_new_n3669_));
AND2X2 AND2X2_2549 ( .A(core__abc_22172_new_n1921_), .B(core__abc_22172_new_n1938_), .Y(core__abc_22172_new_n3673_));
AND2X2 AND2X2_255 ( .A(_abc_19873_new_n916_), .B(core_key_82_), .Y(_abc_19873_new_n1325_));
AND2X2 AND2X2_2550 ( .A(core__abc_22172_new_n3542_), .B(core__abc_22172_new_n3673_), .Y(core__abc_22172_new_n3674_));
AND2X2 AND2X2_2551 ( .A(core__abc_22172_new_n3415_), .B(core__abc_22172_new_n3674_), .Y(core__abc_22172_new_n3675_));
AND2X2 AND2X2_2552 ( .A(core__abc_22172_new_n3541_), .B(core__abc_22172_new_n3673_), .Y(core__abc_22172_new_n3676_));
AND2X2 AND2X2_2553 ( .A(core__abc_22172_new_n1935_), .B(core__abc_22172_new_n1919_), .Y(core__abc_22172_new_n3677_));
AND2X2 AND2X2_2554 ( .A(core__abc_22172_new_n3416_), .B(core__abc_22172_new_n3674_), .Y(core__abc_22172_new_n3681_));
AND2X2 AND2X2_2555 ( .A(core__abc_22172_new_n3013_), .B(core__abc_22172_new_n3681_), .Y(core__abc_22172_new_n3682_));
AND2X2 AND2X2_2556 ( .A(core__abc_22172_new_n3683_), .B(core__abc_22172_new_n1955_), .Y(core__abc_22172_new_n3684_));
AND2X2 AND2X2_2557 ( .A(core__abc_22172_new_n3685_), .B(core__abc_22172_new_n1961_), .Y(core__abc_22172_new_n3686_));
AND2X2 AND2X2_2558 ( .A(core__abc_22172_new_n3690_), .B(core__abc_22172_new_n1418_), .Y(core__abc_22172_new_n3691_));
AND2X2 AND2X2_2559 ( .A(core__abc_22172_new_n3073_), .B(core__abc_22172_new_n1415_), .Y(core__abc_22172_new_n3692_));
AND2X2 AND2X2_256 ( .A(_abc_19873_new_n930_), .B(word0_reg_18_), .Y(_abc_19873_new_n1328_));
AND2X2 AND2X2_2560 ( .A(core__abc_22172_new_n3695_), .B(core__abc_22172_new_n3696_), .Y(core__abc_22172_new_n3697_));
AND2X2 AND2X2_2561 ( .A(core__abc_22172_new_n3688_), .B(core__abc_22172_new_n3698_), .Y(core__abc_22172_new_n3699_));
AND2X2 AND2X2_2562 ( .A(core__abc_22172_new_n3687_), .B(core__abc_22172_new_n3697_), .Y(core__abc_22172_new_n3700_));
AND2X2 AND2X2_2563 ( .A(core__abc_22172_new_n3672_), .B(core__abc_22172_new_n3701_), .Y(core__abc_22172_new_n3702_));
AND2X2 AND2X2_2564 ( .A(core__abc_22172_new_n3671_), .B(core__abc_22172_new_n3703_), .Y(core__abc_22172_new_n3704_));
AND2X2 AND2X2_2565 ( .A(core__abc_22172_new_n3707_), .B(core__abc_22172_new_n2146_), .Y(core__abc_22172_new_n3709_));
AND2X2 AND2X2_2566 ( .A(core__abc_22172_new_n3710_), .B(core__abc_22172_new_n3708_), .Y(core__abc_22172_new_n3711_));
AND2X2 AND2X2_2567 ( .A(core__abc_22172_new_n3712_), .B(core_v3_reg_35_), .Y(core__abc_22172_new_n3713_));
AND2X2 AND2X2_2568 ( .A(core__abc_22172_new_n3714_), .B(core__abc_22172_new_n3715_), .Y(core__abc_22172_new_n3716_));
AND2X2 AND2X2_2569 ( .A(core__abc_22172_new_n3719_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n3720_));
AND2X2 AND2X2_257 ( .A(_abc_19873_new_n907_), .B(word1_reg_18_), .Y(_abc_19873_new_n1329_));
AND2X2 AND2X2_2570 ( .A(core__abc_22172_new_n3720_), .B(core__abc_22172_new_n3718_), .Y(core__abc_22172_new_n3721_));
AND2X2 AND2X2_2571 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n3722_), .Y(core__abc_22172_new_n3723_));
AND2X2 AND2X2_2572 ( .A(core_v3_reg_8_), .B(core_mi_8_), .Y(core__abc_22172_new_n3724_));
AND2X2 AND2X2_2573 ( .A(core__abc_22172_new_n3725_), .B(core__abc_22172_new_n3726_), .Y(core__abc_22172_new_n3727_));
AND2X2 AND2X2_2574 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n3727_), .Y(core__abc_22172_new_n3728_));
AND2X2 AND2X2_2575 ( .A(core__abc_22172_new_n3732_), .B(reset_n), .Y(core__abc_22172_new_n3733_));
AND2X2 AND2X2_2576 ( .A(core__abc_22172_new_n3731_), .B(core__abc_22172_new_n3733_), .Y(core__0v3_reg_63_0__8_));
AND2X2 AND2X2_2577 ( .A(core__abc_22172_new_n3737_), .B(core__abc_22172_new_n1954_), .Y(core__abc_22172_new_n3738_));
AND2X2 AND2X2_2578 ( .A(core__abc_22172_new_n3738_), .B(core__abc_22172_new_n1978_), .Y(core__abc_22172_new_n3739_));
AND2X2 AND2X2_2579 ( .A(core__abc_22172_new_n3740_), .B(core__abc_22172_new_n3741_), .Y(core__abc_22172_new_n3742_));
AND2X2 AND2X2_258 ( .A(_abc_19873_new_n919_), .B(core_mi_50_), .Y(_abc_19873_new_n1331_));
AND2X2 AND2X2_2580 ( .A(core__abc_22172_new_n3745_), .B(core__abc_22172_new_n1435_), .Y(core__abc_22172_new_n3746_));
AND2X2 AND2X2_2581 ( .A(core__abc_22172_new_n3744_), .B(core__abc_22172_new_n1432_), .Y(core__abc_22172_new_n3747_));
AND2X2 AND2X2_2582 ( .A(core__abc_22172_new_n3748_), .B(core__abc_22172_new_n3743_), .Y(core__abc_22172_new_n3749_));
AND2X2 AND2X2_2583 ( .A(core__abc_22172_new_n3750_), .B(core_v3_reg_57_), .Y(core__abc_22172_new_n3751_));
AND2X2 AND2X2_2584 ( .A(core__abc_22172_new_n3742_), .B(core__abc_22172_new_n3753_), .Y(core__abc_22172_new_n3754_));
AND2X2 AND2X2_2585 ( .A(core__abc_22172_new_n3755_), .B(core__abc_22172_new_n3756_), .Y(core__abc_22172_new_n3757_));
AND2X2 AND2X2_2586 ( .A(core__abc_22172_new_n3758_), .B(core__abc_22172_new_n3736_), .Y(core__abc_22172_new_n3759_));
AND2X2 AND2X2_2587 ( .A(core__abc_22172_new_n3735_), .B(core__abc_22172_new_n3759_), .Y(core__abc_22172_new_n3760_));
AND2X2 AND2X2_2588 ( .A(core__abc_22172_new_n3757_), .B(core__abc_22172_new_n3699_), .Y(core__abc_22172_new_n3762_));
AND2X2 AND2X2_2589 ( .A(core__abc_22172_new_n3757_), .B(core__abc_22172_new_n3703_), .Y(core__abc_22172_new_n3764_));
AND2X2 AND2X2_259 ( .A(_abc_19873_new_n1335_), .B(_abc_19873_new_n937_), .Y(\read_data[18] ));
AND2X2 AND2X2_2590 ( .A(core__abc_22172_new_n3671_), .B(core__abc_22172_new_n3764_), .Y(core__abc_22172_new_n3765_));
AND2X2 AND2X2_2591 ( .A(core__abc_22172_new_n3766_), .B(core__abc_22172_new_n3763_), .Y(core__abc_22172_new_n3767_));
AND2X2 AND2X2_2592 ( .A(core__abc_22172_new_n3761_), .B(core__abc_22172_new_n3767_), .Y(core__abc_22172_new_n3768_));
AND2X2 AND2X2_2593 ( .A(core__abc_22172_new_n2129_), .B(core__abc_22172_new_n2146_), .Y(core__abc_22172_new_n3770_));
AND2X2 AND2X2_2594 ( .A(core__abc_22172_new_n3579_), .B(core__abc_22172_new_n3770_), .Y(core__abc_22172_new_n3771_));
AND2X2 AND2X2_2595 ( .A(core__abc_22172_new_n3511_), .B(core__abc_22172_new_n3771_), .Y(core__abc_22172_new_n3772_));
AND2X2 AND2X2_2596 ( .A(core__abc_22172_new_n3633_), .B(core__abc_22172_new_n3770_), .Y(core__abc_22172_new_n3773_));
AND2X2 AND2X2_2597 ( .A(core__abc_22172_new_n2143_), .B(core__abc_22172_new_n2127_), .Y(core__abc_22172_new_n3774_));
AND2X2 AND2X2_2598 ( .A(core__abc_22172_new_n3778_), .B(core__abc_22172_new_n2166_), .Y(core__abc_22172_new_n3779_));
AND2X2 AND2X2_2599 ( .A(core__abc_22172_new_n3777_), .B(core__abc_22172_new_n2163_), .Y(core__abc_22172_new_n3780_));
AND2X2 AND2X2_26 ( .A(_abc_19873_new_n891_), .B(\addr[5] ), .Y(_abc_19873_new_n905_));
AND2X2 AND2X2_260 ( .A(_abc_19873_new_n881_), .B(core_key_115_), .Y(_abc_19873_new_n1337_));
AND2X2 AND2X2_2600 ( .A(core__abc_22172_new_n3783_), .B(core__abc_22172_new_n3784_), .Y(core__abc_22172_new_n3785_));
AND2X2 AND2X2_2601 ( .A(core__abc_22172_new_n3789_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n3790_));
AND2X2 AND2X2_2602 ( .A(core__abc_22172_new_n3790_), .B(core__abc_22172_new_n3787_), .Y(core__abc_22172_new_n3791_));
AND2X2 AND2X2_2603 ( .A(core__abc_22172_new_n3214_), .B(core_key_73_), .Y(core__abc_22172_new_n3792_));
AND2X2 AND2X2_2604 ( .A(core_v3_reg_9_), .B(core_mi_9_), .Y(core__abc_22172_new_n3793_));
AND2X2 AND2X2_2605 ( .A(core__abc_22172_new_n3794_), .B(core__abc_22172_new_n3795_), .Y(core__abc_22172_new_n3796_));
AND2X2 AND2X2_2606 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n3796_), .Y(core__abc_22172_new_n3797_));
AND2X2 AND2X2_2607 ( .A(core__abc_22172_new_n3801_), .B(reset_n), .Y(core__abc_22172_new_n3802_));
AND2X2 AND2X2_2608 ( .A(core__abc_22172_new_n3800_), .B(core__abc_22172_new_n3802_), .Y(core__0v3_reg_63_0__9_));
AND2X2 AND2X2_2609 ( .A(core__abc_22172_new_n3766_), .B(core__abc_22172_new_n3805_), .Y(core__abc_22172_new_n3806_));
AND2X2 AND2X2_261 ( .A(_abc_19873_new_n888_), .B(core_mi_19_), .Y(_abc_19873_new_n1338_));
AND2X2 AND2X2_2610 ( .A(core__abc_22172_new_n1955_), .B(core__abc_22172_new_n1972_), .Y(core__abc_22172_new_n3808_));
AND2X2 AND2X2_2611 ( .A(core__abc_22172_new_n3683_), .B(core__abc_22172_new_n3808_), .Y(core__abc_22172_new_n3809_));
AND2X2 AND2X2_2612 ( .A(core__abc_22172_new_n1954_), .B(core__abc_22172_new_n1971_), .Y(core__abc_22172_new_n3811_));
AND2X2 AND2X2_2613 ( .A(core__abc_22172_new_n3814_), .B(core__abc_22172_new_n1989_), .Y(core__abc_22172_new_n3815_));
AND2X2 AND2X2_2614 ( .A(core__abc_22172_new_n3816_), .B(core__abc_22172_new_n1995_), .Y(core__abc_22172_new_n3817_));
AND2X2 AND2X2_2615 ( .A(core__abc_22172_new_n3073_), .B(core__abc_22172_new_n3077_), .Y(core__abc_22172_new_n3820_));
AND2X2 AND2X2_2616 ( .A(core__abc_22172_new_n3821_), .B(core__abc_22172_new_n3084_), .Y(core__abc_22172_new_n3822_));
AND2X2 AND2X2_2617 ( .A(core__abc_22172_new_n3822_), .B(core__abc_22172_new_n1452_), .Y(core__abc_22172_new_n3823_));
AND2X2 AND2X2_2618 ( .A(core__abc_22172_new_n3828_), .B(core__abc_22172_new_n3829_), .Y(core__abc_22172_new_n3830_));
AND2X2 AND2X2_2619 ( .A(core__abc_22172_new_n3818_), .B(core__abc_22172_new_n3830_), .Y(core__abc_22172_new_n3831_));
AND2X2 AND2X2_262 ( .A(_abc_19873_new_n916_), .B(core_key_83_), .Y(_abc_19873_new_n1340_));
AND2X2 AND2X2_2620 ( .A(core__abc_22172_new_n3832_), .B(core__abc_22172_new_n3833_), .Y(core__abc_22172_new_n3834_));
AND2X2 AND2X2_2621 ( .A(core__abc_22172_new_n3807_), .B(core__abc_22172_new_n3836_), .Y(core__abc_22172_new_n3837_));
AND2X2 AND2X2_2622 ( .A(core__abc_22172_new_n3806_), .B(core__abc_22172_new_n3835_), .Y(core__abc_22172_new_n3838_));
AND2X2 AND2X2_2623 ( .A(core__abc_22172_new_n3842_), .B(core__abc_22172_new_n2183_), .Y(core__abc_22172_new_n3843_));
AND2X2 AND2X2_2624 ( .A(core__abc_22172_new_n3841_), .B(core__abc_22172_new_n2181_), .Y(core__abc_22172_new_n3844_));
AND2X2 AND2X2_2625 ( .A(core__abc_22172_new_n3845_), .B(core_v3_reg_37_), .Y(core__abc_22172_new_n3847_));
AND2X2 AND2X2_2626 ( .A(core__abc_22172_new_n3848_), .B(core__abc_22172_new_n3846_), .Y(core__abc_22172_new_n3849_));
AND2X2 AND2X2_2627 ( .A(core__abc_22172_new_n3852_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n3853_));
AND2X2 AND2X2_2628 ( .A(core__abc_22172_new_n3853_), .B(core__abc_22172_new_n3851_), .Y(core__abc_22172_new_n3854_));
AND2X2 AND2X2_2629 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n3855_), .Y(core__abc_22172_new_n3856_));
AND2X2 AND2X2_263 ( .A(_abc_19873_new_n925_), .B(word2_reg_19_), .Y(_abc_19873_new_n1343_));
AND2X2 AND2X2_2630 ( .A(core_v3_reg_10_), .B(core_mi_10_), .Y(core__abc_22172_new_n3857_));
AND2X2 AND2X2_2631 ( .A(core__abc_22172_new_n3858_), .B(core__abc_22172_new_n3859_), .Y(core__abc_22172_new_n3860_));
AND2X2 AND2X2_2632 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n3860_), .Y(core__abc_22172_new_n3861_));
AND2X2 AND2X2_2633 ( .A(core__abc_22172_new_n3865_), .B(reset_n), .Y(core__abc_22172_new_n3866_));
AND2X2 AND2X2_2634 ( .A(core__abc_22172_new_n3864_), .B(core__abc_22172_new_n3866_), .Y(core__0v3_reg_63_0__10_));
AND2X2 AND2X2_2635 ( .A(core__abc_22172_new_n3871_), .B(core__abc_22172_new_n2012_), .Y(core__abc_22172_new_n3872_));
AND2X2 AND2X2_2636 ( .A(core__abc_22172_new_n3870_), .B(core__abc_22172_new_n2006_), .Y(core__abc_22172_new_n3873_));
AND2X2 AND2X2_2637 ( .A(core__abc_22172_new_n3824_), .B(core__abc_22172_new_n1447_), .Y(core__abc_22172_new_n3876_));
AND2X2 AND2X2_2638 ( .A(core__abc_22172_new_n3876_), .B(core__abc_22172_new_n1469_), .Y(core__abc_22172_new_n3877_));
AND2X2 AND2X2_2639 ( .A(core__abc_22172_new_n3878_), .B(core__abc_22172_new_n3879_), .Y(core__abc_22172_new_n3880_));
AND2X2 AND2X2_264 ( .A(_abc_19873_new_n907_), .B(word1_reg_19_), .Y(_abc_19873_new_n1344_));
AND2X2 AND2X2_2640 ( .A(core__abc_22172_new_n3881_), .B(core_v3_reg_59_), .Y(core__abc_22172_new_n3882_));
AND2X2 AND2X2_2641 ( .A(core__abc_22172_new_n3883_), .B(core__abc_22172_new_n3884_), .Y(core__abc_22172_new_n3885_));
AND2X2 AND2X2_2642 ( .A(core__abc_22172_new_n3887_), .B(core__abc_22172_new_n3888_), .Y(core__abc_22172_new_n3889_));
AND2X2 AND2X2_2643 ( .A(core__abc_22172_new_n3869_), .B(core__abc_22172_new_n3890_), .Y(core__abc_22172_new_n3891_));
AND2X2 AND2X2_2644 ( .A(core__abc_22172_new_n3868_), .B(core__abc_22172_new_n3889_), .Y(core__abc_22172_new_n3892_));
AND2X2 AND2X2_2645 ( .A(core__abc_22172_new_n2163_), .B(core__abc_22172_new_n2181_), .Y(core__abc_22172_new_n3896_));
AND2X2 AND2X2_2646 ( .A(core__abc_22172_new_n3777_), .B(core__abc_22172_new_n3896_), .Y(core__abc_22172_new_n3897_));
AND2X2 AND2X2_2647 ( .A(core__abc_22172_new_n2181_), .B(core__abc_22172_new_n2161_), .Y(core__abc_22172_new_n3898_));
AND2X2 AND2X2_2648 ( .A(core__abc_22172_new_n3900_), .B(core__abc_22172_new_n2197_), .Y(core__abc_22172_new_n3901_));
AND2X2 AND2X2_2649 ( .A(core__abc_22172_new_n3902_), .B(core__abc_22172_new_n2200_), .Y(core__abc_22172_new_n3903_));
AND2X2 AND2X2_265 ( .A(_abc_19873_new_n912_), .B(word3_reg_19_), .Y(_abc_19873_new_n1345_));
AND2X2 AND2X2_2650 ( .A(core__abc_22172_new_n3906_), .B(core__abc_22172_new_n3907_), .Y(core__abc_22172_new_n3908_));
AND2X2 AND2X2_2651 ( .A(core__abc_22172_new_n3911_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n3912_));
AND2X2 AND2X2_2652 ( .A(core__abc_22172_new_n3912_), .B(core__abc_22172_new_n3910_), .Y(core__abc_22172_new_n3913_));
AND2X2 AND2X2_2653 ( .A(core__abc_22172_new_n3214_), .B(core_key_75_), .Y(core__abc_22172_new_n3914_));
AND2X2 AND2X2_2654 ( .A(core_v3_reg_11_), .B(core_mi_11_), .Y(core__abc_22172_new_n3915_));
AND2X2 AND2X2_2655 ( .A(core__abc_22172_new_n3916_), .B(core__abc_22172_new_n3917_), .Y(core__abc_22172_new_n3918_));
AND2X2 AND2X2_2656 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n3918_), .Y(core__abc_22172_new_n3919_));
AND2X2 AND2X2_2657 ( .A(core__abc_22172_new_n3923_), .B(reset_n), .Y(core__abc_22172_new_n3924_));
AND2X2 AND2X2_2658 ( .A(core__abc_22172_new_n3922_), .B(core__abc_22172_new_n3924_), .Y(core__0v3_reg_63_0__11_));
AND2X2 AND2X2_2659 ( .A(core__abc_22172_new_n3889_), .B(core__abc_22172_new_n3836_), .Y(core__abc_22172_new_n3926_));
AND2X2 AND2X2_266 ( .A(_abc_19873_new_n919_), .B(core_mi_51_), .Y(_abc_19873_new_n1348_));
AND2X2 AND2X2_2660 ( .A(core__abc_22172_new_n3926_), .B(core__abc_22172_new_n3804_), .Y(core__abc_22172_new_n3927_));
AND2X2 AND2X2_2661 ( .A(core__abc_22172_new_n3887_), .B(core__abc_22172_new_n3834_), .Y(core__abc_22172_new_n3929_));
AND2X2 AND2X2_2662 ( .A(core__abc_22172_new_n3926_), .B(core__abc_22172_new_n3764_), .Y(core__abc_22172_new_n3932_));
AND2X2 AND2X2_2663 ( .A(core__abc_22172_new_n3671_), .B(core__abc_22172_new_n3932_), .Y(core__abc_22172_new_n3933_));
AND2X2 AND2X2_2664 ( .A(core__abc_22172_new_n1989_), .B(core__abc_22172_new_n2006_), .Y(core__abc_22172_new_n3935_));
AND2X2 AND2X2_2665 ( .A(core__abc_22172_new_n3813_), .B(core__abc_22172_new_n3935_), .Y(core__abc_22172_new_n3936_));
AND2X2 AND2X2_2666 ( .A(core__abc_22172_new_n2003_), .B(core__abc_22172_new_n1987_), .Y(core__abc_22172_new_n3937_));
AND2X2 AND2X2_2667 ( .A(core__abc_22172_new_n3808_), .B(core__abc_22172_new_n3935_), .Y(core__abc_22172_new_n3940_));
AND2X2 AND2X2_2668 ( .A(core__abc_22172_new_n3683_), .B(core__abc_22172_new_n3940_), .Y(core__abc_22172_new_n3941_));
AND2X2 AND2X2_2669 ( .A(core__abc_22172_new_n3942_), .B(core__abc_22172_new_n2023_), .Y(core__abc_22172_new_n3943_));
AND2X2 AND2X2_267 ( .A(_abc_19873_new_n930_), .B(word0_reg_19_), .Y(_abc_19873_new_n1349_));
AND2X2 AND2X2_2670 ( .A(core__abc_22172_new_n3944_), .B(core__abc_22172_new_n2029_), .Y(core__abc_22172_new_n3945_));
AND2X2 AND2X2_2671 ( .A(core__abc_22172_new_n3073_), .B(core__abc_22172_new_n3079_), .Y(core__abc_22172_new_n3948_));
AND2X2 AND2X2_2672 ( .A(core__abc_22172_new_n3949_), .B(core__abc_22172_new_n1483_), .Y(core__abc_22172_new_n3950_));
AND2X2 AND2X2_2673 ( .A(core__abc_22172_new_n3951_), .B(core__abc_22172_new_n1486_), .Y(core__abc_22172_new_n3952_));
AND2X2 AND2X2_2674 ( .A(core__abc_22172_new_n3955_), .B(core__abc_22172_new_n3956_), .Y(core__abc_22172_new_n3957_));
AND2X2 AND2X2_2675 ( .A(core__abc_22172_new_n3946_), .B(core__abc_22172_new_n3957_), .Y(core__abc_22172_new_n3958_));
AND2X2 AND2X2_2676 ( .A(core__abc_22172_new_n3959_), .B(core__abc_22172_new_n3960_), .Y(core__abc_22172_new_n3961_));
AND2X2 AND2X2_2677 ( .A(core__abc_22172_new_n3934_), .B(core__abc_22172_new_n3963_), .Y(core__abc_22172_new_n3964_));
AND2X2 AND2X2_2678 ( .A(core__abc_22172_new_n3965_), .B(core__abc_22172_new_n3966_), .Y(core__abc_22172_new_n3967_));
AND2X2 AND2X2_2679 ( .A(core__abc_22172_new_n3969_), .B(core__abc_22172_new_n2217_), .Y(core__abc_22172_new_n3970_));
AND2X2 AND2X2_268 ( .A(_abc_19873_new_n928_), .B(core_key_51_), .Y(_abc_19873_new_n1351_));
AND2X2 AND2X2_2680 ( .A(core__abc_22172_new_n3968_), .B(core__abc_22172_new_n2214_), .Y(core__abc_22172_new_n3971_));
AND2X2 AND2X2_2681 ( .A(core__abc_22172_new_n3972_), .B(core_v3_reg_39_), .Y(core__abc_22172_new_n3973_));
AND2X2 AND2X2_2682 ( .A(core__abc_22172_new_n3979_), .B(core__abc_22172_new_n3974_), .Y(core__abc_22172_new_n3980_));
AND2X2 AND2X2_2683 ( .A(core__abc_22172_new_n3981_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n3982_));
AND2X2 AND2X2_2684 ( .A(core__abc_22172_new_n3982_), .B(core__abc_22172_new_n3977_), .Y(core__abc_22172_new_n3983_));
AND2X2 AND2X2_2685 ( .A(core__abc_22172_new_n3214_), .B(core_key_76_), .Y(core__abc_22172_new_n3984_));
AND2X2 AND2X2_2686 ( .A(core_v3_reg_12_), .B(core_mi_12_), .Y(core__abc_22172_new_n3985_));
AND2X2 AND2X2_2687 ( .A(core__abc_22172_new_n3986_), .B(core__abc_22172_new_n3987_), .Y(core__abc_22172_new_n3988_));
AND2X2 AND2X2_2688 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n3988_), .Y(core__abc_22172_new_n3989_));
AND2X2 AND2X2_2689 ( .A(core__abc_22172_new_n3993_), .B(reset_n), .Y(core__abc_22172_new_n3994_));
AND2X2 AND2X2_269 ( .A(_abc_19873_new_n901_), .B(core_key_19_), .Y(_abc_19873_new_n1352_));
AND2X2 AND2X2_2690 ( .A(core__abc_22172_new_n3992_), .B(core__abc_22172_new_n3994_), .Y(core__0v3_reg_63_0__12_));
AND2X2 AND2X2_2691 ( .A(core__abc_22172_new_n3998_), .B(core__abc_22172_new_n2046_), .Y(core__abc_22172_new_n3999_));
AND2X2 AND2X2_2692 ( .A(core__abc_22172_new_n3997_), .B(core__abc_22172_new_n2040_), .Y(core__abc_22172_new_n4000_));
AND2X2 AND2X2_2693 ( .A(core__abc_22172_new_n4005_), .B(core__abc_22172_new_n1503_), .Y(core__abc_22172_new_n4006_));
AND2X2 AND2X2_2694 ( .A(core__abc_22172_new_n4004_), .B(core__abc_22172_new_n1500_), .Y(core__abc_22172_new_n4007_));
AND2X2 AND2X2_2695 ( .A(core__abc_22172_new_n4008_), .B(core__abc_22172_new_n4003_), .Y(core__abc_22172_new_n4009_));
AND2X2 AND2X2_2696 ( .A(core__abc_22172_new_n4010_), .B(core_v3_reg_61_), .Y(core__abc_22172_new_n4011_));
AND2X2 AND2X2_2697 ( .A(core__abc_22172_new_n4014_), .B(core__abc_22172_new_n4015_), .Y(core__abc_22172_new_n4016_));
AND2X2 AND2X2_2698 ( .A(core__abc_22172_new_n4017_), .B(core__abc_22172_new_n3996_), .Y(core__abc_22172_new_n4018_));
AND2X2 AND2X2_2699 ( .A(core__abc_22172_new_n3965_), .B(core__abc_22172_new_n4018_), .Y(core__abc_22172_new_n4019_));
AND2X2 AND2X2_27 ( .A(_abc_19873_new_n872_), .B(_abc_19873_new_n905_), .Y(_abc_19873_new_n906_));
AND2X2 AND2X2_270 ( .A(_abc_19873_new_n1356_), .B(_abc_19873_new_n937_), .Y(\read_data[19] ));
AND2X2 AND2X2_2700 ( .A(core__abc_22172_new_n4016_), .B(core__abc_22172_new_n3961_), .Y(core__abc_22172_new_n4021_));
AND2X2 AND2X2_2701 ( .A(core__abc_22172_new_n4016_), .B(core__abc_22172_new_n3963_), .Y(core__abc_22172_new_n4023_));
AND2X2 AND2X2_2702 ( .A(core__abc_22172_new_n3934_), .B(core__abc_22172_new_n4023_), .Y(core__abc_22172_new_n4024_));
AND2X2 AND2X2_2703 ( .A(core__abc_22172_new_n4025_), .B(core__abc_22172_new_n4022_), .Y(core__abc_22172_new_n4026_));
AND2X2 AND2X2_2704 ( .A(core__abc_22172_new_n4020_), .B(core__abc_22172_new_n4026_), .Y(core__abc_22172_new_n4027_));
AND2X2 AND2X2_2705 ( .A(core__abc_22172_new_n2211_), .B(core__abc_22172_new_n2195_), .Y(core__abc_22172_new_n4029_));
AND2X2 AND2X2_2706 ( .A(core__abc_22172_new_n2197_), .B(core__abc_22172_new_n2214_), .Y(core__abc_22172_new_n4031_));
AND2X2 AND2X2_2707 ( .A(core__abc_22172_new_n3899_), .B(core__abc_22172_new_n4031_), .Y(core__abc_22172_new_n4032_));
AND2X2 AND2X2_2708 ( .A(core__abc_22172_new_n3897_), .B(core__abc_22172_new_n4031_), .Y(core__abc_22172_new_n4034_));
AND2X2 AND2X2_2709 ( .A(core__abc_22172_new_n4035_), .B(core__abc_22172_new_n2231_), .Y(core__abc_22172_new_n4036_));
AND2X2 AND2X2_271 ( .A(_abc_19873_new_n912_), .B(word3_reg_20_), .Y(_abc_19873_new_n1358_));
AND2X2 AND2X2_2710 ( .A(core__abc_22172_new_n4037_), .B(core__abc_22172_new_n2234_), .Y(core__abc_22172_new_n4038_));
AND2X2 AND2X2_2711 ( .A(core__abc_22172_new_n4041_), .B(core__abc_22172_new_n4043_), .Y(core__abc_22172_new_n4044_));
AND2X2 AND2X2_2712 ( .A(core__abc_22172_new_n4047_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n4048_));
AND2X2 AND2X2_2713 ( .A(core__abc_22172_new_n4048_), .B(core__abc_22172_new_n4046_), .Y(core__abc_22172_new_n4049_));
AND2X2 AND2X2_2714 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n4050_), .Y(core__abc_22172_new_n4051_));
AND2X2 AND2X2_2715 ( .A(core_v3_reg_13_), .B(core_mi_13_), .Y(core__abc_22172_new_n4052_));
AND2X2 AND2X2_2716 ( .A(core__abc_22172_new_n4053_), .B(core__abc_22172_new_n4054_), .Y(core__abc_22172_new_n4055_));
AND2X2 AND2X2_2717 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n4055_), .Y(core__abc_22172_new_n4056_));
AND2X2 AND2X2_2718 ( .A(core__abc_22172_new_n4060_), .B(reset_n), .Y(core__abc_22172_new_n4061_));
AND2X2 AND2X2_2719 ( .A(core__abc_22172_new_n4059_), .B(core__abc_22172_new_n4061_), .Y(core__0v3_reg_63_0__13_));
AND2X2 AND2X2_272 ( .A(_abc_19873_new_n901_), .B(core_key_20_), .Y(_abc_19873_new_n1359_));
AND2X2 AND2X2_2720 ( .A(core__abc_22172_new_n4025_), .B(core__abc_22172_new_n4065_), .Y(core__abc_22172_new_n4066_));
AND2X2 AND2X2_2721 ( .A(core__abc_22172_new_n2022_), .B(core__abc_22172_new_n2039_), .Y(core__abc_22172_new_n4069_));
AND2X2 AND2X2_2722 ( .A(core__abc_22172_new_n2023_), .B(core__abc_22172_new_n2040_), .Y(core__abc_22172_new_n4072_));
AND2X2 AND2X2_2723 ( .A(core__abc_22172_new_n3942_), .B(core__abc_22172_new_n4072_), .Y(core__abc_22172_new_n4073_));
AND2X2 AND2X2_2724 ( .A(core__abc_22172_new_n4074_), .B(core__abc_22172_new_n2057_), .Y(core__abc_22172_new_n4075_));
AND2X2 AND2X2_2725 ( .A(core__abc_22172_new_n4076_), .B(core__abc_22172_new_n2063_), .Y(core__abc_22172_new_n4077_));
AND2X2 AND2X2_2726 ( .A(core__abc_22172_new_n3949_), .B(core__abc_22172_new_n3075_), .Y(core__abc_22172_new_n4080_));
AND2X2 AND2X2_2727 ( .A(core__abc_22172_new_n4082_), .B(core__abc_22172_new_n1520_), .Y(core__abc_22172_new_n4083_));
AND2X2 AND2X2_2728 ( .A(core__abc_22172_new_n4081_), .B(core__abc_22172_new_n1517_), .Y(core__abc_22172_new_n4084_));
AND2X2 AND2X2_2729 ( .A(core__abc_22172_new_n4087_), .B(core__abc_22172_new_n4088_), .Y(core__abc_22172_new_n4089_));
AND2X2 AND2X2_273 ( .A(_abc_19873_new_n925_), .B(word2_reg_20_), .Y(_abc_19873_new_n1360_));
AND2X2 AND2X2_2730 ( .A(core__abc_22172_new_n4078_), .B(core__abc_22172_new_n4089_), .Y(core__abc_22172_new_n4090_));
AND2X2 AND2X2_2731 ( .A(core__abc_22172_new_n4091_), .B(core__abc_22172_new_n4092_), .Y(core__abc_22172_new_n4093_));
AND2X2 AND2X2_2732 ( .A(core__abc_22172_new_n4067_), .B(core__abc_22172_new_n4093_), .Y(core__abc_22172_new_n4094_));
AND2X2 AND2X2_2733 ( .A(core__abc_22172_new_n4066_), .B(core__abc_22172_new_n4095_), .Y(core__abc_22172_new_n4096_));
AND2X2 AND2X2_2734 ( .A(core__abc_22172_new_n4100_), .B(core__abc_22172_new_n2251_), .Y(core__abc_22172_new_n4101_));
AND2X2 AND2X2_2735 ( .A(core__abc_22172_new_n4099_), .B(core__abc_22172_new_n2248_), .Y(core__abc_22172_new_n4102_));
AND2X2 AND2X2_2736 ( .A(core__abc_22172_new_n4104_), .B(core_v3_reg_41_), .Y(core__abc_22172_new_n4105_));
AND2X2 AND2X2_2737 ( .A(core__abc_22172_new_n4103_), .B(core__abc_22172_new_n4106_), .Y(core__abc_22172_new_n4107_));
AND2X2 AND2X2_2738 ( .A(core__abc_22172_new_n4111_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n4112_));
AND2X2 AND2X2_2739 ( .A(core__abc_22172_new_n4112_), .B(core__abc_22172_new_n4110_), .Y(core__abc_22172_new_n4113_));
AND2X2 AND2X2_274 ( .A(_abc_19873_new_n881_), .B(core_key_116_), .Y(_abc_19873_new_n1363_));
AND2X2 AND2X2_2740 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n4114_), .Y(core__abc_22172_new_n4115_));
AND2X2 AND2X2_2741 ( .A(core_v3_reg_14_), .B(core_mi_14_), .Y(core__abc_22172_new_n4116_));
AND2X2 AND2X2_2742 ( .A(core__abc_22172_new_n4117_), .B(core__abc_22172_new_n4118_), .Y(core__abc_22172_new_n4119_));
AND2X2 AND2X2_2743 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n4119_), .Y(core__abc_22172_new_n4120_));
AND2X2 AND2X2_2744 ( .A(core__abc_22172_new_n4124_), .B(reset_n), .Y(core__abc_22172_new_n4125_));
AND2X2 AND2X2_2745 ( .A(core__abc_22172_new_n4123_), .B(core__abc_22172_new_n4125_), .Y(core__0v3_reg_63_0__14_));
AND2X2 AND2X2_2746 ( .A(core__abc_22172_new_n4130_), .B(core__abc_22172_new_n2074_), .Y(core__abc_22172_new_n4132_));
AND2X2 AND2X2_2747 ( .A(core__abc_22172_new_n4133_), .B(core__abc_22172_new_n4131_), .Y(core__abc_22172_new_n4134_));
AND2X2 AND2X2_2748 ( .A(core__abc_22172_new_n4136_), .B(core__abc_22172_new_n1537_), .Y(core__abc_22172_new_n4137_));
AND2X2 AND2X2_2749 ( .A(core__abc_22172_new_n4135_), .B(core__abc_22172_new_n1534_), .Y(core__abc_22172_new_n4138_));
AND2X2 AND2X2_275 ( .A(_abc_19873_new_n888_), .B(core_mi_20_), .Y(_abc_19873_new_n1364_));
AND2X2 AND2X2_2750 ( .A(core__abc_22172_new_n4139_), .B(core_v3_reg_63_), .Y(core__abc_22172_new_n4140_));
AND2X2 AND2X2_2751 ( .A(core__abc_22172_new_n4141_), .B(core__abc_22172_new_n4142_), .Y(core__abc_22172_new_n4143_));
AND2X2 AND2X2_2752 ( .A(core__abc_22172_new_n4148_), .B(core__abc_22172_new_n4145_), .Y(core__abc_22172_new_n4149_));
AND2X2 AND2X2_2753 ( .A(core__abc_22172_new_n4129_), .B(core__abc_22172_new_n4150_), .Y(core__abc_22172_new_n4151_));
AND2X2 AND2X2_2754 ( .A(core__abc_22172_new_n4128_), .B(core__abc_22172_new_n4149_), .Y(core__abc_22172_new_n4152_));
AND2X2 AND2X2_2755 ( .A(core__abc_22172_new_n2231_), .B(core__abc_22172_new_n2248_), .Y(core__abc_22172_new_n4156_));
AND2X2 AND2X2_2756 ( .A(core__abc_22172_new_n4035_), .B(core__abc_22172_new_n4156_), .Y(core__abc_22172_new_n4157_));
AND2X2 AND2X2_2757 ( .A(core__abc_22172_new_n2248_), .B(core__abc_22172_new_n2229_), .Y(core__abc_22172_new_n4158_));
AND2X2 AND2X2_2758 ( .A(core__abc_22172_new_n4161_), .B(core__abc_22172_new_n2268_), .Y(core__abc_22172_new_n4162_));
AND2X2 AND2X2_2759 ( .A(core__abc_22172_new_n4160_), .B(core__abc_22172_new_n2265_), .Y(core__abc_22172_new_n4163_));
AND2X2 AND2X2_276 ( .A(_abc_19873_new_n928_), .B(core_key_52_), .Y(_abc_19873_new_n1366_));
AND2X2 AND2X2_2760 ( .A(core__abc_22172_new_n4166_), .B(core__abc_22172_new_n4167_), .Y(core__abc_22172_new_n4168_));
AND2X2 AND2X2_2761 ( .A(core__abc_22172_new_n4171_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n4172_));
AND2X2 AND2X2_2762 ( .A(core__abc_22172_new_n4172_), .B(core__abc_22172_new_n4170_), .Y(core__abc_22172_new_n4173_));
AND2X2 AND2X2_2763 ( .A(core__abc_22172_new_n3214_), .B(core_key_79_), .Y(core__abc_22172_new_n4174_));
AND2X2 AND2X2_2764 ( .A(core_v3_reg_15_), .B(core_mi_15_), .Y(core__abc_22172_new_n4175_));
AND2X2 AND2X2_2765 ( .A(core__abc_22172_new_n4176_), .B(core__abc_22172_new_n4177_), .Y(core__abc_22172_new_n4178_));
AND2X2 AND2X2_2766 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n4178_), .Y(core__abc_22172_new_n4179_));
AND2X2 AND2X2_2767 ( .A(core__abc_22172_new_n4183_), .B(reset_n), .Y(core__abc_22172_new_n4184_));
AND2X2 AND2X2_2768 ( .A(core__abc_22172_new_n4182_), .B(core__abc_22172_new_n4184_), .Y(core__0v3_reg_63_0__15_));
AND2X2 AND2X2_2769 ( .A(core__abc_22172_new_n3217_), .B(core_v3_reg_16_), .Y(core__abc_22172_new_n4186_));
AND2X2 AND2X2_277 ( .A(_abc_19873_new_n916_), .B(core_key_84_), .Y(_abc_19873_new_n1367_));
AND2X2 AND2X2_2770 ( .A(core__abc_22172_new_n4149_), .B(core__abc_22172_new_n4093_), .Y(core__abc_22172_new_n4188_));
AND2X2 AND2X2_2771 ( .A(core__abc_22172_new_n4188_), .B(core__abc_22172_new_n4023_), .Y(core__abc_22172_new_n4189_));
AND2X2 AND2X2_2772 ( .A(core__abc_22172_new_n4189_), .B(core__abc_22172_new_n3932_), .Y(core__abc_22172_new_n4190_));
AND2X2 AND2X2_2773 ( .A(core__abc_22172_new_n4190_), .B(core__abc_22172_new_n3671_), .Y(core__abc_22172_new_n4191_));
AND2X2 AND2X2_2774 ( .A(core__abc_22172_new_n4189_), .B(core__abc_22172_new_n3931_), .Y(core__abc_22172_new_n4192_));
AND2X2 AND2X2_2775 ( .A(core__abc_22172_new_n4188_), .B(core__abc_22172_new_n4064_), .Y(core__abc_22172_new_n4193_));
AND2X2 AND2X2_2776 ( .A(core__abc_22172_new_n4145_), .B(core__abc_22172_new_n4127_), .Y(core__abc_22172_new_n4195_));
AND2X2 AND2X2_2777 ( .A(core__abc_22172_new_n2057_), .B(core__abc_22172_new_n2074_), .Y(core__abc_22172_new_n4200_));
AND2X2 AND2X2_2778 ( .A(core__abc_22172_new_n4072_), .B(core__abc_22172_new_n4200_), .Y(core__abc_22172_new_n4201_));
AND2X2 AND2X2_2779 ( .A(core__abc_22172_new_n3940_), .B(core__abc_22172_new_n4201_), .Y(core__abc_22172_new_n4202_));
AND2X2 AND2X2_278 ( .A(_abc_19873_new_n930_), .B(word0_reg_20_), .Y(_abc_19873_new_n1370_));
AND2X2 AND2X2_2780 ( .A(core__abc_22172_new_n3680_), .B(core__abc_22172_new_n4202_), .Y(core__abc_22172_new_n4203_));
AND2X2 AND2X2_2781 ( .A(core__abc_22172_new_n3939_), .B(core__abc_22172_new_n4201_), .Y(core__abc_22172_new_n4204_));
AND2X2 AND2X2_2782 ( .A(core__abc_22172_new_n4071_), .B(core__abc_22172_new_n4200_), .Y(core__abc_22172_new_n4205_));
AND2X2 AND2X2_2783 ( .A(core__abc_22172_new_n2071_), .B(core__abc_22172_new_n2055_), .Y(core__abc_22172_new_n4206_));
AND2X2 AND2X2_2784 ( .A(core__abc_22172_new_n3681_), .B(core__abc_22172_new_n4202_), .Y(core__abc_22172_new_n4211_));
AND2X2 AND2X2_2785 ( .A(core__abc_22172_new_n3013_), .B(core__abc_22172_new_n4211_), .Y(core__abc_22172_new_n4212_));
AND2X2 AND2X2_2786 ( .A(core__abc_22172_new_n4213_), .B(core__abc_22172_new_n2091_), .Y(core__abc_22172_new_n4214_));
AND2X2 AND2X2_2787 ( .A(core__abc_22172_new_n4217_), .B(core__abc_22172_new_n4215_), .Y(core__abc_22172_new_n4218_));
AND2X2 AND2X2_2788 ( .A(core__abc_22172_new_n4218_), .B(core__abc_22172_new_n2097_), .Y(core__abc_22172_new_n4219_));
AND2X2 AND2X2_2789 ( .A(core__abc_22172_new_n4221_), .B(core__abc_22172_new_n1554_), .Y(core__abc_22172_new_n4222_));
AND2X2 AND2X2_279 ( .A(_abc_19873_new_n907_), .B(word1_reg_20_), .Y(_abc_19873_new_n1371_));
AND2X2 AND2X2_2790 ( .A(core__abc_22172_new_n3099_), .B(core__abc_22172_new_n1551_), .Y(core__abc_22172_new_n4223_));
AND2X2 AND2X2_2791 ( .A(core__abc_22172_new_n4226_), .B(core__abc_22172_new_n4227_), .Y(core__abc_22172_new_n4228_));
AND2X2 AND2X2_2792 ( .A(core__abc_22172_new_n4229_), .B(core__abc_22172_new_n4220_), .Y(core__abc_22172_new_n4230_));
AND2X2 AND2X2_2793 ( .A(core__abc_22172_new_n4231_), .B(core__abc_22172_new_n4228_), .Y(core__abc_22172_new_n4232_));
AND2X2 AND2X2_2794 ( .A(core__abc_22172_new_n4199_), .B(core__abc_22172_new_n4234_), .Y(core__abc_22172_new_n4235_));
AND2X2 AND2X2_2795 ( .A(core__abc_22172_new_n4236_), .B(core__abc_22172_new_n4233_), .Y(core__abc_22172_new_n4237_));
AND2X2 AND2X2_2796 ( .A(core__abc_22172_new_n4240_), .B(core__abc_22172_new_n2264_), .Y(core__abc_22172_new_n4241_));
AND2X2 AND2X2_2797 ( .A(core__abc_22172_new_n4241_), .B(core__abc_22172_new_n2285_), .Y(core__abc_22172_new_n4242_));
AND2X2 AND2X2_2798 ( .A(core__abc_22172_new_n4245_), .B(core_v3_reg_43_), .Y(core__abc_22172_new_n4246_));
AND2X2 AND2X2_2799 ( .A(core__abc_22172_new_n4248_), .B(core__abc_22172_new_n4243_), .Y(core__abc_22172_new_n4249_));
AND2X2 AND2X2_28 ( .A(_abc_19873_new_n904_), .B(_abc_19873_new_n906_), .Y(_abc_19873_new_n907_));
AND2X2 AND2X2_280 ( .A(_abc_19873_new_n919_), .B(core_mi_52_), .Y(_abc_19873_new_n1373_));
AND2X2 AND2X2_2800 ( .A(core__abc_22172_new_n4249_), .B(core__abc_22172_new_n4247_), .Y(core__abc_22172_new_n4250_));
AND2X2 AND2X2_2801 ( .A(core__abc_22172_new_n4254_), .B(core__abc_22172_new_n4253_), .Y(core__abc_22172_new_n4255_));
AND2X2 AND2X2_2802 ( .A(core__abc_22172_new_n4252_), .B(core__abc_22172_new_n4256_), .Y(core__abc_22172_new_n4257_));
AND2X2 AND2X2_2803 ( .A(core__abc_22172_new_n4257_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n4258_));
AND2X2 AND2X2_2804 ( .A(core__abc_22172_new_n3214_), .B(core_key_80_), .Y(core__abc_22172_new_n4259_));
AND2X2 AND2X2_2805 ( .A(core_v3_reg_16_), .B(core_mi_16_), .Y(core__abc_22172_new_n4261_));
AND2X2 AND2X2_2806 ( .A(core__abc_22172_new_n4262_), .B(core__abc_22172_new_n4260_), .Y(core__abc_22172_new_n4263_));
AND2X2 AND2X2_2807 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n4263_), .Y(core__abc_22172_new_n4264_));
AND2X2 AND2X2_2808 ( .A(core__abc_22172_new_n4266_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n4267_));
AND2X2 AND2X2_2809 ( .A(core__abc_22172_new_n4268_), .B(reset_n), .Y(core__0v3_reg_63_0__16_));
AND2X2 AND2X2_281 ( .A(_abc_19873_new_n1377_), .B(_abc_19873_new_n937_), .Y(\read_data[20] ));
AND2X2 AND2X2_2810 ( .A(core__abc_22172_new_n2109_), .B(core__abc_22172_new_n2090_), .Y(core__abc_22172_new_n4273_));
AND2X2 AND2X2_2811 ( .A(core__abc_22172_new_n4272_), .B(core__abc_22172_new_n4273_), .Y(core__abc_22172_new_n4274_));
AND2X2 AND2X2_2812 ( .A(core__abc_22172_new_n2108_), .B(core__abc_22172_new_n2089_), .Y(core__abc_22172_new_n4276_));
AND2X2 AND2X2_2813 ( .A(core__abc_22172_new_n2091_), .B(core__abc_22172_new_n2108_), .Y(core__abc_22172_new_n4278_));
AND2X2 AND2X2_2814 ( .A(core__abc_22172_new_n4280_), .B(core__abc_22172_new_n4277_), .Y(core__abc_22172_new_n4281_));
AND2X2 AND2X2_2815 ( .A(core__abc_22172_new_n4275_), .B(core__abc_22172_new_n4281_), .Y(core__abc_22172_new_n4282_));
AND2X2 AND2X2_2816 ( .A(core__abc_22172_new_n4284_), .B(core__abc_22172_new_n1571_), .Y(core__abc_22172_new_n4285_));
AND2X2 AND2X2_2817 ( .A(core__abc_22172_new_n4283_), .B(core__abc_22172_new_n1568_), .Y(core__abc_22172_new_n4286_));
AND2X2 AND2X2_2818 ( .A(core__abc_22172_new_n4287_), .B(core_v3_reg_1_), .Y(core__abc_22172_new_n4288_));
AND2X2 AND2X2_2819 ( .A(core__abc_22172_new_n4289_), .B(core__abc_22172_new_n1281_), .Y(core__abc_22172_new_n4290_));
AND2X2 AND2X2_282 ( .A(_abc_19873_new_n925_), .B(word2_reg_21_), .Y(_abc_19873_new_n1379_));
AND2X2 AND2X2_2820 ( .A(core__abc_22172_new_n4282_), .B(core__abc_22172_new_n4291_), .Y(core__abc_22172_new_n4292_));
AND2X2 AND2X2_2821 ( .A(core__abc_22172_new_n4293_), .B(core__abc_22172_new_n4294_), .Y(core__abc_22172_new_n4295_));
AND2X2 AND2X2_2822 ( .A(core__abc_22172_new_n4296_), .B(core__abc_22172_new_n4271_), .Y(core__abc_22172_new_n4297_));
AND2X2 AND2X2_2823 ( .A(core__abc_22172_new_n4270_), .B(core__abc_22172_new_n4297_), .Y(core__abc_22172_new_n4298_));
AND2X2 AND2X2_2824 ( .A(core__abc_22172_new_n4295_), .B(core__abc_22172_new_n4232_), .Y(core__abc_22172_new_n4300_));
AND2X2 AND2X2_2825 ( .A(core__abc_22172_new_n4295_), .B(core__abc_22172_new_n4234_), .Y(core__abc_22172_new_n4302_));
AND2X2 AND2X2_2826 ( .A(core__abc_22172_new_n4199_), .B(core__abc_22172_new_n4302_), .Y(core__abc_22172_new_n4303_));
AND2X2 AND2X2_2827 ( .A(core__abc_22172_new_n4304_), .B(core__abc_22172_new_n4301_), .Y(core__abc_22172_new_n4305_));
AND2X2 AND2X2_2828 ( .A(core__abc_22172_new_n4299_), .B(core__abc_22172_new_n4305_), .Y(core__abc_22172_new_n4306_));
AND2X2 AND2X2_2829 ( .A(core__abc_22172_new_n4163_), .B(core__abc_22172_new_n2282_), .Y(core__abc_22172_new_n4308_));
AND2X2 AND2X2_283 ( .A(_abc_19873_new_n901_), .B(core_key_21_), .Y(_abc_19873_new_n1380_));
AND2X2 AND2X2_2830 ( .A(core__abc_22172_new_n2282_), .B(core__abc_22172_new_n2263_), .Y(core__abc_22172_new_n4309_));
AND2X2 AND2X2_2831 ( .A(core__abc_22172_new_n4311_), .B(core__abc_22172_new_n2299_), .Y(core__abc_22172_new_n4312_));
AND2X2 AND2X2_2832 ( .A(core__abc_22172_new_n4313_), .B(core__abc_22172_new_n2302_), .Y(core__abc_22172_new_n4314_));
AND2X2 AND2X2_2833 ( .A(core__abc_22172_new_n4317_), .B(core__abc_22172_new_n4319_), .Y(core__abc_22172_new_n4320_));
AND2X2 AND2X2_2834 ( .A(core__abc_22172_new_n4323_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n4324_));
AND2X2 AND2X2_2835 ( .A(core__abc_22172_new_n4324_), .B(core__abc_22172_new_n4322_), .Y(core__abc_22172_new_n4325_));
AND2X2 AND2X2_2836 ( .A(core__abc_22172_new_n3214_), .B(core_key_81_), .Y(core__abc_22172_new_n4326_));
AND2X2 AND2X2_2837 ( .A(core_v3_reg_17_), .B(core_mi_17_), .Y(core__abc_22172_new_n4327_));
AND2X2 AND2X2_2838 ( .A(core__abc_22172_new_n4328_), .B(core__abc_22172_new_n4329_), .Y(core__abc_22172_new_n4330_));
AND2X2 AND2X2_2839 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n4330_), .Y(core__abc_22172_new_n4331_));
AND2X2 AND2X2_284 ( .A(_abc_19873_new_n928_), .B(core_key_53_), .Y(_abc_19873_new_n1381_));
AND2X2 AND2X2_2840 ( .A(core__abc_22172_new_n4335_), .B(reset_n), .Y(core__abc_22172_new_n4336_));
AND2X2 AND2X2_2841 ( .A(core__abc_22172_new_n4334_), .B(core__abc_22172_new_n4336_), .Y(core__0v3_reg_63_0__17_));
AND2X2 AND2X2_2842 ( .A(core__abc_22172_new_n4304_), .B(core__abc_22172_new_n4339_), .Y(core__abc_22172_new_n4340_));
AND2X2 AND2X2_2843 ( .A(core__abc_22172_new_n4277_), .B(core__abc_22172_new_n2106_), .Y(core__abc_22172_new_n4342_));
AND2X2 AND2X2_2844 ( .A(core__abc_22172_new_n4280_), .B(core__abc_22172_new_n4342_), .Y(core__abc_22172_new_n4343_));
AND2X2 AND2X2_2845 ( .A(core__abc_22172_new_n4343_), .B(core__abc_22172_new_n2131_), .Y(core__abc_22172_new_n4345_));
AND2X2 AND2X2_2846 ( .A(core__abc_22172_new_n4346_), .B(core__abc_22172_new_n4344_), .Y(core__abc_22172_new_n4347_));
AND2X2 AND2X2_2847 ( .A(core__abc_22172_new_n3099_), .B(core__abc_22172_new_n3111_), .Y(core__abc_22172_new_n4348_));
AND2X2 AND2X2_2848 ( .A(core__abc_22172_new_n4349_), .B(core__abc_22172_new_n1585_), .Y(core__abc_22172_new_n4350_));
AND2X2 AND2X2_2849 ( .A(core__abc_22172_new_n4351_), .B(core__abc_22172_new_n4352_), .Y(core__abc_22172_new_n4353_));
AND2X2 AND2X2_285 ( .A(_abc_19873_new_n881_), .B(core_key_117_), .Y(_abc_19873_new_n1383_));
AND2X2 AND2X2_2850 ( .A(core__abc_22172_new_n4356_), .B(core__abc_22172_new_n4354_), .Y(core__abc_22172_new_n4357_));
AND2X2 AND2X2_2851 ( .A(core__abc_22172_new_n4347_), .B(core__abc_22172_new_n4358_), .Y(core__abc_22172_new_n4359_));
AND2X2 AND2X2_2852 ( .A(core__abc_22172_new_n4360_), .B(core__abc_22172_new_n4357_), .Y(core__abc_22172_new_n4361_));
AND2X2 AND2X2_2853 ( .A(core__abc_22172_new_n4341_), .B(core__abc_22172_new_n4363_), .Y(core__abc_22172_new_n4364_));
AND2X2 AND2X2_2854 ( .A(core__abc_22172_new_n4340_), .B(core__abc_22172_new_n4362_), .Y(core__abc_22172_new_n4365_));
AND2X2 AND2X2_2855 ( .A(core__abc_22172_new_n4367_), .B(core__abc_22172_new_n2319_), .Y(core__abc_22172_new_n4368_));
AND2X2 AND2X2_2856 ( .A(core__abc_22172_new_n4369_), .B(core__abc_22172_new_n4370_), .Y(core__abc_22172_new_n4371_));
AND2X2 AND2X2_2857 ( .A(core__abc_22172_new_n4372_), .B(core_v3_reg_45_), .Y(core__abc_22172_new_n4373_));
AND2X2 AND2X2_2858 ( .A(core__abc_22172_new_n4371_), .B(core__abc_22172_new_n4374_), .Y(core__abc_22172_new_n4375_));
AND2X2 AND2X2_2859 ( .A(core__abc_22172_new_n4379_), .B(core__abc_22172_new_n4380_), .Y(core__abc_22172_new_n4381_));
AND2X2 AND2X2_286 ( .A(_abc_19873_new_n916_), .B(core_key_85_), .Y(_abc_19873_new_n1384_));
AND2X2 AND2X2_2860 ( .A(core__abc_22172_new_n4382_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n4383_));
AND2X2 AND2X2_2861 ( .A(core__abc_22172_new_n4383_), .B(core__abc_22172_new_n4377_), .Y(core__abc_22172_new_n4384_));
AND2X2 AND2X2_2862 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n4385_), .Y(core__abc_22172_new_n4386_));
AND2X2 AND2X2_2863 ( .A(core_v3_reg_18_), .B(core_mi_18_), .Y(core__abc_22172_new_n4387_));
AND2X2 AND2X2_2864 ( .A(core__abc_22172_new_n4388_), .B(core__abc_22172_new_n4389_), .Y(core__abc_22172_new_n4390_));
AND2X2 AND2X2_2865 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n4390_), .Y(core__abc_22172_new_n4391_));
AND2X2 AND2X2_2866 ( .A(core__abc_22172_new_n4395_), .B(reset_n), .Y(core__abc_22172_new_n4396_));
AND2X2 AND2X2_2867 ( .A(core__abc_22172_new_n4394_), .B(core__abc_22172_new_n4396_), .Y(core__0v3_reg_63_0__18_));
AND2X2 AND2X2_2868 ( .A(core__abc_22172_new_n4344_), .B(core__abc_22172_new_n2124_), .Y(core__abc_22172_new_n4399_));
AND2X2 AND2X2_2869 ( .A(core__abc_22172_new_n4399_), .B(core__abc_22172_new_n2148_), .Y(core__abc_22172_new_n4400_));
AND2X2 AND2X2_287 ( .A(_abc_19873_new_n912_), .B(word3_reg_21_), .Y(_abc_19873_new_n1388_));
AND2X2 AND2X2_2870 ( .A(core__abc_22172_new_n4401_), .B(core__abc_22172_new_n4402_), .Y(core__abc_22172_new_n4403_));
AND2X2 AND2X2_2871 ( .A(core__abc_22172_new_n4351_), .B(core__abc_22172_new_n1583_), .Y(core__abc_22172_new_n4404_));
AND2X2 AND2X2_2872 ( .A(core__abc_22172_new_n4404_), .B(core__abc_22172_new_n1605_), .Y(core__abc_22172_new_n4405_));
AND2X2 AND2X2_2873 ( .A(core__abc_22172_new_n4406_), .B(core__abc_22172_new_n4407_), .Y(core__abc_22172_new_n4408_));
AND2X2 AND2X2_2874 ( .A(core__abc_22172_new_n4409_), .B(core_v3_reg_3_), .Y(core__abc_22172_new_n4410_));
AND2X2 AND2X2_2875 ( .A(core__abc_22172_new_n4408_), .B(core__abc_22172_new_n1320_), .Y(core__abc_22172_new_n4411_));
AND2X2 AND2X2_2876 ( .A(core__abc_22172_new_n4403_), .B(core__abc_22172_new_n4412_), .Y(core__abc_22172_new_n4413_));
AND2X2 AND2X2_2877 ( .A(core__abc_22172_new_n4414_), .B(core__abc_22172_new_n4415_), .Y(core__abc_22172_new_n4416_));
AND2X2 AND2X2_2878 ( .A(core__abc_22172_new_n4398_), .B(core__abc_22172_new_n4416_), .Y(core__abc_22172_new_n4417_));
AND2X2 AND2X2_2879 ( .A(core__abc_22172_new_n4418_), .B(core__abc_22172_new_n4419_), .Y(core__abc_22172_new_n4420_));
AND2X2 AND2X2_288 ( .A(_abc_19873_new_n907_), .B(word1_reg_21_), .Y(_abc_19873_new_n1389_));
AND2X2 AND2X2_2880 ( .A(core__abc_22172_new_n4423_), .B(core__abc_22172_new_n2313_), .Y(core__abc_22172_new_n4424_));
AND2X2 AND2X2_2881 ( .A(core__abc_22172_new_n4424_), .B(core__abc_22172_new_n2333_), .Y(core__abc_22172_new_n4426_));
AND2X2 AND2X2_2882 ( .A(core__abc_22172_new_n4427_), .B(core__abc_22172_new_n4425_), .Y(core__abc_22172_new_n4428_));
AND2X2 AND2X2_2883 ( .A(core__abc_22172_new_n4429_), .B(core__abc_22172_new_n4422_), .Y(core__abc_22172_new_n4430_));
AND2X2 AND2X2_2884 ( .A(core__abc_22172_new_n4428_), .B(core_v3_reg_46_), .Y(core__abc_22172_new_n4431_));
AND2X2 AND2X2_2885 ( .A(core__abc_22172_new_n4435_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n4436_));
AND2X2 AND2X2_2886 ( .A(core__abc_22172_new_n4436_), .B(core__abc_22172_new_n4433_), .Y(core__abc_22172_new_n4437_));
AND2X2 AND2X2_2887 ( .A(core__abc_22172_new_n3214_), .B(core_key_83_), .Y(core__abc_22172_new_n4438_));
AND2X2 AND2X2_2888 ( .A(core_v3_reg_19_), .B(core_mi_19_), .Y(core__abc_22172_new_n4439_));
AND2X2 AND2X2_2889 ( .A(core__abc_22172_new_n4440_), .B(core__abc_22172_new_n4441_), .Y(core__abc_22172_new_n4442_));
AND2X2 AND2X2_289 ( .A(_abc_19873_new_n930_), .B(word0_reg_21_), .Y(_abc_19873_new_n1390_));
AND2X2 AND2X2_2890 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n4442_), .Y(core__abc_22172_new_n4443_));
AND2X2 AND2X2_2891 ( .A(core__abc_22172_new_n4447_), .B(reset_n), .Y(core__abc_22172_new_n4448_));
AND2X2 AND2X2_2892 ( .A(core__abc_22172_new_n4446_), .B(core__abc_22172_new_n4448_), .Y(core__0v3_reg_63_0__19_));
AND2X2 AND2X2_2893 ( .A(core__abc_22172_new_n4416_), .B(core__abc_22172_new_n4363_), .Y(core__abc_22172_new_n4450_));
AND2X2 AND2X2_2894 ( .A(core__abc_22172_new_n4450_), .B(core__abc_22172_new_n4338_), .Y(core__abc_22172_new_n4451_));
AND2X2 AND2X2_2895 ( .A(core__abc_22172_new_n4452_), .B(core__abc_22172_new_n4415_), .Y(core__abc_22172_new_n4453_));
AND2X2 AND2X2_2896 ( .A(core__abc_22172_new_n4450_), .B(core__abc_22172_new_n4302_), .Y(core__abc_22172_new_n4455_));
AND2X2 AND2X2_2897 ( .A(core__abc_22172_new_n4199_), .B(core__abc_22172_new_n4455_), .Y(core__abc_22172_new_n4456_));
AND2X2 AND2X2_2898 ( .A(core__abc_22172_new_n2125_), .B(core__abc_22172_new_n2142_), .Y(core__abc_22172_new_n4458_));
AND2X2 AND2X2_2899 ( .A(core__abc_22172_new_n2139_), .B(core__abc_22172_new_n2123_), .Y(core__abc_22172_new_n4461_));
AND2X2 AND2X2_29 ( .A(_abc_19873_new_n907_), .B(word1_reg_0_), .Y(_abc_19873_new_n908_));
AND2X2 AND2X2_290 ( .A(_abc_19873_new_n888_), .B(core_mi_21_), .Y(_abc_19873_new_n1393_));
AND2X2 AND2X2_2900 ( .A(core__abc_22172_new_n4460_), .B(core__abc_22172_new_n4463_), .Y(core__abc_22172_new_n4464_));
AND2X2 AND2X2_2901 ( .A(core__abc_22172_new_n4278_), .B(core__abc_22172_new_n4458_), .Y(core__abc_22172_new_n4466_));
AND2X2 AND2X2_2902 ( .A(core__abc_22172_new_n4213_), .B(core__abc_22172_new_n4466_), .Y(core__abc_22172_new_n4467_));
AND2X2 AND2X2_2903 ( .A(core__abc_22172_new_n4468_), .B(core__abc_22172_new_n2159_), .Y(core__abc_22172_new_n4469_));
AND2X2 AND2X2_2904 ( .A(core__abc_22172_new_n4470_), .B(core__abc_22172_new_n2165_), .Y(core__abc_22172_new_n4471_));
AND2X2 AND2X2_2905 ( .A(core__abc_22172_new_n3099_), .B(core__abc_22172_new_n3112_), .Y(core__abc_22172_new_n4474_));
AND2X2 AND2X2_2906 ( .A(core__abc_22172_new_n4475_), .B(core__abc_22172_new_n1619_), .Y(core__abc_22172_new_n4476_));
AND2X2 AND2X2_2907 ( .A(core__abc_22172_new_n4477_), .B(core__abc_22172_new_n1622_), .Y(core__abc_22172_new_n4478_));
AND2X2 AND2X2_2908 ( .A(core__abc_22172_new_n4481_), .B(core__abc_22172_new_n4482_), .Y(core__abc_22172_new_n4483_));
AND2X2 AND2X2_2909 ( .A(core__abc_22172_new_n4473_), .B(core__abc_22172_new_n4484_), .Y(core__abc_22172_new_n4485_));
AND2X2 AND2X2_291 ( .A(_abc_19873_new_n919_), .B(core_mi_53_), .Y(_abc_19873_new_n1394_));
AND2X2 AND2X2_2910 ( .A(core__abc_22172_new_n4472_), .B(core__abc_22172_new_n4483_), .Y(core__abc_22172_new_n4486_));
AND2X2 AND2X2_2911 ( .A(core__abc_22172_new_n4457_), .B(core__abc_22172_new_n4488_), .Y(core__abc_22172_new_n4489_));
AND2X2 AND2X2_2912 ( .A(core__abc_22172_new_n4490_), .B(core__abc_22172_new_n4491_), .Y(core__abc_22172_new_n4492_));
AND2X2 AND2X2_2913 ( .A(core__abc_22172_new_n4494_), .B(core__abc_22172_new_n2352_), .Y(core__abc_22172_new_n4496_));
AND2X2 AND2X2_2914 ( .A(core__abc_22172_new_n4497_), .B(core__abc_22172_new_n4495_), .Y(core__abc_22172_new_n4498_));
AND2X2 AND2X2_2915 ( .A(core__abc_22172_new_n4502_), .B(core__abc_22172_new_n4499_), .Y(core__abc_22172_new_n4503_));
AND2X2 AND2X2_2916 ( .A(core__abc_22172_new_n4506_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n4507_));
AND2X2 AND2X2_2917 ( .A(core__abc_22172_new_n4507_), .B(core__abc_22172_new_n4505_), .Y(core__abc_22172_new_n4508_));
AND2X2 AND2X2_2918 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n4509_), .Y(core__abc_22172_new_n4510_));
AND2X2 AND2X2_2919 ( .A(core_v3_reg_20_), .B(core_mi_20_), .Y(core__abc_22172_new_n4511_));
AND2X2 AND2X2_292 ( .A(_abc_19873_new_n1398_), .B(_abc_19873_new_n937_), .Y(\read_data[21] ));
AND2X2 AND2X2_2920 ( .A(core__abc_22172_new_n4512_), .B(core__abc_22172_new_n4513_), .Y(core__abc_22172_new_n4514_));
AND2X2 AND2X2_2921 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n4514_), .Y(core__abc_22172_new_n4515_));
AND2X2 AND2X2_2922 ( .A(core__abc_22172_new_n4519_), .B(reset_n), .Y(core__abc_22172_new_n4520_));
AND2X2 AND2X2_2923 ( .A(core__abc_22172_new_n4518_), .B(core__abc_22172_new_n4520_), .Y(core__0v3_reg_63_0__20_));
AND2X2 AND2X2_2924 ( .A(core__abc_22172_new_n4523_), .B(core__abc_22172_new_n2177_), .Y(core__abc_22172_new_n4524_));
AND2X2 AND2X2_2925 ( .A(core__abc_22172_new_n4522_), .B(core__abc_22172_new_n2176_), .Y(core__abc_22172_new_n4525_));
AND2X2 AND2X2_2926 ( .A(core__abc_22172_new_n4528_), .B(core__abc_22172_new_n1636_), .Y(core__abc_22172_new_n4530_));
AND2X2 AND2X2_2927 ( .A(core__abc_22172_new_n4531_), .B(core__abc_22172_new_n4529_), .Y(core__abc_22172_new_n4532_));
AND2X2 AND2X2_2928 ( .A(core__abc_22172_new_n4533_), .B(core_v3_reg_5_), .Y(core__abc_22172_new_n4534_));
AND2X2 AND2X2_2929 ( .A(core__abc_22172_new_n4532_), .B(core__abc_22172_new_n1357_), .Y(core__abc_22172_new_n4535_));
AND2X2 AND2X2_293 ( .A(_abc_19873_new_n881_), .B(core_key_118_), .Y(_abc_19873_new_n1400_));
AND2X2 AND2X2_2930 ( .A(core__abc_22172_new_n4537_), .B(core__abc_22172_new_n4539_), .Y(core__abc_22172_new_n4540_));
AND2X2 AND2X2_2931 ( .A(core__abc_22172_new_n4490_), .B(core__abc_22172_new_n4542_), .Y(core__abc_22172_new_n4543_));
AND2X2 AND2X2_2932 ( .A(core__abc_22172_new_n4543_), .B(core__abc_22172_new_n4541_), .Y(core__abc_22172_new_n4544_));
AND2X2 AND2X2_2933 ( .A(core__abc_22172_new_n4550_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n4551_));
AND2X2 AND2X2_2934 ( .A(core__abc_22172_new_n4551_), .B(core__abc_22172_new_n4549_), .Y(core__abc_22172_new_n4552_));
AND2X2 AND2X2_2935 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n4553_), .Y(core__abc_22172_new_n4554_));
AND2X2 AND2X2_2936 ( .A(core_v3_reg_21_), .B(core_mi_21_), .Y(core__abc_22172_new_n4555_));
AND2X2 AND2X2_2937 ( .A(core__abc_22172_new_n4556_), .B(core__abc_22172_new_n4557_), .Y(core__abc_22172_new_n4558_));
AND2X2 AND2X2_2938 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n4558_), .Y(core__abc_22172_new_n4559_));
AND2X2 AND2X2_2939 ( .A(core__abc_22172_new_n4563_), .B(reset_n), .Y(core__abc_22172_new_n4564_));
AND2X2 AND2X2_294 ( .A(_abc_19873_new_n888_), .B(core_mi_22_), .Y(_abc_19873_new_n1401_));
AND2X2 AND2X2_2940 ( .A(core__abc_22172_new_n4562_), .B(core__abc_22172_new_n4564_), .Y(core__0v3_reg_63_0__21_));
AND2X2 AND2X2_2941 ( .A(core__abc_22172_new_n4540_), .B(core__abc_22172_new_n4488_), .Y(core__abc_22172_new_n4567_));
AND2X2 AND2X2_2942 ( .A(core__abc_22172_new_n4457_), .B(core__abc_22172_new_n4567_), .Y(core__abc_22172_new_n4568_));
AND2X2 AND2X2_2943 ( .A(core__abc_22172_new_n4570_), .B(core__abc_22172_new_n4537_), .Y(core__abc_22172_new_n4571_));
AND2X2 AND2X2_2944 ( .A(core__abc_22172_new_n2159_), .B(core__abc_22172_new_n2176_), .Y(core__abc_22172_new_n4573_));
AND2X2 AND2X2_2945 ( .A(core__abc_22172_new_n4468_), .B(core__abc_22172_new_n4573_), .Y(core__abc_22172_new_n4574_));
AND2X2 AND2X2_2946 ( .A(core__abc_22172_new_n2158_), .B(core__abc_22172_new_n2174_), .Y(core__abc_22172_new_n4576_));
AND2X2 AND2X2_2947 ( .A(core__abc_22172_new_n4579_), .B(core__abc_22172_new_n2193_), .Y(core__abc_22172_new_n4580_));
AND2X2 AND2X2_2948 ( .A(core__abc_22172_new_n4581_), .B(core__abc_22172_new_n2199_), .Y(core__abc_22172_new_n4582_));
AND2X2 AND2X2_2949 ( .A(core__abc_22172_new_n4475_), .B(core__abc_22172_new_n3108_), .Y(core__abc_22172_new_n4584_));
AND2X2 AND2X2_295 ( .A(_abc_19873_new_n916_), .B(core_key_86_), .Y(_abc_19873_new_n1403_));
AND2X2 AND2X2_2950 ( .A(core__abc_22172_new_n4585_), .B(core__abc_22172_new_n1653_), .Y(core__abc_22172_new_n4586_));
AND2X2 AND2X2_2951 ( .A(core__abc_22172_new_n4587_), .B(core__abc_22172_new_n1656_), .Y(core__abc_22172_new_n4588_));
AND2X2 AND2X2_2952 ( .A(core__abc_22172_new_n4591_), .B(core__abc_22172_new_n4592_), .Y(core__abc_22172_new_n4593_));
AND2X2 AND2X2_2953 ( .A(core__abc_22172_new_n4583_), .B(core__abc_22172_new_n4594_), .Y(core__abc_22172_new_n4595_));
AND2X2 AND2X2_2954 ( .A(core__abc_22172_new_n4596_), .B(core__abc_22172_new_n4597_), .Y(core__abc_22172_new_n4598_));
AND2X2 AND2X2_2955 ( .A(core__abc_22172_new_n4572_), .B(core__abc_22172_new_n4598_), .Y(core__abc_22172_new_n4599_));
AND2X2 AND2X2_2956 ( .A(core__abc_22172_new_n4600_), .B(core__abc_22172_new_n4601_), .Y(core__abc_22172_new_n4602_));
AND2X2 AND2X2_2957 ( .A(core__abc_22172_new_n4605_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n4606_));
AND2X2 AND2X2_2958 ( .A(core__abc_22172_new_n4606_), .B(core__abc_22172_new_n4603_), .Y(core__abc_22172_new_n4607_));
AND2X2 AND2X2_2959 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n4608_), .Y(core__abc_22172_new_n4609_));
AND2X2 AND2X2_296 ( .A(_abc_19873_new_n925_), .B(word2_reg_22_), .Y(_abc_19873_new_n1406_));
AND2X2 AND2X2_2960 ( .A(core_v3_reg_22_), .B(core_mi_22_), .Y(core__abc_22172_new_n4610_));
AND2X2 AND2X2_2961 ( .A(core__abc_22172_new_n4611_), .B(core__abc_22172_new_n4612_), .Y(core__abc_22172_new_n4613_));
AND2X2 AND2X2_2962 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n4613_), .Y(core__abc_22172_new_n4614_));
AND2X2 AND2X2_2963 ( .A(core__abc_22172_new_n4618_), .B(reset_n), .Y(core__abc_22172_new_n4619_));
AND2X2 AND2X2_2964 ( .A(core__abc_22172_new_n4617_), .B(core__abc_22172_new_n4619_), .Y(core__0v3_reg_63_0__22_));
AND2X2 AND2X2_2965 ( .A(core__abc_22172_new_n4600_), .B(core__abc_22172_new_n4597_), .Y(core__abc_22172_new_n4621_));
AND2X2 AND2X2_2966 ( .A(core__abc_22172_new_n4622_), .B(core__abc_22172_new_n2210_), .Y(core__abc_22172_new_n4624_));
AND2X2 AND2X2_2967 ( .A(core__abc_22172_new_n4625_), .B(core__abc_22172_new_n4623_), .Y(core__abc_22172_new_n4626_));
AND2X2 AND2X2_2968 ( .A(core__abc_22172_new_n4628_), .B(core__abc_22172_new_n1673_), .Y(core__abc_22172_new_n4629_));
AND2X2 AND2X2_2969 ( .A(core__abc_22172_new_n4627_), .B(core__abc_22172_new_n1670_), .Y(core__abc_22172_new_n4630_));
AND2X2 AND2X2_297 ( .A(_abc_19873_new_n907_), .B(word1_reg_22_), .Y(_abc_19873_new_n1407_));
AND2X2 AND2X2_2970 ( .A(core__abc_22172_new_n4631_), .B(core_v3_reg_7_), .Y(core__abc_22172_new_n4632_));
AND2X2 AND2X2_2971 ( .A(core__abc_22172_new_n4633_), .B(core__abc_22172_new_n1395_), .Y(core__abc_22172_new_n4634_));
AND2X2 AND2X2_2972 ( .A(core__abc_22172_new_n4640_), .B(core__abc_22172_new_n4636_), .Y(core__abc_22172_new_n4641_));
AND2X2 AND2X2_2973 ( .A(core__abc_22172_new_n4621_), .B(core__abc_22172_new_n4642_), .Y(core__abc_22172_new_n4643_));
AND2X2 AND2X2_2974 ( .A(core__abc_22172_new_n4644_), .B(core__abc_22172_new_n4645_), .Y(core__abc_22172_new_n4646_));
AND2X2 AND2X2_2975 ( .A(core__abc_22172_new_n4649_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n4650_));
AND2X2 AND2X2_2976 ( .A(core__abc_22172_new_n4650_), .B(core__abc_22172_new_n4647_), .Y(core__abc_22172_new_n4651_));
AND2X2 AND2X2_2977 ( .A(core__abc_22172_new_n3214_), .B(core_key_87_), .Y(core__abc_22172_new_n4652_));
AND2X2 AND2X2_2978 ( .A(core_v3_reg_23_), .B(core_mi_23_), .Y(core__abc_22172_new_n4653_));
AND2X2 AND2X2_2979 ( .A(core__abc_22172_new_n4654_), .B(core__abc_22172_new_n4655_), .Y(core__abc_22172_new_n4656_));
AND2X2 AND2X2_298 ( .A(_abc_19873_new_n912_), .B(word3_reg_22_), .Y(_abc_19873_new_n1408_));
AND2X2 AND2X2_2980 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n4656_), .Y(core__abc_22172_new_n4657_));
AND2X2 AND2X2_2981 ( .A(core__abc_22172_new_n4661_), .B(reset_n), .Y(core__abc_22172_new_n4662_));
AND2X2 AND2X2_2982 ( .A(core__abc_22172_new_n4660_), .B(core__abc_22172_new_n4662_), .Y(core__0v3_reg_63_0__23_));
AND2X2 AND2X2_2983 ( .A(core__abc_22172_new_n4641_), .B(core__abc_22172_new_n4598_), .Y(core__abc_22172_new_n4664_));
AND2X2 AND2X2_2984 ( .A(core__abc_22172_new_n4664_), .B(core__abc_22172_new_n4567_), .Y(core__abc_22172_new_n4665_));
AND2X2 AND2X2_2985 ( .A(core__abc_22172_new_n4665_), .B(core__abc_22172_new_n4454_), .Y(core__abc_22172_new_n4666_));
AND2X2 AND2X2_2986 ( .A(core__abc_22172_new_n4664_), .B(core__abc_22172_new_n4571_), .Y(core__abc_22172_new_n4667_));
AND2X2 AND2X2_2987 ( .A(core__abc_22172_new_n4636_), .B(core__abc_22172_new_n4669_), .Y(core__abc_22172_new_n4670_));
AND2X2 AND2X2_2988 ( .A(core__abc_22172_new_n4665_), .B(core__abc_22172_new_n4455_), .Y(core__abc_22172_new_n4674_));
AND2X2 AND2X2_2989 ( .A(core__abc_22172_new_n4199_), .B(core__abc_22172_new_n4674_), .Y(core__abc_22172_new_n4675_));
AND2X2 AND2X2_299 ( .A(_abc_19873_new_n919_), .B(core_mi_54_), .Y(_abc_19873_new_n1411_));
AND2X2 AND2X2_2990 ( .A(core__abc_22172_new_n2193_), .B(core__abc_22172_new_n2210_), .Y(core__abc_22172_new_n4677_));
AND2X2 AND2X2_2991 ( .A(core__abc_22172_new_n4573_), .B(core__abc_22172_new_n4677_), .Y(core__abc_22172_new_n4678_));
AND2X2 AND2X2_2992 ( .A(core__abc_22172_new_n4466_), .B(core__abc_22172_new_n4678_), .Y(core__abc_22172_new_n4679_));
AND2X2 AND2X2_2993 ( .A(core__abc_22172_new_n4213_), .B(core__abc_22172_new_n4679_), .Y(core__abc_22172_new_n4680_));
AND2X2 AND2X2_2994 ( .A(core__abc_22172_new_n4465_), .B(core__abc_22172_new_n4678_), .Y(core__abc_22172_new_n4681_));
AND2X2 AND2X2_2995 ( .A(core__abc_22172_new_n4578_), .B(core__abc_22172_new_n4677_), .Y(core__abc_22172_new_n4682_));
AND2X2 AND2X2_2996 ( .A(core__abc_22172_new_n2207_), .B(core__abc_22172_new_n2191_), .Y(core__abc_22172_new_n4683_));
AND2X2 AND2X2_2997 ( .A(core__abc_22172_new_n4687_), .B(core__abc_22172_new_n2227_), .Y(core__abc_22172_new_n4688_));
AND2X2 AND2X2_2998 ( .A(core__abc_22172_new_n4690_), .B(core__abc_22172_new_n4691_), .Y(core__abc_22172_new_n4692_));
AND2X2 AND2X2_2999 ( .A(core__abc_22172_new_n4692_), .B(core__abc_22172_new_n2233_), .Y(core__abc_22172_new_n4693_));
AND2X2 AND2X2_3 ( .A(_abc_19873_new_n872_), .B(_abc_19873_new_n874_), .Y(_abc_19873_new_n875_));
AND2X2 AND2X2_30 ( .A(_abc_19873_new_n880_), .B(_abc_19873_new_n906_), .Y(_abc_19873_new_n912_));
AND2X2 AND2X2_300 ( .A(_abc_19873_new_n930_), .B(word0_reg_22_), .Y(_abc_19873_new_n1412_));
AND2X2 AND2X2_3000 ( .A(core__abc_22172_new_n3099_), .B(core__abc_22172_new_n3113_), .Y(core__abc_22172_new_n4695_));
AND2X2 AND2X2_3001 ( .A(core__abc_22172_new_n4696_), .B(core__abc_22172_new_n1687_), .Y(core__abc_22172_new_n4697_));
AND2X2 AND2X2_3002 ( .A(core__abc_22172_new_n4698_), .B(core__abc_22172_new_n1690_), .Y(core__abc_22172_new_n4699_));
AND2X2 AND2X2_3003 ( .A(core__abc_22172_new_n4702_), .B(core__abc_22172_new_n4704_), .Y(core__abc_22172_new_n4705_));
AND2X2 AND2X2_3004 ( .A(core__abc_22172_new_n4706_), .B(core__abc_22172_new_n4694_), .Y(core__abc_22172_new_n4707_));
AND2X2 AND2X2_3005 ( .A(core__abc_22172_new_n4708_), .B(core__abc_22172_new_n4705_), .Y(core__abc_22172_new_n4709_));
AND2X2 AND2X2_3006 ( .A(core__abc_22172_new_n4676_), .B(core__abc_22172_new_n4711_), .Y(core__abc_22172_new_n4712_));
AND2X2 AND2X2_3007 ( .A(core__abc_22172_new_n4713_), .B(core__abc_22172_new_n4710_), .Y(core__abc_22172_new_n4714_));
AND2X2 AND2X2_3008 ( .A(core__abc_22172_new_n4718_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n4719_));
AND2X2 AND2X2_3009 ( .A(core__abc_22172_new_n4719_), .B(core__abc_22172_new_n4716_), .Y(core__abc_22172_new_n4720_));
AND2X2 AND2X2_301 ( .A(_abc_19873_new_n928_), .B(core_key_54_), .Y(_abc_19873_new_n1414_));
AND2X2 AND2X2_3010 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n4721_), .Y(core__abc_22172_new_n4722_));
AND2X2 AND2X2_3011 ( .A(core_v3_reg_24_), .B(core_mi_24_), .Y(core__abc_22172_new_n4723_));
AND2X2 AND2X2_3012 ( .A(core__abc_22172_new_n4724_), .B(core__abc_22172_new_n4725_), .Y(core__abc_22172_new_n4726_));
AND2X2 AND2X2_3013 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n4726_), .Y(core__abc_22172_new_n4727_));
AND2X2 AND2X2_3014 ( .A(core__abc_22172_new_n4731_), .B(reset_n), .Y(core__abc_22172_new_n4732_));
AND2X2 AND2X2_3015 ( .A(core__abc_22172_new_n4730_), .B(core__abc_22172_new_n4732_), .Y(core__0v3_reg_63_0__24_));
AND2X2 AND2X2_3016 ( .A(core__abc_22172_new_n4735_), .B(core__abc_22172_new_n2250_), .Y(core__abc_22172_new_n4736_));
AND2X2 AND2X2_3017 ( .A(core__abc_22172_new_n4734_), .B(core__abc_22172_new_n2244_), .Y(core__abc_22172_new_n4737_));
AND2X2 AND2X2_3018 ( .A(core__abc_22172_new_n4740_), .B(core__abc_22172_new_n1707_), .Y(core__abc_22172_new_n4741_));
AND2X2 AND2X2_3019 ( .A(core__abc_22172_new_n4739_), .B(core__abc_22172_new_n1704_), .Y(core__abc_22172_new_n4742_));
AND2X2 AND2X2_302 ( .A(_abc_19873_new_n901_), .B(core_key_22_), .Y(_abc_19873_new_n1415_));
AND2X2 AND2X2_3020 ( .A(core__abc_22172_new_n4743_), .B(core_v3_reg_9_), .Y(core__abc_22172_new_n4744_));
AND2X2 AND2X2_3021 ( .A(core__abc_22172_new_n4745_), .B(core__abc_22172_new_n4746_), .Y(core__abc_22172_new_n4747_));
AND2X2 AND2X2_3022 ( .A(core__abc_22172_new_n4738_), .B(core__abc_22172_new_n4747_), .Y(core__abc_22172_new_n4748_));
AND2X2 AND2X2_3023 ( .A(core__abc_22172_new_n4749_), .B(core__abc_22172_new_n4750_), .Y(core__abc_22172_new_n4751_));
AND2X2 AND2X2_3024 ( .A(core__abc_22172_new_n4754_), .B(core__abc_22172_new_n4753_), .Y(core__abc_22172_new_n4755_));
AND2X2 AND2X2_3025 ( .A(core__abc_22172_new_n4755_), .B(core__abc_22172_new_n4752_), .Y(core__abc_22172_new_n4756_));
AND2X2 AND2X2_3026 ( .A(core__abc_22172_new_n4762_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n4763_));
AND2X2 AND2X2_3027 ( .A(core__abc_22172_new_n4763_), .B(core__abc_22172_new_n4761_), .Y(core__abc_22172_new_n4764_));
AND2X2 AND2X2_3028 ( .A(core__abc_22172_new_n3214_), .B(core_key_89_), .Y(core__abc_22172_new_n4765_));
AND2X2 AND2X2_3029 ( .A(core_v3_reg_25_), .B(core_mi_25_), .Y(core__abc_22172_new_n4766_));
AND2X2 AND2X2_303 ( .A(_abc_19873_new_n1419_), .B(_abc_19873_new_n937_), .Y(\read_data[22] ));
AND2X2 AND2X2_3030 ( .A(core__abc_22172_new_n4767_), .B(core__abc_22172_new_n4768_), .Y(core__abc_22172_new_n4769_));
AND2X2 AND2X2_3031 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n4769_), .Y(core__abc_22172_new_n4770_));
AND2X2 AND2X2_3032 ( .A(core__abc_22172_new_n4774_), .B(reset_n), .Y(core__abc_22172_new_n4775_));
AND2X2 AND2X2_3033 ( .A(core__abc_22172_new_n4773_), .B(core__abc_22172_new_n4775_), .Y(core__0v3_reg_63_0__25_));
AND2X2 AND2X2_3034 ( .A(core__abc_22172_new_n4777_), .B(core__abc_22172_new_n4711_), .Y(core__abc_22172_new_n4778_));
AND2X2 AND2X2_3035 ( .A(core__abc_22172_new_n4676_), .B(core__abc_22172_new_n4778_), .Y(core__abc_22172_new_n4779_));
AND2X2 AND2X2_3036 ( .A(core__abc_22172_new_n4781_), .B(core__abc_22172_new_n4780_), .Y(core__abc_22172_new_n4782_));
AND2X2 AND2X2_3037 ( .A(core__abc_22172_new_n2227_), .B(core__abc_22172_new_n2244_), .Y(core__abc_22172_new_n4784_));
AND2X2 AND2X2_3038 ( .A(core__abc_22172_new_n4687_), .B(core__abc_22172_new_n4784_), .Y(core__abc_22172_new_n4785_));
AND2X2 AND2X2_3039 ( .A(core__abc_22172_new_n2244_), .B(core__abc_22172_new_n2225_), .Y(core__abc_22172_new_n4786_));
AND2X2 AND2X2_304 ( .A(_abc_19873_new_n881_), .B(core_key_119_), .Y(_abc_19873_new_n1421_));
AND2X2 AND2X2_3040 ( .A(core__abc_22172_new_n4788_), .B(core__abc_22172_new_n2261_), .Y(core__abc_22172_new_n4789_));
AND2X2 AND2X2_3041 ( .A(core__abc_22172_new_n4790_), .B(core__abc_22172_new_n2267_), .Y(core__abc_22172_new_n4791_));
AND2X2 AND2X2_3042 ( .A(core__abc_22172_new_n4696_), .B(core__abc_22172_new_n3104_), .Y(core__abc_22172_new_n4795_));
AND2X2 AND2X2_3043 ( .A(core__abc_22172_new_n4797_), .B(core__abc_22172_new_n1724_), .Y(core__abc_22172_new_n4798_));
AND2X2 AND2X2_3044 ( .A(core__abc_22172_new_n4796_), .B(core__abc_22172_new_n1721_), .Y(core__abc_22172_new_n4799_));
AND2X2 AND2X2_3045 ( .A(core__abc_22172_new_n4802_), .B(core__abc_22172_new_n4803_), .Y(core__abc_22172_new_n4804_));
AND2X2 AND2X2_3046 ( .A(core__abc_22172_new_n4793_), .B(core__abc_22172_new_n4805_), .Y(core__abc_22172_new_n4806_));
AND2X2 AND2X2_3047 ( .A(core__abc_22172_new_n4792_), .B(core__abc_22172_new_n4804_), .Y(core__abc_22172_new_n4807_));
AND2X2 AND2X2_3048 ( .A(core__abc_22172_new_n4783_), .B(core__abc_22172_new_n4809_), .Y(core__abc_22172_new_n4810_));
AND2X2 AND2X2_3049 ( .A(core__abc_22172_new_n4811_), .B(core__abc_22172_new_n4812_), .Y(core__abc_22172_new_n4813_));
AND2X2 AND2X2_305 ( .A(_abc_19873_new_n916_), .B(core_key_87_), .Y(_abc_19873_new_n1422_));
AND2X2 AND2X2_3050 ( .A(core__abc_22172_new_n4816_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n4817_));
AND2X2 AND2X2_3051 ( .A(core__abc_22172_new_n4817_), .B(core__abc_22172_new_n4815_), .Y(core__abc_22172_new_n4818_));
AND2X2 AND2X2_3052 ( .A(core__abc_22172_new_n3214_), .B(core_key_90_), .Y(core__abc_22172_new_n4819_));
AND2X2 AND2X2_3053 ( .A(core_v3_reg_26_), .B(core_mi_26_), .Y(core__abc_22172_new_n4820_));
AND2X2 AND2X2_3054 ( .A(core__abc_22172_new_n4821_), .B(core__abc_22172_new_n4822_), .Y(core__abc_22172_new_n4823_));
AND2X2 AND2X2_3055 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n4823_), .Y(core__abc_22172_new_n4824_));
AND2X2 AND2X2_3056 ( .A(core__abc_22172_new_n4828_), .B(reset_n), .Y(core__abc_22172_new_n4829_));
AND2X2 AND2X2_3057 ( .A(core__abc_22172_new_n4827_), .B(core__abc_22172_new_n4829_), .Y(core__0v3_reg_63_0__26_));
AND2X2 AND2X2_3058 ( .A(core__abc_22172_new_n4811_), .B(core__abc_22172_new_n4831_), .Y(core__abc_22172_new_n4832_));
AND2X2 AND2X2_3059 ( .A(core__abc_22172_new_n4834_), .B(core__abc_22172_new_n2284_), .Y(core__abc_22172_new_n4835_));
AND2X2 AND2X2_306 ( .A(_abc_19873_new_n925_), .B(word2_reg_23_), .Y(_abc_19873_new_n1424_));
AND2X2 AND2X2_3060 ( .A(core__abc_22172_new_n4833_), .B(core__abc_22172_new_n2278_), .Y(core__abc_22172_new_n4836_));
AND2X2 AND2X2_3061 ( .A(core__abc_22172_new_n4839_), .B(core__abc_22172_new_n1741_), .Y(core__abc_22172_new_n4840_));
AND2X2 AND2X2_3062 ( .A(core__abc_22172_new_n4838_), .B(core__abc_22172_new_n1738_), .Y(core__abc_22172_new_n4841_));
AND2X2 AND2X2_3063 ( .A(core__abc_22172_new_n4842_), .B(core_v3_reg_11_), .Y(core__abc_22172_new_n4843_));
AND2X2 AND2X2_3064 ( .A(core__abc_22172_new_n4844_), .B(core__abc_22172_new_n4845_), .Y(core__abc_22172_new_n4846_));
AND2X2 AND2X2_3065 ( .A(core__abc_22172_new_n4837_), .B(core__abc_22172_new_n4846_), .Y(core__abc_22172_new_n4847_));
AND2X2 AND2X2_3066 ( .A(core__abc_22172_new_n4848_), .B(core__abc_22172_new_n4849_), .Y(core__abc_22172_new_n4850_));
AND2X2 AND2X2_3067 ( .A(core__abc_22172_new_n4832_), .B(core__abc_22172_new_n4851_), .Y(core__abc_22172_new_n4852_));
AND2X2 AND2X2_3068 ( .A(core__abc_22172_new_n4853_), .B(core__abc_22172_new_n4854_), .Y(core__abc_22172_new_n4855_));
AND2X2 AND2X2_3069 ( .A(core__abc_22172_new_n4858_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n4859_));
AND2X2 AND2X2_307 ( .A(_abc_19873_new_n907_), .B(word1_reg_23_), .Y(_abc_19873_new_n1425_));
AND2X2 AND2X2_3070 ( .A(core__abc_22172_new_n4859_), .B(core__abc_22172_new_n4856_), .Y(core__abc_22172_new_n4860_));
AND2X2 AND2X2_3071 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n4861_), .Y(core__abc_22172_new_n4862_));
AND2X2 AND2X2_3072 ( .A(core_v3_reg_27_), .B(core_mi_27_), .Y(core__abc_22172_new_n4863_));
AND2X2 AND2X2_3073 ( .A(core__abc_22172_new_n4864_), .B(core__abc_22172_new_n4865_), .Y(core__abc_22172_new_n4866_));
AND2X2 AND2X2_3074 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n4866_), .Y(core__abc_22172_new_n4867_));
AND2X2 AND2X2_3075 ( .A(core__abc_22172_new_n4871_), .B(reset_n), .Y(core__abc_22172_new_n4872_));
AND2X2 AND2X2_3076 ( .A(core__abc_22172_new_n4870_), .B(core__abc_22172_new_n4872_), .Y(core__0v3_reg_63_0__27_));
AND2X2 AND2X2_3077 ( .A(core__abc_22172_new_n3217_), .B(core_v3_reg_28_), .Y(core__abc_22172_new_n4874_));
AND2X2 AND2X2_3078 ( .A(core__abc_22172_new_n4875_), .B(core__abc_22172_new_n4876_), .Y(core__abc_22172_new_n4877_));
AND2X2 AND2X2_3079 ( .A(core__abc_22172_new_n4877_), .B(core__abc_22172_new_n4809_), .Y(core__abc_22172_new_n4878_));
AND2X2 AND2X2_308 ( .A(_abc_19873_new_n930_), .B(word0_reg_23_), .Y(_abc_19873_new_n1426_));
AND2X2 AND2X2_3080 ( .A(core__abc_22172_new_n4878_), .B(core__abc_22172_new_n4782_), .Y(core__abc_22172_new_n4879_));
AND2X2 AND2X2_3081 ( .A(core__abc_22172_new_n4875_), .B(core__abc_22172_new_n4806_), .Y(core__abc_22172_new_n4880_));
AND2X2 AND2X2_3082 ( .A(core__abc_22172_new_n4878_), .B(core__abc_22172_new_n4778_), .Y(core__abc_22172_new_n4883_));
AND2X2 AND2X2_3083 ( .A(core__abc_22172_new_n4676_), .B(core__abc_22172_new_n4883_), .Y(core__abc_22172_new_n4884_));
AND2X2 AND2X2_3084 ( .A(core__abc_22172_new_n2261_), .B(core__abc_22172_new_n2278_), .Y(core__abc_22172_new_n4886_));
AND2X2 AND2X2_3085 ( .A(core__abc_22172_new_n4784_), .B(core__abc_22172_new_n4886_), .Y(core__abc_22172_new_n4887_));
AND2X2 AND2X2_3086 ( .A(core__abc_22172_new_n4687_), .B(core__abc_22172_new_n4887_), .Y(core__abc_22172_new_n4888_));
AND2X2 AND2X2_3087 ( .A(core__abc_22172_new_n4787_), .B(core__abc_22172_new_n4886_), .Y(core__abc_22172_new_n4889_));
AND2X2 AND2X2_3088 ( .A(core__abc_22172_new_n2275_), .B(core__abc_22172_new_n2259_), .Y(core__abc_22172_new_n4890_));
AND2X2 AND2X2_3089 ( .A(core__abc_22172_new_n4893_), .B(core__abc_22172_new_n2295_), .Y(core__abc_22172_new_n4894_));
AND2X2 AND2X2_309 ( .A(_abc_19873_new_n912_), .B(word3_reg_23_), .Y(_abc_19873_new_n1430_));
AND2X2 AND2X2_3090 ( .A(core__abc_22172_new_n4896_), .B(core__abc_22172_new_n4897_), .Y(core__abc_22172_new_n4898_));
AND2X2 AND2X2_3091 ( .A(core__abc_22172_new_n4898_), .B(core__abc_22172_new_n2301_), .Y(core__abc_22172_new_n4899_));
AND2X2 AND2X2_3092 ( .A(core__abc_22172_new_n4696_), .B(core__abc_22172_new_n3105_), .Y(core__abc_22172_new_n4903_));
AND2X2 AND2X2_3093 ( .A(core__abc_22172_new_n4904_), .B(core__abc_22172_new_n1755_), .Y(core__abc_22172_new_n4905_));
AND2X2 AND2X2_3094 ( .A(core__abc_22172_new_n4906_), .B(core__abc_22172_new_n1758_), .Y(core__abc_22172_new_n4907_));
AND2X2 AND2X2_3095 ( .A(core__abc_22172_new_n4910_), .B(core__abc_22172_new_n4911_), .Y(core__abc_22172_new_n4912_));
AND2X2 AND2X2_3096 ( .A(core__abc_22172_new_n4901_), .B(core__abc_22172_new_n4913_), .Y(core__abc_22172_new_n4914_));
AND2X2 AND2X2_3097 ( .A(core__abc_22172_new_n4900_), .B(core__abc_22172_new_n4912_), .Y(core__abc_22172_new_n4915_));
AND2X2 AND2X2_3098 ( .A(core__abc_22172_new_n4885_), .B(core__abc_22172_new_n4917_), .Y(core__abc_22172_new_n4918_));
AND2X2 AND2X2_3099 ( .A(core__abc_22172_new_n4919_), .B(core__abc_22172_new_n4920_), .Y(core__abc_22172_new_n4921_));
AND2X2 AND2X2_31 ( .A(_abc_19873_new_n912_), .B(word3_reg_0_), .Y(_abc_19873_new_n913_));
AND2X2 AND2X2_310 ( .A(_abc_19873_new_n928_), .B(core_key_55_), .Y(_abc_19873_new_n1431_));
AND2X2 AND2X2_3100 ( .A(core__abc_22172_new_n4923_), .B(core__abc_22172_new_n4924_), .Y(core__abc_22172_new_n4925_));
AND2X2 AND2X2_3101 ( .A(core__abc_22172_new_n4925_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n4926_));
AND2X2 AND2X2_3102 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n4927_), .Y(core__abc_22172_new_n4928_));
AND2X2 AND2X2_3103 ( .A(core_v3_reg_28_), .B(core_mi_28_), .Y(core__abc_22172_new_n4930_));
AND2X2 AND2X2_3104 ( .A(core__abc_22172_new_n4931_), .B(core__abc_22172_new_n4929_), .Y(core__abc_22172_new_n4932_));
AND2X2 AND2X2_3105 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n4932_), .Y(core__abc_22172_new_n4933_));
AND2X2 AND2X2_3106 ( .A(core__abc_22172_new_n4935_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n4936_));
AND2X2 AND2X2_3107 ( .A(core__abc_22172_new_n4937_), .B(reset_n), .Y(core__0v3_reg_63_0__28_));
AND2X2 AND2X2_3108 ( .A(core__abc_22172_new_n4919_), .B(core__abc_22172_new_n4939_), .Y(core__abc_22172_new_n4940_));
AND2X2 AND2X2_3109 ( .A(core__abc_22172_new_n4943_), .B(core__abc_22172_new_n2318_), .Y(core__abc_22172_new_n4944_));
AND2X2 AND2X2_311 ( .A(_abc_19873_new_n901_), .B(core_key_23_), .Y(_abc_19873_new_n1432_));
AND2X2 AND2X2_3110 ( .A(core__abc_22172_new_n4942_), .B(core__abc_22172_new_n2312_), .Y(core__abc_22172_new_n4945_));
AND2X2 AND2X2_3111 ( .A(core__abc_22172_new_n4948_), .B(core__abc_22172_new_n1775_), .Y(core__abc_22172_new_n4949_));
AND2X2 AND2X2_3112 ( .A(core__abc_22172_new_n4947_), .B(core__abc_22172_new_n1772_), .Y(core__abc_22172_new_n4950_));
AND2X2 AND2X2_3113 ( .A(core__abc_22172_new_n4951_), .B(core_v3_reg_13_), .Y(core__abc_22172_new_n4952_));
AND2X2 AND2X2_3114 ( .A(core__abc_22172_new_n4953_), .B(core__abc_22172_new_n4954_), .Y(core__abc_22172_new_n4955_));
AND2X2 AND2X2_3115 ( .A(core__abc_22172_new_n4946_), .B(core__abc_22172_new_n4955_), .Y(core__abc_22172_new_n4956_));
AND2X2 AND2X2_3116 ( .A(core__abc_22172_new_n4958_), .B(core__abc_22172_new_n4959_), .Y(core__abc_22172_new_n4960_));
AND2X2 AND2X2_3117 ( .A(core__abc_22172_new_n4961_), .B(core__abc_22172_new_n4957_), .Y(core__abc_22172_new_n4962_));
AND2X2 AND2X2_3118 ( .A(core__abc_22172_new_n4941_), .B(core__abc_22172_new_n4963_), .Y(core__abc_22172_new_n4964_));
AND2X2 AND2X2_3119 ( .A(core__abc_22172_new_n4940_), .B(core__abc_22172_new_n4962_), .Y(core__abc_22172_new_n4965_));
AND2X2 AND2X2_312 ( .A(_abc_19873_new_n888_), .B(core_mi_23_), .Y(_abc_19873_new_n1434_));
AND2X2 AND2X2_3120 ( .A(core__abc_22172_new_n4969_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n4970_));
AND2X2 AND2X2_3121 ( .A(core__abc_22172_new_n4970_), .B(core__abc_22172_new_n4967_), .Y(core__abc_22172_new_n4971_));
AND2X2 AND2X2_3122 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n4972_), .Y(core__abc_22172_new_n4973_));
AND2X2 AND2X2_3123 ( .A(core_v3_reg_29_), .B(core_mi_29_), .Y(core__abc_22172_new_n4974_));
AND2X2 AND2X2_3124 ( .A(core__abc_22172_new_n4975_), .B(core__abc_22172_new_n4976_), .Y(core__abc_22172_new_n4977_));
AND2X2 AND2X2_3125 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n4977_), .Y(core__abc_22172_new_n4978_));
AND2X2 AND2X2_3126 ( .A(core__abc_22172_new_n4982_), .B(reset_n), .Y(core__abc_22172_new_n4983_));
AND2X2 AND2X2_3127 ( .A(core__abc_22172_new_n4981_), .B(core__abc_22172_new_n4983_), .Y(core__0v3_reg_63_0__29_));
AND2X2 AND2X2_3128 ( .A(core__abc_22172_new_n2295_), .B(core__abc_22172_new_n2312_), .Y(core__abc_22172_new_n4985_));
AND2X2 AND2X2_3129 ( .A(core__abc_22172_new_n4893_), .B(core__abc_22172_new_n4985_), .Y(core__abc_22172_new_n4986_));
AND2X2 AND2X2_313 ( .A(_abc_19873_new_n919_), .B(core_mi_55_), .Y(_abc_19873_new_n1435_));
AND2X2 AND2X2_3130 ( .A(core__abc_22172_new_n2312_), .B(core__abc_22172_new_n2293_), .Y(core__abc_22172_new_n4987_));
AND2X2 AND2X2_3131 ( .A(core__abc_22172_new_n4989_), .B(core__abc_22172_new_n2329_), .Y(core__abc_22172_new_n4990_));
AND2X2 AND2X2_3132 ( .A(core__abc_22172_new_n4992_), .B(core__abc_22172_new_n4993_), .Y(core__abc_22172_new_n4994_));
AND2X2 AND2X2_3133 ( .A(core__abc_22172_new_n4994_), .B(core__abc_22172_new_n2335_), .Y(core__abc_22172_new_n4995_));
AND2X2 AND2X2_3134 ( .A(core__abc_22172_new_n4904_), .B(core__abc_22172_new_n3101_), .Y(core__abc_22172_new_n4998_));
AND2X2 AND2X2_3135 ( .A(core__abc_22172_new_n4999_), .B(core__abc_22172_new_n1789_), .Y(core__abc_22172_new_n5000_));
AND2X2 AND2X2_3136 ( .A(core__abc_22172_new_n5001_), .B(core__abc_22172_new_n1792_), .Y(core__abc_22172_new_n5002_));
AND2X2 AND2X2_3137 ( .A(core__abc_22172_new_n5005_), .B(core__abc_22172_new_n5006_), .Y(core__abc_22172_new_n5007_));
AND2X2 AND2X2_3138 ( .A(core__abc_22172_new_n4996_), .B(core__abc_22172_new_n5007_), .Y(core__abc_22172_new_n5008_));
AND2X2 AND2X2_3139 ( .A(core__abc_22172_new_n5009_), .B(core__abc_22172_new_n5010_), .Y(core__abc_22172_new_n5011_));
AND2X2 AND2X2_314 ( .A(_abc_19873_new_n1439_), .B(_abc_19873_new_n937_), .Y(\read_data[23] ));
AND2X2 AND2X2_3140 ( .A(core__abc_22172_new_n4961_), .B(core__abc_22172_new_n4939_), .Y(core__abc_22172_new_n5014_));
AND2X2 AND2X2_3141 ( .A(core__abc_22172_new_n4919_), .B(core__abc_22172_new_n5014_), .Y(core__abc_22172_new_n5015_));
AND2X2 AND2X2_3142 ( .A(core__abc_22172_new_n5017_), .B(core__abc_22172_new_n5013_), .Y(core__abc_22172_new_n5018_));
AND2X2 AND2X2_3143 ( .A(core__abc_22172_new_n5016_), .B(core__abc_22172_new_n5012_), .Y(core__abc_22172_new_n5019_));
AND2X2 AND2X2_3144 ( .A(core__abc_22172_new_n5023_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n5024_));
AND2X2 AND2X2_3145 ( .A(core__abc_22172_new_n5024_), .B(core__abc_22172_new_n5021_), .Y(core__abc_22172_new_n5025_));
AND2X2 AND2X2_3146 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n5026_), .Y(core__abc_22172_new_n5027_));
AND2X2 AND2X2_3147 ( .A(core_v3_reg_30_), .B(core_mi_30_), .Y(core__abc_22172_new_n5028_));
AND2X2 AND2X2_3148 ( .A(core__abc_22172_new_n5029_), .B(core__abc_22172_new_n5030_), .Y(core__abc_22172_new_n5031_));
AND2X2 AND2X2_3149 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n5031_), .Y(core__abc_22172_new_n5032_));
AND2X2 AND2X2_315 ( .A(_abc_19873_new_n881_), .B(core_key_120_), .Y(_abc_19873_new_n1441_));
AND2X2 AND2X2_3150 ( .A(core__abc_22172_new_n5036_), .B(reset_n), .Y(core__abc_22172_new_n5037_));
AND2X2 AND2X2_3151 ( .A(core__abc_22172_new_n5035_), .B(core__abc_22172_new_n5037_), .Y(core__0v3_reg_63_0__30_));
AND2X2 AND2X2_3152 ( .A(core__abc_22172_new_n5042_), .B(core__abc_22172_new_n2328_), .Y(core__abc_22172_new_n5043_));
AND2X2 AND2X2_3153 ( .A(core__abc_22172_new_n5044_), .B(core__abc_22172_new_n5041_), .Y(core__abc_22172_new_n5045_));
AND2X2 AND2X2_3154 ( .A(core__abc_22172_new_n5047_), .B(core__abc_22172_new_n1809_), .Y(core__abc_22172_new_n5048_));
AND2X2 AND2X2_3155 ( .A(core__abc_22172_new_n5046_), .B(core__abc_22172_new_n1806_), .Y(core__abc_22172_new_n5049_));
AND2X2 AND2X2_3156 ( .A(core__abc_22172_new_n5050_), .B(core_v3_reg_15_), .Y(core__abc_22172_new_n5051_));
AND2X2 AND2X2_3157 ( .A(core__abc_22172_new_n5053_), .B(core__abc_22172_new_n5052_), .Y(core__abc_22172_new_n5054_));
AND2X2 AND2X2_3158 ( .A(core__abc_22172_new_n5043_), .B(core__abc_22172_new_n2347_), .Y(core__abc_22172_new_n5057_));
AND2X2 AND2X2_3159 ( .A(core__abc_22172_new_n5040_), .B(core__abc_22172_new_n2348_), .Y(core__abc_22172_new_n5058_));
AND2X2 AND2X2_316 ( .A(_abc_19873_new_n888_), .B(core_mi_24_), .Y(_abc_19873_new_n1442_));
AND2X2 AND2X2_3160 ( .A(core__abc_22172_new_n5060_), .B(core__abc_22172_new_n5061_), .Y(core__abc_22172_new_n5062_));
AND2X2 AND2X2_3161 ( .A(core__abc_22172_new_n5056_), .B(core__abc_22172_new_n5063_), .Y(core__abc_22172_new_n5064_));
AND2X2 AND2X2_3162 ( .A(core__abc_22172_new_n5039_), .B(core__abc_22172_new_n5064_), .Y(core__abc_22172_new_n5065_));
AND2X2 AND2X2_3163 ( .A(core__abc_22172_new_n5066_), .B(core__abc_22172_new_n5067_), .Y(core__abc_22172_new_n5068_));
AND2X2 AND2X2_3164 ( .A(core__abc_22172_new_n5071_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n5072_));
AND2X2 AND2X2_3165 ( .A(core__abc_22172_new_n5072_), .B(core__abc_22172_new_n5069_), .Y(core__abc_22172_new_n5073_));
AND2X2 AND2X2_3166 ( .A(core__abc_22172_new_n3214_), .B(core_key_95_), .Y(core__abc_22172_new_n5074_));
AND2X2 AND2X2_3167 ( .A(core_v3_reg_31_), .B(core_mi_31_), .Y(core__abc_22172_new_n5075_));
AND2X2 AND2X2_3168 ( .A(core__abc_22172_new_n5076_), .B(core__abc_22172_new_n5077_), .Y(core__abc_22172_new_n5078_));
AND2X2 AND2X2_3169 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n5078_), .Y(core__abc_22172_new_n5079_));
AND2X2 AND2X2_317 ( .A(_abc_19873_new_n916_), .B(core_key_88_), .Y(_abc_19873_new_n1444_));
AND2X2 AND2X2_3170 ( .A(core__abc_22172_new_n5083_), .B(reset_n), .Y(core__abc_22172_new_n5084_));
AND2X2 AND2X2_3171 ( .A(core__abc_22172_new_n5082_), .B(core__abc_22172_new_n5084_), .Y(core__0v3_reg_63_0__31_));
AND2X2 AND2X2_3172 ( .A(core__abc_22172_new_n3217_), .B(core_v3_reg_32_), .Y(core__abc_22172_new_n5086_));
AND2X2 AND2X2_3173 ( .A(core__abc_22172_new_n4962_), .B(core__abc_22172_new_n4917_), .Y(core__abc_22172_new_n5087_));
AND2X2 AND2X2_3174 ( .A(core__abc_22172_new_n5064_), .B(core__abc_22172_new_n5013_), .Y(core__abc_22172_new_n5088_));
AND2X2 AND2X2_3175 ( .A(core__abc_22172_new_n5088_), .B(core__abc_22172_new_n5087_), .Y(core__abc_22172_new_n5089_));
AND2X2 AND2X2_3176 ( .A(core__abc_22172_new_n5089_), .B(core__abc_22172_new_n4883_), .Y(core__abc_22172_new_n5090_));
AND2X2 AND2X2_3177 ( .A(core__abc_22172_new_n5090_), .B(core__abc_22172_new_n4674_), .Y(core__abc_22172_new_n5091_));
AND2X2 AND2X2_3178 ( .A(core__abc_22172_new_n5091_), .B(core__abc_22172_new_n4199_), .Y(core__abc_22172_new_n5092_));
AND2X2 AND2X2_3179 ( .A(core__abc_22172_new_n5090_), .B(core__abc_22172_new_n4673_), .Y(core__abc_22172_new_n5093_));
AND2X2 AND2X2_318 ( .A(_abc_19873_new_n925_), .B(word2_reg_24_), .Y(_abc_19873_new_n1447_));
AND2X2 AND2X2_3180 ( .A(core__abc_22172_new_n5089_), .B(core__abc_22172_new_n4882_), .Y(core__abc_22172_new_n5094_));
AND2X2 AND2X2_3181 ( .A(core__abc_22172_new_n5095_), .B(core__abc_22172_new_n4957_), .Y(core__abc_22172_new_n5096_));
AND2X2 AND2X2_3182 ( .A(core__abc_22172_new_n5088_), .B(core__abc_22172_new_n5096_), .Y(core__abc_22172_new_n5097_));
AND2X2 AND2X2_3183 ( .A(core__abc_22172_new_n5045_), .B(core__abc_22172_new_n5055_), .Y(core__abc_22172_new_n5098_));
AND2X2 AND2X2_3184 ( .A(core__abc_22172_new_n5099_), .B(core__abc_22172_new_n5056_), .Y(core__abc_22172_new_n5100_));
AND2X2 AND2X2_3185 ( .A(core__abc_22172_new_n5106_), .B(core__abc_22172_new_n1826_), .Y(core__abc_22172_new_n5107_));
AND2X2 AND2X2_3186 ( .A(core__abc_22172_new_n3153_), .B(core__abc_22172_new_n1823_), .Y(core__abc_22172_new_n5108_));
AND2X2 AND2X2_3187 ( .A(core__abc_22172_new_n5111_), .B(core__abc_22172_new_n5112_), .Y(core__abc_22172_new_n5113_));
AND2X2 AND2X2_3188 ( .A(core__abc_22172_new_n5114_), .B(core__abc_22172_new_n1260_), .Y(core__abc_22172_new_n5115_));
AND2X2 AND2X2_3189 ( .A(core__abc_22172_new_n5113_), .B(core__abc_22172_new_n1268_), .Y(core__abc_22172_new_n5116_));
AND2X2 AND2X2_319 ( .A(_abc_19873_new_n907_), .B(word1_reg_24_), .Y(_abc_19873_new_n1448_));
AND2X2 AND2X2_3190 ( .A(core__abc_22172_new_n5104_), .B(core__abc_22172_new_n5118_), .Y(core__abc_22172_new_n5119_));
AND2X2 AND2X2_3191 ( .A(core__abc_22172_new_n5124_), .B(core__abc_22172_new_n5125_), .Y(core__abc_22172_new_n5126_));
AND2X2 AND2X2_3192 ( .A(core__abc_22172_new_n5059_), .B(core__abc_22172_new_n5062_), .Y(core__abc_22172_new_n5128_));
AND2X2 AND2X2_3193 ( .A(core__abc_22172_new_n5134_), .B(core__abc_22172_new_n5135_), .Y(core__abc_22172_new_n5136_));
AND2X2 AND2X2_3194 ( .A(core__abc_22172_new_n5132_), .B(core__abc_22172_new_n5136_), .Y(core__abc_22172_new_n5137_));
AND2X2 AND2X2_3195 ( .A(core__abc_22172_new_n5121_), .B(core__abc_22172_new_n5137_), .Y(core__abc_22172_new_n5138_));
AND2X2 AND2X2_3196 ( .A(core__abc_22172_new_n5120_), .B(core__abc_22172_new_n5138_), .Y(core__abc_22172_new_n5139_));
AND2X2 AND2X2_3197 ( .A(core__abc_22172_new_n5139_), .B(core__abc_22172_new_n5117_), .Y(core__abc_22172_new_n5140_));
AND2X2 AND2X2_3198 ( .A(core__abc_22172_new_n5141_), .B(core__abc_22172_new_n3886_), .Y(core__abc_22172_new_n5142_));
AND2X2 AND2X2_3199 ( .A(core__abc_22172_new_n5143_), .B(core__abc_22172_new_n3885_), .Y(core__abc_22172_new_n5144_));
AND2X2 AND2X2_32 ( .A(_abc_19873_new_n883_), .B(\addr[1] ), .Y(_abc_19873_new_n914_));
AND2X2 AND2X2_320 ( .A(_abc_19873_new_n912_), .B(word3_reg_24_), .Y(_abc_19873_new_n1449_));
AND2X2 AND2X2_3200 ( .A(core__abc_22172_new_n5145_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n5146_));
AND2X2 AND2X2_3201 ( .A(core__abc_22172_new_n3214_), .B(core_key_96_), .Y(core__abc_22172_new_n5147_));
AND2X2 AND2X2_3202 ( .A(core_v3_reg_32_), .B(core_mi_32_), .Y(core__abc_22172_new_n5149_));
AND2X2 AND2X2_3203 ( .A(core__abc_22172_new_n5150_), .B(core__abc_22172_new_n5148_), .Y(core__abc_22172_new_n5151_));
AND2X2 AND2X2_3204 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n5151_), .Y(core__abc_22172_new_n5152_));
AND2X2 AND2X2_3205 ( .A(core__abc_22172_new_n5154_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n5155_));
AND2X2 AND2X2_3206 ( .A(core__abc_22172_new_n5156_), .B(reset_n), .Y(core__0v3_reg_63_0__32_));
AND2X2 AND2X2_3207 ( .A(core__abc_22172_new_n3217_), .B(core_v3_reg_33_), .Y(core__abc_22172_new_n5158_));
AND2X2 AND2X2_3208 ( .A(core__abc_22172_new_n1289_), .B(core__abc_22172_new_n1259_), .Y(core__abc_22172_new_n5161_));
AND2X2 AND2X2_3209 ( .A(core__abc_22172_new_n5165_), .B(core__abc_22172_new_n1843_), .Y(core__abc_22172_new_n5166_));
AND2X2 AND2X2_321 ( .A(_abc_19873_new_n919_), .B(core_mi_56_), .Y(_abc_19873_new_n1452_));
AND2X2 AND2X2_3210 ( .A(core__abc_22172_new_n5164_), .B(core__abc_22172_new_n1840_), .Y(core__abc_22172_new_n5167_));
AND2X2 AND2X2_3211 ( .A(core__abc_22172_new_n5168_), .B(core_v3_reg_17_), .Y(core__abc_22172_new_n5169_));
AND2X2 AND2X2_3212 ( .A(core__abc_22172_new_n5170_), .B(core__abc_22172_new_n5171_), .Y(core__abc_22172_new_n5172_));
AND2X2 AND2X2_3213 ( .A(core__abc_22172_new_n5173_), .B(core__abc_22172_new_n5163_), .Y(core__abc_22172_new_n5174_));
AND2X2 AND2X2_3214 ( .A(core__abc_22172_new_n5172_), .B(core__abc_22172_new_n5162_), .Y(core__abc_22172_new_n5176_));
AND2X2 AND2X2_3215 ( .A(core__abc_22172_new_n5175_), .B(core__abc_22172_new_n5177_), .Y(core__abc_22172_new_n5178_));
AND2X2 AND2X2_3216 ( .A(core__abc_22172_new_n5180_), .B(core__abc_22172_new_n5181_), .Y(core__abc_22172_new_n5182_));
AND2X2 AND2X2_3217 ( .A(core__abc_22172_new_n5183_), .B(core__abc_22172_new_n3960_), .Y(core__abc_22172_new_n5184_));
AND2X2 AND2X2_3218 ( .A(core__abc_22172_new_n5182_), .B(core__abc_22172_new_n3957_), .Y(core__abc_22172_new_n5185_));
AND2X2 AND2X2_3219 ( .A(core__abc_22172_new_n5186_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n5187_));
AND2X2 AND2X2_322 ( .A(_abc_19873_new_n930_), .B(word0_reg_24_), .Y(_abc_19873_new_n1453_));
AND2X2 AND2X2_3220 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n5188_), .Y(core__abc_22172_new_n5189_));
AND2X2 AND2X2_3221 ( .A(core_v3_reg_33_), .B(core_mi_33_), .Y(core__abc_22172_new_n5191_));
AND2X2 AND2X2_3222 ( .A(core__abc_22172_new_n5192_), .B(core__abc_22172_new_n5190_), .Y(core__abc_22172_new_n5193_));
AND2X2 AND2X2_3223 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n5193_), .Y(core__abc_22172_new_n5194_));
AND2X2 AND2X2_3224 ( .A(core__abc_22172_new_n5196_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n5197_));
AND2X2 AND2X2_3225 ( .A(core__abc_22172_new_n5198_), .B(reset_n), .Y(core__0v3_reg_63_0__33_));
AND2X2 AND2X2_3226 ( .A(core__abc_22172_new_n3217_), .B(core_v3_reg_34_), .Y(core__abc_22172_new_n5200_));
AND2X2 AND2X2_3227 ( .A(core__abc_22172_new_n5201_), .B(core__abc_22172_new_n5177_), .Y(core__abc_22172_new_n5202_));
AND2X2 AND2X2_3228 ( .A(core__abc_22172_new_n5178_), .B(core__abc_22172_new_n5118_), .Y(core__abc_22172_new_n5203_));
AND2X2 AND2X2_3229 ( .A(core__abc_22172_new_n5104_), .B(core__abc_22172_new_n5203_), .Y(core__abc_22172_new_n5204_));
AND2X2 AND2X2_323 ( .A(_abc_19873_new_n928_), .B(core_key_56_), .Y(_abc_19873_new_n1455_));
AND2X2 AND2X2_3230 ( .A(core__abc_22172_new_n2919_), .B(core__abc_22172_new_n1299_), .Y(core__abc_22172_new_n5206_));
AND2X2 AND2X2_3231 ( .A(core__abc_22172_new_n3016_), .B(core__abc_22172_new_n1300_), .Y(core__abc_22172_new_n5207_));
AND2X2 AND2X2_3232 ( .A(core__abc_22172_new_n5212_), .B(core__abc_22172_new_n3164_), .Y(core__abc_22172_new_n5213_));
AND2X2 AND2X2_3233 ( .A(core__abc_22172_new_n5214_), .B(core__abc_22172_new_n1857_), .Y(core__abc_22172_new_n5215_));
AND2X2 AND2X2_3234 ( .A(core__abc_22172_new_n5213_), .B(core__abc_22172_new_n1860_), .Y(core__abc_22172_new_n5216_));
AND2X2 AND2X2_3235 ( .A(core__abc_22172_new_n5219_), .B(core__abc_22172_new_n5220_), .Y(core__abc_22172_new_n5221_));
AND2X2 AND2X2_3236 ( .A(core__abc_22172_new_n5222_), .B(core__abc_22172_new_n5209_), .Y(core__abc_22172_new_n5223_));
AND2X2 AND2X2_3237 ( .A(core__abc_22172_new_n5221_), .B(core__abc_22172_new_n5208_), .Y(core__abc_22172_new_n5224_));
AND2X2 AND2X2_3238 ( .A(core__abc_22172_new_n5205_), .B(core__abc_22172_new_n5226_), .Y(core__abc_22172_new_n5227_));
AND2X2 AND2X2_3239 ( .A(core__abc_22172_new_n5228_), .B(core__abc_22172_new_n5229_), .Y(core__abc_22172_new_n5230_));
AND2X2 AND2X2_324 ( .A(_abc_19873_new_n901_), .B(core_key_24_), .Y(_abc_19873_new_n1456_));
AND2X2 AND2X2_3240 ( .A(core__abc_22172_new_n5232_), .B(core__abc_22172_new_n5233_), .Y(core__abc_22172_new_n5234_));
AND2X2 AND2X2_3241 ( .A(core__abc_22172_new_n5234_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n5235_));
AND2X2 AND2X2_3242 ( .A(core__abc_22172_new_n3214_), .B(core_key_98_), .Y(core__abc_22172_new_n5236_));
AND2X2 AND2X2_3243 ( .A(core_v3_reg_34_), .B(core_mi_34_), .Y(core__abc_22172_new_n5238_));
AND2X2 AND2X2_3244 ( .A(core__abc_22172_new_n5239_), .B(core__abc_22172_new_n5237_), .Y(core__abc_22172_new_n5240_));
AND2X2 AND2X2_3245 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n5240_), .Y(core__abc_22172_new_n5241_));
AND2X2 AND2X2_3246 ( .A(core__abc_22172_new_n5243_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n5244_));
AND2X2 AND2X2_3247 ( .A(core__abc_22172_new_n5245_), .B(reset_n), .Y(core__0v3_reg_63_0__34_));
AND2X2 AND2X2_3248 ( .A(core__abc_22172_new_n5228_), .B(core__abc_22172_new_n5248_), .Y(core__abc_22172_new_n5249_));
AND2X2 AND2X2_3249 ( .A(core__abc_22172_new_n5251_), .B(core__abc_22172_new_n1325_), .Y(core__abc_22172_new_n5252_));
AND2X2 AND2X2_325 ( .A(_abc_19873_new_n1460_), .B(_abc_19873_new_n937_), .Y(\read_data[24] ));
AND2X2 AND2X2_3250 ( .A(core__abc_22172_new_n5250_), .B(core__abc_22172_new_n1317_), .Y(core__abc_22172_new_n5253_));
AND2X2 AND2X2_3251 ( .A(core__abc_22172_new_n5255_), .B(core__abc_22172_new_n1874_), .Y(core__abc_22172_new_n5257_));
AND2X2 AND2X2_3252 ( .A(core__abc_22172_new_n5258_), .B(core__abc_22172_new_n5256_), .Y(core__abc_22172_new_n5259_));
AND2X2 AND2X2_3253 ( .A(core__abc_22172_new_n5260_), .B(core_v3_reg_19_), .Y(core__abc_22172_new_n5261_));
AND2X2 AND2X2_3254 ( .A(core__abc_22172_new_n5262_), .B(core__abc_22172_new_n5263_), .Y(core__abc_22172_new_n5264_));
AND2X2 AND2X2_3255 ( .A(core__abc_22172_new_n5264_), .B(core__abc_22172_new_n5254_), .Y(core__abc_22172_new_n5267_));
AND2X2 AND2X2_3256 ( .A(core__abc_22172_new_n5271_), .B(core__abc_22172_new_n5265_), .Y(core__abc_22172_new_n5272_));
AND2X2 AND2X2_3257 ( .A(core__abc_22172_new_n5273_), .B(core__abc_22172_new_n5269_), .Y(core__abc_22172_new_n5274_));
AND2X2 AND2X2_3258 ( .A(core__abc_22172_new_n5277_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n5278_));
AND2X2 AND2X2_3259 ( .A(core__abc_22172_new_n5278_), .B(core__abc_22172_new_n5275_), .Y(core__abc_22172_new_n5279_));
AND2X2 AND2X2_326 ( .A(_abc_19873_new_n881_), .B(core_key_121_), .Y(_abc_19873_new_n1462_));
AND2X2 AND2X2_3260 ( .A(core__abc_22172_new_n3214_), .B(core_key_99_), .Y(core__abc_22172_new_n5280_));
AND2X2 AND2X2_3261 ( .A(core_v3_reg_35_), .B(core_mi_35_), .Y(core__abc_22172_new_n5281_));
AND2X2 AND2X2_3262 ( .A(core__abc_22172_new_n5282_), .B(core__abc_22172_new_n5283_), .Y(core__abc_22172_new_n5284_));
AND2X2 AND2X2_3263 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n5284_), .Y(core__abc_22172_new_n5285_));
AND2X2 AND2X2_3264 ( .A(core__abc_22172_new_n5289_), .B(reset_n), .Y(core__abc_22172_new_n5290_));
AND2X2 AND2X2_3265 ( .A(core__abc_22172_new_n5288_), .B(core__abc_22172_new_n5290_), .Y(core__0v3_reg_63_0__35_));
AND2X2 AND2X2_3266 ( .A(core__abc_22172_new_n3217_), .B(core_v3_reg_36_), .Y(core__abc_22172_new_n5292_));
AND2X2 AND2X2_3267 ( .A(core__abc_22172_new_n5272_), .B(core__abc_22172_new_n5226_), .Y(core__abc_22172_new_n5293_));
AND2X2 AND2X2_3268 ( .A(core__abc_22172_new_n5293_), .B(core__abc_22172_new_n5202_), .Y(core__abc_22172_new_n5294_));
AND2X2 AND2X2_3269 ( .A(core__abc_22172_new_n5295_), .B(core__abc_22172_new_n5265_), .Y(core__abc_22172_new_n5296_));
AND2X2 AND2X2_327 ( .A(_abc_19873_new_n888_), .B(core_mi_25_), .Y(_abc_19873_new_n1463_));
AND2X2 AND2X2_3270 ( .A(core__abc_22172_new_n5293_), .B(core__abc_22172_new_n5203_), .Y(core__abc_22172_new_n5299_));
AND2X2 AND2X2_3271 ( .A(core__abc_22172_new_n5104_), .B(core__abc_22172_new_n5299_), .Y(core__abc_22172_new_n5300_));
AND2X2 AND2X2_3272 ( .A(core__abc_22172_new_n2924_), .B(core__abc_22172_new_n1335_), .Y(core__abc_22172_new_n5302_));
AND2X2 AND2X2_3273 ( .A(core__abc_22172_new_n3020_), .B(core__abc_22172_new_n1343_), .Y(core__abc_22172_new_n5303_));
AND2X2 AND2X2_3274 ( .A(core__abc_22172_new_n3153_), .B(core__abc_22172_new_n3159_), .Y(core__abc_22172_new_n5307_));
AND2X2 AND2X2_3275 ( .A(core__abc_22172_new_n5308_), .B(core__abc_22172_new_n1891_), .Y(core__abc_22172_new_n5309_));
AND2X2 AND2X2_3276 ( .A(core__abc_22172_new_n5310_), .B(core__abc_22172_new_n1894_), .Y(core__abc_22172_new_n5311_));
AND2X2 AND2X2_3277 ( .A(core__abc_22172_new_n5314_), .B(core__abc_22172_new_n5315_), .Y(core__abc_22172_new_n5316_));
AND2X2 AND2X2_3278 ( .A(core__abc_22172_new_n5317_), .B(core__abc_22172_new_n5305_), .Y(core__abc_22172_new_n5318_));
AND2X2 AND2X2_3279 ( .A(core__abc_22172_new_n5316_), .B(core__abc_22172_new_n5304_), .Y(core__abc_22172_new_n5319_));
AND2X2 AND2X2_328 ( .A(_abc_19873_new_n916_), .B(core_key_89_), .Y(_abc_19873_new_n1465_));
AND2X2 AND2X2_3280 ( .A(core__abc_22172_new_n5301_), .B(core__abc_22172_new_n5321_), .Y(core__abc_22172_new_n5322_));
AND2X2 AND2X2_3281 ( .A(core__abc_22172_new_n5323_), .B(core__abc_22172_new_n5324_), .Y(core__abc_22172_new_n5325_));
AND2X2 AND2X2_3282 ( .A(core__abc_22172_new_n5328_), .B(core__abc_22172_new_n5326_), .Y(core__abc_22172_new_n5329_));
AND2X2 AND2X2_3283 ( .A(core__abc_22172_new_n5329_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n5330_));
AND2X2 AND2X2_3284 ( .A(core__abc_22172_new_n3214_), .B(core_key_100_), .Y(core__abc_22172_new_n5331_));
AND2X2 AND2X2_3285 ( .A(core_v3_reg_36_), .B(core_mi_36_), .Y(core__abc_22172_new_n5333_));
AND2X2 AND2X2_3286 ( .A(core__abc_22172_new_n5334_), .B(core__abc_22172_new_n5332_), .Y(core__abc_22172_new_n5335_));
AND2X2 AND2X2_3287 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n5335_), .Y(core__abc_22172_new_n5336_));
AND2X2 AND2X2_3288 ( .A(core__abc_22172_new_n5338_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n5339_));
AND2X2 AND2X2_3289 ( .A(core__abc_22172_new_n5340_), .B(reset_n), .Y(core__0v3_reg_63_0__36_));
AND2X2 AND2X2_329 ( .A(_abc_19873_new_n925_), .B(word2_reg_25_), .Y(_abc_19873_new_n1468_));
AND2X2 AND2X2_3290 ( .A(core__abc_22172_new_n3217_), .B(core_v3_reg_37_), .Y(core__abc_22172_new_n5342_));
AND2X2 AND2X2_3291 ( .A(core__abc_22172_new_n5345_), .B(core__abc_22172_new_n1362_), .Y(core__abc_22172_new_n5346_));
AND2X2 AND2X2_3292 ( .A(core__abc_22172_new_n5344_), .B(core__abc_22172_new_n1353_), .Y(core__abc_22172_new_n5347_));
AND2X2 AND2X2_3293 ( .A(core__abc_22172_new_n5350_), .B(core__abc_22172_new_n1911_), .Y(core__abc_22172_new_n5351_));
AND2X2 AND2X2_3294 ( .A(core__abc_22172_new_n5349_), .B(core__abc_22172_new_n1908_), .Y(core__abc_22172_new_n5352_));
AND2X2 AND2X2_3295 ( .A(core__abc_22172_new_n5353_), .B(core_v3_reg_21_), .Y(core__abc_22172_new_n5354_));
AND2X2 AND2X2_3296 ( .A(core__abc_22172_new_n5355_), .B(core__abc_22172_new_n5356_), .Y(core__abc_22172_new_n5357_));
AND2X2 AND2X2_3297 ( .A(core__abc_22172_new_n5357_), .B(core__abc_22172_new_n5348_), .Y(core__abc_22172_new_n5358_));
AND2X2 AND2X2_3298 ( .A(core__abc_22172_new_n5361_), .B(core__abc_22172_new_n5343_), .Y(core__abc_22172_new_n5362_));
AND2X2 AND2X2_3299 ( .A(core__abc_22172_new_n5323_), .B(core__abc_22172_new_n5362_), .Y(core__abc_22172_new_n5363_));
AND2X2 AND2X2_33 ( .A(_abc_19873_new_n879_), .B(_abc_19873_new_n914_), .Y(_abc_19873_new_n915_));
AND2X2 AND2X2_330 ( .A(_abc_19873_new_n907_), .B(word1_reg_25_), .Y(_abc_19873_new_n1469_));
AND2X2 AND2X2_3300 ( .A(core__abc_22172_new_n5365_), .B(core__abc_22172_new_n5318_), .Y(core__abc_22172_new_n5366_));
AND2X2 AND2X2_3301 ( .A(core__abc_22172_new_n5365_), .B(core__abc_22172_new_n5321_), .Y(core__abc_22172_new_n5368_));
AND2X2 AND2X2_3302 ( .A(core__abc_22172_new_n5301_), .B(core__abc_22172_new_n5368_), .Y(core__abc_22172_new_n5369_));
AND2X2 AND2X2_3303 ( .A(core__abc_22172_new_n5370_), .B(core__abc_22172_new_n5367_), .Y(core__abc_22172_new_n5371_));
AND2X2 AND2X2_3304 ( .A(core__abc_22172_new_n5364_), .B(core__abc_22172_new_n5371_), .Y(core__abc_22172_new_n5372_));
AND2X2 AND2X2_3305 ( .A(core__abc_22172_new_n5372_), .B(core__abc_22172_new_n4229_), .Y(core__abc_22172_new_n5373_));
AND2X2 AND2X2_3306 ( .A(core__abc_22172_new_n5374_), .B(core__abc_22172_new_n4228_), .Y(core__abc_22172_new_n5375_));
AND2X2 AND2X2_3307 ( .A(core__abc_22172_new_n5376_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n5377_));
AND2X2 AND2X2_3308 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n5378_), .Y(core__abc_22172_new_n5379_));
AND2X2 AND2X2_3309 ( .A(core_v3_reg_37_), .B(core_mi_37_), .Y(core__abc_22172_new_n5381_));
AND2X2 AND2X2_331 ( .A(_abc_19873_new_n912_), .B(word3_reg_25_), .Y(_abc_19873_new_n1470_));
AND2X2 AND2X2_3310 ( .A(core__abc_22172_new_n5382_), .B(core__abc_22172_new_n5380_), .Y(core__abc_22172_new_n5383_));
AND2X2 AND2X2_3311 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n5383_), .Y(core__abc_22172_new_n5384_));
AND2X2 AND2X2_3312 ( .A(core__abc_22172_new_n5386_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n5387_));
AND2X2 AND2X2_3313 ( .A(core__abc_22172_new_n5388_), .B(reset_n), .Y(core__0v3_reg_63_0__37_));
AND2X2 AND2X2_3314 ( .A(core__abc_22172_new_n3217_), .B(core_v3_reg_38_), .Y(core__abc_22172_new_n5390_));
AND2X2 AND2X2_3315 ( .A(core__abc_22172_new_n5370_), .B(core__abc_22172_new_n5392_), .Y(core__abc_22172_new_n5393_));
AND2X2 AND2X2_3316 ( .A(core__abc_22172_new_n2924_), .B(core__abc_22172_new_n2926_), .Y(core__abc_22172_new_n5395_));
AND2X2 AND2X2_3317 ( .A(core__abc_22172_new_n5396_), .B(core__abc_22172_new_n1373_), .Y(core__abc_22172_new_n5397_));
AND2X2 AND2X2_3318 ( .A(core__abc_22172_new_n5398_), .B(core__abc_22172_new_n5399_), .Y(core__abc_22172_new_n5400_));
AND2X2 AND2X2_3319 ( .A(core__abc_22172_new_n5308_), .B(core__abc_22172_new_n3155_), .Y(core__abc_22172_new_n5402_));
AND2X2 AND2X2_332 ( .A(_abc_19873_new_n919_), .B(core_mi_57_), .Y(_abc_19873_new_n1473_));
AND2X2 AND2X2_3320 ( .A(core__abc_22172_new_n5404_), .B(core__abc_22172_new_n1928_), .Y(core__abc_22172_new_n5405_));
AND2X2 AND2X2_3321 ( .A(core__abc_22172_new_n5403_), .B(core__abc_22172_new_n1925_), .Y(core__abc_22172_new_n5406_));
AND2X2 AND2X2_3322 ( .A(core__abc_22172_new_n5409_), .B(core__abc_22172_new_n5411_), .Y(core__abc_22172_new_n5412_));
AND2X2 AND2X2_3323 ( .A(core__abc_22172_new_n5413_), .B(core__abc_22172_new_n5401_), .Y(core__abc_22172_new_n5414_));
AND2X2 AND2X2_3324 ( .A(core__abc_22172_new_n5412_), .B(core__abc_22172_new_n5400_), .Y(core__abc_22172_new_n5415_));
AND2X2 AND2X2_3325 ( .A(core__abc_22172_new_n5394_), .B(core__abc_22172_new_n5417_), .Y(core__abc_22172_new_n5418_));
AND2X2 AND2X2_3326 ( .A(core__abc_22172_new_n5393_), .B(core__abc_22172_new_n5416_), .Y(core__abc_22172_new_n5419_));
AND2X2 AND2X2_3327 ( .A(core__abc_22172_new_n5420_), .B(core__abc_22172_new_n4291_), .Y(core__abc_22172_new_n5421_));
AND2X2 AND2X2_3328 ( .A(core__abc_22172_new_n5423_), .B(core__abc_22172_new_n5422_), .Y(core__abc_22172_new_n5424_));
AND2X2 AND2X2_3329 ( .A(core__abc_22172_new_n5425_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n5426_));
AND2X2 AND2X2_333 ( .A(_abc_19873_new_n930_), .B(word0_reg_25_), .Y(_abc_19873_new_n1474_));
AND2X2 AND2X2_3330 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n5427_), .Y(core__abc_22172_new_n5428_));
AND2X2 AND2X2_3331 ( .A(core_v3_reg_38_), .B(core_mi_38_), .Y(core__abc_22172_new_n5430_));
AND2X2 AND2X2_3332 ( .A(core__abc_22172_new_n5431_), .B(core__abc_22172_new_n5429_), .Y(core__abc_22172_new_n5432_));
AND2X2 AND2X2_3333 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n5432_), .Y(core__abc_22172_new_n5433_));
AND2X2 AND2X2_3334 ( .A(core__abc_22172_new_n5435_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n5436_));
AND2X2 AND2X2_3335 ( .A(core__abc_22172_new_n5437_), .B(reset_n), .Y(core__0v3_reg_63_0__38_));
AND2X2 AND2X2_3336 ( .A(core__abc_22172_new_n5398_), .B(core__abc_22172_new_n1372_), .Y(core__abc_22172_new_n5440_));
AND2X2 AND2X2_3337 ( .A(core__abc_22172_new_n5440_), .B(core__abc_22172_new_n1400_), .Y(core__abc_22172_new_n5441_));
AND2X2 AND2X2_3338 ( .A(core__abc_22172_new_n5442_), .B(core__abc_22172_new_n5443_), .Y(core__abc_22172_new_n5444_));
AND2X2 AND2X2_3339 ( .A(core__abc_22172_new_n5446_), .B(core__abc_22172_new_n1945_), .Y(core__abc_22172_new_n5447_));
AND2X2 AND2X2_334 ( .A(_abc_19873_new_n928_), .B(core_key_57_), .Y(_abc_19873_new_n1476_));
AND2X2 AND2X2_3340 ( .A(core__abc_22172_new_n5445_), .B(core__abc_22172_new_n1942_), .Y(core__abc_22172_new_n5448_));
AND2X2 AND2X2_3341 ( .A(core__abc_22172_new_n5449_), .B(core_v3_reg_23_), .Y(core__abc_22172_new_n5450_));
AND2X2 AND2X2_3342 ( .A(core__abc_22172_new_n5451_), .B(core__abc_22172_new_n5452_), .Y(core__abc_22172_new_n5453_));
AND2X2 AND2X2_3343 ( .A(core__abc_22172_new_n5454_), .B(core__abc_22172_new_n5444_), .Y(core__abc_22172_new_n5455_));
AND2X2 AND2X2_3344 ( .A(core__abc_22172_new_n5456_), .B(core__abc_22172_new_n5457_), .Y(core__abc_22172_new_n5458_));
AND2X2 AND2X2_3345 ( .A(core__abc_22172_new_n5463_), .B(core__abc_22172_new_n5459_), .Y(core__abc_22172_new_n5464_));
AND2X2 AND2X2_3346 ( .A(core__abc_22172_new_n5467_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n5468_));
AND2X2 AND2X2_3347 ( .A(core__abc_22172_new_n5468_), .B(core__abc_22172_new_n5466_), .Y(core__abc_22172_new_n5469_));
AND2X2 AND2X2_3348 ( .A(core__abc_22172_new_n3214_), .B(core_key_103_), .Y(core__abc_22172_new_n5470_));
AND2X2 AND2X2_3349 ( .A(core_v3_reg_39_), .B(core_mi_39_), .Y(core__abc_22172_new_n5471_));
AND2X2 AND2X2_335 ( .A(_abc_19873_new_n901_), .B(core_key_25_), .Y(_abc_19873_new_n1477_));
AND2X2 AND2X2_3350 ( .A(core__abc_22172_new_n5472_), .B(core__abc_22172_new_n5473_), .Y(core__abc_22172_new_n5474_));
AND2X2 AND2X2_3351 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n5474_), .Y(core__abc_22172_new_n5475_));
AND2X2 AND2X2_3352 ( .A(core__abc_22172_new_n5479_), .B(reset_n), .Y(core__abc_22172_new_n5480_));
AND2X2 AND2X2_3353 ( .A(core__abc_22172_new_n5478_), .B(core__abc_22172_new_n5480_), .Y(core__0v3_reg_63_0__39_));
AND2X2 AND2X2_3354 ( .A(core__abc_22172_new_n3217_), .B(core_v3_reg_40_), .Y(core__abc_22172_new_n5482_));
AND2X2 AND2X2_3355 ( .A(core__abc_22172_new_n5458_), .B(core__abc_22172_new_n5417_), .Y(core__abc_22172_new_n5483_));
AND2X2 AND2X2_3356 ( .A(core__abc_22172_new_n5483_), .B(core__abc_22172_new_n5368_), .Y(core__abc_22172_new_n5484_));
AND2X2 AND2X2_3357 ( .A(core__abc_22172_new_n5298_), .B(core__abc_22172_new_n5484_), .Y(core__abc_22172_new_n5485_));
AND2X2 AND2X2_3358 ( .A(core__abc_22172_new_n5483_), .B(core__abc_22172_new_n5391_), .Y(core__abc_22172_new_n5486_));
AND2X2 AND2X2_3359 ( .A(core__abc_22172_new_n5487_), .B(core__abc_22172_new_n5457_), .Y(core__abc_22172_new_n5488_));
AND2X2 AND2X2_336 ( .A(_abc_19873_new_n1481_), .B(_abc_19873_new_n937_), .Y(\read_data[25] ));
AND2X2 AND2X2_3360 ( .A(core__abc_22172_new_n5484_), .B(core__abc_22172_new_n5299_), .Y(core__abc_22172_new_n5491_));
AND2X2 AND2X2_3361 ( .A(core__abc_22172_new_n5104_), .B(core__abc_22172_new_n5491_), .Y(core__abc_22172_new_n5492_));
AND2X2 AND2X2_3362 ( .A(core__abc_22172_new_n2935_), .B(core__abc_22172_new_n1411_), .Y(core__abc_22172_new_n5494_));
AND2X2 AND2X2_3363 ( .A(core__abc_22172_new_n3024_), .B(core__abc_22172_new_n1417_), .Y(core__abc_22172_new_n5495_));
AND2X2 AND2X2_3364 ( .A(core__abc_22172_new_n3180_), .B(core__abc_22172_new_n1959_), .Y(core__abc_22172_new_n5499_));
AND2X2 AND2X2_3365 ( .A(core__abc_22172_new_n5500_), .B(core__abc_22172_new_n1962_), .Y(core__abc_22172_new_n5501_));
AND2X2 AND2X2_3366 ( .A(core__abc_22172_new_n5504_), .B(core__abc_22172_new_n5505_), .Y(core__abc_22172_new_n5506_));
AND2X2 AND2X2_3367 ( .A(core__abc_22172_new_n5507_), .B(core__abc_22172_new_n5497_), .Y(core__abc_22172_new_n5508_));
AND2X2 AND2X2_3368 ( .A(core__abc_22172_new_n5506_), .B(core__abc_22172_new_n5496_), .Y(core__abc_22172_new_n5509_));
AND2X2 AND2X2_3369 ( .A(core__abc_22172_new_n5493_), .B(core__abc_22172_new_n5511_), .Y(core__abc_22172_new_n5512_));
AND2X2 AND2X2_337 ( .A(_abc_19873_new_n881_), .B(core_key_122_), .Y(_abc_19873_new_n1483_));
AND2X2 AND2X2_3370 ( .A(core__abc_22172_new_n5515_), .B(core__abc_22172_new_n5513_), .Y(core__abc_22172_new_n5516_));
AND2X2 AND2X2_3371 ( .A(core__abc_22172_new_n5516_), .B(core__abc_22172_new_n5510_), .Y(core__abc_22172_new_n5517_));
AND2X2 AND2X2_3372 ( .A(core__abc_22172_new_n5518_), .B(core__abc_22172_new_n4412_), .Y(core__abc_22172_new_n5519_));
AND2X2 AND2X2_3373 ( .A(core__abc_22172_new_n5521_), .B(core__abc_22172_new_n5520_), .Y(core__abc_22172_new_n5522_));
AND2X2 AND2X2_3374 ( .A(core__abc_22172_new_n5523_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n5524_));
AND2X2 AND2X2_3375 ( .A(core__abc_22172_new_n3214_), .B(core_key_104_), .Y(core__abc_22172_new_n5525_));
AND2X2 AND2X2_3376 ( .A(core_v3_reg_40_), .B(core_mi_40_), .Y(core__abc_22172_new_n5527_));
AND2X2 AND2X2_3377 ( .A(core__abc_22172_new_n5528_), .B(core__abc_22172_new_n5526_), .Y(core__abc_22172_new_n5529_));
AND2X2 AND2X2_3378 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n5529_), .Y(core__abc_22172_new_n5530_));
AND2X2 AND2X2_3379 ( .A(core__abc_22172_new_n5532_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n5533_));
AND2X2 AND2X2_338 ( .A(_abc_19873_new_n916_), .B(core_key_90_), .Y(_abc_19873_new_n1484_));
AND2X2 AND2X2_3380 ( .A(core__abc_22172_new_n5534_), .B(reset_n), .Y(core__0v3_reg_63_0__40_));
AND2X2 AND2X2_3381 ( .A(core__abc_22172_new_n3217_), .B(core_v3_reg_41_), .Y(core__abc_22172_new_n5536_));
AND2X2 AND2X2_3382 ( .A(core__abc_22172_new_n5538_), .B(core__abc_22172_new_n5537_), .Y(core__abc_22172_new_n5539_));
AND2X2 AND2X2_3383 ( .A(core__abc_22172_new_n5542_), .B(core__abc_22172_new_n1434_), .Y(core__abc_22172_new_n5543_));
AND2X2 AND2X2_3384 ( .A(core__abc_22172_new_n5541_), .B(core__abc_22172_new_n1428_), .Y(core__abc_22172_new_n5544_));
AND2X2 AND2X2_3385 ( .A(core__abc_22172_new_n5549_), .B(core__abc_22172_new_n1979_), .Y(core__abc_22172_new_n5550_));
AND2X2 AND2X2_3386 ( .A(core__abc_22172_new_n5548_), .B(core__abc_22172_new_n1976_), .Y(core__abc_22172_new_n5551_));
AND2X2 AND2X2_3387 ( .A(core__abc_22172_new_n5552_), .B(core__abc_22172_new_n5547_), .Y(core__abc_22172_new_n5553_));
AND2X2 AND2X2_3388 ( .A(core__abc_22172_new_n5554_), .B(core_v3_reg_25_), .Y(core__abc_22172_new_n5555_));
AND2X2 AND2X2_3389 ( .A(core__abc_22172_new_n5557_), .B(core__abc_22172_new_n5546_), .Y(core__abc_22172_new_n5558_));
AND2X2 AND2X2_339 ( .A(_abc_19873_new_n925_), .B(word2_reg_26_), .Y(_abc_19873_new_n1486_));
AND2X2 AND2X2_3390 ( .A(core__abc_22172_new_n5556_), .B(core__abc_22172_new_n5545_), .Y(core__abc_22172_new_n5560_));
AND2X2 AND2X2_3391 ( .A(core__abc_22172_new_n5559_), .B(core__abc_22172_new_n5561_), .Y(core__abc_22172_new_n5562_));
AND2X2 AND2X2_3392 ( .A(core__abc_22172_new_n5563_), .B(core__abc_22172_new_n5565_), .Y(core__abc_22172_new_n5566_));
AND2X2 AND2X2_3393 ( .A(core__abc_22172_new_n5568_), .B(core__abc_22172_new_n5569_), .Y(core__abc_22172_new_n5570_));
AND2X2 AND2X2_3394 ( .A(core__abc_22172_new_n5570_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n5571_));
AND2X2 AND2X2_3395 ( .A(core__abc_22172_new_n3214_), .B(core_key_105_), .Y(core__abc_22172_new_n5572_));
AND2X2 AND2X2_3396 ( .A(core_v3_reg_41_), .B(core_mi_41_), .Y(core__abc_22172_new_n5574_));
AND2X2 AND2X2_3397 ( .A(core__abc_22172_new_n5575_), .B(core__abc_22172_new_n5573_), .Y(core__abc_22172_new_n5576_));
AND2X2 AND2X2_3398 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n5576_), .Y(core__abc_22172_new_n5577_));
AND2X2 AND2X2_3399 ( .A(core__abc_22172_new_n5579_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n5580_));
AND2X2 AND2X2_34 ( .A(_abc_19873_new_n875_), .B(_abc_19873_new_n915_), .Y(_abc_19873_new_n916_));
AND2X2 AND2X2_340 ( .A(_abc_19873_new_n907_), .B(word1_reg_26_), .Y(_abc_19873_new_n1487_));
AND2X2 AND2X2_3400 ( .A(core__abc_22172_new_n5581_), .B(reset_n), .Y(core__0v3_reg_63_0__41_));
AND2X2 AND2X2_3401 ( .A(core__abc_22172_new_n3217_), .B(core_v3_reg_42_), .Y(core__abc_22172_new_n5583_));
AND2X2 AND2X2_3402 ( .A(core__abc_22172_new_n2935_), .B(core__abc_22172_new_n2939_), .Y(core__abc_22172_new_n5584_));
AND2X2 AND2X2_3403 ( .A(core__abc_22172_new_n5585_), .B(core__abc_22172_new_n1445_), .Y(core__abc_22172_new_n5586_));
AND2X2 AND2X2_3404 ( .A(core__abc_22172_new_n5587_), .B(core__abc_22172_new_n1451_), .Y(core__abc_22172_new_n5588_));
AND2X2 AND2X2_3405 ( .A(core__abc_22172_new_n5592_), .B(core__abc_22172_new_n1996_), .Y(core__abc_22172_new_n5593_));
AND2X2 AND2X2_3406 ( .A(core__abc_22172_new_n5596_), .B(core__abc_22172_new_n5597_), .Y(core__abc_22172_new_n5598_));
AND2X2 AND2X2_3407 ( .A(core__abc_22172_new_n5599_), .B(core__abc_22172_new_n5590_), .Y(core__abc_22172_new_n5600_));
AND2X2 AND2X2_3408 ( .A(core__abc_22172_new_n5598_), .B(core__abc_22172_new_n5589_), .Y(core__abc_22172_new_n5601_));
AND2X2 AND2X2_3409 ( .A(core__abc_22172_new_n5538_), .B(core__abc_22172_new_n5604_), .Y(core__abc_22172_new_n5605_));
AND2X2 AND2X2_341 ( .A(_abc_19873_new_n930_), .B(word0_reg_26_), .Y(_abc_19873_new_n1488_));
AND2X2 AND2X2_3410 ( .A(core__abc_22172_new_n5606_), .B(core__abc_22172_new_n5602_), .Y(core__abc_22172_new_n5608_));
AND2X2 AND2X2_3411 ( .A(core__abc_22172_new_n5609_), .B(core__abc_22172_new_n5607_), .Y(core__abc_22172_new_n5610_));
AND2X2 AND2X2_3412 ( .A(core__abc_22172_new_n5613_), .B(core__abc_22172_new_n5611_), .Y(core__abc_22172_new_n5614_));
AND2X2 AND2X2_3413 ( .A(core__abc_22172_new_n5614_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n5615_));
AND2X2 AND2X2_3414 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n5616_), .Y(core__abc_22172_new_n5617_));
AND2X2 AND2X2_3415 ( .A(core_v3_reg_42_), .B(core_mi_42_), .Y(core__abc_22172_new_n5619_));
AND2X2 AND2X2_3416 ( .A(core__abc_22172_new_n5620_), .B(core__abc_22172_new_n5618_), .Y(core__abc_22172_new_n5621_));
AND2X2 AND2X2_3417 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n5621_), .Y(core__abc_22172_new_n5622_));
AND2X2 AND2X2_3418 ( .A(core__abc_22172_new_n5624_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n5625_));
AND2X2 AND2X2_3419 ( .A(core__abc_22172_new_n5626_), .B(reset_n), .Y(core__0v3_reg_63_0__42_));
AND2X2 AND2X2_342 ( .A(_abc_19873_new_n912_), .B(word3_reg_26_), .Y(_abc_19873_new_n1492_));
AND2X2 AND2X2_3420 ( .A(core__abc_22172_new_n5607_), .B(core__abc_22172_new_n5628_), .Y(core__abc_22172_new_n5629_));
AND2X2 AND2X2_3421 ( .A(core__abc_22172_new_n5630_), .B(core__abc_22172_new_n1462_), .Y(core__abc_22172_new_n5632_));
AND2X2 AND2X2_3422 ( .A(core__abc_22172_new_n5633_), .B(core__abc_22172_new_n5631_), .Y(core__abc_22172_new_n5634_));
AND2X2 AND2X2_3423 ( .A(core__abc_22172_new_n3194_), .B(core__abc_22172_new_n5634_), .Y(core__abc_22172_new_n5635_));
AND2X2 AND2X2_3424 ( .A(core__abc_22172_new_n3193_), .B(core__abc_22172_new_n5636_), .Y(core__abc_22172_new_n5637_));
AND2X2 AND2X2_3425 ( .A(core__abc_22172_new_n5642_), .B(core__abc_22172_new_n5639_), .Y(core__abc_22172_new_n5643_));
AND2X2 AND2X2_3426 ( .A(core__abc_22172_new_n5646_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n5647_));
AND2X2 AND2X2_3427 ( .A(core__abc_22172_new_n5647_), .B(core__abc_22172_new_n5645_), .Y(core__abc_22172_new_n5648_));
AND2X2 AND2X2_3428 ( .A(core__abc_22172_new_n3214_), .B(core_key_107_), .Y(core__abc_22172_new_n5649_));
AND2X2 AND2X2_3429 ( .A(core_v3_reg_43_), .B(core_mi_43_), .Y(core__abc_22172_new_n5650_));
AND2X2 AND2X2_343 ( .A(_abc_19873_new_n928_), .B(core_key_58_), .Y(_abc_19873_new_n1493_));
AND2X2 AND2X2_3430 ( .A(core__abc_22172_new_n5651_), .B(core__abc_22172_new_n5652_), .Y(core__abc_22172_new_n5653_));
AND2X2 AND2X2_3431 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n5653_), .Y(core__abc_22172_new_n5654_));
AND2X2 AND2X2_3432 ( .A(core__abc_22172_new_n5658_), .B(reset_n), .Y(core__abc_22172_new_n5659_));
AND2X2 AND2X2_3433 ( .A(core__abc_22172_new_n5657_), .B(core__abc_22172_new_n5659_), .Y(core__0v3_reg_63_0__43_));
AND2X2 AND2X2_3434 ( .A(core__abc_22172_new_n3217_), .B(core_v3_reg_44_), .Y(core__abc_22172_new_n5661_));
AND2X2 AND2X2_3435 ( .A(core__abc_22172_new_n5603_), .B(core__abc_22172_new_n5561_), .Y(core__abc_22172_new_n5662_));
AND2X2 AND2X2_3436 ( .A(core__abc_22172_new_n5641_), .B(core__abc_22172_new_n5663_), .Y(core__abc_22172_new_n5664_));
AND2X2 AND2X2_3437 ( .A(core__abc_22172_new_n5664_), .B(core__abc_22172_new_n5662_), .Y(core__abc_22172_new_n5665_));
AND2X2 AND2X2_3438 ( .A(core__abc_22172_new_n5666_), .B(core__abc_22172_new_n5667_), .Y(core__abc_22172_new_n5668_));
AND2X2 AND2X2_3439 ( .A(core__abc_22172_new_n5562_), .B(core__abc_22172_new_n5511_), .Y(core__abc_22172_new_n5671_));
AND2X2 AND2X2_344 ( .A(_abc_19873_new_n901_), .B(core_key_26_), .Y(_abc_19873_new_n1494_));
AND2X2 AND2X2_3440 ( .A(core__abc_22172_new_n5664_), .B(core__abc_22172_new_n5671_), .Y(core__abc_22172_new_n5672_));
AND2X2 AND2X2_3441 ( .A(core__abc_22172_new_n5493_), .B(core__abc_22172_new_n5672_), .Y(core__abc_22172_new_n5673_));
AND2X2 AND2X2_3442 ( .A(core__abc_22172_new_n2935_), .B(core__abc_22172_new_n2941_), .Y(core__abc_22172_new_n5675_));
AND2X2 AND2X2_3443 ( .A(core__abc_22172_new_n5676_), .B(core__abc_22172_new_n1479_), .Y(core__abc_22172_new_n5677_));
AND2X2 AND2X2_3444 ( .A(core__abc_22172_new_n5678_), .B(core__abc_22172_new_n1485_), .Y(core__abc_22172_new_n5679_));
AND2X2 AND2X2_3445 ( .A(core__abc_22172_new_n3273_), .B(core__abc_22172_new_n5681_), .Y(core__abc_22172_new_n5682_));
AND2X2 AND2X2_3446 ( .A(core__abc_22172_new_n3272_), .B(core__abc_22172_new_n5680_), .Y(core__abc_22172_new_n5683_));
AND2X2 AND2X2_3447 ( .A(core__abc_22172_new_n5674_), .B(core__abc_22172_new_n5685_), .Y(core__abc_22172_new_n5686_));
AND2X2 AND2X2_3448 ( .A(core__abc_22172_new_n5687_), .B(core__abc_22172_new_n5668_), .Y(core__abc_22172_new_n5688_));
AND2X2 AND2X2_3449 ( .A(core__abc_22172_new_n5690_), .B(core__abc_22172_new_n5688_), .Y(core__abc_22172_new_n5691_));
AND2X2 AND2X2_345 ( .A(_abc_19873_new_n919_), .B(core_mi_58_), .Y(_abc_19873_new_n1496_));
AND2X2 AND2X2_3450 ( .A(core__abc_22172_new_n5691_), .B(core__abc_22172_new_n5684_), .Y(core__abc_22172_new_n5692_));
AND2X2 AND2X2_3451 ( .A(core__abc_22172_new_n5693_), .B(core__abc_22172_new_n4635_), .Y(core__abc_22172_new_n5694_));
AND2X2 AND2X2_3452 ( .A(core__abc_22172_new_n5695_), .B(core__abc_22172_new_n4639_), .Y(core__abc_22172_new_n5696_));
AND2X2 AND2X2_3453 ( .A(core__abc_22172_new_n5697_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n5698_));
AND2X2 AND2X2_3454 ( .A(core__abc_22172_new_n3214_), .B(core_key_108_), .Y(core__abc_22172_new_n5699_));
AND2X2 AND2X2_3455 ( .A(core_v3_reg_44_), .B(core_mi_44_), .Y(core__abc_22172_new_n5701_));
AND2X2 AND2X2_3456 ( .A(core__abc_22172_new_n5702_), .B(core__abc_22172_new_n5700_), .Y(core__abc_22172_new_n5703_));
AND2X2 AND2X2_3457 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n5703_), .Y(core__abc_22172_new_n5704_));
AND2X2 AND2X2_3458 ( .A(core__abc_22172_new_n5706_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n5707_));
AND2X2 AND2X2_3459 ( .A(core__abc_22172_new_n5708_), .B(reset_n), .Y(core__0v3_reg_63_0__44_));
AND2X2 AND2X2_346 ( .A(_abc_19873_new_n888_), .B(core_mi_26_), .Y(_abc_19873_new_n1497_));
AND2X2 AND2X2_3460 ( .A(core__abc_22172_new_n3217_), .B(core_v3_reg_45_), .Y(core__abc_22172_new_n5710_));
AND2X2 AND2X2_3461 ( .A(core__abc_22172_new_n5713_), .B(core__abc_22172_new_n1502_), .Y(core__abc_22172_new_n5714_));
AND2X2 AND2X2_3462 ( .A(core__abc_22172_new_n5712_), .B(core__abc_22172_new_n1496_), .Y(core__abc_22172_new_n5715_));
AND2X2 AND2X2_3463 ( .A(core__abc_22172_new_n3330_), .B(core__abc_22172_new_n5717_), .Y(core__abc_22172_new_n5718_));
AND2X2 AND2X2_3464 ( .A(core__abc_22172_new_n3329_), .B(core__abc_22172_new_n5716_), .Y(core__abc_22172_new_n5719_));
AND2X2 AND2X2_3465 ( .A(core__abc_22172_new_n5724_), .B(core__abc_22172_new_n5722_), .Y(core__abc_22172_new_n5725_));
AND2X2 AND2X2_3466 ( .A(core__abc_22172_new_n5725_), .B(core__abc_22172_new_n4706_), .Y(core__abc_22172_new_n5726_));
AND2X2 AND2X2_3467 ( .A(core__abc_22172_new_n5727_), .B(core__abc_22172_new_n4705_), .Y(core__abc_22172_new_n5728_));
AND2X2 AND2X2_3468 ( .A(core__abc_22172_new_n5729_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n5730_));
AND2X2 AND2X2_3469 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n5731_), .Y(core__abc_22172_new_n5732_));
AND2X2 AND2X2_347 ( .A(_abc_19873_new_n1501_), .B(_abc_19873_new_n937_), .Y(\read_data[26] ));
AND2X2 AND2X2_3470 ( .A(core_v3_reg_45_), .B(core_mi_45_), .Y(core__abc_22172_new_n5734_));
AND2X2 AND2X2_3471 ( .A(core__abc_22172_new_n5735_), .B(core__abc_22172_new_n5733_), .Y(core__abc_22172_new_n5736_));
AND2X2 AND2X2_3472 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n5736_), .Y(core__abc_22172_new_n5737_));
AND2X2 AND2X2_3473 ( .A(core__abc_22172_new_n5739_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n5740_));
AND2X2 AND2X2_3474 ( .A(core__abc_22172_new_n5741_), .B(reset_n), .Y(core__0v3_reg_63_0__45_));
AND2X2 AND2X2_3475 ( .A(core__abc_22172_new_n3217_), .B(core_v3_reg_46_), .Y(core__abc_22172_new_n5743_));
AND2X2 AND2X2_3476 ( .A(core__abc_22172_new_n5721_), .B(core__abc_22172_new_n5685_), .Y(core__abc_22172_new_n5744_));
AND2X2 AND2X2_3477 ( .A(core__abc_22172_new_n5674_), .B(core__abc_22172_new_n5744_), .Y(core__abc_22172_new_n5745_));
AND2X2 AND2X2_3478 ( .A(core__abc_22172_new_n5747_), .B(core__abc_22172_new_n5746_), .Y(core__abc_22172_new_n5748_));
AND2X2 AND2X2_3479 ( .A(core__abc_22172_new_n5676_), .B(core__abc_22172_new_n2937_), .Y(core__abc_22172_new_n5750_));
AND2X2 AND2X2_348 ( .A(_abc_19873_new_n881_), .B(core_key_123_), .Y(_abc_19873_new_n1503_));
AND2X2 AND2X2_3480 ( .A(core__abc_22172_new_n5751_), .B(core__abc_22172_new_n1513_), .Y(core__abc_22172_new_n5752_));
AND2X2 AND2X2_3481 ( .A(core__abc_22172_new_n5753_), .B(core__abc_22172_new_n5754_), .Y(core__abc_22172_new_n5755_));
AND2X2 AND2X2_3482 ( .A(core__abc_22172_new_n3395_), .B(core__abc_22172_new_n5756_), .Y(core__abc_22172_new_n5757_));
AND2X2 AND2X2_3483 ( .A(core__abc_22172_new_n3363_), .B(core__abc_22172_new_n5755_), .Y(core__abc_22172_new_n5758_));
AND2X2 AND2X2_3484 ( .A(core__abc_22172_new_n5749_), .B(core__abc_22172_new_n5760_), .Y(core__abc_22172_new_n5761_));
AND2X2 AND2X2_3485 ( .A(core__abc_22172_new_n5763_), .B(core__abc_22172_new_n5764_), .Y(core__abc_22172_new_n5765_));
AND2X2 AND2X2_3486 ( .A(core__abc_22172_new_n5765_), .B(core__abc_22172_new_n5759_), .Y(core__abc_22172_new_n5766_));
AND2X2 AND2X2_3487 ( .A(core__abc_22172_new_n5767_), .B(core__abc_22172_new_n4750_), .Y(core__abc_22172_new_n5768_));
AND2X2 AND2X2_3488 ( .A(core__abc_22172_new_n5769_), .B(core__abc_22172_new_n4747_), .Y(core__abc_22172_new_n5770_));
AND2X2 AND2X2_3489 ( .A(core__abc_22172_new_n5771_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n5772_));
AND2X2 AND2X2_349 ( .A(_abc_19873_new_n916_), .B(core_key_91_), .Y(_abc_19873_new_n1504_));
AND2X2 AND2X2_3490 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n5773_), .Y(core__abc_22172_new_n5774_));
AND2X2 AND2X2_3491 ( .A(core_v3_reg_46_), .B(core_mi_46_), .Y(core__abc_22172_new_n5776_));
AND2X2 AND2X2_3492 ( .A(core__abc_22172_new_n5777_), .B(core__abc_22172_new_n5775_), .Y(core__abc_22172_new_n5778_));
AND2X2 AND2X2_3493 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n5778_), .Y(core__abc_22172_new_n5779_));
AND2X2 AND2X2_3494 ( .A(core__abc_22172_new_n5781_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n5782_));
AND2X2 AND2X2_3495 ( .A(core__abc_22172_new_n5783_), .B(reset_n), .Y(core__0v3_reg_63_0__46_));
AND2X2 AND2X2_3496 ( .A(core__abc_22172_new_n3217_), .B(core_v3_reg_47_), .Y(core__abc_22172_new_n5785_));
AND2X2 AND2X2_3497 ( .A(core__abc_22172_new_n5787_), .B(core__abc_22172_new_n1530_), .Y(core__abc_22172_new_n5789_));
AND2X2 AND2X2_3498 ( .A(core__abc_22172_new_n5790_), .B(core__abc_22172_new_n5788_), .Y(core__abc_22172_new_n5791_));
AND2X2 AND2X2_3499 ( .A(core__abc_22172_new_n3452_), .B(core__abc_22172_new_n5791_), .Y(core__abc_22172_new_n5792_));
AND2X2 AND2X2_35 ( .A(_abc_19873_new_n916_), .B(core_key_64_), .Y(_abc_19873_new_n917_));
AND2X2 AND2X2_350 ( .A(_abc_19873_new_n912_), .B(word3_reg_27_), .Y(_abc_19873_new_n1506_));
AND2X2 AND2X2_3500 ( .A(core__abc_22172_new_n3457_), .B(core__abc_22172_new_n5793_), .Y(core__abc_22172_new_n5794_));
AND2X2 AND2X2_3501 ( .A(core__abc_22172_new_n5798_), .B(core__abc_22172_new_n5797_), .Y(core__abc_22172_new_n5799_));
AND2X2 AND2X2_3502 ( .A(core__abc_22172_new_n5801_), .B(core__abc_22172_new_n5800_), .Y(core__abc_22172_new_n5802_));
AND2X2 AND2X2_3503 ( .A(core__abc_22172_new_n5803_), .B(core__abc_22172_new_n5796_), .Y(core__abc_22172_new_n5804_));
AND2X2 AND2X2_3504 ( .A(core__abc_22172_new_n5807_), .B(core__abc_22172_new_n5806_), .Y(core__abc_22172_new_n5808_));
AND2X2 AND2X2_3505 ( .A(core__abc_22172_new_n5805_), .B(core__abc_22172_new_n5809_), .Y(core__abc_22172_new_n5810_));
AND2X2 AND2X2_3506 ( .A(core__abc_22172_new_n5810_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n5811_));
AND2X2 AND2X2_3507 ( .A(core__abc_22172_new_n3214_), .B(core_key_111_), .Y(core__abc_22172_new_n5812_));
AND2X2 AND2X2_3508 ( .A(core_v3_reg_47_), .B(core_mi_47_), .Y(core__abc_22172_new_n5814_));
AND2X2 AND2X2_3509 ( .A(core__abc_22172_new_n5815_), .B(core__abc_22172_new_n5813_), .Y(core__abc_22172_new_n5816_));
AND2X2 AND2X2_351 ( .A(_abc_19873_new_n907_), .B(word1_reg_27_), .Y(_abc_19873_new_n1507_));
AND2X2 AND2X2_3510 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n5816_), .Y(core__abc_22172_new_n5817_));
AND2X2 AND2X2_3511 ( .A(core__abc_22172_new_n5819_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n5820_));
AND2X2 AND2X2_3512 ( .A(core__abc_22172_new_n5821_), .B(reset_n), .Y(core__0v3_reg_63_0__47_));
AND2X2 AND2X2_3513 ( .A(core__abc_22172_new_n3217_), .B(core_v3_reg_48_), .Y(core__abc_22172_new_n5823_));
AND2X2 AND2X2_3514 ( .A(core__abc_22172_new_n5802_), .B(core__abc_22172_new_n5760_), .Y(core__abc_22172_new_n5824_));
AND2X2 AND2X2_3515 ( .A(core__abc_22172_new_n5824_), .B(core__abc_22172_new_n5744_), .Y(core__abc_22172_new_n5825_));
AND2X2 AND2X2_3516 ( .A(core__abc_22172_new_n5825_), .B(core__abc_22172_new_n5672_), .Y(core__abc_22172_new_n5826_));
AND2X2 AND2X2_3517 ( .A(core__abc_22172_new_n5826_), .B(core__abc_22172_new_n5491_), .Y(core__abc_22172_new_n5827_));
AND2X2 AND2X2_3518 ( .A(core__abc_22172_new_n5104_), .B(core__abc_22172_new_n5827_), .Y(core__abc_22172_new_n5828_));
AND2X2 AND2X2_3519 ( .A(core__abc_22172_new_n5490_), .B(core__abc_22172_new_n5826_), .Y(core__abc_22172_new_n5829_));
AND2X2 AND2X2_352 ( .A(_abc_19873_new_n930_), .B(word0_reg_27_), .Y(_abc_19873_new_n1508_));
AND2X2 AND2X2_3520 ( .A(core__abc_22172_new_n5670_), .B(core__abc_22172_new_n5825_), .Y(core__abc_22172_new_n5830_));
AND2X2 AND2X2_3521 ( .A(core__abc_22172_new_n5824_), .B(core__abc_22172_new_n5748_), .Y(core__abc_22172_new_n5831_));
AND2X2 AND2X2_3522 ( .A(core__abc_22172_new_n5832_), .B(core__abc_22172_new_n5801_), .Y(core__abc_22172_new_n5833_));
AND2X2 AND2X2_3523 ( .A(core__abc_22172_new_n2960_), .B(core__abc_22172_new_n1547_), .Y(core__abc_22172_new_n5838_));
AND2X2 AND2X2_3524 ( .A(core__abc_22172_new_n3028_), .B(core__abc_22172_new_n1553_), .Y(core__abc_22172_new_n5839_));
AND2X2 AND2X2_3525 ( .A(core__abc_22172_new_n3520_), .B(core__abc_22172_new_n5841_), .Y(core__abc_22172_new_n5842_));
AND2X2 AND2X2_3526 ( .A(core__abc_22172_new_n3519_), .B(core__abc_22172_new_n5840_), .Y(core__abc_22172_new_n5843_));
AND2X2 AND2X2_3527 ( .A(core__abc_22172_new_n5837_), .B(core__abc_22172_new_n5845_), .Y(core__abc_22172_new_n5846_));
AND2X2 AND2X2_3528 ( .A(core__abc_22172_new_n5851_), .B(core__abc_22172_new_n5850_), .Y(core__abc_22172_new_n5852_));
AND2X2 AND2X2_3529 ( .A(core__abc_22172_new_n5852_), .B(core__abc_22172_new_n5849_), .Y(core__abc_22172_new_n5853_));
AND2X2 AND2X2_353 ( .A(_abc_19873_new_n925_), .B(word2_reg_27_), .Y(_abc_19873_new_n1512_));
AND2X2 AND2X2_3530 ( .A(core__abc_22172_new_n5848_), .B(core__abc_22172_new_n5853_), .Y(core__abc_22172_new_n5854_));
AND2X2 AND2X2_3531 ( .A(core__abc_22172_new_n5854_), .B(core__abc_22172_new_n5844_), .Y(core__abc_22172_new_n5855_));
AND2X2 AND2X2_3532 ( .A(core__abc_22172_new_n5856_), .B(core__abc_22172_new_n4849_), .Y(core__abc_22172_new_n5857_));
AND2X2 AND2X2_3533 ( .A(core__abc_22172_new_n5858_), .B(core__abc_22172_new_n4846_), .Y(core__abc_22172_new_n5859_));
AND2X2 AND2X2_3534 ( .A(core__abc_22172_new_n5860_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n5861_));
AND2X2 AND2X2_3535 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n5862_), .Y(core__abc_22172_new_n5863_));
AND2X2 AND2X2_3536 ( .A(core_v3_reg_48_), .B(core_mi_48_), .Y(core__abc_22172_new_n5865_));
AND2X2 AND2X2_3537 ( .A(core__abc_22172_new_n5866_), .B(core__abc_22172_new_n5864_), .Y(core__abc_22172_new_n5867_));
AND2X2 AND2X2_3538 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n5867_), .Y(core__abc_22172_new_n5868_));
AND2X2 AND2X2_3539 ( .A(core__abc_22172_new_n5870_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n5871_));
AND2X2 AND2X2_354 ( .A(_abc_19873_new_n928_), .B(core_key_59_), .Y(_abc_19873_new_n1513_));
AND2X2 AND2X2_3540 ( .A(core__abc_22172_new_n5872_), .B(reset_n), .Y(core__0v3_reg_63_0__48_));
AND2X2 AND2X2_3541 ( .A(core__abc_22172_new_n3217_), .B(core_v3_reg_49_), .Y(core__abc_22172_new_n5874_));
AND2X2 AND2X2_3542 ( .A(core__abc_22172_new_n5878_), .B(core__abc_22172_new_n1570_), .Y(core__abc_22172_new_n5879_));
AND2X2 AND2X2_3543 ( .A(core__abc_22172_new_n5877_), .B(core__abc_22172_new_n1564_), .Y(core__abc_22172_new_n5880_));
AND2X2 AND2X2_3544 ( .A(core__abc_22172_new_n3586_), .B(core__abc_22172_new_n5881_), .Y(core__abc_22172_new_n5884_));
AND2X2 AND2X2_3545 ( .A(core__abc_22172_new_n5885_), .B(core__abc_22172_new_n5876_), .Y(core__abc_22172_new_n5886_));
AND2X2 AND2X2_3546 ( .A(core__abc_22172_new_n5875_), .B(core__abc_22172_new_n5886_), .Y(core__abc_22172_new_n5887_));
AND2X2 AND2X2_3547 ( .A(core__abc_22172_new_n5889_), .B(core__abc_22172_new_n5842_), .Y(core__abc_22172_new_n5890_));
AND2X2 AND2X2_3548 ( .A(core__abc_22172_new_n5889_), .B(core__abc_22172_new_n5845_), .Y(core__abc_22172_new_n5892_));
AND2X2 AND2X2_3549 ( .A(core__abc_22172_new_n5894_), .B(core__abc_22172_new_n5891_), .Y(core__abc_22172_new_n5895_));
AND2X2 AND2X2_355 ( .A(_abc_19873_new_n901_), .B(core_key_27_), .Y(_abc_19873_new_n1514_));
AND2X2 AND2X2_3550 ( .A(core__abc_22172_new_n5888_), .B(core__abc_22172_new_n5895_), .Y(core__abc_22172_new_n5896_));
AND2X2 AND2X2_3551 ( .A(core__abc_22172_new_n5897_), .B(core__abc_22172_new_n4913_), .Y(core__abc_22172_new_n5898_));
AND2X2 AND2X2_3552 ( .A(core__abc_22172_new_n5896_), .B(core__abc_22172_new_n4912_), .Y(core__abc_22172_new_n5899_));
AND2X2 AND2X2_3553 ( .A(core__abc_22172_new_n5900_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n5901_));
AND2X2 AND2X2_3554 ( .A(core__abc_22172_new_n3214_), .B(core_key_113_), .Y(core__abc_22172_new_n5902_));
AND2X2 AND2X2_3555 ( .A(core_v3_reg_49_), .B(core_mi_49_), .Y(core__abc_22172_new_n5904_));
AND2X2 AND2X2_3556 ( .A(core__abc_22172_new_n5905_), .B(core__abc_22172_new_n5903_), .Y(core__abc_22172_new_n5906_));
AND2X2 AND2X2_3557 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n5906_), .Y(core__abc_22172_new_n5907_));
AND2X2 AND2X2_3558 ( .A(core__abc_22172_new_n5909_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n5910_));
AND2X2 AND2X2_3559 ( .A(core__abc_22172_new_n5911_), .B(reset_n), .Y(core__0v3_reg_63_0__49_));
AND2X2 AND2X2_356 ( .A(_abc_19873_new_n919_), .B(core_mi_59_), .Y(_abc_19873_new_n1516_));
AND2X2 AND2X2_3560 ( .A(core__abc_22172_new_n3217_), .B(core_v3_reg_50_), .Y(core__abc_22172_new_n5913_));
AND2X2 AND2X2_3561 ( .A(core__abc_22172_new_n5891_), .B(core__abc_22172_new_n5882_), .Y(core__abc_22172_new_n5914_));
AND2X2 AND2X2_3562 ( .A(core__abc_22172_new_n5894_), .B(core__abc_22172_new_n5914_), .Y(core__abc_22172_new_n5915_));
AND2X2 AND2X2_3563 ( .A(core__abc_22172_new_n2960_), .B(core__abc_22172_new_n2971_), .Y(core__abc_22172_new_n5916_));
AND2X2 AND2X2_3564 ( .A(core__abc_22172_new_n5917_), .B(core__abc_22172_new_n1581_), .Y(core__abc_22172_new_n5918_));
AND2X2 AND2X2_3565 ( .A(core__abc_22172_new_n5919_), .B(core__abc_22172_new_n5920_), .Y(core__abc_22172_new_n5921_));
AND2X2 AND2X2_3566 ( .A(core__abc_22172_new_n3643_), .B(core__abc_22172_new_n5921_), .Y(core__abc_22172_new_n5922_));
AND2X2 AND2X2_3567 ( .A(core__abc_22172_new_n3642_), .B(core__abc_22172_new_n5923_), .Y(core__abc_22172_new_n5924_));
AND2X2 AND2X2_3568 ( .A(core__abc_22172_new_n5915_), .B(core__abc_22172_new_n5925_), .Y(core__abc_22172_new_n5928_));
AND2X2 AND2X2_3569 ( .A(core__abc_22172_new_n5929_), .B(core__abc_22172_new_n4959_), .Y(core__abc_22172_new_n5930_));
AND2X2 AND2X2_357 ( .A(_abc_19873_new_n888_), .B(core_mi_27_), .Y(_abc_19873_new_n1517_));
AND2X2 AND2X2_3570 ( .A(core__abc_22172_new_n5931_), .B(core__abc_22172_new_n4955_), .Y(core__abc_22172_new_n5932_));
AND2X2 AND2X2_3571 ( .A(core__abc_22172_new_n5933_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n5934_));
AND2X2 AND2X2_3572 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n5935_), .Y(core__abc_22172_new_n5936_));
AND2X2 AND2X2_3573 ( .A(core_v3_reg_50_), .B(core_mi_50_), .Y(core__abc_22172_new_n5938_));
AND2X2 AND2X2_3574 ( .A(core__abc_22172_new_n5939_), .B(core__abc_22172_new_n5937_), .Y(core__abc_22172_new_n5940_));
AND2X2 AND2X2_3575 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n5940_), .Y(core__abc_22172_new_n5941_));
AND2X2 AND2X2_3576 ( .A(core__abc_22172_new_n5943_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n5944_));
AND2X2 AND2X2_3577 ( .A(core__abc_22172_new_n5945_), .B(reset_n), .Y(core__0v3_reg_63_0__50_));
AND2X2 AND2X2_3578 ( .A(core__abc_22172_new_n3217_), .B(core_v3_reg_51_), .Y(core__abc_22172_new_n5947_));
AND2X2 AND2X2_3579 ( .A(core__abc_22172_new_n5926_), .B(core__abc_22172_new_n5948_), .Y(core__abc_22172_new_n5949_));
AND2X2 AND2X2_358 ( .A(_abc_19873_new_n1521_), .B(_abc_19873_new_n937_), .Y(\read_data[27] ));
AND2X2 AND2X2_3580 ( .A(core__abc_22172_new_n5950_), .B(core__abc_22172_new_n1598_), .Y(core__abc_22172_new_n5952_));
AND2X2 AND2X2_3581 ( .A(core__abc_22172_new_n5953_), .B(core__abc_22172_new_n5951_), .Y(core__abc_22172_new_n5954_));
AND2X2 AND2X2_3582 ( .A(core__abc_22172_new_n3716_), .B(core__abc_22172_new_n5955_), .Y(core__abc_22172_new_n5957_));
AND2X2 AND2X2_3583 ( .A(core__abc_22172_new_n5958_), .B(core__abc_22172_new_n5956_), .Y(core__abc_22172_new_n5959_));
AND2X2 AND2X2_3584 ( .A(core__abc_22172_new_n5949_), .B(core__abc_22172_new_n5960_), .Y(core__abc_22172_new_n5961_));
AND2X2 AND2X2_3585 ( .A(core__abc_22172_new_n5962_), .B(core__abc_22172_new_n5963_), .Y(core__abc_22172_new_n5964_));
AND2X2 AND2X2_3586 ( .A(core__abc_22172_new_n5964_), .B(core__abc_22172_new_n5007_), .Y(core__abc_22172_new_n5965_));
AND2X2 AND2X2_3587 ( .A(core__abc_22172_new_n5966_), .B(core__abc_22172_new_n5010_), .Y(core__abc_22172_new_n5967_));
AND2X2 AND2X2_3588 ( .A(core__abc_22172_new_n5968_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n5969_));
AND2X2 AND2X2_3589 ( .A(core__abc_22172_new_n3214_), .B(core_key_115_), .Y(core__abc_22172_new_n5970_));
AND2X2 AND2X2_359 ( .A(_abc_19873_new_n881_), .B(core_key_124_), .Y(_abc_19873_new_n1523_));
AND2X2 AND2X2_3590 ( .A(core_v3_reg_51_), .B(core_mi_51_), .Y(core__abc_22172_new_n5972_));
AND2X2 AND2X2_3591 ( .A(core__abc_22172_new_n5973_), .B(core__abc_22172_new_n5971_), .Y(core__abc_22172_new_n5974_));
AND2X2 AND2X2_3592 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n5974_), .Y(core__abc_22172_new_n5975_));
AND2X2 AND2X2_3593 ( .A(core__abc_22172_new_n5977_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n5978_));
AND2X2 AND2X2_3594 ( .A(core__abc_22172_new_n5979_), .B(reset_n), .Y(core__0v3_reg_63_0__51_));
AND2X2 AND2X2_3595 ( .A(core__abc_22172_new_n3217_), .B(core_v3_reg_52_), .Y(core__abc_22172_new_n5981_));
AND2X2 AND2X2_3596 ( .A(core__abc_22172_new_n5959_), .B(core__abc_22172_new_n5983_), .Y(core__abc_22172_new_n5984_));
AND2X2 AND2X2_3597 ( .A(core__abc_22172_new_n5984_), .B(core__abc_22172_new_n5982_), .Y(core__abc_22172_new_n5985_));
AND2X2 AND2X2_3598 ( .A(core__abc_22172_new_n5986_), .B(core__abc_22172_new_n5956_), .Y(core__abc_22172_new_n5987_));
AND2X2 AND2X2_3599 ( .A(core__abc_22172_new_n5984_), .B(core__abc_22172_new_n5892_), .Y(core__abc_22172_new_n5990_));
AND2X2 AND2X2_36 ( .A(_abc_19873_new_n886_), .B(_abc_19873_new_n903_), .Y(_abc_19873_new_n918_));
AND2X2 AND2X2_360 ( .A(_abc_19873_new_n888_), .B(core_mi_28_), .Y(_abc_19873_new_n1524_));
AND2X2 AND2X2_3600 ( .A(core__abc_22172_new_n5837_), .B(core__abc_22172_new_n5990_), .Y(core__abc_22172_new_n5991_));
AND2X2 AND2X2_3601 ( .A(core__abc_22172_new_n2960_), .B(core__abc_22172_new_n2973_), .Y(core__abc_22172_new_n5993_));
AND2X2 AND2X2_3602 ( .A(core__abc_22172_new_n5994_), .B(core__abc_22172_new_n1615_), .Y(core__abc_22172_new_n5995_));
AND2X2 AND2X2_3603 ( .A(core__abc_22172_new_n5996_), .B(core__abc_22172_new_n1621_), .Y(core__abc_22172_new_n5997_));
AND2X2 AND2X2_3604 ( .A(core__abc_22172_new_n3786_), .B(core__abc_22172_new_n5999_), .Y(core__abc_22172_new_n6000_));
AND2X2 AND2X2_3605 ( .A(core__abc_22172_new_n3785_), .B(core__abc_22172_new_n5998_), .Y(core__abc_22172_new_n6001_));
AND2X2 AND2X2_3606 ( .A(core__abc_22172_new_n5992_), .B(core__abc_22172_new_n6003_), .Y(core__abc_22172_new_n6004_));
AND2X2 AND2X2_3607 ( .A(core__abc_22172_new_n6007_), .B(core__abc_22172_new_n6005_), .Y(core__abc_22172_new_n6008_));
AND2X2 AND2X2_3608 ( .A(core__abc_22172_new_n6008_), .B(core__abc_22172_new_n6002_), .Y(core__abc_22172_new_n6009_));
AND2X2 AND2X2_3609 ( .A(core__abc_22172_new_n6010_), .B(core__abc_22172_new_n5055_), .Y(core__abc_22172_new_n6011_));
AND2X2 AND2X2_361 ( .A(_abc_19873_new_n916_), .B(core_key_92_), .Y(_abc_19873_new_n1526_));
AND2X2 AND2X2_3610 ( .A(core__abc_22172_new_n6012_), .B(core__abc_22172_new_n5062_), .Y(core__abc_22172_new_n6013_));
AND2X2 AND2X2_3611 ( .A(core__abc_22172_new_n6014_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n6015_));
AND2X2 AND2X2_3612 ( .A(core__abc_22172_new_n3214_), .B(core_key_116_), .Y(core__abc_22172_new_n6016_));
AND2X2 AND2X2_3613 ( .A(core_v3_reg_52_), .B(core_mi_52_), .Y(core__abc_22172_new_n6018_));
AND2X2 AND2X2_3614 ( .A(core__abc_22172_new_n6019_), .B(core__abc_22172_new_n6017_), .Y(core__abc_22172_new_n6020_));
AND2X2 AND2X2_3615 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n6020_), .Y(core__abc_22172_new_n6021_));
AND2X2 AND2X2_3616 ( .A(core__abc_22172_new_n6023_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n6024_));
AND2X2 AND2X2_3617 ( .A(core__abc_22172_new_n6025_), .B(reset_n), .Y(core__0v3_reg_63_0__52_));
AND2X2 AND2X2_3618 ( .A(core__abc_22172_new_n3217_), .B(core_v3_reg_53_), .Y(core__abc_22172_new_n6027_));
AND2X2 AND2X2_3619 ( .A(core__abc_22172_new_n6030_), .B(core__abc_22172_new_n1638_), .Y(core__abc_22172_new_n6031_));
AND2X2 AND2X2_362 ( .A(_abc_19873_new_n925_), .B(word2_reg_28_), .Y(_abc_19873_new_n1529_));
AND2X2 AND2X2_3620 ( .A(core__abc_22172_new_n6029_), .B(core__abc_22172_new_n1632_), .Y(core__abc_22172_new_n6032_));
AND2X2 AND2X2_3621 ( .A(core__abc_22172_new_n3850_), .B(core__abc_22172_new_n6034_), .Y(core__abc_22172_new_n6035_));
AND2X2 AND2X2_3622 ( .A(core__abc_22172_new_n3849_), .B(core__abc_22172_new_n6033_), .Y(core__abc_22172_new_n6036_));
AND2X2 AND2X2_3623 ( .A(core__abc_22172_new_n6041_), .B(core__abc_22172_new_n6039_), .Y(core__abc_22172_new_n6042_));
AND2X2 AND2X2_3624 ( .A(core__abc_22172_new_n6044_), .B(core__abc_22172_new_n6045_), .Y(core__abc_22172_new_n6046_));
AND2X2 AND2X2_3625 ( .A(core__abc_22172_new_n6046_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n6047_));
AND2X2 AND2X2_3626 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n6048_), .Y(core__abc_22172_new_n6049_));
AND2X2 AND2X2_3627 ( .A(core_v3_reg_53_), .B(core_mi_53_), .Y(core__abc_22172_new_n6051_));
AND2X2 AND2X2_3628 ( .A(core__abc_22172_new_n6052_), .B(core__abc_22172_new_n6050_), .Y(core__abc_22172_new_n6053_));
AND2X2 AND2X2_3629 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n6053_), .Y(core__abc_22172_new_n6054_));
AND2X2 AND2X2_363 ( .A(_abc_19873_new_n907_), .B(word1_reg_28_), .Y(_abc_19873_new_n1530_));
AND2X2 AND2X2_3630 ( .A(core__abc_22172_new_n6056_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n6057_));
AND2X2 AND2X2_3631 ( .A(core__abc_22172_new_n6058_), .B(reset_n), .Y(core__0v3_reg_63_0__53_));
AND2X2 AND2X2_3632 ( .A(core__abc_22172_new_n3217_), .B(core_v3_reg_54_), .Y(core__abc_22172_new_n6060_));
AND2X2 AND2X2_3633 ( .A(core__abc_22172_new_n6038_), .B(core__abc_22172_new_n6003_), .Y(core__abc_22172_new_n6061_));
AND2X2 AND2X2_3634 ( .A(core__abc_22172_new_n5992_), .B(core__abc_22172_new_n6061_), .Y(core__abc_22172_new_n6062_));
AND2X2 AND2X2_3635 ( .A(core__abc_22172_new_n6064_), .B(core__abc_22172_new_n6063_), .Y(core__abc_22172_new_n6065_));
AND2X2 AND2X2_3636 ( .A(core__abc_22172_new_n5994_), .B(core__abc_22172_new_n2969_), .Y(core__abc_22172_new_n6067_));
AND2X2 AND2X2_3637 ( .A(core__abc_22172_new_n6068_), .B(core__abc_22172_new_n1649_), .Y(core__abc_22172_new_n6069_));
AND2X2 AND2X2_3638 ( .A(core__abc_22172_new_n6070_), .B(core__abc_22172_new_n1655_), .Y(core__abc_22172_new_n6071_));
AND2X2 AND2X2_3639 ( .A(core__abc_22172_new_n3909_), .B(core__abc_22172_new_n6073_), .Y(core__abc_22172_new_n6074_));
AND2X2 AND2X2_364 ( .A(_abc_19873_new_n912_), .B(word3_reg_28_), .Y(_abc_19873_new_n1531_));
AND2X2 AND2X2_3640 ( .A(core__abc_22172_new_n3908_), .B(core__abc_22172_new_n6072_), .Y(core__abc_22172_new_n6075_));
AND2X2 AND2X2_3641 ( .A(core__abc_22172_new_n6066_), .B(core__abc_22172_new_n6077_), .Y(core__abc_22172_new_n6078_));
AND2X2 AND2X2_3642 ( .A(core__abc_22172_new_n6080_), .B(core__abc_22172_new_n6081_), .Y(core__abc_22172_new_n6082_));
AND2X2 AND2X2_3643 ( .A(core__abc_22172_new_n6082_), .B(core__abc_22172_new_n6076_), .Y(core__abc_22172_new_n6083_));
AND2X2 AND2X2_3644 ( .A(core__abc_22172_new_n6084_), .B(core__abc_22172_new_n5173_), .Y(core__abc_22172_new_n6085_));
AND2X2 AND2X2_3645 ( .A(core__abc_22172_new_n6086_), .B(core__abc_22172_new_n5172_), .Y(core__abc_22172_new_n6087_));
AND2X2 AND2X2_3646 ( .A(core__abc_22172_new_n6088_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n6089_));
AND2X2 AND2X2_3647 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n6090_), .Y(core__abc_22172_new_n6091_));
AND2X2 AND2X2_3648 ( .A(core_v3_reg_54_), .B(core_mi_54_), .Y(core__abc_22172_new_n6093_));
AND2X2 AND2X2_3649 ( .A(core__abc_22172_new_n6094_), .B(core__abc_22172_new_n6092_), .Y(core__abc_22172_new_n6095_));
AND2X2 AND2X2_365 ( .A(_abc_19873_new_n919_), .B(core_mi_60_), .Y(_abc_19873_new_n1534_));
AND2X2 AND2X2_3650 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n6095_), .Y(core__abc_22172_new_n6096_));
AND2X2 AND2X2_3651 ( .A(core__abc_22172_new_n6098_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n6099_));
AND2X2 AND2X2_3652 ( .A(core__abc_22172_new_n6100_), .B(reset_n), .Y(core__0v3_reg_63_0__54_));
AND2X2 AND2X2_3653 ( .A(core__abc_22172_new_n3217_), .B(core_v3_reg_55_), .Y(core__abc_22172_new_n6102_));
AND2X2 AND2X2_3654 ( .A(core__abc_22172_new_n6105_), .B(core__abc_22172_new_n1672_), .Y(core__abc_22172_new_n6106_));
AND2X2 AND2X2_3655 ( .A(core__abc_22172_new_n6104_), .B(core__abc_22172_new_n1666_), .Y(core__abc_22172_new_n6107_));
AND2X2 AND2X2_3656 ( .A(core__abc_22172_new_n3976_), .B(core__abc_22172_new_n6109_), .Y(core__abc_22172_new_n6110_));
AND2X2 AND2X2_3657 ( .A(core__abc_22172_new_n3980_), .B(core__abc_22172_new_n6108_), .Y(core__abc_22172_new_n6111_));
AND2X2 AND2X2_3658 ( .A(core__abc_22172_new_n6115_), .B(core__abc_22172_new_n6114_), .Y(core__abc_22172_new_n6116_));
AND2X2 AND2X2_3659 ( .A(core__abc_22172_new_n6118_), .B(core__abc_22172_new_n6117_), .Y(core__abc_22172_new_n6119_));
AND2X2 AND2X2_366 ( .A(_abc_19873_new_n930_), .B(word0_reg_28_), .Y(_abc_19873_new_n1535_));
AND2X2 AND2X2_3660 ( .A(core__abc_22172_new_n6120_), .B(core__abc_22172_new_n6113_), .Y(core__abc_22172_new_n6121_));
AND2X2 AND2X2_3661 ( .A(core__abc_22172_new_n6124_), .B(core__abc_22172_new_n6123_), .Y(core__abc_22172_new_n6125_));
AND2X2 AND2X2_3662 ( .A(core__abc_22172_new_n6122_), .B(core__abc_22172_new_n6126_), .Y(core__abc_22172_new_n6127_));
AND2X2 AND2X2_3663 ( .A(core__abc_22172_new_n6127_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n6128_));
AND2X2 AND2X2_3664 ( .A(core__abc_22172_new_n3214_), .B(core_key_119_), .Y(core__abc_22172_new_n6129_));
AND2X2 AND2X2_3665 ( .A(core_v3_reg_55_), .B(core_mi_55_), .Y(core__abc_22172_new_n6131_));
AND2X2 AND2X2_3666 ( .A(core__abc_22172_new_n6132_), .B(core__abc_22172_new_n6130_), .Y(core__abc_22172_new_n6133_));
AND2X2 AND2X2_3667 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n6133_), .Y(core__abc_22172_new_n6134_));
AND2X2 AND2X2_3668 ( .A(core__abc_22172_new_n6136_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n6137_));
AND2X2 AND2X2_3669 ( .A(core__abc_22172_new_n6138_), .B(reset_n), .Y(core__0v3_reg_63_0__55_));
AND2X2 AND2X2_367 ( .A(_abc_19873_new_n928_), .B(core_key_60_), .Y(_abc_19873_new_n1537_));
AND2X2 AND2X2_3670 ( .A(core__abc_22172_new_n3217_), .B(core_v3_reg_56_), .Y(core__abc_22172_new_n6140_));
AND2X2 AND2X2_3671 ( .A(core__abc_22172_new_n6119_), .B(core__abc_22172_new_n6077_), .Y(core__abc_22172_new_n6142_));
AND2X2 AND2X2_3672 ( .A(core__abc_22172_new_n6142_), .B(core__abc_22172_new_n6061_), .Y(core__abc_22172_new_n6143_));
AND2X2 AND2X2_3673 ( .A(core__abc_22172_new_n6143_), .B(core__abc_22172_new_n5990_), .Y(core__abc_22172_new_n6144_));
AND2X2 AND2X2_3674 ( .A(core__abc_22172_new_n5837_), .B(core__abc_22172_new_n6144_), .Y(core__abc_22172_new_n6145_));
AND2X2 AND2X2_3675 ( .A(core__abc_22172_new_n6143_), .B(core__abc_22172_new_n5989_), .Y(core__abc_22172_new_n6146_));
AND2X2 AND2X2_3676 ( .A(core__abc_22172_new_n6142_), .B(core__abc_22172_new_n6065_), .Y(core__abc_22172_new_n6147_));
AND2X2 AND2X2_3677 ( .A(core__abc_22172_new_n6148_), .B(core__abc_22172_new_n6117_), .Y(core__abc_22172_new_n6149_));
AND2X2 AND2X2_3678 ( .A(core__abc_22172_new_n2960_), .B(core__abc_22172_new_n2974_), .Y(core__abc_22172_new_n6154_));
AND2X2 AND2X2_3679 ( .A(core__abc_22172_new_n6155_), .B(core__abc_22172_new_n1683_), .Y(core__abc_22172_new_n6156_));
AND2X2 AND2X2_368 ( .A(_abc_19873_new_n901_), .B(core_key_28_), .Y(_abc_19873_new_n1538_));
AND2X2 AND2X2_3680 ( .A(core__abc_22172_new_n6157_), .B(core__abc_22172_new_n1689_), .Y(core__abc_22172_new_n6158_));
AND2X2 AND2X2_3681 ( .A(core__abc_22172_new_n4044_), .B(core__abc_22172_new_n6160_), .Y(core__abc_22172_new_n6161_));
AND2X2 AND2X2_3682 ( .A(core__abc_22172_new_n4045_), .B(core__abc_22172_new_n6159_), .Y(core__abc_22172_new_n6162_));
AND2X2 AND2X2_3683 ( .A(core__abc_22172_new_n6153_), .B(core__abc_22172_new_n6164_), .Y(core__abc_22172_new_n6165_));
AND2X2 AND2X2_3684 ( .A(core__abc_22172_new_n6171_), .B(core__abc_22172_new_n6149_), .Y(core__abc_22172_new_n6172_));
AND2X2 AND2X2_3685 ( .A(core__abc_22172_new_n6170_), .B(core__abc_22172_new_n6172_), .Y(core__abc_22172_new_n6173_));
AND2X2 AND2X2_3686 ( .A(core__abc_22172_new_n6169_), .B(core__abc_22172_new_n6173_), .Y(core__abc_22172_new_n6174_));
AND2X2 AND2X2_3687 ( .A(core__abc_22172_new_n6174_), .B(core__abc_22172_new_n6163_), .Y(core__abc_22172_new_n6175_));
AND2X2 AND2X2_3688 ( .A(core__abc_22172_new_n6176_), .B(core__abc_22172_new_n6141_), .Y(core__abc_22172_new_n6177_));
AND2X2 AND2X2_3689 ( .A(core__abc_22172_new_n6178_), .B(core__abc_22172_new_n5264_), .Y(core__abc_22172_new_n6179_));
AND2X2 AND2X2_369 ( .A(_abc_19873_new_n1542_), .B(_abc_19873_new_n937_), .Y(\read_data[28] ));
AND2X2 AND2X2_3690 ( .A(core__abc_22172_new_n6180_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n6181_));
AND2X2 AND2X2_3691 ( .A(core__abc_22172_new_n3214_), .B(core_key_120_), .Y(core__abc_22172_new_n6182_));
AND2X2 AND2X2_3692 ( .A(core_v3_reg_56_), .B(core_mi_56_), .Y(core__abc_22172_new_n6184_));
AND2X2 AND2X2_3693 ( .A(core__abc_22172_new_n6185_), .B(core__abc_22172_new_n6183_), .Y(core__abc_22172_new_n6186_));
AND2X2 AND2X2_3694 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n6186_), .Y(core__abc_22172_new_n6187_));
AND2X2 AND2X2_3695 ( .A(core__abc_22172_new_n6189_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n6190_));
AND2X2 AND2X2_3696 ( .A(core__abc_22172_new_n6191_), .B(reset_n), .Y(core__0v3_reg_63_0__56_));
AND2X2 AND2X2_3697 ( .A(core__abc_22172_new_n3217_), .B(core_v3_reg_57_), .Y(core__abc_22172_new_n6193_));
AND2X2 AND2X2_3698 ( .A(core__abc_22172_new_n6196_), .B(core__abc_22172_new_n1706_), .Y(core__abc_22172_new_n6197_));
AND2X2 AND2X2_3699 ( .A(core__abc_22172_new_n6195_), .B(core__abc_22172_new_n1700_), .Y(core__abc_22172_new_n6198_));
AND2X2 AND2X2_37 ( .A(_abc_19873_new_n875_), .B(_abc_19873_new_n918_), .Y(_abc_19873_new_n919_));
AND2X2 AND2X2_370 ( .A(_abc_19873_new_n928_), .B(core_key_61_), .Y(_abc_19873_new_n1544_));
AND2X2 AND2X2_3700 ( .A(core__abc_22172_new_n4109_), .B(core__abc_22172_new_n6200_), .Y(core__abc_22172_new_n6201_));
AND2X2 AND2X2_3701 ( .A(core__abc_22172_new_n4108_), .B(core__abc_22172_new_n6199_), .Y(core__abc_22172_new_n6202_));
AND2X2 AND2X2_3702 ( .A(core__abc_22172_new_n6207_), .B(core__abc_22172_new_n6205_), .Y(core__abc_22172_new_n6208_));
AND2X2 AND2X2_3703 ( .A(core__abc_22172_new_n6210_), .B(core__abc_22172_new_n6211_), .Y(core__abc_22172_new_n6212_));
AND2X2 AND2X2_3704 ( .A(core__abc_22172_new_n6212_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n6213_));
AND2X2 AND2X2_3705 ( .A(core__abc_22172_new_n3214_), .B(core_key_121_), .Y(core__abc_22172_new_n6214_));
AND2X2 AND2X2_3706 ( .A(core_v3_reg_57_), .B(core_mi_57_), .Y(core__abc_22172_new_n6216_));
AND2X2 AND2X2_3707 ( .A(core__abc_22172_new_n6217_), .B(core__abc_22172_new_n6215_), .Y(core__abc_22172_new_n6218_));
AND2X2 AND2X2_3708 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n6218_), .Y(core__abc_22172_new_n6219_));
AND2X2 AND2X2_3709 ( .A(core__abc_22172_new_n6221_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n6222_));
AND2X2 AND2X2_371 ( .A(_abc_19873_new_n901_), .B(core_key_29_), .Y(_abc_19873_new_n1545_));
AND2X2 AND2X2_3710 ( .A(core__abc_22172_new_n6223_), .B(reset_n), .Y(core__0v3_reg_63_0__57_));
AND2X2 AND2X2_3711 ( .A(core__abc_22172_new_n3217_), .B(core_v3_reg_58_), .Y(core__abc_22172_new_n6225_));
AND2X2 AND2X2_3712 ( .A(core__abc_22172_new_n6227_), .B(core__abc_22172_new_n6229_), .Y(core__abc_22172_new_n6230_));
AND2X2 AND2X2_3713 ( .A(core__abc_22172_new_n6204_), .B(core__abc_22172_new_n6164_), .Y(core__abc_22172_new_n6232_));
AND2X2 AND2X2_3714 ( .A(core__abc_22172_new_n6153_), .B(core__abc_22172_new_n6232_), .Y(core__abc_22172_new_n6233_));
AND2X2 AND2X2_3715 ( .A(core__abc_22172_new_n6236_), .B(core__abc_22172_new_n2996_), .Y(core__abc_22172_new_n6237_));
AND2X2 AND2X2_3716 ( .A(core__abc_22172_new_n6237_), .B(core__abc_22172_new_n1723_), .Y(core__abc_22172_new_n6240_));
AND2X2 AND2X2_3717 ( .A(core__abc_22172_new_n4169_), .B(core__abc_22172_new_n6242_), .Y(core__abc_22172_new_n6243_));
AND2X2 AND2X2_3718 ( .A(core__abc_22172_new_n4168_), .B(core__abc_22172_new_n6241_), .Y(core__abc_22172_new_n6244_));
AND2X2 AND2X2_3719 ( .A(core__abc_22172_new_n6234_), .B(core__abc_22172_new_n6246_), .Y(core__abc_22172_new_n6247_));
AND2X2 AND2X2_372 ( .A(_abc_19873_new_n916_), .B(core_key_93_), .Y(_abc_19873_new_n1547_));
AND2X2 AND2X2_3720 ( .A(core__abc_22172_new_n6248_), .B(core__abc_22172_new_n6249_), .Y(core__abc_22172_new_n6250_));
AND2X2 AND2X2_3721 ( .A(core__abc_22172_new_n6251_), .B(core__abc_22172_new_n6226_), .Y(core__abc_22172_new_n6252_));
AND2X2 AND2X2_3722 ( .A(core__abc_22172_new_n6250_), .B(core__abc_22172_new_n5357_), .Y(core__abc_22172_new_n6253_));
AND2X2 AND2X2_3723 ( .A(core__abc_22172_new_n6254_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n6255_));
AND2X2 AND2X2_3724 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n6256_), .Y(core__abc_22172_new_n6257_));
AND2X2 AND2X2_3725 ( .A(core_v3_reg_58_), .B(core_mi_58_), .Y(core__abc_22172_new_n6259_));
AND2X2 AND2X2_3726 ( .A(core__abc_22172_new_n6260_), .B(core__abc_22172_new_n6258_), .Y(core__abc_22172_new_n6261_));
AND2X2 AND2X2_3727 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n6261_), .Y(core__abc_22172_new_n6262_));
AND2X2 AND2X2_3728 ( .A(core__abc_22172_new_n6264_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n6265_));
AND2X2 AND2X2_3729 ( .A(core__abc_22172_new_n6266_), .B(reset_n), .Y(core__0v3_reg_63_0__58_));
AND2X2 AND2X2_373 ( .A(_abc_19873_new_n881_), .B(core_key_125_), .Y(_abc_19873_new_n1548_));
AND2X2 AND2X2_3730 ( .A(core__abc_22172_new_n6248_), .B(core__abc_22172_new_n6268_), .Y(core__abc_22172_new_n6269_));
AND2X2 AND2X2_3731 ( .A(core__abc_22172_new_n6238_), .B(core__abc_22172_new_n1716_), .Y(core__abc_22172_new_n6271_));
AND2X2 AND2X2_3732 ( .A(core__abc_22172_new_n6271_), .B(core__abc_22172_new_n1740_), .Y(core__abc_22172_new_n6272_));
AND2X2 AND2X2_3733 ( .A(core__abc_22172_new_n6273_), .B(core__abc_22172_new_n6274_), .Y(core__abc_22172_new_n6275_));
AND2X2 AND2X2_3734 ( .A(core__abc_22172_new_n6277_), .B(core__abc_22172_new_n6278_), .Y(core__abc_22172_new_n6279_));
AND2X2 AND2X2_3735 ( .A(core__abc_22172_new_n4251_), .B(core__abc_22172_new_n6275_), .Y(core__abc_22172_new_n6281_));
AND2X2 AND2X2_3736 ( .A(core__abc_22172_new_n4255_), .B(core__abc_22172_new_n6276_), .Y(core__abc_22172_new_n6282_));
AND2X2 AND2X2_3737 ( .A(core__abc_22172_new_n6280_), .B(core__abc_22172_new_n6284_), .Y(core__abc_22172_new_n6285_));
AND2X2 AND2X2_3738 ( .A(core__abc_22172_new_n6288_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n6289_));
AND2X2 AND2X2_3739 ( .A(core__abc_22172_new_n6289_), .B(core__abc_22172_new_n6287_), .Y(core__abc_22172_new_n6290_));
AND2X2 AND2X2_374 ( .A(_abc_19873_new_n930_), .B(word0_reg_29_), .Y(_abc_19873_new_n1551_));
AND2X2 AND2X2_3740 ( .A(core__abc_22172_new_n3214_), .B(core_key_123_), .Y(core__abc_22172_new_n6291_));
AND2X2 AND2X2_3741 ( .A(core_v3_reg_59_), .B(core_mi_59_), .Y(core__abc_22172_new_n6292_));
AND2X2 AND2X2_3742 ( .A(core__abc_22172_new_n6293_), .B(core__abc_22172_new_n6294_), .Y(core__abc_22172_new_n6295_));
AND2X2 AND2X2_3743 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n6295_), .Y(core__abc_22172_new_n6296_));
AND2X2 AND2X2_3744 ( .A(core__abc_22172_new_n6300_), .B(reset_n), .Y(core__abc_22172_new_n6301_));
AND2X2 AND2X2_3745 ( .A(core__abc_22172_new_n6299_), .B(core__abc_22172_new_n6301_), .Y(core__0v3_reg_63_0__59_));
AND2X2 AND2X2_3746 ( .A(core__abc_22172_new_n3217_), .B(core_v3_reg_60_), .Y(core__abc_22172_new_n6303_));
AND2X2 AND2X2_3747 ( .A(core__abc_22172_new_n6279_), .B(core__abc_22172_new_n6246_), .Y(core__abc_22172_new_n6304_));
AND2X2 AND2X2_3748 ( .A(core__abc_22172_new_n6304_), .B(core__abc_22172_new_n6232_), .Y(core__abc_22172_new_n6305_));
AND2X2 AND2X2_3749 ( .A(core__abc_22172_new_n6153_), .B(core__abc_22172_new_n6305_), .Y(core__abc_22172_new_n6306_));
AND2X2 AND2X2_375 ( .A(_abc_19873_new_n907_), .B(word1_reg_29_), .Y(_abc_19873_new_n1552_));
AND2X2 AND2X2_3750 ( .A(core__abc_22172_new_n6304_), .B(core__abc_22172_new_n6231_), .Y(core__abc_22172_new_n6307_));
AND2X2 AND2X2_3751 ( .A(core__abc_22172_new_n6308_), .B(core__abc_22172_new_n6277_), .Y(core__abc_22172_new_n6309_));
AND2X2 AND2X2_3752 ( .A(core__abc_22172_new_n6155_), .B(core__abc_22172_new_n2966_), .Y(core__abc_22172_new_n6313_));
AND2X2 AND2X2_3753 ( .A(core__abc_22172_new_n6314_), .B(core__abc_22172_new_n1751_), .Y(core__abc_22172_new_n6315_));
AND2X2 AND2X2_3754 ( .A(core__abc_22172_new_n6316_), .B(core__abc_22172_new_n1757_), .Y(core__abc_22172_new_n6317_));
AND2X2 AND2X2_3755 ( .A(core__abc_22172_new_n4320_), .B(core__abc_22172_new_n6319_), .Y(core__abc_22172_new_n6320_));
AND2X2 AND2X2_3756 ( .A(core__abc_22172_new_n4321_), .B(core__abc_22172_new_n6318_), .Y(core__abc_22172_new_n6321_));
AND2X2 AND2X2_3757 ( .A(core__abc_22172_new_n6312_), .B(core__abc_22172_new_n6323_), .Y(core__abc_22172_new_n6324_));
AND2X2 AND2X2_3758 ( .A(core__abc_22172_new_n6329_), .B(core__abc_22172_new_n6309_), .Y(core__abc_22172_new_n6330_));
AND2X2 AND2X2_3759 ( .A(core__abc_22172_new_n6328_), .B(core__abc_22172_new_n6330_), .Y(core__abc_22172_new_n6331_));
AND2X2 AND2X2_376 ( .A(_abc_19873_new_n925_), .B(word2_reg_29_), .Y(_abc_19873_new_n1554_));
AND2X2 AND2X2_3760 ( .A(core__abc_22172_new_n6331_), .B(core__abc_22172_new_n6322_), .Y(core__abc_22172_new_n6332_));
AND2X2 AND2X2_3761 ( .A(core__abc_22172_new_n6333_), .B(core__abc_22172_new_n5454_), .Y(core__abc_22172_new_n6334_));
AND2X2 AND2X2_3762 ( .A(core__abc_22172_new_n6335_), .B(core__abc_22172_new_n5453_), .Y(core__abc_22172_new_n6336_));
AND2X2 AND2X2_3763 ( .A(core__abc_22172_new_n6337_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n6338_));
AND2X2 AND2X2_3764 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n6339_), .Y(core__abc_22172_new_n6340_));
AND2X2 AND2X2_3765 ( .A(core_v3_reg_60_), .B(core_mi_60_), .Y(core__abc_22172_new_n6342_));
AND2X2 AND2X2_3766 ( .A(core__abc_22172_new_n6343_), .B(core__abc_22172_new_n6341_), .Y(core__abc_22172_new_n6344_));
AND2X2 AND2X2_3767 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n6344_), .Y(core__abc_22172_new_n6345_));
AND2X2 AND2X2_3768 ( .A(core__abc_22172_new_n6347_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n6348_));
AND2X2 AND2X2_3769 ( .A(core__abc_22172_new_n6349_), .B(reset_n), .Y(core__0v3_reg_63_0__60_));
AND2X2 AND2X2_377 ( .A(_abc_19873_new_n912_), .B(word3_reg_29_), .Y(_abc_19873_new_n1555_));
AND2X2 AND2X2_3770 ( .A(core__abc_22172_new_n3217_), .B(core_v3_reg_61_), .Y(core__abc_22172_new_n6351_));
AND2X2 AND2X2_3771 ( .A(core__abc_22172_new_n6354_), .B(core__abc_22172_new_n1774_), .Y(core__abc_22172_new_n6355_));
AND2X2 AND2X2_3772 ( .A(core__abc_22172_new_n6353_), .B(core__abc_22172_new_n1768_), .Y(core__abc_22172_new_n6356_));
AND2X2 AND2X2_3773 ( .A(core__abc_22172_new_n4381_), .B(core__abc_22172_new_n6358_), .Y(core__abc_22172_new_n6359_));
AND2X2 AND2X2_3774 ( .A(core__abc_22172_new_n4376_), .B(core__abc_22172_new_n6357_), .Y(core__abc_22172_new_n6360_));
AND2X2 AND2X2_3775 ( .A(core__abc_22172_new_n6364_), .B(core__abc_22172_new_n6363_), .Y(core__abc_22172_new_n6365_));
AND2X2 AND2X2_3776 ( .A(core__abc_22172_new_n6367_), .B(core__abc_22172_new_n6366_), .Y(core__abc_22172_new_n6368_));
AND2X2 AND2X2_3777 ( .A(core__abc_22172_new_n6369_), .B(core__abc_22172_new_n6362_), .Y(core__abc_22172_new_n6370_));
AND2X2 AND2X2_3778 ( .A(core__abc_22172_new_n6373_), .B(core__abc_22172_new_n6372_), .Y(core__abc_22172_new_n6374_));
AND2X2 AND2X2_3779 ( .A(core__abc_22172_new_n6371_), .B(core__abc_22172_new_n6375_), .Y(core__abc_22172_new_n6376_));
AND2X2 AND2X2_378 ( .A(_abc_19873_new_n888_), .B(core_mi_29_), .Y(_abc_19873_new_n1558_));
AND2X2 AND2X2_3780 ( .A(core__abc_22172_new_n6376_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n6377_));
AND2X2 AND2X2_3781 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n6378_), .Y(core__abc_22172_new_n6379_));
AND2X2 AND2X2_3782 ( .A(core_v3_reg_61_), .B(core_mi_61_), .Y(core__abc_22172_new_n6381_));
AND2X2 AND2X2_3783 ( .A(core__abc_22172_new_n6382_), .B(core__abc_22172_new_n6380_), .Y(core__abc_22172_new_n6383_));
AND2X2 AND2X2_3784 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n6383_), .Y(core__abc_22172_new_n6384_));
AND2X2 AND2X2_3785 ( .A(core__abc_22172_new_n6386_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n6387_));
AND2X2 AND2X2_3786 ( .A(core__abc_22172_new_n6388_), .B(reset_n), .Y(core__0v3_reg_63_0__61_));
AND2X2 AND2X2_3787 ( .A(core__abc_22172_new_n3217_), .B(core_v3_reg_62_), .Y(core__abc_22172_new_n6390_));
AND2X2 AND2X2_3788 ( .A(core__abc_22172_new_n6367_), .B(core__abc_22172_new_n6320_), .Y(core__abc_22172_new_n6393_));
AND2X2 AND2X2_3789 ( .A(core__abc_22172_new_n6392_), .B(core__abc_22172_new_n6395_), .Y(core__abc_22172_new_n6396_));
AND2X2 AND2X2_379 ( .A(_abc_19873_new_n919_), .B(core_mi_61_), .Y(_abc_19873_new_n1559_));
AND2X2 AND2X2_3790 ( .A(core__abc_22172_new_n6314_), .B(core__abc_22172_new_n2962_), .Y(core__abc_22172_new_n6397_));
AND2X2 AND2X2_3791 ( .A(core__abc_22172_new_n6398_), .B(core__abc_22172_new_n1785_), .Y(core__abc_22172_new_n6399_));
AND2X2 AND2X2_3792 ( .A(core__abc_22172_new_n6400_), .B(core__abc_22172_new_n1791_), .Y(core__abc_22172_new_n6401_));
AND2X2 AND2X2_3793 ( .A(core__abc_22172_new_n4434_), .B(core__abc_22172_new_n6403_), .Y(core__abc_22172_new_n6404_));
AND2X2 AND2X2_3794 ( .A(core__abc_22172_new_n4432_), .B(core__abc_22172_new_n6402_), .Y(core__abc_22172_new_n6405_));
AND2X2 AND2X2_3795 ( .A(core__abc_22172_new_n6396_), .B(core__abc_22172_new_n6406_), .Y(core__abc_22172_new_n6407_));
AND2X2 AND2X2_3796 ( .A(core__abc_22172_new_n6368_), .B(core__abc_22172_new_n6323_), .Y(core__abc_22172_new_n6408_));
AND2X2 AND2X2_3797 ( .A(core__abc_22172_new_n6312_), .B(core__abc_22172_new_n6408_), .Y(core__abc_22172_new_n6409_));
AND2X2 AND2X2_3798 ( .A(core__abc_22172_new_n6410_), .B(core__abc_22172_new_n6411_), .Y(core__abc_22172_new_n6412_));
AND2X2 AND2X2_3799 ( .A(core__abc_22172_new_n6416_), .B(core__abc_22172_new_n6415_), .Y(core__abc_22172_new_n6417_));
AND2X2 AND2X2_38 ( .A(_abc_19873_new_n919_), .B(core_mi_32_), .Y(_abc_19873_new_n920_));
AND2X2 AND2X2_380 ( .A(_abc_19873_new_n1563_), .B(_abc_19873_new_n937_), .Y(\read_data[29] ));
AND2X2 AND2X2_3800 ( .A(core__abc_22172_new_n6414_), .B(core__abc_22172_new_n6418_), .Y(core__abc_22172_new_n6419_));
AND2X2 AND2X2_3801 ( .A(core__abc_22172_new_n6419_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n6420_));
AND2X2 AND2X2_3802 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n6421_), .Y(core__abc_22172_new_n6422_));
AND2X2 AND2X2_3803 ( .A(core_v3_reg_62_), .B(core_mi_62_), .Y(core__abc_22172_new_n6424_));
AND2X2 AND2X2_3804 ( .A(core__abc_22172_new_n6425_), .B(core__abc_22172_new_n6423_), .Y(core__abc_22172_new_n6426_));
AND2X2 AND2X2_3805 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n6426_), .Y(core__abc_22172_new_n6427_));
AND2X2 AND2X2_3806 ( .A(core__abc_22172_new_n6429_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n6430_));
AND2X2 AND2X2_3807 ( .A(core__abc_22172_new_n6431_), .B(reset_n), .Y(core__0v3_reg_63_0__62_));
AND2X2 AND2X2_3808 ( .A(core__abc_22172_new_n6435_), .B(core__abc_22172_new_n1808_), .Y(core__abc_22172_new_n6436_));
AND2X2 AND2X2_3809 ( .A(core__abc_22172_new_n6434_), .B(core__abc_22172_new_n1802_), .Y(core__abc_22172_new_n6437_));
AND2X2 AND2X2_381 ( .A(_abc_19873_new_n881_), .B(core_key_126_), .Y(_abc_19873_new_n1565_));
AND2X2 AND2X2_3810 ( .A(core__abc_22172_new_n4504_), .B(core__abc_22172_new_n6439_), .Y(core__abc_22172_new_n6440_));
AND2X2 AND2X2_3811 ( .A(core__abc_22172_new_n4503_), .B(core__abc_22172_new_n6438_), .Y(core__abc_22172_new_n6441_));
AND2X2 AND2X2_3812 ( .A(core__abc_22172_new_n6416_), .B(core__abc_22172_new_n6444_), .Y(core__abc_22172_new_n6445_));
AND2X2 AND2X2_3813 ( .A(core__abc_22172_new_n6447_), .B(core__abc_22172_new_n6443_), .Y(core__abc_22172_new_n6448_));
AND2X2 AND2X2_3814 ( .A(core__abc_22172_new_n6451_), .B(core__abc_22172_new_n6450_), .Y(core__abc_22172_new_n6452_));
AND2X2 AND2X2_3815 ( .A(core__abc_22172_new_n6453_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n6454_));
AND2X2 AND2X2_3816 ( .A(core__abc_22172_new_n6454_), .B(core__abc_22172_new_n6449_), .Y(core__abc_22172_new_n6455_));
AND2X2 AND2X2_3817 ( .A(core__abc_22172_new_n3214_), .B(core_key_127_), .Y(core__abc_22172_new_n6456_));
AND2X2 AND2X2_3818 ( .A(core_v3_reg_63_), .B(core_mi_63_), .Y(core__abc_22172_new_n6457_));
AND2X2 AND2X2_3819 ( .A(core__abc_22172_new_n6458_), .B(core__abc_22172_new_n6459_), .Y(core__abc_22172_new_n6460_));
AND2X2 AND2X2_382 ( .A(_abc_19873_new_n888_), .B(core_mi_30_), .Y(_abc_19873_new_n1566_));
AND2X2 AND2X2_3820 ( .A(core__abc_22172_new_n2660_), .B(core__abc_22172_new_n6460_), .Y(core__abc_22172_new_n6461_));
AND2X2 AND2X2_3821 ( .A(core__abc_22172_new_n6465_), .B(reset_n), .Y(core__abc_22172_new_n6466_));
AND2X2 AND2X2_3822 ( .A(core__abc_22172_new_n6464_), .B(core__abc_22172_new_n6466_), .Y(core__0v3_reg_63_0__63_));
AND2X2 AND2X2_3823 ( .A(core__abc_22172_new_n6438_), .B(core__abc_22172_new_n6468_), .Y(core__abc_22172_new_n6469_));
AND2X2 AND2X2_3824 ( .A(core__abc_22172_new_n6439_), .B(core_v1_reg_18_), .Y(core__abc_22172_new_n6470_));
AND2X2 AND2X2_3825 ( .A(core__abc_22172_new_n6471_), .B(core__abc_22172_new_n5050_), .Y(core__abc_22172_new_n6473_));
AND2X2 AND2X2_3826 ( .A(core__abc_22172_new_n6474_), .B(core__abc_22172_new_n6472_), .Y(core__abc_22172_new_n6475_));
AND2X2 AND2X2_3827 ( .A(core__abc_22172_new_n6477_), .B(core__abc_22172_new_n6478_), .Y(core__abc_22172_new_n6479_));
AND2X2 AND2X2_3828 ( .A(core__abc_22172_new_n6482_), .B(core__abc_22172_new_n6480_), .Y(core__abc_22172_new_n6483_));
AND2X2 AND2X2_3829 ( .A(core__abc_22172_new_n6475_), .B(core__abc_22172_new_n6483_), .Y(core__abc_22172_new_n6484_));
AND2X2 AND2X2_383 ( .A(_abc_19873_new_n916_), .B(core_key_94_), .Y(_abc_19873_new_n1568_));
AND2X2 AND2X2_3830 ( .A(core__abc_22172_new_n6357_), .B(core__abc_22172_new_n6486_), .Y(core__abc_22172_new_n6487_));
AND2X2 AND2X2_3831 ( .A(core__abc_22172_new_n6358_), .B(core_v1_reg_16_), .Y(core__abc_22172_new_n6488_));
AND2X2 AND2X2_3832 ( .A(core__abc_22172_new_n6490_), .B(core__abc_22172_new_n6485_), .Y(core__abc_22172_new_n6491_));
AND2X2 AND2X2_3833 ( .A(core__abc_22172_new_n6489_), .B(core__abc_22172_new_n4951_), .Y(core__abc_22172_new_n6493_));
AND2X2 AND2X2_3834 ( .A(core__abc_22172_new_n6492_), .B(core__abc_22172_new_n6494_), .Y(core__abc_22172_new_n6495_));
AND2X2 AND2X2_3835 ( .A(core__abc_22172_new_n6497_), .B(core__abc_22172_new_n6498_), .Y(core__abc_22172_new_n6499_));
AND2X2 AND2X2_3836 ( .A(core__abc_22172_new_n6500_), .B(core__abc_22172_new_n4909_), .Y(core__abc_22172_new_n6501_));
AND2X2 AND2X2_3837 ( .A(core__abc_22172_new_n6499_), .B(core__abc_22172_new_n4908_), .Y(core__abc_22172_new_n6502_));
AND2X2 AND2X2_3838 ( .A(core__abc_22172_new_n6495_), .B(core__abc_22172_new_n6504_), .Y(core__abc_22172_new_n6505_));
AND2X2 AND2X2_3839 ( .A(core__abc_22172_new_n6484_), .B(core__abc_22172_new_n6505_), .Y(core__abc_22172_new_n6506_));
AND2X2 AND2X2_384 ( .A(_abc_19873_new_n925_), .B(word2_reg_30_), .Y(_abc_19873_new_n1571_));
AND2X2 AND2X2_3840 ( .A(core__abc_22172_new_n6275_), .B(core_v1_reg_14_), .Y(core__abc_22172_new_n6508_));
AND2X2 AND2X2_3841 ( .A(core__abc_22172_new_n6509_), .B(core__abc_22172_new_n6507_), .Y(core__abc_22172_new_n6510_));
AND2X2 AND2X2_3842 ( .A(core__abc_22172_new_n6512_), .B(core__abc_22172_new_n6514_), .Y(core__abc_22172_new_n6515_));
AND2X2 AND2X2_3843 ( .A(core__abc_22172_new_n6517_), .B(core__abc_22172_new_n6518_), .Y(core__abc_22172_new_n6519_));
AND2X2 AND2X2_3844 ( .A(core__abc_22172_new_n6520_), .B(core__abc_22172_new_n4801_), .Y(core__abc_22172_new_n6521_));
AND2X2 AND2X2_3845 ( .A(core__abc_22172_new_n6519_), .B(core__abc_22172_new_n4800_), .Y(core__abc_22172_new_n6522_));
AND2X2 AND2X2_3846 ( .A(core__abc_22172_new_n6515_), .B(core__abc_22172_new_n6524_), .Y(core__abc_22172_new_n6525_));
AND2X2 AND2X2_3847 ( .A(core__abc_22172_new_n6199_), .B(core__abc_22172_new_n6527_), .Y(core__abc_22172_new_n6528_));
AND2X2 AND2X2_3848 ( .A(core__abc_22172_new_n6200_), .B(core_v1_reg_12_), .Y(core__abc_22172_new_n6529_));
AND2X2 AND2X2_3849 ( .A(core__abc_22172_new_n6531_), .B(core__abc_22172_new_n6526_), .Y(core__abc_22172_new_n6532_));
AND2X2 AND2X2_385 ( .A(_abc_19873_new_n907_), .B(word1_reg_30_), .Y(_abc_19873_new_n1572_));
AND2X2 AND2X2_3850 ( .A(core__abc_22172_new_n6535_), .B(core__abc_22172_new_n6536_), .Y(core__abc_22172_new_n6537_));
AND2X2 AND2X2_3851 ( .A(core__abc_22172_new_n6538_), .B(core__abc_22172_new_n4701_), .Y(core__abc_22172_new_n6539_));
AND2X2 AND2X2_3852 ( .A(core__abc_22172_new_n6530_), .B(core__abc_22172_new_n4743_), .Y(core__abc_22172_new_n6541_));
AND2X2 AND2X2_3853 ( .A(core__abc_22172_new_n6533_), .B(core__abc_22172_new_n6542_), .Y(core__abc_22172_new_n6543_));
AND2X2 AND2X2_3854 ( .A(core__abc_22172_new_n6525_), .B(core__abc_22172_new_n6544_), .Y(core__abc_22172_new_n6545_));
AND2X2 AND2X2_3855 ( .A(core__abc_22172_new_n6512_), .B(core__abc_22172_new_n6547_), .Y(core__abc_22172_new_n6548_));
AND2X2 AND2X2_3856 ( .A(core__abc_22172_new_n6506_), .B(core__abc_22172_new_n6551_), .Y(core__abc_22172_new_n6552_));
AND2X2 AND2X2_3857 ( .A(core__abc_22172_new_n6553_), .B(core__abc_22172_new_n6494_), .Y(core__abc_22172_new_n6554_));
AND2X2 AND2X2_3858 ( .A(core__abc_22172_new_n6484_), .B(core__abc_22172_new_n6554_), .Y(core__abc_22172_new_n6555_));
AND2X2 AND2X2_3859 ( .A(core__abc_22172_new_n6474_), .B(core__abc_22172_new_n6557_), .Y(core__abc_22172_new_n6558_));
AND2X2 AND2X2_386 ( .A(_abc_19873_new_n912_), .B(word3_reg_30_), .Y(_abc_19873_new_n1573_));
AND2X2 AND2X2_3860 ( .A(core__abc_22172_new_n6533_), .B(core__abc_22172_new_n6562_), .Y(core__abc_22172_new_n6563_));
AND2X2 AND2X2_3861 ( .A(core__abc_22172_new_n6537_), .B(core__abc_22172_new_n4700_), .Y(core__abc_22172_new_n6564_));
AND2X2 AND2X2_3862 ( .A(core__abc_22172_new_n6563_), .B(core__abc_22172_new_n6566_), .Y(core__abc_22172_new_n6567_));
AND2X2 AND2X2_3863 ( .A(core__abc_22172_new_n6525_), .B(core__abc_22172_new_n6567_), .Y(core__abc_22172_new_n6568_));
AND2X2 AND2X2_3864 ( .A(core__abc_22172_new_n6506_), .B(core__abc_22172_new_n6568_), .Y(core__abc_22172_new_n6569_));
AND2X2 AND2X2_3865 ( .A(core__abc_22172_new_n6108_), .B(core__abc_22172_new_n6570_), .Y(core__abc_22172_new_n6571_));
AND2X2 AND2X2_3866 ( .A(core__abc_22172_new_n6572_), .B(core__abc_22172_new_n6573_), .Y(core__abc_22172_new_n6574_));
AND2X2 AND2X2_3867 ( .A(core__abc_22172_new_n6576_), .B(core__abc_22172_new_n6577_), .Y(core__abc_22172_new_n6578_));
AND2X2 AND2X2_3868 ( .A(core__abc_22172_new_n6580_), .B(core__abc_22172_new_n6581_), .Y(core__abc_22172_new_n6582_));
AND2X2 AND2X2_3869 ( .A(core__abc_22172_new_n6583_), .B(core__abc_22172_new_n4590_), .Y(core__abc_22172_new_n6584_));
AND2X2 AND2X2_387 ( .A(_abc_19873_new_n919_), .B(core_mi_62_), .Y(_abc_19873_new_n1576_));
AND2X2 AND2X2_3870 ( .A(core__abc_22172_new_n6582_), .B(core__abc_22172_new_n4589_), .Y(core__abc_22172_new_n6585_));
AND2X2 AND2X2_3871 ( .A(core__abc_22172_new_n6578_), .B(core__abc_22172_new_n6587_), .Y(core__abc_22172_new_n6588_));
AND2X2 AND2X2_3872 ( .A(core__abc_22172_new_n6033_), .B(core__abc_22172_new_n6589_), .Y(core__abc_22172_new_n6590_));
AND2X2 AND2X2_3873 ( .A(core__abc_22172_new_n6034_), .B(core_v1_reg_8_), .Y(core__abc_22172_new_n6591_));
AND2X2 AND2X2_3874 ( .A(core__abc_22172_new_n6592_), .B(core__abc_22172_new_n4533_), .Y(core__abc_22172_new_n6594_));
AND2X2 AND2X2_3875 ( .A(core__abc_22172_new_n6595_), .B(core__abc_22172_new_n6593_), .Y(core__abc_22172_new_n6596_));
AND2X2 AND2X2_3876 ( .A(core__abc_22172_new_n6598_), .B(core__abc_22172_new_n6599_), .Y(core__abc_22172_new_n6600_));
AND2X2 AND2X2_3877 ( .A(core__abc_22172_new_n6601_), .B(core__abc_22172_new_n4480_), .Y(core__abc_22172_new_n6602_));
AND2X2 AND2X2_3878 ( .A(core__abc_22172_new_n6600_), .B(core__abc_22172_new_n4479_), .Y(core__abc_22172_new_n6603_));
AND2X2 AND2X2_3879 ( .A(core__abc_22172_new_n6596_), .B(core__abc_22172_new_n6605_), .Y(core__abc_22172_new_n6606_));
AND2X2 AND2X2_388 ( .A(_abc_19873_new_n930_), .B(word0_reg_30_), .Y(_abc_19873_new_n1577_));
AND2X2 AND2X2_3880 ( .A(core__abc_22172_new_n6588_), .B(core__abc_22172_new_n6606_), .Y(core__abc_22172_new_n6607_));
AND2X2 AND2X2_3881 ( .A(core__abc_22172_new_n6610_), .B(core__abc_22172_new_n6609_), .Y(core__abc_22172_new_n6611_));
AND2X2 AND2X2_3882 ( .A(core__abc_22172_new_n6612_), .B(core__abc_22172_new_n4353_), .Y(core__abc_22172_new_n6613_));
AND2X2 AND2X2_3883 ( .A(core__abc_22172_new_n6611_), .B(core__abc_22172_new_n4355_), .Y(core__abc_22172_new_n6614_));
AND2X2 AND2X2_3884 ( .A(core__abc_22172_new_n5955_), .B(core__abc_22172_new_n6617_), .Y(core__abc_22172_new_n6618_));
AND2X2 AND2X2_3885 ( .A(core__abc_22172_new_n5954_), .B(core_v1_reg_6_), .Y(core__abc_22172_new_n6619_));
AND2X2 AND2X2_3886 ( .A(core__abc_22172_new_n6623_), .B(core__abc_22172_new_n6621_), .Y(core__abc_22172_new_n6624_));
AND2X2 AND2X2_3887 ( .A(core__abc_22172_new_n6624_), .B(core__abc_22172_new_n6616_), .Y(core__abc_22172_new_n6625_));
AND2X2 AND2X2_3888 ( .A(core__abc_22172_new_n5881_), .B(core__abc_22172_new_n6626_), .Y(core__abc_22172_new_n6627_));
AND2X2 AND2X2_3889 ( .A(core__abc_22172_new_n6628_), .B(core__abc_22172_new_n6629_), .Y(core__abc_22172_new_n6630_));
AND2X2 AND2X2_389 ( .A(_abc_19873_new_n928_), .B(core_key_62_), .Y(_abc_19873_new_n1579_));
AND2X2 AND2X2_3890 ( .A(core__abc_22172_new_n6630_), .B(core__abc_22172_new_n4289_), .Y(core__abc_22172_new_n6631_));
AND2X2 AND2X2_3891 ( .A(core__abc_22172_new_n6634_), .B(core__abc_22172_new_n6635_), .Y(core__abc_22172_new_n6636_));
AND2X2 AND2X2_3892 ( .A(core__abc_22172_new_n6637_), .B(core__abc_22172_new_n4225_), .Y(core__abc_22172_new_n6638_));
AND2X2 AND2X2_3893 ( .A(core__abc_22172_new_n6640_), .B(core__abc_22172_new_n4287_), .Y(core__abc_22172_new_n6641_));
AND2X2 AND2X2_3894 ( .A(core__abc_22172_new_n6642_), .B(core__abc_22172_new_n6632_), .Y(core__abc_22172_new_n6643_));
AND2X2 AND2X2_3895 ( .A(core__abc_22172_new_n6625_), .B(core__abc_22172_new_n6644_), .Y(core__abc_22172_new_n6645_));
AND2X2 AND2X2_3896 ( .A(core__abc_22172_new_n6621_), .B(core__abc_22172_new_n6646_), .Y(core__abc_22172_new_n6647_));
AND2X2 AND2X2_3897 ( .A(core__abc_22172_new_n6648_), .B(core__abc_22172_new_n6623_), .Y(core__abc_22172_new_n6649_));
AND2X2 AND2X2_3898 ( .A(core__abc_22172_new_n6607_), .B(core__abc_22172_new_n6650_), .Y(core__abc_22172_new_n6651_));
AND2X2 AND2X2_3899 ( .A(core__abc_22172_new_n6593_), .B(core__abc_22172_new_n6652_), .Y(core__abc_22172_new_n6653_));
AND2X2 AND2X2_39 ( .A(_abc_19873_new_n893_), .B(_abc_19873_new_n918_), .Y(_abc_19873_new_n923_));
AND2X2 AND2X2_390 ( .A(_abc_19873_new_n901_), .B(core_key_30_), .Y(_abc_19873_new_n1580_));
AND2X2 AND2X2_3900 ( .A(core__abc_22172_new_n6588_), .B(core__abc_22172_new_n6655_), .Y(core__abc_22172_new_n6656_));
AND2X2 AND2X2_3901 ( .A(core__abc_22172_new_n6577_), .B(core__abc_22172_new_n6584_), .Y(core__abc_22172_new_n6658_));
AND2X2 AND2X2_3902 ( .A(core__abc_22172_new_n5793_), .B(core__abc_22172_new_n6662_), .Y(core__abc_22172_new_n6663_));
AND2X2 AND2X2_3903 ( .A(core__abc_22172_new_n5791_), .B(core_v1_reg_2_), .Y(core__abc_22172_new_n6664_));
AND2X2 AND2X2_3904 ( .A(core__abc_22172_new_n6669_), .B(core__abc_22172_new_n6666_), .Y(core__abc_22172_new_n6670_));
AND2X2 AND2X2_3905 ( .A(core__abc_22172_new_n6672_), .B(core__abc_22172_new_n6671_), .Y(core__abc_22172_new_n6673_));
AND2X2 AND2X2_3906 ( .A(core__abc_22172_new_n6674_), .B(core__abc_22172_new_n4086_), .Y(core__abc_22172_new_n6675_));
AND2X2 AND2X2_3907 ( .A(core__abc_22172_new_n6673_), .B(core__abc_22172_new_n4085_), .Y(core__abc_22172_new_n6676_));
AND2X2 AND2X2_3908 ( .A(core__abc_22172_new_n6670_), .B(core__abc_22172_new_n6678_), .Y(core__abc_22172_new_n6679_));
AND2X2 AND2X2_3909 ( .A(core__abc_22172_new_n5716_), .B(core__abc_22172_new_n6680_), .Y(core__abc_22172_new_n6681_));
AND2X2 AND2X2_391 ( .A(_abc_19873_new_n1584_), .B(_abc_19873_new_n937_), .Y(\read_data[30] ));
AND2X2 AND2X2_3910 ( .A(core__abc_22172_new_n5717_), .B(core_v1_reg_0_), .Y(core__abc_22172_new_n6682_));
AND2X2 AND2X2_3911 ( .A(core__abc_22172_new_n6683_), .B(core__abc_22172_new_n4008_), .Y(core__abc_22172_new_n6684_));
AND2X2 AND2X2_3912 ( .A(core__abc_22172_new_n6686_), .B(core__abc_22172_new_n4010_), .Y(core__abc_22172_new_n6687_));
AND2X2 AND2X2_3913 ( .A(core__abc_22172_new_n6689_), .B(core__abc_22172_new_n6690_), .Y(core__abc_22172_new_n6691_));
AND2X2 AND2X2_3914 ( .A(core__abc_22172_new_n6692_), .B(core__abc_22172_new_n3954_), .Y(core__abc_22172_new_n6693_));
AND2X2 AND2X2_3915 ( .A(core__abc_22172_new_n6688_), .B(core__abc_22172_new_n6694_), .Y(core__abc_22172_new_n6695_));
AND2X2 AND2X2_3916 ( .A(core__abc_22172_new_n6696_), .B(core__abc_22172_new_n6685_), .Y(core__abc_22172_new_n6697_));
AND2X2 AND2X2_3917 ( .A(core__abc_22172_new_n6679_), .B(core__abc_22172_new_n6697_), .Y(core__abc_22172_new_n6698_));
AND2X2 AND2X2_3918 ( .A(core__abc_22172_new_n6669_), .B(core__abc_22172_new_n6675_), .Y(core__abc_22172_new_n6700_));
AND2X2 AND2X2_3919 ( .A(core__abc_22172_new_n6688_), .B(core__abc_22172_new_n6685_), .Y(core__abc_22172_new_n6703_));
AND2X2 AND2X2_392 ( .A(_abc_19873_new_n881_), .B(core_key_127_), .Y(_abc_19873_new_n1586_));
AND2X2 AND2X2_3920 ( .A(core__abc_22172_new_n6691_), .B(core__abc_22172_new_n3953_), .Y(core__abc_22172_new_n6704_));
AND2X2 AND2X2_3921 ( .A(core__abc_22172_new_n6703_), .B(core__abc_22172_new_n6706_), .Y(core__abc_22172_new_n6707_));
AND2X2 AND2X2_3922 ( .A(core__abc_22172_new_n6679_), .B(core__abc_22172_new_n6707_), .Y(core__abc_22172_new_n6708_));
AND2X2 AND2X2_3923 ( .A(core__abc_22172_new_n5634_), .B(core_v1_reg_62_), .Y(core__abc_22172_new_n6710_));
AND2X2 AND2X2_3924 ( .A(core__abc_22172_new_n6711_), .B(core__abc_22172_new_n6709_), .Y(core__abc_22172_new_n6712_));
AND2X2 AND2X2_3925 ( .A(core__abc_22172_new_n6718_), .B(core__abc_22172_new_n6719_), .Y(core__abc_22172_new_n6720_));
AND2X2 AND2X2_3926 ( .A(core__abc_22172_new_n6721_), .B(core__abc_22172_new_n3827_), .Y(core__abc_22172_new_n6722_));
AND2X2 AND2X2_3927 ( .A(core__abc_22172_new_n6716_), .B(core__abc_22172_new_n6722_), .Y(core__abc_22172_new_n6723_));
AND2X2 AND2X2_3928 ( .A(core__abc_22172_new_n6714_), .B(core__abc_22172_new_n6716_), .Y(core__abc_22172_new_n6725_));
AND2X2 AND2X2_3929 ( .A(core__abc_22172_new_n6720_), .B(core__abc_22172_new_n3826_), .Y(core__abc_22172_new_n6726_));
AND2X2 AND2X2_393 ( .A(_abc_19873_new_n916_), .B(core_key_95_), .Y(_abc_19873_new_n1587_));
AND2X2 AND2X2_3930 ( .A(core__abc_22172_new_n6725_), .B(core__abc_22172_new_n6728_), .Y(core__abc_22172_new_n6729_));
AND2X2 AND2X2_3931 ( .A(core__abc_22172_new_n5545_), .B(core__abc_22172_new_n6730_), .Y(core__abc_22172_new_n6731_));
AND2X2 AND2X2_3932 ( .A(core__abc_22172_new_n5546_), .B(core_v1_reg_60_), .Y(core__abc_22172_new_n6732_));
AND2X2 AND2X2_3933 ( .A(core__abc_22172_new_n6733_), .B(core__abc_22172_new_n3748_), .Y(core__abc_22172_new_n6736_));
AND2X2 AND2X2_3934 ( .A(core__abc_22172_new_n6739_), .B(core__abc_22172_new_n6740_), .Y(core__abc_22172_new_n6741_));
AND2X2 AND2X2_3935 ( .A(core__abc_22172_new_n6742_), .B(core__abc_22172_new_n3694_), .Y(core__abc_22172_new_n6743_));
AND2X2 AND2X2_3936 ( .A(core__abc_22172_new_n6737_), .B(core__abc_22172_new_n6743_), .Y(core__abc_22172_new_n6744_));
AND2X2 AND2X2_3937 ( .A(core__abc_22172_new_n6729_), .B(core__abc_22172_new_n6745_), .Y(core__abc_22172_new_n6746_));
AND2X2 AND2X2_3938 ( .A(core__abc_22172_new_n5444_), .B(core_v1_reg_58_), .Y(core__abc_22172_new_n6749_));
AND2X2 AND2X2_3939 ( .A(core__abc_22172_new_n6750_), .B(core__abc_22172_new_n6748_), .Y(core__abc_22172_new_n6751_));
AND2X2 AND2X2_394 ( .A(_abc_19873_new_n912_), .B(word3_reg_31_), .Y(_abc_19873_new_n1589_));
AND2X2 AND2X2_3940 ( .A(core__abc_22172_new_n6751_), .B(core__abc_22172_new_n3618_), .Y(core__abc_22172_new_n6752_));
AND2X2 AND2X2_3941 ( .A(core__abc_22172_new_n6756_), .B(core__abc_22172_new_n6755_), .Y(core__abc_22172_new_n6757_));
AND2X2 AND2X2_3942 ( .A(core__abc_22172_new_n6758_), .B(core__abc_22172_new_n3557_), .Y(core__abc_22172_new_n6759_));
AND2X2 AND2X2_3943 ( .A(core__abc_22172_new_n6753_), .B(core__abc_22172_new_n6759_), .Y(core__abc_22172_new_n6760_));
AND2X2 AND2X2_3944 ( .A(core__abc_22172_new_n6762_), .B(core__abc_22172_new_n6753_), .Y(core__abc_22172_new_n6763_));
AND2X2 AND2X2_3945 ( .A(core__abc_22172_new_n6757_), .B(core__abc_22172_new_n3556_), .Y(core__abc_22172_new_n6764_));
AND2X2 AND2X2_3946 ( .A(core__abc_22172_new_n6763_), .B(core__abc_22172_new_n6766_), .Y(core__abc_22172_new_n6767_));
AND2X2 AND2X2_3947 ( .A(core__abc_22172_new_n5348_), .B(core__abc_22172_new_n6768_), .Y(core__abc_22172_new_n6769_));
AND2X2 AND2X2_3948 ( .A(core__abc_22172_new_n6770_), .B(core_v1_reg_56_), .Y(core__abc_22172_new_n6771_));
AND2X2 AND2X2_3949 ( .A(core__abc_22172_new_n6773_), .B(core__abc_22172_new_n3488_), .Y(core__abc_22172_new_n6774_));
AND2X2 AND2X2_395 ( .A(_abc_19873_new_n907_), .B(word1_reg_31_), .Y(_abc_19873_new_n1590_));
AND2X2 AND2X2_3950 ( .A(core__abc_22172_new_n6772_), .B(core__abc_22172_new_n3486_), .Y(core__abc_22172_new_n6775_));
AND2X2 AND2X2_3951 ( .A(core__abc_22172_new_n6778_), .B(core__abc_22172_new_n6779_), .Y(core__abc_22172_new_n6780_));
AND2X2 AND2X2_3952 ( .A(core__abc_22172_new_n6781_), .B(core__abc_22172_new_n3428_), .Y(core__abc_22172_new_n6782_));
AND2X2 AND2X2_3953 ( .A(core__abc_22172_new_n5254_), .B(core__abc_22172_new_n6783_), .Y(core__abc_22172_new_n6784_));
AND2X2 AND2X2_3954 ( .A(core__abc_22172_new_n6785_), .B(core_v1_reg_54_), .Y(core__abc_22172_new_n6786_));
AND2X2 AND2X2_3955 ( .A(core__abc_22172_new_n6788_), .B(core__abc_22172_new_n3376_), .Y(core__abc_22172_new_n6789_));
AND2X2 AND2X2_3956 ( .A(core__abc_22172_new_n6792_), .B(core__abc_22172_new_n6793_), .Y(core__abc_22172_new_n6794_));
AND2X2 AND2X2_3957 ( .A(core__abc_22172_new_n6798_), .B(core__abc_22172_new_n6799_), .Y(core__abc_22172_new_n6800_));
AND2X2 AND2X2_3958 ( .A(core__abc_22172_new_n1268_), .B(core_v1_reg_51_), .Y(core__abc_22172_new_n6803_));
AND2X2 AND2X2_3959 ( .A(core__abc_22172_new_n6804_), .B(core__abc_22172_new_n6805_), .Y(core__abc_22172_new_n6806_));
AND2X2 AND2X2_396 ( .A(_abc_19873_new_n930_), .B(word0_reg_31_), .Y(_abc_19873_new_n1591_));
AND2X2 AND2X2_3960 ( .A(core__abc_22172_new_n6807_), .B(core__abc_22172_new_n1266_), .Y(core__abc_22172_new_n6808_));
AND2X2 AND2X2_3961 ( .A(core__abc_22172_new_n6810_), .B(core__abc_22172_new_n6801_), .Y(core__abc_22172_new_n6811_));
AND2X2 AND2X2_3962 ( .A(core__abc_22172_new_n6811_), .B(core__abc_22172_new_n6808_), .Y(core__abc_22172_new_n6812_));
AND2X2 AND2X2_3963 ( .A(core__abc_22172_new_n6815_), .B(core__abc_22172_new_n6795_), .Y(core__abc_22172_new_n6816_));
AND2X2 AND2X2_3964 ( .A(core__abc_22172_new_n6813_), .B(core__abc_22172_new_n6816_), .Y(core__abc_22172_new_n6817_));
AND2X2 AND2X2_3965 ( .A(core__abc_22172_new_n6818_), .B(core__abc_22172_new_n6790_), .Y(core__abc_22172_new_n6819_));
AND2X2 AND2X2_3966 ( .A(core__abc_22172_new_n6780_), .B(core__abc_22172_new_n3426_), .Y(core__abc_22172_new_n6821_));
AND2X2 AND2X2_3967 ( .A(core__abc_22172_new_n6820_), .B(core__abc_22172_new_n6823_), .Y(core__abc_22172_new_n6824_));
AND2X2 AND2X2_3968 ( .A(core__abc_22172_new_n6825_), .B(core__abc_22172_new_n6776_), .Y(core__abc_22172_new_n6826_));
AND2X2 AND2X2_3969 ( .A(core__abc_22172_new_n6827_), .B(core__abc_22172_new_n6767_), .Y(core__abc_22172_new_n6828_));
AND2X2 AND2X2_397 ( .A(_abc_19873_new_n925_), .B(word2_reg_31_), .Y(_abc_19873_new_n1595_));
AND2X2 AND2X2_3970 ( .A(core__abc_22172_new_n6737_), .B(core__abc_22172_new_n6734_), .Y(core__abc_22172_new_n6830_));
AND2X2 AND2X2_3971 ( .A(core__abc_22172_new_n6741_), .B(core__abc_22172_new_n3693_), .Y(core__abc_22172_new_n6831_));
AND2X2 AND2X2_3972 ( .A(core__abc_22172_new_n6830_), .B(core__abc_22172_new_n6833_), .Y(core__abc_22172_new_n6834_));
AND2X2 AND2X2_3973 ( .A(core__abc_22172_new_n6729_), .B(core__abc_22172_new_n6834_), .Y(core__abc_22172_new_n6835_));
AND2X2 AND2X2_3974 ( .A(core__abc_22172_new_n6829_), .B(core__abc_22172_new_n6835_), .Y(core__abc_22172_new_n6836_));
AND2X2 AND2X2_3975 ( .A(core__abc_22172_new_n6837_), .B(core__abc_22172_new_n6708_), .Y(core__abc_22172_new_n6838_));
AND2X2 AND2X2_3976 ( .A(core__abc_22172_new_n6840_), .B(core__abc_22172_new_n6632_), .Y(core__abc_22172_new_n6841_));
AND2X2 AND2X2_3977 ( .A(core__abc_22172_new_n6636_), .B(core__abc_22172_new_n4224_), .Y(core__abc_22172_new_n6842_));
AND2X2 AND2X2_3978 ( .A(core__abc_22172_new_n6841_), .B(core__abc_22172_new_n6844_), .Y(core__abc_22172_new_n6845_));
AND2X2 AND2X2_3979 ( .A(core__abc_22172_new_n6625_), .B(core__abc_22172_new_n6845_), .Y(core__abc_22172_new_n6846_));
AND2X2 AND2X2_398 ( .A(_abc_19873_new_n928_), .B(core_key_63_), .Y(_abc_19873_new_n1596_));
AND2X2 AND2X2_3980 ( .A(core__abc_22172_new_n6607_), .B(core__abc_22172_new_n6846_), .Y(core__abc_22172_new_n6847_));
AND2X2 AND2X2_3981 ( .A(core__abc_22172_new_n6847_), .B(core__abc_22172_new_n6839_), .Y(core__abc_22172_new_n6848_));
AND2X2 AND2X2_3982 ( .A(core__abc_22172_new_n6849_), .B(core__abc_22172_new_n6569_), .Y(core__abc_22172_new_n6850_));
AND2X2 AND2X2_3983 ( .A(core__abc_22172_new_n6853_), .B(core__abc_22172_new_n6854_), .Y(core__abc_22172_new_n6855_));
AND2X2 AND2X2_3984 ( .A(core__abc_22172_new_n6856_), .B(core__abc_22172_new_n5110_), .Y(core__abc_22172_new_n6857_));
AND2X2 AND2X2_3985 ( .A(core__abc_22172_new_n6855_), .B(core__abc_22172_new_n5109_), .Y(core__abc_22172_new_n6858_));
AND2X2 AND2X2_3986 ( .A(core__abc_22172_new_n6851_), .B(core__abc_22172_new_n6860_), .Y(core__abc_22172_new_n6861_));
AND2X2 AND2X2_3987 ( .A(core__abc_22172_new_n6862_), .B(core__abc_22172_new_n6859_), .Y(core__abc_22172_new_n6863_));
AND2X2 AND2X2_3988 ( .A(core__abc_22172_new_n6865_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n6866_));
AND2X2 AND2X2_3989 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n6867_), .Y(core__abc_22172_new_n6868_));
AND2X2 AND2X2_399 ( .A(_abc_19873_new_n901_), .B(core_key_31_), .Y(_abc_19873_new_n1597_));
AND2X2 AND2X2_3990 ( .A(core__abc_22172_new_n6869_), .B(core__abc_22172_new_n6871_), .Y(core__abc_22172_new_n6872_));
AND2X2 AND2X2_3991 ( .A(core__abc_22172_new_n3196_), .B(core__abc_22172_new_n6872_), .Y(core__abc_22172_new_n6873_));
AND2X2 AND2X2_3992 ( .A(core__abc_22172_new_n6875_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n6876_));
AND2X2 AND2X2_3993 ( .A(core__abc_22172_new_n6878_), .B(core__abc_22172_new_n3197_), .Y(core__abc_22172_new_n6879_));
AND2X2 AND2X2_3994 ( .A(core__abc_22172_new_n6880_), .B(core_v2_reg_0_), .Y(core__abc_22172_new_n6881_));
AND2X2 AND2X2_3995 ( .A(core__abc_22172_new_n6882_), .B(reset_n), .Y(core__0v2_reg_63_0__0_));
AND2X2 AND2X2_3996 ( .A(core__abc_22172_new_n3239_), .B(core__abc_22172_new_n6885_), .Y(core__abc_22172_new_n6886_));
AND2X2 AND2X2_3997 ( .A(core__abc_22172_new_n6887_), .B(core__abc_22172_new_n6888_), .Y(core__abc_22172_new_n6889_));
AND2X2 AND2X2_3998 ( .A(core__abc_22172_new_n6889_), .B(core__abc_22172_new_n6884_), .Y(core__abc_22172_new_n6890_));
AND2X2 AND2X2_3999 ( .A(core__abc_22172_new_n6891_), .B(core__abc_22172_new_n5168_), .Y(core__abc_22172_new_n6892_));
AND2X2 AND2X2_4 ( .A(\addr[0] ), .B(\addr[1] ), .Y(_abc_19873_new_n876_));
AND2X2 AND2X2_40 ( .A(_abc_19873_new_n923_), .B(core_ready), .Y(_abc_19873_new_n924_));
AND2X2 AND2X2_400 ( .A(_abc_19873_new_n888_), .B(core_mi_31_), .Y(_abc_19873_new_n1599_));
AND2X2 AND2X2_4000 ( .A(core__abc_22172_new_n6895_), .B(core__abc_22172_new_n6894_), .Y(core__abc_22172_new_n6896_));
AND2X2 AND2X2_4001 ( .A(core__abc_22172_new_n6896_), .B(core__abc_22172_new_n6893_), .Y(core__abc_22172_new_n6897_));
AND2X2 AND2X2_4002 ( .A(core__abc_22172_new_n6901_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n6902_));
AND2X2 AND2X2_4003 ( .A(core__abc_22172_new_n3214_), .B(core_key_1_), .Y(core__abc_22172_new_n6903_));
AND2X2 AND2X2_4004 ( .A(core__abc_22172_new_n3196_), .B(core__abc_22172_new_n1280_), .Y(core__abc_22172_new_n6904_));
AND2X2 AND2X2_4005 ( .A(core__abc_22172_new_n6906_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n6907_));
AND2X2 AND2X2_4006 ( .A(core__abc_22172_new_n6880_), .B(core_v2_reg_1_), .Y(core__abc_22172_new_n6908_));
AND2X2 AND2X2_4007 ( .A(core__abc_22172_new_n6909_), .B(reset_n), .Y(core__0v2_reg_63_0__1_));
AND2X2 AND2X2_4008 ( .A(core__abc_22172_new_n6911_), .B(core__abc_22172_new_n6860_), .Y(core__abc_22172_new_n6912_));
AND2X2 AND2X2_4009 ( .A(core__abc_22172_new_n6851_), .B(core__abc_22172_new_n6912_), .Y(core__abc_22172_new_n6913_));
AND2X2 AND2X2_401 ( .A(_abc_19873_new_n919_), .B(core_mi_63_), .Y(_abc_19873_new_n1600_));
AND2X2 AND2X2_4010 ( .A(core__abc_22172_new_n6911_), .B(core__abc_22172_new_n6857_), .Y(core__abc_22172_new_n6914_));
AND2X2 AND2X2_4011 ( .A(core__abc_22172_new_n6919_), .B(core__abc_22172_new_n6918_), .Y(core__abc_22172_new_n6920_));
AND2X2 AND2X2_4012 ( .A(core__abc_22172_new_n6920_), .B(core__abc_22172_new_n5217_), .Y(core__abc_22172_new_n6921_));
AND2X2 AND2X2_4013 ( .A(core__abc_22172_new_n6922_), .B(core__abc_22172_new_n5218_), .Y(core__abc_22172_new_n6923_));
AND2X2 AND2X2_4014 ( .A(core__abc_22172_new_n6916_), .B(core__abc_22172_new_n6925_), .Y(core__abc_22172_new_n6926_));
AND2X2 AND2X2_4015 ( .A(core__abc_22172_new_n6927_), .B(core__abc_22172_new_n6928_), .Y(core__abc_22172_new_n6929_));
AND2X2 AND2X2_4016 ( .A(core__abc_22172_new_n6929_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n6930_));
AND2X2 AND2X2_4017 ( .A(core__abc_22172_new_n3214_), .B(core_key_2_), .Y(core__abc_22172_new_n6931_));
AND2X2 AND2X2_4018 ( .A(core__abc_22172_new_n3196_), .B(core__abc_22172_new_n1302_), .Y(core__abc_22172_new_n6932_));
AND2X2 AND2X2_4019 ( .A(core__abc_22172_new_n6934_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n6935_));
AND2X2 AND2X2_402 ( .A(_abc_19873_new_n1604_), .B(_abc_19873_new_n937_), .Y(\read_data[31] ));
AND2X2 AND2X2_4020 ( .A(core__abc_22172_new_n6880_), .B(core_v2_reg_2_), .Y(core__abc_22172_new_n6936_));
AND2X2 AND2X2_4021 ( .A(core__abc_22172_new_n6937_), .B(reset_n), .Y(core__0v2_reg_63_0__2_));
AND2X2 AND2X2_4022 ( .A(core__abc_22172_new_n6927_), .B(core__abc_22172_new_n6939_), .Y(core__abc_22172_new_n6940_));
AND2X2 AND2X2_4023 ( .A(core__abc_22172_new_n3369_), .B(core_v1_reg_22_), .Y(core__abc_22172_new_n6942_));
AND2X2 AND2X2_4024 ( .A(core__abc_22172_new_n6943_), .B(core__abc_22172_new_n6941_), .Y(core__abc_22172_new_n6944_));
AND2X2 AND2X2_4025 ( .A(core__abc_22172_new_n6944_), .B(core__abc_22172_new_n5259_), .Y(core__abc_22172_new_n6945_));
AND2X2 AND2X2_4026 ( .A(core__abc_22172_new_n6946_), .B(core__abc_22172_new_n5260_), .Y(core__abc_22172_new_n6947_));
AND2X2 AND2X2_4027 ( .A(core__abc_22172_new_n6940_), .B(core__abc_22172_new_n6948_), .Y(core__abc_22172_new_n6949_));
AND2X2 AND2X2_4028 ( .A(core__abc_22172_new_n6950_), .B(core__abc_22172_new_n6951_), .Y(core__abc_22172_new_n6952_));
AND2X2 AND2X2_4029 ( .A(core__abc_22172_new_n6952_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n6953_));
AND2X2 AND2X2_403 ( .A(core_siphash_valid_reg), .B(core_siphash_word_96_), .Y(_abc_19873_new_n1606_));
AND2X2 AND2X2_4030 ( .A(core__abc_22172_new_n3214_), .B(core_key_3_), .Y(core__abc_22172_new_n6954_));
AND2X2 AND2X2_4031 ( .A(core__abc_22172_new_n3196_), .B(core__abc_22172_new_n1319_), .Y(core__abc_22172_new_n6955_));
AND2X2 AND2X2_4032 ( .A(core__abc_22172_new_n6957_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n6958_));
AND2X2 AND2X2_4033 ( .A(core__abc_22172_new_n6880_), .B(core_v2_reg_3_), .Y(core__abc_22172_new_n6959_));
AND2X2 AND2X2_4034 ( .A(core__abc_22172_new_n6960_), .B(reset_n), .Y(core__0v2_reg_63_0__3_));
AND2X2 AND2X2_4035 ( .A(core__abc_22172_new_n6963_), .B(core__abc_22172_new_n6964_), .Y(core__abc_22172_new_n6965_));
AND2X2 AND2X2_4036 ( .A(core__abc_22172_new_n6965_), .B(core__abc_22172_new_n5312_), .Y(core__abc_22172_new_n6966_));
AND2X2 AND2X2_4037 ( .A(core__abc_22172_new_n6967_), .B(core__abc_22172_new_n5313_), .Y(core__abc_22172_new_n6968_));
AND2X2 AND2X2_4038 ( .A(core__abc_22172_new_n6971_), .B(core__abc_22172_new_n6939_), .Y(core__abc_22172_new_n6972_));
AND2X2 AND2X2_4039 ( .A(core__abc_22172_new_n6927_), .B(core__abc_22172_new_n6972_), .Y(core__abc_22172_new_n6973_));
AND2X2 AND2X2_404 ( .A(_abc_19873_new_n1607_), .B(word3_reg_0_), .Y(_abc_19873_new_n1608_));
AND2X2 AND2X2_4040 ( .A(core__abc_22172_new_n6975_), .B(core__abc_22172_new_n6970_), .Y(core__abc_22172_new_n6976_));
AND2X2 AND2X2_4041 ( .A(core__abc_22172_new_n6974_), .B(core__abc_22172_new_n6969_), .Y(core__abc_22172_new_n6977_));
AND2X2 AND2X2_4042 ( .A(core__abc_22172_new_n6979_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n6980_));
AND2X2 AND2X2_4043 ( .A(core__abc_22172_new_n3214_), .B(core_key_4_), .Y(core__abc_22172_new_n6981_));
AND2X2 AND2X2_4044 ( .A(core__abc_22172_new_n6982_), .B(core__abc_22172_new_n6983_), .Y(core__abc_22172_new_n6984_));
AND2X2 AND2X2_4045 ( .A(core__abc_22172_new_n3196_), .B(core__abc_22172_new_n6984_), .Y(core__abc_22172_new_n6985_));
AND2X2 AND2X2_4046 ( .A(core__abc_22172_new_n6987_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n6988_));
AND2X2 AND2X2_4047 ( .A(core__abc_22172_new_n6880_), .B(core_v2_reg_4_), .Y(core__abc_22172_new_n6989_));
AND2X2 AND2X2_4048 ( .A(core__abc_22172_new_n6990_), .B(reset_n), .Y(core__0v2_reg_63_0__4_));
AND2X2 AND2X2_4049 ( .A(core__abc_22172_new_n6994_), .B(core__abc_22172_new_n6993_), .Y(core__abc_22172_new_n6995_));
AND2X2 AND2X2_405 ( .A(_abc_19873_new_n1609_), .B(reset_n), .Y(_0word3_reg_31_0__0_));
AND2X2 AND2X2_4050 ( .A(core__abc_22172_new_n3480_), .B(core_v1_reg_24_), .Y(core__abc_22172_new_n6996_));
AND2X2 AND2X2_4051 ( .A(core__abc_22172_new_n6997_), .B(core__abc_22172_new_n5353_), .Y(core__abc_22172_new_n6998_));
AND2X2 AND2X2_4052 ( .A(core__abc_22172_new_n6999_), .B(core__abc_22172_new_n7000_), .Y(core__abc_22172_new_n7001_));
AND2X2 AND2X2_4053 ( .A(core__abc_22172_new_n6992_), .B(core__abc_22172_new_n7002_), .Y(core__abc_22172_new_n7003_));
AND2X2 AND2X2_4054 ( .A(core__abc_22172_new_n7004_), .B(core__abc_22172_new_n7005_), .Y(core__abc_22172_new_n7006_));
AND2X2 AND2X2_4055 ( .A(core__abc_22172_new_n7007_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n7008_));
AND2X2 AND2X2_4056 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n7009_), .Y(core__abc_22172_new_n7010_));
AND2X2 AND2X2_4057 ( .A(core__abc_22172_new_n3196_), .B(core__abc_22172_new_n1356_), .Y(core__abc_22172_new_n7011_));
AND2X2 AND2X2_4058 ( .A(core__abc_22172_new_n7013_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n7014_));
AND2X2 AND2X2_4059 ( .A(core__abc_22172_new_n6880_), .B(core_v2_reg_5_), .Y(core__abc_22172_new_n7015_));
AND2X2 AND2X2_406 ( .A(core_siphash_valid_reg), .B(core_siphash_word_97_), .Y(_abc_19873_new_n1611_));
AND2X2 AND2X2_4060 ( .A(core__abc_22172_new_n7016_), .B(reset_n), .Y(core__0v2_reg_63_0__5_));
AND2X2 AND2X2_4061 ( .A(core__abc_22172_new_n7019_), .B(core__abc_22172_new_n7020_), .Y(core__abc_22172_new_n7021_));
AND2X2 AND2X2_4062 ( .A(core__abc_22172_new_n7021_), .B(core__abc_22172_new_n5407_), .Y(core__abc_22172_new_n7022_));
AND2X2 AND2X2_4063 ( .A(core__abc_22172_new_n7023_), .B(core__abc_22172_new_n5408_), .Y(core__abc_22172_new_n7024_));
AND2X2 AND2X2_4064 ( .A(core__abc_22172_new_n7000_), .B(core__abc_22172_new_n7026_), .Y(core__abc_22172_new_n7027_));
AND2X2 AND2X2_4065 ( .A(core__abc_22172_new_n7001_), .B(core__abc_22172_new_n6970_), .Y(core__abc_22172_new_n7029_));
AND2X2 AND2X2_4066 ( .A(core__abc_22172_new_n7031_), .B(core__abc_22172_new_n7028_), .Y(core__abc_22172_new_n7032_));
AND2X2 AND2X2_4067 ( .A(core__abc_22172_new_n7032_), .B(core__abc_22172_new_n7025_), .Y(core__abc_22172_new_n7035_));
AND2X2 AND2X2_4068 ( .A(core__abc_22172_new_n7037_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n7038_));
AND2X2 AND2X2_4069 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n7039_), .Y(core__abc_22172_new_n7040_));
AND2X2 AND2X2_407 ( .A(_abc_19873_new_n1607_), .B(word3_reg_1_), .Y(_abc_19873_new_n1612_));
AND2X2 AND2X2_4070 ( .A(core__abc_22172_new_n3196_), .B(core__abc_22172_new_n1375_), .Y(core__abc_22172_new_n7041_));
AND2X2 AND2X2_4071 ( .A(core__abc_22172_new_n7043_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n7044_));
AND2X2 AND2X2_4072 ( .A(core__abc_22172_new_n6880_), .B(core_v2_reg_6_), .Y(core__abc_22172_new_n7045_));
AND2X2 AND2X2_4073 ( .A(core__abc_22172_new_n7046_), .B(reset_n), .Y(core__0v2_reg_63_0__6_));
AND2X2 AND2X2_4074 ( .A(core__abc_22172_new_n7033_), .B(core__abc_22172_new_n7048_), .Y(core__abc_22172_new_n7049_));
AND2X2 AND2X2_4075 ( .A(core__abc_22172_new_n3609_), .B(core__abc_22172_new_n7051_), .Y(core__abc_22172_new_n7052_));
AND2X2 AND2X2_4076 ( .A(core__abc_22172_new_n3610_), .B(core_v1_reg_26_), .Y(core__abc_22172_new_n7053_));
AND2X2 AND2X2_4077 ( .A(core__abc_22172_new_n7055_), .B(core__abc_22172_new_n7050_), .Y(core__abc_22172_new_n7056_));
AND2X2 AND2X2_4078 ( .A(core__abc_22172_new_n7054_), .B(core__abc_22172_new_n5449_), .Y(core__abc_22172_new_n7057_));
AND2X2 AND2X2_4079 ( .A(core__abc_22172_new_n7049_), .B(core__abc_22172_new_n7058_), .Y(core__abc_22172_new_n7059_));
AND2X2 AND2X2_408 ( .A(_abc_19873_new_n1613_), .B(reset_n), .Y(_0word3_reg_31_0__1_));
AND2X2 AND2X2_4080 ( .A(core__abc_22172_new_n7060_), .B(core__abc_22172_new_n7061_), .Y(core__abc_22172_new_n7062_));
AND2X2 AND2X2_4081 ( .A(core__abc_22172_new_n7062_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n7063_));
AND2X2 AND2X2_4082 ( .A(core__abc_22172_new_n3214_), .B(core_key_7_), .Y(core__abc_22172_new_n7064_));
AND2X2 AND2X2_4083 ( .A(core__abc_22172_new_n3196_), .B(core__abc_22172_new_n1394_), .Y(core__abc_22172_new_n7065_));
AND2X2 AND2X2_4084 ( .A(core__abc_22172_new_n7067_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n7068_));
AND2X2 AND2X2_4085 ( .A(core__abc_22172_new_n6880_), .B(core_v2_reg_7_), .Y(core__abc_22172_new_n7069_));
AND2X2 AND2X2_4086 ( .A(core__abc_22172_new_n7070_), .B(reset_n), .Y(core__0v2_reg_63_0__7_));
AND2X2 AND2X2_4087 ( .A(core__abc_22172_new_n7073_), .B(core__abc_22172_new_n6912_), .Y(core__abc_22172_new_n7074_));
AND2X2 AND2X2_4088 ( .A(core__abc_22172_new_n7077_), .B(core__abc_22172_new_n7074_), .Y(core__abc_22172_new_n7078_));
AND2X2 AND2X2_4089 ( .A(core__abc_22172_new_n6851_), .B(core__abc_22172_new_n7078_), .Y(core__abc_22172_new_n7079_));
AND2X2 AND2X2_409 ( .A(core_siphash_valid_reg), .B(core_siphash_word_98_), .Y(_abc_19873_new_n1615_));
AND2X2 AND2X2_4090 ( .A(core__abc_22172_new_n7073_), .B(core__abc_22172_new_n6915_), .Y(core__abc_22172_new_n7081_));
AND2X2 AND2X2_4091 ( .A(core__abc_22172_new_n7082_), .B(core__abc_22172_new_n7080_), .Y(core__abc_22172_new_n7083_));
AND2X2 AND2X2_4092 ( .A(core__abc_22172_new_n7086_), .B(core__abc_22172_new_n7085_), .Y(core__abc_22172_new_n7087_));
AND2X2 AND2X2_4093 ( .A(core__abc_22172_new_n7089_), .B(core__abc_22172_new_n7088_), .Y(core__abc_22172_new_n7090_));
AND2X2 AND2X2_4094 ( .A(core__abc_22172_new_n7084_), .B(core__abc_22172_new_n7090_), .Y(core__abc_22172_new_n7091_));
AND2X2 AND2X2_4095 ( .A(core__abc_22172_new_n7095_), .B(core__abc_22172_new_n7096_), .Y(core__abc_22172_new_n7097_));
AND2X2 AND2X2_4096 ( .A(core__abc_22172_new_n7097_), .B(core__abc_22172_new_n5502_), .Y(core__abc_22172_new_n7098_));
AND2X2 AND2X2_4097 ( .A(core__abc_22172_new_n7099_), .B(core__abc_22172_new_n5503_), .Y(core__abc_22172_new_n7100_));
AND2X2 AND2X2_4098 ( .A(core__abc_22172_new_n7093_), .B(core__abc_22172_new_n7102_), .Y(core__abc_22172_new_n7103_));
AND2X2 AND2X2_4099 ( .A(core__abc_22172_new_n7104_), .B(core__abc_22172_new_n7101_), .Y(core__abc_22172_new_n7105_));
AND2X2 AND2X2_41 ( .A(_abc_19873_new_n906_), .B(_abc_19873_new_n915_), .Y(_abc_19873_new_n925_));
AND2X2 AND2X2_410 ( .A(_abc_19873_new_n1607_), .B(word3_reg_2_), .Y(_abc_19873_new_n1616_));
AND2X2 AND2X2_4100 ( .A(core__abc_22172_new_n7107_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n7108_));
AND2X2 AND2X2_4101 ( .A(core__abc_22172_new_n3214_), .B(core_key_8_), .Y(core__abc_22172_new_n7109_));
AND2X2 AND2X2_4102 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_8_), .Y(core__abc_22172_new_n7110_));
AND2X2 AND2X2_4103 ( .A(core__abc_22172_new_n7115_), .B(reset_n), .Y(core__abc_22172_new_n7116_));
AND2X2 AND2X2_4104 ( .A(core__abc_22172_new_n7113_), .B(core__abc_22172_new_n7116_), .Y(core__0v2_reg_63_0__8_));
AND2X2 AND2X2_4105 ( .A(core__abc_22172_new_n7119_), .B(core__abc_22172_new_n7118_), .Y(core__abc_22172_new_n7120_));
AND2X2 AND2X2_4106 ( .A(core__abc_22172_new_n3742_), .B(core_v1_reg_28_), .Y(core__abc_22172_new_n7121_));
AND2X2 AND2X2_4107 ( .A(core__abc_22172_new_n7122_), .B(core__abc_22172_new_n5552_), .Y(core__abc_22172_new_n7124_));
AND2X2 AND2X2_4108 ( .A(core__abc_22172_new_n7125_), .B(core__abc_22172_new_n7123_), .Y(core__abc_22172_new_n7126_));
AND2X2 AND2X2_4109 ( .A(core__abc_22172_new_n7129_), .B(core__abc_22172_new_n7128_), .Y(core__abc_22172_new_n7130_));
AND2X2 AND2X2_411 ( .A(_abc_19873_new_n1617_), .B(reset_n), .Y(_0word3_reg_31_0__2_));
AND2X2 AND2X2_4110 ( .A(core__abc_22172_new_n7130_), .B(core__abc_22172_new_n7127_), .Y(core__abc_22172_new_n7131_));
AND2X2 AND2X2_4111 ( .A(core__abc_22172_new_n7135_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n7136_));
AND2X2 AND2X2_4112 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n7137_), .Y(core__abc_22172_new_n7138_));
AND2X2 AND2X2_4113 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_9_), .Y(core__abc_22172_new_n7139_));
AND2X2 AND2X2_4114 ( .A(core__abc_22172_new_n7143_), .B(reset_n), .Y(core__abc_22172_new_n7144_));
AND2X2 AND2X2_4115 ( .A(core__abc_22172_new_n7142_), .B(core__abc_22172_new_n7144_), .Y(core__0v2_reg_63_0__9_));
AND2X2 AND2X2_4116 ( .A(core__abc_22172_new_n7126_), .B(core__abc_22172_new_n7102_), .Y(core__abc_22172_new_n7146_));
AND2X2 AND2X2_4117 ( .A(core__abc_22172_new_n7093_), .B(core__abc_22172_new_n7146_), .Y(core__abc_22172_new_n7147_));
AND2X2 AND2X2_4118 ( .A(core__abc_22172_new_n7148_), .B(core__abc_22172_new_n7123_), .Y(core__abc_22172_new_n7149_));
AND2X2 AND2X2_4119 ( .A(core__abc_22172_new_n7153_), .B(core__abc_22172_new_n7154_), .Y(core__abc_22172_new_n7155_));
AND2X2 AND2X2_412 ( .A(core_siphash_valid_reg), .B(core_siphash_word_99_), .Y(_abc_19873_new_n1619_));
AND2X2 AND2X2_4120 ( .A(core__abc_22172_new_n7156_), .B(core__abc_22172_new_n5595_), .Y(core__abc_22172_new_n7157_));
AND2X2 AND2X2_4121 ( .A(core__abc_22172_new_n7155_), .B(core__abc_22172_new_n5594_), .Y(core__abc_22172_new_n7158_));
AND2X2 AND2X2_4122 ( .A(core__abc_22172_new_n7151_), .B(core__abc_22172_new_n7160_), .Y(core__abc_22172_new_n7161_));
AND2X2 AND2X2_4123 ( .A(core__abc_22172_new_n7162_), .B(core__abc_22172_new_n7163_), .Y(core__abc_22172_new_n7164_));
AND2X2 AND2X2_4124 ( .A(core__abc_22172_new_n7164_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n7165_));
AND2X2 AND2X2_4125 ( .A(core__abc_22172_new_n3214_), .B(core_key_10_), .Y(core__abc_22172_new_n7166_));
AND2X2 AND2X2_4126 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_10_), .Y(core__abc_22172_new_n7167_));
AND2X2 AND2X2_4127 ( .A(core__abc_22172_new_n7171_), .B(reset_n), .Y(core__abc_22172_new_n7172_));
AND2X2 AND2X2_4128 ( .A(core__abc_22172_new_n7170_), .B(core__abc_22172_new_n7172_), .Y(core__0v2_reg_63_0__10_));
AND2X2 AND2X2_4129 ( .A(core__abc_22172_new_n7162_), .B(core__abc_22172_new_n7174_), .Y(core__abc_22172_new_n7175_));
AND2X2 AND2X2_413 ( .A(_abc_19873_new_n1607_), .B(word3_reg_3_), .Y(_abc_19873_new_n1620_));
AND2X2 AND2X2_4130 ( .A(core__abc_22172_new_n3874_), .B(core__abc_22172_new_n7176_), .Y(core__abc_22172_new_n7177_));
AND2X2 AND2X2_4131 ( .A(core__abc_22172_new_n3875_), .B(core_v1_reg_30_), .Y(core__abc_22172_new_n7178_));
AND2X2 AND2X2_4132 ( .A(core__abc_22172_new_n7179_), .B(core__abc_22172_new_n3189_), .Y(core__abc_22172_new_n7181_));
AND2X2 AND2X2_4133 ( .A(core__abc_22172_new_n7182_), .B(core__abc_22172_new_n7180_), .Y(core__abc_22172_new_n7183_));
AND2X2 AND2X2_4134 ( .A(core__abc_22172_new_n7175_), .B(core__abc_22172_new_n7184_), .Y(core__abc_22172_new_n7185_));
AND2X2 AND2X2_4135 ( .A(core__abc_22172_new_n7186_), .B(core__abc_22172_new_n7187_), .Y(core__abc_22172_new_n7188_));
AND2X2 AND2X2_4136 ( .A(core__abc_22172_new_n7188_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n7189_));
AND2X2 AND2X2_4137 ( .A(core__abc_22172_new_n3214_), .B(core_key_11_), .Y(core__abc_22172_new_n7190_));
AND2X2 AND2X2_4138 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_11_), .Y(core__abc_22172_new_n7191_));
AND2X2 AND2X2_4139 ( .A(core__abc_22172_new_n7195_), .B(reset_n), .Y(core__abc_22172_new_n7196_));
AND2X2 AND2X2_414 ( .A(_abc_19873_new_n1621_), .B(reset_n), .Y(_0word3_reg_31_0__3_));
AND2X2 AND2X2_4140 ( .A(core__abc_22172_new_n7194_), .B(core__abc_22172_new_n7196_), .Y(core__0v2_reg_63_0__11_));
AND2X2 AND2X2_4141 ( .A(core__abc_22172_new_n7183_), .B(core__abc_22172_new_n7160_), .Y(core__abc_22172_new_n7198_));
AND2X2 AND2X2_4142 ( .A(core__abc_22172_new_n7198_), .B(core__abc_22172_new_n7150_), .Y(core__abc_22172_new_n7199_));
AND2X2 AND2X2_4143 ( .A(core__abc_22172_new_n7182_), .B(core__abc_22172_new_n7157_), .Y(core__abc_22172_new_n7201_));
AND2X2 AND2X2_4144 ( .A(core__abc_22172_new_n7198_), .B(core__abc_22172_new_n7146_), .Y(core__abc_22172_new_n7204_));
AND2X2 AND2X2_4145 ( .A(core__abc_22172_new_n7093_), .B(core__abc_22172_new_n7204_), .Y(core__abc_22172_new_n7205_));
AND2X2 AND2X2_4146 ( .A(core__abc_22172_new_n7208_), .B(core__abc_22172_new_n7209_), .Y(core__abc_22172_new_n7210_));
AND2X2 AND2X2_4147 ( .A(core__abc_22172_new_n7211_), .B(core__abc_22172_new_n3269_), .Y(core__abc_22172_new_n7212_));
AND2X2 AND2X2_4148 ( .A(core__abc_22172_new_n7210_), .B(core__abc_22172_new_n3268_), .Y(core__abc_22172_new_n7213_));
AND2X2 AND2X2_4149 ( .A(core__abc_22172_new_n7206_), .B(core__abc_22172_new_n7215_), .Y(core__abc_22172_new_n7216_));
AND2X2 AND2X2_415 ( .A(core_siphash_valid_reg), .B(core_siphash_word_100_), .Y(_abc_19873_new_n1623_));
AND2X2 AND2X2_4150 ( .A(core__abc_22172_new_n7217_), .B(core__abc_22172_new_n7214_), .Y(core__abc_22172_new_n7218_));
AND2X2 AND2X2_4151 ( .A(core__abc_22172_new_n7220_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n7221_));
AND2X2 AND2X2_4152 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n7222_), .Y(core__abc_22172_new_n7223_));
AND2X2 AND2X2_4153 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_12_), .Y(core__abc_22172_new_n7224_));
AND2X2 AND2X2_4154 ( .A(core__abc_22172_new_n7228_), .B(reset_n), .Y(core__abc_22172_new_n7229_));
AND2X2 AND2X2_4155 ( .A(core__abc_22172_new_n7227_), .B(core__abc_22172_new_n7229_), .Y(core__0v2_reg_63_0__12_));
AND2X2 AND2X2_4156 ( .A(core__abc_22172_new_n4001_), .B(core__abc_22172_new_n7233_), .Y(core__abc_22172_new_n7234_));
AND2X2 AND2X2_4157 ( .A(core__abc_22172_new_n4002_), .B(core_v1_reg_32_), .Y(core__abc_22172_new_n7235_));
AND2X2 AND2X2_4158 ( .A(core__abc_22172_new_n7237_), .B(core__abc_22172_new_n7232_), .Y(core__abc_22172_new_n7238_));
AND2X2 AND2X2_4159 ( .A(core__abc_22172_new_n7236_), .B(core__abc_22172_new_n3325_), .Y(core__abc_22172_new_n7239_));
AND2X2 AND2X2_416 ( .A(_abc_19873_new_n1607_), .B(word3_reg_4_), .Y(_abc_19873_new_n1624_));
AND2X2 AND2X2_4160 ( .A(core__abc_22172_new_n7231_), .B(core__abc_22172_new_n7240_), .Y(core__abc_22172_new_n7241_));
AND2X2 AND2X2_4161 ( .A(core__abc_22172_new_n7242_), .B(core__abc_22172_new_n7243_), .Y(core__abc_22172_new_n7244_));
AND2X2 AND2X2_4162 ( .A(core__abc_22172_new_n7245_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n7246_));
AND2X2 AND2X2_4163 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n7247_), .Y(core__abc_22172_new_n7248_));
AND2X2 AND2X2_4164 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_13_), .Y(core__abc_22172_new_n7249_));
AND2X2 AND2X2_4165 ( .A(core__abc_22172_new_n7253_), .B(reset_n), .Y(core__abc_22172_new_n7254_));
AND2X2 AND2X2_4166 ( .A(core__abc_22172_new_n7252_), .B(core__abc_22172_new_n7254_), .Y(core__0v2_reg_63_0__13_));
AND2X2 AND2X2_4167 ( .A(core__abc_22172_new_n7257_), .B(core__abc_22172_new_n7256_), .Y(core__abc_22172_new_n7258_));
AND2X2 AND2X2_4168 ( .A(core__abc_22172_new_n7243_), .B(core__abc_22172_new_n7215_), .Y(core__abc_22172_new_n7260_));
AND2X2 AND2X2_4169 ( .A(core__abc_22172_new_n7262_), .B(core__abc_22172_new_n7259_), .Y(core__abc_22172_new_n7263_));
AND2X2 AND2X2_417 ( .A(_abc_19873_new_n1625_), .B(reset_n), .Y(_0word3_reg_31_0__4_));
AND2X2 AND2X2_4170 ( .A(core__abc_22172_new_n7267_), .B(core__abc_22172_new_n7268_), .Y(core__abc_22172_new_n7269_));
AND2X2 AND2X2_4171 ( .A(core__abc_22172_new_n7269_), .B(core__abc_22172_new_n3358_), .Y(core__abc_22172_new_n7270_));
AND2X2 AND2X2_4172 ( .A(core__abc_22172_new_n7271_), .B(core__abc_22172_new_n3359_), .Y(core__abc_22172_new_n7272_));
AND2X2 AND2X2_4173 ( .A(core__abc_22172_new_n7264_), .B(core__abc_22172_new_n7274_), .Y(core__abc_22172_new_n7275_));
AND2X2 AND2X2_4174 ( .A(core__abc_22172_new_n7263_), .B(core__abc_22172_new_n7273_), .Y(core__abc_22172_new_n7276_));
AND2X2 AND2X2_4175 ( .A(core__abc_22172_new_n7278_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n7279_));
AND2X2 AND2X2_4176 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n7280_), .Y(core__abc_22172_new_n7281_));
AND2X2 AND2X2_4177 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_14_), .Y(core__abc_22172_new_n7282_));
AND2X2 AND2X2_4178 ( .A(core__abc_22172_new_n7286_), .B(reset_n), .Y(core__abc_22172_new_n7287_));
AND2X2 AND2X2_4179 ( .A(core__abc_22172_new_n7285_), .B(core__abc_22172_new_n7287_), .Y(core__0v2_reg_63_0__14_));
AND2X2 AND2X2_418 ( .A(core_siphash_valid_reg), .B(core_siphash_word_101_), .Y(_abc_19873_new_n1627_));
AND2X2 AND2X2_4180 ( .A(core__abc_22172_new_n4134_), .B(core_v1_reg_34_), .Y(core__abc_22172_new_n7292_));
AND2X2 AND2X2_4181 ( .A(core__abc_22172_new_n7293_), .B(core__abc_22172_new_n7291_), .Y(core__abc_22172_new_n7294_));
AND2X2 AND2X2_4182 ( .A(core__abc_22172_new_n7294_), .B(core__abc_22172_new_n3450_), .Y(core__abc_22172_new_n7295_));
AND2X2 AND2X2_4183 ( .A(core__abc_22172_new_n7297_), .B(core__abc_22172_new_n3447_), .Y(core__abc_22172_new_n7298_));
AND2X2 AND2X2_4184 ( .A(core__abc_22172_new_n7290_), .B(core__abc_22172_new_n7299_), .Y(core__abc_22172_new_n7300_));
AND2X2 AND2X2_4185 ( .A(core__abc_22172_new_n7301_), .B(core__abc_22172_new_n7302_), .Y(core__abc_22172_new_n7303_));
AND2X2 AND2X2_4186 ( .A(core__abc_22172_new_n7289_), .B(core__abc_22172_new_n7303_), .Y(core__abc_22172_new_n7304_));
AND2X2 AND2X2_4187 ( .A(core__abc_22172_new_n7306_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n7307_));
AND2X2 AND2X2_4188 ( .A(core__abc_22172_new_n3214_), .B(core_key_15_), .Y(core__abc_22172_new_n7308_));
AND2X2 AND2X2_4189 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_15_), .Y(core__abc_22172_new_n7309_));
AND2X2 AND2X2_419 ( .A(_abc_19873_new_n1607_), .B(word3_reg_5_), .Y(_abc_19873_new_n1628_));
AND2X2 AND2X2_4190 ( .A(core__abc_22172_new_n7313_), .B(reset_n), .Y(core__abc_22172_new_n7314_));
AND2X2 AND2X2_4191 ( .A(core__abc_22172_new_n7312_), .B(core__abc_22172_new_n7314_), .Y(core__0v2_reg_63_0__15_));
AND2X2 AND2X2_4192 ( .A(core__abc_22172_new_n7302_), .B(core__abc_22172_new_n7272_), .Y(core__abc_22172_new_n7321_));
AND2X2 AND2X2_4193 ( .A(core__abc_22172_new_n7320_), .B(core__abc_22172_new_n7323_), .Y(core__abc_22172_new_n7324_));
AND2X2 AND2X2_4194 ( .A(core__abc_22172_new_n7319_), .B(core__abc_22172_new_n7324_), .Y(core__abc_22172_new_n7325_));
AND2X2 AND2X2_4195 ( .A(core__abc_22172_new_n7328_), .B(core__abc_22172_new_n7325_), .Y(core__abc_22172_new_n7329_));
AND2X2 AND2X2_4196 ( .A(core__abc_22172_new_n7303_), .B(core__abc_22172_new_n7274_), .Y(core__abc_22172_new_n7330_));
AND2X2 AND2X2_4197 ( .A(core__abc_22172_new_n7330_), .B(core__abc_22172_new_n7260_), .Y(core__abc_22172_new_n7331_));
AND2X2 AND2X2_4198 ( .A(core__abc_22172_new_n7331_), .B(core__abc_22172_new_n7204_), .Y(core__abc_22172_new_n7332_));
AND2X2 AND2X2_4199 ( .A(core__abc_22172_new_n7332_), .B(core__abc_22172_new_n7078_), .Y(core__abc_22172_new_n7333_));
AND2X2 AND2X2_42 ( .A(_abc_19873_new_n925_), .B(word2_reg_0_), .Y(_abc_19873_new_n926_));
AND2X2 AND2X2_420 ( .A(_abc_19873_new_n1629_), .B(reset_n), .Y(_0word3_reg_31_0__5_));
AND2X2 AND2X2_4200 ( .A(core__abc_22172_new_n7333_), .B(core__abc_22172_new_n6851_), .Y(core__abc_22172_new_n7334_));
AND2X2 AND2X2_4201 ( .A(core__abc_22172_new_n7335_), .B(core__abc_22172_new_n7329_), .Y(core__abc_22172_new_n7336_));
AND2X2 AND2X2_4202 ( .A(core__abc_22172_new_n7339_), .B(core__abc_22172_new_n7340_), .Y(core__abc_22172_new_n7341_));
AND2X2 AND2X2_4203 ( .A(core__abc_22172_new_n3516_), .B(core__abc_22172_new_n7342_), .Y(core__abc_22172_new_n7343_));
AND2X2 AND2X2_4204 ( .A(core__abc_22172_new_n3515_), .B(core__abc_22172_new_n7341_), .Y(core__abc_22172_new_n7344_));
AND2X2 AND2X2_4205 ( .A(core__abc_22172_new_n7337_), .B(core__abc_22172_new_n7346_), .Y(core__abc_22172_new_n7347_));
AND2X2 AND2X2_4206 ( .A(core__abc_22172_new_n7336_), .B(core__abc_22172_new_n7345_), .Y(core__abc_22172_new_n7348_));
AND2X2 AND2X2_4207 ( .A(core__abc_22172_new_n7350_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n7351_));
AND2X2 AND2X2_4208 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n7352_), .Y(core__abc_22172_new_n7353_));
AND2X2 AND2X2_4209 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_16_), .Y(core__abc_22172_new_n7354_));
AND2X2 AND2X2_421 ( .A(core_siphash_valid_reg), .B(core_siphash_word_102_), .Y(_abc_19873_new_n1631_));
AND2X2 AND2X2_4210 ( .A(core__abc_22172_new_n7358_), .B(reset_n), .Y(core__abc_22172_new_n7359_));
AND2X2 AND2X2_4211 ( .A(core__abc_22172_new_n7357_), .B(core__abc_22172_new_n7359_), .Y(core__0v2_reg_63_0__16_));
AND2X2 AND2X2_4212 ( .A(core__abc_22172_new_n7362_), .B(core__abc_22172_new_n7361_), .Y(core__abc_22172_new_n7363_));
AND2X2 AND2X2_4213 ( .A(core__abc_22172_new_n7365_), .B(core__abc_22172_new_n7364_), .Y(core__abc_22172_new_n7366_));
AND2X2 AND2X2_4214 ( .A(core__abc_22172_new_n4282_), .B(core_v1_reg_36_), .Y(core__abc_22172_new_n7367_));
AND2X2 AND2X2_4215 ( .A(core__abc_22172_new_n3584_), .B(core__abc_22172_new_n7369_), .Y(core__abc_22172_new_n7370_));
AND2X2 AND2X2_4216 ( .A(core__abc_22172_new_n3582_), .B(core__abc_22172_new_n7368_), .Y(core__abc_22172_new_n7372_));
AND2X2 AND2X2_4217 ( .A(core__abc_22172_new_n7371_), .B(core__abc_22172_new_n7373_), .Y(core__abc_22172_new_n7374_));
AND2X2 AND2X2_4218 ( .A(core__abc_22172_new_n7378_), .B(core__abc_22172_new_n7375_), .Y(core__abc_22172_new_n7379_));
AND2X2 AND2X2_4219 ( .A(core__abc_22172_new_n7380_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n7381_));
AND2X2 AND2X2_422 ( .A(_abc_19873_new_n1607_), .B(word3_reg_6_), .Y(_abc_19873_new_n1632_));
AND2X2 AND2X2_4220 ( .A(core__abc_22172_new_n3214_), .B(core_key_17_), .Y(core__abc_22172_new_n7382_));
AND2X2 AND2X2_4221 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_17_), .Y(core__abc_22172_new_n7383_));
AND2X2 AND2X2_4222 ( .A(core__abc_22172_new_n7387_), .B(reset_n), .Y(core__abc_22172_new_n7388_));
AND2X2 AND2X2_4223 ( .A(core__abc_22172_new_n7386_), .B(core__abc_22172_new_n7388_), .Y(core__0v2_reg_63_0__17_));
AND2X2 AND2X2_4224 ( .A(core__abc_22172_new_n7392_), .B(core__abc_22172_new_n7391_), .Y(core__abc_22172_new_n7393_));
AND2X2 AND2X2_4225 ( .A(core__abc_22172_new_n3639_), .B(core__abc_22172_new_n7394_), .Y(core__abc_22172_new_n7395_));
AND2X2 AND2X2_4226 ( .A(core__abc_22172_new_n3638_), .B(core__abc_22172_new_n7393_), .Y(core__abc_22172_new_n7396_));
AND2X2 AND2X2_4227 ( .A(core__abc_22172_new_n7371_), .B(core__abc_22172_new_n7361_), .Y(core__abc_22172_new_n7399_));
AND2X2 AND2X2_4228 ( .A(core__abc_22172_new_n7362_), .B(core__abc_22172_new_n7399_), .Y(core__abc_22172_new_n7400_));
AND2X2 AND2X2_4229 ( .A(core__abc_22172_new_n7402_), .B(core__abc_22172_new_n7398_), .Y(core__abc_22172_new_n7403_));
AND2X2 AND2X2_423 ( .A(_abc_19873_new_n1633_), .B(reset_n), .Y(_0word3_reg_31_0__6_));
AND2X2 AND2X2_4230 ( .A(core__abc_22172_new_n7401_), .B(core__abc_22172_new_n7397_), .Y(core__abc_22172_new_n7404_));
AND2X2 AND2X2_4231 ( .A(core__abc_22172_new_n7406_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n7407_));
AND2X2 AND2X2_4232 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n7408_), .Y(core__abc_22172_new_n7409_));
AND2X2 AND2X2_4233 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_18_), .Y(core__abc_22172_new_n7410_));
AND2X2 AND2X2_4234 ( .A(core__abc_22172_new_n7414_), .B(reset_n), .Y(core__abc_22172_new_n7415_));
AND2X2 AND2X2_4235 ( .A(core__abc_22172_new_n7413_), .B(core__abc_22172_new_n7415_), .Y(core__0v2_reg_63_0__18_));
AND2X2 AND2X2_4236 ( .A(core__abc_22172_new_n7419_), .B(core__abc_22172_new_n7418_), .Y(core__abc_22172_new_n7420_));
AND2X2 AND2X2_4237 ( .A(core__abc_22172_new_n4403_), .B(core_v1_reg_38_), .Y(core__abc_22172_new_n7421_));
AND2X2 AND2X2_4238 ( .A(core__abc_22172_new_n3711_), .B(core__abc_22172_new_n7423_), .Y(core__abc_22172_new_n7424_));
AND2X2 AND2X2_4239 ( .A(core__abc_22172_new_n3712_), .B(core__abc_22172_new_n7422_), .Y(core__abc_22172_new_n7426_));
AND2X2 AND2X2_424 ( .A(core_siphash_valid_reg), .B(core_siphash_word_103_), .Y(_abc_19873_new_n1635_));
AND2X2 AND2X2_4240 ( .A(core__abc_22172_new_n7427_), .B(core__abc_22172_new_n7425_), .Y(core__abc_22172_new_n7428_));
AND2X2 AND2X2_4241 ( .A(core__abc_22172_new_n7432_), .B(core__abc_22172_new_n7429_), .Y(core__abc_22172_new_n7433_));
AND2X2 AND2X2_4242 ( .A(core__abc_22172_new_n7433_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n7434_));
AND2X2 AND2X2_4243 ( .A(core__abc_22172_new_n3214_), .B(core_key_19_), .Y(core__abc_22172_new_n7435_));
AND2X2 AND2X2_4244 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_19_), .Y(core__abc_22172_new_n7436_));
AND2X2 AND2X2_4245 ( .A(core__abc_22172_new_n7440_), .B(reset_n), .Y(core__abc_22172_new_n7441_));
AND2X2 AND2X2_4246 ( .A(core__abc_22172_new_n7439_), .B(core__abc_22172_new_n7441_), .Y(core__0v2_reg_63_0__19_));
AND2X2 AND2X2_4247 ( .A(core__abc_22172_new_n7427_), .B(core__abc_22172_new_n7443_), .Y(core__abc_22172_new_n7444_));
AND2X2 AND2X2_4248 ( .A(core__abc_22172_new_n7428_), .B(core__abc_22172_new_n7398_), .Y(core__abc_22172_new_n7447_));
AND2X2 AND2X2_4249 ( .A(core__abc_22172_new_n7449_), .B(core__abc_22172_new_n7445_), .Y(core__abc_22172_new_n7450_));
AND2X2 AND2X2_425 ( .A(_abc_19873_new_n1607_), .B(word3_reg_7_), .Y(_abc_19873_new_n1636_));
AND2X2 AND2X2_4250 ( .A(core__abc_22172_new_n7374_), .B(core__abc_22172_new_n7346_), .Y(core__abc_22172_new_n7451_));
AND2X2 AND2X2_4251 ( .A(core__abc_22172_new_n7447_), .B(core__abc_22172_new_n7451_), .Y(core__abc_22172_new_n7452_));
AND2X2 AND2X2_4252 ( .A(core__abc_22172_new_n7454_), .B(core__abc_22172_new_n7450_), .Y(core__abc_22172_new_n7455_));
AND2X2 AND2X2_4253 ( .A(core__abc_22172_new_n7457_), .B(core__abc_22172_new_n7458_), .Y(core__abc_22172_new_n7459_));
AND2X2 AND2X2_4254 ( .A(core__abc_22172_new_n3782_), .B(core__abc_22172_new_n7460_), .Y(core__abc_22172_new_n7461_));
AND2X2 AND2X2_4255 ( .A(core__abc_22172_new_n3781_), .B(core__abc_22172_new_n7459_), .Y(core__abc_22172_new_n7462_));
AND2X2 AND2X2_4256 ( .A(core__abc_22172_new_n7455_), .B(core__abc_22172_new_n7463_), .Y(core__abc_22172_new_n7466_));
AND2X2 AND2X2_4257 ( .A(core__abc_22172_new_n7468_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n7469_));
AND2X2 AND2X2_4258 ( .A(core__abc_22172_new_n3214_), .B(core_key_20_), .Y(core__abc_22172_new_n7470_));
AND2X2 AND2X2_4259 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_20_), .Y(core__abc_22172_new_n7471_));
AND2X2 AND2X2_426 ( .A(_abc_19873_new_n1637_), .B(reset_n), .Y(_0word3_reg_31_0__7_));
AND2X2 AND2X2_4260 ( .A(core__abc_22172_new_n7475_), .B(reset_n), .Y(core__abc_22172_new_n7476_));
AND2X2 AND2X2_4261 ( .A(core__abc_22172_new_n7474_), .B(core__abc_22172_new_n7476_), .Y(core__0v2_reg_63_0__20_));
AND2X2 AND2X2_4262 ( .A(core__abc_22172_new_n7464_), .B(core__abc_22172_new_n7478_), .Y(core__abc_22172_new_n7479_));
AND2X2 AND2X2_4263 ( .A(core__abc_22172_new_n4526_), .B(core__abc_22172_new_n7482_), .Y(core__abc_22172_new_n7483_));
AND2X2 AND2X2_4264 ( .A(core__abc_22172_new_n4527_), .B(core_v1_reg_40_), .Y(core__abc_22172_new_n7484_));
AND2X2 AND2X2_4265 ( .A(core__abc_22172_new_n7481_), .B(core__abc_22172_new_n7486_), .Y(core__abc_22172_new_n7487_));
AND2X2 AND2X2_4266 ( .A(core__abc_22172_new_n3845_), .B(core__abc_22172_new_n7485_), .Y(core__abc_22172_new_n7489_));
AND2X2 AND2X2_4267 ( .A(core__abc_22172_new_n7488_), .B(core__abc_22172_new_n7490_), .Y(core__abc_22172_new_n7491_));
AND2X2 AND2X2_4268 ( .A(core__abc_22172_new_n7492_), .B(core__abc_22172_new_n7494_), .Y(core__abc_22172_new_n7495_));
AND2X2 AND2X2_4269 ( .A(core__abc_22172_new_n7495_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n7496_));
AND2X2 AND2X2_427 ( .A(core_siphash_valid_reg), .B(core_siphash_word_104_), .Y(_abc_19873_new_n1639_));
AND2X2 AND2X2_4270 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n7497_), .Y(core__abc_22172_new_n7498_));
AND2X2 AND2X2_4271 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_21_), .Y(core__abc_22172_new_n7499_));
AND2X2 AND2X2_4272 ( .A(core__abc_22172_new_n7503_), .B(reset_n), .Y(core__abc_22172_new_n7504_));
AND2X2 AND2X2_4273 ( .A(core__abc_22172_new_n7502_), .B(core__abc_22172_new_n7504_), .Y(core__0v2_reg_63_0__21_));
AND2X2 AND2X2_4274 ( .A(core__abc_22172_new_n7508_), .B(core__abc_22172_new_n7509_), .Y(core__abc_22172_new_n7510_));
AND2X2 AND2X2_4275 ( .A(core__abc_22172_new_n3905_), .B(core__abc_22172_new_n7511_), .Y(core__abc_22172_new_n7512_));
AND2X2 AND2X2_4276 ( .A(core__abc_22172_new_n3904_), .B(core__abc_22172_new_n7510_), .Y(core__abc_22172_new_n7513_));
AND2X2 AND2X2_4277 ( .A(core__abc_22172_new_n7488_), .B(core__abc_22172_new_n7478_), .Y(core__abc_22172_new_n7517_));
AND2X2 AND2X2_4278 ( .A(core__abc_22172_new_n7516_), .B(core__abc_22172_new_n7518_), .Y(core__abc_22172_new_n7519_));
AND2X2 AND2X2_4279 ( .A(core__abc_22172_new_n7519_), .B(core__abc_22172_new_n7514_), .Y(core__abc_22172_new_n7522_));
AND2X2 AND2X2_428 ( .A(_abc_19873_new_n1607_), .B(word3_reg_8_), .Y(_abc_19873_new_n1640_));
AND2X2 AND2X2_4280 ( .A(core__abc_22172_new_n7524_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n7525_));
AND2X2 AND2X2_4281 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n7526_), .Y(core__abc_22172_new_n7527_));
AND2X2 AND2X2_4282 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_22_), .Y(core__abc_22172_new_n7528_));
AND2X2 AND2X2_4283 ( .A(core__abc_22172_new_n7532_), .B(reset_n), .Y(core__abc_22172_new_n7533_));
AND2X2 AND2X2_4284 ( .A(core__abc_22172_new_n7531_), .B(core__abc_22172_new_n7533_), .Y(core__0v2_reg_63_0__22_));
AND2X2 AND2X2_4285 ( .A(core__abc_22172_new_n7520_), .B(core__abc_22172_new_n7535_), .Y(core__abc_22172_new_n7536_));
AND2X2 AND2X2_4286 ( .A(core__abc_22172_new_n4638_), .B(core__abc_22172_new_n7538_), .Y(core__abc_22172_new_n7539_));
AND2X2 AND2X2_4287 ( .A(core__abc_22172_new_n4626_), .B(core_v1_reg_42_), .Y(core__abc_22172_new_n7540_));
AND2X2 AND2X2_4288 ( .A(core__abc_22172_new_n7537_), .B(core__abc_22172_new_n7542_), .Y(core__abc_22172_new_n7543_));
AND2X2 AND2X2_4289 ( .A(core__abc_22172_new_n3972_), .B(core__abc_22172_new_n7541_), .Y(core__abc_22172_new_n7545_));
AND2X2 AND2X2_429 ( .A(_abc_19873_new_n1641_), .B(reset_n), .Y(_0word3_reg_31_0__8_));
AND2X2 AND2X2_4290 ( .A(core__abc_22172_new_n7544_), .B(core__abc_22172_new_n7546_), .Y(core__abc_22172_new_n7547_));
AND2X2 AND2X2_4291 ( .A(core__abc_22172_new_n7536_), .B(core__abc_22172_new_n7548_), .Y(core__abc_22172_new_n7549_));
AND2X2 AND2X2_4292 ( .A(core__abc_22172_new_n7550_), .B(core__abc_22172_new_n7547_), .Y(core__abc_22172_new_n7551_));
AND2X2 AND2X2_4293 ( .A(core__abc_22172_new_n7553_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n7554_));
AND2X2 AND2X2_4294 ( .A(core__abc_22172_new_n3214_), .B(core_key_23_), .Y(core__abc_22172_new_n7555_));
AND2X2 AND2X2_4295 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_23_), .Y(core__abc_22172_new_n7556_));
AND2X2 AND2X2_4296 ( .A(core__abc_22172_new_n7560_), .B(reset_n), .Y(core__abc_22172_new_n7561_));
AND2X2 AND2X2_4297 ( .A(core__abc_22172_new_n7559_), .B(core__abc_22172_new_n7561_), .Y(core__0v2_reg_63_0__23_));
AND2X2 AND2X2_4298 ( .A(core__abc_22172_new_n7547_), .B(core__abc_22172_new_n7565_), .Y(core__abc_22172_new_n7566_));
AND2X2 AND2X2_4299 ( .A(core__abc_22172_new_n7566_), .B(core__abc_22172_new_n7564_), .Y(core__abc_22172_new_n7567_));
AND2X2 AND2X2_43 ( .A(_abc_19873_new_n875_), .B(_abc_19873_new_n904_), .Y(_abc_19873_new_n928_));
AND2X2 AND2X2_430 ( .A(core_siphash_valid_reg), .B(core_siphash_word_105_), .Y(_abc_19873_new_n1643_));
AND2X2 AND2X2_4300 ( .A(core__abc_22172_new_n7563_), .B(core__abc_22172_new_n7567_), .Y(core__abc_22172_new_n7568_));
AND2X2 AND2X2_4301 ( .A(core__abc_22172_new_n7566_), .B(core__abc_22172_new_n7569_), .Y(core__abc_22172_new_n7570_));
AND2X2 AND2X2_4302 ( .A(core__abc_22172_new_n7546_), .B(core__abc_22172_new_n7512_), .Y(core__abc_22172_new_n7571_));
AND2X2 AND2X2_4303 ( .A(core__abc_22172_new_n7567_), .B(core__abc_22172_new_n7452_), .Y(core__abc_22172_new_n7575_));
AND2X2 AND2X2_4304 ( .A(core__abc_22172_new_n7337_), .B(core__abc_22172_new_n7575_), .Y(core__abc_22172_new_n7576_));
AND2X2 AND2X2_4305 ( .A(core__abc_22172_new_n7579_), .B(core__abc_22172_new_n7580_), .Y(core__abc_22172_new_n7581_));
AND2X2 AND2X2_4306 ( .A(core__abc_22172_new_n4040_), .B(core__abc_22172_new_n7582_), .Y(core__abc_22172_new_n7583_));
AND2X2 AND2X2_4307 ( .A(core__abc_22172_new_n4039_), .B(core__abc_22172_new_n7581_), .Y(core__abc_22172_new_n7584_));
AND2X2 AND2X2_4308 ( .A(core__abc_22172_new_n7577_), .B(core__abc_22172_new_n7586_), .Y(core__abc_22172_new_n7587_));
AND2X2 AND2X2_4309 ( .A(core__abc_22172_new_n7588_), .B(core__abc_22172_new_n7585_), .Y(core__abc_22172_new_n7589_));
AND2X2 AND2X2_431 ( .A(_abc_19873_new_n1607_), .B(word3_reg_9_), .Y(_abc_19873_new_n1644_));
AND2X2 AND2X2_4310 ( .A(core__abc_22172_new_n7591_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n7592_));
AND2X2 AND2X2_4311 ( .A(core__abc_22172_new_n3214_), .B(core_key_24_), .Y(core__abc_22172_new_n7593_));
AND2X2 AND2X2_4312 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_24_), .Y(core__abc_22172_new_n7594_));
AND2X2 AND2X2_4313 ( .A(core__abc_22172_new_n7598_), .B(reset_n), .Y(core__abc_22172_new_n7599_));
AND2X2 AND2X2_4314 ( .A(core__abc_22172_new_n7597_), .B(core__abc_22172_new_n7599_), .Y(core__0v2_reg_63_0__24_));
AND2X2 AND2X2_4315 ( .A(core__abc_22172_new_n4749_), .B(core_v1_reg_44_), .Y(core__abc_22172_new_n7602_));
AND2X2 AND2X2_4316 ( .A(core__abc_22172_new_n7603_), .B(core__abc_22172_new_n7604_), .Y(core__abc_22172_new_n7605_));
AND2X2 AND2X2_4317 ( .A(core__abc_22172_new_n4104_), .B(core__abc_22172_new_n7605_), .Y(core__abc_22172_new_n7606_));
AND2X2 AND2X2_4318 ( .A(core__abc_22172_new_n4103_), .B(core__abc_22172_new_n7608_), .Y(core__abc_22172_new_n7609_));
AND2X2 AND2X2_4319 ( .A(core__abc_22172_new_n7607_), .B(core__abc_22172_new_n7610_), .Y(core__abc_22172_new_n7611_));
AND2X2 AND2X2_432 ( .A(_abc_19873_new_n1645_), .B(reset_n), .Y(_0word3_reg_31_0__9_));
AND2X2 AND2X2_4320 ( .A(core__abc_22172_new_n7615_), .B(core__abc_22172_new_n7612_), .Y(core__abc_22172_new_n7616_));
AND2X2 AND2X2_4321 ( .A(core__abc_22172_new_n7616_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n7617_));
AND2X2 AND2X2_4322 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n7618_), .Y(core__abc_22172_new_n7619_));
AND2X2 AND2X2_4323 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_25_), .Y(core__abc_22172_new_n7620_));
AND2X2 AND2X2_4324 ( .A(core__abc_22172_new_n7624_), .B(reset_n), .Y(core__abc_22172_new_n7625_));
AND2X2 AND2X2_4325 ( .A(core__abc_22172_new_n7623_), .B(core__abc_22172_new_n7625_), .Y(core__0v2_reg_63_0__25_));
AND2X2 AND2X2_4326 ( .A(core__abc_22172_new_n7628_), .B(core__abc_22172_new_n7629_), .Y(core__abc_22172_new_n7630_));
AND2X2 AND2X2_4327 ( .A(core__abc_22172_new_n4165_), .B(core__abc_22172_new_n7631_), .Y(core__abc_22172_new_n7632_));
AND2X2 AND2X2_4328 ( .A(core__abc_22172_new_n4164_), .B(core__abc_22172_new_n7630_), .Y(core__abc_22172_new_n7633_));
AND2X2 AND2X2_4329 ( .A(core__abc_22172_new_n7611_), .B(core__abc_22172_new_n7586_), .Y(core__abc_22172_new_n7636_));
AND2X2 AND2X2_433 ( .A(core_siphash_valid_reg), .B(core_siphash_word_106_), .Y(_abc_19873_new_n1647_));
AND2X2 AND2X2_4330 ( .A(core__abc_22172_new_n7577_), .B(core__abc_22172_new_n7636_), .Y(core__abc_22172_new_n7637_));
AND2X2 AND2X2_4331 ( .A(core__abc_22172_new_n7607_), .B(core__abc_22172_new_n7638_), .Y(core__abc_22172_new_n7639_));
AND2X2 AND2X2_4332 ( .A(core__abc_22172_new_n7642_), .B(core__abc_22172_new_n7635_), .Y(core__abc_22172_new_n7643_));
AND2X2 AND2X2_4333 ( .A(core__abc_22172_new_n7644_), .B(core__abc_22172_new_n7645_), .Y(core__abc_22172_new_n7646_));
AND2X2 AND2X2_4334 ( .A(core__abc_22172_new_n7646_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n7647_));
AND2X2 AND2X2_4335 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n7648_), .Y(core__abc_22172_new_n7649_));
AND2X2 AND2X2_4336 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_26_), .Y(core__abc_22172_new_n7650_));
AND2X2 AND2X2_4337 ( .A(core__abc_22172_new_n7654_), .B(reset_n), .Y(core__abc_22172_new_n7655_));
AND2X2 AND2X2_4338 ( .A(core__abc_22172_new_n7653_), .B(core__abc_22172_new_n7655_), .Y(core__0v2_reg_63_0__26_));
AND2X2 AND2X2_4339 ( .A(core__abc_22172_new_n7644_), .B(core__abc_22172_new_n7657_), .Y(core__abc_22172_new_n7658_));
AND2X2 AND2X2_434 ( .A(_abc_19873_new_n1607_), .B(word3_reg_10_), .Y(_abc_19873_new_n1648_));
AND2X2 AND2X2_4340 ( .A(core__abc_22172_new_n4837_), .B(core__abc_22172_new_n7660_), .Y(core__abc_22172_new_n7661_));
AND2X2 AND2X2_4341 ( .A(core__abc_22172_new_n4848_), .B(core_v1_reg_46_), .Y(core__abc_22172_new_n7662_));
AND2X2 AND2X2_4342 ( .A(core__abc_22172_new_n4249_), .B(core__abc_22172_new_n7664_), .Y(core__abc_22172_new_n7665_));
AND2X2 AND2X2_4343 ( .A(core__abc_22172_new_n4245_), .B(core__abc_22172_new_n7663_), .Y(core__abc_22172_new_n7666_));
AND2X2 AND2X2_4344 ( .A(core__abc_22172_new_n7669_), .B(core__abc_22172_new_n7670_), .Y(core__abc_22172_new_n7671_));
AND2X2 AND2X2_4345 ( .A(core__abc_22172_new_n7671_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n7672_));
AND2X2 AND2X2_4346 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n7673_), .Y(core__abc_22172_new_n7674_));
AND2X2 AND2X2_4347 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_27_), .Y(core__abc_22172_new_n7675_));
AND2X2 AND2X2_4348 ( .A(core__abc_22172_new_n7679_), .B(reset_n), .Y(core__abc_22172_new_n7680_));
AND2X2 AND2X2_4349 ( .A(core__abc_22172_new_n7678_), .B(core__abc_22172_new_n7680_), .Y(core__0v2_reg_63_0__27_));
AND2X2 AND2X2_435 ( .A(_abc_19873_new_n1649_), .B(reset_n), .Y(_0word3_reg_31_0__10_));
AND2X2 AND2X2_4350 ( .A(core__abc_22172_new_n7668_), .B(core__abc_22172_new_n7635_), .Y(core__abc_22172_new_n7682_));
AND2X2 AND2X2_4351 ( .A(core__abc_22172_new_n7682_), .B(core__abc_22172_new_n7636_), .Y(core__abc_22172_new_n7683_));
AND2X2 AND2X2_4352 ( .A(core__abc_22172_new_n7577_), .B(core__abc_22172_new_n7683_), .Y(core__abc_22172_new_n7684_));
AND2X2 AND2X2_4353 ( .A(core__abc_22172_new_n7682_), .B(core__abc_22172_new_n7641_), .Y(core__abc_22172_new_n7685_));
AND2X2 AND2X2_4354 ( .A(core__abc_22172_new_n7668_), .B(core__abc_22172_new_n7632_), .Y(core__abc_22172_new_n7686_));
AND2X2 AND2X2_4355 ( .A(core__abc_22172_new_n7692_), .B(core__abc_22172_new_n7693_), .Y(core__abc_22172_new_n7694_));
AND2X2 AND2X2_4356 ( .A(core__abc_22172_new_n4316_), .B(core__abc_22172_new_n7695_), .Y(core__abc_22172_new_n7696_));
AND2X2 AND2X2_4357 ( .A(core__abc_22172_new_n4315_), .B(core__abc_22172_new_n7694_), .Y(core__abc_22172_new_n7697_));
AND2X2 AND2X2_4358 ( .A(core__abc_22172_new_n7690_), .B(core__abc_22172_new_n7698_), .Y(core__abc_22172_new_n7699_));
AND2X2 AND2X2_4359 ( .A(core__abc_22172_new_n7689_), .B(core__abc_22172_new_n7700_), .Y(core__abc_22172_new_n7701_));
AND2X2 AND2X2_436 ( .A(core_siphash_valid_reg), .B(core_siphash_word_107_), .Y(_abc_19873_new_n1651_));
AND2X2 AND2X2_4360 ( .A(core__abc_22172_new_n7703_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n7704_));
AND2X2 AND2X2_4361 ( .A(core__abc_22172_new_n3214_), .B(core_key_28_), .Y(core__abc_22172_new_n7705_));
AND2X2 AND2X2_4362 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_28_), .Y(core__abc_22172_new_n7706_));
AND2X2 AND2X2_4363 ( .A(core__abc_22172_new_n7710_), .B(reset_n), .Y(core__abc_22172_new_n7711_));
AND2X2 AND2X2_4364 ( .A(core__abc_22172_new_n7709_), .B(core__abc_22172_new_n7711_), .Y(core__0v2_reg_63_0__28_));
AND2X2 AND2X2_4365 ( .A(core__abc_22172_new_n4958_), .B(core__abc_22172_new_n7713_), .Y(core__abc_22172_new_n7714_));
AND2X2 AND2X2_4366 ( .A(core__abc_22172_new_n4946_), .B(core_v1_reg_48_), .Y(core__abc_22172_new_n7715_));
AND2X2 AND2X2_4367 ( .A(core__abc_22172_new_n4372_), .B(core__abc_22172_new_n7716_), .Y(core__abc_22172_new_n7717_));
AND2X2 AND2X2_4368 ( .A(core__abc_22172_new_n4371_), .B(core__abc_22172_new_n7718_), .Y(core__abc_22172_new_n7719_));
AND2X2 AND2X2_4369 ( .A(core__abc_22172_new_n7722_), .B(core__abc_22172_new_n7720_), .Y(core__abc_22172_new_n7723_));
AND2X2 AND2X2_437 ( .A(_abc_19873_new_n1607_), .B(word3_reg_11_), .Y(_abc_19873_new_n1652_));
AND2X2 AND2X2_4370 ( .A(core__abc_22172_new_n7721_), .B(core__abc_22172_new_n7724_), .Y(core__abc_22172_new_n7725_));
AND2X2 AND2X2_4371 ( .A(core__abc_22172_new_n7727_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n7728_));
AND2X2 AND2X2_4372 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n7729_), .Y(core__abc_22172_new_n7730_));
AND2X2 AND2X2_4373 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_29_), .Y(core__abc_22172_new_n7731_));
AND2X2 AND2X2_4374 ( .A(core__abc_22172_new_n7735_), .B(reset_n), .Y(core__abc_22172_new_n7736_));
AND2X2 AND2X2_4375 ( .A(core__abc_22172_new_n7734_), .B(core__abc_22172_new_n7736_), .Y(core__0v2_reg_63_0__29_));
AND2X2 AND2X2_4376 ( .A(core__abc_22172_new_n7724_), .B(core__abc_22172_new_n7700_), .Y(core__abc_22172_new_n7738_));
AND2X2 AND2X2_4377 ( .A(core__abc_22172_new_n7689_), .B(core__abc_22172_new_n7738_), .Y(core__abc_22172_new_n7739_));
AND2X2 AND2X2_4378 ( .A(core__abc_22172_new_n7724_), .B(core__abc_22172_new_n7696_), .Y(core__abc_22172_new_n7740_));
AND2X2 AND2X2_4379 ( .A(core__abc_22172_new_n7745_), .B(core__abc_22172_new_n7746_), .Y(core__abc_22172_new_n7747_));
AND2X2 AND2X2_438 ( .A(_abc_19873_new_n1653_), .B(reset_n), .Y(_0word3_reg_31_0__11_));
AND2X2 AND2X2_4380 ( .A(core__abc_22172_new_n4428_), .B(core__abc_22172_new_n7748_), .Y(core__abc_22172_new_n7749_));
AND2X2 AND2X2_4381 ( .A(core__abc_22172_new_n4429_), .B(core__abc_22172_new_n7747_), .Y(core__abc_22172_new_n7750_));
AND2X2 AND2X2_4382 ( .A(core__abc_22172_new_n7743_), .B(core__abc_22172_new_n7751_), .Y(core__abc_22172_new_n7752_));
AND2X2 AND2X2_4383 ( .A(core__abc_22172_new_n7742_), .B(core__abc_22172_new_n7753_), .Y(core__abc_22172_new_n7754_));
AND2X2 AND2X2_4384 ( .A(core__abc_22172_new_n7756_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n7757_));
AND2X2 AND2X2_4385 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n7758_), .Y(core__abc_22172_new_n7759_));
AND2X2 AND2X2_4386 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_30_), .Y(core__abc_22172_new_n7760_));
AND2X2 AND2X2_4387 ( .A(core__abc_22172_new_n7764_), .B(reset_n), .Y(core__abc_22172_new_n7765_));
AND2X2 AND2X2_4388 ( .A(core__abc_22172_new_n7763_), .B(core__abc_22172_new_n7765_), .Y(core__0v2_reg_63_0__30_));
AND2X2 AND2X2_4389 ( .A(core__abc_22172_new_n5059_), .B(core__abc_22172_new_n7768_), .Y(core__abc_22172_new_n7769_));
AND2X2 AND2X2_439 ( .A(core_siphash_valid_reg), .B(core_siphash_word_108_), .Y(_abc_19873_new_n1655_));
AND2X2 AND2X2_4390 ( .A(core__abc_22172_new_n5045_), .B(core_v1_reg_50_), .Y(core__abc_22172_new_n7770_));
AND2X2 AND2X2_4391 ( .A(core__abc_22172_new_n7774_), .B(core__abc_22172_new_n7773_), .Y(core__abc_22172_new_n7775_));
AND2X2 AND2X2_4392 ( .A(core__abc_22172_new_n7779_), .B(core__abc_22172_new_n7776_), .Y(core__abc_22172_new_n7780_));
AND2X2 AND2X2_4393 ( .A(core__abc_22172_new_n7780_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n7781_));
AND2X2 AND2X2_4394 ( .A(core__abc_22172_new_n3214_), .B(core_key_31_), .Y(core__abc_22172_new_n7782_));
AND2X2 AND2X2_4395 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_31_), .Y(core__abc_22172_new_n7783_));
AND2X2 AND2X2_4396 ( .A(core__abc_22172_new_n7787_), .B(reset_n), .Y(core__abc_22172_new_n7788_));
AND2X2 AND2X2_4397 ( .A(core__abc_22172_new_n7786_), .B(core__abc_22172_new_n7788_), .Y(core__0v2_reg_63_0__31_));
AND2X2 AND2X2_4398 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n7790_), .Y(core__abc_22172_new_n7791_));
AND2X2 AND2X2_4399 ( .A(core__abc_22172_new_n6806_), .B(core__abc_22172_new_n1265_), .Y(core__abc_22172_new_n7792_));
AND2X2 AND2X2_44 ( .A(_abc_19873_new_n928_), .B(core_key_32_), .Y(_abc_19873_new_n929_));
AND2X2 AND2X2_440 ( .A(_abc_19873_new_n1607_), .B(word3_reg_12_), .Y(_abc_19873_new_n1656_));
AND2X2 AND2X2_4400 ( .A(core__abc_22172_new_n3205_), .B(core__abc_22172_new_n7794_), .Y(core__abc_22172_new_n7795_));
AND2X2 AND2X2_4401 ( .A(core__abc_22172_new_n7114_), .B(core__abc_22172_new_n7796_), .Y(core__abc_22172_new_n7797_));
AND2X2 AND2X2_4402 ( .A(core__abc_22172_new_n7798_), .B(core_v2_reg_32_), .Y(core__abc_22172_new_n7799_));
AND2X2 AND2X2_4403 ( .A(core__abc_22172_new_n7800_), .B(reset_n), .Y(core__0v2_reg_63_0__32_));
AND2X2 AND2X2_4404 ( .A(core__abc_22172_new_n7798_), .B(core_v2_reg_33_), .Y(core__abc_22172_new_n7802_));
AND2X2 AND2X2_4405 ( .A(core__abc_22172_new_n3214_), .B(core_key_33_), .Y(core__abc_22172_new_n7803_));
AND2X2 AND2X2_4406 ( .A(core__abc_22172_new_n7804_), .B(core__abc_22172_new_n7805_), .Y(core__abc_22172_new_n7806_));
AND2X2 AND2X2_4407 ( .A(core__abc_22172_new_n7806_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n7807_));
AND2X2 AND2X2_4408 ( .A(core__abc_22172_new_n7114_), .B(core__abc_22172_new_n7808_), .Y(core__abc_22172_new_n7809_));
AND2X2 AND2X2_4409 ( .A(core__abc_22172_new_n7810_), .B(reset_n), .Y(core__0v2_reg_63_0__33_));
AND2X2 AND2X2_441 ( .A(_abc_19873_new_n1657_), .B(reset_n), .Y(_0word3_reg_31_0__12_));
AND2X2 AND2X2_4410 ( .A(core__abc_22172_new_n7812_), .B(core__abc_22172_new_n7813_), .Y(core__abc_22172_new_n7814_));
AND2X2 AND2X2_4411 ( .A(core__abc_22172_new_n7814_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n7815_));
AND2X2 AND2X2_4412 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n7816_), .Y(core__abc_22172_new_n7817_));
AND2X2 AND2X2_4413 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_34_), .Y(core__abc_22172_new_n7818_));
AND2X2 AND2X2_4414 ( .A(core__abc_22172_new_n7822_), .B(reset_n), .Y(core__abc_22172_new_n7823_));
AND2X2 AND2X2_4415 ( .A(core__abc_22172_new_n7823_), .B(core__abc_22172_new_n7821_), .Y(core__0v2_reg_63_0__34_));
AND2X2 AND2X2_4416 ( .A(core__abc_22172_new_n7826_), .B(core__abc_22172_new_n6790_), .Y(core__abc_22172_new_n7827_));
AND2X2 AND2X2_4417 ( .A(core__abc_22172_new_n7828_), .B(core__abc_22172_new_n7825_), .Y(core__abc_22172_new_n7829_));
AND2X2 AND2X2_4418 ( .A(core__abc_22172_new_n7827_), .B(core__abc_22172_new_n6818_), .Y(core__abc_22172_new_n7830_));
AND2X2 AND2X2_4419 ( .A(core__abc_22172_new_n7832_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n7833_));
AND2X2 AND2X2_442 ( .A(core_siphash_valid_reg), .B(core_siphash_word_109_), .Y(_abc_19873_new_n1659_));
AND2X2 AND2X2_4420 ( .A(core__abc_22172_new_n3214_), .B(core_key_35_), .Y(core__abc_22172_new_n7834_));
AND2X2 AND2X2_4421 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_35_), .Y(core__abc_22172_new_n7835_));
AND2X2 AND2X2_4422 ( .A(core__abc_22172_new_n7839_), .B(reset_n), .Y(core__abc_22172_new_n7840_));
AND2X2 AND2X2_4423 ( .A(core__abc_22172_new_n7838_), .B(core__abc_22172_new_n7840_), .Y(core__0v2_reg_63_0__35_));
AND2X2 AND2X2_4424 ( .A(core__abc_22172_new_n7842_), .B(core__abc_22172_new_n7843_), .Y(core__abc_22172_new_n7844_));
AND2X2 AND2X2_4425 ( .A(core__abc_22172_new_n7844_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n7845_));
AND2X2 AND2X2_4426 ( .A(core__abc_22172_new_n3214_), .B(core_key_36_), .Y(core__abc_22172_new_n7846_));
AND2X2 AND2X2_4427 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_36_), .Y(core__abc_22172_new_n7847_));
AND2X2 AND2X2_4428 ( .A(core__abc_22172_new_n7851_), .B(reset_n), .Y(core__abc_22172_new_n7852_));
AND2X2 AND2X2_4429 ( .A(core__abc_22172_new_n7850_), .B(core__abc_22172_new_n7852_), .Y(core__0v2_reg_63_0__36_));
AND2X2 AND2X2_443 ( .A(_abc_19873_new_n1607_), .B(word3_reg_13_), .Y(_abc_19873_new_n1660_));
AND2X2 AND2X2_4430 ( .A(core__abc_22172_new_n7855_), .B(core__abc_22172_new_n6776_), .Y(core__abc_22172_new_n7856_));
AND2X2 AND2X2_4431 ( .A(core__abc_22172_new_n7854_), .B(core__abc_22172_new_n7856_), .Y(core__abc_22172_new_n7857_));
AND2X2 AND2X2_4432 ( .A(core__abc_22172_new_n7858_), .B(core__abc_22172_new_n7859_), .Y(core__abc_22172_new_n7860_));
AND2X2 AND2X2_4433 ( .A(core__abc_22172_new_n7861_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n7862_));
AND2X2 AND2X2_4434 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n7863_), .Y(core__abc_22172_new_n7864_));
AND2X2 AND2X2_4435 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_37_), .Y(core__abc_22172_new_n7865_));
AND2X2 AND2X2_4436 ( .A(core__abc_22172_new_n7869_), .B(reset_n), .Y(core__abc_22172_new_n7870_));
AND2X2 AND2X2_4437 ( .A(core__abc_22172_new_n7868_), .B(core__abc_22172_new_n7870_), .Y(core__0v2_reg_63_0__37_));
AND2X2 AND2X2_4438 ( .A(core__abc_22172_new_n6827_), .B(core__abc_22172_new_n6766_), .Y(core__abc_22172_new_n7872_));
AND2X2 AND2X2_4439 ( .A(core__abc_22172_new_n7873_), .B(core__abc_22172_new_n7874_), .Y(core__abc_22172_new_n7875_));
AND2X2 AND2X2_444 ( .A(_abc_19873_new_n1661_), .B(reset_n), .Y(_0word3_reg_31_0__13_));
AND2X2 AND2X2_4440 ( .A(core__abc_22172_new_n7875_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n7876_));
AND2X2 AND2X2_4441 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n7877_), .Y(core__abc_22172_new_n7878_));
AND2X2 AND2X2_4442 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_38_), .Y(core__abc_22172_new_n7879_));
AND2X2 AND2X2_4443 ( .A(core__abc_22172_new_n7883_), .B(reset_n), .Y(core__abc_22172_new_n7884_));
AND2X2 AND2X2_4444 ( .A(core__abc_22172_new_n7882_), .B(core__abc_22172_new_n7884_), .Y(core__0v2_reg_63_0__38_));
AND2X2 AND2X2_4445 ( .A(core__abc_22172_new_n7890_), .B(core__abc_22172_new_n7887_), .Y(core__abc_22172_new_n7891_));
AND2X2 AND2X2_4446 ( .A(core__abc_22172_new_n7891_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n7892_));
AND2X2 AND2X2_4447 ( .A(core__abc_22172_new_n3214_), .B(core_key_39_), .Y(core__abc_22172_new_n7893_));
AND2X2 AND2X2_4448 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_39_), .Y(core__abc_22172_new_n7894_));
AND2X2 AND2X2_4449 ( .A(core__abc_22172_new_n7898_), .B(reset_n), .Y(core__abc_22172_new_n7899_));
AND2X2 AND2X2_445 ( .A(core_siphash_valid_reg), .B(core_siphash_word_110_), .Y(_abc_19873_new_n1663_));
AND2X2 AND2X2_4450 ( .A(core__abc_22172_new_n7897_), .B(core__abc_22172_new_n7899_), .Y(core__0v2_reg_63_0__39_));
AND2X2 AND2X2_4451 ( .A(core__abc_22172_new_n6829_), .B(core__abc_22172_new_n6833_), .Y(core__abc_22172_new_n7901_));
AND2X2 AND2X2_4452 ( .A(core__abc_22172_new_n7902_), .B(core__abc_22172_new_n7903_), .Y(core__abc_22172_new_n7904_));
AND2X2 AND2X2_4453 ( .A(core__abc_22172_new_n7904_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n7905_));
AND2X2 AND2X2_4454 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n7906_), .Y(core__abc_22172_new_n7907_));
AND2X2 AND2X2_4455 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_40_), .Y(core__abc_22172_new_n7908_));
AND2X2 AND2X2_4456 ( .A(core__abc_22172_new_n7912_), .B(reset_n), .Y(core__abc_22172_new_n7913_));
AND2X2 AND2X2_4457 ( .A(core__abc_22172_new_n7911_), .B(core__abc_22172_new_n7913_), .Y(core__0v2_reg_63_0__40_));
AND2X2 AND2X2_4458 ( .A(core__abc_22172_new_n7917_), .B(core__abc_22172_new_n7915_), .Y(core__abc_22172_new_n7918_));
AND2X2 AND2X2_4459 ( .A(core__abc_22172_new_n7916_), .B(core__abc_22172_new_n6830_), .Y(core__abc_22172_new_n7919_));
AND2X2 AND2X2_446 ( .A(_abc_19873_new_n1607_), .B(word3_reg_14_), .Y(_abc_19873_new_n1664_));
AND2X2 AND2X2_4460 ( .A(core__abc_22172_new_n7921_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n7922_));
AND2X2 AND2X2_4461 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n7923_), .Y(core__abc_22172_new_n7924_));
AND2X2 AND2X2_4462 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_41_), .Y(core__abc_22172_new_n7925_));
AND2X2 AND2X2_4463 ( .A(core__abc_22172_new_n7929_), .B(reset_n), .Y(core__abc_22172_new_n7930_));
AND2X2 AND2X2_4464 ( .A(core__abc_22172_new_n7928_), .B(core__abc_22172_new_n7930_), .Y(core__0v2_reg_63_0__41_));
AND2X2 AND2X2_4465 ( .A(core__abc_22172_new_n6829_), .B(core__abc_22172_new_n6834_), .Y(core__abc_22172_new_n7932_));
AND2X2 AND2X2_4466 ( .A(core__abc_22172_new_n7933_), .B(core__abc_22172_new_n6728_), .Y(core__abc_22172_new_n7934_));
AND2X2 AND2X2_4467 ( .A(core__abc_22172_new_n7935_), .B(core__abc_22172_new_n7936_), .Y(core__abc_22172_new_n7937_));
AND2X2 AND2X2_4468 ( .A(core__abc_22172_new_n7937_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n7938_));
AND2X2 AND2X2_4469 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n7939_), .Y(core__abc_22172_new_n7940_));
AND2X2 AND2X2_447 ( .A(_abc_19873_new_n1665_), .B(reset_n), .Y(_0word3_reg_31_0__14_));
AND2X2 AND2X2_4470 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_42_), .Y(core__abc_22172_new_n7941_));
AND2X2 AND2X2_4471 ( .A(core__abc_22172_new_n7945_), .B(reset_n), .Y(core__abc_22172_new_n7946_));
AND2X2 AND2X2_4472 ( .A(core__abc_22172_new_n7944_), .B(core__abc_22172_new_n7946_), .Y(core__0v2_reg_63_0__42_));
AND2X2 AND2X2_4473 ( .A(core__abc_22172_new_n7950_), .B(core__abc_22172_new_n7948_), .Y(core__abc_22172_new_n7951_));
AND2X2 AND2X2_4474 ( .A(core__abc_22172_new_n7949_), .B(core__abc_22172_new_n6725_), .Y(core__abc_22172_new_n7952_));
AND2X2 AND2X2_4475 ( .A(core__abc_22172_new_n7954_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n7955_));
AND2X2 AND2X2_4476 ( .A(core__abc_22172_new_n3214_), .B(core_key_43_), .Y(core__abc_22172_new_n7956_));
AND2X2 AND2X2_4477 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_43_), .Y(core__abc_22172_new_n7957_));
AND2X2 AND2X2_4478 ( .A(core__abc_22172_new_n7961_), .B(reset_n), .Y(core__abc_22172_new_n7962_));
AND2X2 AND2X2_4479 ( .A(core__abc_22172_new_n7960_), .B(core__abc_22172_new_n7962_), .Y(core__0v2_reg_63_0__43_));
AND2X2 AND2X2_448 ( .A(core_siphash_valid_reg), .B(core_siphash_word_111_), .Y(_abc_19873_new_n1667_));
AND2X2 AND2X2_4480 ( .A(core__abc_22172_new_n6837_), .B(core__abc_22172_new_n6706_), .Y(core__abc_22172_new_n7964_));
AND2X2 AND2X2_4481 ( .A(core__abc_22172_new_n7965_), .B(core__abc_22172_new_n7966_), .Y(core__abc_22172_new_n7967_));
AND2X2 AND2X2_4482 ( .A(core__abc_22172_new_n7967_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n7968_));
AND2X2 AND2X2_4483 ( .A(core__abc_22172_new_n3214_), .B(core_key_44_), .Y(core__abc_22172_new_n7969_));
AND2X2 AND2X2_4484 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_44_), .Y(core__abc_22172_new_n7970_));
AND2X2 AND2X2_4485 ( .A(core__abc_22172_new_n7974_), .B(reset_n), .Y(core__abc_22172_new_n7975_));
AND2X2 AND2X2_4486 ( .A(core__abc_22172_new_n7973_), .B(core__abc_22172_new_n7975_), .Y(core__0v2_reg_63_0__44_));
AND2X2 AND2X2_4487 ( .A(core__abc_22172_new_n7965_), .B(core__abc_22172_new_n6694_), .Y(core__abc_22172_new_n7978_));
AND2X2 AND2X2_4488 ( .A(core__abc_22172_new_n7979_), .B(core__abc_22172_new_n7977_), .Y(core__abc_22172_new_n7980_));
AND2X2 AND2X2_4489 ( .A(core__abc_22172_new_n7978_), .B(core__abc_22172_new_n6703_), .Y(core__abc_22172_new_n7981_));
AND2X2 AND2X2_449 ( .A(_abc_19873_new_n1607_), .B(word3_reg_15_), .Y(_abc_19873_new_n1668_));
AND2X2 AND2X2_4490 ( .A(core__abc_22172_new_n7982_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n7983_));
AND2X2 AND2X2_4491 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n7984_), .Y(core__abc_22172_new_n7985_));
AND2X2 AND2X2_4492 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_45_), .Y(core__abc_22172_new_n7986_));
AND2X2 AND2X2_4493 ( .A(core__abc_22172_new_n7990_), .B(reset_n), .Y(core__abc_22172_new_n7991_));
AND2X2 AND2X2_4494 ( .A(core__abc_22172_new_n7989_), .B(core__abc_22172_new_n7991_), .Y(core__0v2_reg_63_0__45_));
AND2X2 AND2X2_4495 ( .A(core__abc_22172_new_n7965_), .B(core__abc_22172_new_n6695_), .Y(core__abc_22172_new_n7993_));
AND2X2 AND2X2_4496 ( .A(core__abc_22172_new_n7994_), .B(core__abc_22172_new_n6677_), .Y(core__abc_22172_new_n7995_));
AND2X2 AND2X2_4497 ( .A(core__abc_22172_new_n7999_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8000_));
AND2X2 AND2X2_4498 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n8001_), .Y(core__abc_22172_new_n8002_));
AND2X2 AND2X2_4499 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_46_), .Y(core__abc_22172_new_n8003_));
AND2X2 AND2X2_45 ( .A(_abc_19873_new_n900_), .B(_abc_19873_new_n906_), .Y(_abc_19873_new_n930_));
AND2X2 AND2X2_450 ( .A(_abc_19873_new_n1669_), .B(reset_n), .Y(_0word3_reg_31_0__15_));
AND2X2 AND2X2_4500 ( .A(core__abc_22172_new_n8007_), .B(reset_n), .Y(core__abc_22172_new_n8008_));
AND2X2 AND2X2_4501 ( .A(core__abc_22172_new_n8006_), .B(core__abc_22172_new_n8008_), .Y(core__0v2_reg_63_0__46_));
AND2X2 AND2X2_4502 ( .A(core__abc_22172_new_n8012_), .B(core__abc_22172_new_n8010_), .Y(core__abc_22172_new_n8013_));
AND2X2 AND2X2_4503 ( .A(core__abc_22172_new_n8011_), .B(core__abc_22172_new_n6670_), .Y(core__abc_22172_new_n8014_));
AND2X2 AND2X2_4504 ( .A(core__abc_22172_new_n8016_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8017_));
AND2X2 AND2X2_4505 ( .A(core__abc_22172_new_n3214_), .B(core_key_47_), .Y(core__abc_22172_new_n8018_));
AND2X2 AND2X2_4506 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_47_), .Y(core__abc_22172_new_n8019_));
AND2X2 AND2X2_4507 ( .A(core__abc_22172_new_n8023_), .B(reset_n), .Y(core__abc_22172_new_n8024_));
AND2X2 AND2X2_4508 ( .A(core__abc_22172_new_n8022_), .B(core__abc_22172_new_n8024_), .Y(core__0v2_reg_63_0__47_));
AND2X2 AND2X2_4509 ( .A(core__abc_22172_new_n8026_), .B(core__abc_22172_new_n6843_), .Y(core__abc_22172_new_n8027_));
AND2X2 AND2X2_451 ( .A(core_siphash_valid_reg), .B(core_siphash_word_112_), .Y(_abc_19873_new_n1671_));
AND2X2 AND2X2_4510 ( .A(core__abc_22172_new_n6839_), .B(core__abc_22172_new_n6844_), .Y(core__abc_22172_new_n8028_));
AND2X2 AND2X2_4511 ( .A(core__abc_22172_new_n8030_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8031_));
AND2X2 AND2X2_4512 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n8032_), .Y(core__abc_22172_new_n8033_));
AND2X2 AND2X2_4513 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_48_), .Y(core__abc_22172_new_n8034_));
AND2X2 AND2X2_4514 ( .A(core__abc_22172_new_n8038_), .B(reset_n), .Y(core__abc_22172_new_n8039_));
AND2X2 AND2X2_4515 ( .A(core__abc_22172_new_n8037_), .B(core__abc_22172_new_n8039_), .Y(core__0v2_reg_63_0__48_));
AND2X2 AND2X2_4516 ( .A(core__abc_22172_new_n8042_), .B(core__abc_22172_new_n8041_), .Y(core__abc_22172_new_n8043_));
AND2X2 AND2X2_4517 ( .A(core__abc_22172_new_n8044_), .B(core__abc_22172_new_n6841_), .Y(core__abc_22172_new_n8045_));
AND2X2 AND2X2_4518 ( .A(core__abc_22172_new_n8046_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8047_));
AND2X2 AND2X2_4519 ( .A(core__abc_22172_new_n3214_), .B(core_key_49_), .Y(core__abc_22172_new_n8048_));
AND2X2 AND2X2_452 ( .A(_abc_19873_new_n1607_), .B(word3_reg_16_), .Y(_abc_19873_new_n1672_));
AND2X2 AND2X2_4520 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_49_), .Y(core__abc_22172_new_n8049_));
AND2X2 AND2X2_4521 ( .A(core__abc_22172_new_n8053_), .B(reset_n), .Y(core__abc_22172_new_n8054_));
AND2X2 AND2X2_4522 ( .A(core__abc_22172_new_n8052_), .B(core__abc_22172_new_n8054_), .Y(core__0v2_reg_63_0__49_));
AND2X2 AND2X2_4523 ( .A(core__abc_22172_new_n6839_), .B(core__abc_22172_new_n6845_), .Y(core__abc_22172_new_n8056_));
AND2X2 AND2X2_4524 ( .A(core__abc_22172_new_n8057_), .B(core__abc_22172_new_n6616_), .Y(core__abc_22172_new_n8058_));
AND2X2 AND2X2_4525 ( .A(core__abc_22172_new_n8059_), .B(core__abc_22172_new_n8060_), .Y(core__abc_22172_new_n8061_));
AND2X2 AND2X2_4526 ( .A(core__abc_22172_new_n8061_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8062_));
AND2X2 AND2X2_4527 ( .A(core__abc_22172_new_n3214_), .B(core_key_50_), .Y(core__abc_22172_new_n8063_));
AND2X2 AND2X2_4528 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_50_), .Y(core__abc_22172_new_n8064_));
AND2X2 AND2X2_4529 ( .A(core__abc_22172_new_n8068_), .B(reset_n), .Y(core__abc_22172_new_n8069_));
AND2X2 AND2X2_453 ( .A(_abc_19873_new_n1673_), .B(reset_n), .Y(_0word3_reg_31_0__16_));
AND2X2 AND2X2_4530 ( .A(core__abc_22172_new_n8067_), .B(core__abc_22172_new_n8069_), .Y(core__0v2_reg_63_0__50_));
AND2X2 AND2X2_4531 ( .A(core__abc_22172_new_n8059_), .B(core__abc_22172_new_n6646_), .Y(core__abc_22172_new_n8072_));
AND2X2 AND2X2_4532 ( .A(core__abc_22172_new_n8072_), .B(core__abc_22172_new_n8071_), .Y(core__abc_22172_new_n8073_));
AND2X2 AND2X2_4533 ( .A(core__abc_22172_new_n8074_), .B(core__abc_22172_new_n8075_), .Y(core__abc_22172_new_n8076_));
AND2X2 AND2X2_4534 ( .A(core__abc_22172_new_n8076_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8077_));
AND2X2 AND2X2_4535 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n8078_), .Y(core__abc_22172_new_n8079_));
AND2X2 AND2X2_4536 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_51_), .Y(core__abc_22172_new_n8080_));
AND2X2 AND2X2_4537 ( .A(core__abc_22172_new_n8084_), .B(reset_n), .Y(core__abc_22172_new_n8085_));
AND2X2 AND2X2_4538 ( .A(core__abc_22172_new_n8083_), .B(core__abc_22172_new_n8085_), .Y(core__0v2_reg_63_0__51_));
AND2X2 AND2X2_4539 ( .A(core__abc_22172_new_n8059_), .B(core__abc_22172_new_n6647_), .Y(core__abc_22172_new_n8087_));
AND2X2 AND2X2_454 ( .A(core_siphash_valid_reg), .B(core_siphash_word_113_), .Y(_abc_19873_new_n1675_));
AND2X2 AND2X2_4540 ( .A(core__abc_22172_new_n8088_), .B(core__abc_22172_new_n6623_), .Y(core__abc_22172_new_n8089_));
AND2X2 AND2X2_4541 ( .A(core__abc_22172_new_n8089_), .B(core__abc_22172_new_n6605_), .Y(core__abc_22172_new_n8090_));
AND2X2 AND2X2_4542 ( .A(core__abc_22172_new_n8091_), .B(core__abc_22172_new_n6604_), .Y(core__abc_22172_new_n8092_));
AND2X2 AND2X2_4543 ( .A(core__abc_22172_new_n8094_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8095_));
AND2X2 AND2X2_4544 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n8096_), .Y(core__abc_22172_new_n8097_));
AND2X2 AND2X2_4545 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_52_), .Y(core__abc_22172_new_n8098_));
AND2X2 AND2X2_4546 ( .A(core__abc_22172_new_n8102_), .B(reset_n), .Y(core__abc_22172_new_n8103_));
AND2X2 AND2X2_4547 ( .A(core__abc_22172_new_n8101_), .B(core__abc_22172_new_n8103_), .Y(core__0v2_reg_63_0__52_));
AND2X2 AND2X2_4548 ( .A(core__abc_22172_new_n8106_), .B(core__abc_22172_new_n8105_), .Y(core__abc_22172_new_n8107_));
AND2X2 AND2X2_4549 ( .A(core__abc_22172_new_n8108_), .B(core__abc_22172_new_n8109_), .Y(core__abc_22172_new_n8110_));
AND2X2 AND2X2_455 ( .A(_abc_19873_new_n1607_), .B(word3_reg_17_), .Y(_abc_19873_new_n1676_));
AND2X2 AND2X2_4550 ( .A(core__abc_22172_new_n8111_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8112_));
AND2X2 AND2X2_4551 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n8113_), .Y(core__abc_22172_new_n8114_));
AND2X2 AND2X2_4552 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_53_), .Y(core__abc_22172_new_n8115_));
AND2X2 AND2X2_4553 ( .A(core__abc_22172_new_n8119_), .B(reset_n), .Y(core__abc_22172_new_n8120_));
AND2X2 AND2X2_4554 ( .A(core__abc_22172_new_n8118_), .B(core__abc_22172_new_n8120_), .Y(core__0v2_reg_63_0__53_));
AND2X2 AND2X2_4555 ( .A(core__abc_22172_new_n8089_), .B(core__abc_22172_new_n6606_), .Y(core__abc_22172_new_n8122_));
AND2X2 AND2X2_4556 ( .A(core__abc_22172_new_n8123_), .B(core__abc_22172_new_n6587_), .Y(core__abc_22172_new_n8124_));
AND2X2 AND2X2_4557 ( .A(core__abc_22172_new_n8125_), .B(core__abc_22172_new_n8126_), .Y(core__abc_22172_new_n8127_));
AND2X2 AND2X2_4558 ( .A(core__abc_22172_new_n8127_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8128_));
AND2X2 AND2X2_4559 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n8129_), .Y(core__abc_22172_new_n8130_));
AND2X2 AND2X2_456 ( .A(_abc_19873_new_n1677_), .B(reset_n), .Y(_0word3_reg_31_0__17_));
AND2X2 AND2X2_4560 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_54_), .Y(core__abc_22172_new_n8131_));
AND2X2 AND2X2_4561 ( .A(core__abc_22172_new_n8135_), .B(reset_n), .Y(core__abc_22172_new_n8136_));
AND2X2 AND2X2_4562 ( .A(core__abc_22172_new_n8134_), .B(core__abc_22172_new_n8136_), .Y(core__0v2_reg_63_0__54_));
AND2X2 AND2X2_4563 ( .A(core__abc_22172_new_n8140_), .B(core__abc_22172_new_n8138_), .Y(core__abc_22172_new_n8141_));
AND2X2 AND2X2_4564 ( .A(core__abc_22172_new_n8139_), .B(core__abc_22172_new_n6578_), .Y(core__abc_22172_new_n8142_));
AND2X2 AND2X2_4565 ( .A(core__abc_22172_new_n8144_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8145_));
AND2X2 AND2X2_4566 ( .A(core__abc_22172_new_n3214_), .B(core_key_55_), .Y(core__abc_22172_new_n8146_));
AND2X2 AND2X2_4567 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_55_), .Y(core__abc_22172_new_n8147_));
AND2X2 AND2X2_4568 ( .A(core__abc_22172_new_n8151_), .B(reset_n), .Y(core__abc_22172_new_n8152_));
AND2X2 AND2X2_4569 ( .A(core__abc_22172_new_n8150_), .B(core__abc_22172_new_n8152_), .Y(core__0v2_reg_63_0__55_));
AND2X2 AND2X2_457 ( .A(core_siphash_valid_reg), .B(core_siphash_word_114_), .Y(_abc_19873_new_n1679_));
AND2X2 AND2X2_4570 ( .A(core__abc_22172_new_n8154_), .B(core__abc_22172_new_n6565_), .Y(core__abc_22172_new_n8155_));
AND2X2 AND2X2_4571 ( .A(core__abc_22172_new_n6849_), .B(core__abc_22172_new_n6566_), .Y(core__abc_22172_new_n8156_));
AND2X2 AND2X2_4572 ( .A(core__abc_22172_new_n8158_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8159_));
AND2X2 AND2X2_4573 ( .A(core__abc_22172_new_n3214_), .B(core_key_56_), .Y(core__abc_22172_new_n8160_));
AND2X2 AND2X2_4574 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_56_), .Y(core__abc_22172_new_n8161_));
AND2X2 AND2X2_4575 ( .A(core__abc_22172_new_n8165_), .B(reset_n), .Y(core__abc_22172_new_n8166_));
AND2X2 AND2X2_4576 ( .A(core__abc_22172_new_n8164_), .B(core__abc_22172_new_n8166_), .Y(core__0v2_reg_63_0__56_));
AND2X2 AND2X2_4577 ( .A(core__abc_22172_new_n8169_), .B(core__abc_22172_new_n6540_), .Y(core__abc_22172_new_n8170_));
AND2X2 AND2X2_4578 ( .A(core__abc_22172_new_n8170_), .B(core__abc_22172_new_n8168_), .Y(core__abc_22172_new_n8171_));
AND2X2 AND2X2_4579 ( .A(core__abc_22172_new_n8172_), .B(core__abc_22172_new_n8173_), .Y(core__abc_22172_new_n8174_));
AND2X2 AND2X2_458 ( .A(_abc_19873_new_n1607_), .B(word3_reg_18_), .Y(_abc_19873_new_n1680_));
AND2X2 AND2X2_4580 ( .A(core__abc_22172_new_n8174_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8175_));
AND2X2 AND2X2_4581 ( .A(core__abc_22172_new_n3214_), .B(core_key_57_), .Y(core__abc_22172_new_n8176_));
AND2X2 AND2X2_4582 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_57_), .Y(core__abc_22172_new_n8177_));
AND2X2 AND2X2_4583 ( .A(core__abc_22172_new_n8181_), .B(reset_n), .Y(core__abc_22172_new_n8182_));
AND2X2 AND2X2_4584 ( .A(core__abc_22172_new_n8180_), .B(core__abc_22172_new_n8182_), .Y(core__0v2_reg_63_0__57_));
AND2X2 AND2X2_4585 ( .A(core__abc_22172_new_n6849_), .B(core__abc_22172_new_n6567_), .Y(core__abc_22172_new_n8184_));
AND2X2 AND2X2_4586 ( .A(core__abc_22172_new_n8185_), .B(core__abc_22172_new_n6524_), .Y(core__abc_22172_new_n8186_));
AND2X2 AND2X2_4587 ( .A(core__abc_22172_new_n8187_), .B(core__abc_22172_new_n8188_), .Y(core__abc_22172_new_n8189_));
AND2X2 AND2X2_4588 ( .A(core__abc_22172_new_n8189_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8190_));
AND2X2 AND2X2_4589 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n8191_), .Y(core__abc_22172_new_n8192_));
AND2X2 AND2X2_459 ( .A(_abc_19873_new_n1681_), .B(reset_n), .Y(_0word3_reg_31_0__18_));
AND2X2 AND2X2_4590 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_58_), .Y(core__abc_22172_new_n8193_));
AND2X2 AND2X2_4591 ( .A(core__abc_22172_new_n8197_), .B(reset_n), .Y(core__abc_22172_new_n8198_));
AND2X2 AND2X2_4592 ( .A(core__abc_22172_new_n8196_), .B(core__abc_22172_new_n8198_), .Y(core__0v2_reg_63_0__58_));
AND2X2 AND2X2_4593 ( .A(core__abc_22172_new_n8187_), .B(core__abc_22172_new_n6547_), .Y(core__abc_22172_new_n8201_));
AND2X2 AND2X2_4594 ( .A(core__abc_22172_new_n8202_), .B(core__abc_22172_new_n8200_), .Y(core__abc_22172_new_n8203_));
AND2X2 AND2X2_4595 ( .A(core__abc_22172_new_n8201_), .B(core__abc_22172_new_n6515_), .Y(core__abc_22172_new_n8204_));
AND2X2 AND2X2_4596 ( .A(core__abc_22172_new_n8205_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8206_));
AND2X2 AND2X2_4597 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n8207_), .Y(core__abc_22172_new_n8208_));
AND2X2 AND2X2_4598 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_59_), .Y(core__abc_22172_new_n8209_));
AND2X2 AND2X2_4599 ( .A(core__abc_22172_new_n8213_), .B(reset_n), .Y(core__abc_22172_new_n8214_));
AND2X2 AND2X2_46 ( .A(_abc_19873_new_n930_), .B(word0_reg_0_), .Y(_abc_19873_new_n931_));
AND2X2 AND2X2_460 ( .A(core_siphash_valid_reg), .B(core_siphash_word_115_), .Y(_abc_19873_new_n1683_));
AND2X2 AND2X2_4600 ( .A(core__abc_22172_new_n8212_), .B(core__abc_22172_new_n8214_), .Y(core__0v2_reg_63_0__59_));
AND2X2 AND2X2_4601 ( .A(core__abc_22172_new_n8202_), .B(core__abc_22172_new_n6514_), .Y(core__abc_22172_new_n8216_));
AND2X2 AND2X2_4602 ( .A(core__abc_22172_new_n8217_), .B(core__abc_22172_new_n6512_), .Y(core__abc_22172_new_n8218_));
AND2X2 AND2X2_4603 ( .A(core__abc_22172_new_n8219_), .B(core__abc_22172_new_n6504_), .Y(core__abc_22172_new_n8220_));
AND2X2 AND2X2_4604 ( .A(core__abc_22172_new_n8218_), .B(core__abc_22172_new_n6503_), .Y(core__abc_22172_new_n8221_));
AND2X2 AND2X2_4605 ( .A(core__abc_22172_new_n8223_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8224_));
AND2X2 AND2X2_4606 ( .A(core__abc_22172_new_n3214_), .B(core_key_60_), .Y(core__abc_22172_new_n8225_));
AND2X2 AND2X2_4607 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_60_), .Y(core__abc_22172_new_n8226_));
AND2X2 AND2X2_4608 ( .A(core__abc_22172_new_n8230_), .B(reset_n), .Y(core__abc_22172_new_n8231_));
AND2X2 AND2X2_4609 ( .A(core__abc_22172_new_n8229_), .B(core__abc_22172_new_n8231_), .Y(core__0v2_reg_63_0__60_));
AND2X2 AND2X2_461 ( .A(_abc_19873_new_n1607_), .B(word3_reg_19_), .Y(_abc_19873_new_n1684_));
AND2X2 AND2X2_4610 ( .A(core__abc_22172_new_n8234_), .B(core__abc_22172_new_n8233_), .Y(core__abc_22172_new_n8235_));
AND2X2 AND2X2_4611 ( .A(core__abc_22172_new_n8236_), .B(core__abc_22172_new_n8237_), .Y(core__abc_22172_new_n8238_));
AND2X2 AND2X2_4612 ( .A(core__abc_22172_new_n8239_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8240_));
AND2X2 AND2X2_4613 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n8241_), .Y(core__abc_22172_new_n8242_));
AND2X2 AND2X2_4614 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_61_), .Y(core__abc_22172_new_n8243_));
AND2X2 AND2X2_4615 ( .A(core__abc_22172_new_n8247_), .B(reset_n), .Y(core__abc_22172_new_n8248_));
AND2X2 AND2X2_4616 ( .A(core__abc_22172_new_n8246_), .B(core__abc_22172_new_n8248_), .Y(core__0v2_reg_63_0__61_));
AND2X2 AND2X2_4617 ( .A(core__abc_22172_new_n8219_), .B(core__abc_22172_new_n6505_), .Y(core__abc_22172_new_n8250_));
AND2X2 AND2X2_4618 ( .A(core__abc_22172_new_n8251_), .B(core__abc_22172_new_n6483_), .Y(core__abc_22172_new_n8252_));
AND2X2 AND2X2_4619 ( .A(core__abc_22172_new_n8253_), .B(core__abc_22172_new_n8254_), .Y(core__abc_22172_new_n8255_));
AND2X2 AND2X2_462 ( .A(_abc_19873_new_n1685_), .B(reset_n), .Y(_0word3_reg_31_0__19_));
AND2X2 AND2X2_4620 ( .A(core__abc_22172_new_n8255_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8256_));
AND2X2 AND2X2_4621 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n8257_), .Y(core__abc_22172_new_n8258_));
AND2X2 AND2X2_4622 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_62_), .Y(core__abc_22172_new_n8259_));
AND2X2 AND2X2_4623 ( .A(core__abc_22172_new_n8263_), .B(reset_n), .Y(core__abc_22172_new_n8264_));
AND2X2 AND2X2_4624 ( .A(core__abc_22172_new_n8262_), .B(core__abc_22172_new_n8264_), .Y(core__0v2_reg_63_0__62_));
AND2X2 AND2X2_4625 ( .A(core__abc_22172_new_n8253_), .B(core__abc_22172_new_n6480_), .Y(core__abc_22172_new_n8267_));
AND2X2 AND2X2_4626 ( .A(core__abc_22172_new_n8267_), .B(core__abc_22172_new_n8266_), .Y(core__abc_22172_new_n8268_));
AND2X2 AND2X2_4627 ( .A(core__abc_22172_new_n8272_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8273_));
AND2X2 AND2X2_4628 ( .A(core__abc_22172_new_n3214_), .B(core_key_63_), .Y(core__abc_22172_new_n8274_));
AND2X2 AND2X2_4629 ( .A(core__abc_22172_new_n3196_), .B(core_v2_reg_63_), .Y(core__abc_22172_new_n8275_));
AND2X2 AND2X2_463 ( .A(core_siphash_valid_reg), .B(core_siphash_word_116_), .Y(_abc_19873_new_n1687_));
AND2X2 AND2X2_4630 ( .A(core__abc_22172_new_n8279_), .B(reset_n), .Y(core__abc_22172_new_n8280_));
AND2X2 AND2X2_4631 ( .A(core__abc_22172_new_n8278_), .B(core__abc_22172_new_n8280_), .Y(core__0v2_reg_63_0__63_));
AND2X2 AND2X2_4632 ( .A(core__abc_22172_new_n3213_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n8282_));
AND2X2 AND2X2_4633 ( .A(core__abc_22172_new_n8283_), .B(core_v1_reg_0_), .Y(core__abc_22172_new_n8284_));
AND2X2 AND2X2_4634 ( .A(core__abc_22172_new_n7297_), .B(core__abc_22172_new_n7795_), .Y(core__abc_22172_new_n8285_));
AND2X2 AND2X2_4635 ( .A(core__abc_22172_new_n3205_), .B(core__abc_22172_new_n7793_), .Y(core__abc_22172_new_n8286_));
AND2X2 AND2X2_4636 ( .A(core__abc_22172_new_n7294_), .B(core__abc_22172_new_n8286_), .Y(core__abc_22172_new_n8287_));
AND2X2 AND2X2_4637 ( .A(core__abc_22172_new_n1218_), .B(core_siphash_ctrl_reg_5_), .Y(core__abc_22172_new_n8288_));
AND2X2 AND2X2_4638 ( .A(core__abc_22172_new_n3198_), .B(core__abc_22172_new_n8288_), .Y(core__abc_22172_new_n8289_));
AND2X2 AND2X2_4639 ( .A(core__abc_22172_new_n8289_), .B(core__abc_22172_new_n6680_), .Y(core__abc_22172_new_n8290_));
AND2X2 AND2X2_464 ( .A(_abc_19873_new_n1607_), .B(word3_reg_20_), .Y(_abc_19873_new_n1688_));
AND2X2 AND2X2_4640 ( .A(core__abc_22172_new_n8293_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n8294_));
AND2X2 AND2X2_4641 ( .A(core__abc_22172_new_n8295_), .B(reset_n), .Y(core__0v1_reg_63_0__0_));
AND2X2 AND2X2_4642 ( .A(core__abc_22172_new_n8299_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8300_));
AND2X2 AND2X2_4643 ( .A(core__abc_22172_new_n8300_), .B(core__abc_22172_new_n8297_), .Y(core__abc_22172_new_n8301_));
AND2X2 AND2X2_4644 ( .A(core_key_65_), .B(core_long), .Y(core__abc_22172_new_n8303_));
AND2X2 AND2X2_4645 ( .A(core__abc_22172_new_n8304_), .B(core__abc_22172_new_n8302_), .Y(core__abc_22172_new_n8305_));
AND2X2 AND2X2_4646 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n8305_), .Y(core__abc_22172_new_n8306_));
AND2X2 AND2X2_4647 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_1_), .Y(core__abc_22172_new_n8307_));
AND2X2 AND2X2_4648 ( .A(core__abc_22172_new_n8311_), .B(reset_n), .Y(core__abc_22172_new_n8312_));
AND2X2 AND2X2_4649 ( .A(core__abc_22172_new_n8310_), .B(core__abc_22172_new_n8312_), .Y(core__0v1_reg_63_0__1_));
AND2X2 AND2X2_465 ( .A(_abc_19873_new_n1689_), .B(reset_n), .Y(_0word3_reg_31_0__20_));
AND2X2 AND2X2_4650 ( .A(core__abc_22172_new_n8283_), .B(core_v1_reg_2_), .Y(core__abc_22172_new_n8314_));
AND2X2 AND2X2_4651 ( .A(core__abc_22172_new_n8315_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8316_));
AND2X2 AND2X2_4652 ( .A(core__abc_22172_new_n7369_), .B(core__abc_22172_new_n8316_), .Y(core__abc_22172_new_n8317_));
AND2X2 AND2X2_4653 ( .A(core__abc_22172_new_n7368_), .B(core__abc_22172_new_n7815_), .Y(core__abc_22172_new_n8318_));
AND2X2 AND2X2_4654 ( .A(core__abc_22172_new_n8320_), .B(core__abc_22172_new_n8321_), .Y(core__abc_22172_new_n8322_));
AND2X2 AND2X2_4655 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n8322_), .Y(core__abc_22172_new_n8323_));
AND2X2 AND2X2_4656 ( .A(core__abc_22172_new_n8289_), .B(core__abc_22172_new_n6662_), .Y(core__abc_22172_new_n8324_));
AND2X2 AND2X2_4657 ( .A(core__abc_22172_new_n8327_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n8328_));
AND2X2 AND2X2_4658 ( .A(core__abc_22172_new_n8329_), .B(reset_n), .Y(core__0v1_reg_63_0__2_));
AND2X2 AND2X2_4659 ( .A(core__abc_22172_new_n8283_), .B(core_v1_reg_3_), .Y(core__abc_22172_new_n8331_));
AND2X2 AND2X2_466 ( .A(core_siphash_valid_reg), .B(core_siphash_word_117_), .Y(_abc_19873_new_n1691_));
AND2X2 AND2X2_4660 ( .A(core__abc_22172_new_n7831_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8333_));
AND2X2 AND2X2_4661 ( .A(core__abc_22172_new_n8332_), .B(core__abc_22172_new_n8334_), .Y(core__abc_22172_new_n8335_));
AND2X2 AND2X2_4662 ( .A(core__abc_22172_new_n8336_), .B(core__abc_22172_new_n8338_), .Y(core__abc_22172_new_n8339_));
AND2X2 AND2X2_4663 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n8339_), .Y(core__abc_22172_new_n8340_));
AND2X2 AND2X2_4664 ( .A(core__abc_22172_new_n8289_), .B(core__abc_22172_new_n6633_), .Y(core__abc_22172_new_n8341_));
AND2X2 AND2X2_4665 ( .A(core__abc_22172_new_n8343_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n8344_));
AND2X2 AND2X2_4666 ( .A(core__abc_22172_new_n8345_), .B(reset_n), .Y(core__0v1_reg_63_0__3_));
AND2X2 AND2X2_4667 ( .A(core__abc_22172_new_n8283_), .B(core_v1_reg_4_), .Y(core__abc_22172_new_n8347_));
AND2X2 AND2X2_4668 ( .A(core__abc_22172_new_n8348_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8349_));
AND2X2 AND2X2_4669 ( .A(core__abc_22172_new_n7423_), .B(core__abc_22172_new_n8349_), .Y(core__abc_22172_new_n8350_));
AND2X2 AND2X2_467 ( .A(_abc_19873_new_n1607_), .B(word3_reg_21_), .Y(_abc_19873_new_n1692_));
AND2X2 AND2X2_4670 ( .A(core__abc_22172_new_n7422_), .B(core__abc_22172_new_n7845_), .Y(core__abc_22172_new_n8351_));
AND2X2 AND2X2_4671 ( .A(core__abc_22172_new_n3214_), .B(core_key_68_), .Y(core__abc_22172_new_n8352_));
AND2X2 AND2X2_4672 ( .A(core__abc_22172_new_n8289_), .B(core__abc_22172_new_n6626_), .Y(core__abc_22172_new_n8353_));
AND2X2 AND2X2_4673 ( .A(core__abc_22172_new_n8356_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n8357_));
AND2X2 AND2X2_4674 ( .A(core__abc_22172_new_n8358_), .B(reset_n), .Y(core__0v1_reg_63_0__4_));
AND2X2 AND2X2_4675 ( .A(core__abc_22172_new_n7860_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8360_));
AND2X2 AND2X2_4676 ( .A(core__abc_22172_new_n8362_), .B(core__abc_22172_new_n8361_), .Y(core__abc_22172_new_n8363_));
AND2X2 AND2X2_4677 ( .A(core__abc_22172_new_n8364_), .B(core__abc_22172_new_n8365_), .Y(core__abc_22172_new_n8366_));
AND2X2 AND2X2_4678 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n8366_), .Y(core__abc_22172_new_n8367_));
AND2X2 AND2X2_4679 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_5_), .Y(core__abc_22172_new_n8368_));
AND2X2 AND2X2_468 ( .A(_abc_19873_new_n1693_), .B(reset_n), .Y(_0word3_reg_31_0__21_));
AND2X2 AND2X2_4680 ( .A(core__abc_22172_new_n8372_), .B(reset_n), .Y(core__abc_22172_new_n8373_));
AND2X2 AND2X2_4681 ( .A(core__abc_22172_new_n8371_), .B(core__abc_22172_new_n8373_), .Y(core__0v1_reg_63_0__5_));
AND2X2 AND2X2_4682 ( .A(core__abc_22172_new_n8283_), .B(core_v1_reg_6_), .Y(core__abc_22172_new_n8375_));
AND2X2 AND2X2_4683 ( .A(core__abc_22172_new_n7485_), .B(core__abc_22172_new_n7876_), .Y(core__abc_22172_new_n8376_));
AND2X2 AND2X2_4684 ( .A(core__abc_22172_new_n8377_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8378_));
AND2X2 AND2X2_4685 ( .A(core__abc_22172_new_n7486_), .B(core__abc_22172_new_n8378_), .Y(core__abc_22172_new_n8379_));
AND2X2 AND2X2_4686 ( .A(core__abc_22172_new_n8380_), .B(core__abc_22172_new_n8381_), .Y(core__abc_22172_new_n8382_));
AND2X2 AND2X2_4687 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n8382_), .Y(core__abc_22172_new_n8383_));
AND2X2 AND2X2_4688 ( .A(core__abc_22172_new_n8289_), .B(core__abc_22172_new_n6617_), .Y(core__abc_22172_new_n8384_));
AND2X2 AND2X2_4689 ( .A(core__abc_22172_new_n8387_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n8388_));
AND2X2 AND2X2_469 ( .A(core_siphash_valid_reg), .B(core_siphash_word_118_), .Y(_abc_19873_new_n1695_));
AND2X2 AND2X2_4690 ( .A(core__abc_22172_new_n8389_), .B(reset_n), .Y(core__0v1_reg_63_0__6_));
AND2X2 AND2X2_4691 ( .A(core__abc_22172_new_n8283_), .B(core_v1_reg_7_), .Y(core__abc_22172_new_n8391_));
AND2X2 AND2X2_4692 ( .A(core__abc_22172_new_n8393_), .B(core__abc_22172_new_n8394_), .Y(core__abc_22172_new_n8395_));
AND2X2 AND2X2_4693 ( .A(core__abc_22172_new_n8395_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8396_));
AND2X2 AND2X2_4694 ( .A(core_key_71_), .B(core_long), .Y(core__abc_22172_new_n8397_));
AND2X2 AND2X2_4695 ( .A(core__abc_22172_new_n8398_), .B(core__abc_22172_new_n8399_), .Y(core__abc_22172_new_n8400_));
AND2X2 AND2X2_4696 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n8400_), .Y(core__abc_22172_new_n8401_));
AND2X2 AND2X2_4697 ( .A(core__abc_22172_new_n8289_), .B(core__abc_22172_new_n6597_), .Y(core__abc_22172_new_n8402_));
AND2X2 AND2X2_4698 ( .A(core__abc_22172_new_n8404_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n8405_));
AND2X2 AND2X2_4699 ( .A(core__abc_22172_new_n8406_), .B(reset_n), .Y(core__0v1_reg_63_0__7_));
AND2X2 AND2X2_47 ( .A(_abc_19873_new_n936_), .B(cs), .Y(_abc_19873_new_n937_));
AND2X2 AND2X2_470 ( .A(_abc_19873_new_n1607_), .B(word3_reg_22_), .Y(_abc_19873_new_n1696_));
AND2X2 AND2X2_4700 ( .A(core__abc_22172_new_n8408_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8409_));
AND2X2 AND2X2_4701 ( .A(core__abc_22172_new_n8411_), .B(core__abc_22172_new_n8410_), .Y(core__abc_22172_new_n8412_));
AND2X2 AND2X2_4702 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_8_), .Y(core__abc_22172_new_n8413_));
AND2X2 AND2X2_4703 ( .A(core__abc_22172_new_n8417_), .B(reset_n), .Y(core__abc_22172_new_n8418_));
AND2X2 AND2X2_4704 ( .A(core__abc_22172_new_n8416_), .B(core__abc_22172_new_n8418_), .Y(core__0v1_reg_63_0__8_));
AND2X2 AND2X2_4705 ( .A(core__abc_22172_new_n8421_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8422_));
AND2X2 AND2X2_4706 ( .A(core__abc_22172_new_n8422_), .B(core__abc_22172_new_n8420_), .Y(core__abc_22172_new_n8423_));
AND2X2 AND2X2_4707 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n8424_), .Y(core__abc_22172_new_n8425_));
AND2X2 AND2X2_4708 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_9_), .Y(core__abc_22172_new_n8426_));
AND2X2 AND2X2_4709 ( .A(core__abc_22172_new_n8430_), .B(reset_n), .Y(core__abc_22172_new_n8431_));
AND2X2 AND2X2_471 ( .A(_abc_19873_new_n1697_), .B(reset_n), .Y(_0word3_reg_31_0__22_));
AND2X2 AND2X2_4710 ( .A(core__abc_22172_new_n8429_), .B(core__abc_22172_new_n8431_), .Y(core__0v1_reg_63_0__9_));
AND2X2 AND2X2_4711 ( .A(core__abc_22172_new_n8435_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8436_));
AND2X2 AND2X2_4712 ( .A(core__abc_22172_new_n8436_), .B(core__abc_22172_new_n8434_), .Y(core__abc_22172_new_n8437_));
AND2X2 AND2X2_4713 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_10_), .Y(core__abc_22172_new_n8438_));
AND2X2 AND2X2_4714 ( .A(core__abc_22172_new_n8442_), .B(reset_n), .Y(core__abc_22172_new_n8443_));
AND2X2 AND2X2_4715 ( .A(core__abc_22172_new_n8441_), .B(core__abc_22172_new_n8443_), .Y(core__0v1_reg_63_0__10_));
AND2X2 AND2X2_4716 ( .A(core__abc_22172_new_n8446_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8447_));
AND2X2 AND2X2_4717 ( .A(core__abc_22172_new_n8447_), .B(core__abc_22172_new_n8445_), .Y(core__abc_22172_new_n8448_));
AND2X2 AND2X2_4718 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n8449_), .Y(core__abc_22172_new_n8450_));
AND2X2 AND2X2_4719 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_11_), .Y(core__abc_22172_new_n8451_));
AND2X2 AND2X2_472 ( .A(core_siphash_valid_reg), .B(core_siphash_word_119_), .Y(_abc_19873_new_n1699_));
AND2X2 AND2X2_4720 ( .A(core__abc_22172_new_n8455_), .B(reset_n), .Y(core__abc_22172_new_n8456_));
AND2X2 AND2X2_4721 ( .A(core__abc_22172_new_n8454_), .B(core__abc_22172_new_n8456_), .Y(core__0v1_reg_63_0__11_));
AND2X2 AND2X2_4722 ( .A(core__abc_22172_new_n8460_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8461_));
AND2X2 AND2X2_4723 ( .A(core__abc_22172_new_n8461_), .B(core__abc_22172_new_n8459_), .Y(core__abc_22172_new_n8462_));
AND2X2 AND2X2_4724 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_12_), .Y(core__abc_22172_new_n8463_));
AND2X2 AND2X2_4725 ( .A(core__abc_22172_new_n8467_), .B(reset_n), .Y(core__abc_22172_new_n8468_));
AND2X2 AND2X2_4726 ( .A(core__abc_22172_new_n8466_), .B(core__abc_22172_new_n8468_), .Y(core__0v1_reg_63_0__12_));
AND2X2 AND2X2_4727 ( .A(core__abc_22172_new_n8472_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8473_));
AND2X2 AND2X2_4728 ( .A(core__abc_22172_new_n8473_), .B(core__abc_22172_new_n8470_), .Y(core__abc_22172_new_n8474_));
AND2X2 AND2X2_4729 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_13_), .Y(core__abc_22172_new_n8475_));
AND2X2 AND2X2_473 ( .A(_abc_19873_new_n1607_), .B(word3_reg_23_), .Y(_abc_19873_new_n1700_));
AND2X2 AND2X2_4730 ( .A(core__abc_22172_new_n8479_), .B(reset_n), .Y(core__abc_22172_new_n8480_));
AND2X2 AND2X2_4731 ( .A(core__abc_22172_new_n8478_), .B(core__abc_22172_new_n8480_), .Y(core__0v1_reg_63_0__13_));
AND2X2 AND2X2_4732 ( .A(core__abc_22172_new_n8483_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8484_));
AND2X2 AND2X2_4733 ( .A(core__abc_22172_new_n8484_), .B(core__abc_22172_new_n8482_), .Y(core__abc_22172_new_n8485_));
AND2X2 AND2X2_4734 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_14_), .Y(core__abc_22172_new_n8486_));
AND2X2 AND2X2_4735 ( .A(core__abc_22172_new_n8490_), .B(reset_n), .Y(core__abc_22172_new_n8491_));
AND2X2 AND2X2_4736 ( .A(core__abc_22172_new_n8489_), .B(core__abc_22172_new_n8491_), .Y(core__0v1_reg_63_0__14_));
AND2X2 AND2X2_4737 ( .A(core__abc_22172_new_n8494_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8495_));
AND2X2 AND2X2_4738 ( .A(core__abc_22172_new_n8495_), .B(core__abc_22172_new_n8493_), .Y(core__abc_22172_new_n8496_));
AND2X2 AND2X2_4739 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_15_), .Y(core__abc_22172_new_n8497_));
AND2X2 AND2X2_474 ( .A(_abc_19873_new_n1701_), .B(reset_n), .Y(_0word3_reg_31_0__23_));
AND2X2 AND2X2_4740 ( .A(core__abc_22172_new_n8501_), .B(reset_n), .Y(core__abc_22172_new_n8502_));
AND2X2 AND2X2_4741 ( .A(core__abc_22172_new_n8500_), .B(core__abc_22172_new_n8502_), .Y(core__0v1_reg_63_0__15_));
AND2X2 AND2X2_4742 ( .A(core__abc_22172_new_n8505_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8506_));
AND2X2 AND2X2_4743 ( .A(core__abc_22172_new_n8506_), .B(core__abc_22172_new_n8504_), .Y(core__abc_22172_new_n8507_));
AND2X2 AND2X2_4744 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_16_), .Y(core__abc_22172_new_n8508_));
AND2X2 AND2X2_4745 ( .A(core__abc_22172_new_n8512_), .B(reset_n), .Y(core__abc_22172_new_n8513_));
AND2X2 AND2X2_4746 ( .A(core__abc_22172_new_n8511_), .B(core__abc_22172_new_n8513_), .Y(core__0v1_reg_63_0__16_));
AND2X2 AND2X2_4747 ( .A(core__abc_22172_new_n8517_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8518_));
AND2X2 AND2X2_4748 ( .A(core__abc_22172_new_n8518_), .B(core__abc_22172_new_n8516_), .Y(core__abc_22172_new_n8519_));
AND2X2 AND2X2_4749 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_17_), .Y(core__abc_22172_new_n8520_));
AND2X2 AND2X2_475 ( .A(core_siphash_valid_reg), .B(core_siphash_word_120_), .Y(_abc_19873_new_n1703_));
AND2X2 AND2X2_4750 ( .A(core__abc_22172_new_n8524_), .B(reset_n), .Y(core__abc_22172_new_n8525_));
AND2X2 AND2X2_4751 ( .A(core__abc_22172_new_n8523_), .B(core__abc_22172_new_n8525_), .Y(core__0v1_reg_63_0__17_));
AND2X2 AND2X2_4752 ( .A(core__abc_22172_new_n8529_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8530_));
AND2X2 AND2X2_4753 ( .A(core__abc_22172_new_n8530_), .B(core__abc_22172_new_n8528_), .Y(core__abc_22172_new_n8531_));
AND2X2 AND2X2_4754 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_18_), .Y(core__abc_22172_new_n8532_));
AND2X2 AND2X2_4755 ( .A(core__abc_22172_new_n8536_), .B(reset_n), .Y(core__abc_22172_new_n8537_));
AND2X2 AND2X2_4756 ( .A(core__abc_22172_new_n8535_), .B(core__abc_22172_new_n8537_), .Y(core__0v1_reg_63_0__18_));
AND2X2 AND2X2_4757 ( .A(core__abc_22172_new_n8541_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8542_));
AND2X2 AND2X2_4758 ( .A(core__abc_22172_new_n8542_), .B(core__abc_22172_new_n8540_), .Y(core__abc_22172_new_n8543_));
AND2X2 AND2X2_4759 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_19_), .Y(core__abc_22172_new_n8544_));
AND2X2 AND2X2_476 ( .A(_abc_19873_new_n1607_), .B(word3_reg_24_), .Y(_abc_19873_new_n1704_));
AND2X2 AND2X2_4760 ( .A(core__abc_22172_new_n8548_), .B(reset_n), .Y(core__abc_22172_new_n8549_));
AND2X2 AND2X2_4761 ( .A(core__abc_22172_new_n8547_), .B(core__abc_22172_new_n8549_), .Y(core__0v1_reg_63_0__19_));
AND2X2 AND2X2_4762 ( .A(core__abc_22172_new_n8552_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8553_));
AND2X2 AND2X2_4763 ( .A(core__abc_22172_new_n8553_), .B(core__abc_22172_new_n8551_), .Y(core__abc_22172_new_n8554_));
AND2X2 AND2X2_4764 ( .A(core__abc_22172_new_n3214_), .B(core_key_84_), .Y(core__abc_22172_new_n8555_));
AND2X2 AND2X2_4765 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_20_), .Y(core__abc_22172_new_n8556_));
AND2X2 AND2X2_4766 ( .A(core__abc_22172_new_n8560_), .B(reset_n), .Y(core__abc_22172_new_n8561_));
AND2X2 AND2X2_4767 ( .A(core__abc_22172_new_n8559_), .B(core__abc_22172_new_n8561_), .Y(core__0v1_reg_63_0__20_));
AND2X2 AND2X2_4768 ( .A(core__abc_22172_new_n8564_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8565_));
AND2X2 AND2X2_4769 ( .A(core__abc_22172_new_n8565_), .B(core__abc_22172_new_n8563_), .Y(core__abc_22172_new_n8566_));
AND2X2 AND2X2_477 ( .A(_abc_19873_new_n1705_), .B(reset_n), .Y(_0word3_reg_31_0__24_));
AND2X2 AND2X2_4770 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_21_), .Y(core__abc_22172_new_n8567_));
AND2X2 AND2X2_4771 ( .A(core__abc_22172_new_n8571_), .B(reset_n), .Y(core__abc_22172_new_n8572_));
AND2X2 AND2X2_4772 ( .A(core__abc_22172_new_n8570_), .B(core__abc_22172_new_n8572_), .Y(core__0v1_reg_63_0__21_));
AND2X2 AND2X2_4773 ( .A(core__abc_22172_new_n8576_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8577_));
AND2X2 AND2X2_4774 ( .A(core__abc_22172_new_n8577_), .B(core__abc_22172_new_n8575_), .Y(core__abc_22172_new_n8578_));
AND2X2 AND2X2_4775 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_22_), .Y(core__abc_22172_new_n8579_));
AND2X2 AND2X2_4776 ( .A(core__abc_22172_new_n8583_), .B(reset_n), .Y(core__abc_22172_new_n8584_));
AND2X2 AND2X2_4777 ( .A(core__abc_22172_new_n8582_), .B(core__abc_22172_new_n8584_), .Y(core__0v1_reg_63_0__22_));
AND2X2 AND2X2_4778 ( .A(core__abc_22172_new_n8587_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8588_));
AND2X2 AND2X2_4779 ( .A(core__abc_22172_new_n8588_), .B(core__abc_22172_new_n8586_), .Y(core__abc_22172_new_n8589_));
AND2X2 AND2X2_478 ( .A(core_siphash_valid_reg), .B(core_siphash_word_121_), .Y(_abc_19873_new_n1707_));
AND2X2 AND2X2_4780 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_23_), .Y(core__abc_22172_new_n8590_));
AND2X2 AND2X2_4781 ( .A(core__abc_22172_new_n8594_), .B(reset_n), .Y(core__abc_22172_new_n8595_));
AND2X2 AND2X2_4782 ( .A(core__abc_22172_new_n8593_), .B(core__abc_22172_new_n8595_), .Y(core__0v1_reg_63_0__23_));
AND2X2 AND2X2_4783 ( .A(core__abc_22172_new_n8599_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8600_));
AND2X2 AND2X2_4784 ( .A(core__abc_22172_new_n8600_), .B(core__abc_22172_new_n8598_), .Y(core__abc_22172_new_n8601_));
AND2X2 AND2X2_4785 ( .A(core__abc_22172_new_n3214_), .B(core_key_88_), .Y(core__abc_22172_new_n8602_));
AND2X2 AND2X2_4786 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_24_), .Y(core__abc_22172_new_n8603_));
AND2X2 AND2X2_4787 ( .A(core__abc_22172_new_n8607_), .B(reset_n), .Y(core__abc_22172_new_n8608_));
AND2X2 AND2X2_4788 ( .A(core__abc_22172_new_n8606_), .B(core__abc_22172_new_n8608_), .Y(core__0v1_reg_63_0__24_));
AND2X2 AND2X2_4789 ( .A(core__abc_22172_new_n8612_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8613_));
AND2X2 AND2X2_479 ( .A(_abc_19873_new_n1607_), .B(word3_reg_25_), .Y(_abc_19873_new_n1708_));
AND2X2 AND2X2_4790 ( .A(core__abc_22172_new_n8613_), .B(core__abc_22172_new_n8611_), .Y(core__abc_22172_new_n8614_));
AND2X2 AND2X2_4791 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n8615_), .Y(core__abc_22172_new_n8616_));
AND2X2 AND2X2_4792 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_25_), .Y(core__abc_22172_new_n8617_));
AND2X2 AND2X2_4793 ( .A(core__abc_22172_new_n8621_), .B(reset_n), .Y(core__abc_22172_new_n8622_));
AND2X2 AND2X2_4794 ( .A(core__abc_22172_new_n8620_), .B(core__abc_22172_new_n8622_), .Y(core__0v1_reg_63_0__25_));
AND2X2 AND2X2_4795 ( .A(core__abc_22172_new_n8627_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8628_));
AND2X2 AND2X2_4796 ( .A(core__abc_22172_new_n8628_), .B(core__abc_22172_new_n8625_), .Y(core__abc_22172_new_n8629_));
AND2X2 AND2X2_4797 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n8630_), .Y(core__abc_22172_new_n8631_));
AND2X2 AND2X2_4798 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_26_), .Y(core__abc_22172_new_n8632_));
AND2X2 AND2X2_4799 ( .A(core__abc_22172_new_n8636_), .B(reset_n), .Y(core__abc_22172_new_n8637_));
AND2X2 AND2X2_48 ( .A(_abc_19873_new_n935_), .B(_abc_19873_new_n937_), .Y(\read_data[0] ));
AND2X2 AND2X2_480 ( .A(_abc_19873_new_n1709_), .B(reset_n), .Y(_0word3_reg_31_0__25_));
AND2X2 AND2X2_4800 ( .A(core__abc_22172_new_n8635_), .B(core__abc_22172_new_n8637_), .Y(core__0v1_reg_63_0__26_));
AND2X2 AND2X2_4801 ( .A(core__abc_22172_new_n8641_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8642_));
AND2X2 AND2X2_4802 ( .A(core__abc_22172_new_n8642_), .B(core__abc_22172_new_n8640_), .Y(core__abc_22172_new_n8643_));
AND2X2 AND2X2_4803 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_27_), .Y(core__abc_22172_new_n8644_));
AND2X2 AND2X2_4804 ( .A(core__abc_22172_new_n8648_), .B(reset_n), .Y(core__abc_22172_new_n8649_));
AND2X2 AND2X2_4805 ( .A(core__abc_22172_new_n8647_), .B(core__abc_22172_new_n8649_), .Y(core__0v1_reg_63_0__27_));
AND2X2 AND2X2_4806 ( .A(core__abc_22172_new_n8652_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8653_));
AND2X2 AND2X2_4807 ( .A(core__abc_22172_new_n8653_), .B(core__abc_22172_new_n8651_), .Y(core__abc_22172_new_n8654_));
AND2X2 AND2X2_4808 ( .A(core__abc_22172_new_n3214_), .B(core_key_92_), .Y(core__abc_22172_new_n8655_));
AND2X2 AND2X2_4809 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_28_), .Y(core__abc_22172_new_n8656_));
AND2X2 AND2X2_481 ( .A(core_siphash_valid_reg), .B(core_siphash_word_122_), .Y(_abc_19873_new_n1711_));
AND2X2 AND2X2_4810 ( .A(core__abc_22172_new_n8660_), .B(reset_n), .Y(core__abc_22172_new_n8661_));
AND2X2 AND2X2_4811 ( .A(core__abc_22172_new_n8659_), .B(core__abc_22172_new_n8661_), .Y(core__0v1_reg_63_0__28_));
AND2X2 AND2X2_4812 ( .A(core__abc_22172_new_n8664_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8665_));
AND2X2 AND2X2_4813 ( .A(core__abc_22172_new_n8665_), .B(core__abc_22172_new_n8663_), .Y(core__abc_22172_new_n8666_));
AND2X2 AND2X2_4814 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_29_), .Y(core__abc_22172_new_n8667_));
AND2X2 AND2X2_4815 ( .A(core__abc_22172_new_n8671_), .B(reset_n), .Y(core__abc_22172_new_n8672_));
AND2X2 AND2X2_4816 ( .A(core__abc_22172_new_n8670_), .B(core__abc_22172_new_n8672_), .Y(core__0v1_reg_63_0__29_));
AND2X2 AND2X2_4817 ( .A(core__abc_22172_new_n8676_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8677_));
AND2X2 AND2X2_4818 ( .A(core__abc_22172_new_n8677_), .B(core__abc_22172_new_n8675_), .Y(core__abc_22172_new_n8678_));
AND2X2 AND2X2_4819 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_30_), .Y(core__abc_22172_new_n8679_));
AND2X2 AND2X2_482 ( .A(_abc_19873_new_n1607_), .B(word3_reg_26_), .Y(_abc_19873_new_n1712_));
AND2X2 AND2X2_4820 ( .A(core__abc_22172_new_n8683_), .B(reset_n), .Y(core__abc_22172_new_n8684_));
AND2X2 AND2X2_4821 ( .A(core__abc_22172_new_n8682_), .B(core__abc_22172_new_n8684_), .Y(core__0v1_reg_63_0__30_));
AND2X2 AND2X2_4822 ( .A(core__abc_22172_new_n8687_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8688_));
AND2X2 AND2X2_4823 ( .A(core__abc_22172_new_n8688_), .B(core__abc_22172_new_n8686_), .Y(core__abc_22172_new_n8689_));
AND2X2 AND2X2_4824 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_31_), .Y(core__abc_22172_new_n8690_));
AND2X2 AND2X2_4825 ( .A(core__abc_22172_new_n8694_), .B(reset_n), .Y(core__abc_22172_new_n8695_));
AND2X2 AND2X2_4826 ( .A(core__abc_22172_new_n8693_), .B(core__abc_22172_new_n8695_), .Y(core__0v1_reg_63_0__31_));
AND2X2 AND2X2_4827 ( .A(core__abc_22172_new_n8698_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8699_));
AND2X2 AND2X2_4828 ( .A(core__abc_22172_new_n8699_), .B(core__abc_22172_new_n8697_), .Y(core__abc_22172_new_n8700_));
AND2X2 AND2X2_4829 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n8701_), .Y(core__abc_22172_new_n8702_));
AND2X2 AND2X2_483 ( .A(_abc_19873_new_n1713_), .B(reset_n), .Y(_0word3_reg_31_0__26_));
AND2X2 AND2X2_4830 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_32_), .Y(core__abc_22172_new_n8703_));
AND2X2 AND2X2_4831 ( .A(core__abc_22172_new_n8707_), .B(reset_n), .Y(core__abc_22172_new_n8708_));
AND2X2 AND2X2_4832 ( .A(core__abc_22172_new_n8706_), .B(core__abc_22172_new_n8708_), .Y(core__0v1_reg_63_0__32_));
AND2X2 AND2X2_4833 ( .A(core__abc_22172_new_n8711_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8712_));
AND2X2 AND2X2_4834 ( .A(core__abc_22172_new_n8712_), .B(core__abc_22172_new_n8710_), .Y(core__abc_22172_new_n8713_));
AND2X2 AND2X2_4835 ( .A(core__abc_22172_new_n3214_), .B(core_key_97_), .Y(core__abc_22172_new_n8714_));
AND2X2 AND2X2_4836 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_33_), .Y(core__abc_22172_new_n8715_));
AND2X2 AND2X2_4837 ( .A(core__abc_22172_new_n8719_), .B(reset_n), .Y(core__abc_22172_new_n8720_));
AND2X2 AND2X2_4838 ( .A(core__abc_22172_new_n8718_), .B(core__abc_22172_new_n8720_), .Y(core__0v1_reg_63_0__33_));
AND2X2 AND2X2_4839 ( .A(core__abc_22172_new_n8724_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8725_));
AND2X2 AND2X2_484 ( .A(core_siphash_valid_reg), .B(core_siphash_word_123_), .Y(_abc_19873_new_n1715_));
AND2X2 AND2X2_4840 ( .A(core__abc_22172_new_n8725_), .B(core__abc_22172_new_n8723_), .Y(core__abc_22172_new_n8726_));
AND2X2 AND2X2_4841 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_34_), .Y(core__abc_22172_new_n8727_));
AND2X2 AND2X2_4842 ( .A(core__abc_22172_new_n8731_), .B(reset_n), .Y(core__abc_22172_new_n8732_));
AND2X2 AND2X2_4843 ( .A(core__abc_22172_new_n8730_), .B(core__abc_22172_new_n8732_), .Y(core__0v1_reg_63_0__34_));
AND2X2 AND2X2_4844 ( .A(core__abc_22172_new_n8736_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8737_));
AND2X2 AND2X2_4845 ( .A(core__abc_22172_new_n8737_), .B(core__abc_22172_new_n8735_), .Y(core__abc_22172_new_n8738_));
AND2X2 AND2X2_4846 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_35_), .Y(core__abc_22172_new_n8739_));
AND2X2 AND2X2_4847 ( .A(core__abc_22172_new_n8743_), .B(reset_n), .Y(core__abc_22172_new_n8744_));
AND2X2 AND2X2_4848 ( .A(core__abc_22172_new_n8742_), .B(core__abc_22172_new_n8744_), .Y(core__0v1_reg_63_0__35_));
AND2X2 AND2X2_4849 ( .A(core__abc_22172_new_n8747_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8748_));
AND2X2 AND2X2_485 ( .A(_abc_19873_new_n1607_), .B(word3_reg_27_), .Y(_abc_19873_new_n1716_));
AND2X2 AND2X2_4850 ( .A(core__abc_22172_new_n8748_), .B(core__abc_22172_new_n8746_), .Y(core__abc_22172_new_n8749_));
AND2X2 AND2X2_4851 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_36_), .Y(core__abc_22172_new_n8750_));
AND2X2 AND2X2_4852 ( .A(core__abc_22172_new_n8754_), .B(reset_n), .Y(core__abc_22172_new_n8755_));
AND2X2 AND2X2_4853 ( .A(core__abc_22172_new_n8753_), .B(core__abc_22172_new_n8755_), .Y(core__0v1_reg_63_0__36_));
AND2X2 AND2X2_4854 ( .A(core__abc_22172_new_n8758_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8759_));
AND2X2 AND2X2_4855 ( .A(core__abc_22172_new_n8759_), .B(core__abc_22172_new_n8757_), .Y(core__abc_22172_new_n8760_));
AND2X2 AND2X2_4856 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_37_), .Y(core__abc_22172_new_n8761_));
AND2X2 AND2X2_4857 ( .A(core__abc_22172_new_n8765_), .B(reset_n), .Y(core__abc_22172_new_n8766_));
AND2X2 AND2X2_4858 ( .A(core__abc_22172_new_n8764_), .B(core__abc_22172_new_n8766_), .Y(core__0v1_reg_63_0__37_));
AND2X2 AND2X2_4859 ( .A(core__abc_22172_new_n8770_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8771_));
AND2X2 AND2X2_486 ( .A(_abc_19873_new_n1717_), .B(reset_n), .Y(_0word3_reg_31_0__27_));
AND2X2 AND2X2_4860 ( .A(core__abc_22172_new_n8771_), .B(core__abc_22172_new_n8768_), .Y(core__abc_22172_new_n8772_));
AND2X2 AND2X2_4861 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_38_), .Y(core__abc_22172_new_n8773_));
AND2X2 AND2X2_4862 ( .A(core__abc_22172_new_n8777_), .B(reset_n), .Y(core__abc_22172_new_n8778_));
AND2X2 AND2X2_4863 ( .A(core__abc_22172_new_n8776_), .B(core__abc_22172_new_n8778_), .Y(core__0v1_reg_63_0__38_));
AND2X2 AND2X2_4864 ( .A(core__abc_22172_new_n8782_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8783_));
AND2X2 AND2X2_4865 ( .A(core__abc_22172_new_n8783_), .B(core__abc_22172_new_n8781_), .Y(core__abc_22172_new_n8784_));
AND2X2 AND2X2_4866 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_39_), .Y(core__abc_22172_new_n8785_));
AND2X2 AND2X2_4867 ( .A(core__abc_22172_new_n8789_), .B(reset_n), .Y(core__abc_22172_new_n8790_));
AND2X2 AND2X2_4868 ( .A(core__abc_22172_new_n8788_), .B(core__abc_22172_new_n8790_), .Y(core__0v1_reg_63_0__39_));
AND2X2 AND2X2_4869 ( .A(core__abc_22172_new_n8793_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8794_));
AND2X2 AND2X2_487 ( .A(core_siphash_valid_reg), .B(core_siphash_word_124_), .Y(_abc_19873_new_n1719_));
AND2X2 AND2X2_4870 ( .A(core__abc_22172_new_n8794_), .B(core__abc_22172_new_n8792_), .Y(core__abc_22172_new_n8795_));
AND2X2 AND2X2_4871 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_40_), .Y(core__abc_22172_new_n8796_));
AND2X2 AND2X2_4872 ( .A(core__abc_22172_new_n8800_), .B(reset_n), .Y(core__abc_22172_new_n8801_));
AND2X2 AND2X2_4873 ( .A(core__abc_22172_new_n8799_), .B(core__abc_22172_new_n8801_), .Y(core__0v1_reg_63_0__40_));
AND2X2 AND2X2_4874 ( .A(core__abc_22172_new_n8804_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8805_));
AND2X2 AND2X2_4875 ( .A(core__abc_22172_new_n8805_), .B(core__abc_22172_new_n8803_), .Y(core__abc_22172_new_n8806_));
AND2X2 AND2X2_4876 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n8807_), .Y(core__abc_22172_new_n8808_));
AND2X2 AND2X2_4877 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_41_), .Y(core__abc_22172_new_n8809_));
AND2X2 AND2X2_4878 ( .A(core__abc_22172_new_n8813_), .B(reset_n), .Y(core__abc_22172_new_n8814_));
AND2X2 AND2X2_4879 ( .A(core__abc_22172_new_n8812_), .B(core__abc_22172_new_n8814_), .Y(core__0v1_reg_63_0__41_));
AND2X2 AND2X2_488 ( .A(_abc_19873_new_n1607_), .B(word3_reg_28_), .Y(_abc_19873_new_n1720_));
AND2X2 AND2X2_4880 ( .A(core__abc_22172_new_n8818_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8819_));
AND2X2 AND2X2_4881 ( .A(core__abc_22172_new_n8819_), .B(core__abc_22172_new_n8817_), .Y(core__abc_22172_new_n8820_));
AND2X2 AND2X2_4882 ( .A(core__abc_22172_new_n3214_), .B(core_key_106_), .Y(core__abc_22172_new_n8821_));
AND2X2 AND2X2_4883 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_42_), .Y(core__abc_22172_new_n8822_));
AND2X2 AND2X2_4884 ( .A(core__abc_22172_new_n8826_), .B(reset_n), .Y(core__abc_22172_new_n8827_));
AND2X2 AND2X2_4885 ( .A(core__abc_22172_new_n8825_), .B(core__abc_22172_new_n8827_), .Y(core__0v1_reg_63_0__42_));
AND2X2 AND2X2_4886 ( .A(core__abc_22172_new_n8831_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8832_));
AND2X2 AND2X2_4887 ( .A(core__abc_22172_new_n8832_), .B(core__abc_22172_new_n8830_), .Y(core__abc_22172_new_n8833_));
AND2X2 AND2X2_4888 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_43_), .Y(core__abc_22172_new_n8834_));
AND2X2 AND2X2_4889 ( .A(core__abc_22172_new_n8838_), .B(reset_n), .Y(core__abc_22172_new_n8839_));
AND2X2 AND2X2_489 ( .A(_abc_19873_new_n1721_), .B(reset_n), .Y(_0word3_reg_31_0__28_));
AND2X2 AND2X2_4890 ( .A(core__abc_22172_new_n8837_), .B(core__abc_22172_new_n8839_), .Y(core__0v1_reg_63_0__43_));
AND2X2 AND2X2_4891 ( .A(core__abc_22172_new_n8842_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8843_));
AND2X2 AND2X2_4892 ( .A(core__abc_22172_new_n8843_), .B(core__abc_22172_new_n8841_), .Y(core__abc_22172_new_n8844_));
AND2X2 AND2X2_4893 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n8845_), .Y(core__abc_22172_new_n8846_));
AND2X2 AND2X2_4894 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_44_), .Y(core__abc_22172_new_n8847_));
AND2X2 AND2X2_4895 ( .A(core__abc_22172_new_n8851_), .B(reset_n), .Y(core__abc_22172_new_n8852_));
AND2X2 AND2X2_4896 ( .A(core__abc_22172_new_n8850_), .B(core__abc_22172_new_n8852_), .Y(core__0v1_reg_63_0__44_));
AND2X2 AND2X2_4897 ( .A(core__abc_22172_new_n8856_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8857_));
AND2X2 AND2X2_4898 ( .A(core__abc_22172_new_n8857_), .B(core__abc_22172_new_n8855_), .Y(core__abc_22172_new_n8858_));
AND2X2 AND2X2_4899 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_45_), .Y(core__abc_22172_new_n8859_));
AND2X2 AND2X2_49 ( .A(_abc_19873_new_n881_), .B(core_key_97_), .Y(_abc_19873_new_n939_));
AND2X2 AND2X2_490 ( .A(core_siphash_valid_reg), .B(core_siphash_word_125_), .Y(_abc_19873_new_n1723_));
AND2X2 AND2X2_4900 ( .A(core__abc_22172_new_n8863_), .B(reset_n), .Y(core__abc_22172_new_n8864_));
AND2X2 AND2X2_4901 ( .A(core__abc_22172_new_n8862_), .B(core__abc_22172_new_n8864_), .Y(core__0v1_reg_63_0__45_));
AND2X2 AND2X2_4902 ( .A(core__abc_22172_new_n8867_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8868_));
AND2X2 AND2X2_4903 ( .A(core__abc_22172_new_n8868_), .B(core__abc_22172_new_n8866_), .Y(core__abc_22172_new_n8869_));
AND2X2 AND2X2_4904 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_46_), .Y(core__abc_22172_new_n8870_));
AND2X2 AND2X2_4905 ( .A(core__abc_22172_new_n8874_), .B(reset_n), .Y(core__abc_22172_new_n8875_));
AND2X2 AND2X2_4906 ( .A(core__abc_22172_new_n8873_), .B(core__abc_22172_new_n8875_), .Y(core__0v1_reg_63_0__46_));
AND2X2 AND2X2_4907 ( .A(core__abc_22172_new_n8878_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8879_));
AND2X2 AND2X2_4908 ( .A(core__abc_22172_new_n8879_), .B(core__abc_22172_new_n8877_), .Y(core__abc_22172_new_n8880_));
AND2X2 AND2X2_4909 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_47_), .Y(core__abc_22172_new_n8881_));
AND2X2 AND2X2_491 ( .A(_abc_19873_new_n1607_), .B(word3_reg_29_), .Y(_abc_19873_new_n1724_));
AND2X2 AND2X2_4910 ( .A(core__abc_22172_new_n8885_), .B(reset_n), .Y(core__abc_22172_new_n8886_));
AND2X2 AND2X2_4911 ( .A(core__abc_22172_new_n8884_), .B(core__abc_22172_new_n8886_), .Y(core__0v1_reg_63_0__47_));
AND2X2 AND2X2_4912 ( .A(core__abc_22172_new_n8890_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8891_));
AND2X2 AND2X2_4913 ( .A(core__abc_22172_new_n8891_), .B(core__abc_22172_new_n8888_), .Y(core__abc_22172_new_n8892_));
AND2X2 AND2X2_4914 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_48_), .Y(core__abc_22172_new_n8893_));
AND2X2 AND2X2_4915 ( .A(core__abc_22172_new_n8897_), .B(reset_n), .Y(core__abc_22172_new_n8898_));
AND2X2 AND2X2_4916 ( .A(core__abc_22172_new_n8896_), .B(core__abc_22172_new_n8898_), .Y(core__0v1_reg_63_0__48_));
AND2X2 AND2X2_4917 ( .A(core__abc_22172_new_n8901_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8902_));
AND2X2 AND2X2_4918 ( .A(core__abc_22172_new_n8902_), .B(core__abc_22172_new_n8900_), .Y(core__abc_22172_new_n8903_));
AND2X2 AND2X2_4919 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n8904_), .Y(core__abc_22172_new_n8905_));
AND2X2 AND2X2_492 ( .A(_abc_19873_new_n1725_), .B(reset_n), .Y(_0word3_reg_31_0__29_));
AND2X2 AND2X2_4920 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_49_), .Y(core__abc_22172_new_n8906_));
AND2X2 AND2X2_4921 ( .A(core__abc_22172_new_n8910_), .B(reset_n), .Y(core__abc_22172_new_n8911_));
AND2X2 AND2X2_4922 ( .A(core__abc_22172_new_n8909_), .B(core__abc_22172_new_n8911_), .Y(core__0v1_reg_63_0__49_));
AND2X2 AND2X2_4923 ( .A(core__abc_22172_new_n8914_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8915_));
AND2X2 AND2X2_4924 ( .A(core__abc_22172_new_n8915_), .B(core__abc_22172_new_n8913_), .Y(core__abc_22172_new_n8916_));
AND2X2 AND2X2_4925 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_50_), .Y(core__abc_22172_new_n8917_));
AND2X2 AND2X2_4926 ( .A(core__abc_22172_new_n8921_), .B(reset_n), .Y(core__abc_22172_new_n8922_));
AND2X2 AND2X2_4927 ( .A(core__abc_22172_new_n8920_), .B(core__abc_22172_new_n8922_), .Y(core__0v1_reg_63_0__50_));
AND2X2 AND2X2_4928 ( .A(core__abc_22172_new_n8926_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8927_));
AND2X2 AND2X2_4929 ( .A(core__abc_22172_new_n8927_), .B(core__abc_22172_new_n8925_), .Y(core__abc_22172_new_n8928_));
AND2X2 AND2X2_493 ( .A(core_siphash_valid_reg), .B(core_siphash_word_126_), .Y(_abc_19873_new_n1727_));
AND2X2 AND2X2_4930 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n8929_), .Y(core__abc_22172_new_n8930_));
AND2X2 AND2X2_4931 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_51_), .Y(core__abc_22172_new_n8931_));
AND2X2 AND2X2_4932 ( .A(core__abc_22172_new_n8935_), .B(reset_n), .Y(core__abc_22172_new_n8936_));
AND2X2 AND2X2_4933 ( .A(core__abc_22172_new_n8934_), .B(core__abc_22172_new_n8936_), .Y(core__0v1_reg_63_0__51_));
AND2X2 AND2X2_4934 ( .A(core__abc_22172_new_n8939_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8940_));
AND2X2 AND2X2_4935 ( .A(core__abc_22172_new_n8940_), .B(core__abc_22172_new_n8938_), .Y(core__abc_22172_new_n8941_));
AND2X2 AND2X2_4936 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_52_), .Y(core__abc_22172_new_n8942_));
AND2X2 AND2X2_4937 ( .A(core__abc_22172_new_n8946_), .B(reset_n), .Y(core__abc_22172_new_n8947_));
AND2X2 AND2X2_4938 ( .A(core__abc_22172_new_n8945_), .B(core__abc_22172_new_n8947_), .Y(core__0v1_reg_63_0__52_));
AND2X2 AND2X2_4939 ( .A(core__abc_22172_new_n8951_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8952_));
AND2X2 AND2X2_494 ( .A(_abc_19873_new_n1607_), .B(word3_reg_30_), .Y(_abc_19873_new_n1728_));
AND2X2 AND2X2_4940 ( .A(core__abc_22172_new_n8952_), .B(core__abc_22172_new_n8950_), .Y(core__abc_22172_new_n8953_));
AND2X2 AND2X2_4941 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_53_), .Y(core__abc_22172_new_n8954_));
AND2X2 AND2X2_4942 ( .A(core__abc_22172_new_n8958_), .B(reset_n), .Y(core__abc_22172_new_n8959_));
AND2X2 AND2X2_4943 ( .A(core__abc_22172_new_n8957_), .B(core__abc_22172_new_n8959_), .Y(core__0v1_reg_63_0__53_));
AND2X2 AND2X2_4944 ( .A(core__abc_22172_new_n8963_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8964_));
AND2X2 AND2X2_4945 ( .A(core__abc_22172_new_n8964_), .B(core__abc_22172_new_n8961_), .Y(core__abc_22172_new_n8965_));
AND2X2 AND2X2_4946 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_54_), .Y(core__abc_22172_new_n8966_));
AND2X2 AND2X2_4947 ( .A(core__abc_22172_new_n8970_), .B(reset_n), .Y(core__abc_22172_new_n8971_));
AND2X2 AND2X2_4948 ( .A(core__abc_22172_new_n8969_), .B(core__abc_22172_new_n8971_), .Y(core__0v1_reg_63_0__54_));
AND2X2 AND2X2_4949 ( .A(core__abc_22172_new_n8974_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8975_));
AND2X2 AND2X2_495 ( .A(_abc_19873_new_n1729_), .B(reset_n), .Y(_0word3_reg_31_0__30_));
AND2X2 AND2X2_4950 ( .A(core__abc_22172_new_n8975_), .B(core__abc_22172_new_n8973_), .Y(core__abc_22172_new_n8976_));
AND2X2 AND2X2_4951 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_55_), .Y(core__abc_22172_new_n8977_));
AND2X2 AND2X2_4952 ( .A(core__abc_22172_new_n8981_), .B(reset_n), .Y(core__abc_22172_new_n8982_));
AND2X2 AND2X2_4953 ( .A(core__abc_22172_new_n8980_), .B(core__abc_22172_new_n8982_), .Y(core__0v1_reg_63_0__55_));
AND2X2 AND2X2_4954 ( .A(core__abc_22172_new_n8985_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8986_));
AND2X2 AND2X2_4955 ( .A(core__abc_22172_new_n8986_), .B(core__abc_22172_new_n8984_), .Y(core__abc_22172_new_n8987_));
AND2X2 AND2X2_4956 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_56_), .Y(core__abc_22172_new_n8988_));
AND2X2 AND2X2_4957 ( .A(core__abc_22172_new_n8992_), .B(reset_n), .Y(core__abc_22172_new_n8993_));
AND2X2 AND2X2_4958 ( .A(core__abc_22172_new_n8991_), .B(core__abc_22172_new_n8993_), .Y(core__0v1_reg_63_0__56_));
AND2X2 AND2X2_4959 ( .A(core__abc_22172_new_n8997_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n8998_));
AND2X2 AND2X2_496 ( .A(core_siphash_valid_reg), .B(core_siphash_word_127_), .Y(_abc_19873_new_n1731_));
AND2X2 AND2X2_4960 ( .A(core__abc_22172_new_n8998_), .B(core__abc_22172_new_n8996_), .Y(core__abc_22172_new_n8999_));
AND2X2 AND2X2_4961 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_57_), .Y(core__abc_22172_new_n9000_));
AND2X2 AND2X2_4962 ( .A(core__abc_22172_new_n9004_), .B(reset_n), .Y(core__abc_22172_new_n9005_));
AND2X2 AND2X2_4963 ( .A(core__abc_22172_new_n9003_), .B(core__abc_22172_new_n9005_), .Y(core__0v1_reg_63_0__57_));
AND2X2 AND2X2_4964 ( .A(core__abc_22172_new_n9010_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9011_));
AND2X2 AND2X2_4965 ( .A(core__abc_22172_new_n9011_), .B(core__abc_22172_new_n9008_), .Y(core__abc_22172_new_n9012_));
AND2X2 AND2X2_4966 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_58_), .Y(core__abc_22172_new_n9013_));
AND2X2 AND2X2_4967 ( .A(core__abc_22172_new_n9017_), .B(reset_n), .Y(core__abc_22172_new_n9018_));
AND2X2 AND2X2_4968 ( .A(core__abc_22172_new_n9016_), .B(core__abc_22172_new_n9018_), .Y(core__0v1_reg_63_0__58_));
AND2X2 AND2X2_4969 ( .A(core__abc_22172_new_n9022_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9023_));
AND2X2 AND2X2_497 ( .A(_abc_19873_new_n1607_), .B(word3_reg_31_), .Y(_abc_19873_new_n1732_));
AND2X2 AND2X2_4970 ( .A(core__abc_22172_new_n9023_), .B(core__abc_22172_new_n9021_), .Y(core__abc_22172_new_n9024_));
AND2X2 AND2X2_4971 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_59_), .Y(core__abc_22172_new_n9025_));
AND2X2 AND2X2_4972 ( .A(core__abc_22172_new_n9029_), .B(reset_n), .Y(core__abc_22172_new_n9030_));
AND2X2 AND2X2_4973 ( .A(core__abc_22172_new_n9028_), .B(core__abc_22172_new_n9030_), .Y(core__0v1_reg_63_0__59_));
AND2X2 AND2X2_4974 ( .A(core__abc_22172_new_n9034_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9035_));
AND2X2 AND2X2_4975 ( .A(core__abc_22172_new_n9035_), .B(core__abc_22172_new_n9032_), .Y(core__abc_22172_new_n9036_));
AND2X2 AND2X2_4976 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_60_), .Y(core__abc_22172_new_n9037_));
AND2X2 AND2X2_4977 ( .A(core__abc_22172_new_n2623_), .B(core_key_124_), .Y(core__abc_22172_new_n9038_));
AND2X2 AND2X2_4978 ( .A(core__abc_22172_new_n9042_), .B(reset_n), .Y(core__abc_22172_new_n9043_));
AND2X2 AND2X2_4979 ( .A(core__abc_22172_new_n9041_), .B(core__abc_22172_new_n9043_), .Y(core__0v1_reg_63_0__60_));
AND2X2 AND2X2_498 ( .A(_abc_19873_new_n1733_), .B(reset_n), .Y(_0word3_reg_31_0__31_));
AND2X2 AND2X2_4980 ( .A(core__abc_22172_new_n9046_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9047_));
AND2X2 AND2X2_4981 ( .A(core__abc_22172_new_n9047_), .B(core__abc_22172_new_n9045_), .Y(core__abc_22172_new_n9048_));
AND2X2 AND2X2_4982 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_61_), .Y(core__abc_22172_new_n9049_));
AND2X2 AND2X2_4983 ( .A(core__abc_22172_new_n9053_), .B(reset_n), .Y(core__abc_22172_new_n9054_));
AND2X2 AND2X2_4984 ( .A(core__abc_22172_new_n9052_), .B(core__abc_22172_new_n9054_), .Y(core__0v1_reg_63_0__61_));
AND2X2 AND2X2_4985 ( .A(core__abc_22172_new_n9057_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9058_));
AND2X2 AND2X2_4986 ( .A(core__abc_22172_new_n9058_), .B(core__abc_22172_new_n9056_), .Y(core__abc_22172_new_n9059_));
AND2X2 AND2X2_4987 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_62_), .Y(core__abc_22172_new_n9060_));
AND2X2 AND2X2_4988 ( .A(core__abc_22172_new_n9064_), .B(reset_n), .Y(core__abc_22172_new_n9065_));
AND2X2 AND2X2_4989 ( .A(core__abc_22172_new_n9063_), .B(core__abc_22172_new_n9065_), .Y(core__0v1_reg_63_0__62_));
AND2X2 AND2X2_499 ( .A(core_siphash_valid_reg), .B(core_siphash_word_64_), .Y(_abc_19873_new_n1735_));
AND2X2 AND2X2_4990 ( .A(core__abc_22172_new_n9069_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9070_));
AND2X2 AND2X2_4991 ( .A(core__abc_22172_new_n9070_), .B(core__abc_22172_new_n9068_), .Y(core__abc_22172_new_n9071_));
AND2X2 AND2X2_4992 ( .A(core__abc_22172_new_n8289_), .B(core_v1_reg_63_), .Y(core__abc_22172_new_n9072_));
AND2X2 AND2X2_4993 ( .A(core__abc_22172_new_n9076_), .B(reset_n), .Y(core__abc_22172_new_n9077_));
AND2X2 AND2X2_4994 ( .A(core__abc_22172_new_n9075_), .B(core__abc_22172_new_n9077_), .Y(core__0v1_reg_63_0__63_));
AND2X2 AND2X2_4995 ( .A(core__abc_22172_new_n2630_), .B(core__abc_22172_new_n2623_), .Y(core__abc_22172_new_n9079_));
AND2X2 AND2X2_4996 ( .A(core__abc_22172_new_n3199_), .B(core__abc_22172_new_n9079_), .Y(core__abc_22172_new_n9080_));
AND2X2 AND2X2_4997 ( .A(core__abc_22172_new_n6878_), .B(core__abc_22172_new_n9081_), .Y(core__abc_22172_new_n9082_));
AND2X2 AND2X2_4998 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_0_), .Y(core__abc_22172_new_n9084_));
AND2X2 AND2X2_4999 ( .A(core__abc_22172_new_n3044_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9085_));
AND2X2 AND2X2_5 ( .A(_abc_19873_new_n877_), .B(_abc_19873_new_n878_), .Y(_abc_19873_new_n879_));
AND2X2 AND2X2_50 ( .A(_abc_19873_new_n888_), .B(core_mi_1_), .Y(_abc_19873_new_n940_));
AND2X2 AND2X2_500 ( .A(_abc_19873_new_n1607_), .B(word2_reg_0_), .Y(_abc_19873_new_n1736_));
AND2X2 AND2X2_5000 ( .A(core_v0_reg_0_), .B(core_mi_reg_0_), .Y(core__abc_22172_new_n9087_));
AND2X2 AND2X2_5001 ( .A(core__abc_22172_new_n9088_), .B(core__abc_22172_new_n9086_), .Y(core__abc_22172_new_n9089_));
AND2X2 AND2X2_5002 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9089_), .Y(core__abc_22172_new_n9090_));
AND2X2 AND2X2_5003 ( .A(core__abc_22172_new_n9092_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9093_));
AND2X2 AND2X2_5004 ( .A(core__abc_22172_new_n9094_), .B(reset_n), .Y(core__0v0_reg_63_0__0_));
AND2X2 AND2X2_5005 ( .A(core__abc_22172_new_n3255_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9096_));
AND2X2 AND2X2_5006 ( .A(core_v0_reg_1_), .B(core_mi_reg_1_), .Y(core__abc_22172_new_n9098_));
AND2X2 AND2X2_5007 ( .A(core__abc_22172_new_n9099_), .B(core__abc_22172_new_n9097_), .Y(core__abc_22172_new_n9100_));
AND2X2 AND2X2_5008 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9100_), .Y(core__abc_22172_new_n9101_));
AND2X2 AND2X2_5009 ( .A(core__abc_22172_new_n9103_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9104_));
AND2X2 AND2X2_501 ( .A(_abc_19873_new_n1737_), .B(reset_n), .Y(_0word2_reg_31_0__0_));
AND2X2 AND2X2_5010 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_1_), .Y(core__abc_22172_new_n9105_));
AND2X2 AND2X2_5011 ( .A(core__abc_22172_new_n9106_), .B(reset_n), .Y(core__0v0_reg_63_0__1_));
AND2X2 AND2X2_5012 ( .A(core__abc_22172_new_n3320_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9108_));
AND2X2 AND2X2_5013 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n9109_), .Y(core__abc_22172_new_n9110_));
AND2X2 AND2X2_5014 ( .A(core_v0_reg_2_), .B(core_mi_reg_2_), .Y(core__abc_22172_new_n9112_));
AND2X2 AND2X2_5015 ( .A(core__abc_22172_new_n9113_), .B(core__abc_22172_new_n9111_), .Y(core__abc_22172_new_n9114_));
AND2X2 AND2X2_5016 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9114_), .Y(core__abc_22172_new_n9115_));
AND2X2 AND2X2_5017 ( .A(core__abc_22172_new_n9117_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9118_));
AND2X2 AND2X2_5018 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_2_), .Y(core__abc_22172_new_n9119_));
AND2X2 AND2X2_5019 ( .A(core__abc_22172_new_n9120_), .B(reset_n), .Y(core__0v0_reg_63_0__2_));
AND2X2 AND2X2_502 ( .A(core_siphash_valid_reg), .B(core_siphash_word_65_), .Y(_abc_19873_new_n1739_));
AND2X2 AND2X2_5020 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_3_), .Y(core__abc_22172_new_n9122_));
AND2X2 AND2X2_5021 ( .A(core__abc_22172_new_n3393_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9123_));
AND2X2 AND2X2_5022 ( .A(core_v0_reg_3_), .B(core_mi_reg_3_), .Y(core__abc_22172_new_n9125_));
AND2X2 AND2X2_5023 ( .A(core__abc_22172_new_n9126_), .B(core__abc_22172_new_n9124_), .Y(core__abc_22172_new_n9127_));
AND2X2 AND2X2_5024 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9127_), .Y(core__abc_22172_new_n9128_));
AND2X2 AND2X2_5025 ( .A(core__abc_22172_new_n9130_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9131_));
AND2X2 AND2X2_5026 ( .A(core__abc_22172_new_n9132_), .B(reset_n), .Y(core__0v0_reg_63_0__3_));
AND2X2 AND2X2_5027 ( .A(core__abc_22172_new_n3442_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9134_));
AND2X2 AND2X2_5028 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n9135_), .Y(core__abc_22172_new_n9136_));
AND2X2 AND2X2_5029 ( .A(core_v0_reg_4_), .B(core_mi_reg_4_), .Y(core__abc_22172_new_n9138_));
AND2X2 AND2X2_503 ( .A(_abc_19873_new_n1607_), .B(word2_reg_1_), .Y(_abc_19873_new_n1740_));
AND2X2 AND2X2_5030 ( .A(core__abc_22172_new_n9139_), .B(core__abc_22172_new_n9137_), .Y(core__abc_22172_new_n9140_));
AND2X2 AND2X2_5031 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9140_), .Y(core__abc_22172_new_n9141_));
AND2X2 AND2X2_5032 ( .A(core__abc_22172_new_n9143_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9144_));
AND2X2 AND2X2_5033 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_4_), .Y(core__abc_22172_new_n9145_));
AND2X2 AND2X2_5034 ( .A(core__abc_22172_new_n9146_), .B(reset_n), .Y(core__0v0_reg_63_0__4_));
AND2X2 AND2X2_5035 ( .A(core__abc_22172_new_n3500_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9148_));
AND2X2 AND2X2_5036 ( .A(core_v0_reg_5_), .B(core_mi_reg_5_), .Y(core__abc_22172_new_n9150_));
AND2X2 AND2X2_5037 ( .A(core__abc_22172_new_n9151_), .B(core__abc_22172_new_n9149_), .Y(core__abc_22172_new_n9152_));
AND2X2 AND2X2_5038 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9152_), .Y(core__abc_22172_new_n9153_));
AND2X2 AND2X2_5039 ( .A(core__abc_22172_new_n9155_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9156_));
AND2X2 AND2X2_504 ( .A(_abc_19873_new_n1741_), .B(reset_n), .Y(_0word2_reg_31_0__1_));
AND2X2 AND2X2_5040 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_5_), .Y(core__abc_22172_new_n9157_));
AND2X2 AND2X2_5041 ( .A(core__abc_22172_new_n9158_), .B(reset_n), .Y(core__0v0_reg_63_0__5_));
AND2X2 AND2X2_5042 ( .A(core__abc_22172_new_n3573_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9160_));
AND2X2 AND2X2_5043 ( .A(core_v0_reg_6_), .B(core_mi_reg_6_), .Y(core__abc_22172_new_n9162_));
AND2X2 AND2X2_5044 ( .A(core__abc_22172_new_n9163_), .B(core__abc_22172_new_n9161_), .Y(core__abc_22172_new_n9164_));
AND2X2 AND2X2_5045 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9164_), .Y(core__abc_22172_new_n9165_));
AND2X2 AND2X2_5046 ( .A(core__abc_22172_new_n9167_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9168_));
AND2X2 AND2X2_5047 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_6_), .Y(core__abc_22172_new_n9169_));
AND2X2 AND2X2_5048 ( .A(core__abc_22172_new_n9170_), .B(reset_n), .Y(core__0v0_reg_63_0__6_));
AND2X2 AND2X2_5049 ( .A(core__abc_22172_new_n3631_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9172_));
AND2X2 AND2X2_505 ( .A(core_siphash_valid_reg), .B(core_siphash_word_66_), .Y(_abc_19873_new_n1743_));
AND2X2 AND2X2_5050 ( .A(core_v0_reg_7_), .B(core_mi_reg_7_), .Y(core__abc_22172_new_n9174_));
AND2X2 AND2X2_5051 ( .A(core__abc_22172_new_n9175_), .B(core__abc_22172_new_n9173_), .Y(core__abc_22172_new_n9176_));
AND2X2 AND2X2_5052 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9176_), .Y(core__abc_22172_new_n9177_));
AND2X2 AND2X2_5053 ( .A(core__abc_22172_new_n9179_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9180_));
AND2X2 AND2X2_5054 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_7_), .Y(core__abc_22172_new_n9181_));
AND2X2 AND2X2_5055 ( .A(core__abc_22172_new_n9182_), .B(reset_n), .Y(core__0v0_reg_63_0__7_));
AND2X2 AND2X2_5056 ( .A(core__abc_22172_new_n3706_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9184_));
AND2X2 AND2X2_5057 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n9185_), .Y(core__abc_22172_new_n9186_));
AND2X2 AND2X2_5058 ( .A(core_v0_reg_8_), .B(core_mi_reg_8_), .Y(core__abc_22172_new_n9188_));
AND2X2 AND2X2_5059 ( .A(core__abc_22172_new_n9189_), .B(core__abc_22172_new_n9187_), .Y(core__abc_22172_new_n9190_));
AND2X2 AND2X2_506 ( .A(_abc_19873_new_n1607_), .B(word2_reg_2_), .Y(_abc_19873_new_n1744_));
AND2X2 AND2X2_5060 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9190_), .Y(core__abc_22172_new_n9191_));
AND2X2 AND2X2_5061 ( .A(core__abc_22172_new_n9193_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9194_));
AND2X2 AND2X2_5062 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_8_), .Y(core__abc_22172_new_n9195_));
AND2X2 AND2X2_5063 ( .A(core__abc_22172_new_n9196_), .B(reset_n), .Y(core__0v0_reg_63_0__8_));
AND2X2 AND2X2_5064 ( .A(core__abc_22172_new_n3768_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9198_));
AND2X2 AND2X2_5065 ( .A(core__abc_22172_new_n3214_), .B(core_key_9_), .Y(core__abc_22172_new_n9199_));
AND2X2 AND2X2_5066 ( .A(core_v0_reg_9_), .B(core_mi_reg_9_), .Y(core__abc_22172_new_n9201_));
AND2X2 AND2X2_5067 ( .A(core__abc_22172_new_n9202_), .B(core__abc_22172_new_n9200_), .Y(core__abc_22172_new_n9203_));
AND2X2 AND2X2_5068 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9203_), .Y(core__abc_22172_new_n9204_));
AND2X2 AND2X2_5069 ( .A(core__abc_22172_new_n9206_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9207_));
AND2X2 AND2X2_507 ( .A(_abc_19873_new_n1745_), .B(reset_n), .Y(_0word2_reg_31_0__2_));
AND2X2 AND2X2_5070 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_9_), .Y(core__abc_22172_new_n9208_));
AND2X2 AND2X2_5071 ( .A(core__abc_22172_new_n9209_), .B(reset_n), .Y(core__0v0_reg_63_0__9_));
AND2X2 AND2X2_5072 ( .A(core__abc_22172_new_n3840_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9211_));
AND2X2 AND2X2_5073 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n9212_), .Y(core__abc_22172_new_n9213_));
AND2X2 AND2X2_5074 ( .A(core_v0_reg_10_), .B(core_mi_reg_10_), .Y(core__abc_22172_new_n9215_));
AND2X2 AND2X2_5075 ( .A(core__abc_22172_new_n9216_), .B(core__abc_22172_new_n9214_), .Y(core__abc_22172_new_n9217_));
AND2X2 AND2X2_5076 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9217_), .Y(core__abc_22172_new_n9218_));
AND2X2 AND2X2_5077 ( .A(core__abc_22172_new_n9220_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9221_));
AND2X2 AND2X2_5078 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_10_), .Y(core__abc_22172_new_n9222_));
AND2X2 AND2X2_5079 ( .A(core__abc_22172_new_n9223_), .B(reset_n), .Y(core__0v0_reg_63_0__10_));
AND2X2 AND2X2_508 ( .A(core_siphash_valid_reg), .B(core_siphash_word_67_), .Y(_abc_19873_new_n1747_));
AND2X2 AND2X2_5080 ( .A(core__abc_22172_new_n3894_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9225_));
AND2X2 AND2X2_5081 ( .A(core_v0_reg_11_), .B(core_mi_reg_11_), .Y(core__abc_22172_new_n9227_));
AND2X2 AND2X2_5082 ( .A(core__abc_22172_new_n9228_), .B(core__abc_22172_new_n9226_), .Y(core__abc_22172_new_n9229_));
AND2X2 AND2X2_5083 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9229_), .Y(core__abc_22172_new_n9230_));
AND2X2 AND2X2_5084 ( .A(core__abc_22172_new_n9232_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9233_));
AND2X2 AND2X2_5085 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_11_), .Y(core__abc_22172_new_n9234_));
AND2X2 AND2X2_5086 ( .A(core__abc_22172_new_n9235_), .B(reset_n), .Y(core__0v0_reg_63_0__11_));
AND2X2 AND2X2_5087 ( .A(core__abc_22172_new_n3967_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9237_));
AND2X2 AND2X2_5088 ( .A(core__abc_22172_new_n3214_), .B(core_key_12_), .Y(core__abc_22172_new_n9238_));
AND2X2 AND2X2_5089 ( .A(core_v0_reg_12_), .B(core_mi_reg_12_), .Y(core__abc_22172_new_n9240_));
AND2X2 AND2X2_509 ( .A(_abc_19873_new_n1607_), .B(word2_reg_3_), .Y(_abc_19873_new_n1748_));
AND2X2 AND2X2_5090 ( .A(core__abc_22172_new_n9241_), .B(core__abc_22172_new_n9239_), .Y(core__abc_22172_new_n9242_));
AND2X2 AND2X2_5091 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9242_), .Y(core__abc_22172_new_n9243_));
AND2X2 AND2X2_5092 ( .A(core__abc_22172_new_n9245_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9246_));
AND2X2 AND2X2_5093 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_12_), .Y(core__abc_22172_new_n9247_));
AND2X2 AND2X2_5094 ( .A(core__abc_22172_new_n9248_), .B(reset_n), .Y(core__0v0_reg_63_0__12_));
AND2X2 AND2X2_5095 ( .A(core__abc_22172_new_n4027_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9250_));
AND2X2 AND2X2_5096 ( .A(core_v0_reg_13_), .B(core_mi_reg_13_), .Y(core__abc_22172_new_n9252_));
AND2X2 AND2X2_5097 ( .A(core__abc_22172_new_n9253_), .B(core__abc_22172_new_n9251_), .Y(core__abc_22172_new_n9254_));
AND2X2 AND2X2_5098 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9254_), .Y(core__abc_22172_new_n9255_));
AND2X2 AND2X2_5099 ( .A(core__abc_22172_new_n9257_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9258_));
AND2X2 AND2X2_51 ( .A(_abc_19873_new_n894_), .B(core_compress), .Y(_abc_19873_new_n942_));
AND2X2 AND2X2_510 ( .A(_abc_19873_new_n1749_), .B(reset_n), .Y(_0word2_reg_31_0__3_));
AND2X2 AND2X2_5100 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_13_), .Y(core__abc_22172_new_n9259_));
AND2X2 AND2X2_5101 ( .A(core__abc_22172_new_n9260_), .B(reset_n), .Y(core__0v0_reg_63_0__13_));
AND2X2 AND2X2_5102 ( .A(core__abc_22172_new_n4098_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9262_));
AND2X2 AND2X2_5103 ( .A(core_v0_reg_14_), .B(core_mi_reg_14_), .Y(core__abc_22172_new_n9264_));
AND2X2 AND2X2_5104 ( .A(core__abc_22172_new_n9265_), .B(core__abc_22172_new_n9263_), .Y(core__abc_22172_new_n9266_));
AND2X2 AND2X2_5105 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9266_), .Y(core__abc_22172_new_n9267_));
AND2X2 AND2X2_5106 ( .A(core__abc_22172_new_n9269_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9270_));
AND2X2 AND2X2_5107 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_14_), .Y(core__abc_22172_new_n9271_));
AND2X2 AND2X2_5108 ( .A(core__abc_22172_new_n9272_), .B(reset_n), .Y(core__0v0_reg_63_0__14_));
AND2X2 AND2X2_5109 ( .A(core__abc_22172_new_n4154_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9274_));
AND2X2 AND2X2_511 ( .A(core_siphash_valid_reg), .B(core_siphash_word_68_), .Y(_abc_19873_new_n1751_));
AND2X2 AND2X2_5110 ( .A(core_v0_reg_15_), .B(core_mi_reg_15_), .Y(core__abc_22172_new_n9276_));
AND2X2 AND2X2_5111 ( .A(core__abc_22172_new_n9277_), .B(core__abc_22172_new_n9275_), .Y(core__abc_22172_new_n9278_));
AND2X2 AND2X2_5112 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9278_), .Y(core__abc_22172_new_n9279_));
AND2X2 AND2X2_5113 ( .A(core__abc_22172_new_n9281_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9282_));
AND2X2 AND2X2_5114 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_15_), .Y(core__abc_22172_new_n9283_));
AND2X2 AND2X2_5115 ( .A(core__abc_22172_new_n9284_), .B(reset_n), .Y(core__0v0_reg_63_0__15_));
AND2X2 AND2X2_5116 ( .A(core__abc_22172_new_n4239_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9286_));
AND2X2 AND2X2_5117 ( .A(core_v0_reg_16_), .B(core_mi_reg_16_), .Y(core__abc_22172_new_n9288_));
AND2X2 AND2X2_5118 ( .A(core__abc_22172_new_n9289_), .B(core__abc_22172_new_n9287_), .Y(core__abc_22172_new_n9290_));
AND2X2 AND2X2_5119 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9290_), .Y(core__abc_22172_new_n9291_));
AND2X2 AND2X2_512 ( .A(_abc_19873_new_n1607_), .B(word2_reg_4_), .Y(_abc_19873_new_n1752_));
AND2X2 AND2X2_5120 ( .A(core__abc_22172_new_n9293_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9294_));
AND2X2 AND2X2_5121 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_16_), .Y(core__abc_22172_new_n9295_));
AND2X2 AND2X2_5122 ( .A(core__abc_22172_new_n9296_), .B(reset_n), .Y(core__0v0_reg_63_0__16_));
AND2X2 AND2X2_5123 ( .A(core__abc_22172_new_n4306_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9298_));
AND2X2 AND2X2_5124 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n9299_), .Y(core__abc_22172_new_n9300_));
AND2X2 AND2X2_5125 ( .A(core_v0_reg_17_), .B(core_mi_reg_17_), .Y(core__abc_22172_new_n9302_));
AND2X2 AND2X2_5126 ( .A(core__abc_22172_new_n9303_), .B(core__abc_22172_new_n9301_), .Y(core__abc_22172_new_n9304_));
AND2X2 AND2X2_5127 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9304_), .Y(core__abc_22172_new_n9305_));
AND2X2 AND2X2_5128 ( .A(core__abc_22172_new_n9307_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9308_));
AND2X2 AND2X2_5129 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_17_), .Y(core__abc_22172_new_n9309_));
AND2X2 AND2X2_513 ( .A(_abc_19873_new_n1753_), .B(reset_n), .Y(_0word2_reg_31_0__4_));
AND2X2 AND2X2_5130 ( .A(core__abc_22172_new_n9310_), .B(reset_n), .Y(core__0v0_reg_63_0__17_));
AND2X2 AND2X2_5131 ( .A(core__abc_22172_new_n4378_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9312_));
AND2X2 AND2X2_5132 ( .A(core__abc_22172_new_n3214_), .B(core_key_18_), .Y(core__abc_22172_new_n9313_));
AND2X2 AND2X2_5133 ( .A(core_v0_reg_18_), .B(core_mi_reg_18_), .Y(core__abc_22172_new_n9315_));
AND2X2 AND2X2_5134 ( .A(core__abc_22172_new_n9316_), .B(core__abc_22172_new_n9314_), .Y(core__abc_22172_new_n9317_));
AND2X2 AND2X2_5135 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9317_), .Y(core__abc_22172_new_n9318_));
AND2X2 AND2X2_5136 ( .A(core__abc_22172_new_n9320_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9321_));
AND2X2 AND2X2_5137 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_18_), .Y(core__abc_22172_new_n9322_));
AND2X2 AND2X2_5138 ( .A(core__abc_22172_new_n9323_), .B(reset_n), .Y(core__0v0_reg_63_0__18_));
AND2X2 AND2X2_5139 ( .A(core__abc_22172_new_n4420_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9325_));
AND2X2 AND2X2_514 ( .A(core_siphash_valid_reg), .B(core_siphash_word_69_), .Y(_abc_19873_new_n1755_));
AND2X2 AND2X2_5140 ( .A(core_v0_reg_19_), .B(core_mi_reg_19_), .Y(core__abc_22172_new_n9327_));
AND2X2 AND2X2_5141 ( .A(core__abc_22172_new_n9328_), .B(core__abc_22172_new_n9326_), .Y(core__abc_22172_new_n9329_));
AND2X2 AND2X2_5142 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9329_), .Y(core__abc_22172_new_n9330_));
AND2X2 AND2X2_5143 ( .A(core__abc_22172_new_n9332_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9333_));
AND2X2 AND2X2_5144 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_19_), .Y(core__abc_22172_new_n9334_));
AND2X2 AND2X2_5145 ( .A(core__abc_22172_new_n9335_), .B(reset_n), .Y(core__0v0_reg_63_0__19_));
AND2X2 AND2X2_5146 ( .A(core__abc_22172_new_n4492_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9337_));
AND2X2 AND2X2_5147 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n9338_), .Y(core__abc_22172_new_n9339_));
AND2X2 AND2X2_5148 ( .A(core_v0_reg_20_), .B(core_mi_reg_20_), .Y(core__abc_22172_new_n9341_));
AND2X2 AND2X2_5149 ( .A(core__abc_22172_new_n9342_), .B(core__abc_22172_new_n9340_), .Y(core__abc_22172_new_n9343_));
AND2X2 AND2X2_515 ( .A(_abc_19873_new_n1607_), .B(word2_reg_5_), .Y(_abc_19873_new_n1756_));
AND2X2 AND2X2_5150 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9343_), .Y(core__abc_22172_new_n9344_));
AND2X2 AND2X2_5151 ( .A(core__abc_22172_new_n9346_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9347_));
AND2X2 AND2X2_5152 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_20_), .Y(core__abc_22172_new_n9348_));
AND2X2 AND2X2_5153 ( .A(core__abc_22172_new_n9349_), .B(reset_n), .Y(core__0v0_reg_63_0__20_));
AND2X2 AND2X2_5154 ( .A(core__abc_22172_new_n4548_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9351_));
AND2X2 AND2X2_5155 ( .A(core_v0_reg_21_), .B(core_mi_reg_21_), .Y(core__abc_22172_new_n9353_));
AND2X2 AND2X2_5156 ( .A(core__abc_22172_new_n9354_), .B(core__abc_22172_new_n9352_), .Y(core__abc_22172_new_n9355_));
AND2X2 AND2X2_5157 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9355_), .Y(core__abc_22172_new_n9356_));
AND2X2 AND2X2_5158 ( .A(core__abc_22172_new_n9358_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9359_));
AND2X2 AND2X2_5159 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_21_), .Y(core__abc_22172_new_n9360_));
AND2X2 AND2X2_516 ( .A(_abc_19873_new_n1757_), .B(reset_n), .Y(_0word2_reg_31_0__5_));
AND2X2 AND2X2_5160 ( .A(core__abc_22172_new_n9361_), .B(reset_n), .Y(core__0v0_reg_63_0__21_));
AND2X2 AND2X2_5161 ( .A(core__abc_22172_new_n4602_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9363_));
AND2X2 AND2X2_5162 ( .A(core_v0_reg_22_), .B(core_mi_reg_22_), .Y(core__abc_22172_new_n9365_));
AND2X2 AND2X2_5163 ( .A(core__abc_22172_new_n9366_), .B(core__abc_22172_new_n9364_), .Y(core__abc_22172_new_n9367_));
AND2X2 AND2X2_5164 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9367_), .Y(core__abc_22172_new_n9368_));
AND2X2 AND2X2_5165 ( .A(core__abc_22172_new_n9370_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9371_));
AND2X2 AND2X2_5166 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_22_), .Y(core__abc_22172_new_n9372_));
AND2X2 AND2X2_5167 ( .A(core__abc_22172_new_n9373_), .B(reset_n), .Y(core__0v0_reg_63_0__22_));
AND2X2 AND2X2_5168 ( .A(core__abc_22172_new_n4646_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9375_));
AND2X2 AND2X2_5169 ( .A(core_v0_reg_23_), .B(core_mi_reg_23_), .Y(core__abc_22172_new_n9377_));
AND2X2 AND2X2_517 ( .A(core_siphash_valid_reg), .B(core_siphash_word_70_), .Y(_abc_19873_new_n1759_));
AND2X2 AND2X2_5170 ( .A(core__abc_22172_new_n9378_), .B(core__abc_22172_new_n9376_), .Y(core__abc_22172_new_n9379_));
AND2X2 AND2X2_5171 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9379_), .Y(core__abc_22172_new_n9380_));
AND2X2 AND2X2_5172 ( .A(core__abc_22172_new_n9382_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9383_));
AND2X2 AND2X2_5173 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_23_), .Y(core__abc_22172_new_n9384_));
AND2X2 AND2X2_5174 ( .A(core__abc_22172_new_n9385_), .B(reset_n), .Y(core__0v0_reg_63_0__23_));
AND2X2 AND2X2_5175 ( .A(core__abc_22172_new_n4717_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9387_));
AND2X2 AND2X2_5176 ( .A(core_v0_reg_24_), .B(core_mi_reg_24_), .Y(core__abc_22172_new_n9389_));
AND2X2 AND2X2_5177 ( .A(core__abc_22172_new_n9390_), .B(core__abc_22172_new_n9388_), .Y(core__abc_22172_new_n9391_));
AND2X2 AND2X2_5178 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9391_), .Y(core__abc_22172_new_n9392_));
AND2X2 AND2X2_5179 ( .A(core__abc_22172_new_n9394_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9395_));
AND2X2 AND2X2_518 ( .A(_abc_19873_new_n1607_), .B(word2_reg_6_), .Y(_abc_19873_new_n1760_));
AND2X2 AND2X2_5180 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_24_), .Y(core__abc_22172_new_n9396_));
AND2X2 AND2X2_5181 ( .A(core__abc_22172_new_n9397_), .B(reset_n), .Y(core__0v0_reg_63_0__24_));
AND2X2 AND2X2_5182 ( .A(core__abc_22172_new_n4760_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9399_));
AND2X2 AND2X2_5183 ( .A(core__abc_22172_new_n3214_), .B(core_key_25_), .Y(core__abc_22172_new_n9400_));
AND2X2 AND2X2_5184 ( .A(core_v0_reg_25_), .B(core_mi_reg_25_), .Y(core__abc_22172_new_n9402_));
AND2X2 AND2X2_5185 ( .A(core__abc_22172_new_n9403_), .B(core__abc_22172_new_n9401_), .Y(core__abc_22172_new_n9404_));
AND2X2 AND2X2_5186 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9404_), .Y(core__abc_22172_new_n9405_));
AND2X2 AND2X2_5187 ( .A(core__abc_22172_new_n9407_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9408_));
AND2X2 AND2X2_5188 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_25_), .Y(core__abc_22172_new_n9409_));
AND2X2 AND2X2_5189 ( .A(core__abc_22172_new_n9410_), .B(reset_n), .Y(core__0v0_reg_63_0__25_));
AND2X2 AND2X2_519 ( .A(_abc_19873_new_n1761_), .B(reset_n), .Y(_0word2_reg_31_0__6_));
AND2X2 AND2X2_5190 ( .A(core__abc_22172_new_n4813_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9412_));
AND2X2 AND2X2_5191 ( .A(core__abc_22172_new_n3214_), .B(core_key_26_), .Y(core__abc_22172_new_n9413_));
AND2X2 AND2X2_5192 ( .A(core_v0_reg_26_), .B(core_mi_reg_26_), .Y(core__abc_22172_new_n9415_));
AND2X2 AND2X2_5193 ( .A(core__abc_22172_new_n9416_), .B(core__abc_22172_new_n9414_), .Y(core__abc_22172_new_n9417_));
AND2X2 AND2X2_5194 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9417_), .Y(core__abc_22172_new_n9418_));
AND2X2 AND2X2_5195 ( .A(core__abc_22172_new_n9420_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9421_));
AND2X2 AND2X2_5196 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_26_), .Y(core__abc_22172_new_n9422_));
AND2X2 AND2X2_5197 ( .A(core__abc_22172_new_n9423_), .B(reset_n), .Y(core__0v0_reg_63_0__26_));
AND2X2 AND2X2_5198 ( .A(core__abc_22172_new_n4855_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9425_));
AND2X2 AND2X2_5199 ( .A(core__abc_22172_new_n3214_), .B(core_key_27_), .Y(core__abc_22172_new_n9426_));
AND2X2 AND2X2_52 ( .A(_abc_19873_new_n897_), .B(core_compression_rounds_1_), .Y(_abc_19873_new_n943_));
AND2X2 AND2X2_520 ( .A(core_siphash_valid_reg), .B(core_siphash_word_71_), .Y(_abc_19873_new_n1763_));
AND2X2 AND2X2_5200 ( .A(core_v0_reg_27_), .B(core_mi_reg_27_), .Y(core__abc_22172_new_n9428_));
AND2X2 AND2X2_5201 ( .A(core__abc_22172_new_n9429_), .B(core__abc_22172_new_n9427_), .Y(core__abc_22172_new_n9430_));
AND2X2 AND2X2_5202 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9430_), .Y(core__abc_22172_new_n9431_));
AND2X2 AND2X2_5203 ( .A(core__abc_22172_new_n9433_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9434_));
AND2X2 AND2X2_5204 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_27_), .Y(core__abc_22172_new_n9435_));
AND2X2 AND2X2_5205 ( .A(core__abc_22172_new_n9436_), .B(reset_n), .Y(core__0v0_reg_63_0__27_));
AND2X2 AND2X2_5206 ( .A(core__abc_22172_new_n4921_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9438_));
AND2X2 AND2X2_5207 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n9439_), .Y(core__abc_22172_new_n9440_));
AND2X2 AND2X2_5208 ( .A(core_v0_reg_28_), .B(core_mi_reg_28_), .Y(core__abc_22172_new_n9442_));
AND2X2 AND2X2_5209 ( .A(core__abc_22172_new_n9443_), .B(core__abc_22172_new_n9441_), .Y(core__abc_22172_new_n9444_));
AND2X2 AND2X2_521 ( .A(_abc_19873_new_n1607_), .B(word2_reg_7_), .Y(_abc_19873_new_n1764_));
AND2X2 AND2X2_5210 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9444_), .Y(core__abc_22172_new_n9445_));
AND2X2 AND2X2_5211 ( .A(core__abc_22172_new_n9447_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9448_));
AND2X2 AND2X2_5212 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_28_), .Y(core__abc_22172_new_n9449_));
AND2X2 AND2X2_5213 ( .A(core__abc_22172_new_n9450_), .B(reset_n), .Y(core__0v0_reg_63_0__28_));
AND2X2 AND2X2_5214 ( .A(core__abc_22172_new_n4966_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9452_));
AND2X2 AND2X2_5215 ( .A(core_v0_reg_29_), .B(core_mi_reg_29_), .Y(core__abc_22172_new_n9454_));
AND2X2 AND2X2_5216 ( .A(core__abc_22172_new_n9455_), .B(core__abc_22172_new_n9453_), .Y(core__abc_22172_new_n9456_));
AND2X2 AND2X2_5217 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9456_), .Y(core__abc_22172_new_n9457_));
AND2X2 AND2X2_5218 ( .A(core__abc_22172_new_n9459_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9460_));
AND2X2 AND2X2_5219 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_29_), .Y(core__abc_22172_new_n9461_));
AND2X2 AND2X2_522 ( .A(_abc_19873_new_n1765_), .B(reset_n), .Y(_0word2_reg_31_0__7_));
AND2X2 AND2X2_5220 ( .A(core__abc_22172_new_n9462_), .B(reset_n), .Y(core__0v0_reg_63_0__29_));
AND2X2 AND2X2_5221 ( .A(core__abc_22172_new_n5022_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9464_));
AND2X2 AND2X2_5222 ( .A(core_v0_reg_30_), .B(core_mi_reg_30_), .Y(core__abc_22172_new_n9466_));
AND2X2 AND2X2_5223 ( .A(core__abc_22172_new_n9467_), .B(core__abc_22172_new_n9465_), .Y(core__abc_22172_new_n9468_));
AND2X2 AND2X2_5224 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9468_), .Y(core__abc_22172_new_n9469_));
AND2X2 AND2X2_5225 ( .A(core__abc_22172_new_n9471_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9472_));
AND2X2 AND2X2_5226 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_30_), .Y(core__abc_22172_new_n9473_));
AND2X2 AND2X2_5227 ( .A(core__abc_22172_new_n9474_), .B(reset_n), .Y(core__0v0_reg_63_0__30_));
AND2X2 AND2X2_5228 ( .A(core__abc_22172_new_n5068_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9476_));
AND2X2 AND2X2_5229 ( .A(core_v0_reg_31_), .B(core_mi_reg_31_), .Y(core__abc_22172_new_n9478_));
AND2X2 AND2X2_523 ( .A(core_siphash_valid_reg), .B(core_siphash_word_72_), .Y(_abc_19873_new_n1767_));
AND2X2 AND2X2_5230 ( .A(core__abc_22172_new_n9479_), .B(core__abc_22172_new_n9477_), .Y(core__abc_22172_new_n9480_));
AND2X2 AND2X2_5231 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9480_), .Y(core__abc_22172_new_n9481_));
AND2X2 AND2X2_5232 ( .A(core__abc_22172_new_n9483_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9484_));
AND2X2 AND2X2_5233 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_31_), .Y(core__abc_22172_new_n9485_));
AND2X2 AND2X2_5234 ( .A(core__abc_22172_new_n9486_), .B(reset_n), .Y(core__0v0_reg_63_0__31_));
AND2X2 AND2X2_5235 ( .A(core__abc_22172_new_n5143_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9488_));
AND2X2 AND2X2_5236 ( .A(core_v0_reg_32_), .B(core_mi_reg_32_), .Y(core__abc_22172_new_n9490_));
AND2X2 AND2X2_5237 ( .A(core__abc_22172_new_n9491_), .B(core__abc_22172_new_n9489_), .Y(core__abc_22172_new_n9492_));
AND2X2 AND2X2_5238 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9492_), .Y(core__abc_22172_new_n9493_));
AND2X2 AND2X2_5239 ( .A(core__abc_22172_new_n9495_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9496_));
AND2X2 AND2X2_524 ( .A(_abc_19873_new_n1607_), .B(word2_reg_8_), .Y(_abc_19873_new_n1768_));
AND2X2 AND2X2_5240 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_32_), .Y(core__abc_22172_new_n9497_));
AND2X2 AND2X2_5241 ( .A(core__abc_22172_new_n9498_), .B(reset_n), .Y(core__0v0_reg_63_0__32_));
AND2X2 AND2X2_5242 ( .A(core__abc_22172_new_n5182_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9500_));
AND2X2 AND2X2_5243 ( .A(core_v0_reg_33_), .B(core_mi_reg_33_), .Y(core__abc_22172_new_n9502_));
AND2X2 AND2X2_5244 ( .A(core__abc_22172_new_n9503_), .B(core__abc_22172_new_n9501_), .Y(core__abc_22172_new_n9504_));
AND2X2 AND2X2_5245 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9504_), .Y(core__abc_22172_new_n9505_));
AND2X2 AND2X2_5246 ( .A(core__abc_22172_new_n9507_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9508_));
AND2X2 AND2X2_5247 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_33_), .Y(core__abc_22172_new_n9509_));
AND2X2 AND2X2_5248 ( .A(core__abc_22172_new_n9510_), .B(reset_n), .Y(core__0v0_reg_63_0__33_));
AND2X2 AND2X2_5249 ( .A(core__abc_22172_new_n5230_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9512_));
AND2X2 AND2X2_525 ( .A(_abc_19873_new_n1769_), .B(reset_n), .Y(_0word2_reg_31_0__8_));
AND2X2 AND2X2_5250 ( .A(core_v0_reg_34_), .B(core_mi_reg_34_), .Y(core__abc_22172_new_n9514_));
AND2X2 AND2X2_5251 ( .A(core__abc_22172_new_n9515_), .B(core__abc_22172_new_n9513_), .Y(core__abc_22172_new_n9516_));
AND2X2 AND2X2_5252 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9516_), .Y(core__abc_22172_new_n9517_));
AND2X2 AND2X2_5253 ( .A(core__abc_22172_new_n9519_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9520_));
AND2X2 AND2X2_5254 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_34_), .Y(core__abc_22172_new_n9521_));
AND2X2 AND2X2_5255 ( .A(core__abc_22172_new_n9522_), .B(reset_n), .Y(core__0v0_reg_63_0__34_));
AND2X2 AND2X2_5256 ( .A(core__abc_22172_new_n5274_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9524_));
AND2X2 AND2X2_5257 ( .A(core_v0_reg_35_), .B(core_mi_reg_35_), .Y(core__abc_22172_new_n9526_));
AND2X2 AND2X2_5258 ( .A(core__abc_22172_new_n9527_), .B(core__abc_22172_new_n9525_), .Y(core__abc_22172_new_n9528_));
AND2X2 AND2X2_5259 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9528_), .Y(core__abc_22172_new_n9529_));
AND2X2 AND2X2_526 ( .A(core_siphash_valid_reg), .B(core_siphash_word_73_), .Y(_abc_19873_new_n1771_));
AND2X2 AND2X2_5260 ( .A(core__abc_22172_new_n9531_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9532_));
AND2X2 AND2X2_5261 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_35_), .Y(core__abc_22172_new_n9533_));
AND2X2 AND2X2_5262 ( .A(core__abc_22172_new_n9534_), .B(reset_n), .Y(core__0v0_reg_63_0__35_));
AND2X2 AND2X2_5263 ( .A(core__abc_22172_new_n5325_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9536_));
AND2X2 AND2X2_5264 ( .A(core_v0_reg_36_), .B(core_mi_reg_36_), .Y(core__abc_22172_new_n9538_));
AND2X2 AND2X2_5265 ( .A(core__abc_22172_new_n9539_), .B(core__abc_22172_new_n9537_), .Y(core__abc_22172_new_n9540_));
AND2X2 AND2X2_5266 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9540_), .Y(core__abc_22172_new_n9541_));
AND2X2 AND2X2_5267 ( .A(core__abc_22172_new_n9543_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9544_));
AND2X2 AND2X2_5268 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_36_), .Y(core__abc_22172_new_n9545_));
AND2X2 AND2X2_5269 ( .A(core__abc_22172_new_n9546_), .B(reset_n), .Y(core__0v0_reg_63_0__36_));
AND2X2 AND2X2_527 ( .A(_abc_19873_new_n1607_), .B(word2_reg_9_), .Y(_abc_19873_new_n1772_));
AND2X2 AND2X2_5270 ( .A(core__abc_22172_new_n5372_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9548_));
AND2X2 AND2X2_5271 ( .A(core_v0_reg_37_), .B(core_mi_reg_37_), .Y(core__abc_22172_new_n9550_));
AND2X2 AND2X2_5272 ( .A(core__abc_22172_new_n9551_), .B(core__abc_22172_new_n9549_), .Y(core__abc_22172_new_n9552_));
AND2X2 AND2X2_5273 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9552_), .Y(core__abc_22172_new_n9553_));
AND2X2 AND2X2_5274 ( .A(core__abc_22172_new_n9555_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9556_));
AND2X2 AND2X2_5275 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_37_), .Y(core__abc_22172_new_n9557_));
AND2X2 AND2X2_5276 ( .A(core__abc_22172_new_n9558_), .B(reset_n), .Y(core__0v0_reg_63_0__37_));
AND2X2 AND2X2_5277 ( .A(core__abc_22172_new_n5423_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9560_));
AND2X2 AND2X2_5278 ( .A(core_v0_reg_38_), .B(core_mi_reg_38_), .Y(core__abc_22172_new_n9562_));
AND2X2 AND2X2_5279 ( .A(core__abc_22172_new_n9563_), .B(core__abc_22172_new_n9561_), .Y(core__abc_22172_new_n9564_));
AND2X2 AND2X2_528 ( .A(_abc_19873_new_n1773_), .B(reset_n), .Y(_0word2_reg_31_0__9_));
AND2X2 AND2X2_5280 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9564_), .Y(core__abc_22172_new_n9565_));
AND2X2 AND2X2_5281 ( .A(core__abc_22172_new_n9567_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9568_));
AND2X2 AND2X2_5282 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_38_), .Y(core__abc_22172_new_n9569_));
AND2X2 AND2X2_5283 ( .A(core__abc_22172_new_n9570_), .B(reset_n), .Y(core__0v0_reg_63_0__38_));
AND2X2 AND2X2_5284 ( .A(core__abc_22172_new_n5464_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9572_));
AND2X2 AND2X2_5285 ( .A(core_v0_reg_39_), .B(core_mi_reg_39_), .Y(core__abc_22172_new_n9574_));
AND2X2 AND2X2_5286 ( .A(core__abc_22172_new_n9575_), .B(core__abc_22172_new_n9573_), .Y(core__abc_22172_new_n9576_));
AND2X2 AND2X2_5287 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9576_), .Y(core__abc_22172_new_n9577_));
AND2X2 AND2X2_5288 ( .A(core__abc_22172_new_n9579_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9580_));
AND2X2 AND2X2_5289 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_39_), .Y(core__abc_22172_new_n9581_));
AND2X2 AND2X2_529 ( .A(core_siphash_valid_reg), .B(core_siphash_word_74_), .Y(_abc_19873_new_n1775_));
AND2X2 AND2X2_5290 ( .A(core__abc_22172_new_n9582_), .B(reset_n), .Y(core__0v0_reg_63_0__39_));
AND2X2 AND2X2_5291 ( .A(core__abc_22172_new_n5521_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9584_));
AND2X2 AND2X2_5292 ( .A(core_v0_reg_40_), .B(core_mi_reg_40_), .Y(core__abc_22172_new_n9586_));
AND2X2 AND2X2_5293 ( .A(core__abc_22172_new_n9587_), .B(core__abc_22172_new_n9585_), .Y(core__abc_22172_new_n9588_));
AND2X2 AND2X2_5294 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9588_), .Y(core__abc_22172_new_n9589_));
AND2X2 AND2X2_5295 ( .A(core__abc_22172_new_n9591_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9592_));
AND2X2 AND2X2_5296 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_40_), .Y(core__abc_22172_new_n9593_));
AND2X2 AND2X2_5297 ( .A(core__abc_22172_new_n9594_), .B(reset_n), .Y(core__0v0_reg_63_0__40_));
AND2X2 AND2X2_5298 ( .A(core__abc_22172_new_n5566_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9596_));
AND2X2 AND2X2_5299 ( .A(core__abc_22172_new_n3214_), .B(core_key_41_), .Y(core__abc_22172_new_n9597_));
AND2X2 AND2X2_53 ( .A(_abc_19873_new_n901_), .B(core_key_1_), .Y(_abc_19873_new_n945_));
AND2X2 AND2X2_530 ( .A(_abc_19873_new_n1607_), .B(word2_reg_10_), .Y(_abc_19873_new_n1776_));
AND2X2 AND2X2_5300 ( .A(core_v0_reg_41_), .B(core_mi_reg_41_), .Y(core__abc_22172_new_n9599_));
AND2X2 AND2X2_5301 ( .A(core__abc_22172_new_n9600_), .B(core__abc_22172_new_n9598_), .Y(core__abc_22172_new_n9601_));
AND2X2 AND2X2_5302 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9601_), .Y(core__abc_22172_new_n9602_));
AND2X2 AND2X2_5303 ( .A(core__abc_22172_new_n9604_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9605_));
AND2X2 AND2X2_5304 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_41_), .Y(core__abc_22172_new_n9606_));
AND2X2 AND2X2_5305 ( .A(core__abc_22172_new_n9607_), .B(reset_n), .Y(core__0v0_reg_63_0__41_));
AND2X2 AND2X2_5306 ( .A(core__abc_22172_new_n5610_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9609_));
AND2X2 AND2X2_5307 ( .A(core_v0_reg_42_), .B(core_mi_reg_42_), .Y(core__abc_22172_new_n9611_));
AND2X2 AND2X2_5308 ( .A(core__abc_22172_new_n9612_), .B(core__abc_22172_new_n9610_), .Y(core__abc_22172_new_n9613_));
AND2X2 AND2X2_5309 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9613_), .Y(core__abc_22172_new_n9614_));
AND2X2 AND2X2_531 ( .A(_abc_19873_new_n1777_), .B(reset_n), .Y(_0word2_reg_31_0__10_));
AND2X2 AND2X2_5310 ( .A(core__abc_22172_new_n9616_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9617_));
AND2X2 AND2X2_5311 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_42_), .Y(core__abc_22172_new_n9618_));
AND2X2 AND2X2_5312 ( .A(core__abc_22172_new_n9619_), .B(reset_n), .Y(core__0v0_reg_63_0__42_));
AND2X2 AND2X2_5313 ( .A(core__abc_22172_new_n5643_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9621_));
AND2X2 AND2X2_5314 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n9622_), .Y(core__abc_22172_new_n9623_));
AND2X2 AND2X2_5315 ( .A(core_v0_reg_43_), .B(core_mi_reg_43_), .Y(core__abc_22172_new_n9625_));
AND2X2 AND2X2_5316 ( .A(core__abc_22172_new_n9626_), .B(core__abc_22172_new_n9624_), .Y(core__abc_22172_new_n9627_));
AND2X2 AND2X2_5317 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9627_), .Y(core__abc_22172_new_n9628_));
AND2X2 AND2X2_5318 ( .A(core__abc_22172_new_n9630_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9631_));
AND2X2 AND2X2_5319 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_43_), .Y(core__abc_22172_new_n9632_));
AND2X2 AND2X2_532 ( .A(core_siphash_valid_reg), .B(core_siphash_word_75_), .Y(_abc_19873_new_n1779_));
AND2X2 AND2X2_5320 ( .A(core__abc_22172_new_n9633_), .B(reset_n), .Y(core__0v0_reg_63_0__43_));
AND2X2 AND2X2_5321 ( .A(core__abc_22172_new_n5695_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9635_));
AND2X2 AND2X2_5322 ( .A(core_v0_reg_44_), .B(core_mi_reg_44_), .Y(core__abc_22172_new_n9637_));
AND2X2 AND2X2_5323 ( .A(core__abc_22172_new_n9638_), .B(core__abc_22172_new_n9636_), .Y(core__abc_22172_new_n9639_));
AND2X2 AND2X2_5324 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9639_), .Y(core__abc_22172_new_n9640_));
AND2X2 AND2X2_5325 ( .A(core__abc_22172_new_n9642_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9643_));
AND2X2 AND2X2_5326 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_44_), .Y(core__abc_22172_new_n9644_));
AND2X2 AND2X2_5327 ( .A(core__abc_22172_new_n9645_), .B(reset_n), .Y(core__0v0_reg_63_0__44_));
AND2X2 AND2X2_5328 ( .A(core__abc_22172_new_n5725_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9647_));
AND2X2 AND2X2_5329 ( .A(core_v0_reg_45_), .B(core_mi_reg_45_), .Y(core__abc_22172_new_n9649_));
AND2X2 AND2X2_533 ( .A(_abc_19873_new_n1607_), .B(word2_reg_11_), .Y(_abc_19873_new_n1780_));
AND2X2 AND2X2_5330 ( .A(core__abc_22172_new_n9650_), .B(core__abc_22172_new_n9648_), .Y(core__abc_22172_new_n9651_));
AND2X2 AND2X2_5331 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9651_), .Y(core__abc_22172_new_n9652_));
AND2X2 AND2X2_5332 ( .A(core__abc_22172_new_n9654_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9655_));
AND2X2 AND2X2_5333 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_45_), .Y(core__abc_22172_new_n9656_));
AND2X2 AND2X2_5334 ( .A(core__abc_22172_new_n9657_), .B(reset_n), .Y(core__0v0_reg_63_0__45_));
AND2X2 AND2X2_5335 ( .A(core__abc_22172_new_n5769_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9659_));
AND2X2 AND2X2_5336 ( .A(core_v0_reg_46_), .B(core_mi_reg_46_), .Y(core__abc_22172_new_n9661_));
AND2X2 AND2X2_5337 ( .A(core__abc_22172_new_n9662_), .B(core__abc_22172_new_n9660_), .Y(core__abc_22172_new_n9663_));
AND2X2 AND2X2_5338 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9663_), .Y(core__abc_22172_new_n9664_));
AND2X2 AND2X2_5339 ( .A(core__abc_22172_new_n9666_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9667_));
AND2X2 AND2X2_534 ( .A(_abc_19873_new_n1781_), .B(reset_n), .Y(_0word2_reg_31_0__11_));
AND2X2 AND2X2_5340 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_46_), .Y(core__abc_22172_new_n9668_));
AND2X2 AND2X2_5341 ( .A(core__abc_22172_new_n9669_), .B(reset_n), .Y(core__0v0_reg_63_0__46_));
AND2X2 AND2X2_5342 ( .A(core__abc_22172_new_n5808_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9671_));
AND2X2 AND2X2_5343 ( .A(core_v0_reg_47_), .B(core_mi_reg_47_), .Y(core__abc_22172_new_n9673_));
AND2X2 AND2X2_5344 ( .A(core__abc_22172_new_n9674_), .B(core__abc_22172_new_n9672_), .Y(core__abc_22172_new_n9675_));
AND2X2 AND2X2_5345 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9675_), .Y(core__abc_22172_new_n9676_));
AND2X2 AND2X2_5346 ( .A(core__abc_22172_new_n9678_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9679_));
AND2X2 AND2X2_5347 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_47_), .Y(core__abc_22172_new_n9680_));
AND2X2 AND2X2_5348 ( .A(core__abc_22172_new_n9681_), .B(reset_n), .Y(core__0v0_reg_63_0__47_));
AND2X2 AND2X2_5349 ( .A(core__abc_22172_new_n5858_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9683_));
AND2X2 AND2X2_535 ( .A(core_siphash_valid_reg), .B(core_siphash_word_76_), .Y(_abc_19873_new_n1783_));
AND2X2 AND2X2_5350 ( .A(core_v0_reg_48_), .B(core_mi_reg_48_), .Y(core__abc_22172_new_n9685_));
AND2X2 AND2X2_5351 ( .A(core__abc_22172_new_n9686_), .B(core__abc_22172_new_n9684_), .Y(core__abc_22172_new_n9687_));
AND2X2 AND2X2_5352 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9687_), .Y(core__abc_22172_new_n9688_));
AND2X2 AND2X2_5353 ( .A(core__abc_22172_new_n9690_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9691_));
AND2X2 AND2X2_5354 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_48_), .Y(core__abc_22172_new_n9692_));
AND2X2 AND2X2_5355 ( .A(core__abc_22172_new_n9693_), .B(reset_n), .Y(core__0v0_reg_63_0__48_));
AND2X2 AND2X2_5356 ( .A(core__abc_22172_new_n5896_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9695_));
AND2X2 AND2X2_5357 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n9696_), .Y(core__abc_22172_new_n9697_));
AND2X2 AND2X2_5358 ( .A(core_v0_reg_49_), .B(core_mi_reg_49_), .Y(core__abc_22172_new_n9699_));
AND2X2 AND2X2_5359 ( .A(core__abc_22172_new_n9700_), .B(core__abc_22172_new_n9698_), .Y(core__abc_22172_new_n9701_));
AND2X2 AND2X2_536 ( .A(_abc_19873_new_n1607_), .B(word2_reg_12_), .Y(_abc_19873_new_n1784_));
AND2X2 AND2X2_5360 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9701_), .Y(core__abc_22172_new_n9702_));
AND2X2 AND2X2_5361 ( .A(core__abc_22172_new_n9704_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9705_));
AND2X2 AND2X2_5362 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_49_), .Y(core__abc_22172_new_n9706_));
AND2X2 AND2X2_5363 ( .A(core__abc_22172_new_n9707_), .B(reset_n), .Y(core__0v0_reg_63_0__49_));
AND2X2 AND2X2_5364 ( .A(core__abc_22172_new_n5931_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9709_));
AND2X2 AND2X2_5365 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n9710_), .Y(core__abc_22172_new_n9711_));
AND2X2 AND2X2_5366 ( .A(core_v0_reg_50_), .B(core_mi_reg_50_), .Y(core__abc_22172_new_n9713_));
AND2X2 AND2X2_5367 ( .A(core__abc_22172_new_n9714_), .B(core__abc_22172_new_n9712_), .Y(core__abc_22172_new_n9715_));
AND2X2 AND2X2_5368 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9715_), .Y(core__abc_22172_new_n9716_));
AND2X2 AND2X2_5369 ( .A(core__abc_22172_new_n9718_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9719_));
AND2X2 AND2X2_537 ( .A(_abc_19873_new_n1785_), .B(reset_n), .Y(_0word2_reg_31_0__12_));
AND2X2 AND2X2_5370 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_50_), .Y(core__abc_22172_new_n9720_));
AND2X2 AND2X2_5371 ( .A(core__abc_22172_new_n9721_), .B(reset_n), .Y(core__0v0_reg_63_0__50_));
AND2X2 AND2X2_5372 ( .A(core__abc_22172_new_n5964_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9723_));
AND2X2 AND2X2_5373 ( .A(core_v0_reg_51_), .B(core_mi_reg_51_), .Y(core__abc_22172_new_n9725_));
AND2X2 AND2X2_5374 ( .A(core__abc_22172_new_n9726_), .B(core__abc_22172_new_n9724_), .Y(core__abc_22172_new_n9727_));
AND2X2 AND2X2_5375 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9727_), .Y(core__abc_22172_new_n9728_));
AND2X2 AND2X2_5376 ( .A(core__abc_22172_new_n9730_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9731_));
AND2X2 AND2X2_5377 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_51_), .Y(core__abc_22172_new_n9732_));
AND2X2 AND2X2_5378 ( .A(core__abc_22172_new_n9733_), .B(reset_n), .Y(core__0v0_reg_63_0__51_));
AND2X2 AND2X2_5379 ( .A(core__abc_22172_new_n6012_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9735_));
AND2X2 AND2X2_538 ( .A(core_siphash_valid_reg), .B(core_siphash_word_77_), .Y(_abc_19873_new_n1787_));
AND2X2 AND2X2_5380 ( .A(core__abc_22172_new_n3214_), .B(core_key_52_), .Y(core__abc_22172_new_n9736_));
AND2X2 AND2X2_5381 ( .A(core_v0_reg_52_), .B(core_mi_reg_52_), .Y(core__abc_22172_new_n9738_));
AND2X2 AND2X2_5382 ( .A(core__abc_22172_new_n9739_), .B(core__abc_22172_new_n9737_), .Y(core__abc_22172_new_n9740_));
AND2X2 AND2X2_5383 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9740_), .Y(core__abc_22172_new_n9741_));
AND2X2 AND2X2_5384 ( .A(core__abc_22172_new_n9743_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9744_));
AND2X2 AND2X2_5385 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_52_), .Y(core__abc_22172_new_n9745_));
AND2X2 AND2X2_5386 ( .A(core__abc_22172_new_n9746_), .B(reset_n), .Y(core__0v0_reg_63_0__52_));
AND2X2 AND2X2_5387 ( .A(core__abc_22172_new_n6042_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9748_));
AND2X2 AND2X2_5388 ( .A(core_v0_reg_53_), .B(core_mi_reg_53_), .Y(core__abc_22172_new_n9750_));
AND2X2 AND2X2_5389 ( .A(core__abc_22172_new_n9751_), .B(core__abc_22172_new_n9749_), .Y(core__abc_22172_new_n9752_));
AND2X2 AND2X2_539 ( .A(_abc_19873_new_n1607_), .B(word2_reg_13_), .Y(_abc_19873_new_n1788_));
AND2X2 AND2X2_5390 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9752_), .Y(core__abc_22172_new_n9753_));
AND2X2 AND2X2_5391 ( .A(core__abc_22172_new_n9755_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9756_));
AND2X2 AND2X2_5392 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_53_), .Y(core__abc_22172_new_n9757_));
AND2X2 AND2X2_5393 ( .A(core__abc_22172_new_n9758_), .B(reset_n), .Y(core__0v0_reg_63_0__53_));
AND2X2 AND2X2_5394 ( .A(core__abc_22172_new_n6086_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9760_));
AND2X2 AND2X2_5395 ( .A(core_v0_reg_54_), .B(core_mi_reg_54_), .Y(core__abc_22172_new_n9762_));
AND2X2 AND2X2_5396 ( .A(core__abc_22172_new_n9763_), .B(core__abc_22172_new_n9761_), .Y(core__abc_22172_new_n9764_));
AND2X2 AND2X2_5397 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9764_), .Y(core__abc_22172_new_n9765_));
AND2X2 AND2X2_5398 ( .A(core__abc_22172_new_n9767_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9768_));
AND2X2 AND2X2_5399 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_54_), .Y(core__abc_22172_new_n9769_));
AND2X2 AND2X2_54 ( .A(_abc_19873_new_n907_), .B(word1_reg_1_), .Y(_abc_19873_new_n946_));
AND2X2 AND2X2_540 ( .A(_abc_19873_new_n1789_), .B(reset_n), .Y(_0word2_reg_31_0__13_));
AND2X2 AND2X2_5400 ( .A(core__abc_22172_new_n9770_), .B(reset_n), .Y(core__0v0_reg_63_0__54_));
AND2X2 AND2X2_5401 ( .A(core__abc_22172_new_n6125_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9772_));
AND2X2 AND2X2_5402 ( .A(core_v0_reg_55_), .B(core_mi_reg_55_), .Y(core__abc_22172_new_n9774_));
AND2X2 AND2X2_5403 ( .A(core__abc_22172_new_n9775_), .B(core__abc_22172_new_n9773_), .Y(core__abc_22172_new_n9776_));
AND2X2 AND2X2_5404 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9776_), .Y(core__abc_22172_new_n9777_));
AND2X2 AND2X2_5405 ( .A(core__abc_22172_new_n9779_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9780_));
AND2X2 AND2X2_5406 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_55_), .Y(core__abc_22172_new_n9781_));
AND2X2 AND2X2_5407 ( .A(core__abc_22172_new_n9782_), .B(reset_n), .Y(core__0v0_reg_63_0__55_));
AND2X2 AND2X2_5408 ( .A(core__abc_22172_new_n6178_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9784_));
AND2X2 AND2X2_5409 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n9785_), .Y(core__abc_22172_new_n9786_));
AND2X2 AND2X2_541 ( .A(core_siphash_valid_reg), .B(core_siphash_word_78_), .Y(_abc_19873_new_n1791_));
AND2X2 AND2X2_5410 ( .A(core_v0_reg_56_), .B(core_mi_reg_56_), .Y(core__abc_22172_new_n9788_));
AND2X2 AND2X2_5411 ( .A(core__abc_22172_new_n9789_), .B(core__abc_22172_new_n9787_), .Y(core__abc_22172_new_n9790_));
AND2X2 AND2X2_5412 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9790_), .Y(core__abc_22172_new_n9791_));
AND2X2 AND2X2_5413 ( .A(core__abc_22172_new_n9793_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9794_));
AND2X2 AND2X2_5414 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_56_), .Y(core__abc_22172_new_n9795_));
AND2X2 AND2X2_5415 ( .A(core__abc_22172_new_n9796_), .B(reset_n), .Y(core__0v0_reg_63_0__56_));
AND2X2 AND2X2_5416 ( .A(core__abc_22172_new_n6208_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9798_));
AND2X2 AND2X2_5417 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n9799_), .Y(core__abc_22172_new_n9800_));
AND2X2 AND2X2_5418 ( .A(core_v0_reg_57_), .B(core_mi_reg_57_), .Y(core__abc_22172_new_n9802_));
AND2X2 AND2X2_5419 ( .A(core__abc_22172_new_n9803_), .B(core__abc_22172_new_n9801_), .Y(core__abc_22172_new_n9804_));
AND2X2 AND2X2_542 ( .A(_abc_19873_new_n1607_), .B(word2_reg_14_), .Y(_abc_19873_new_n1792_));
AND2X2 AND2X2_5420 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9804_), .Y(core__abc_22172_new_n9805_));
AND2X2 AND2X2_5421 ( .A(core__abc_22172_new_n9807_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9808_));
AND2X2 AND2X2_5422 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_57_), .Y(core__abc_22172_new_n9809_));
AND2X2 AND2X2_5423 ( .A(core__abc_22172_new_n9810_), .B(reset_n), .Y(core__0v0_reg_63_0__57_));
AND2X2 AND2X2_5424 ( .A(core__abc_22172_new_n6250_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9812_));
AND2X2 AND2X2_5425 ( .A(core__abc_22172_new_n3214_), .B(core_key_58_), .Y(core__abc_22172_new_n9813_));
AND2X2 AND2X2_5426 ( .A(core_v0_reg_58_), .B(core_mi_reg_58_), .Y(core__abc_22172_new_n9815_));
AND2X2 AND2X2_5427 ( .A(core__abc_22172_new_n9816_), .B(core__abc_22172_new_n9814_), .Y(core__abc_22172_new_n9817_));
AND2X2 AND2X2_5428 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9817_), .Y(core__abc_22172_new_n9818_));
AND2X2 AND2X2_5429 ( .A(core__abc_22172_new_n9820_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9821_));
AND2X2 AND2X2_543 ( .A(_abc_19873_new_n1793_), .B(reset_n), .Y(_0word2_reg_31_0__14_));
AND2X2 AND2X2_5430 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_58_), .Y(core__abc_22172_new_n9822_));
AND2X2 AND2X2_5431 ( .A(core__abc_22172_new_n9823_), .B(reset_n), .Y(core__0v0_reg_63_0__58_));
AND2X2 AND2X2_5432 ( .A(core__abc_22172_new_n6285_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9825_));
AND2X2 AND2X2_5433 ( .A(core__abc_22172_new_n3214_), .B(core_key_59_), .Y(core__abc_22172_new_n9826_));
AND2X2 AND2X2_5434 ( .A(core_v0_reg_59_), .B(core_mi_reg_59_), .Y(core__abc_22172_new_n9828_));
AND2X2 AND2X2_5435 ( .A(core__abc_22172_new_n9829_), .B(core__abc_22172_new_n9827_), .Y(core__abc_22172_new_n9830_));
AND2X2 AND2X2_5436 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9830_), .Y(core__abc_22172_new_n9831_));
AND2X2 AND2X2_5437 ( .A(core__abc_22172_new_n9833_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9834_));
AND2X2 AND2X2_5438 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_59_), .Y(core__abc_22172_new_n9835_));
AND2X2 AND2X2_5439 ( .A(core__abc_22172_new_n9836_), .B(reset_n), .Y(core__0v0_reg_63_0__59_));
AND2X2 AND2X2_544 ( .A(core_siphash_valid_reg), .B(core_siphash_word_79_), .Y(_abc_19873_new_n1795_));
AND2X2 AND2X2_5440 ( .A(core__abc_22172_new_n6335_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9838_));
AND2X2 AND2X2_5441 ( .A(core__abc_22172_new_n3214_), .B(core__abc_22172_new_n9839_), .Y(core__abc_22172_new_n9840_));
AND2X2 AND2X2_5442 ( .A(core_v0_reg_60_), .B(core_mi_reg_60_), .Y(core__abc_22172_new_n9842_));
AND2X2 AND2X2_5443 ( .A(core__abc_22172_new_n9843_), .B(core__abc_22172_new_n9841_), .Y(core__abc_22172_new_n9844_));
AND2X2 AND2X2_5444 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9844_), .Y(core__abc_22172_new_n9845_));
AND2X2 AND2X2_5445 ( .A(core__abc_22172_new_n9847_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9848_));
AND2X2 AND2X2_5446 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_60_), .Y(core__abc_22172_new_n9849_));
AND2X2 AND2X2_5447 ( .A(core__abc_22172_new_n9850_), .B(reset_n), .Y(core__0v0_reg_63_0__60_));
AND2X2 AND2X2_5448 ( .A(core__abc_22172_new_n6374_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9852_));
AND2X2 AND2X2_5449 ( .A(core_v0_reg_61_), .B(core_mi_reg_61_), .Y(core__abc_22172_new_n9854_));
AND2X2 AND2X2_545 ( .A(_abc_19873_new_n1607_), .B(word2_reg_15_), .Y(_abc_19873_new_n1796_));
AND2X2 AND2X2_5450 ( .A(core__abc_22172_new_n9855_), .B(core__abc_22172_new_n9853_), .Y(core__abc_22172_new_n9856_));
AND2X2 AND2X2_5451 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9856_), .Y(core__abc_22172_new_n9857_));
AND2X2 AND2X2_5452 ( .A(core__abc_22172_new_n9859_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9860_));
AND2X2 AND2X2_5453 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_61_), .Y(core__abc_22172_new_n9861_));
AND2X2 AND2X2_5454 ( .A(core__abc_22172_new_n9862_), .B(reset_n), .Y(core__0v0_reg_63_0__61_));
AND2X2 AND2X2_5455 ( .A(core__abc_22172_new_n6417_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9864_));
AND2X2 AND2X2_5456 ( .A(core_v0_reg_62_), .B(core_mi_reg_62_), .Y(core__abc_22172_new_n9866_));
AND2X2 AND2X2_5457 ( .A(core__abc_22172_new_n9867_), .B(core__abc_22172_new_n9865_), .Y(core__abc_22172_new_n9868_));
AND2X2 AND2X2_5458 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9868_), .Y(core__abc_22172_new_n9869_));
AND2X2 AND2X2_5459 ( .A(core__abc_22172_new_n9871_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9872_));
AND2X2 AND2X2_546 ( .A(_abc_19873_new_n1797_), .B(reset_n), .Y(_0word2_reg_31_0__15_));
AND2X2 AND2X2_5460 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_62_), .Y(core__abc_22172_new_n9873_));
AND2X2 AND2X2_5461 ( .A(core__abc_22172_new_n9874_), .B(reset_n), .Y(core__0v0_reg_63_0__62_));
AND2X2 AND2X2_5462 ( .A(core__abc_22172_new_n6448_), .B(core__abc_22172_new_n3205_), .Y(core__abc_22172_new_n9876_));
AND2X2 AND2X2_5463 ( .A(core_v0_reg_63_), .B(core_mi_reg_63_), .Y(core__abc_22172_new_n9878_));
AND2X2 AND2X2_5464 ( .A(core__abc_22172_new_n9879_), .B(core__abc_22172_new_n9877_), .Y(core__abc_22172_new_n9880_));
AND2X2 AND2X2_5465 ( .A(core__abc_22172_new_n9080_), .B(core__abc_22172_new_n9880_), .Y(core__abc_22172_new_n9881_));
AND2X2 AND2X2_5466 ( .A(core__abc_22172_new_n9883_), .B(core__abc_22172_new_n4187_), .Y(core__abc_22172_new_n9884_));
AND2X2 AND2X2_5467 ( .A(core__abc_22172_new_n9083_), .B(core_v0_reg_63_), .Y(core__abc_22172_new_n9885_));
AND2X2 AND2X2_5468 ( .A(core__abc_22172_new_n9886_), .B(reset_n), .Y(core__0v0_reg_63_0__63_));
AND2X2 AND2X2_5469 ( .A(core__abc_22172_new_n1222_), .B(reset_n), .Y(core__abc_22172_new_n9888_));
AND2X2 AND2X2_547 ( .A(core_siphash_valid_reg), .B(core_siphash_word_80_), .Y(_abc_19873_new_n1799_));
AND2X2 AND2X2_5470 ( .A(core__abc_22172_new_n9888_), .B(core__abc_22172_new_n1212_), .Y(core__abc_15204_auto_fsm_map_cc_118_implement_pattern_cache_1474));
AND2X2 AND2X2_5471 ( .A(core__abc_22172_new_n9888_), .B(core__abc_22172_new_n1165_), .Y(core__abc_22172_new_n9890_));
AND2X2 AND2X2_5472 ( .A(core__abc_22172_new_n9890_), .B(core_siphash_ctrl_reg_6_), .Y(core__abc_22172_new_n9891_));
AND2X2 AND2X2_5473 ( .A(core__abc_22172_new_n9891_), .B(core__abc_22172_new_n6870_), .Y(core__abc_15204_auto_fsm_map_cc_118_implement_pattern_cache_1470));
AND2X2 AND2X2_5474 ( .A(core__abc_22172_new_n9891_), .B(core_long), .Y(core__abc_15204_auto_fsm_map_cc_118_implement_pattern_cache_1496));
AND2X2 AND2X2_5475 ( .A(core__abc_22172_new_n9890_), .B(core_siphash_ctrl_reg_3_), .Y(core__abc_15204_auto_fsm_map_cc_118_implement_pattern_cache_1509));
AND2X2 AND2X2_5476 ( .A(core__abc_22172_new_n9896_), .B(core_siphash_valid_reg), .Y(core__abc_22172_new_n9897_));
AND2X2 AND2X2_5477 ( .A(core__abc_22172_new_n9898_), .B(reset_n), .Y(core__0siphash_valid_reg_0_0_));
AND2X2 AND2X2_548 ( .A(_abc_19873_new_n1607_), .B(word2_reg_16_), .Y(_abc_19873_new_n1800_));
AND2X2 AND2X2_549 ( .A(_abc_19873_new_n1801_), .B(reset_n), .Y(_0word2_reg_31_0__16_));
AND2X2 AND2X2_55 ( .A(_abc_19873_new_n912_), .B(word3_reg_1_), .Y(_abc_19873_new_n950_));
AND2X2 AND2X2_550 ( .A(core_siphash_valid_reg), .B(core_siphash_word_81_), .Y(_abc_19873_new_n1803_));
AND2X2 AND2X2_551 ( .A(_abc_19873_new_n1607_), .B(word2_reg_17_), .Y(_abc_19873_new_n1804_));
AND2X2 AND2X2_552 ( .A(_abc_19873_new_n1805_), .B(reset_n), .Y(_0word2_reg_31_0__17_));
AND2X2 AND2X2_553 ( .A(core_siphash_valid_reg), .B(core_siphash_word_82_), .Y(_abc_19873_new_n1807_));
AND2X2 AND2X2_554 ( .A(_abc_19873_new_n1607_), .B(word2_reg_18_), .Y(_abc_19873_new_n1808_));
AND2X2 AND2X2_555 ( .A(_abc_19873_new_n1809_), .B(reset_n), .Y(_0word2_reg_31_0__18_));
AND2X2 AND2X2_556 ( .A(core_siphash_valid_reg), .B(core_siphash_word_83_), .Y(_abc_19873_new_n1811_));
AND2X2 AND2X2_557 ( .A(_abc_19873_new_n1607_), .B(word2_reg_19_), .Y(_abc_19873_new_n1812_));
AND2X2 AND2X2_558 ( .A(_abc_19873_new_n1813_), .B(reset_n), .Y(_0word2_reg_31_0__19_));
AND2X2 AND2X2_559 ( .A(core_siphash_valid_reg), .B(core_siphash_word_84_), .Y(_abc_19873_new_n1815_));
AND2X2 AND2X2_56 ( .A(_abc_19873_new_n916_), .B(core_key_65_), .Y(_abc_19873_new_n951_));
AND2X2 AND2X2_560 ( .A(_abc_19873_new_n1607_), .B(word2_reg_20_), .Y(_abc_19873_new_n1816_));
AND2X2 AND2X2_561 ( .A(_abc_19873_new_n1817_), .B(reset_n), .Y(_0word2_reg_31_0__20_));
AND2X2 AND2X2_562 ( .A(core_siphash_valid_reg), .B(core_siphash_word_85_), .Y(_abc_19873_new_n1819_));
AND2X2 AND2X2_563 ( .A(_abc_19873_new_n1607_), .B(word2_reg_21_), .Y(_abc_19873_new_n1820_));
AND2X2 AND2X2_564 ( .A(_abc_19873_new_n1821_), .B(reset_n), .Y(_0word2_reg_31_0__21_));
AND2X2 AND2X2_565 ( .A(core_siphash_valid_reg), .B(core_siphash_word_86_), .Y(_abc_19873_new_n1823_));
AND2X2 AND2X2_566 ( .A(_abc_19873_new_n1607_), .B(word2_reg_22_), .Y(_abc_19873_new_n1824_));
AND2X2 AND2X2_567 ( .A(_abc_19873_new_n1825_), .B(reset_n), .Y(_0word2_reg_31_0__22_));
AND2X2 AND2X2_568 ( .A(core_siphash_valid_reg), .B(core_siphash_word_87_), .Y(_abc_19873_new_n1827_));
AND2X2 AND2X2_569 ( .A(_abc_19873_new_n1607_), .B(word2_reg_23_), .Y(_abc_19873_new_n1828_));
AND2X2 AND2X2_57 ( .A(_abc_19873_new_n919_), .B(core_mi_33_), .Y(_abc_19873_new_n952_));
AND2X2 AND2X2_570 ( .A(_abc_19873_new_n1829_), .B(reset_n), .Y(_0word2_reg_31_0__23_));
AND2X2 AND2X2_571 ( .A(core_siphash_valid_reg), .B(core_siphash_word_88_), .Y(_abc_19873_new_n1831_));
AND2X2 AND2X2_572 ( .A(_abc_19873_new_n1607_), .B(word2_reg_24_), .Y(_abc_19873_new_n1832_));
AND2X2 AND2X2_573 ( .A(_abc_19873_new_n1833_), .B(reset_n), .Y(_0word2_reg_31_0__24_));
AND2X2 AND2X2_574 ( .A(core_siphash_valid_reg), .B(core_siphash_word_89_), .Y(_abc_19873_new_n1835_));
AND2X2 AND2X2_575 ( .A(_abc_19873_new_n1607_), .B(word2_reg_25_), .Y(_abc_19873_new_n1836_));
AND2X2 AND2X2_576 ( .A(_abc_19873_new_n1837_), .B(reset_n), .Y(_0word2_reg_31_0__25_));
AND2X2 AND2X2_577 ( .A(core_siphash_valid_reg), .B(core_siphash_word_90_), .Y(_abc_19873_new_n1839_));
AND2X2 AND2X2_578 ( .A(_abc_19873_new_n1607_), .B(word2_reg_26_), .Y(_abc_19873_new_n1840_));
AND2X2 AND2X2_579 ( .A(_abc_19873_new_n1841_), .B(reset_n), .Y(_0word2_reg_31_0__26_));
AND2X2 AND2X2_58 ( .A(_abc_19873_new_n923_), .B(core_siphash_valid_reg), .Y(_abc_19873_new_n955_));
AND2X2 AND2X2_580 ( .A(core_siphash_valid_reg), .B(core_siphash_word_91_), .Y(_abc_19873_new_n1843_));
AND2X2 AND2X2_581 ( .A(_abc_19873_new_n1607_), .B(word2_reg_27_), .Y(_abc_19873_new_n1844_));
AND2X2 AND2X2_582 ( .A(_abc_19873_new_n1845_), .B(reset_n), .Y(_0word2_reg_31_0__27_));
AND2X2 AND2X2_583 ( .A(core_siphash_valid_reg), .B(core_siphash_word_92_), .Y(_abc_19873_new_n1847_));
AND2X2 AND2X2_584 ( .A(_abc_19873_new_n1607_), .B(word2_reg_28_), .Y(_abc_19873_new_n1848_));
AND2X2 AND2X2_585 ( .A(_abc_19873_new_n1849_), .B(reset_n), .Y(_0word2_reg_31_0__28_));
AND2X2 AND2X2_586 ( .A(core_siphash_valid_reg), .B(core_siphash_word_93_), .Y(_abc_19873_new_n1851_));
AND2X2 AND2X2_587 ( .A(_abc_19873_new_n1607_), .B(word2_reg_29_), .Y(_abc_19873_new_n1852_));
AND2X2 AND2X2_588 ( .A(_abc_19873_new_n1853_), .B(reset_n), .Y(_0word2_reg_31_0__29_));
AND2X2 AND2X2_589 ( .A(core_siphash_valid_reg), .B(core_siphash_word_94_), .Y(_abc_19873_new_n1855_));
AND2X2 AND2X2_59 ( .A(_abc_19873_new_n925_), .B(word2_reg_1_), .Y(_abc_19873_new_n956_));
AND2X2 AND2X2_590 ( .A(_abc_19873_new_n1607_), .B(word2_reg_30_), .Y(_abc_19873_new_n1856_));
AND2X2 AND2X2_591 ( .A(_abc_19873_new_n1857_), .B(reset_n), .Y(_0word2_reg_31_0__30_));
AND2X2 AND2X2_592 ( .A(core_siphash_valid_reg), .B(core_siphash_word_95_), .Y(_abc_19873_new_n1859_));
AND2X2 AND2X2_593 ( .A(_abc_19873_new_n1607_), .B(word2_reg_31_), .Y(_abc_19873_new_n1860_));
AND2X2 AND2X2_594 ( .A(_abc_19873_new_n1861_), .B(reset_n), .Y(_0word2_reg_31_0__31_));
AND2X2 AND2X2_595 ( .A(core_siphash_valid_reg), .B(core_siphash_word_32_), .Y(_abc_19873_new_n1863_));
AND2X2 AND2X2_596 ( .A(_abc_19873_new_n1607_), .B(word1_reg_0_), .Y(_abc_19873_new_n1864_));
AND2X2 AND2X2_597 ( .A(_abc_19873_new_n1865_), .B(reset_n), .Y(_0word1_reg_31_0__0_));
AND2X2 AND2X2_598 ( .A(core_siphash_valid_reg), .B(core_siphash_word_33_), .Y(_abc_19873_new_n1867_));
AND2X2 AND2X2_599 ( .A(_abc_19873_new_n1607_), .B(word1_reg_1_), .Y(_abc_19873_new_n1868_));
AND2X2 AND2X2_6 ( .A(_abc_19873_new_n879_), .B(_abc_19873_new_n876_), .Y(_abc_19873_new_n880_));
AND2X2 AND2X2_60 ( .A(_abc_19873_new_n928_), .B(core_key_33_), .Y(_abc_19873_new_n958_));
AND2X2 AND2X2_600 ( .A(_abc_19873_new_n1869_), .B(reset_n), .Y(_0word1_reg_31_0__1_));
AND2X2 AND2X2_601 ( .A(core_siphash_valid_reg), .B(core_siphash_word_34_), .Y(_abc_19873_new_n1871_));
AND2X2 AND2X2_602 ( .A(_abc_19873_new_n1607_), .B(word1_reg_2_), .Y(_abc_19873_new_n1872_));
AND2X2 AND2X2_603 ( .A(_abc_19873_new_n1873_), .B(reset_n), .Y(_0word1_reg_31_0__2_));
AND2X2 AND2X2_604 ( .A(core_siphash_valid_reg), .B(core_siphash_word_35_), .Y(_abc_19873_new_n1875_));
AND2X2 AND2X2_605 ( .A(_abc_19873_new_n1607_), .B(word1_reg_3_), .Y(_abc_19873_new_n1876_));
AND2X2 AND2X2_606 ( .A(_abc_19873_new_n1877_), .B(reset_n), .Y(_0word1_reg_31_0__3_));
AND2X2 AND2X2_607 ( .A(core_siphash_valid_reg), .B(core_siphash_word_36_), .Y(_abc_19873_new_n1879_));
AND2X2 AND2X2_608 ( .A(_abc_19873_new_n1607_), .B(word1_reg_4_), .Y(_abc_19873_new_n1880_));
AND2X2 AND2X2_609 ( .A(_abc_19873_new_n1881_), .B(reset_n), .Y(_0word1_reg_31_0__4_));
AND2X2 AND2X2_61 ( .A(_abc_19873_new_n930_), .B(word0_reg_1_), .Y(_abc_19873_new_n959_));
AND2X2 AND2X2_610 ( .A(core_siphash_valid_reg), .B(core_siphash_word_37_), .Y(_abc_19873_new_n1883_));
AND2X2 AND2X2_611 ( .A(_abc_19873_new_n1607_), .B(word1_reg_5_), .Y(_abc_19873_new_n1884_));
AND2X2 AND2X2_612 ( .A(_abc_19873_new_n1885_), .B(reset_n), .Y(_0word1_reg_31_0__5_));
AND2X2 AND2X2_613 ( .A(core_siphash_valid_reg), .B(core_siphash_word_38_), .Y(_abc_19873_new_n1887_));
AND2X2 AND2X2_614 ( .A(_abc_19873_new_n1607_), .B(word1_reg_6_), .Y(_abc_19873_new_n1888_));
AND2X2 AND2X2_615 ( .A(_abc_19873_new_n1889_), .B(reset_n), .Y(_0word1_reg_31_0__6_));
AND2X2 AND2X2_616 ( .A(core_siphash_valid_reg), .B(core_siphash_word_39_), .Y(_abc_19873_new_n1891_));
AND2X2 AND2X2_617 ( .A(_abc_19873_new_n1607_), .B(word1_reg_7_), .Y(_abc_19873_new_n1892_));
AND2X2 AND2X2_618 ( .A(_abc_19873_new_n1893_), .B(reset_n), .Y(_0word1_reg_31_0__7_));
AND2X2 AND2X2_619 ( .A(core_siphash_valid_reg), .B(core_siphash_word_40_), .Y(_abc_19873_new_n1895_));
AND2X2 AND2X2_62 ( .A(_abc_19873_new_n963_), .B(_abc_19873_new_n937_), .Y(\read_data[1] ));
AND2X2 AND2X2_620 ( .A(_abc_19873_new_n1607_), .B(word1_reg_8_), .Y(_abc_19873_new_n1896_));
AND2X2 AND2X2_621 ( .A(_abc_19873_new_n1897_), .B(reset_n), .Y(_0word1_reg_31_0__8_));
AND2X2 AND2X2_622 ( .A(core_siphash_valid_reg), .B(core_siphash_word_41_), .Y(_abc_19873_new_n1899_));
AND2X2 AND2X2_623 ( .A(_abc_19873_new_n1607_), .B(word1_reg_9_), .Y(_abc_19873_new_n1900_));
AND2X2 AND2X2_624 ( .A(_abc_19873_new_n1901_), .B(reset_n), .Y(_0word1_reg_31_0__9_));
AND2X2 AND2X2_625 ( .A(core_siphash_valid_reg), .B(core_siphash_word_42_), .Y(_abc_19873_new_n1903_));
AND2X2 AND2X2_626 ( .A(_abc_19873_new_n1607_), .B(word1_reg_10_), .Y(_abc_19873_new_n1904_));
AND2X2 AND2X2_627 ( .A(_abc_19873_new_n1905_), .B(reset_n), .Y(_0word1_reg_31_0__10_));
AND2X2 AND2X2_628 ( .A(core_siphash_valid_reg), .B(core_siphash_word_43_), .Y(_abc_19873_new_n1907_));
AND2X2 AND2X2_629 ( .A(_abc_19873_new_n1607_), .B(word1_reg_11_), .Y(_abc_19873_new_n1908_));
AND2X2 AND2X2_63 ( .A(_abc_19873_new_n925_), .B(word2_reg_2_), .Y(_abc_19873_new_n965_));
AND2X2 AND2X2_630 ( .A(_abc_19873_new_n1909_), .B(reset_n), .Y(_0word1_reg_31_0__11_));
AND2X2 AND2X2_631 ( .A(core_siphash_valid_reg), .B(core_siphash_word_44_), .Y(_abc_19873_new_n1911_));
AND2X2 AND2X2_632 ( .A(_abc_19873_new_n1607_), .B(word1_reg_12_), .Y(_abc_19873_new_n1912_));
AND2X2 AND2X2_633 ( .A(_abc_19873_new_n1913_), .B(reset_n), .Y(_0word1_reg_31_0__12_));
AND2X2 AND2X2_634 ( .A(core_siphash_valid_reg), .B(core_siphash_word_45_), .Y(_abc_19873_new_n1915_));
AND2X2 AND2X2_635 ( .A(_abc_19873_new_n1607_), .B(word1_reg_13_), .Y(_abc_19873_new_n1916_));
AND2X2 AND2X2_636 ( .A(_abc_19873_new_n1917_), .B(reset_n), .Y(_0word1_reg_31_0__13_));
AND2X2 AND2X2_637 ( .A(core_siphash_valid_reg), .B(core_siphash_word_46_), .Y(_abc_19873_new_n1919_));
AND2X2 AND2X2_638 ( .A(_abc_19873_new_n1607_), .B(word1_reg_14_), .Y(_abc_19873_new_n1920_));
AND2X2 AND2X2_639 ( .A(_abc_19873_new_n1921_), .B(reset_n), .Y(_0word1_reg_31_0__14_));
AND2X2 AND2X2_64 ( .A(_abc_19873_new_n916_), .B(core_key_66_), .Y(_abc_19873_new_n966_));
AND2X2 AND2X2_640 ( .A(core_siphash_valid_reg), .B(core_siphash_word_47_), .Y(_abc_19873_new_n1923_));
AND2X2 AND2X2_641 ( .A(_abc_19873_new_n1607_), .B(word1_reg_15_), .Y(_abc_19873_new_n1924_));
AND2X2 AND2X2_642 ( .A(_abc_19873_new_n1925_), .B(reset_n), .Y(_0word1_reg_31_0__15_));
AND2X2 AND2X2_643 ( .A(core_siphash_valid_reg), .B(core_siphash_word_48_), .Y(_abc_19873_new_n1927_));
AND2X2 AND2X2_644 ( .A(_abc_19873_new_n1607_), .B(word1_reg_16_), .Y(_abc_19873_new_n1928_));
AND2X2 AND2X2_645 ( .A(_abc_19873_new_n1929_), .B(reset_n), .Y(_0word1_reg_31_0__16_));
AND2X2 AND2X2_646 ( .A(core_siphash_valid_reg), .B(core_siphash_word_49_), .Y(_abc_19873_new_n1931_));
AND2X2 AND2X2_647 ( .A(_abc_19873_new_n1607_), .B(word1_reg_17_), .Y(_abc_19873_new_n1932_));
AND2X2 AND2X2_648 ( .A(_abc_19873_new_n1933_), .B(reset_n), .Y(_0word1_reg_31_0__17_));
AND2X2 AND2X2_649 ( .A(core_siphash_valid_reg), .B(core_siphash_word_50_), .Y(_abc_19873_new_n1935_));
AND2X2 AND2X2_65 ( .A(_abc_19873_new_n881_), .B(core_key_98_), .Y(_abc_19873_new_n967_));
AND2X2 AND2X2_650 ( .A(_abc_19873_new_n1607_), .B(word1_reg_18_), .Y(_abc_19873_new_n1936_));
AND2X2 AND2X2_651 ( .A(_abc_19873_new_n1937_), .B(reset_n), .Y(_0word1_reg_31_0__18_));
AND2X2 AND2X2_652 ( .A(core_siphash_valid_reg), .B(core_siphash_word_51_), .Y(_abc_19873_new_n1939_));
AND2X2 AND2X2_653 ( .A(_abc_19873_new_n1607_), .B(word1_reg_19_), .Y(_abc_19873_new_n1940_));
AND2X2 AND2X2_654 ( .A(_abc_19873_new_n1941_), .B(reset_n), .Y(_0word1_reg_31_0__19_));
AND2X2 AND2X2_655 ( .A(core_siphash_valid_reg), .B(core_siphash_word_52_), .Y(_abc_19873_new_n1943_));
AND2X2 AND2X2_656 ( .A(_abc_19873_new_n1607_), .B(word1_reg_20_), .Y(_abc_19873_new_n1944_));
AND2X2 AND2X2_657 ( .A(_abc_19873_new_n1945_), .B(reset_n), .Y(_0word1_reg_31_0__20_));
AND2X2 AND2X2_658 ( .A(core_siphash_valid_reg), .B(core_siphash_word_53_), .Y(_abc_19873_new_n1947_));
AND2X2 AND2X2_659 ( .A(_abc_19873_new_n1607_), .B(word1_reg_21_), .Y(_abc_19873_new_n1948_));
AND2X2 AND2X2_66 ( .A(_abc_19873_new_n928_), .B(core_key_34_), .Y(_abc_19873_new_n969_));
AND2X2 AND2X2_660 ( .A(_abc_19873_new_n1949_), .B(reset_n), .Y(_0word1_reg_31_0__21_));
AND2X2 AND2X2_661 ( .A(core_siphash_valid_reg), .B(core_siphash_word_54_), .Y(_abc_19873_new_n1951_));
AND2X2 AND2X2_662 ( .A(_abc_19873_new_n1607_), .B(word1_reg_22_), .Y(_abc_19873_new_n1952_));
AND2X2 AND2X2_663 ( .A(_abc_19873_new_n1953_), .B(reset_n), .Y(_0word1_reg_31_0__22_));
AND2X2 AND2X2_664 ( .A(core_siphash_valid_reg), .B(core_siphash_word_55_), .Y(_abc_19873_new_n1955_));
AND2X2 AND2X2_665 ( .A(_abc_19873_new_n1607_), .B(word1_reg_23_), .Y(_abc_19873_new_n1956_));
AND2X2 AND2X2_666 ( .A(_abc_19873_new_n1957_), .B(reset_n), .Y(_0word1_reg_31_0__23_));
AND2X2 AND2X2_667 ( .A(core_siphash_valid_reg), .B(core_siphash_word_56_), .Y(_abc_19873_new_n1959_));
AND2X2 AND2X2_668 ( .A(_abc_19873_new_n1607_), .B(word1_reg_24_), .Y(_abc_19873_new_n1960_));
AND2X2 AND2X2_669 ( .A(_abc_19873_new_n1961_), .B(reset_n), .Y(_0word1_reg_31_0__24_));
AND2X2 AND2X2_67 ( .A(_abc_19873_new_n901_), .B(core_key_2_), .Y(_abc_19873_new_n970_));
AND2X2 AND2X2_670 ( .A(core_siphash_valid_reg), .B(core_siphash_word_57_), .Y(_abc_19873_new_n1963_));
AND2X2 AND2X2_671 ( .A(_abc_19873_new_n1607_), .B(word1_reg_25_), .Y(_abc_19873_new_n1964_));
AND2X2 AND2X2_672 ( .A(_abc_19873_new_n1965_), .B(reset_n), .Y(_0word1_reg_31_0__25_));
AND2X2 AND2X2_673 ( .A(core_siphash_valid_reg), .B(core_siphash_word_58_), .Y(_abc_19873_new_n1967_));
AND2X2 AND2X2_674 ( .A(_abc_19873_new_n1607_), .B(word1_reg_26_), .Y(_abc_19873_new_n1968_));
AND2X2 AND2X2_675 ( .A(_abc_19873_new_n1969_), .B(reset_n), .Y(_0word1_reg_31_0__26_));
AND2X2 AND2X2_676 ( .A(core_siphash_valid_reg), .B(core_siphash_word_59_), .Y(_abc_19873_new_n1971_));
AND2X2 AND2X2_677 ( .A(_abc_19873_new_n1607_), .B(word1_reg_27_), .Y(_abc_19873_new_n1972_));
AND2X2 AND2X2_678 ( .A(_abc_19873_new_n1973_), .B(reset_n), .Y(_0word1_reg_31_0__27_));
AND2X2 AND2X2_679 ( .A(core_siphash_valid_reg), .B(core_siphash_word_60_), .Y(_abc_19873_new_n1975_));
AND2X2 AND2X2_68 ( .A(_abc_19873_new_n930_), .B(word0_reg_2_), .Y(_abc_19873_new_n974_));
AND2X2 AND2X2_680 ( .A(_abc_19873_new_n1607_), .B(word1_reg_28_), .Y(_abc_19873_new_n1976_));
AND2X2 AND2X2_681 ( .A(_abc_19873_new_n1977_), .B(reset_n), .Y(_0word1_reg_31_0__28_));
AND2X2 AND2X2_682 ( .A(core_siphash_valid_reg), .B(core_siphash_word_61_), .Y(_abc_19873_new_n1979_));
AND2X2 AND2X2_683 ( .A(_abc_19873_new_n1607_), .B(word1_reg_29_), .Y(_abc_19873_new_n1980_));
AND2X2 AND2X2_684 ( .A(_abc_19873_new_n1981_), .B(reset_n), .Y(_0word1_reg_31_0__29_));
AND2X2 AND2X2_685 ( .A(core_siphash_valid_reg), .B(core_siphash_word_62_), .Y(_abc_19873_new_n1983_));
AND2X2 AND2X2_686 ( .A(_abc_19873_new_n1607_), .B(word1_reg_30_), .Y(_abc_19873_new_n1984_));
AND2X2 AND2X2_687 ( .A(_abc_19873_new_n1985_), .B(reset_n), .Y(_0word1_reg_31_0__30_));
AND2X2 AND2X2_688 ( .A(core_siphash_valid_reg), .B(core_siphash_word_63_), .Y(_abc_19873_new_n1987_));
AND2X2 AND2X2_689 ( .A(_abc_19873_new_n1607_), .B(word1_reg_31_), .Y(_abc_19873_new_n1988_));
AND2X2 AND2X2_69 ( .A(_abc_19873_new_n907_), .B(word1_reg_2_), .Y(_abc_19873_new_n975_));
AND2X2 AND2X2_690 ( .A(_abc_19873_new_n1989_), .B(reset_n), .Y(_0word1_reg_31_0__31_));
AND2X2 AND2X2_691 ( .A(core_siphash_valid_reg), .B(core_siphash_word_0_), .Y(_abc_19873_new_n1991_));
AND2X2 AND2X2_692 ( .A(_abc_19873_new_n1607_), .B(word0_reg_0_), .Y(_abc_19873_new_n1992_));
AND2X2 AND2X2_693 ( .A(_abc_19873_new_n1993_), .B(reset_n), .Y(_0word0_reg_31_0__0_));
AND2X2 AND2X2_694 ( .A(core_siphash_valid_reg), .B(core_siphash_word_1_), .Y(_abc_19873_new_n1995_));
AND2X2 AND2X2_695 ( .A(_abc_19873_new_n1607_), .B(word0_reg_1_), .Y(_abc_19873_new_n1996_));
AND2X2 AND2X2_696 ( .A(_abc_19873_new_n1997_), .B(reset_n), .Y(_0word0_reg_31_0__1_));
AND2X2 AND2X2_697 ( .A(core_siphash_valid_reg), .B(core_siphash_word_2_), .Y(_abc_19873_new_n1999_));
AND2X2 AND2X2_698 ( .A(_abc_19873_new_n1607_), .B(word0_reg_2_), .Y(_abc_19873_new_n2000_));
AND2X2 AND2X2_699 ( .A(_abc_19873_new_n2001_), .B(reset_n), .Y(_0word0_reg_31_0__2_));
AND2X2 AND2X2_7 ( .A(_abc_19873_new_n875_), .B(_abc_19873_new_n880_), .Y(_abc_19873_new_n881_));
AND2X2 AND2X2_70 ( .A(_abc_19873_new_n912_), .B(word3_reg_2_), .Y(_abc_19873_new_n977_));
AND2X2 AND2X2_700 ( .A(core_siphash_valid_reg), .B(core_siphash_word_3_), .Y(_abc_19873_new_n2003_));
AND2X2 AND2X2_701 ( .A(_abc_19873_new_n1607_), .B(word0_reg_3_), .Y(_abc_19873_new_n2004_));
AND2X2 AND2X2_702 ( .A(_abc_19873_new_n2005_), .B(reset_n), .Y(_0word0_reg_31_0__3_));
AND2X2 AND2X2_703 ( .A(core_siphash_valid_reg), .B(core_siphash_word_4_), .Y(_abc_19873_new_n2007_));
AND2X2 AND2X2_704 ( .A(_abc_19873_new_n1607_), .B(word0_reg_4_), .Y(_abc_19873_new_n2008_));
AND2X2 AND2X2_705 ( .A(_abc_19873_new_n2009_), .B(reset_n), .Y(_0word0_reg_31_0__4_));
AND2X2 AND2X2_706 ( .A(core_siphash_valid_reg), .B(core_siphash_word_5_), .Y(_abc_19873_new_n2011_));
AND2X2 AND2X2_707 ( .A(_abc_19873_new_n1607_), .B(word0_reg_5_), .Y(_abc_19873_new_n2012_));
AND2X2 AND2X2_708 ( .A(_abc_19873_new_n2013_), .B(reset_n), .Y(_0word0_reg_31_0__5_));
AND2X2 AND2X2_709 ( .A(core_siphash_valid_reg), .B(core_siphash_word_6_), .Y(_abc_19873_new_n2015_));
AND2X2 AND2X2_71 ( .A(_abc_19873_new_n919_), .B(core_mi_34_), .Y(_abc_19873_new_n979_));
AND2X2 AND2X2_710 ( .A(_abc_19873_new_n1607_), .B(word0_reg_6_), .Y(_abc_19873_new_n2016_));
AND2X2 AND2X2_711 ( .A(_abc_19873_new_n2017_), .B(reset_n), .Y(_0word0_reg_31_0__6_));
AND2X2 AND2X2_712 ( .A(core_siphash_valid_reg), .B(core_siphash_word_7_), .Y(_abc_19873_new_n2019_));
AND2X2 AND2X2_713 ( .A(_abc_19873_new_n1607_), .B(word0_reg_7_), .Y(_abc_19873_new_n2020_));
AND2X2 AND2X2_714 ( .A(_abc_19873_new_n2021_), .B(reset_n), .Y(_0word0_reg_31_0__7_));
AND2X2 AND2X2_715 ( .A(core_siphash_valid_reg), .B(core_siphash_word_8_), .Y(_abc_19873_new_n2023_));
AND2X2 AND2X2_716 ( .A(_abc_19873_new_n1607_), .B(word0_reg_8_), .Y(_abc_19873_new_n2024_));
AND2X2 AND2X2_717 ( .A(_abc_19873_new_n2025_), .B(reset_n), .Y(_0word0_reg_31_0__8_));
AND2X2 AND2X2_718 ( .A(core_siphash_valid_reg), .B(core_siphash_word_9_), .Y(_abc_19873_new_n2027_));
AND2X2 AND2X2_719 ( .A(_abc_19873_new_n1607_), .B(word0_reg_9_), .Y(_abc_19873_new_n2028_));
AND2X2 AND2X2_72 ( .A(_abc_19873_new_n888_), .B(core_mi_2_), .Y(_abc_19873_new_n980_));
AND2X2 AND2X2_720 ( .A(_abc_19873_new_n2029_), .B(reset_n), .Y(_0word0_reg_31_0__9_));
AND2X2 AND2X2_721 ( .A(core_siphash_valid_reg), .B(core_siphash_word_10_), .Y(_abc_19873_new_n2031_));
AND2X2 AND2X2_722 ( .A(_abc_19873_new_n1607_), .B(word0_reg_10_), .Y(_abc_19873_new_n2032_));
AND2X2 AND2X2_723 ( .A(_abc_19873_new_n2033_), .B(reset_n), .Y(_0word0_reg_31_0__10_));
AND2X2 AND2X2_724 ( .A(core_siphash_valid_reg), .B(core_siphash_word_11_), .Y(_abc_19873_new_n2035_));
AND2X2 AND2X2_725 ( .A(_abc_19873_new_n1607_), .B(word0_reg_11_), .Y(_abc_19873_new_n2036_));
AND2X2 AND2X2_726 ( .A(_abc_19873_new_n2037_), .B(reset_n), .Y(_0word0_reg_31_0__11_));
AND2X2 AND2X2_727 ( .A(core_siphash_valid_reg), .B(core_siphash_word_12_), .Y(_abc_19873_new_n2039_));
AND2X2 AND2X2_728 ( .A(_abc_19873_new_n1607_), .B(word0_reg_12_), .Y(_abc_19873_new_n2040_));
AND2X2 AND2X2_729 ( .A(_abc_19873_new_n2041_), .B(reset_n), .Y(_0word0_reg_31_0__12_));
AND2X2 AND2X2_73 ( .A(_abc_19873_new_n897_), .B(core_compression_rounds_2_), .Y(_abc_19873_new_n982_));
AND2X2 AND2X2_730 ( .A(core_siphash_valid_reg), .B(core_siphash_word_13_), .Y(_abc_19873_new_n2043_));
AND2X2 AND2X2_731 ( .A(_abc_19873_new_n1607_), .B(word0_reg_13_), .Y(_abc_19873_new_n2044_));
AND2X2 AND2X2_732 ( .A(_abc_19873_new_n2045_), .B(reset_n), .Y(_0word0_reg_31_0__13_));
AND2X2 AND2X2_733 ( .A(core_siphash_valid_reg), .B(core_siphash_word_14_), .Y(_abc_19873_new_n2047_));
AND2X2 AND2X2_734 ( .A(_abc_19873_new_n1607_), .B(word0_reg_14_), .Y(_abc_19873_new_n2048_));
AND2X2 AND2X2_735 ( .A(_abc_19873_new_n2049_), .B(reset_n), .Y(_0word0_reg_31_0__14_));
AND2X2 AND2X2_736 ( .A(core_siphash_valid_reg), .B(core_siphash_word_15_), .Y(_abc_19873_new_n2051_));
AND2X2 AND2X2_737 ( .A(_abc_19873_new_n1607_), .B(word0_reg_15_), .Y(_abc_19873_new_n2052_));
AND2X2 AND2X2_738 ( .A(_abc_19873_new_n2053_), .B(reset_n), .Y(_0word0_reg_31_0__15_));
AND2X2 AND2X2_739 ( .A(core_siphash_valid_reg), .B(core_siphash_word_16_), .Y(_abc_19873_new_n2055_));
AND2X2 AND2X2_74 ( .A(_abc_19873_new_n894_), .B(core_finalize), .Y(_abc_19873_new_n983_));
AND2X2 AND2X2_740 ( .A(_abc_19873_new_n1607_), .B(word0_reg_16_), .Y(_abc_19873_new_n2056_));
AND2X2 AND2X2_741 ( .A(_abc_19873_new_n2057_), .B(reset_n), .Y(_0word0_reg_31_0__16_));
AND2X2 AND2X2_742 ( .A(core_siphash_valid_reg), .B(core_siphash_word_17_), .Y(_abc_19873_new_n2059_));
AND2X2 AND2X2_743 ( .A(_abc_19873_new_n1607_), .B(word0_reg_17_), .Y(_abc_19873_new_n2060_));
AND2X2 AND2X2_744 ( .A(_abc_19873_new_n2061_), .B(reset_n), .Y(_0word0_reg_31_0__17_));
AND2X2 AND2X2_745 ( .A(core_siphash_valid_reg), .B(core_siphash_word_18_), .Y(_abc_19873_new_n2063_));
AND2X2 AND2X2_746 ( .A(_abc_19873_new_n1607_), .B(word0_reg_18_), .Y(_abc_19873_new_n2064_));
AND2X2 AND2X2_747 ( .A(_abc_19873_new_n2065_), .B(reset_n), .Y(_0word0_reg_31_0__18_));
AND2X2 AND2X2_748 ( .A(core_siphash_valid_reg), .B(core_siphash_word_19_), .Y(_abc_19873_new_n2067_));
AND2X2 AND2X2_749 ( .A(_abc_19873_new_n1607_), .B(word0_reg_19_), .Y(_abc_19873_new_n2068_));
AND2X2 AND2X2_75 ( .A(_abc_19873_new_n987_), .B(_abc_19873_new_n937_), .Y(\read_data[2] ));
AND2X2 AND2X2_750 ( .A(_abc_19873_new_n2069_), .B(reset_n), .Y(_0word0_reg_31_0__19_));
AND2X2 AND2X2_751 ( .A(core_siphash_valid_reg), .B(core_siphash_word_20_), .Y(_abc_19873_new_n2071_));
AND2X2 AND2X2_752 ( .A(_abc_19873_new_n1607_), .B(word0_reg_20_), .Y(_abc_19873_new_n2072_));
AND2X2 AND2X2_753 ( .A(_abc_19873_new_n2073_), .B(reset_n), .Y(_0word0_reg_31_0__20_));
AND2X2 AND2X2_754 ( .A(core_siphash_valid_reg), .B(core_siphash_word_21_), .Y(_abc_19873_new_n2075_));
AND2X2 AND2X2_755 ( .A(_abc_19873_new_n1607_), .B(word0_reg_21_), .Y(_abc_19873_new_n2076_));
AND2X2 AND2X2_756 ( .A(_abc_19873_new_n2077_), .B(reset_n), .Y(_0word0_reg_31_0__21_));
AND2X2 AND2X2_757 ( .A(core_siphash_valid_reg), .B(core_siphash_word_22_), .Y(_abc_19873_new_n2079_));
AND2X2 AND2X2_758 ( .A(_abc_19873_new_n1607_), .B(word0_reg_22_), .Y(_abc_19873_new_n2080_));
AND2X2 AND2X2_759 ( .A(_abc_19873_new_n2081_), .B(reset_n), .Y(_0word0_reg_31_0__22_));
AND2X2 AND2X2_76 ( .A(_abc_19873_new_n912_), .B(word3_reg_3_), .Y(_abc_19873_new_n989_));
AND2X2 AND2X2_760 ( .A(core_siphash_valid_reg), .B(core_siphash_word_23_), .Y(_abc_19873_new_n2083_));
AND2X2 AND2X2_761 ( .A(_abc_19873_new_n1607_), .B(word0_reg_23_), .Y(_abc_19873_new_n2084_));
AND2X2 AND2X2_762 ( .A(_abc_19873_new_n2085_), .B(reset_n), .Y(_0word0_reg_31_0__23_));
AND2X2 AND2X2_763 ( .A(core_siphash_valid_reg), .B(core_siphash_word_24_), .Y(_abc_19873_new_n2087_));
AND2X2 AND2X2_764 ( .A(_abc_19873_new_n1607_), .B(word0_reg_24_), .Y(_abc_19873_new_n2088_));
AND2X2 AND2X2_765 ( .A(_abc_19873_new_n2089_), .B(reset_n), .Y(_0word0_reg_31_0__24_));
AND2X2 AND2X2_766 ( .A(core_siphash_valid_reg), .B(core_siphash_word_25_), .Y(_abc_19873_new_n2091_));
AND2X2 AND2X2_767 ( .A(_abc_19873_new_n1607_), .B(word0_reg_25_), .Y(_abc_19873_new_n2092_));
AND2X2 AND2X2_768 ( .A(_abc_19873_new_n2093_), .B(reset_n), .Y(_0word0_reg_31_0__25_));
AND2X2 AND2X2_769 ( .A(core_siphash_valid_reg), .B(core_siphash_word_26_), .Y(_abc_19873_new_n2095_));
AND2X2 AND2X2_77 ( .A(_abc_19873_new_n888_), .B(core_mi_3_), .Y(_abc_19873_new_n990_));
AND2X2 AND2X2_770 ( .A(_abc_19873_new_n1607_), .B(word0_reg_26_), .Y(_abc_19873_new_n2096_));
AND2X2 AND2X2_771 ( .A(_abc_19873_new_n2097_), .B(reset_n), .Y(_0word0_reg_31_0__26_));
AND2X2 AND2X2_772 ( .A(core_siphash_valid_reg), .B(core_siphash_word_27_), .Y(_abc_19873_new_n2099_));
AND2X2 AND2X2_773 ( .A(_abc_19873_new_n1607_), .B(word0_reg_27_), .Y(_abc_19873_new_n2100_));
AND2X2 AND2X2_774 ( .A(_abc_19873_new_n2101_), .B(reset_n), .Y(_0word0_reg_31_0__27_));
AND2X2 AND2X2_775 ( .A(core_siphash_valid_reg), .B(core_siphash_word_28_), .Y(_abc_19873_new_n2103_));
AND2X2 AND2X2_776 ( .A(_abc_19873_new_n1607_), .B(word0_reg_28_), .Y(_abc_19873_new_n2104_));
AND2X2 AND2X2_777 ( .A(_abc_19873_new_n2105_), .B(reset_n), .Y(_0word0_reg_31_0__28_));
AND2X2 AND2X2_778 ( .A(core_siphash_valid_reg), .B(core_siphash_word_29_), .Y(_abc_19873_new_n2107_));
AND2X2 AND2X2_779 ( .A(_abc_19873_new_n1607_), .B(word0_reg_29_), .Y(_abc_19873_new_n2108_));
AND2X2 AND2X2_78 ( .A(_abc_19873_new_n919_), .B(core_mi_35_), .Y(_abc_19873_new_n991_));
AND2X2 AND2X2_780 ( .A(_abc_19873_new_n2109_), .B(reset_n), .Y(_0word0_reg_31_0__29_));
AND2X2 AND2X2_781 ( .A(core_siphash_valid_reg), .B(core_siphash_word_30_), .Y(_abc_19873_new_n2111_));
AND2X2 AND2X2_782 ( .A(_abc_19873_new_n1607_), .B(word0_reg_30_), .Y(_abc_19873_new_n2112_));
AND2X2 AND2X2_783 ( .A(_abc_19873_new_n2113_), .B(reset_n), .Y(_0word0_reg_31_0__30_));
AND2X2 AND2X2_784 ( .A(core_siphash_valid_reg), .B(core_siphash_word_31_), .Y(_abc_19873_new_n2115_));
AND2X2 AND2X2_785 ( .A(_abc_19873_new_n1607_), .B(word0_reg_31_), .Y(_abc_19873_new_n2116_));
AND2X2 AND2X2_786 ( .A(_abc_19873_new_n2117_), .B(reset_n), .Y(_0word0_reg_31_0__31_));
AND2X2 AND2X2_787 ( .A(we), .B(cs), .Y(_abc_19873_new_n2119_));
AND2X2 AND2X2_788 ( .A(_abc_19873_new_n919_), .B(_abc_19873_new_n2119_), .Y(_abc_19873_new_n2120_));
AND2X2 AND2X2_789 ( .A(_abc_19873_new_n2120_), .B(_abc_19873_new_n2122_), .Y(_abc_19873_new_n2123_));
AND2X2 AND2X2_79 ( .A(_abc_19873_new_n897_), .B(core_compression_rounds_3_), .Y(_abc_19873_new_n993_));
AND2X2 AND2X2_790 ( .A(_abc_19873_new_n2124_), .B(_abc_19873_new_n2121_), .Y(_abc_19873_new_n2125_));
AND2X2 AND2X2_791 ( .A(_abc_19873_new_n2125_), .B(reset_n), .Y(_0mi1_reg_31_0__0_));
AND2X2 AND2X2_792 ( .A(_abc_19873_new_n2120_), .B(_abc_19873_new_n2128_), .Y(_abc_19873_new_n2129_));
AND2X2 AND2X2_793 ( .A(_abc_19873_new_n2130_), .B(_abc_19873_new_n2127_), .Y(_abc_19873_new_n2131_));
AND2X2 AND2X2_794 ( .A(_abc_19873_new_n2131_), .B(reset_n), .Y(_0mi1_reg_31_0__1_));
AND2X2 AND2X2_795 ( .A(_abc_19873_new_n2120_), .B(_abc_19873_new_n2134_), .Y(_abc_19873_new_n2135_));
AND2X2 AND2X2_796 ( .A(_abc_19873_new_n2136_), .B(_abc_19873_new_n2133_), .Y(_abc_19873_new_n2137_));
AND2X2 AND2X2_797 ( .A(_abc_19873_new_n2137_), .B(reset_n), .Y(_0mi1_reg_31_0__2_));
AND2X2 AND2X2_798 ( .A(_abc_19873_new_n2120_), .B(_abc_19873_new_n2140_), .Y(_abc_19873_new_n2141_));
AND2X2 AND2X2_799 ( .A(_abc_19873_new_n2142_), .B(_abc_19873_new_n2139_), .Y(_abc_19873_new_n2143_));
AND2X2 AND2X2_8 ( .A(_abc_19873_new_n881_), .B(core_key_96_), .Y(_abc_19873_new_n882_));
AND2X2 AND2X2_80 ( .A(_abc_19873_new_n893_), .B(_abc_19873_new_n900_), .Y(_abc_19873_new_n994_));
AND2X2 AND2X2_800 ( .A(_abc_19873_new_n2143_), .B(reset_n), .Y(_0mi1_reg_31_0__3_));
AND2X2 AND2X2_801 ( .A(_abc_19873_new_n2120_), .B(_abc_19873_new_n2146_), .Y(_abc_19873_new_n2147_));
AND2X2 AND2X2_802 ( .A(_abc_19873_new_n2148_), .B(_abc_19873_new_n2145_), .Y(_abc_19873_new_n2149_));
AND2X2 AND2X2_803 ( .A(_abc_19873_new_n2149_), .B(reset_n), .Y(_0mi1_reg_31_0__4_));
AND2X2 AND2X2_804 ( .A(_abc_19873_new_n2120_), .B(_abc_19873_new_n2152_), .Y(_abc_19873_new_n2153_));
AND2X2 AND2X2_805 ( .A(_abc_19873_new_n2154_), .B(_abc_19873_new_n2151_), .Y(_abc_19873_new_n2155_));
AND2X2 AND2X2_806 ( .A(_abc_19873_new_n2155_), .B(reset_n), .Y(_0mi1_reg_31_0__5_));
AND2X2 AND2X2_807 ( .A(_abc_19873_new_n2120_), .B(_abc_19873_new_n2158_), .Y(_abc_19873_new_n2159_));
AND2X2 AND2X2_808 ( .A(_abc_19873_new_n2160_), .B(_abc_19873_new_n2157_), .Y(_abc_19873_new_n2161_));
AND2X2 AND2X2_809 ( .A(_abc_19873_new_n2161_), .B(reset_n), .Y(_0mi1_reg_31_0__6_));
AND2X2 AND2X2_81 ( .A(_abc_19873_new_n925_), .B(word2_reg_3_), .Y(_abc_19873_new_n998_));
AND2X2 AND2X2_810 ( .A(_abc_19873_new_n2120_), .B(_abc_19873_new_n2164_), .Y(_abc_19873_new_n2165_));
AND2X2 AND2X2_811 ( .A(_abc_19873_new_n2166_), .B(_abc_19873_new_n2163_), .Y(_abc_19873_new_n2167_));
AND2X2 AND2X2_812 ( .A(_abc_19873_new_n2167_), .B(reset_n), .Y(_0mi1_reg_31_0__7_));
AND2X2 AND2X2_813 ( .A(_abc_19873_new_n2120_), .B(_abc_19873_new_n2170_), .Y(_abc_19873_new_n2171_));
AND2X2 AND2X2_814 ( .A(_abc_19873_new_n2172_), .B(_abc_19873_new_n2169_), .Y(_abc_19873_new_n2173_));
AND2X2 AND2X2_815 ( .A(_abc_19873_new_n2173_), .B(reset_n), .Y(_0mi1_reg_31_0__8_));
AND2X2 AND2X2_816 ( .A(_abc_19873_new_n2120_), .B(_abc_19873_new_n2176_), .Y(_abc_19873_new_n2177_));
AND2X2 AND2X2_817 ( .A(_abc_19873_new_n2178_), .B(_abc_19873_new_n2175_), .Y(_abc_19873_new_n2179_));
AND2X2 AND2X2_818 ( .A(_abc_19873_new_n2179_), .B(reset_n), .Y(_0mi1_reg_31_0__9_));
AND2X2 AND2X2_819 ( .A(_abc_19873_new_n2120_), .B(_abc_19873_new_n2182_), .Y(_abc_19873_new_n2183_));
AND2X2 AND2X2_82 ( .A(_abc_19873_new_n930_), .B(word0_reg_3_), .Y(_abc_19873_new_n999_));
AND2X2 AND2X2_820 ( .A(_abc_19873_new_n2184_), .B(_abc_19873_new_n2181_), .Y(_abc_19873_new_n2185_));
AND2X2 AND2X2_821 ( .A(_abc_19873_new_n2185_), .B(reset_n), .Y(_0mi1_reg_31_0__10_));
AND2X2 AND2X2_822 ( .A(_abc_19873_new_n2120_), .B(_abc_19873_new_n2188_), .Y(_abc_19873_new_n2189_));
AND2X2 AND2X2_823 ( .A(_abc_19873_new_n2190_), .B(_abc_19873_new_n2187_), .Y(_abc_19873_new_n2191_));
AND2X2 AND2X2_824 ( .A(_abc_19873_new_n2191_), .B(reset_n), .Y(_0mi1_reg_31_0__11_));
AND2X2 AND2X2_825 ( .A(_abc_19873_new_n2120_), .B(_abc_19873_new_n2194_), .Y(_abc_19873_new_n2195_));
AND2X2 AND2X2_826 ( .A(_abc_19873_new_n2196_), .B(_abc_19873_new_n2193_), .Y(_abc_19873_new_n2197_));
AND2X2 AND2X2_827 ( .A(_abc_19873_new_n2197_), .B(reset_n), .Y(_0mi1_reg_31_0__12_));
AND2X2 AND2X2_828 ( .A(_abc_19873_new_n2120_), .B(_abc_19873_new_n2200_), .Y(_abc_19873_new_n2201_));
AND2X2 AND2X2_829 ( .A(_abc_19873_new_n2202_), .B(_abc_19873_new_n2199_), .Y(_abc_19873_new_n2203_));
AND2X2 AND2X2_83 ( .A(_abc_19873_new_n907_), .B(word1_reg_3_), .Y(_abc_19873_new_n1000_));
AND2X2 AND2X2_830 ( .A(_abc_19873_new_n2203_), .B(reset_n), .Y(_0mi1_reg_31_0__13_));
AND2X2 AND2X2_831 ( .A(_abc_19873_new_n2120_), .B(_abc_19873_new_n2206_), .Y(_abc_19873_new_n2207_));
AND2X2 AND2X2_832 ( .A(_abc_19873_new_n2208_), .B(_abc_19873_new_n2205_), .Y(_abc_19873_new_n2209_));
AND2X2 AND2X2_833 ( .A(_abc_19873_new_n2209_), .B(reset_n), .Y(_0mi1_reg_31_0__14_));
AND2X2 AND2X2_834 ( .A(_abc_19873_new_n2120_), .B(_abc_19873_new_n2212_), .Y(_abc_19873_new_n2213_));
AND2X2 AND2X2_835 ( .A(_abc_19873_new_n2214_), .B(_abc_19873_new_n2211_), .Y(_abc_19873_new_n2215_));
AND2X2 AND2X2_836 ( .A(_abc_19873_new_n2215_), .B(reset_n), .Y(_0mi1_reg_31_0__15_));
AND2X2 AND2X2_837 ( .A(_abc_19873_new_n2120_), .B(_abc_19873_new_n2218_), .Y(_abc_19873_new_n2219_));
AND2X2 AND2X2_838 ( .A(_abc_19873_new_n2220_), .B(_abc_19873_new_n2217_), .Y(_abc_19873_new_n2221_));
AND2X2 AND2X2_839 ( .A(_abc_19873_new_n2221_), .B(reset_n), .Y(_0mi1_reg_31_0__16_));
AND2X2 AND2X2_84 ( .A(_abc_19873_new_n928_), .B(core_key_35_), .Y(_abc_19873_new_n1003_));
AND2X2 AND2X2_840 ( .A(_abc_19873_new_n2120_), .B(_abc_19873_new_n2224_), .Y(_abc_19873_new_n2225_));
AND2X2 AND2X2_841 ( .A(_abc_19873_new_n2226_), .B(_abc_19873_new_n2223_), .Y(_abc_19873_new_n2227_));
AND2X2 AND2X2_842 ( .A(_abc_19873_new_n2227_), .B(reset_n), .Y(_0mi1_reg_31_0__17_));
AND2X2 AND2X2_843 ( .A(_abc_19873_new_n2120_), .B(_abc_19873_new_n2230_), .Y(_abc_19873_new_n2231_));
AND2X2 AND2X2_844 ( .A(_abc_19873_new_n2232_), .B(_abc_19873_new_n2229_), .Y(_abc_19873_new_n2233_));
AND2X2 AND2X2_845 ( .A(_abc_19873_new_n2233_), .B(reset_n), .Y(_0mi1_reg_31_0__18_));
AND2X2 AND2X2_846 ( .A(_abc_19873_new_n2120_), .B(_abc_19873_new_n2236_), .Y(_abc_19873_new_n2237_));
AND2X2 AND2X2_847 ( .A(_abc_19873_new_n2238_), .B(_abc_19873_new_n2235_), .Y(_abc_19873_new_n2239_));
AND2X2 AND2X2_848 ( .A(_abc_19873_new_n2239_), .B(reset_n), .Y(_0mi1_reg_31_0__19_));
AND2X2 AND2X2_849 ( .A(_abc_19873_new_n2120_), .B(_abc_19873_new_n2242_), .Y(_abc_19873_new_n2243_));
AND2X2 AND2X2_85 ( .A(_abc_19873_new_n901_), .B(core_key_3_), .Y(_abc_19873_new_n1004_));
AND2X2 AND2X2_850 ( .A(_abc_19873_new_n2244_), .B(_abc_19873_new_n2241_), .Y(_abc_19873_new_n2245_));
AND2X2 AND2X2_851 ( .A(_abc_19873_new_n2245_), .B(reset_n), .Y(_0mi1_reg_31_0__20_));
AND2X2 AND2X2_852 ( .A(_abc_19873_new_n2120_), .B(_abc_19873_new_n2248_), .Y(_abc_19873_new_n2249_));
AND2X2 AND2X2_853 ( .A(_abc_19873_new_n2250_), .B(_abc_19873_new_n2247_), .Y(_abc_19873_new_n2251_));
AND2X2 AND2X2_854 ( .A(_abc_19873_new_n2251_), .B(reset_n), .Y(_0mi1_reg_31_0__21_));
AND2X2 AND2X2_855 ( .A(_abc_19873_new_n2120_), .B(_abc_19873_new_n2254_), .Y(_abc_19873_new_n2255_));
AND2X2 AND2X2_856 ( .A(_abc_19873_new_n2256_), .B(_abc_19873_new_n2253_), .Y(_abc_19873_new_n2257_));
AND2X2 AND2X2_857 ( .A(_abc_19873_new_n2257_), .B(reset_n), .Y(_0mi1_reg_31_0__22_));
AND2X2 AND2X2_858 ( .A(_abc_19873_new_n2120_), .B(_abc_19873_new_n2260_), .Y(_abc_19873_new_n2261_));
AND2X2 AND2X2_859 ( .A(_abc_19873_new_n2262_), .B(_abc_19873_new_n2259_), .Y(_abc_19873_new_n2263_));
AND2X2 AND2X2_86 ( .A(_abc_19873_new_n881_), .B(core_key_99_), .Y(_abc_19873_new_n1006_));
AND2X2 AND2X2_860 ( .A(_abc_19873_new_n2263_), .B(reset_n), .Y(_0mi1_reg_31_0__23_));
AND2X2 AND2X2_861 ( .A(_abc_19873_new_n2120_), .B(_abc_19873_new_n2266_), .Y(_abc_19873_new_n2267_));
AND2X2 AND2X2_862 ( .A(_abc_19873_new_n2268_), .B(_abc_19873_new_n2265_), .Y(_abc_19873_new_n2269_));
AND2X2 AND2X2_863 ( .A(_abc_19873_new_n2269_), .B(reset_n), .Y(_0mi1_reg_31_0__24_));
AND2X2 AND2X2_864 ( .A(_abc_19873_new_n2120_), .B(_abc_19873_new_n2272_), .Y(_abc_19873_new_n2273_));
AND2X2 AND2X2_865 ( .A(_abc_19873_new_n2274_), .B(_abc_19873_new_n2271_), .Y(_abc_19873_new_n2275_));
AND2X2 AND2X2_866 ( .A(_abc_19873_new_n2275_), .B(reset_n), .Y(_0mi1_reg_31_0__25_));
AND2X2 AND2X2_867 ( .A(_abc_19873_new_n2120_), .B(_abc_19873_new_n2278_), .Y(_abc_19873_new_n2279_));
AND2X2 AND2X2_868 ( .A(_abc_19873_new_n2280_), .B(_abc_19873_new_n2277_), .Y(_abc_19873_new_n2281_));
AND2X2 AND2X2_869 ( .A(_abc_19873_new_n2281_), .B(reset_n), .Y(_0mi1_reg_31_0__26_));
AND2X2 AND2X2_87 ( .A(_abc_19873_new_n916_), .B(core_key_67_), .Y(_abc_19873_new_n1007_));
AND2X2 AND2X2_870 ( .A(_abc_19873_new_n2120_), .B(_abc_19873_new_n2284_), .Y(_abc_19873_new_n2285_));
AND2X2 AND2X2_871 ( .A(_abc_19873_new_n2286_), .B(_abc_19873_new_n2283_), .Y(_abc_19873_new_n2287_));
AND2X2 AND2X2_872 ( .A(_abc_19873_new_n2287_), .B(reset_n), .Y(_0mi1_reg_31_0__27_));
AND2X2 AND2X2_873 ( .A(_abc_19873_new_n2120_), .B(_abc_19873_new_n2290_), .Y(_abc_19873_new_n2291_));
AND2X2 AND2X2_874 ( .A(_abc_19873_new_n2292_), .B(_abc_19873_new_n2289_), .Y(_abc_19873_new_n2293_));
AND2X2 AND2X2_875 ( .A(_abc_19873_new_n2293_), .B(reset_n), .Y(_0mi1_reg_31_0__28_));
AND2X2 AND2X2_876 ( .A(_abc_19873_new_n2120_), .B(_abc_19873_new_n2296_), .Y(_abc_19873_new_n2297_));
AND2X2 AND2X2_877 ( .A(_abc_19873_new_n2298_), .B(_abc_19873_new_n2295_), .Y(_abc_19873_new_n2299_));
AND2X2 AND2X2_878 ( .A(_abc_19873_new_n2299_), .B(reset_n), .Y(_0mi1_reg_31_0__29_));
AND2X2 AND2X2_879 ( .A(_abc_19873_new_n2120_), .B(_abc_19873_new_n2302_), .Y(_abc_19873_new_n2303_));
AND2X2 AND2X2_88 ( .A(_abc_19873_new_n1011_), .B(_abc_19873_new_n937_), .Y(\read_data[3] ));
AND2X2 AND2X2_880 ( .A(_abc_19873_new_n2304_), .B(_abc_19873_new_n2301_), .Y(_abc_19873_new_n2305_));
AND2X2 AND2X2_881 ( .A(_abc_19873_new_n2305_), .B(reset_n), .Y(_0mi1_reg_31_0__30_));
AND2X2 AND2X2_882 ( .A(_abc_19873_new_n2120_), .B(_abc_19873_new_n2308_), .Y(_abc_19873_new_n2309_));
AND2X2 AND2X2_883 ( .A(_abc_19873_new_n2310_), .B(_abc_19873_new_n2307_), .Y(_abc_19873_new_n2311_));
AND2X2 AND2X2_884 ( .A(_abc_19873_new_n2311_), .B(reset_n), .Y(_0mi1_reg_31_0__31_));
AND2X2 AND2X2_885 ( .A(_abc_19873_new_n888_), .B(_abc_19873_new_n2119_), .Y(_abc_19873_new_n2313_));
AND2X2 AND2X2_886 ( .A(_abc_19873_new_n2313_), .B(_abc_19873_new_n2122_), .Y(_abc_19873_new_n2315_));
AND2X2 AND2X2_887 ( .A(_abc_19873_new_n2316_), .B(reset_n), .Y(_abc_19873_new_n2317_));
AND2X2 AND2X2_888 ( .A(_abc_19873_new_n2317_), .B(_abc_19873_new_n2314_), .Y(_0mi0_reg_31_0__0_));
AND2X2 AND2X2_889 ( .A(_abc_19873_new_n2313_), .B(_abc_19873_new_n2128_), .Y(_abc_19873_new_n2320_));
AND2X2 AND2X2_89 ( .A(_abc_19873_new_n912_), .B(word3_reg_4_), .Y(_abc_19873_new_n1013_));
AND2X2 AND2X2_890 ( .A(_abc_19873_new_n2321_), .B(reset_n), .Y(_abc_19873_new_n2322_));
AND2X2 AND2X2_891 ( .A(_abc_19873_new_n2322_), .B(_abc_19873_new_n2319_), .Y(_0mi0_reg_31_0__1_));
AND2X2 AND2X2_892 ( .A(_abc_19873_new_n2313_), .B(_abc_19873_new_n2134_), .Y(_abc_19873_new_n2325_));
AND2X2 AND2X2_893 ( .A(_abc_19873_new_n2326_), .B(reset_n), .Y(_abc_19873_new_n2327_));
AND2X2 AND2X2_894 ( .A(_abc_19873_new_n2327_), .B(_abc_19873_new_n2324_), .Y(_0mi0_reg_31_0__2_));
AND2X2 AND2X2_895 ( .A(_abc_19873_new_n2313_), .B(_abc_19873_new_n2140_), .Y(_abc_19873_new_n2330_));
AND2X2 AND2X2_896 ( .A(_abc_19873_new_n2331_), .B(reset_n), .Y(_abc_19873_new_n2332_));
AND2X2 AND2X2_897 ( .A(_abc_19873_new_n2332_), .B(_abc_19873_new_n2329_), .Y(_0mi0_reg_31_0__3_));
AND2X2 AND2X2_898 ( .A(_abc_19873_new_n2313_), .B(_abc_19873_new_n2146_), .Y(_abc_19873_new_n2335_));
AND2X2 AND2X2_899 ( .A(_abc_19873_new_n2336_), .B(reset_n), .Y(_abc_19873_new_n2337_));
AND2X2 AND2X2_9 ( .A(_abc_19873_new_n883_), .B(_abc_19873_new_n884_), .Y(_abc_19873_new_n885_));
AND2X2 AND2X2_90 ( .A(_abc_19873_new_n888_), .B(core_mi_4_), .Y(_abc_19873_new_n1014_));
AND2X2 AND2X2_900 ( .A(_abc_19873_new_n2337_), .B(_abc_19873_new_n2334_), .Y(_0mi0_reg_31_0__4_));
AND2X2 AND2X2_901 ( .A(_abc_19873_new_n2313_), .B(_abc_19873_new_n2152_), .Y(_abc_19873_new_n2340_));
AND2X2 AND2X2_902 ( .A(_abc_19873_new_n2341_), .B(reset_n), .Y(_abc_19873_new_n2342_));
AND2X2 AND2X2_903 ( .A(_abc_19873_new_n2342_), .B(_abc_19873_new_n2339_), .Y(_0mi0_reg_31_0__5_));
AND2X2 AND2X2_904 ( .A(_abc_19873_new_n2313_), .B(_abc_19873_new_n2158_), .Y(_abc_19873_new_n2345_));
AND2X2 AND2X2_905 ( .A(_abc_19873_new_n2346_), .B(reset_n), .Y(_abc_19873_new_n2347_));
AND2X2 AND2X2_906 ( .A(_abc_19873_new_n2347_), .B(_abc_19873_new_n2344_), .Y(_0mi0_reg_31_0__6_));
AND2X2 AND2X2_907 ( .A(_abc_19873_new_n2313_), .B(_abc_19873_new_n2164_), .Y(_abc_19873_new_n2350_));
AND2X2 AND2X2_908 ( .A(_abc_19873_new_n2351_), .B(reset_n), .Y(_abc_19873_new_n2352_));
AND2X2 AND2X2_909 ( .A(_abc_19873_new_n2352_), .B(_abc_19873_new_n2349_), .Y(_0mi0_reg_31_0__7_));
AND2X2 AND2X2_91 ( .A(_abc_19873_new_n919_), .B(core_mi_36_), .Y(_abc_19873_new_n1015_));
AND2X2 AND2X2_910 ( .A(_abc_19873_new_n2313_), .B(_abc_19873_new_n2170_), .Y(_abc_19873_new_n2355_));
AND2X2 AND2X2_911 ( .A(_abc_19873_new_n2356_), .B(reset_n), .Y(_abc_19873_new_n2357_));
AND2X2 AND2X2_912 ( .A(_abc_19873_new_n2357_), .B(_abc_19873_new_n2354_), .Y(_0mi0_reg_31_0__8_));
AND2X2 AND2X2_913 ( .A(_abc_19873_new_n2313_), .B(_abc_19873_new_n2176_), .Y(_abc_19873_new_n2360_));
AND2X2 AND2X2_914 ( .A(_abc_19873_new_n2361_), .B(reset_n), .Y(_abc_19873_new_n2362_));
AND2X2 AND2X2_915 ( .A(_abc_19873_new_n2362_), .B(_abc_19873_new_n2359_), .Y(_0mi0_reg_31_0__9_));
AND2X2 AND2X2_916 ( .A(_abc_19873_new_n2313_), .B(_abc_19873_new_n2182_), .Y(_abc_19873_new_n2365_));
AND2X2 AND2X2_917 ( .A(_abc_19873_new_n2366_), .B(reset_n), .Y(_abc_19873_new_n2367_));
AND2X2 AND2X2_918 ( .A(_abc_19873_new_n2367_), .B(_abc_19873_new_n2364_), .Y(_0mi0_reg_31_0__10_));
AND2X2 AND2X2_919 ( .A(_abc_19873_new_n2313_), .B(_abc_19873_new_n2188_), .Y(_abc_19873_new_n2370_));
AND2X2 AND2X2_92 ( .A(_abc_19873_new_n897_), .B(core_final_rounds_0_), .Y(_abc_19873_new_n1017_));
AND2X2 AND2X2_920 ( .A(_abc_19873_new_n2371_), .B(reset_n), .Y(_abc_19873_new_n2372_));
AND2X2 AND2X2_921 ( .A(_abc_19873_new_n2372_), .B(_abc_19873_new_n2369_), .Y(_0mi0_reg_31_0__11_));
AND2X2 AND2X2_922 ( .A(_abc_19873_new_n2313_), .B(_abc_19873_new_n2194_), .Y(_abc_19873_new_n2375_));
AND2X2 AND2X2_923 ( .A(_abc_19873_new_n2376_), .B(reset_n), .Y(_abc_19873_new_n2377_));
AND2X2 AND2X2_924 ( .A(_abc_19873_new_n2377_), .B(_abc_19873_new_n2374_), .Y(_0mi0_reg_31_0__12_));
AND2X2 AND2X2_925 ( .A(_abc_19873_new_n2313_), .B(_abc_19873_new_n2200_), .Y(_abc_19873_new_n2380_));
AND2X2 AND2X2_926 ( .A(_abc_19873_new_n2381_), .B(reset_n), .Y(_abc_19873_new_n2382_));
AND2X2 AND2X2_927 ( .A(_abc_19873_new_n2382_), .B(_abc_19873_new_n2379_), .Y(_0mi0_reg_31_0__13_));
AND2X2 AND2X2_928 ( .A(_abc_19873_new_n2313_), .B(_abc_19873_new_n2206_), .Y(_abc_19873_new_n2385_));
AND2X2 AND2X2_929 ( .A(_abc_19873_new_n2386_), .B(reset_n), .Y(_abc_19873_new_n2387_));
AND2X2 AND2X2_93 ( .A(_abc_19873_new_n893_), .B(_abc_19873_new_n915_), .Y(_abc_19873_new_n1018_));
AND2X2 AND2X2_930 ( .A(_abc_19873_new_n2387_), .B(_abc_19873_new_n2384_), .Y(_0mi0_reg_31_0__14_));
AND2X2 AND2X2_931 ( .A(_abc_19873_new_n2313_), .B(_abc_19873_new_n2212_), .Y(_abc_19873_new_n2390_));
AND2X2 AND2X2_932 ( .A(_abc_19873_new_n2391_), .B(reset_n), .Y(_abc_19873_new_n2392_));
AND2X2 AND2X2_933 ( .A(_abc_19873_new_n2392_), .B(_abc_19873_new_n2389_), .Y(_0mi0_reg_31_0__15_));
AND2X2 AND2X2_934 ( .A(_abc_19873_new_n2313_), .B(_abc_19873_new_n2218_), .Y(_abc_19873_new_n2395_));
AND2X2 AND2X2_935 ( .A(_abc_19873_new_n2396_), .B(reset_n), .Y(_abc_19873_new_n2397_));
AND2X2 AND2X2_936 ( .A(_abc_19873_new_n2397_), .B(_abc_19873_new_n2394_), .Y(_0mi0_reg_31_0__16_));
AND2X2 AND2X2_937 ( .A(_abc_19873_new_n2313_), .B(_abc_19873_new_n2224_), .Y(_abc_19873_new_n2400_));
AND2X2 AND2X2_938 ( .A(_abc_19873_new_n2401_), .B(reset_n), .Y(_abc_19873_new_n2402_));
AND2X2 AND2X2_939 ( .A(_abc_19873_new_n2402_), .B(_abc_19873_new_n2399_), .Y(_0mi0_reg_31_0__17_));
AND2X2 AND2X2_94 ( .A(_abc_19873_new_n925_), .B(word2_reg_4_), .Y(_abc_19873_new_n1022_));
AND2X2 AND2X2_940 ( .A(_abc_19873_new_n2313_), .B(_abc_19873_new_n2230_), .Y(_abc_19873_new_n2405_));
AND2X2 AND2X2_941 ( .A(_abc_19873_new_n2406_), .B(reset_n), .Y(_abc_19873_new_n2407_));
AND2X2 AND2X2_942 ( .A(_abc_19873_new_n2407_), .B(_abc_19873_new_n2404_), .Y(_0mi0_reg_31_0__18_));
AND2X2 AND2X2_943 ( .A(_abc_19873_new_n2313_), .B(_abc_19873_new_n2236_), .Y(_abc_19873_new_n2410_));
AND2X2 AND2X2_944 ( .A(_abc_19873_new_n2411_), .B(reset_n), .Y(_abc_19873_new_n2412_));
AND2X2 AND2X2_945 ( .A(_abc_19873_new_n2412_), .B(_abc_19873_new_n2409_), .Y(_0mi0_reg_31_0__19_));
AND2X2 AND2X2_946 ( .A(_abc_19873_new_n2313_), .B(_abc_19873_new_n2242_), .Y(_abc_19873_new_n2415_));
AND2X2 AND2X2_947 ( .A(_abc_19873_new_n2416_), .B(reset_n), .Y(_abc_19873_new_n2417_));
AND2X2 AND2X2_948 ( .A(_abc_19873_new_n2417_), .B(_abc_19873_new_n2414_), .Y(_0mi0_reg_31_0__20_));
AND2X2 AND2X2_949 ( .A(_abc_19873_new_n2313_), .B(_abc_19873_new_n2248_), .Y(_abc_19873_new_n2420_));
AND2X2 AND2X2_95 ( .A(_abc_19873_new_n930_), .B(word0_reg_4_), .Y(_abc_19873_new_n1023_));
AND2X2 AND2X2_950 ( .A(_abc_19873_new_n2421_), .B(reset_n), .Y(_abc_19873_new_n2422_));
AND2X2 AND2X2_951 ( .A(_abc_19873_new_n2422_), .B(_abc_19873_new_n2419_), .Y(_0mi0_reg_31_0__21_));
AND2X2 AND2X2_952 ( .A(_abc_19873_new_n2313_), .B(_abc_19873_new_n2254_), .Y(_abc_19873_new_n2425_));
AND2X2 AND2X2_953 ( .A(_abc_19873_new_n2426_), .B(reset_n), .Y(_abc_19873_new_n2427_));
AND2X2 AND2X2_954 ( .A(_abc_19873_new_n2427_), .B(_abc_19873_new_n2424_), .Y(_0mi0_reg_31_0__22_));
AND2X2 AND2X2_955 ( .A(_abc_19873_new_n2313_), .B(_abc_19873_new_n2260_), .Y(_abc_19873_new_n2430_));
AND2X2 AND2X2_956 ( .A(_abc_19873_new_n2431_), .B(reset_n), .Y(_abc_19873_new_n2432_));
AND2X2 AND2X2_957 ( .A(_abc_19873_new_n2432_), .B(_abc_19873_new_n2429_), .Y(_0mi0_reg_31_0__23_));
AND2X2 AND2X2_958 ( .A(_abc_19873_new_n2313_), .B(_abc_19873_new_n2266_), .Y(_abc_19873_new_n2435_));
AND2X2 AND2X2_959 ( .A(_abc_19873_new_n2436_), .B(reset_n), .Y(_abc_19873_new_n2437_));
AND2X2 AND2X2_96 ( .A(_abc_19873_new_n907_), .B(word1_reg_4_), .Y(_abc_19873_new_n1024_));
AND2X2 AND2X2_960 ( .A(_abc_19873_new_n2437_), .B(_abc_19873_new_n2434_), .Y(_0mi0_reg_31_0__24_));
AND2X2 AND2X2_961 ( .A(_abc_19873_new_n2313_), .B(_abc_19873_new_n2272_), .Y(_abc_19873_new_n2440_));
AND2X2 AND2X2_962 ( .A(_abc_19873_new_n2441_), .B(reset_n), .Y(_abc_19873_new_n2442_));
AND2X2 AND2X2_963 ( .A(_abc_19873_new_n2442_), .B(_abc_19873_new_n2439_), .Y(_0mi0_reg_31_0__25_));
AND2X2 AND2X2_964 ( .A(_abc_19873_new_n2313_), .B(_abc_19873_new_n2278_), .Y(_abc_19873_new_n2445_));
AND2X2 AND2X2_965 ( .A(_abc_19873_new_n2446_), .B(reset_n), .Y(_abc_19873_new_n2447_));
AND2X2 AND2X2_966 ( .A(_abc_19873_new_n2447_), .B(_abc_19873_new_n2444_), .Y(_0mi0_reg_31_0__26_));
AND2X2 AND2X2_967 ( .A(_abc_19873_new_n2313_), .B(_abc_19873_new_n2284_), .Y(_abc_19873_new_n2450_));
AND2X2 AND2X2_968 ( .A(_abc_19873_new_n2451_), .B(reset_n), .Y(_abc_19873_new_n2452_));
AND2X2 AND2X2_969 ( .A(_abc_19873_new_n2452_), .B(_abc_19873_new_n2449_), .Y(_0mi0_reg_31_0__27_));
AND2X2 AND2X2_97 ( .A(_abc_19873_new_n901_), .B(core_key_4_), .Y(_abc_19873_new_n1027_));
AND2X2 AND2X2_970 ( .A(_abc_19873_new_n2313_), .B(_abc_19873_new_n2290_), .Y(_abc_19873_new_n2455_));
AND2X2 AND2X2_971 ( .A(_abc_19873_new_n2456_), .B(reset_n), .Y(_abc_19873_new_n2457_));
AND2X2 AND2X2_972 ( .A(_abc_19873_new_n2457_), .B(_abc_19873_new_n2454_), .Y(_0mi0_reg_31_0__28_));
AND2X2 AND2X2_973 ( .A(_abc_19873_new_n2313_), .B(_abc_19873_new_n2296_), .Y(_abc_19873_new_n2460_));
AND2X2 AND2X2_974 ( .A(_abc_19873_new_n2461_), .B(reset_n), .Y(_abc_19873_new_n2462_));
AND2X2 AND2X2_975 ( .A(_abc_19873_new_n2462_), .B(_abc_19873_new_n2459_), .Y(_0mi0_reg_31_0__29_));
AND2X2 AND2X2_976 ( .A(_abc_19873_new_n2313_), .B(_abc_19873_new_n2302_), .Y(_abc_19873_new_n2465_));
AND2X2 AND2X2_977 ( .A(_abc_19873_new_n2466_), .B(reset_n), .Y(_abc_19873_new_n2467_));
AND2X2 AND2X2_978 ( .A(_abc_19873_new_n2467_), .B(_abc_19873_new_n2464_), .Y(_0mi0_reg_31_0__30_));
AND2X2 AND2X2_979 ( .A(_abc_19873_new_n2313_), .B(_abc_19873_new_n2308_), .Y(_abc_19873_new_n2470_));
AND2X2 AND2X2_98 ( .A(_abc_19873_new_n928_), .B(core_key_36_), .Y(_abc_19873_new_n1028_));
AND2X2 AND2X2_980 ( .A(_abc_19873_new_n2471_), .B(reset_n), .Y(_abc_19873_new_n2472_));
AND2X2 AND2X2_981 ( .A(_abc_19873_new_n2472_), .B(_abc_19873_new_n2469_), .Y(_0mi0_reg_31_0__31_));
AND2X2 AND2X2_982 ( .A(_abc_19873_new_n881_), .B(_abc_19873_new_n2119_), .Y(_abc_19873_new_n2474_));
AND2X2 AND2X2_983 ( .A(_abc_19873_new_n2474_), .B(_abc_19873_new_n2122_), .Y(_abc_19873_new_n2476_));
AND2X2 AND2X2_984 ( .A(_abc_19873_new_n2477_), .B(reset_n), .Y(_abc_19873_new_n2478_));
AND2X2 AND2X2_985 ( .A(_abc_19873_new_n2478_), .B(_abc_19873_new_n2475_), .Y(_0key3_reg_31_0__0_));
AND2X2 AND2X2_986 ( .A(_abc_19873_new_n2474_), .B(_abc_19873_new_n2128_), .Y(_abc_19873_new_n2481_));
AND2X2 AND2X2_987 ( .A(_abc_19873_new_n2482_), .B(reset_n), .Y(_abc_19873_new_n2483_));
AND2X2 AND2X2_988 ( .A(_abc_19873_new_n2483_), .B(_abc_19873_new_n2480_), .Y(_0key3_reg_31_0__1_));
AND2X2 AND2X2_989 ( .A(_abc_19873_new_n2474_), .B(_abc_19873_new_n2134_), .Y(_abc_19873_new_n2486_));
AND2X2 AND2X2_99 ( .A(_abc_19873_new_n881_), .B(core_key_100_), .Y(_abc_19873_new_n1030_));
AND2X2 AND2X2_990 ( .A(_abc_19873_new_n2487_), .B(reset_n), .Y(_abc_19873_new_n2488_));
AND2X2 AND2X2_991 ( .A(_abc_19873_new_n2488_), .B(_abc_19873_new_n2485_), .Y(_0key3_reg_31_0__2_));
AND2X2 AND2X2_992 ( .A(_abc_19873_new_n2474_), .B(_abc_19873_new_n2140_), .Y(_abc_19873_new_n2491_));
AND2X2 AND2X2_993 ( .A(_abc_19873_new_n2492_), .B(reset_n), .Y(_abc_19873_new_n2493_));
AND2X2 AND2X2_994 ( .A(_abc_19873_new_n2493_), .B(_abc_19873_new_n2490_), .Y(_0key3_reg_31_0__3_));
AND2X2 AND2X2_995 ( .A(_abc_19873_new_n2474_), .B(_abc_19873_new_n2146_), .Y(_abc_19873_new_n2496_));
AND2X2 AND2X2_996 ( .A(_abc_19873_new_n2497_), .B(reset_n), .Y(_abc_19873_new_n2498_));
AND2X2 AND2X2_997 ( .A(_abc_19873_new_n2498_), .B(_abc_19873_new_n2495_), .Y(_0key3_reg_31_0__4_));
AND2X2 AND2X2_998 ( .A(_abc_19873_new_n2474_), .B(_abc_19873_new_n2152_), .Y(_abc_19873_new_n2501_));
AND2X2 AND2X2_999 ( .A(_abc_19873_new_n2502_), .B(reset_n), .Y(_abc_19873_new_n2503_));
DFFPOSX1 DFFPOSX1_1 ( .CLK(clk), .D(_0ctrl_reg_2_0__0_), .Q(core_initalize));
DFFPOSX1 DFFPOSX1_10 ( .CLK(clk), .D(_0param_reg_7_0__5_), .Q(core_final_rounds_1_));
DFFPOSX1 DFFPOSX1_100 ( .CLK(clk), .D(_0key2_reg_31_0__23_), .Q(core_key_87_));
DFFPOSX1 DFFPOSX1_101 ( .CLK(clk), .D(_0key2_reg_31_0__24_), .Q(core_key_88_));
DFFPOSX1 DFFPOSX1_102 ( .CLK(clk), .D(_0key2_reg_31_0__25_), .Q(core_key_89_));
DFFPOSX1 DFFPOSX1_103 ( .CLK(clk), .D(_0key2_reg_31_0__26_), .Q(core_key_90_));
DFFPOSX1 DFFPOSX1_104 ( .CLK(clk), .D(_0key2_reg_31_0__27_), .Q(core_key_91_));
DFFPOSX1 DFFPOSX1_105 ( .CLK(clk), .D(_0key2_reg_31_0__28_), .Q(core_key_92_));
DFFPOSX1 DFFPOSX1_106 ( .CLK(clk), .D(_0key2_reg_31_0__29_), .Q(core_key_93_));
DFFPOSX1 DFFPOSX1_107 ( .CLK(clk), .D(_0key2_reg_31_0__30_), .Q(core_key_94_));
DFFPOSX1 DFFPOSX1_108 ( .CLK(clk), .D(_0key2_reg_31_0__31_), .Q(core_key_95_));
DFFPOSX1 DFFPOSX1_109 ( .CLK(clk), .D(_0key3_reg_31_0__0_), .Q(core_key_96_));
DFFPOSX1 DFFPOSX1_11 ( .CLK(clk), .D(_0param_reg_7_0__6_), .Q(core_final_rounds_2_));
DFFPOSX1 DFFPOSX1_110 ( .CLK(clk), .D(_0key3_reg_31_0__1_), .Q(core_key_97_));
DFFPOSX1 DFFPOSX1_111 ( .CLK(clk), .D(_0key3_reg_31_0__2_), .Q(core_key_98_));
DFFPOSX1 DFFPOSX1_112 ( .CLK(clk), .D(_0key3_reg_31_0__3_), .Q(core_key_99_));
DFFPOSX1 DFFPOSX1_113 ( .CLK(clk), .D(_0key3_reg_31_0__4_), .Q(core_key_100_));
DFFPOSX1 DFFPOSX1_114 ( .CLK(clk), .D(_0key3_reg_31_0__5_), .Q(core_key_101_));
DFFPOSX1 DFFPOSX1_115 ( .CLK(clk), .D(_0key3_reg_31_0__6_), .Q(core_key_102_));
DFFPOSX1 DFFPOSX1_116 ( .CLK(clk), .D(_0key3_reg_31_0__7_), .Q(core_key_103_));
DFFPOSX1 DFFPOSX1_117 ( .CLK(clk), .D(_0key3_reg_31_0__8_), .Q(core_key_104_));
DFFPOSX1 DFFPOSX1_118 ( .CLK(clk), .D(_0key3_reg_31_0__9_), .Q(core_key_105_));
DFFPOSX1 DFFPOSX1_119 ( .CLK(clk), .D(_0key3_reg_31_0__10_), .Q(core_key_106_));
DFFPOSX1 DFFPOSX1_12 ( .CLK(clk), .D(_0param_reg_7_0__7_), .Q(core_final_rounds_3_));
DFFPOSX1 DFFPOSX1_120 ( .CLK(clk), .D(_0key3_reg_31_0__11_), .Q(core_key_107_));
DFFPOSX1 DFFPOSX1_121 ( .CLK(clk), .D(_0key3_reg_31_0__12_), .Q(core_key_108_));
DFFPOSX1 DFFPOSX1_122 ( .CLK(clk), .D(_0key3_reg_31_0__13_), .Q(core_key_109_));
DFFPOSX1 DFFPOSX1_123 ( .CLK(clk), .D(_0key3_reg_31_0__14_), .Q(core_key_110_));
DFFPOSX1 DFFPOSX1_124 ( .CLK(clk), .D(_0key3_reg_31_0__15_), .Q(core_key_111_));
DFFPOSX1 DFFPOSX1_125 ( .CLK(clk), .D(_0key3_reg_31_0__16_), .Q(core_key_112_));
DFFPOSX1 DFFPOSX1_126 ( .CLK(clk), .D(_0key3_reg_31_0__17_), .Q(core_key_113_));
DFFPOSX1 DFFPOSX1_127 ( .CLK(clk), .D(_0key3_reg_31_0__18_), .Q(core_key_114_));
DFFPOSX1 DFFPOSX1_128 ( .CLK(clk), .D(_0key3_reg_31_0__19_), .Q(core_key_115_));
DFFPOSX1 DFFPOSX1_129 ( .CLK(clk), .D(_0key3_reg_31_0__20_), .Q(core_key_116_));
DFFPOSX1 DFFPOSX1_13 ( .CLK(clk), .D(_0key0_reg_31_0__0_), .Q(core_key_0_));
DFFPOSX1 DFFPOSX1_130 ( .CLK(clk), .D(_0key3_reg_31_0__21_), .Q(core_key_117_));
DFFPOSX1 DFFPOSX1_131 ( .CLK(clk), .D(_0key3_reg_31_0__22_), .Q(core_key_118_));
DFFPOSX1 DFFPOSX1_132 ( .CLK(clk), .D(_0key3_reg_31_0__23_), .Q(core_key_119_));
DFFPOSX1 DFFPOSX1_133 ( .CLK(clk), .D(_0key3_reg_31_0__24_), .Q(core_key_120_));
DFFPOSX1 DFFPOSX1_134 ( .CLK(clk), .D(_0key3_reg_31_0__25_), .Q(core_key_121_));
DFFPOSX1 DFFPOSX1_135 ( .CLK(clk), .D(_0key3_reg_31_0__26_), .Q(core_key_122_));
DFFPOSX1 DFFPOSX1_136 ( .CLK(clk), .D(_0key3_reg_31_0__27_), .Q(core_key_123_));
DFFPOSX1 DFFPOSX1_137 ( .CLK(clk), .D(_0key3_reg_31_0__28_), .Q(core_key_124_));
DFFPOSX1 DFFPOSX1_138 ( .CLK(clk), .D(_0key3_reg_31_0__29_), .Q(core_key_125_));
DFFPOSX1 DFFPOSX1_139 ( .CLK(clk), .D(_0key3_reg_31_0__30_), .Q(core_key_126_));
DFFPOSX1 DFFPOSX1_14 ( .CLK(clk), .D(_0key0_reg_31_0__1_), .Q(core_key_1_));
DFFPOSX1 DFFPOSX1_140 ( .CLK(clk), .D(_0key3_reg_31_0__31_), .Q(core_key_127_));
DFFPOSX1 DFFPOSX1_141 ( .CLK(clk), .D(_0mi0_reg_31_0__0_), .Q(core_mi_0_));
DFFPOSX1 DFFPOSX1_142 ( .CLK(clk), .D(_0mi0_reg_31_0__1_), .Q(core_mi_1_));
DFFPOSX1 DFFPOSX1_143 ( .CLK(clk), .D(_0mi0_reg_31_0__2_), .Q(core_mi_2_));
DFFPOSX1 DFFPOSX1_144 ( .CLK(clk), .D(_0mi0_reg_31_0__3_), .Q(core_mi_3_));
DFFPOSX1 DFFPOSX1_145 ( .CLK(clk), .D(_0mi0_reg_31_0__4_), .Q(core_mi_4_));
DFFPOSX1 DFFPOSX1_146 ( .CLK(clk), .D(_0mi0_reg_31_0__5_), .Q(core_mi_5_));
DFFPOSX1 DFFPOSX1_147 ( .CLK(clk), .D(_0mi0_reg_31_0__6_), .Q(core_mi_6_));
DFFPOSX1 DFFPOSX1_148 ( .CLK(clk), .D(_0mi0_reg_31_0__7_), .Q(core_mi_7_));
DFFPOSX1 DFFPOSX1_149 ( .CLK(clk), .D(_0mi0_reg_31_0__8_), .Q(core_mi_8_));
DFFPOSX1 DFFPOSX1_15 ( .CLK(clk), .D(_0key0_reg_31_0__2_), .Q(core_key_2_));
DFFPOSX1 DFFPOSX1_150 ( .CLK(clk), .D(_0mi0_reg_31_0__9_), .Q(core_mi_9_));
DFFPOSX1 DFFPOSX1_151 ( .CLK(clk), .D(_0mi0_reg_31_0__10_), .Q(core_mi_10_));
DFFPOSX1 DFFPOSX1_152 ( .CLK(clk), .D(_0mi0_reg_31_0__11_), .Q(core_mi_11_));
DFFPOSX1 DFFPOSX1_153 ( .CLK(clk), .D(_0mi0_reg_31_0__12_), .Q(core_mi_12_));
DFFPOSX1 DFFPOSX1_154 ( .CLK(clk), .D(_0mi0_reg_31_0__13_), .Q(core_mi_13_));
DFFPOSX1 DFFPOSX1_155 ( .CLK(clk), .D(_0mi0_reg_31_0__14_), .Q(core_mi_14_));
DFFPOSX1 DFFPOSX1_156 ( .CLK(clk), .D(_0mi0_reg_31_0__15_), .Q(core_mi_15_));
DFFPOSX1 DFFPOSX1_157 ( .CLK(clk), .D(_0mi0_reg_31_0__16_), .Q(core_mi_16_));
DFFPOSX1 DFFPOSX1_158 ( .CLK(clk), .D(_0mi0_reg_31_0__17_), .Q(core_mi_17_));
DFFPOSX1 DFFPOSX1_159 ( .CLK(clk), .D(_0mi0_reg_31_0__18_), .Q(core_mi_18_));
DFFPOSX1 DFFPOSX1_16 ( .CLK(clk), .D(_0key0_reg_31_0__3_), .Q(core_key_3_));
DFFPOSX1 DFFPOSX1_160 ( .CLK(clk), .D(_0mi0_reg_31_0__19_), .Q(core_mi_19_));
DFFPOSX1 DFFPOSX1_161 ( .CLK(clk), .D(_0mi0_reg_31_0__20_), .Q(core_mi_20_));
DFFPOSX1 DFFPOSX1_162 ( .CLK(clk), .D(_0mi0_reg_31_0__21_), .Q(core_mi_21_));
DFFPOSX1 DFFPOSX1_163 ( .CLK(clk), .D(_0mi0_reg_31_0__22_), .Q(core_mi_22_));
DFFPOSX1 DFFPOSX1_164 ( .CLK(clk), .D(_0mi0_reg_31_0__23_), .Q(core_mi_23_));
DFFPOSX1 DFFPOSX1_165 ( .CLK(clk), .D(_0mi0_reg_31_0__24_), .Q(core_mi_24_));
DFFPOSX1 DFFPOSX1_166 ( .CLK(clk), .D(_0mi0_reg_31_0__25_), .Q(core_mi_25_));
DFFPOSX1 DFFPOSX1_167 ( .CLK(clk), .D(_0mi0_reg_31_0__26_), .Q(core_mi_26_));
DFFPOSX1 DFFPOSX1_168 ( .CLK(clk), .D(_0mi0_reg_31_0__27_), .Q(core_mi_27_));
DFFPOSX1 DFFPOSX1_169 ( .CLK(clk), .D(_0mi0_reg_31_0__28_), .Q(core_mi_28_));
DFFPOSX1 DFFPOSX1_17 ( .CLK(clk), .D(_0key0_reg_31_0__4_), .Q(core_key_4_));
DFFPOSX1 DFFPOSX1_170 ( .CLK(clk), .D(_0mi0_reg_31_0__29_), .Q(core_mi_29_));
DFFPOSX1 DFFPOSX1_171 ( .CLK(clk), .D(_0mi0_reg_31_0__30_), .Q(core_mi_30_));
DFFPOSX1 DFFPOSX1_172 ( .CLK(clk), .D(_0mi0_reg_31_0__31_), .Q(core_mi_31_));
DFFPOSX1 DFFPOSX1_173 ( .CLK(clk), .D(_0mi1_reg_31_0__0_), .Q(core_mi_32_));
DFFPOSX1 DFFPOSX1_174 ( .CLK(clk), .D(_0mi1_reg_31_0__1_), .Q(core_mi_33_));
DFFPOSX1 DFFPOSX1_175 ( .CLK(clk), .D(_0mi1_reg_31_0__2_), .Q(core_mi_34_));
DFFPOSX1 DFFPOSX1_176 ( .CLK(clk), .D(_0mi1_reg_31_0__3_), .Q(core_mi_35_));
DFFPOSX1 DFFPOSX1_177 ( .CLK(clk), .D(_0mi1_reg_31_0__4_), .Q(core_mi_36_));
DFFPOSX1 DFFPOSX1_178 ( .CLK(clk), .D(_0mi1_reg_31_0__5_), .Q(core_mi_37_));
DFFPOSX1 DFFPOSX1_179 ( .CLK(clk), .D(_0mi1_reg_31_0__6_), .Q(core_mi_38_));
DFFPOSX1 DFFPOSX1_18 ( .CLK(clk), .D(_0key0_reg_31_0__5_), .Q(core_key_5_));
DFFPOSX1 DFFPOSX1_180 ( .CLK(clk), .D(_0mi1_reg_31_0__7_), .Q(core_mi_39_));
DFFPOSX1 DFFPOSX1_181 ( .CLK(clk), .D(_0mi1_reg_31_0__8_), .Q(core_mi_40_));
DFFPOSX1 DFFPOSX1_182 ( .CLK(clk), .D(_0mi1_reg_31_0__9_), .Q(core_mi_41_));
DFFPOSX1 DFFPOSX1_183 ( .CLK(clk), .D(_0mi1_reg_31_0__10_), .Q(core_mi_42_));
DFFPOSX1 DFFPOSX1_184 ( .CLK(clk), .D(_0mi1_reg_31_0__11_), .Q(core_mi_43_));
DFFPOSX1 DFFPOSX1_185 ( .CLK(clk), .D(_0mi1_reg_31_0__12_), .Q(core_mi_44_));
DFFPOSX1 DFFPOSX1_186 ( .CLK(clk), .D(_0mi1_reg_31_0__13_), .Q(core_mi_45_));
DFFPOSX1 DFFPOSX1_187 ( .CLK(clk), .D(_0mi1_reg_31_0__14_), .Q(core_mi_46_));
DFFPOSX1 DFFPOSX1_188 ( .CLK(clk), .D(_0mi1_reg_31_0__15_), .Q(core_mi_47_));
DFFPOSX1 DFFPOSX1_189 ( .CLK(clk), .D(_0mi1_reg_31_0__16_), .Q(core_mi_48_));
DFFPOSX1 DFFPOSX1_19 ( .CLK(clk), .D(_0key0_reg_31_0__6_), .Q(core_key_6_));
DFFPOSX1 DFFPOSX1_190 ( .CLK(clk), .D(_0mi1_reg_31_0__17_), .Q(core_mi_49_));
DFFPOSX1 DFFPOSX1_191 ( .CLK(clk), .D(_0mi1_reg_31_0__18_), .Q(core_mi_50_));
DFFPOSX1 DFFPOSX1_192 ( .CLK(clk), .D(_0mi1_reg_31_0__19_), .Q(core_mi_51_));
DFFPOSX1 DFFPOSX1_193 ( .CLK(clk), .D(_0mi1_reg_31_0__20_), .Q(core_mi_52_));
DFFPOSX1 DFFPOSX1_194 ( .CLK(clk), .D(_0mi1_reg_31_0__21_), .Q(core_mi_53_));
DFFPOSX1 DFFPOSX1_195 ( .CLK(clk), .D(_0mi1_reg_31_0__22_), .Q(core_mi_54_));
DFFPOSX1 DFFPOSX1_196 ( .CLK(clk), .D(_0mi1_reg_31_0__23_), .Q(core_mi_55_));
DFFPOSX1 DFFPOSX1_197 ( .CLK(clk), .D(_0mi1_reg_31_0__24_), .Q(core_mi_56_));
DFFPOSX1 DFFPOSX1_198 ( .CLK(clk), .D(_0mi1_reg_31_0__25_), .Q(core_mi_57_));
DFFPOSX1 DFFPOSX1_199 ( .CLK(clk), .D(_0mi1_reg_31_0__26_), .Q(core_mi_58_));
DFFPOSX1 DFFPOSX1_2 ( .CLK(clk), .D(_0ctrl_reg_2_0__1_), .Q(core_compress));
DFFPOSX1 DFFPOSX1_20 ( .CLK(clk), .D(_0key0_reg_31_0__7_), .Q(core_key_7_));
DFFPOSX1 DFFPOSX1_200 ( .CLK(clk), .D(_0mi1_reg_31_0__27_), .Q(core_mi_59_));
DFFPOSX1 DFFPOSX1_201 ( .CLK(clk), .D(_0mi1_reg_31_0__28_), .Q(core_mi_60_));
DFFPOSX1 DFFPOSX1_202 ( .CLK(clk), .D(_0mi1_reg_31_0__29_), .Q(core_mi_61_));
DFFPOSX1 DFFPOSX1_203 ( .CLK(clk), .D(_0mi1_reg_31_0__30_), .Q(core_mi_62_));
DFFPOSX1 DFFPOSX1_204 ( .CLK(clk), .D(_0mi1_reg_31_0__31_), .Q(core_mi_63_));
DFFPOSX1 DFFPOSX1_205 ( .CLK(clk), .D(_0word0_reg_31_0__0_), .Q(word0_reg_0_));
DFFPOSX1 DFFPOSX1_206 ( .CLK(clk), .D(_0word0_reg_31_0__1_), .Q(word0_reg_1_));
DFFPOSX1 DFFPOSX1_207 ( .CLK(clk), .D(_0word0_reg_31_0__2_), .Q(word0_reg_2_));
DFFPOSX1 DFFPOSX1_208 ( .CLK(clk), .D(_0word0_reg_31_0__3_), .Q(word0_reg_3_));
DFFPOSX1 DFFPOSX1_209 ( .CLK(clk), .D(_0word0_reg_31_0__4_), .Q(word0_reg_4_));
DFFPOSX1 DFFPOSX1_21 ( .CLK(clk), .D(_0key0_reg_31_0__8_), .Q(core_key_8_));
DFFPOSX1 DFFPOSX1_210 ( .CLK(clk), .D(_0word0_reg_31_0__5_), .Q(word0_reg_5_));
DFFPOSX1 DFFPOSX1_211 ( .CLK(clk), .D(_0word0_reg_31_0__6_), .Q(word0_reg_6_));
DFFPOSX1 DFFPOSX1_212 ( .CLK(clk), .D(_0word0_reg_31_0__7_), .Q(word0_reg_7_));
DFFPOSX1 DFFPOSX1_213 ( .CLK(clk), .D(_0word0_reg_31_0__8_), .Q(word0_reg_8_));
DFFPOSX1 DFFPOSX1_214 ( .CLK(clk), .D(_0word0_reg_31_0__9_), .Q(word0_reg_9_));
DFFPOSX1 DFFPOSX1_215 ( .CLK(clk), .D(_0word0_reg_31_0__10_), .Q(word0_reg_10_));
DFFPOSX1 DFFPOSX1_216 ( .CLK(clk), .D(_0word0_reg_31_0__11_), .Q(word0_reg_11_));
DFFPOSX1 DFFPOSX1_217 ( .CLK(clk), .D(_0word0_reg_31_0__12_), .Q(word0_reg_12_));
DFFPOSX1 DFFPOSX1_218 ( .CLK(clk), .D(_0word0_reg_31_0__13_), .Q(word0_reg_13_));
DFFPOSX1 DFFPOSX1_219 ( .CLK(clk), .D(_0word0_reg_31_0__14_), .Q(word0_reg_14_));
DFFPOSX1 DFFPOSX1_22 ( .CLK(clk), .D(_0key0_reg_31_0__9_), .Q(core_key_9_));
DFFPOSX1 DFFPOSX1_220 ( .CLK(clk), .D(_0word0_reg_31_0__15_), .Q(word0_reg_15_));
DFFPOSX1 DFFPOSX1_221 ( .CLK(clk), .D(_0word0_reg_31_0__16_), .Q(word0_reg_16_));
DFFPOSX1 DFFPOSX1_222 ( .CLK(clk), .D(_0word0_reg_31_0__17_), .Q(word0_reg_17_));
DFFPOSX1 DFFPOSX1_223 ( .CLK(clk), .D(_0word0_reg_31_0__18_), .Q(word0_reg_18_));
DFFPOSX1 DFFPOSX1_224 ( .CLK(clk), .D(_0word0_reg_31_0__19_), .Q(word0_reg_19_));
DFFPOSX1 DFFPOSX1_225 ( .CLK(clk), .D(_0word0_reg_31_0__20_), .Q(word0_reg_20_));
DFFPOSX1 DFFPOSX1_226 ( .CLK(clk), .D(_0word0_reg_31_0__21_), .Q(word0_reg_21_));
DFFPOSX1 DFFPOSX1_227 ( .CLK(clk), .D(_0word0_reg_31_0__22_), .Q(word0_reg_22_));
DFFPOSX1 DFFPOSX1_228 ( .CLK(clk), .D(_0word0_reg_31_0__23_), .Q(word0_reg_23_));
DFFPOSX1 DFFPOSX1_229 ( .CLK(clk), .D(_0word0_reg_31_0__24_), .Q(word0_reg_24_));
DFFPOSX1 DFFPOSX1_23 ( .CLK(clk), .D(_0key0_reg_31_0__10_), .Q(core_key_10_));
DFFPOSX1 DFFPOSX1_230 ( .CLK(clk), .D(_0word0_reg_31_0__25_), .Q(word0_reg_25_));
DFFPOSX1 DFFPOSX1_231 ( .CLK(clk), .D(_0word0_reg_31_0__26_), .Q(word0_reg_26_));
DFFPOSX1 DFFPOSX1_232 ( .CLK(clk), .D(_0word0_reg_31_0__27_), .Q(word0_reg_27_));
DFFPOSX1 DFFPOSX1_233 ( .CLK(clk), .D(_0word0_reg_31_0__28_), .Q(word0_reg_28_));
DFFPOSX1 DFFPOSX1_234 ( .CLK(clk), .D(_0word0_reg_31_0__29_), .Q(word0_reg_29_));
DFFPOSX1 DFFPOSX1_235 ( .CLK(clk), .D(_0word0_reg_31_0__30_), .Q(word0_reg_30_));
DFFPOSX1 DFFPOSX1_236 ( .CLK(clk), .D(_0word0_reg_31_0__31_), .Q(word0_reg_31_));
DFFPOSX1 DFFPOSX1_237 ( .CLK(clk), .D(_0word1_reg_31_0__0_), .Q(word1_reg_0_));
DFFPOSX1 DFFPOSX1_238 ( .CLK(clk), .D(_0word1_reg_31_0__1_), .Q(word1_reg_1_));
DFFPOSX1 DFFPOSX1_239 ( .CLK(clk), .D(_0word1_reg_31_0__2_), .Q(word1_reg_2_));
DFFPOSX1 DFFPOSX1_24 ( .CLK(clk), .D(_0key0_reg_31_0__11_), .Q(core_key_11_));
DFFPOSX1 DFFPOSX1_240 ( .CLK(clk), .D(_0word1_reg_31_0__3_), .Q(word1_reg_3_));
DFFPOSX1 DFFPOSX1_241 ( .CLK(clk), .D(_0word1_reg_31_0__4_), .Q(word1_reg_4_));
DFFPOSX1 DFFPOSX1_242 ( .CLK(clk), .D(_0word1_reg_31_0__5_), .Q(word1_reg_5_));
DFFPOSX1 DFFPOSX1_243 ( .CLK(clk), .D(_0word1_reg_31_0__6_), .Q(word1_reg_6_));
DFFPOSX1 DFFPOSX1_244 ( .CLK(clk), .D(_0word1_reg_31_0__7_), .Q(word1_reg_7_));
DFFPOSX1 DFFPOSX1_245 ( .CLK(clk), .D(_0word1_reg_31_0__8_), .Q(word1_reg_8_));
DFFPOSX1 DFFPOSX1_246 ( .CLK(clk), .D(_0word1_reg_31_0__9_), .Q(word1_reg_9_));
DFFPOSX1 DFFPOSX1_247 ( .CLK(clk), .D(_0word1_reg_31_0__10_), .Q(word1_reg_10_));
DFFPOSX1 DFFPOSX1_248 ( .CLK(clk), .D(_0word1_reg_31_0__11_), .Q(word1_reg_11_));
DFFPOSX1 DFFPOSX1_249 ( .CLK(clk), .D(_0word1_reg_31_0__12_), .Q(word1_reg_12_));
DFFPOSX1 DFFPOSX1_25 ( .CLK(clk), .D(_0key0_reg_31_0__12_), .Q(core_key_12_));
DFFPOSX1 DFFPOSX1_250 ( .CLK(clk), .D(_0word1_reg_31_0__13_), .Q(word1_reg_13_));
DFFPOSX1 DFFPOSX1_251 ( .CLK(clk), .D(_0word1_reg_31_0__14_), .Q(word1_reg_14_));
DFFPOSX1 DFFPOSX1_252 ( .CLK(clk), .D(_0word1_reg_31_0__15_), .Q(word1_reg_15_));
DFFPOSX1 DFFPOSX1_253 ( .CLK(clk), .D(_0word1_reg_31_0__16_), .Q(word1_reg_16_));
DFFPOSX1 DFFPOSX1_254 ( .CLK(clk), .D(_0word1_reg_31_0__17_), .Q(word1_reg_17_));
DFFPOSX1 DFFPOSX1_255 ( .CLK(clk), .D(_0word1_reg_31_0__18_), .Q(word1_reg_18_));
DFFPOSX1 DFFPOSX1_256 ( .CLK(clk), .D(_0word1_reg_31_0__19_), .Q(word1_reg_19_));
DFFPOSX1 DFFPOSX1_257 ( .CLK(clk), .D(_0word1_reg_31_0__20_), .Q(word1_reg_20_));
DFFPOSX1 DFFPOSX1_258 ( .CLK(clk), .D(_0word1_reg_31_0__21_), .Q(word1_reg_21_));
DFFPOSX1 DFFPOSX1_259 ( .CLK(clk), .D(_0word1_reg_31_0__22_), .Q(word1_reg_22_));
DFFPOSX1 DFFPOSX1_26 ( .CLK(clk), .D(_0key0_reg_31_0__13_), .Q(core_key_13_));
DFFPOSX1 DFFPOSX1_260 ( .CLK(clk), .D(_0word1_reg_31_0__23_), .Q(word1_reg_23_));
DFFPOSX1 DFFPOSX1_261 ( .CLK(clk), .D(_0word1_reg_31_0__24_), .Q(word1_reg_24_));
DFFPOSX1 DFFPOSX1_262 ( .CLK(clk), .D(_0word1_reg_31_0__25_), .Q(word1_reg_25_));
DFFPOSX1 DFFPOSX1_263 ( .CLK(clk), .D(_0word1_reg_31_0__26_), .Q(word1_reg_26_));
DFFPOSX1 DFFPOSX1_264 ( .CLK(clk), .D(_0word1_reg_31_0__27_), .Q(word1_reg_27_));
DFFPOSX1 DFFPOSX1_265 ( .CLK(clk), .D(_0word1_reg_31_0__28_), .Q(word1_reg_28_));
DFFPOSX1 DFFPOSX1_266 ( .CLK(clk), .D(_0word1_reg_31_0__29_), .Q(word1_reg_29_));
DFFPOSX1 DFFPOSX1_267 ( .CLK(clk), .D(_0word1_reg_31_0__30_), .Q(word1_reg_30_));
DFFPOSX1 DFFPOSX1_268 ( .CLK(clk), .D(_0word1_reg_31_0__31_), .Q(word1_reg_31_));
DFFPOSX1 DFFPOSX1_269 ( .CLK(clk), .D(_0word2_reg_31_0__0_), .Q(word2_reg_0_));
DFFPOSX1 DFFPOSX1_27 ( .CLK(clk), .D(_0key0_reg_31_0__14_), .Q(core_key_14_));
DFFPOSX1 DFFPOSX1_270 ( .CLK(clk), .D(_0word2_reg_31_0__1_), .Q(word2_reg_1_));
DFFPOSX1 DFFPOSX1_271 ( .CLK(clk), .D(_0word2_reg_31_0__2_), .Q(word2_reg_2_));
DFFPOSX1 DFFPOSX1_272 ( .CLK(clk), .D(_0word2_reg_31_0__3_), .Q(word2_reg_3_));
DFFPOSX1 DFFPOSX1_273 ( .CLK(clk), .D(_0word2_reg_31_0__4_), .Q(word2_reg_4_));
DFFPOSX1 DFFPOSX1_274 ( .CLK(clk), .D(_0word2_reg_31_0__5_), .Q(word2_reg_5_));
DFFPOSX1 DFFPOSX1_275 ( .CLK(clk), .D(_0word2_reg_31_0__6_), .Q(word2_reg_6_));
DFFPOSX1 DFFPOSX1_276 ( .CLK(clk), .D(_0word2_reg_31_0__7_), .Q(word2_reg_7_));
DFFPOSX1 DFFPOSX1_277 ( .CLK(clk), .D(_0word2_reg_31_0__8_), .Q(word2_reg_8_));
DFFPOSX1 DFFPOSX1_278 ( .CLK(clk), .D(_0word2_reg_31_0__9_), .Q(word2_reg_9_));
DFFPOSX1 DFFPOSX1_279 ( .CLK(clk), .D(_0word2_reg_31_0__10_), .Q(word2_reg_10_));
DFFPOSX1 DFFPOSX1_28 ( .CLK(clk), .D(_0key0_reg_31_0__15_), .Q(core_key_15_));
DFFPOSX1 DFFPOSX1_280 ( .CLK(clk), .D(_0word2_reg_31_0__11_), .Q(word2_reg_11_));
DFFPOSX1 DFFPOSX1_281 ( .CLK(clk), .D(_0word2_reg_31_0__12_), .Q(word2_reg_12_));
DFFPOSX1 DFFPOSX1_282 ( .CLK(clk), .D(_0word2_reg_31_0__13_), .Q(word2_reg_13_));
DFFPOSX1 DFFPOSX1_283 ( .CLK(clk), .D(_0word2_reg_31_0__14_), .Q(word2_reg_14_));
DFFPOSX1 DFFPOSX1_284 ( .CLK(clk), .D(_0word2_reg_31_0__15_), .Q(word2_reg_15_));
DFFPOSX1 DFFPOSX1_285 ( .CLK(clk), .D(_0word2_reg_31_0__16_), .Q(word2_reg_16_));
DFFPOSX1 DFFPOSX1_286 ( .CLK(clk), .D(_0word2_reg_31_0__17_), .Q(word2_reg_17_));
DFFPOSX1 DFFPOSX1_287 ( .CLK(clk), .D(_0word2_reg_31_0__18_), .Q(word2_reg_18_));
DFFPOSX1 DFFPOSX1_288 ( .CLK(clk), .D(_0word2_reg_31_0__19_), .Q(word2_reg_19_));
DFFPOSX1 DFFPOSX1_289 ( .CLK(clk), .D(_0word2_reg_31_0__20_), .Q(word2_reg_20_));
DFFPOSX1 DFFPOSX1_29 ( .CLK(clk), .D(_0key0_reg_31_0__16_), .Q(core_key_16_));
DFFPOSX1 DFFPOSX1_290 ( .CLK(clk), .D(_0word2_reg_31_0__21_), .Q(word2_reg_21_));
DFFPOSX1 DFFPOSX1_291 ( .CLK(clk), .D(_0word2_reg_31_0__22_), .Q(word2_reg_22_));
DFFPOSX1 DFFPOSX1_292 ( .CLK(clk), .D(_0word2_reg_31_0__23_), .Q(word2_reg_23_));
DFFPOSX1 DFFPOSX1_293 ( .CLK(clk), .D(_0word2_reg_31_0__24_), .Q(word2_reg_24_));
DFFPOSX1 DFFPOSX1_294 ( .CLK(clk), .D(_0word2_reg_31_0__25_), .Q(word2_reg_25_));
DFFPOSX1 DFFPOSX1_295 ( .CLK(clk), .D(_0word2_reg_31_0__26_), .Q(word2_reg_26_));
DFFPOSX1 DFFPOSX1_296 ( .CLK(clk), .D(_0word2_reg_31_0__27_), .Q(word2_reg_27_));
DFFPOSX1 DFFPOSX1_297 ( .CLK(clk), .D(_0word2_reg_31_0__28_), .Q(word2_reg_28_));
DFFPOSX1 DFFPOSX1_298 ( .CLK(clk), .D(_0word2_reg_31_0__29_), .Q(word2_reg_29_));
DFFPOSX1 DFFPOSX1_299 ( .CLK(clk), .D(_0word2_reg_31_0__30_), .Q(word2_reg_30_));
DFFPOSX1 DFFPOSX1_3 ( .CLK(clk), .D(_0ctrl_reg_2_0__2_), .Q(core_finalize));
DFFPOSX1 DFFPOSX1_30 ( .CLK(clk), .D(_0key0_reg_31_0__17_), .Q(core_key_17_));
DFFPOSX1 DFFPOSX1_300 ( .CLK(clk), .D(_0word2_reg_31_0__31_), .Q(word2_reg_31_));
DFFPOSX1 DFFPOSX1_301 ( .CLK(clk), .D(_0word3_reg_31_0__0_), .Q(word3_reg_0_));
DFFPOSX1 DFFPOSX1_302 ( .CLK(clk), .D(_0word3_reg_31_0__1_), .Q(word3_reg_1_));
DFFPOSX1 DFFPOSX1_303 ( .CLK(clk), .D(_0word3_reg_31_0__2_), .Q(word3_reg_2_));
DFFPOSX1 DFFPOSX1_304 ( .CLK(clk), .D(_0word3_reg_31_0__3_), .Q(word3_reg_3_));
DFFPOSX1 DFFPOSX1_305 ( .CLK(clk), .D(_0word3_reg_31_0__4_), .Q(word3_reg_4_));
DFFPOSX1 DFFPOSX1_306 ( .CLK(clk), .D(_0word3_reg_31_0__5_), .Q(word3_reg_5_));
DFFPOSX1 DFFPOSX1_307 ( .CLK(clk), .D(_0word3_reg_31_0__6_), .Q(word3_reg_6_));
DFFPOSX1 DFFPOSX1_308 ( .CLK(clk), .D(_0word3_reg_31_0__7_), .Q(word3_reg_7_));
DFFPOSX1 DFFPOSX1_309 ( .CLK(clk), .D(_0word3_reg_31_0__8_), .Q(word3_reg_8_));
DFFPOSX1 DFFPOSX1_31 ( .CLK(clk), .D(_0key0_reg_31_0__18_), .Q(core_key_18_));
DFFPOSX1 DFFPOSX1_310 ( .CLK(clk), .D(_0word3_reg_31_0__9_), .Q(word3_reg_9_));
DFFPOSX1 DFFPOSX1_311 ( .CLK(clk), .D(_0word3_reg_31_0__10_), .Q(word3_reg_10_));
DFFPOSX1 DFFPOSX1_312 ( .CLK(clk), .D(_0word3_reg_31_0__11_), .Q(word3_reg_11_));
DFFPOSX1 DFFPOSX1_313 ( .CLK(clk), .D(_0word3_reg_31_0__12_), .Q(word3_reg_12_));
DFFPOSX1 DFFPOSX1_314 ( .CLK(clk), .D(_0word3_reg_31_0__13_), .Q(word3_reg_13_));
DFFPOSX1 DFFPOSX1_315 ( .CLK(clk), .D(_0word3_reg_31_0__14_), .Q(word3_reg_14_));
DFFPOSX1 DFFPOSX1_316 ( .CLK(clk), .D(_0word3_reg_31_0__15_), .Q(word3_reg_15_));
DFFPOSX1 DFFPOSX1_317 ( .CLK(clk), .D(_0word3_reg_31_0__16_), .Q(word3_reg_16_));
DFFPOSX1 DFFPOSX1_318 ( .CLK(clk), .D(_0word3_reg_31_0__17_), .Q(word3_reg_17_));
DFFPOSX1 DFFPOSX1_319 ( .CLK(clk), .D(_0word3_reg_31_0__18_), .Q(word3_reg_18_));
DFFPOSX1 DFFPOSX1_32 ( .CLK(clk), .D(_0key0_reg_31_0__19_), .Q(core_key_19_));
DFFPOSX1 DFFPOSX1_320 ( .CLK(clk), .D(_0word3_reg_31_0__19_), .Q(word3_reg_19_));
DFFPOSX1 DFFPOSX1_321 ( .CLK(clk), .D(_0word3_reg_31_0__20_), .Q(word3_reg_20_));
DFFPOSX1 DFFPOSX1_322 ( .CLK(clk), .D(_0word3_reg_31_0__21_), .Q(word3_reg_21_));
DFFPOSX1 DFFPOSX1_323 ( .CLK(clk), .D(_0word3_reg_31_0__22_), .Q(word3_reg_22_));
DFFPOSX1 DFFPOSX1_324 ( .CLK(clk), .D(_0word3_reg_31_0__23_), .Q(word3_reg_23_));
DFFPOSX1 DFFPOSX1_325 ( .CLK(clk), .D(_0word3_reg_31_0__24_), .Q(word3_reg_24_));
DFFPOSX1 DFFPOSX1_326 ( .CLK(clk), .D(_0word3_reg_31_0__25_), .Q(word3_reg_25_));
DFFPOSX1 DFFPOSX1_327 ( .CLK(clk), .D(_0word3_reg_31_0__26_), .Q(word3_reg_26_));
DFFPOSX1 DFFPOSX1_328 ( .CLK(clk), .D(_0word3_reg_31_0__27_), .Q(word3_reg_27_));
DFFPOSX1 DFFPOSX1_329 ( .CLK(clk), .D(_0word3_reg_31_0__28_), .Q(word3_reg_28_));
DFFPOSX1 DFFPOSX1_33 ( .CLK(clk), .D(_0key0_reg_31_0__20_), .Q(core_key_20_));
DFFPOSX1 DFFPOSX1_330 ( .CLK(clk), .D(_0word3_reg_31_0__29_), .Q(word3_reg_29_));
DFFPOSX1 DFFPOSX1_331 ( .CLK(clk), .D(_0word3_reg_31_0__30_), .Q(word3_reg_30_));
DFFPOSX1 DFFPOSX1_332 ( .CLK(clk), .D(_0word3_reg_31_0__31_), .Q(word3_reg_31_));
DFFPOSX1 DFFPOSX1_333 ( .CLK(clk), .D(core__abc_15204_auto_fsm_map_cc_170_map_fsm_1439_0_), .Q(core_siphash_ctrl_reg_0_));
DFFPOSX1 DFFPOSX1_334 ( .CLK(clk), .D(core__abc_15204_auto_fsm_map_cc_118_implement_pattern_cache_1470), .Q(core_siphash_ctrl_reg_1_));
DFFPOSX1 DFFPOSX1_335 ( .CLK(clk), .D(core__abc_15204_auto_fsm_map_cc_118_implement_pattern_cache_1474), .Q(core_siphash_ctrl_reg_2_));
DFFPOSX1 DFFPOSX1_336 ( .CLK(clk), .D(core__abc_15204_auto_fsm_map_cc_170_map_fsm_1439_3_), .Q(core_siphash_ctrl_reg_3_));
DFFPOSX1 DFFPOSX1_337 ( .CLK(clk), .D(core__abc_15204_auto_fsm_map_cc_170_map_fsm_1439_4_), .Q(core_siphash_ctrl_reg_4_));
DFFPOSX1 DFFPOSX1_338 ( .CLK(clk), .D(core__abc_15204_auto_fsm_map_cc_118_implement_pattern_cache_1496), .Q(core_siphash_ctrl_reg_5_));
DFFPOSX1 DFFPOSX1_339 ( .CLK(clk), .D(core__abc_15204_auto_fsm_map_cc_170_map_fsm_1439_6_), .Q(core_siphash_ctrl_reg_6_));
DFFPOSX1 DFFPOSX1_34 ( .CLK(clk), .D(_0key0_reg_31_0__21_), .Q(core_key_21_));
DFFPOSX1 DFFPOSX1_340 ( .CLK(clk), .D(core__abc_15204_auto_fsm_map_cc_118_implement_pattern_cache_1509), .Q(core_siphash_word1_we));
DFFPOSX1 DFFPOSX1_341 ( .CLK(clk), .D(core__0v0_reg_63_0__0_), .Q(core_v0_reg_0_));
DFFPOSX1 DFFPOSX1_342 ( .CLK(clk), .D(core__0v0_reg_63_0__1_), .Q(core_v0_reg_1_));
DFFPOSX1 DFFPOSX1_343 ( .CLK(clk), .D(core__0v0_reg_63_0__2_), .Q(core_v0_reg_2_));
DFFPOSX1 DFFPOSX1_344 ( .CLK(clk), .D(core__0v0_reg_63_0__3_), .Q(core_v0_reg_3_));
DFFPOSX1 DFFPOSX1_345 ( .CLK(clk), .D(core__0v0_reg_63_0__4_), .Q(core_v0_reg_4_));
DFFPOSX1 DFFPOSX1_346 ( .CLK(clk), .D(core__0v0_reg_63_0__5_), .Q(core_v0_reg_5_));
DFFPOSX1 DFFPOSX1_347 ( .CLK(clk), .D(core__0v0_reg_63_0__6_), .Q(core_v0_reg_6_));
DFFPOSX1 DFFPOSX1_348 ( .CLK(clk), .D(core__0v0_reg_63_0__7_), .Q(core_v0_reg_7_));
DFFPOSX1 DFFPOSX1_349 ( .CLK(clk), .D(core__0v0_reg_63_0__8_), .Q(core_v0_reg_8_));
DFFPOSX1 DFFPOSX1_35 ( .CLK(clk), .D(_0key0_reg_31_0__22_), .Q(core_key_22_));
DFFPOSX1 DFFPOSX1_350 ( .CLK(clk), .D(core__0v0_reg_63_0__9_), .Q(core_v0_reg_9_));
DFFPOSX1 DFFPOSX1_351 ( .CLK(clk), .D(core__0v0_reg_63_0__10_), .Q(core_v0_reg_10_));
DFFPOSX1 DFFPOSX1_352 ( .CLK(clk), .D(core__0v0_reg_63_0__11_), .Q(core_v0_reg_11_));
DFFPOSX1 DFFPOSX1_353 ( .CLK(clk), .D(core__0v0_reg_63_0__12_), .Q(core_v0_reg_12_));
DFFPOSX1 DFFPOSX1_354 ( .CLK(clk), .D(core__0v0_reg_63_0__13_), .Q(core_v0_reg_13_));
DFFPOSX1 DFFPOSX1_355 ( .CLK(clk), .D(core__0v0_reg_63_0__14_), .Q(core_v0_reg_14_));
DFFPOSX1 DFFPOSX1_356 ( .CLK(clk), .D(core__0v0_reg_63_0__15_), .Q(core_v0_reg_15_));
DFFPOSX1 DFFPOSX1_357 ( .CLK(clk), .D(core__0v0_reg_63_0__16_), .Q(core_v0_reg_16_));
DFFPOSX1 DFFPOSX1_358 ( .CLK(clk), .D(core__0v0_reg_63_0__17_), .Q(core_v0_reg_17_));
DFFPOSX1 DFFPOSX1_359 ( .CLK(clk), .D(core__0v0_reg_63_0__18_), .Q(core_v0_reg_18_));
DFFPOSX1 DFFPOSX1_36 ( .CLK(clk), .D(_0key0_reg_31_0__23_), .Q(core_key_23_));
DFFPOSX1 DFFPOSX1_360 ( .CLK(clk), .D(core__0v0_reg_63_0__19_), .Q(core_v0_reg_19_));
DFFPOSX1 DFFPOSX1_361 ( .CLK(clk), .D(core__0v0_reg_63_0__20_), .Q(core_v0_reg_20_));
DFFPOSX1 DFFPOSX1_362 ( .CLK(clk), .D(core__0v0_reg_63_0__21_), .Q(core_v0_reg_21_));
DFFPOSX1 DFFPOSX1_363 ( .CLK(clk), .D(core__0v0_reg_63_0__22_), .Q(core_v0_reg_22_));
DFFPOSX1 DFFPOSX1_364 ( .CLK(clk), .D(core__0v0_reg_63_0__23_), .Q(core_v0_reg_23_));
DFFPOSX1 DFFPOSX1_365 ( .CLK(clk), .D(core__0v0_reg_63_0__24_), .Q(core_v0_reg_24_));
DFFPOSX1 DFFPOSX1_366 ( .CLK(clk), .D(core__0v0_reg_63_0__25_), .Q(core_v0_reg_25_));
DFFPOSX1 DFFPOSX1_367 ( .CLK(clk), .D(core__0v0_reg_63_0__26_), .Q(core_v0_reg_26_));
DFFPOSX1 DFFPOSX1_368 ( .CLK(clk), .D(core__0v0_reg_63_0__27_), .Q(core_v0_reg_27_));
DFFPOSX1 DFFPOSX1_369 ( .CLK(clk), .D(core__0v0_reg_63_0__28_), .Q(core_v0_reg_28_));
DFFPOSX1 DFFPOSX1_37 ( .CLK(clk), .D(_0key0_reg_31_0__24_), .Q(core_key_24_));
DFFPOSX1 DFFPOSX1_370 ( .CLK(clk), .D(core__0v0_reg_63_0__29_), .Q(core_v0_reg_29_));
DFFPOSX1 DFFPOSX1_371 ( .CLK(clk), .D(core__0v0_reg_63_0__30_), .Q(core_v0_reg_30_));
DFFPOSX1 DFFPOSX1_372 ( .CLK(clk), .D(core__0v0_reg_63_0__31_), .Q(core_v0_reg_31_));
DFFPOSX1 DFFPOSX1_373 ( .CLK(clk), .D(core__0v0_reg_63_0__32_), .Q(core_v0_reg_32_));
DFFPOSX1 DFFPOSX1_374 ( .CLK(clk), .D(core__0v0_reg_63_0__33_), .Q(core_v0_reg_33_));
DFFPOSX1 DFFPOSX1_375 ( .CLK(clk), .D(core__0v0_reg_63_0__34_), .Q(core_v0_reg_34_));
DFFPOSX1 DFFPOSX1_376 ( .CLK(clk), .D(core__0v0_reg_63_0__35_), .Q(core_v0_reg_35_));
DFFPOSX1 DFFPOSX1_377 ( .CLK(clk), .D(core__0v0_reg_63_0__36_), .Q(core_v0_reg_36_));
DFFPOSX1 DFFPOSX1_378 ( .CLK(clk), .D(core__0v0_reg_63_0__37_), .Q(core_v0_reg_37_));
DFFPOSX1 DFFPOSX1_379 ( .CLK(clk), .D(core__0v0_reg_63_0__38_), .Q(core_v0_reg_38_));
DFFPOSX1 DFFPOSX1_38 ( .CLK(clk), .D(_0key0_reg_31_0__25_), .Q(core_key_25_));
DFFPOSX1 DFFPOSX1_380 ( .CLK(clk), .D(core__0v0_reg_63_0__39_), .Q(core_v0_reg_39_));
DFFPOSX1 DFFPOSX1_381 ( .CLK(clk), .D(core__0v0_reg_63_0__40_), .Q(core_v0_reg_40_));
DFFPOSX1 DFFPOSX1_382 ( .CLK(clk), .D(core__0v0_reg_63_0__41_), .Q(core_v0_reg_41_));
DFFPOSX1 DFFPOSX1_383 ( .CLK(clk), .D(core__0v0_reg_63_0__42_), .Q(core_v0_reg_42_));
DFFPOSX1 DFFPOSX1_384 ( .CLK(clk), .D(core__0v0_reg_63_0__43_), .Q(core_v0_reg_43_));
DFFPOSX1 DFFPOSX1_385 ( .CLK(clk), .D(core__0v0_reg_63_0__44_), .Q(core_v0_reg_44_));
DFFPOSX1 DFFPOSX1_386 ( .CLK(clk), .D(core__0v0_reg_63_0__45_), .Q(core_v0_reg_45_));
DFFPOSX1 DFFPOSX1_387 ( .CLK(clk), .D(core__0v0_reg_63_0__46_), .Q(core_v0_reg_46_));
DFFPOSX1 DFFPOSX1_388 ( .CLK(clk), .D(core__0v0_reg_63_0__47_), .Q(core_v0_reg_47_));
DFFPOSX1 DFFPOSX1_389 ( .CLK(clk), .D(core__0v0_reg_63_0__48_), .Q(core_v0_reg_48_));
DFFPOSX1 DFFPOSX1_39 ( .CLK(clk), .D(_0key0_reg_31_0__26_), .Q(core_key_26_));
DFFPOSX1 DFFPOSX1_390 ( .CLK(clk), .D(core__0v0_reg_63_0__49_), .Q(core_v0_reg_49_));
DFFPOSX1 DFFPOSX1_391 ( .CLK(clk), .D(core__0v0_reg_63_0__50_), .Q(core_v0_reg_50_));
DFFPOSX1 DFFPOSX1_392 ( .CLK(clk), .D(core__0v0_reg_63_0__51_), .Q(core_v0_reg_51_));
DFFPOSX1 DFFPOSX1_393 ( .CLK(clk), .D(core__0v0_reg_63_0__52_), .Q(core_v0_reg_52_));
DFFPOSX1 DFFPOSX1_394 ( .CLK(clk), .D(core__0v0_reg_63_0__53_), .Q(core_v0_reg_53_));
DFFPOSX1 DFFPOSX1_395 ( .CLK(clk), .D(core__0v0_reg_63_0__54_), .Q(core_v0_reg_54_));
DFFPOSX1 DFFPOSX1_396 ( .CLK(clk), .D(core__0v0_reg_63_0__55_), .Q(core_v0_reg_55_));
DFFPOSX1 DFFPOSX1_397 ( .CLK(clk), .D(core__0v0_reg_63_0__56_), .Q(core_v0_reg_56_));
DFFPOSX1 DFFPOSX1_398 ( .CLK(clk), .D(core__0v0_reg_63_0__57_), .Q(core_v0_reg_57_));
DFFPOSX1 DFFPOSX1_399 ( .CLK(clk), .D(core__0v0_reg_63_0__58_), .Q(core_v0_reg_58_));
DFFPOSX1 DFFPOSX1_4 ( .CLK(clk), .D(_0long_reg_0_0_), .Q(core_long));
DFFPOSX1 DFFPOSX1_40 ( .CLK(clk), .D(_0key0_reg_31_0__27_), .Q(core_key_27_));
DFFPOSX1 DFFPOSX1_400 ( .CLK(clk), .D(core__0v0_reg_63_0__59_), .Q(core_v0_reg_59_));
DFFPOSX1 DFFPOSX1_401 ( .CLK(clk), .D(core__0v0_reg_63_0__60_), .Q(core_v0_reg_60_));
DFFPOSX1 DFFPOSX1_402 ( .CLK(clk), .D(core__0v0_reg_63_0__61_), .Q(core_v0_reg_61_));
DFFPOSX1 DFFPOSX1_403 ( .CLK(clk), .D(core__0v0_reg_63_0__62_), .Q(core_v0_reg_62_));
DFFPOSX1 DFFPOSX1_404 ( .CLK(clk), .D(core__0v0_reg_63_0__63_), .Q(core_v0_reg_63_));
DFFPOSX1 DFFPOSX1_405 ( .CLK(clk), .D(core__0v1_reg_63_0__0_), .Q(core_v1_reg_0_));
DFFPOSX1 DFFPOSX1_406 ( .CLK(clk), .D(core__0v1_reg_63_0__1_), .Q(core_v1_reg_1_));
DFFPOSX1 DFFPOSX1_407 ( .CLK(clk), .D(core__0v1_reg_63_0__2_), .Q(core_v1_reg_2_));
DFFPOSX1 DFFPOSX1_408 ( .CLK(clk), .D(core__0v1_reg_63_0__3_), .Q(core_v1_reg_3_));
DFFPOSX1 DFFPOSX1_409 ( .CLK(clk), .D(core__0v1_reg_63_0__4_), .Q(core_v1_reg_4_));
DFFPOSX1 DFFPOSX1_41 ( .CLK(clk), .D(_0key0_reg_31_0__28_), .Q(core_key_28_));
DFFPOSX1 DFFPOSX1_410 ( .CLK(clk), .D(core__0v1_reg_63_0__5_), .Q(core_v1_reg_5_));
DFFPOSX1 DFFPOSX1_411 ( .CLK(clk), .D(core__0v1_reg_63_0__6_), .Q(core_v1_reg_6_));
DFFPOSX1 DFFPOSX1_412 ( .CLK(clk), .D(core__0v1_reg_63_0__7_), .Q(core_v1_reg_7_));
DFFPOSX1 DFFPOSX1_413 ( .CLK(clk), .D(core__0v1_reg_63_0__8_), .Q(core_v1_reg_8_));
DFFPOSX1 DFFPOSX1_414 ( .CLK(clk), .D(core__0v1_reg_63_0__9_), .Q(core_v1_reg_9_));
DFFPOSX1 DFFPOSX1_415 ( .CLK(clk), .D(core__0v1_reg_63_0__10_), .Q(core_v1_reg_10_));
DFFPOSX1 DFFPOSX1_416 ( .CLK(clk), .D(core__0v1_reg_63_0__11_), .Q(core_v1_reg_11_));
DFFPOSX1 DFFPOSX1_417 ( .CLK(clk), .D(core__0v1_reg_63_0__12_), .Q(core_v1_reg_12_));
DFFPOSX1 DFFPOSX1_418 ( .CLK(clk), .D(core__0v1_reg_63_0__13_), .Q(core_v1_reg_13_));
DFFPOSX1 DFFPOSX1_419 ( .CLK(clk), .D(core__0v1_reg_63_0__14_), .Q(core_v1_reg_14_));
DFFPOSX1 DFFPOSX1_42 ( .CLK(clk), .D(_0key0_reg_31_0__29_), .Q(core_key_29_));
DFFPOSX1 DFFPOSX1_420 ( .CLK(clk), .D(core__0v1_reg_63_0__15_), .Q(core_v1_reg_15_));
DFFPOSX1 DFFPOSX1_421 ( .CLK(clk), .D(core__0v1_reg_63_0__16_), .Q(core_v1_reg_16_));
DFFPOSX1 DFFPOSX1_422 ( .CLK(clk), .D(core__0v1_reg_63_0__17_), .Q(core_v1_reg_17_));
DFFPOSX1 DFFPOSX1_423 ( .CLK(clk), .D(core__0v1_reg_63_0__18_), .Q(core_v1_reg_18_));
DFFPOSX1 DFFPOSX1_424 ( .CLK(clk), .D(core__0v1_reg_63_0__19_), .Q(core_v1_reg_19_));
DFFPOSX1 DFFPOSX1_425 ( .CLK(clk), .D(core__0v1_reg_63_0__20_), .Q(core_v1_reg_20_));
DFFPOSX1 DFFPOSX1_426 ( .CLK(clk), .D(core__0v1_reg_63_0__21_), .Q(core_v1_reg_21_));
DFFPOSX1 DFFPOSX1_427 ( .CLK(clk), .D(core__0v1_reg_63_0__22_), .Q(core_v1_reg_22_));
DFFPOSX1 DFFPOSX1_428 ( .CLK(clk), .D(core__0v1_reg_63_0__23_), .Q(core_v1_reg_23_));
DFFPOSX1 DFFPOSX1_429 ( .CLK(clk), .D(core__0v1_reg_63_0__24_), .Q(core_v1_reg_24_));
DFFPOSX1 DFFPOSX1_43 ( .CLK(clk), .D(_0key0_reg_31_0__30_), .Q(core_key_30_));
DFFPOSX1 DFFPOSX1_430 ( .CLK(clk), .D(core__0v1_reg_63_0__25_), .Q(core_v1_reg_25_));
DFFPOSX1 DFFPOSX1_431 ( .CLK(clk), .D(core__0v1_reg_63_0__26_), .Q(core_v1_reg_26_));
DFFPOSX1 DFFPOSX1_432 ( .CLK(clk), .D(core__0v1_reg_63_0__27_), .Q(core_v1_reg_27_));
DFFPOSX1 DFFPOSX1_433 ( .CLK(clk), .D(core__0v1_reg_63_0__28_), .Q(core_v1_reg_28_));
DFFPOSX1 DFFPOSX1_434 ( .CLK(clk), .D(core__0v1_reg_63_0__29_), .Q(core_v1_reg_29_));
DFFPOSX1 DFFPOSX1_435 ( .CLK(clk), .D(core__0v1_reg_63_0__30_), .Q(core_v1_reg_30_));
DFFPOSX1 DFFPOSX1_436 ( .CLK(clk), .D(core__0v1_reg_63_0__31_), .Q(core_v1_reg_31_));
DFFPOSX1 DFFPOSX1_437 ( .CLK(clk), .D(core__0v1_reg_63_0__32_), .Q(core_v1_reg_32_));
DFFPOSX1 DFFPOSX1_438 ( .CLK(clk), .D(core__0v1_reg_63_0__33_), .Q(core_v1_reg_33_));
DFFPOSX1 DFFPOSX1_439 ( .CLK(clk), .D(core__0v1_reg_63_0__34_), .Q(core_v1_reg_34_));
DFFPOSX1 DFFPOSX1_44 ( .CLK(clk), .D(_0key0_reg_31_0__31_), .Q(core_key_31_));
DFFPOSX1 DFFPOSX1_440 ( .CLK(clk), .D(core__0v1_reg_63_0__35_), .Q(core_v1_reg_35_));
DFFPOSX1 DFFPOSX1_441 ( .CLK(clk), .D(core__0v1_reg_63_0__36_), .Q(core_v1_reg_36_));
DFFPOSX1 DFFPOSX1_442 ( .CLK(clk), .D(core__0v1_reg_63_0__37_), .Q(core_v1_reg_37_));
DFFPOSX1 DFFPOSX1_443 ( .CLK(clk), .D(core__0v1_reg_63_0__38_), .Q(core_v1_reg_38_));
DFFPOSX1 DFFPOSX1_444 ( .CLK(clk), .D(core__0v1_reg_63_0__39_), .Q(core_v1_reg_39_));
DFFPOSX1 DFFPOSX1_445 ( .CLK(clk), .D(core__0v1_reg_63_0__40_), .Q(core_v1_reg_40_));
DFFPOSX1 DFFPOSX1_446 ( .CLK(clk), .D(core__0v1_reg_63_0__41_), .Q(core_v1_reg_41_));
DFFPOSX1 DFFPOSX1_447 ( .CLK(clk), .D(core__0v1_reg_63_0__42_), .Q(core_v1_reg_42_));
DFFPOSX1 DFFPOSX1_448 ( .CLK(clk), .D(core__0v1_reg_63_0__43_), .Q(core_v1_reg_43_));
DFFPOSX1 DFFPOSX1_449 ( .CLK(clk), .D(core__0v1_reg_63_0__44_), .Q(core_v1_reg_44_));
DFFPOSX1 DFFPOSX1_45 ( .CLK(clk), .D(_0key1_reg_31_0__0_), .Q(core_key_32_));
DFFPOSX1 DFFPOSX1_450 ( .CLK(clk), .D(core__0v1_reg_63_0__45_), .Q(core_v1_reg_45_));
DFFPOSX1 DFFPOSX1_451 ( .CLK(clk), .D(core__0v1_reg_63_0__46_), .Q(core_v1_reg_46_));
DFFPOSX1 DFFPOSX1_452 ( .CLK(clk), .D(core__0v1_reg_63_0__47_), .Q(core_v1_reg_47_));
DFFPOSX1 DFFPOSX1_453 ( .CLK(clk), .D(core__0v1_reg_63_0__48_), .Q(core_v1_reg_48_));
DFFPOSX1 DFFPOSX1_454 ( .CLK(clk), .D(core__0v1_reg_63_0__49_), .Q(core_v1_reg_49_));
DFFPOSX1 DFFPOSX1_455 ( .CLK(clk), .D(core__0v1_reg_63_0__50_), .Q(core_v1_reg_50_));
DFFPOSX1 DFFPOSX1_456 ( .CLK(clk), .D(core__0v1_reg_63_0__51_), .Q(core_v1_reg_51_));
DFFPOSX1 DFFPOSX1_457 ( .CLK(clk), .D(core__0v1_reg_63_0__52_), .Q(core_v1_reg_52_));
DFFPOSX1 DFFPOSX1_458 ( .CLK(clk), .D(core__0v1_reg_63_0__53_), .Q(core_v1_reg_53_));
DFFPOSX1 DFFPOSX1_459 ( .CLK(clk), .D(core__0v1_reg_63_0__54_), .Q(core_v1_reg_54_));
DFFPOSX1 DFFPOSX1_46 ( .CLK(clk), .D(_0key1_reg_31_0__1_), .Q(core_key_33_));
DFFPOSX1 DFFPOSX1_460 ( .CLK(clk), .D(core__0v1_reg_63_0__55_), .Q(core_v1_reg_55_));
DFFPOSX1 DFFPOSX1_461 ( .CLK(clk), .D(core__0v1_reg_63_0__56_), .Q(core_v1_reg_56_));
DFFPOSX1 DFFPOSX1_462 ( .CLK(clk), .D(core__0v1_reg_63_0__57_), .Q(core_v1_reg_57_));
DFFPOSX1 DFFPOSX1_463 ( .CLK(clk), .D(core__0v1_reg_63_0__58_), .Q(core_v1_reg_58_));
DFFPOSX1 DFFPOSX1_464 ( .CLK(clk), .D(core__0v1_reg_63_0__59_), .Q(core_v1_reg_59_));
DFFPOSX1 DFFPOSX1_465 ( .CLK(clk), .D(core__0v1_reg_63_0__60_), .Q(core_v1_reg_60_));
DFFPOSX1 DFFPOSX1_466 ( .CLK(clk), .D(core__0v1_reg_63_0__61_), .Q(core_v1_reg_61_));
DFFPOSX1 DFFPOSX1_467 ( .CLK(clk), .D(core__0v1_reg_63_0__62_), .Q(core_v1_reg_62_));
DFFPOSX1 DFFPOSX1_468 ( .CLK(clk), .D(core__0v1_reg_63_0__63_), .Q(core_v1_reg_63_));
DFFPOSX1 DFFPOSX1_469 ( .CLK(clk), .D(core__0v2_reg_63_0__0_), .Q(core_v2_reg_0_));
DFFPOSX1 DFFPOSX1_47 ( .CLK(clk), .D(_0key1_reg_31_0__2_), .Q(core_key_34_));
DFFPOSX1 DFFPOSX1_470 ( .CLK(clk), .D(core__0v2_reg_63_0__1_), .Q(core_v2_reg_1_));
DFFPOSX1 DFFPOSX1_471 ( .CLK(clk), .D(core__0v2_reg_63_0__2_), .Q(core_v2_reg_2_));
DFFPOSX1 DFFPOSX1_472 ( .CLK(clk), .D(core__0v2_reg_63_0__3_), .Q(core_v2_reg_3_));
DFFPOSX1 DFFPOSX1_473 ( .CLK(clk), .D(core__0v2_reg_63_0__4_), .Q(core_v2_reg_4_));
DFFPOSX1 DFFPOSX1_474 ( .CLK(clk), .D(core__0v2_reg_63_0__5_), .Q(core_v2_reg_5_));
DFFPOSX1 DFFPOSX1_475 ( .CLK(clk), .D(core__0v2_reg_63_0__6_), .Q(core_v2_reg_6_));
DFFPOSX1 DFFPOSX1_476 ( .CLK(clk), .D(core__0v2_reg_63_0__7_), .Q(core_v2_reg_7_));
DFFPOSX1 DFFPOSX1_477 ( .CLK(clk), .D(core__0v2_reg_63_0__8_), .Q(core_v2_reg_8_));
DFFPOSX1 DFFPOSX1_478 ( .CLK(clk), .D(core__0v2_reg_63_0__9_), .Q(core_v2_reg_9_));
DFFPOSX1 DFFPOSX1_479 ( .CLK(clk), .D(core__0v2_reg_63_0__10_), .Q(core_v2_reg_10_));
DFFPOSX1 DFFPOSX1_48 ( .CLK(clk), .D(_0key1_reg_31_0__3_), .Q(core_key_35_));
DFFPOSX1 DFFPOSX1_480 ( .CLK(clk), .D(core__0v2_reg_63_0__11_), .Q(core_v2_reg_11_));
DFFPOSX1 DFFPOSX1_481 ( .CLK(clk), .D(core__0v2_reg_63_0__12_), .Q(core_v2_reg_12_));
DFFPOSX1 DFFPOSX1_482 ( .CLK(clk), .D(core__0v2_reg_63_0__13_), .Q(core_v2_reg_13_));
DFFPOSX1 DFFPOSX1_483 ( .CLK(clk), .D(core__0v2_reg_63_0__14_), .Q(core_v2_reg_14_));
DFFPOSX1 DFFPOSX1_484 ( .CLK(clk), .D(core__0v2_reg_63_0__15_), .Q(core_v2_reg_15_));
DFFPOSX1 DFFPOSX1_485 ( .CLK(clk), .D(core__0v2_reg_63_0__16_), .Q(core_v2_reg_16_));
DFFPOSX1 DFFPOSX1_486 ( .CLK(clk), .D(core__0v2_reg_63_0__17_), .Q(core_v2_reg_17_));
DFFPOSX1 DFFPOSX1_487 ( .CLK(clk), .D(core__0v2_reg_63_0__18_), .Q(core_v2_reg_18_));
DFFPOSX1 DFFPOSX1_488 ( .CLK(clk), .D(core__0v2_reg_63_0__19_), .Q(core_v2_reg_19_));
DFFPOSX1 DFFPOSX1_489 ( .CLK(clk), .D(core__0v2_reg_63_0__20_), .Q(core_v2_reg_20_));
DFFPOSX1 DFFPOSX1_49 ( .CLK(clk), .D(_0key1_reg_31_0__4_), .Q(core_key_36_));
DFFPOSX1 DFFPOSX1_490 ( .CLK(clk), .D(core__0v2_reg_63_0__21_), .Q(core_v2_reg_21_));
DFFPOSX1 DFFPOSX1_491 ( .CLK(clk), .D(core__0v2_reg_63_0__22_), .Q(core_v2_reg_22_));
DFFPOSX1 DFFPOSX1_492 ( .CLK(clk), .D(core__0v2_reg_63_0__23_), .Q(core_v2_reg_23_));
DFFPOSX1 DFFPOSX1_493 ( .CLK(clk), .D(core__0v2_reg_63_0__24_), .Q(core_v2_reg_24_));
DFFPOSX1 DFFPOSX1_494 ( .CLK(clk), .D(core__0v2_reg_63_0__25_), .Q(core_v2_reg_25_));
DFFPOSX1 DFFPOSX1_495 ( .CLK(clk), .D(core__0v2_reg_63_0__26_), .Q(core_v2_reg_26_));
DFFPOSX1 DFFPOSX1_496 ( .CLK(clk), .D(core__0v2_reg_63_0__27_), .Q(core_v2_reg_27_));
DFFPOSX1 DFFPOSX1_497 ( .CLK(clk), .D(core__0v2_reg_63_0__28_), .Q(core_v2_reg_28_));
DFFPOSX1 DFFPOSX1_498 ( .CLK(clk), .D(core__0v2_reg_63_0__29_), .Q(core_v2_reg_29_));
DFFPOSX1 DFFPOSX1_499 ( .CLK(clk), .D(core__0v2_reg_63_0__30_), .Q(core_v2_reg_30_));
DFFPOSX1 DFFPOSX1_5 ( .CLK(clk), .D(_0param_reg_7_0__0_), .Q(core_compression_rounds_0_));
DFFPOSX1 DFFPOSX1_50 ( .CLK(clk), .D(_0key1_reg_31_0__5_), .Q(core_key_37_));
DFFPOSX1 DFFPOSX1_500 ( .CLK(clk), .D(core__0v2_reg_63_0__31_), .Q(core_v2_reg_31_));
DFFPOSX1 DFFPOSX1_501 ( .CLK(clk), .D(core__0v2_reg_63_0__32_), .Q(core_v2_reg_32_));
DFFPOSX1 DFFPOSX1_502 ( .CLK(clk), .D(core__0v2_reg_63_0__33_), .Q(core_v2_reg_33_));
DFFPOSX1 DFFPOSX1_503 ( .CLK(clk), .D(core__0v2_reg_63_0__34_), .Q(core_v2_reg_34_));
DFFPOSX1 DFFPOSX1_504 ( .CLK(clk), .D(core__0v2_reg_63_0__35_), .Q(core_v2_reg_35_));
DFFPOSX1 DFFPOSX1_505 ( .CLK(clk), .D(core__0v2_reg_63_0__36_), .Q(core_v2_reg_36_));
DFFPOSX1 DFFPOSX1_506 ( .CLK(clk), .D(core__0v2_reg_63_0__37_), .Q(core_v2_reg_37_));
DFFPOSX1 DFFPOSX1_507 ( .CLK(clk), .D(core__0v2_reg_63_0__38_), .Q(core_v2_reg_38_));
DFFPOSX1 DFFPOSX1_508 ( .CLK(clk), .D(core__0v2_reg_63_0__39_), .Q(core_v2_reg_39_));
DFFPOSX1 DFFPOSX1_509 ( .CLK(clk), .D(core__0v2_reg_63_0__40_), .Q(core_v2_reg_40_));
DFFPOSX1 DFFPOSX1_51 ( .CLK(clk), .D(_0key1_reg_31_0__6_), .Q(core_key_38_));
DFFPOSX1 DFFPOSX1_510 ( .CLK(clk), .D(core__0v2_reg_63_0__41_), .Q(core_v2_reg_41_));
DFFPOSX1 DFFPOSX1_511 ( .CLK(clk), .D(core__0v2_reg_63_0__42_), .Q(core_v2_reg_42_));
DFFPOSX1 DFFPOSX1_512 ( .CLK(clk), .D(core__0v2_reg_63_0__43_), .Q(core_v2_reg_43_));
DFFPOSX1 DFFPOSX1_513 ( .CLK(clk), .D(core__0v2_reg_63_0__44_), .Q(core_v2_reg_44_));
DFFPOSX1 DFFPOSX1_514 ( .CLK(clk), .D(core__0v2_reg_63_0__45_), .Q(core_v2_reg_45_));
DFFPOSX1 DFFPOSX1_515 ( .CLK(clk), .D(core__0v2_reg_63_0__46_), .Q(core_v2_reg_46_));
DFFPOSX1 DFFPOSX1_516 ( .CLK(clk), .D(core__0v2_reg_63_0__47_), .Q(core_v2_reg_47_));
DFFPOSX1 DFFPOSX1_517 ( .CLK(clk), .D(core__0v2_reg_63_0__48_), .Q(core_v2_reg_48_));
DFFPOSX1 DFFPOSX1_518 ( .CLK(clk), .D(core__0v2_reg_63_0__49_), .Q(core_v2_reg_49_));
DFFPOSX1 DFFPOSX1_519 ( .CLK(clk), .D(core__0v2_reg_63_0__50_), .Q(core_v2_reg_50_));
DFFPOSX1 DFFPOSX1_52 ( .CLK(clk), .D(_0key1_reg_31_0__7_), .Q(core_key_39_));
DFFPOSX1 DFFPOSX1_520 ( .CLK(clk), .D(core__0v2_reg_63_0__51_), .Q(core_v2_reg_51_));
DFFPOSX1 DFFPOSX1_521 ( .CLK(clk), .D(core__0v2_reg_63_0__52_), .Q(core_v2_reg_52_));
DFFPOSX1 DFFPOSX1_522 ( .CLK(clk), .D(core__0v2_reg_63_0__53_), .Q(core_v2_reg_53_));
DFFPOSX1 DFFPOSX1_523 ( .CLK(clk), .D(core__0v2_reg_63_0__54_), .Q(core_v2_reg_54_));
DFFPOSX1 DFFPOSX1_524 ( .CLK(clk), .D(core__0v2_reg_63_0__55_), .Q(core_v2_reg_55_));
DFFPOSX1 DFFPOSX1_525 ( .CLK(clk), .D(core__0v2_reg_63_0__56_), .Q(core_v2_reg_56_));
DFFPOSX1 DFFPOSX1_526 ( .CLK(clk), .D(core__0v2_reg_63_0__57_), .Q(core_v2_reg_57_));
DFFPOSX1 DFFPOSX1_527 ( .CLK(clk), .D(core__0v2_reg_63_0__58_), .Q(core_v2_reg_58_));
DFFPOSX1 DFFPOSX1_528 ( .CLK(clk), .D(core__0v2_reg_63_0__59_), .Q(core_v2_reg_59_));
DFFPOSX1 DFFPOSX1_529 ( .CLK(clk), .D(core__0v2_reg_63_0__60_), .Q(core_v2_reg_60_));
DFFPOSX1 DFFPOSX1_53 ( .CLK(clk), .D(_0key1_reg_31_0__8_), .Q(core_key_40_));
DFFPOSX1 DFFPOSX1_530 ( .CLK(clk), .D(core__0v2_reg_63_0__61_), .Q(core_v2_reg_61_));
DFFPOSX1 DFFPOSX1_531 ( .CLK(clk), .D(core__0v2_reg_63_0__62_), .Q(core_v2_reg_62_));
DFFPOSX1 DFFPOSX1_532 ( .CLK(clk), .D(core__0v2_reg_63_0__63_), .Q(core_v2_reg_63_));
DFFPOSX1 DFFPOSX1_533 ( .CLK(clk), .D(core__0v3_reg_63_0__0_), .Q(core_v3_reg_0_));
DFFPOSX1 DFFPOSX1_534 ( .CLK(clk), .D(core__0v3_reg_63_0__1_), .Q(core_v3_reg_1_));
DFFPOSX1 DFFPOSX1_535 ( .CLK(clk), .D(core__0v3_reg_63_0__2_), .Q(core_v3_reg_2_));
DFFPOSX1 DFFPOSX1_536 ( .CLK(clk), .D(core__0v3_reg_63_0__3_), .Q(core_v3_reg_3_));
DFFPOSX1 DFFPOSX1_537 ( .CLK(clk), .D(core__0v3_reg_63_0__4_), .Q(core_v3_reg_4_));
DFFPOSX1 DFFPOSX1_538 ( .CLK(clk), .D(core__0v3_reg_63_0__5_), .Q(core_v3_reg_5_));
DFFPOSX1 DFFPOSX1_539 ( .CLK(clk), .D(core__0v3_reg_63_0__6_), .Q(core_v3_reg_6_));
DFFPOSX1 DFFPOSX1_54 ( .CLK(clk), .D(_0key1_reg_31_0__9_), .Q(core_key_41_));
DFFPOSX1 DFFPOSX1_540 ( .CLK(clk), .D(core__0v3_reg_63_0__7_), .Q(core_v3_reg_7_));
DFFPOSX1 DFFPOSX1_541 ( .CLK(clk), .D(core__0v3_reg_63_0__8_), .Q(core_v3_reg_8_));
DFFPOSX1 DFFPOSX1_542 ( .CLK(clk), .D(core__0v3_reg_63_0__9_), .Q(core_v3_reg_9_));
DFFPOSX1 DFFPOSX1_543 ( .CLK(clk), .D(core__0v3_reg_63_0__10_), .Q(core_v3_reg_10_));
DFFPOSX1 DFFPOSX1_544 ( .CLK(clk), .D(core__0v3_reg_63_0__11_), .Q(core_v3_reg_11_));
DFFPOSX1 DFFPOSX1_545 ( .CLK(clk), .D(core__0v3_reg_63_0__12_), .Q(core_v3_reg_12_));
DFFPOSX1 DFFPOSX1_546 ( .CLK(clk), .D(core__0v3_reg_63_0__13_), .Q(core_v3_reg_13_));
DFFPOSX1 DFFPOSX1_547 ( .CLK(clk), .D(core__0v3_reg_63_0__14_), .Q(core_v3_reg_14_));
DFFPOSX1 DFFPOSX1_548 ( .CLK(clk), .D(core__0v3_reg_63_0__15_), .Q(core_v3_reg_15_));
DFFPOSX1 DFFPOSX1_549 ( .CLK(clk), .D(core__0v3_reg_63_0__16_), .Q(core_v3_reg_16_));
DFFPOSX1 DFFPOSX1_55 ( .CLK(clk), .D(_0key1_reg_31_0__10_), .Q(core_key_42_));
DFFPOSX1 DFFPOSX1_550 ( .CLK(clk), .D(core__0v3_reg_63_0__17_), .Q(core_v3_reg_17_));
DFFPOSX1 DFFPOSX1_551 ( .CLK(clk), .D(core__0v3_reg_63_0__18_), .Q(core_v3_reg_18_));
DFFPOSX1 DFFPOSX1_552 ( .CLK(clk), .D(core__0v3_reg_63_0__19_), .Q(core_v3_reg_19_));
DFFPOSX1 DFFPOSX1_553 ( .CLK(clk), .D(core__0v3_reg_63_0__20_), .Q(core_v3_reg_20_));
DFFPOSX1 DFFPOSX1_554 ( .CLK(clk), .D(core__0v3_reg_63_0__21_), .Q(core_v3_reg_21_));
DFFPOSX1 DFFPOSX1_555 ( .CLK(clk), .D(core__0v3_reg_63_0__22_), .Q(core_v3_reg_22_));
DFFPOSX1 DFFPOSX1_556 ( .CLK(clk), .D(core__0v3_reg_63_0__23_), .Q(core_v3_reg_23_));
DFFPOSX1 DFFPOSX1_557 ( .CLK(clk), .D(core__0v3_reg_63_0__24_), .Q(core_v3_reg_24_));
DFFPOSX1 DFFPOSX1_558 ( .CLK(clk), .D(core__0v3_reg_63_0__25_), .Q(core_v3_reg_25_));
DFFPOSX1 DFFPOSX1_559 ( .CLK(clk), .D(core__0v3_reg_63_0__26_), .Q(core_v3_reg_26_));
DFFPOSX1 DFFPOSX1_56 ( .CLK(clk), .D(_0key1_reg_31_0__11_), .Q(core_key_43_));
DFFPOSX1 DFFPOSX1_560 ( .CLK(clk), .D(core__0v3_reg_63_0__27_), .Q(core_v3_reg_27_));
DFFPOSX1 DFFPOSX1_561 ( .CLK(clk), .D(core__0v3_reg_63_0__28_), .Q(core_v3_reg_28_));
DFFPOSX1 DFFPOSX1_562 ( .CLK(clk), .D(core__0v3_reg_63_0__29_), .Q(core_v3_reg_29_));
DFFPOSX1 DFFPOSX1_563 ( .CLK(clk), .D(core__0v3_reg_63_0__30_), .Q(core_v3_reg_30_));
DFFPOSX1 DFFPOSX1_564 ( .CLK(clk), .D(core__0v3_reg_63_0__31_), .Q(core_v3_reg_31_));
DFFPOSX1 DFFPOSX1_565 ( .CLK(clk), .D(core__0v3_reg_63_0__32_), .Q(core_v3_reg_32_));
DFFPOSX1 DFFPOSX1_566 ( .CLK(clk), .D(core__0v3_reg_63_0__33_), .Q(core_v3_reg_33_));
DFFPOSX1 DFFPOSX1_567 ( .CLK(clk), .D(core__0v3_reg_63_0__34_), .Q(core_v3_reg_34_));
DFFPOSX1 DFFPOSX1_568 ( .CLK(clk), .D(core__0v3_reg_63_0__35_), .Q(core_v3_reg_35_));
DFFPOSX1 DFFPOSX1_569 ( .CLK(clk), .D(core__0v3_reg_63_0__36_), .Q(core_v3_reg_36_));
DFFPOSX1 DFFPOSX1_57 ( .CLK(clk), .D(_0key1_reg_31_0__12_), .Q(core_key_44_));
DFFPOSX1 DFFPOSX1_570 ( .CLK(clk), .D(core__0v3_reg_63_0__37_), .Q(core_v3_reg_37_));
DFFPOSX1 DFFPOSX1_571 ( .CLK(clk), .D(core__0v3_reg_63_0__38_), .Q(core_v3_reg_38_));
DFFPOSX1 DFFPOSX1_572 ( .CLK(clk), .D(core__0v3_reg_63_0__39_), .Q(core_v3_reg_39_));
DFFPOSX1 DFFPOSX1_573 ( .CLK(clk), .D(core__0v3_reg_63_0__40_), .Q(core_v3_reg_40_));
DFFPOSX1 DFFPOSX1_574 ( .CLK(clk), .D(core__0v3_reg_63_0__41_), .Q(core_v3_reg_41_));
DFFPOSX1 DFFPOSX1_575 ( .CLK(clk), .D(core__0v3_reg_63_0__42_), .Q(core_v3_reg_42_));
DFFPOSX1 DFFPOSX1_576 ( .CLK(clk), .D(core__0v3_reg_63_0__43_), .Q(core_v3_reg_43_));
DFFPOSX1 DFFPOSX1_577 ( .CLK(clk), .D(core__0v3_reg_63_0__44_), .Q(core_v3_reg_44_));
DFFPOSX1 DFFPOSX1_578 ( .CLK(clk), .D(core__0v3_reg_63_0__45_), .Q(core_v3_reg_45_));
DFFPOSX1 DFFPOSX1_579 ( .CLK(clk), .D(core__0v3_reg_63_0__46_), .Q(core_v3_reg_46_));
DFFPOSX1 DFFPOSX1_58 ( .CLK(clk), .D(_0key1_reg_31_0__13_), .Q(core_key_45_));
DFFPOSX1 DFFPOSX1_580 ( .CLK(clk), .D(core__0v3_reg_63_0__47_), .Q(core_v3_reg_47_));
DFFPOSX1 DFFPOSX1_581 ( .CLK(clk), .D(core__0v3_reg_63_0__48_), .Q(core_v3_reg_48_));
DFFPOSX1 DFFPOSX1_582 ( .CLK(clk), .D(core__0v3_reg_63_0__49_), .Q(core_v3_reg_49_));
DFFPOSX1 DFFPOSX1_583 ( .CLK(clk), .D(core__0v3_reg_63_0__50_), .Q(core_v3_reg_50_));
DFFPOSX1 DFFPOSX1_584 ( .CLK(clk), .D(core__0v3_reg_63_0__51_), .Q(core_v3_reg_51_));
DFFPOSX1 DFFPOSX1_585 ( .CLK(clk), .D(core__0v3_reg_63_0__52_), .Q(core_v3_reg_52_));
DFFPOSX1 DFFPOSX1_586 ( .CLK(clk), .D(core__0v3_reg_63_0__53_), .Q(core_v3_reg_53_));
DFFPOSX1 DFFPOSX1_587 ( .CLK(clk), .D(core__0v3_reg_63_0__54_), .Q(core_v3_reg_54_));
DFFPOSX1 DFFPOSX1_588 ( .CLK(clk), .D(core__0v3_reg_63_0__55_), .Q(core_v3_reg_55_));
DFFPOSX1 DFFPOSX1_589 ( .CLK(clk), .D(core__0v3_reg_63_0__56_), .Q(core_v3_reg_56_));
DFFPOSX1 DFFPOSX1_59 ( .CLK(clk), .D(_0key1_reg_31_0__14_), .Q(core_key_46_));
DFFPOSX1 DFFPOSX1_590 ( .CLK(clk), .D(core__0v3_reg_63_0__57_), .Q(core_v3_reg_57_));
DFFPOSX1 DFFPOSX1_591 ( .CLK(clk), .D(core__0v3_reg_63_0__58_), .Q(core_v3_reg_58_));
DFFPOSX1 DFFPOSX1_592 ( .CLK(clk), .D(core__0v3_reg_63_0__59_), .Q(core_v3_reg_59_));
DFFPOSX1 DFFPOSX1_593 ( .CLK(clk), .D(core__0v3_reg_63_0__60_), .Q(core_v3_reg_60_));
DFFPOSX1 DFFPOSX1_594 ( .CLK(clk), .D(core__0v3_reg_63_0__61_), .Q(core_v3_reg_61_));
DFFPOSX1 DFFPOSX1_595 ( .CLK(clk), .D(core__0v3_reg_63_0__62_), .Q(core_v3_reg_62_));
DFFPOSX1 DFFPOSX1_596 ( .CLK(clk), .D(core__0v3_reg_63_0__63_), .Q(core_v3_reg_63_));
DFFPOSX1 DFFPOSX1_597 ( .CLK(clk), .D(core__0mi_reg_63_0__0_), .Q(core_mi_reg_0_));
DFFPOSX1 DFFPOSX1_598 ( .CLK(clk), .D(core__0mi_reg_63_0__1_), .Q(core_mi_reg_1_));
DFFPOSX1 DFFPOSX1_599 ( .CLK(clk), .D(core__0mi_reg_63_0__2_), .Q(core_mi_reg_2_));
DFFPOSX1 DFFPOSX1_6 ( .CLK(clk), .D(_0param_reg_7_0__1_), .Q(core_compression_rounds_1_));
DFFPOSX1 DFFPOSX1_60 ( .CLK(clk), .D(_0key1_reg_31_0__15_), .Q(core_key_47_));
DFFPOSX1 DFFPOSX1_600 ( .CLK(clk), .D(core__0mi_reg_63_0__3_), .Q(core_mi_reg_3_));
DFFPOSX1 DFFPOSX1_601 ( .CLK(clk), .D(core__0mi_reg_63_0__4_), .Q(core_mi_reg_4_));
DFFPOSX1 DFFPOSX1_602 ( .CLK(clk), .D(core__0mi_reg_63_0__5_), .Q(core_mi_reg_5_));
DFFPOSX1 DFFPOSX1_603 ( .CLK(clk), .D(core__0mi_reg_63_0__6_), .Q(core_mi_reg_6_));
DFFPOSX1 DFFPOSX1_604 ( .CLK(clk), .D(core__0mi_reg_63_0__7_), .Q(core_mi_reg_7_));
DFFPOSX1 DFFPOSX1_605 ( .CLK(clk), .D(core__0mi_reg_63_0__8_), .Q(core_mi_reg_8_));
DFFPOSX1 DFFPOSX1_606 ( .CLK(clk), .D(core__0mi_reg_63_0__9_), .Q(core_mi_reg_9_));
DFFPOSX1 DFFPOSX1_607 ( .CLK(clk), .D(core__0mi_reg_63_0__10_), .Q(core_mi_reg_10_));
DFFPOSX1 DFFPOSX1_608 ( .CLK(clk), .D(core__0mi_reg_63_0__11_), .Q(core_mi_reg_11_));
DFFPOSX1 DFFPOSX1_609 ( .CLK(clk), .D(core__0mi_reg_63_0__12_), .Q(core_mi_reg_12_));
DFFPOSX1 DFFPOSX1_61 ( .CLK(clk), .D(_0key1_reg_31_0__16_), .Q(core_key_48_));
DFFPOSX1 DFFPOSX1_610 ( .CLK(clk), .D(core__0mi_reg_63_0__13_), .Q(core_mi_reg_13_));
DFFPOSX1 DFFPOSX1_611 ( .CLK(clk), .D(core__0mi_reg_63_0__14_), .Q(core_mi_reg_14_));
DFFPOSX1 DFFPOSX1_612 ( .CLK(clk), .D(core__0mi_reg_63_0__15_), .Q(core_mi_reg_15_));
DFFPOSX1 DFFPOSX1_613 ( .CLK(clk), .D(core__0mi_reg_63_0__16_), .Q(core_mi_reg_16_));
DFFPOSX1 DFFPOSX1_614 ( .CLK(clk), .D(core__0mi_reg_63_0__17_), .Q(core_mi_reg_17_));
DFFPOSX1 DFFPOSX1_615 ( .CLK(clk), .D(core__0mi_reg_63_0__18_), .Q(core_mi_reg_18_));
DFFPOSX1 DFFPOSX1_616 ( .CLK(clk), .D(core__0mi_reg_63_0__19_), .Q(core_mi_reg_19_));
DFFPOSX1 DFFPOSX1_617 ( .CLK(clk), .D(core__0mi_reg_63_0__20_), .Q(core_mi_reg_20_));
DFFPOSX1 DFFPOSX1_618 ( .CLK(clk), .D(core__0mi_reg_63_0__21_), .Q(core_mi_reg_21_));
DFFPOSX1 DFFPOSX1_619 ( .CLK(clk), .D(core__0mi_reg_63_0__22_), .Q(core_mi_reg_22_));
DFFPOSX1 DFFPOSX1_62 ( .CLK(clk), .D(_0key1_reg_31_0__17_), .Q(core_key_49_));
DFFPOSX1 DFFPOSX1_620 ( .CLK(clk), .D(core__0mi_reg_63_0__23_), .Q(core_mi_reg_23_));
DFFPOSX1 DFFPOSX1_621 ( .CLK(clk), .D(core__0mi_reg_63_0__24_), .Q(core_mi_reg_24_));
DFFPOSX1 DFFPOSX1_622 ( .CLK(clk), .D(core__0mi_reg_63_0__25_), .Q(core_mi_reg_25_));
DFFPOSX1 DFFPOSX1_623 ( .CLK(clk), .D(core__0mi_reg_63_0__26_), .Q(core_mi_reg_26_));
DFFPOSX1 DFFPOSX1_624 ( .CLK(clk), .D(core__0mi_reg_63_0__27_), .Q(core_mi_reg_27_));
DFFPOSX1 DFFPOSX1_625 ( .CLK(clk), .D(core__0mi_reg_63_0__28_), .Q(core_mi_reg_28_));
DFFPOSX1 DFFPOSX1_626 ( .CLK(clk), .D(core__0mi_reg_63_0__29_), .Q(core_mi_reg_29_));
DFFPOSX1 DFFPOSX1_627 ( .CLK(clk), .D(core__0mi_reg_63_0__30_), .Q(core_mi_reg_30_));
DFFPOSX1 DFFPOSX1_628 ( .CLK(clk), .D(core__0mi_reg_63_0__31_), .Q(core_mi_reg_31_));
DFFPOSX1 DFFPOSX1_629 ( .CLK(clk), .D(core__0mi_reg_63_0__32_), .Q(core_mi_reg_32_));
DFFPOSX1 DFFPOSX1_63 ( .CLK(clk), .D(_0key1_reg_31_0__18_), .Q(core_key_50_));
DFFPOSX1 DFFPOSX1_630 ( .CLK(clk), .D(core__0mi_reg_63_0__33_), .Q(core_mi_reg_33_));
DFFPOSX1 DFFPOSX1_631 ( .CLK(clk), .D(core__0mi_reg_63_0__34_), .Q(core_mi_reg_34_));
DFFPOSX1 DFFPOSX1_632 ( .CLK(clk), .D(core__0mi_reg_63_0__35_), .Q(core_mi_reg_35_));
DFFPOSX1 DFFPOSX1_633 ( .CLK(clk), .D(core__0mi_reg_63_0__36_), .Q(core_mi_reg_36_));
DFFPOSX1 DFFPOSX1_634 ( .CLK(clk), .D(core__0mi_reg_63_0__37_), .Q(core_mi_reg_37_));
DFFPOSX1 DFFPOSX1_635 ( .CLK(clk), .D(core__0mi_reg_63_0__38_), .Q(core_mi_reg_38_));
DFFPOSX1 DFFPOSX1_636 ( .CLK(clk), .D(core__0mi_reg_63_0__39_), .Q(core_mi_reg_39_));
DFFPOSX1 DFFPOSX1_637 ( .CLK(clk), .D(core__0mi_reg_63_0__40_), .Q(core_mi_reg_40_));
DFFPOSX1 DFFPOSX1_638 ( .CLK(clk), .D(core__0mi_reg_63_0__41_), .Q(core_mi_reg_41_));
DFFPOSX1 DFFPOSX1_639 ( .CLK(clk), .D(core__0mi_reg_63_0__42_), .Q(core_mi_reg_42_));
DFFPOSX1 DFFPOSX1_64 ( .CLK(clk), .D(_0key1_reg_31_0__19_), .Q(core_key_51_));
DFFPOSX1 DFFPOSX1_640 ( .CLK(clk), .D(core__0mi_reg_63_0__43_), .Q(core_mi_reg_43_));
DFFPOSX1 DFFPOSX1_641 ( .CLK(clk), .D(core__0mi_reg_63_0__44_), .Q(core_mi_reg_44_));
DFFPOSX1 DFFPOSX1_642 ( .CLK(clk), .D(core__0mi_reg_63_0__45_), .Q(core_mi_reg_45_));
DFFPOSX1 DFFPOSX1_643 ( .CLK(clk), .D(core__0mi_reg_63_0__46_), .Q(core_mi_reg_46_));
DFFPOSX1 DFFPOSX1_644 ( .CLK(clk), .D(core__0mi_reg_63_0__47_), .Q(core_mi_reg_47_));
DFFPOSX1 DFFPOSX1_645 ( .CLK(clk), .D(core__0mi_reg_63_0__48_), .Q(core_mi_reg_48_));
DFFPOSX1 DFFPOSX1_646 ( .CLK(clk), .D(core__0mi_reg_63_0__49_), .Q(core_mi_reg_49_));
DFFPOSX1 DFFPOSX1_647 ( .CLK(clk), .D(core__0mi_reg_63_0__50_), .Q(core_mi_reg_50_));
DFFPOSX1 DFFPOSX1_648 ( .CLK(clk), .D(core__0mi_reg_63_0__51_), .Q(core_mi_reg_51_));
DFFPOSX1 DFFPOSX1_649 ( .CLK(clk), .D(core__0mi_reg_63_0__52_), .Q(core_mi_reg_52_));
DFFPOSX1 DFFPOSX1_65 ( .CLK(clk), .D(_0key1_reg_31_0__20_), .Q(core_key_52_));
DFFPOSX1 DFFPOSX1_650 ( .CLK(clk), .D(core__0mi_reg_63_0__53_), .Q(core_mi_reg_53_));
DFFPOSX1 DFFPOSX1_651 ( .CLK(clk), .D(core__0mi_reg_63_0__54_), .Q(core_mi_reg_54_));
DFFPOSX1 DFFPOSX1_652 ( .CLK(clk), .D(core__0mi_reg_63_0__55_), .Q(core_mi_reg_55_));
DFFPOSX1 DFFPOSX1_653 ( .CLK(clk), .D(core__0mi_reg_63_0__56_), .Q(core_mi_reg_56_));
DFFPOSX1 DFFPOSX1_654 ( .CLK(clk), .D(core__0mi_reg_63_0__57_), .Q(core_mi_reg_57_));
DFFPOSX1 DFFPOSX1_655 ( .CLK(clk), .D(core__0mi_reg_63_0__58_), .Q(core_mi_reg_58_));
DFFPOSX1 DFFPOSX1_656 ( .CLK(clk), .D(core__0mi_reg_63_0__59_), .Q(core_mi_reg_59_));
DFFPOSX1 DFFPOSX1_657 ( .CLK(clk), .D(core__0mi_reg_63_0__60_), .Q(core_mi_reg_60_));
DFFPOSX1 DFFPOSX1_658 ( .CLK(clk), .D(core__0mi_reg_63_0__61_), .Q(core_mi_reg_61_));
DFFPOSX1 DFFPOSX1_659 ( .CLK(clk), .D(core__0mi_reg_63_0__62_), .Q(core_mi_reg_62_));
DFFPOSX1 DFFPOSX1_66 ( .CLK(clk), .D(_0key1_reg_31_0__21_), .Q(core_key_53_));
DFFPOSX1 DFFPOSX1_660 ( .CLK(clk), .D(core__0mi_reg_63_0__63_), .Q(core_mi_reg_63_));
DFFPOSX1 DFFPOSX1_661 ( .CLK(clk), .D(core__0loop_ctr_reg_3_0__0_), .Q(core_loop_ctr_reg_0_));
DFFPOSX1 DFFPOSX1_662 ( .CLK(clk), .D(core__0loop_ctr_reg_3_0__1_), .Q(core_loop_ctr_reg_1_));
DFFPOSX1 DFFPOSX1_663 ( .CLK(clk), .D(core__0loop_ctr_reg_3_0__2_), .Q(core_loop_ctr_reg_2_));
DFFPOSX1 DFFPOSX1_664 ( .CLK(clk), .D(core__0loop_ctr_reg_3_0__3_), .Q(core_loop_ctr_reg_3_));
DFFPOSX1 DFFPOSX1_665 ( .CLK(clk), .D(core__0ready_reg_0_0_), .Q(core_ready));
DFFPOSX1 DFFPOSX1_666 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__0_), .Q(core_siphash_word_0_));
DFFPOSX1 DFFPOSX1_667 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__1_), .Q(core_siphash_word_1_));
DFFPOSX1 DFFPOSX1_668 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__2_), .Q(core_siphash_word_2_));
DFFPOSX1 DFFPOSX1_669 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__3_), .Q(core_siphash_word_3_));
DFFPOSX1 DFFPOSX1_67 ( .CLK(clk), .D(_0key1_reg_31_0__22_), .Q(core_key_54_));
DFFPOSX1 DFFPOSX1_670 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__4_), .Q(core_siphash_word_4_));
DFFPOSX1 DFFPOSX1_671 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__5_), .Q(core_siphash_word_5_));
DFFPOSX1 DFFPOSX1_672 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__6_), .Q(core_siphash_word_6_));
DFFPOSX1 DFFPOSX1_673 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__7_), .Q(core_siphash_word_7_));
DFFPOSX1 DFFPOSX1_674 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__8_), .Q(core_siphash_word_8_));
DFFPOSX1 DFFPOSX1_675 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__9_), .Q(core_siphash_word_9_));
DFFPOSX1 DFFPOSX1_676 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__10_), .Q(core_siphash_word_10_));
DFFPOSX1 DFFPOSX1_677 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__11_), .Q(core_siphash_word_11_));
DFFPOSX1 DFFPOSX1_678 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__12_), .Q(core_siphash_word_12_));
DFFPOSX1 DFFPOSX1_679 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__13_), .Q(core_siphash_word_13_));
DFFPOSX1 DFFPOSX1_68 ( .CLK(clk), .D(_0key1_reg_31_0__23_), .Q(core_key_55_));
DFFPOSX1 DFFPOSX1_680 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__14_), .Q(core_siphash_word_14_));
DFFPOSX1 DFFPOSX1_681 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__15_), .Q(core_siphash_word_15_));
DFFPOSX1 DFFPOSX1_682 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__16_), .Q(core_siphash_word_16_));
DFFPOSX1 DFFPOSX1_683 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__17_), .Q(core_siphash_word_17_));
DFFPOSX1 DFFPOSX1_684 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__18_), .Q(core_siphash_word_18_));
DFFPOSX1 DFFPOSX1_685 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__19_), .Q(core_siphash_word_19_));
DFFPOSX1 DFFPOSX1_686 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__20_), .Q(core_siphash_word_20_));
DFFPOSX1 DFFPOSX1_687 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__21_), .Q(core_siphash_word_21_));
DFFPOSX1 DFFPOSX1_688 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__22_), .Q(core_siphash_word_22_));
DFFPOSX1 DFFPOSX1_689 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__23_), .Q(core_siphash_word_23_));
DFFPOSX1 DFFPOSX1_69 ( .CLK(clk), .D(_0key1_reg_31_0__24_), .Q(core_key_56_));
DFFPOSX1 DFFPOSX1_690 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__24_), .Q(core_siphash_word_24_));
DFFPOSX1 DFFPOSX1_691 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__25_), .Q(core_siphash_word_25_));
DFFPOSX1 DFFPOSX1_692 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__26_), .Q(core_siphash_word_26_));
DFFPOSX1 DFFPOSX1_693 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__27_), .Q(core_siphash_word_27_));
DFFPOSX1 DFFPOSX1_694 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__28_), .Q(core_siphash_word_28_));
DFFPOSX1 DFFPOSX1_695 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__29_), .Q(core_siphash_word_29_));
DFFPOSX1 DFFPOSX1_696 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__30_), .Q(core_siphash_word_30_));
DFFPOSX1 DFFPOSX1_697 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__31_), .Q(core_siphash_word_31_));
DFFPOSX1 DFFPOSX1_698 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__32_), .Q(core_siphash_word_32_));
DFFPOSX1 DFFPOSX1_699 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__33_), .Q(core_siphash_word_33_));
DFFPOSX1 DFFPOSX1_7 ( .CLK(clk), .D(_0param_reg_7_0__2_), .Q(core_compression_rounds_2_));
DFFPOSX1 DFFPOSX1_70 ( .CLK(clk), .D(_0key1_reg_31_0__25_), .Q(core_key_57_));
DFFPOSX1 DFFPOSX1_700 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__34_), .Q(core_siphash_word_34_));
DFFPOSX1 DFFPOSX1_701 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__35_), .Q(core_siphash_word_35_));
DFFPOSX1 DFFPOSX1_702 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__36_), .Q(core_siphash_word_36_));
DFFPOSX1 DFFPOSX1_703 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__37_), .Q(core_siphash_word_37_));
DFFPOSX1 DFFPOSX1_704 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__38_), .Q(core_siphash_word_38_));
DFFPOSX1 DFFPOSX1_705 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__39_), .Q(core_siphash_word_39_));
DFFPOSX1 DFFPOSX1_706 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__40_), .Q(core_siphash_word_40_));
DFFPOSX1 DFFPOSX1_707 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__41_), .Q(core_siphash_word_41_));
DFFPOSX1 DFFPOSX1_708 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__42_), .Q(core_siphash_word_42_));
DFFPOSX1 DFFPOSX1_709 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__43_), .Q(core_siphash_word_43_));
DFFPOSX1 DFFPOSX1_71 ( .CLK(clk), .D(_0key1_reg_31_0__26_), .Q(core_key_58_));
DFFPOSX1 DFFPOSX1_710 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__44_), .Q(core_siphash_word_44_));
DFFPOSX1 DFFPOSX1_711 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__45_), .Q(core_siphash_word_45_));
DFFPOSX1 DFFPOSX1_712 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__46_), .Q(core_siphash_word_46_));
DFFPOSX1 DFFPOSX1_713 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__47_), .Q(core_siphash_word_47_));
DFFPOSX1 DFFPOSX1_714 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__48_), .Q(core_siphash_word_48_));
DFFPOSX1 DFFPOSX1_715 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__49_), .Q(core_siphash_word_49_));
DFFPOSX1 DFFPOSX1_716 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__50_), .Q(core_siphash_word_50_));
DFFPOSX1 DFFPOSX1_717 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__51_), .Q(core_siphash_word_51_));
DFFPOSX1 DFFPOSX1_718 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__52_), .Q(core_siphash_word_52_));
DFFPOSX1 DFFPOSX1_719 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__53_), .Q(core_siphash_word_53_));
DFFPOSX1 DFFPOSX1_72 ( .CLK(clk), .D(_0key1_reg_31_0__27_), .Q(core_key_59_));
DFFPOSX1 DFFPOSX1_720 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__54_), .Q(core_siphash_word_54_));
DFFPOSX1 DFFPOSX1_721 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__55_), .Q(core_siphash_word_55_));
DFFPOSX1 DFFPOSX1_722 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__56_), .Q(core_siphash_word_56_));
DFFPOSX1 DFFPOSX1_723 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__57_), .Q(core_siphash_word_57_));
DFFPOSX1 DFFPOSX1_724 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__58_), .Q(core_siphash_word_58_));
DFFPOSX1 DFFPOSX1_725 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__59_), .Q(core_siphash_word_59_));
DFFPOSX1 DFFPOSX1_726 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__60_), .Q(core_siphash_word_60_));
DFFPOSX1 DFFPOSX1_727 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__61_), .Q(core_siphash_word_61_));
DFFPOSX1 DFFPOSX1_728 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__62_), .Q(core_siphash_word_62_));
DFFPOSX1 DFFPOSX1_729 ( .CLK(clk), .D(core__0siphash_word0_reg_63_0__63_), .Q(core_siphash_word_63_));
DFFPOSX1 DFFPOSX1_73 ( .CLK(clk), .D(_0key1_reg_31_0__28_), .Q(core_key_60_));
DFFPOSX1 DFFPOSX1_730 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__0_), .Q(core_siphash_word_64_));
DFFPOSX1 DFFPOSX1_731 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__1_), .Q(core_siphash_word_65_));
DFFPOSX1 DFFPOSX1_732 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__2_), .Q(core_siphash_word_66_));
DFFPOSX1 DFFPOSX1_733 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__3_), .Q(core_siphash_word_67_));
DFFPOSX1 DFFPOSX1_734 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__4_), .Q(core_siphash_word_68_));
DFFPOSX1 DFFPOSX1_735 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__5_), .Q(core_siphash_word_69_));
DFFPOSX1 DFFPOSX1_736 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__6_), .Q(core_siphash_word_70_));
DFFPOSX1 DFFPOSX1_737 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__7_), .Q(core_siphash_word_71_));
DFFPOSX1 DFFPOSX1_738 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__8_), .Q(core_siphash_word_72_));
DFFPOSX1 DFFPOSX1_739 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__9_), .Q(core_siphash_word_73_));
DFFPOSX1 DFFPOSX1_74 ( .CLK(clk), .D(_0key1_reg_31_0__29_), .Q(core_key_61_));
DFFPOSX1 DFFPOSX1_740 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__10_), .Q(core_siphash_word_74_));
DFFPOSX1 DFFPOSX1_741 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__11_), .Q(core_siphash_word_75_));
DFFPOSX1 DFFPOSX1_742 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__12_), .Q(core_siphash_word_76_));
DFFPOSX1 DFFPOSX1_743 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__13_), .Q(core_siphash_word_77_));
DFFPOSX1 DFFPOSX1_744 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__14_), .Q(core_siphash_word_78_));
DFFPOSX1 DFFPOSX1_745 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__15_), .Q(core_siphash_word_79_));
DFFPOSX1 DFFPOSX1_746 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__16_), .Q(core_siphash_word_80_));
DFFPOSX1 DFFPOSX1_747 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__17_), .Q(core_siphash_word_81_));
DFFPOSX1 DFFPOSX1_748 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__18_), .Q(core_siphash_word_82_));
DFFPOSX1 DFFPOSX1_749 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__19_), .Q(core_siphash_word_83_));
DFFPOSX1 DFFPOSX1_75 ( .CLK(clk), .D(_0key1_reg_31_0__30_), .Q(core_key_62_));
DFFPOSX1 DFFPOSX1_750 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__20_), .Q(core_siphash_word_84_));
DFFPOSX1 DFFPOSX1_751 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__21_), .Q(core_siphash_word_85_));
DFFPOSX1 DFFPOSX1_752 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__22_), .Q(core_siphash_word_86_));
DFFPOSX1 DFFPOSX1_753 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__23_), .Q(core_siphash_word_87_));
DFFPOSX1 DFFPOSX1_754 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__24_), .Q(core_siphash_word_88_));
DFFPOSX1 DFFPOSX1_755 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__25_), .Q(core_siphash_word_89_));
DFFPOSX1 DFFPOSX1_756 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__26_), .Q(core_siphash_word_90_));
DFFPOSX1 DFFPOSX1_757 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__27_), .Q(core_siphash_word_91_));
DFFPOSX1 DFFPOSX1_758 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__28_), .Q(core_siphash_word_92_));
DFFPOSX1 DFFPOSX1_759 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__29_), .Q(core_siphash_word_93_));
DFFPOSX1 DFFPOSX1_76 ( .CLK(clk), .D(_0key1_reg_31_0__31_), .Q(core_key_63_));
DFFPOSX1 DFFPOSX1_760 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__30_), .Q(core_siphash_word_94_));
DFFPOSX1 DFFPOSX1_761 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__31_), .Q(core_siphash_word_95_));
DFFPOSX1 DFFPOSX1_762 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__32_), .Q(core_siphash_word_96_));
DFFPOSX1 DFFPOSX1_763 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__33_), .Q(core_siphash_word_97_));
DFFPOSX1 DFFPOSX1_764 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__34_), .Q(core_siphash_word_98_));
DFFPOSX1 DFFPOSX1_765 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__35_), .Q(core_siphash_word_99_));
DFFPOSX1 DFFPOSX1_766 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__36_), .Q(core_siphash_word_100_));
DFFPOSX1 DFFPOSX1_767 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__37_), .Q(core_siphash_word_101_));
DFFPOSX1 DFFPOSX1_768 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__38_), .Q(core_siphash_word_102_));
DFFPOSX1 DFFPOSX1_769 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__39_), .Q(core_siphash_word_103_));
DFFPOSX1 DFFPOSX1_77 ( .CLK(clk), .D(_0key2_reg_31_0__0_), .Q(core_key_64_));
DFFPOSX1 DFFPOSX1_770 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__40_), .Q(core_siphash_word_104_));
DFFPOSX1 DFFPOSX1_771 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__41_), .Q(core_siphash_word_105_));
DFFPOSX1 DFFPOSX1_772 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__42_), .Q(core_siphash_word_106_));
DFFPOSX1 DFFPOSX1_773 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__43_), .Q(core_siphash_word_107_));
DFFPOSX1 DFFPOSX1_774 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__44_), .Q(core_siphash_word_108_));
DFFPOSX1 DFFPOSX1_775 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__45_), .Q(core_siphash_word_109_));
DFFPOSX1 DFFPOSX1_776 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__46_), .Q(core_siphash_word_110_));
DFFPOSX1 DFFPOSX1_777 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__47_), .Q(core_siphash_word_111_));
DFFPOSX1 DFFPOSX1_778 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__48_), .Q(core_siphash_word_112_));
DFFPOSX1 DFFPOSX1_779 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__49_), .Q(core_siphash_word_113_));
DFFPOSX1 DFFPOSX1_78 ( .CLK(clk), .D(_0key2_reg_31_0__1_), .Q(core_key_65_));
DFFPOSX1 DFFPOSX1_780 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__50_), .Q(core_siphash_word_114_));
DFFPOSX1 DFFPOSX1_781 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__51_), .Q(core_siphash_word_115_));
DFFPOSX1 DFFPOSX1_782 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__52_), .Q(core_siphash_word_116_));
DFFPOSX1 DFFPOSX1_783 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__53_), .Q(core_siphash_word_117_));
DFFPOSX1 DFFPOSX1_784 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__54_), .Q(core_siphash_word_118_));
DFFPOSX1 DFFPOSX1_785 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__55_), .Q(core_siphash_word_119_));
DFFPOSX1 DFFPOSX1_786 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__56_), .Q(core_siphash_word_120_));
DFFPOSX1 DFFPOSX1_787 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__57_), .Q(core_siphash_word_121_));
DFFPOSX1 DFFPOSX1_788 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__58_), .Q(core_siphash_word_122_));
DFFPOSX1 DFFPOSX1_789 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__59_), .Q(core_siphash_word_123_));
DFFPOSX1 DFFPOSX1_79 ( .CLK(clk), .D(_0key2_reg_31_0__2_), .Q(core_key_66_));
DFFPOSX1 DFFPOSX1_790 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__60_), .Q(core_siphash_word_124_));
DFFPOSX1 DFFPOSX1_791 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__61_), .Q(core_siphash_word_125_));
DFFPOSX1 DFFPOSX1_792 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__62_), .Q(core_siphash_word_126_));
DFFPOSX1 DFFPOSX1_793 ( .CLK(clk), .D(core__0siphash_word1_reg_63_0__63_), .Q(core_siphash_word_127_));
DFFPOSX1 DFFPOSX1_794 ( .CLK(clk), .D(core__0siphash_valid_reg_0_0_), .Q(core_siphash_valid_reg));
DFFPOSX1 DFFPOSX1_8 ( .CLK(clk), .D(_0param_reg_7_0__3_), .Q(core_compression_rounds_3_));
DFFPOSX1 DFFPOSX1_80 ( .CLK(clk), .D(_0key2_reg_31_0__3_), .Q(core_key_67_));
DFFPOSX1 DFFPOSX1_81 ( .CLK(clk), .D(_0key2_reg_31_0__4_), .Q(core_key_68_));
DFFPOSX1 DFFPOSX1_82 ( .CLK(clk), .D(_0key2_reg_31_0__5_), .Q(core_key_69_));
DFFPOSX1 DFFPOSX1_83 ( .CLK(clk), .D(_0key2_reg_31_0__6_), .Q(core_key_70_));
DFFPOSX1 DFFPOSX1_84 ( .CLK(clk), .D(_0key2_reg_31_0__7_), .Q(core_key_71_));
DFFPOSX1 DFFPOSX1_85 ( .CLK(clk), .D(_0key2_reg_31_0__8_), .Q(core_key_72_));
DFFPOSX1 DFFPOSX1_86 ( .CLK(clk), .D(_0key2_reg_31_0__9_), .Q(core_key_73_));
DFFPOSX1 DFFPOSX1_87 ( .CLK(clk), .D(_0key2_reg_31_0__10_), .Q(core_key_74_));
DFFPOSX1 DFFPOSX1_88 ( .CLK(clk), .D(_0key2_reg_31_0__11_), .Q(core_key_75_));
DFFPOSX1 DFFPOSX1_89 ( .CLK(clk), .D(_0key2_reg_31_0__12_), .Q(core_key_76_));
DFFPOSX1 DFFPOSX1_9 ( .CLK(clk), .D(_0param_reg_7_0__4_), .Q(core_final_rounds_0_));
DFFPOSX1 DFFPOSX1_90 ( .CLK(clk), .D(_0key2_reg_31_0__13_), .Q(core_key_77_));
DFFPOSX1 DFFPOSX1_91 ( .CLK(clk), .D(_0key2_reg_31_0__14_), .Q(core_key_78_));
DFFPOSX1 DFFPOSX1_92 ( .CLK(clk), .D(_0key2_reg_31_0__15_), .Q(core_key_79_));
DFFPOSX1 DFFPOSX1_93 ( .CLK(clk), .D(_0key2_reg_31_0__16_), .Q(core_key_80_));
DFFPOSX1 DFFPOSX1_94 ( .CLK(clk), .D(_0key2_reg_31_0__17_), .Q(core_key_81_));
DFFPOSX1 DFFPOSX1_95 ( .CLK(clk), .D(_0key2_reg_31_0__18_), .Q(core_key_82_));
DFFPOSX1 DFFPOSX1_96 ( .CLK(clk), .D(_0key2_reg_31_0__19_), .Q(core_key_83_));
DFFPOSX1 DFFPOSX1_97 ( .CLK(clk), .D(_0key2_reg_31_0__20_), .Q(core_key_84_));
DFFPOSX1 DFFPOSX1_98 ( .CLK(clk), .D(_0key2_reg_31_0__21_), .Q(core_key_85_));
DFFPOSX1 DFFPOSX1_99 ( .CLK(clk), .D(_0key2_reg_31_0__22_), .Q(core_key_86_));
INVX1 INVX1_1 ( .A(\addr[7] ), .Y(_abc_19873_new_n870_));
INVX1 INVX1_10 ( .A(core_siphash_valid_reg), .Y(_abc_19873_new_n1607_));
INVX1 INVX1_100 ( .A(_abc_19873_new_n2440_), .Y(_abc_19873_new_n2441_));
INVX1 INVX1_1000 ( .A(core__abc_22172_new_n4806_), .Y(core__abc_22172_new_n4831_));
INVX1 INVX1_1001 ( .A(core__abc_22172_new_n4833_), .Y(core__abc_22172_new_n4834_));
INVX1 INVX1_1002 ( .A(core__abc_22172_new_n4838_), .Y(core__abc_22172_new_n4839_));
INVX1 INVX1_1003 ( .A(core__abc_22172_new_n4843_), .Y(core__abc_22172_new_n4844_));
INVX1 INVX1_1004 ( .A(core__abc_22172_new_n4837_), .Y(core__abc_22172_new_n4848_));
INVX1 INVX1_1005 ( .A(core__abc_22172_new_n4846_), .Y(core__abc_22172_new_n4849_));
INVX1 INVX1_1006 ( .A(core__abc_22172_new_n4852_), .Y(core__abc_22172_new_n4853_));
INVX1 INVX1_1007 ( .A(core__abc_22172_new_n4855_), .Y(core__abc_22172_new_n4857_));
INVX1 INVX1_1008 ( .A(core_key_91_), .Y(core__abc_22172_new_n4861_));
INVX1 INVX1_1009 ( .A(core__abc_22172_new_n4863_), .Y(core__abc_22172_new_n4864_));
INVX1 INVX1_101 ( .A(_abc_19873_new_n2445_), .Y(_abc_19873_new_n2446_));
INVX1 INVX1_1010 ( .A(core__abc_22172_new_n4847_), .Y(core__abc_22172_new_n4875_));
INVX1 INVX1_1011 ( .A(core__abc_22172_new_n4887_), .Y(core__abc_22172_new_n4895_));
INVX1 INVX1_1012 ( .A(core__abc_22172_new_n4892_), .Y(core__abc_22172_new_n4897_));
INVX1 INVX1_1013 ( .A(core__abc_22172_new_n4900_), .Y(core__abc_22172_new_n4901_));
INVX1 INVX1_1014 ( .A(core_v3_reg_12_), .Y(core__abc_22172_new_n4902_));
INVX1 INVX1_1015 ( .A(core__abc_22172_new_n4904_), .Y(core__abc_22172_new_n4906_));
INVX1 INVX1_1016 ( .A(core__abc_22172_new_n4908_), .Y(core__abc_22172_new_n4909_));
INVX1 INVX1_1017 ( .A(core__abc_22172_new_n4912_), .Y(core__abc_22172_new_n4913_));
INVX1 INVX1_1018 ( .A(core__abc_22172_new_n4916_), .Y(core__abc_22172_new_n4917_));
INVX1 INVX1_1019 ( .A(core__abc_22172_new_n4918_), .Y(core__abc_22172_new_n4919_));
INVX1 INVX1_102 ( .A(_abc_19873_new_n2450_), .Y(_abc_19873_new_n2451_));
INVX1 INVX1_1020 ( .A(core__abc_22172_new_n4921_), .Y(core__abc_22172_new_n4922_));
INVX1 INVX1_1021 ( .A(core_key_92_), .Y(core__abc_22172_new_n4927_));
INVX1 INVX1_1022 ( .A(core__abc_22172_new_n4930_), .Y(core__abc_22172_new_n4931_));
INVX1 INVX1_1023 ( .A(core__abc_22172_new_n4914_), .Y(core__abc_22172_new_n4939_));
INVX1 INVX1_1024 ( .A(core__abc_22172_new_n4940_), .Y(core__abc_22172_new_n4941_));
INVX1 INVX1_1025 ( .A(core__abc_22172_new_n4942_), .Y(core__abc_22172_new_n4943_));
INVX1 INVX1_1026 ( .A(core__abc_22172_new_n4947_), .Y(core__abc_22172_new_n4948_));
INVX1 INVX1_1027 ( .A(core__abc_22172_new_n4952_), .Y(core__abc_22172_new_n4953_));
INVX1 INVX1_1028 ( .A(core__abc_22172_new_n4956_), .Y(core__abc_22172_new_n4957_));
INVX1 INVX1_1029 ( .A(core__abc_22172_new_n4946_), .Y(core__abc_22172_new_n4958_));
INVX1 INVX1_103 ( .A(_abc_19873_new_n2455_), .Y(_abc_19873_new_n2456_));
INVX1 INVX1_1030 ( .A(core__abc_22172_new_n4955_), .Y(core__abc_22172_new_n4959_));
INVX1 INVX1_1031 ( .A(core__abc_22172_new_n4960_), .Y(core__abc_22172_new_n4961_));
INVX1 INVX1_1032 ( .A(core__abc_22172_new_n4962_), .Y(core__abc_22172_new_n4963_));
INVX1 INVX1_1033 ( .A(core__abc_22172_new_n4966_), .Y(core__abc_22172_new_n4968_));
INVX1 INVX1_1034 ( .A(core_key_93_), .Y(core__abc_22172_new_n4972_));
INVX1 INVX1_1035 ( .A(core__abc_22172_new_n4974_), .Y(core__abc_22172_new_n4975_));
INVX1 INVX1_1036 ( .A(core__abc_22172_new_n4985_), .Y(core__abc_22172_new_n4991_));
INVX1 INVX1_1037 ( .A(core__abc_22172_new_n4988_), .Y(core__abc_22172_new_n4993_));
INVX1 INVX1_1038 ( .A(core_v3_reg_14_), .Y(core__abc_22172_new_n4997_));
INVX1 INVX1_1039 ( .A(core__abc_22172_new_n4999_), .Y(core__abc_22172_new_n5001_));
INVX1 INVX1_104 ( .A(_abc_19873_new_n2460_), .Y(_abc_19873_new_n2461_));
INVX1 INVX1_1040 ( .A(core__abc_22172_new_n5003_), .Y(core__abc_22172_new_n5004_));
INVX1 INVX1_1041 ( .A(core__abc_22172_new_n4996_), .Y(core__abc_22172_new_n5009_));
INVX1 INVX1_1042 ( .A(core__abc_22172_new_n5007_), .Y(core__abc_22172_new_n5010_));
INVX1 INVX1_1043 ( .A(core__abc_22172_new_n5012_), .Y(core__abc_22172_new_n5013_));
INVX1 INVX1_1044 ( .A(core__abc_22172_new_n5016_), .Y(core__abc_22172_new_n5017_));
INVX1 INVX1_1045 ( .A(core__abc_22172_new_n5020_), .Y(core__abc_22172_new_n5022_));
INVX1 INVX1_1046 ( .A(core_key_94_), .Y(core__abc_22172_new_n5026_));
INVX1 INVX1_1047 ( .A(core__abc_22172_new_n5028_), .Y(core__abc_22172_new_n5029_));
INVX1 INVX1_1048 ( .A(core__abc_22172_new_n5046_), .Y(core__abc_22172_new_n5047_));
INVX1 INVX1_1049 ( .A(core_v3_reg_15_), .Y(core__abc_22172_new_n5052_));
INVX1 INVX1_105 ( .A(_abc_19873_new_n2465_), .Y(_abc_19873_new_n2466_));
INVX1 INVX1_1050 ( .A(core__abc_22172_new_n5050_), .Y(core__abc_22172_new_n5053_));
INVX1 INVX1_1051 ( .A(core__abc_22172_new_n5051_), .Y(core__abc_22172_new_n5060_));
INVX1 INVX1_1052 ( .A(core__abc_22172_new_n5065_), .Y(core__abc_22172_new_n5066_));
INVX1 INVX1_1053 ( .A(core__abc_22172_new_n5068_), .Y(core__abc_22172_new_n5070_));
INVX1 INVX1_1054 ( .A(core__abc_22172_new_n5075_), .Y(core__abc_22172_new_n5076_));
INVX1 INVX1_1055 ( .A(core__abc_22172_new_n5014_), .Y(core__abc_22172_new_n5095_));
INVX1 INVX1_1056 ( .A(core_v3_reg_16_), .Y(core__abc_22172_new_n5105_));
INVX1 INVX1_1057 ( .A(core__abc_22172_new_n3153_), .Y(core__abc_22172_new_n5106_));
INVX1 INVX1_1058 ( .A(core__abc_22172_new_n5109_), .Y(core__abc_22172_new_n5110_));
INVX1 INVX1_1059 ( .A(core__abc_22172_new_n5113_), .Y(core__abc_22172_new_n5114_));
INVX1 INVX1_106 ( .A(_abc_19873_new_n2470_), .Y(_abc_19873_new_n2471_));
INVX1 INVX1_1060 ( .A(core__abc_22172_new_n5117_), .Y(core__abc_22172_new_n5118_));
INVX1 INVX1_1061 ( .A(core__abc_22172_new_n5092_), .Y(core__abc_22172_new_n5120_));
INVX1 INVX1_1062 ( .A(core__abc_22172_new_n5093_), .Y(core__abc_22172_new_n5121_));
INVX1 INVX1_1063 ( .A(core__abc_22172_new_n4782_), .Y(core__abc_22172_new_n5122_));
INVX1 INVX1_1064 ( .A(core__abc_22172_new_n4881_), .Y(core__abc_22172_new_n5125_));
INVX1 INVX1_1065 ( .A(core__abc_22172_new_n5087_), .Y(core__abc_22172_new_n5127_));
INVX1 INVX1_1066 ( .A(core__abc_22172_new_n5100_), .Y(core__abc_22172_new_n5135_));
INVX1 INVX1_1067 ( .A(core__abc_22172_new_n5141_), .Y(core__abc_22172_new_n5143_));
INVX1 INVX1_1068 ( .A(core__abc_22172_new_n5149_), .Y(core__abc_22172_new_n5150_));
INVX1 INVX1_1069 ( .A(core__abc_22172_new_n5159_), .Y(core__abc_22172_new_n5160_));
INVX1 INVX1_107 ( .A(_abc_19873_new_n2476_), .Y(_abc_19873_new_n2477_));
INVX1 INVX1_1070 ( .A(core__abc_22172_new_n5162_), .Y(core__abc_22172_new_n5163_));
INVX1 INVX1_1071 ( .A(core__abc_22172_new_n5164_), .Y(core__abc_22172_new_n5165_));
INVX1 INVX1_1072 ( .A(core__abc_22172_new_n5169_), .Y(core__abc_22172_new_n5170_));
INVX1 INVX1_1073 ( .A(core__abc_22172_new_n5172_), .Y(core__abc_22172_new_n5173_));
INVX1 INVX1_1074 ( .A(core__abc_22172_new_n5174_), .Y(core__abc_22172_new_n5175_));
INVX1 INVX1_1075 ( .A(core__abc_22172_new_n5176_), .Y(core__abc_22172_new_n5177_));
INVX1 INVX1_1076 ( .A(core__abc_22172_new_n5178_), .Y(core__abc_22172_new_n5179_));
INVX1 INVX1_1077 ( .A(core__abc_22172_new_n5182_), .Y(core__abc_22172_new_n5183_));
INVX1 INVX1_1078 ( .A(core_key_97_), .Y(core__abc_22172_new_n5188_));
INVX1 INVX1_1079 ( .A(core__abc_22172_new_n5191_), .Y(core__abc_22172_new_n5192_));
INVX1 INVX1_108 ( .A(_abc_19873_new_n2481_), .Y(_abc_19873_new_n2482_));
INVX1 INVX1_1080 ( .A(core__abc_22172_new_n5208_), .Y(core__abc_22172_new_n5209_));
INVX1 INVX1_1081 ( .A(core_v3_reg_18_), .Y(core__abc_22172_new_n5210_));
INVX1 INVX1_1082 ( .A(core__abc_22172_new_n3157_), .Y(core__abc_22172_new_n5211_));
INVX1 INVX1_1083 ( .A(core__abc_22172_new_n5213_), .Y(core__abc_22172_new_n5214_));
INVX1 INVX1_1084 ( .A(core__abc_22172_new_n5217_), .Y(core__abc_22172_new_n5218_));
INVX1 INVX1_1085 ( .A(core__abc_22172_new_n5221_), .Y(core__abc_22172_new_n5222_));
INVX1 INVX1_1086 ( .A(core__abc_22172_new_n5225_), .Y(core__abc_22172_new_n5226_));
INVX1 INVX1_1087 ( .A(core__abc_22172_new_n5227_), .Y(core__abc_22172_new_n5228_));
INVX1 INVX1_1088 ( .A(core__abc_22172_new_n5230_), .Y(core__abc_22172_new_n5231_));
INVX1 INVX1_1089 ( .A(core__abc_22172_new_n5238_), .Y(core__abc_22172_new_n5239_));
INVX1 INVX1_109 ( .A(_abc_19873_new_n2486_), .Y(_abc_19873_new_n2487_));
INVX1 INVX1_1090 ( .A(core__abc_22172_new_n4089_), .Y(core__abc_22172_new_n5247_));
INVX1 INVX1_1091 ( .A(core__abc_22172_new_n5223_), .Y(core__abc_22172_new_n5248_));
INVX1 INVX1_1092 ( .A(core__abc_22172_new_n5250_), .Y(core__abc_22172_new_n5251_));
INVX1 INVX1_1093 ( .A(core__abc_22172_new_n5257_), .Y(core__abc_22172_new_n5258_));
INVX1 INVX1_1094 ( .A(core__abc_22172_new_n5259_), .Y(core__abc_22172_new_n5260_));
INVX1 INVX1_1095 ( .A(core__abc_22172_new_n5261_), .Y(core__abc_22172_new_n5262_));
INVX1 INVX1_1096 ( .A(core__abc_22172_new_n5265_), .Y(core__abc_22172_new_n5266_));
INVX1 INVX1_1097 ( .A(core__abc_22172_new_n5249_), .Y(core__abc_22172_new_n5270_));
INVX1 INVX1_1098 ( .A(core__abc_22172_new_n5267_), .Y(core__abc_22172_new_n5271_));
INVX1 INVX1_1099 ( .A(core__abc_22172_new_n5274_), .Y(core__abc_22172_new_n5276_));
INVX1 INVX1_11 ( .A(\write_data[0] ), .Y(_abc_19873_new_n2122_));
INVX1 INVX1_110 ( .A(_abc_19873_new_n2491_), .Y(_abc_19873_new_n2492_));
INVX1 INVX1_1100 ( .A(core__abc_22172_new_n5281_), .Y(core__abc_22172_new_n5282_));
INVX1 INVX1_1101 ( .A(core__abc_22172_new_n5296_), .Y(core__abc_22172_new_n5297_));
INVX1 INVX1_1102 ( .A(core__abc_22172_new_n5304_), .Y(core__abc_22172_new_n5305_));
INVX1 INVX1_1103 ( .A(core_v3_reg_20_), .Y(core__abc_22172_new_n5306_));
INVX1 INVX1_1104 ( .A(core__abc_22172_new_n5308_), .Y(core__abc_22172_new_n5310_));
INVX1 INVX1_1105 ( .A(core__abc_22172_new_n5312_), .Y(core__abc_22172_new_n5313_));
INVX1 INVX1_1106 ( .A(core__abc_22172_new_n5316_), .Y(core__abc_22172_new_n5317_));
INVX1 INVX1_1107 ( .A(core__abc_22172_new_n5320_), .Y(core__abc_22172_new_n5321_));
INVX1 INVX1_1108 ( .A(core__abc_22172_new_n5322_), .Y(core__abc_22172_new_n5323_));
INVX1 INVX1_1109 ( .A(core__abc_22172_new_n5325_), .Y(core__abc_22172_new_n5327_));
INVX1 INVX1_111 ( .A(_abc_19873_new_n2496_), .Y(_abc_19873_new_n2497_));
INVX1 INVX1_1110 ( .A(core__abc_22172_new_n5333_), .Y(core__abc_22172_new_n5334_));
INVX1 INVX1_1111 ( .A(core__abc_22172_new_n5318_), .Y(core__abc_22172_new_n5343_));
INVX1 INVX1_1112 ( .A(core__abc_22172_new_n5344_), .Y(core__abc_22172_new_n5345_));
INVX1 INVX1_1113 ( .A(core__abc_22172_new_n5349_), .Y(core__abc_22172_new_n5350_));
INVX1 INVX1_1114 ( .A(core__abc_22172_new_n5354_), .Y(core__abc_22172_new_n5355_));
INVX1 INVX1_1115 ( .A(core__abc_22172_new_n5359_), .Y(core__abc_22172_new_n5360_));
INVX1 INVX1_1116 ( .A(core__abc_22172_new_n5363_), .Y(core__abc_22172_new_n5364_));
INVX1 INVX1_1117 ( .A(core__abc_22172_new_n5361_), .Y(core__abc_22172_new_n5365_));
INVX1 INVX1_1118 ( .A(core__abc_22172_new_n5366_), .Y(core__abc_22172_new_n5367_));
INVX1 INVX1_1119 ( .A(core__abc_22172_new_n5369_), .Y(core__abc_22172_new_n5370_));
INVX1 INVX1_112 ( .A(_abc_19873_new_n2501_), .Y(_abc_19873_new_n2502_));
INVX1 INVX1_1120 ( .A(core__abc_22172_new_n5372_), .Y(core__abc_22172_new_n5374_));
INVX1 INVX1_1121 ( .A(core_key_101_), .Y(core__abc_22172_new_n5378_));
INVX1 INVX1_1122 ( .A(core__abc_22172_new_n5381_), .Y(core__abc_22172_new_n5382_));
INVX1 INVX1_1123 ( .A(core__abc_22172_new_n5391_), .Y(core__abc_22172_new_n5392_));
INVX1 INVX1_1124 ( .A(core__abc_22172_new_n5393_), .Y(core__abc_22172_new_n5394_));
INVX1 INVX1_1125 ( .A(core__abc_22172_new_n5397_), .Y(core__abc_22172_new_n5398_));
INVX1 INVX1_1126 ( .A(core__abc_22172_new_n5400_), .Y(core__abc_22172_new_n5401_));
INVX1 INVX1_1127 ( .A(core__abc_22172_new_n5403_), .Y(core__abc_22172_new_n5404_));
INVX1 INVX1_1128 ( .A(core__abc_22172_new_n5407_), .Y(core__abc_22172_new_n5408_));
INVX1 INVX1_1129 ( .A(core_v3_reg_22_), .Y(core__abc_22172_new_n5410_));
INVX1 INVX1_113 ( .A(_abc_19873_new_n2506_), .Y(_abc_19873_new_n2507_));
INVX1 INVX1_1130 ( .A(core__abc_22172_new_n5412_), .Y(core__abc_22172_new_n5413_));
INVX1 INVX1_1131 ( .A(core__abc_22172_new_n5416_), .Y(core__abc_22172_new_n5417_));
INVX1 INVX1_1132 ( .A(core__abc_22172_new_n4291_), .Y(core__abc_22172_new_n5422_));
INVX1 INVX1_1133 ( .A(core__abc_22172_new_n5420_), .Y(core__abc_22172_new_n5423_));
INVX1 INVX1_1134 ( .A(core_key_102_), .Y(core__abc_22172_new_n5427_));
INVX1 INVX1_1135 ( .A(core__abc_22172_new_n5430_), .Y(core__abc_22172_new_n5431_));
INVX1 INVX1_1136 ( .A(core__abc_22172_new_n5441_), .Y(core__abc_22172_new_n5442_));
INVX1 INVX1_1137 ( .A(core__abc_22172_new_n5445_), .Y(core__abc_22172_new_n5446_));
INVX1 INVX1_1138 ( .A(core__abc_22172_new_n5450_), .Y(core__abc_22172_new_n5451_));
INVX1 INVX1_1139 ( .A(core__abc_22172_new_n5453_), .Y(core__abc_22172_new_n5454_));
INVX1 INVX1_114 ( .A(_abc_19873_new_n2511_), .Y(_abc_19873_new_n2512_));
INVX1 INVX1_1140 ( .A(core__abc_22172_new_n5455_), .Y(core__abc_22172_new_n5456_));
INVX1 INVX1_1141 ( .A(core__abc_22172_new_n5439_), .Y(core__abc_22172_new_n5460_));
INVX1 INVX1_1142 ( .A(core__abc_22172_new_n5457_), .Y(core__abc_22172_new_n5461_));
INVX1 INVX1_1143 ( .A(core__abc_22172_new_n5464_), .Y(core__abc_22172_new_n5465_));
INVX1 INVX1_1144 ( .A(core__abc_22172_new_n5471_), .Y(core__abc_22172_new_n5472_));
INVX1 INVX1_1145 ( .A(core__abc_22172_new_n5496_), .Y(core__abc_22172_new_n5497_));
INVX1 INVX1_1146 ( .A(core_v3_reg_24_), .Y(core__abc_22172_new_n5498_));
INVX1 INVX1_1147 ( .A(core__abc_22172_new_n3180_), .Y(core__abc_22172_new_n5500_));
INVX1 INVX1_1148 ( .A(core__abc_22172_new_n5502_), .Y(core__abc_22172_new_n5503_));
INVX1 INVX1_1149 ( .A(core__abc_22172_new_n5506_), .Y(core__abc_22172_new_n5507_));
INVX1 INVX1_115 ( .A(_abc_19873_new_n2516_), .Y(_abc_19873_new_n2517_));
INVX1 INVX1_1150 ( .A(core__abc_22172_new_n5510_), .Y(core__abc_22172_new_n5511_));
INVX1 INVX1_1151 ( .A(core__abc_22172_new_n5490_), .Y(core__abc_22172_new_n5513_));
INVX1 INVX1_1152 ( .A(core__abc_22172_new_n5491_), .Y(core__abc_22172_new_n5514_));
INVX1 INVX1_1153 ( .A(core__abc_22172_new_n4412_), .Y(core__abc_22172_new_n5520_));
INVX1 INVX1_1154 ( .A(core__abc_22172_new_n5518_), .Y(core__abc_22172_new_n5521_));
INVX1 INVX1_1155 ( .A(core__abc_22172_new_n5527_), .Y(core__abc_22172_new_n5528_));
INVX1 INVX1_1156 ( .A(core__abc_22172_new_n5508_), .Y(core__abc_22172_new_n5537_));
INVX1 INVX1_1157 ( .A(core__abc_22172_new_n5512_), .Y(core__abc_22172_new_n5538_));
INVX1 INVX1_1158 ( .A(core__abc_22172_new_n5539_), .Y(core__abc_22172_new_n5540_));
INVX1 INVX1_1159 ( .A(core__abc_22172_new_n5541_), .Y(core__abc_22172_new_n5542_));
INVX1 INVX1_116 ( .A(_abc_19873_new_n2521_), .Y(_abc_19873_new_n2522_));
INVX1 INVX1_1160 ( .A(core__abc_22172_new_n5545_), .Y(core__abc_22172_new_n5546_));
INVX1 INVX1_1161 ( .A(core_v3_reg_25_), .Y(core__abc_22172_new_n5547_));
INVX1 INVX1_1162 ( .A(core__abc_22172_new_n5548_), .Y(core__abc_22172_new_n5549_));
INVX1 INVX1_1163 ( .A(core__abc_22172_new_n5552_), .Y(core__abc_22172_new_n5554_));
INVX1 INVX1_1164 ( .A(core__abc_22172_new_n5556_), .Y(core__abc_22172_new_n5557_));
INVX1 INVX1_1165 ( .A(core__abc_22172_new_n5558_), .Y(core__abc_22172_new_n5559_));
INVX1 INVX1_1166 ( .A(core__abc_22172_new_n5560_), .Y(core__abc_22172_new_n5561_));
INVX1 INVX1_1167 ( .A(core__abc_22172_new_n5562_), .Y(core__abc_22172_new_n5564_));
INVX1 INVX1_1168 ( .A(core__abc_22172_new_n5566_), .Y(core__abc_22172_new_n5567_));
INVX1 INVX1_1169 ( .A(core__abc_22172_new_n5574_), .Y(core__abc_22172_new_n5575_));
INVX1 INVX1_117 ( .A(_abc_19873_new_n2526_), .Y(_abc_19873_new_n2527_));
INVX1 INVX1_1170 ( .A(core__abc_22172_new_n5585_), .Y(core__abc_22172_new_n5587_));
INVX1 INVX1_1171 ( .A(core__abc_22172_new_n5589_), .Y(core__abc_22172_new_n5590_));
INVX1 INVX1_1172 ( .A(core_v3_reg_26_), .Y(core__abc_22172_new_n5591_));
INVX1 INVX1_1173 ( .A(core__abc_22172_new_n3183_), .Y(core__abc_22172_new_n5592_));
INVX1 INVX1_1174 ( .A(core__abc_22172_new_n5594_), .Y(core__abc_22172_new_n5595_));
INVX1 INVX1_1175 ( .A(core__abc_22172_new_n5598_), .Y(core__abc_22172_new_n5599_));
INVX1 INVX1_1176 ( .A(core__abc_22172_new_n5603_), .Y(core__abc_22172_new_n5604_));
INVX1 INVX1_1177 ( .A(core__abc_22172_new_n5608_), .Y(core__abc_22172_new_n5609_));
INVX1 INVX1_1178 ( .A(core__abc_22172_new_n5610_), .Y(core__abc_22172_new_n5612_));
INVX1 INVX1_1179 ( .A(core_key_106_), .Y(core__abc_22172_new_n5616_));
INVX1 INVX1_118 ( .A(_abc_19873_new_n2531_), .Y(_abc_19873_new_n2532_));
INVX1 INVX1_1180 ( .A(core__abc_22172_new_n5619_), .Y(core__abc_22172_new_n5620_));
INVX1 INVX1_1181 ( .A(core__abc_22172_new_n5600_), .Y(core__abc_22172_new_n5628_));
INVX1 INVX1_1182 ( .A(core__abc_22172_new_n5632_), .Y(core__abc_22172_new_n5633_));
INVX1 INVX1_1183 ( .A(core__abc_22172_new_n5634_), .Y(core__abc_22172_new_n5636_));
INVX1 INVX1_1184 ( .A(core__abc_22172_new_n5629_), .Y(core__abc_22172_new_n5640_));
INVX1 INVX1_1185 ( .A(core__abc_22172_new_n5638_), .Y(core__abc_22172_new_n5641_));
INVX1 INVX1_1186 ( .A(core__abc_22172_new_n5643_), .Y(core__abc_22172_new_n5644_));
INVX1 INVX1_1187 ( .A(core__abc_22172_new_n5650_), .Y(core__abc_22172_new_n5651_));
INVX1 INVX1_1188 ( .A(core__abc_22172_new_n5602_), .Y(core__abc_22172_new_n5663_));
INVX1 INVX1_1189 ( .A(core__abc_22172_new_n5635_), .Y(core__abc_22172_new_n5666_));
INVX1 INVX1_119 ( .A(_abc_19873_new_n2536_), .Y(_abc_19873_new_n2537_));
INVX1 INVX1_1190 ( .A(core__abc_22172_new_n5668_), .Y(core__abc_22172_new_n5669_));
INVX1 INVX1_1191 ( .A(core__abc_22172_new_n5676_), .Y(core__abc_22172_new_n5678_));
INVX1 INVX1_1192 ( .A(core__abc_22172_new_n5680_), .Y(core__abc_22172_new_n5681_));
INVX1 INVX1_1193 ( .A(core__abc_22172_new_n5684_), .Y(core__abc_22172_new_n5685_));
INVX1 INVX1_1194 ( .A(core__abc_22172_new_n5665_), .Y(core__abc_22172_new_n5687_));
INVX1 INVX1_1195 ( .A(core__abc_22172_new_n5672_), .Y(core__abc_22172_new_n5689_));
INVX1 INVX1_1196 ( .A(core__abc_22172_new_n5693_), .Y(core__abc_22172_new_n5695_));
INVX1 INVX1_1197 ( .A(core__abc_22172_new_n5701_), .Y(core__abc_22172_new_n5702_));
INVX1 INVX1_1198 ( .A(core__abc_22172_new_n5712_), .Y(core__abc_22172_new_n5713_));
INVX1 INVX1_1199 ( .A(core__abc_22172_new_n5716_), .Y(core__abc_22172_new_n5717_));
INVX1 INVX1_12 ( .A(_abc_19873_new_n2123_), .Y(_abc_19873_new_n2124_));
INVX1 INVX1_120 ( .A(_abc_19873_new_n2541_), .Y(_abc_19873_new_n2542_));
INVX1 INVX1_1200 ( .A(core__abc_22172_new_n5720_), .Y(core__abc_22172_new_n5721_));
INVX1 INVX1_1201 ( .A(core__abc_22172_new_n5711_), .Y(core__abc_22172_new_n5723_));
INVX1 INVX1_1202 ( .A(core__abc_22172_new_n5725_), .Y(core__abc_22172_new_n5727_));
INVX1 INVX1_1203 ( .A(core_key_109_), .Y(core__abc_22172_new_n5731_));
INVX1 INVX1_1204 ( .A(core__abc_22172_new_n5734_), .Y(core__abc_22172_new_n5735_));
INVX1 INVX1_1205 ( .A(core__abc_22172_new_n5719_), .Y(core__abc_22172_new_n5746_));
INVX1 INVX1_1206 ( .A(core__abc_22172_new_n5752_), .Y(core__abc_22172_new_n5753_));
INVX1 INVX1_1207 ( .A(core__abc_22172_new_n5755_), .Y(core__abc_22172_new_n5756_));
INVX1 INVX1_1208 ( .A(core__abc_22172_new_n5759_), .Y(core__abc_22172_new_n5760_));
INVX1 INVX1_1209 ( .A(core__abc_22172_new_n5744_), .Y(core__abc_22172_new_n5762_));
INVX1 INVX1_121 ( .A(_abc_19873_new_n2546_), .Y(_abc_19873_new_n2547_));
INVX1 INVX1_1210 ( .A(core__abc_22172_new_n5748_), .Y(core__abc_22172_new_n5764_));
INVX1 INVX1_1211 ( .A(core__abc_22172_new_n5767_), .Y(core__abc_22172_new_n5769_));
INVX1 INVX1_1212 ( .A(core_key_110_), .Y(core__abc_22172_new_n5773_));
INVX1 INVX1_1213 ( .A(core__abc_22172_new_n5776_), .Y(core__abc_22172_new_n5777_));
INVX1 INVX1_1214 ( .A(core__abc_22172_new_n5789_), .Y(core__abc_22172_new_n5790_));
INVX1 INVX1_1215 ( .A(core__abc_22172_new_n5791_), .Y(core__abc_22172_new_n5793_));
INVX1 INVX1_1216 ( .A(core__abc_22172_new_n5758_), .Y(core__abc_22172_new_n5797_));
INVX1 INVX1_1217 ( .A(core__abc_22172_new_n5814_), .Y(core__abc_22172_new_n5815_));
INVX1 INVX1_1218 ( .A(core__abc_22172_new_n5840_), .Y(core__abc_22172_new_n5841_));
INVX1 INVX1_1219 ( .A(core__abc_22172_new_n5844_), .Y(core__abc_22172_new_n5845_));
INVX1 INVX1_122 ( .A(_abc_19873_new_n2551_), .Y(_abc_19873_new_n2552_));
INVX1 INVX1_1220 ( .A(core__abc_22172_new_n5827_), .Y(core__abc_22172_new_n5847_));
INVX1 INVX1_1221 ( .A(core__abc_22172_new_n5829_), .Y(core__abc_22172_new_n5849_));
INVX1 INVX1_1222 ( .A(core__abc_22172_new_n5830_), .Y(core__abc_22172_new_n5850_));
INVX1 INVX1_1223 ( .A(core__abc_22172_new_n5834_), .Y(core__abc_22172_new_n5851_));
INVX1 INVX1_1224 ( .A(core__abc_22172_new_n5856_), .Y(core__abc_22172_new_n5858_));
INVX1 INVX1_1225 ( .A(core_key_112_), .Y(core__abc_22172_new_n5862_));
INVX1 INVX1_1226 ( .A(core__abc_22172_new_n5865_), .Y(core__abc_22172_new_n5866_));
INVX1 INVX1_1227 ( .A(core__abc_22172_new_n5846_), .Y(core__abc_22172_new_n5875_));
INVX1 INVX1_1228 ( .A(core__abc_22172_new_n5842_), .Y(core__abc_22172_new_n5876_));
INVX1 INVX1_1229 ( .A(core__abc_22172_new_n5877_), .Y(core__abc_22172_new_n5878_));
INVX1 INVX1_123 ( .A(_abc_19873_new_n2556_), .Y(_abc_19873_new_n2557_));
INVX1 INVX1_1230 ( .A(core__abc_22172_new_n5882_), .Y(core__abc_22172_new_n5883_));
INVX1 INVX1_1231 ( .A(core__abc_22172_new_n5887_), .Y(core__abc_22172_new_n5888_));
INVX1 INVX1_1232 ( .A(core__abc_22172_new_n5885_), .Y(core__abc_22172_new_n5889_));
INVX1 INVX1_1233 ( .A(core__abc_22172_new_n5890_), .Y(core__abc_22172_new_n5891_));
INVX1 INVX1_1234 ( .A(core__abc_22172_new_n5892_), .Y(core__abc_22172_new_n5893_));
INVX1 INVX1_1235 ( .A(core__abc_22172_new_n5896_), .Y(core__abc_22172_new_n5897_));
INVX1 INVX1_1236 ( .A(core__abc_22172_new_n5904_), .Y(core__abc_22172_new_n5905_));
INVX1 INVX1_1237 ( .A(core__abc_22172_new_n5918_), .Y(core__abc_22172_new_n5919_));
INVX1 INVX1_1238 ( .A(core__abc_22172_new_n5921_), .Y(core__abc_22172_new_n5923_));
INVX1 INVX1_1239 ( .A(core__abc_22172_new_n5926_), .Y(core__abc_22172_new_n5927_));
INVX1 INVX1_124 ( .A(_abc_19873_new_n2561_), .Y(_abc_19873_new_n2562_));
INVX1 INVX1_1240 ( .A(core__abc_22172_new_n5929_), .Y(core__abc_22172_new_n5931_));
INVX1 INVX1_1241 ( .A(core_key_114_), .Y(core__abc_22172_new_n5935_));
INVX1 INVX1_1242 ( .A(core__abc_22172_new_n5938_), .Y(core__abc_22172_new_n5939_));
INVX1 INVX1_1243 ( .A(core__abc_22172_new_n5922_), .Y(core__abc_22172_new_n5948_));
INVX1 INVX1_1244 ( .A(core__abc_22172_new_n5952_), .Y(core__abc_22172_new_n5953_));
INVX1 INVX1_1245 ( .A(core__abc_22172_new_n5954_), .Y(core__abc_22172_new_n5955_));
INVX1 INVX1_1246 ( .A(core__abc_22172_new_n5957_), .Y(core__abc_22172_new_n5958_));
INVX1 INVX1_1247 ( .A(core__abc_22172_new_n5959_), .Y(core__abc_22172_new_n5960_));
INVX1 INVX1_1248 ( .A(core__abc_22172_new_n5961_), .Y(core__abc_22172_new_n5962_));
INVX1 INVX1_1249 ( .A(core__abc_22172_new_n5964_), .Y(core__abc_22172_new_n5966_));
INVX1 INVX1_125 ( .A(_abc_19873_new_n2566_), .Y(_abc_19873_new_n2567_));
INVX1 INVX1_1250 ( .A(core__abc_22172_new_n5972_), .Y(core__abc_22172_new_n5973_));
INVX1 INVX1_1251 ( .A(core__abc_22172_new_n5914_), .Y(core__abc_22172_new_n5982_));
INVX1 INVX1_1252 ( .A(core__abc_22172_new_n5925_), .Y(core__abc_22172_new_n5983_));
INVX1 INVX1_1253 ( .A(core__abc_22172_new_n5987_), .Y(core__abc_22172_new_n5988_));
INVX1 INVX1_1254 ( .A(core__abc_22172_new_n5994_), .Y(core__abc_22172_new_n5996_));
INVX1 INVX1_1255 ( .A(core__abc_22172_new_n5998_), .Y(core__abc_22172_new_n5999_));
INVX1 INVX1_1256 ( .A(core__abc_22172_new_n6002_), .Y(core__abc_22172_new_n6003_));
INVX1 INVX1_1257 ( .A(core__abc_22172_new_n5989_), .Y(core__abc_22172_new_n6005_));
INVX1 INVX1_1258 ( .A(core__abc_22172_new_n5990_), .Y(core__abc_22172_new_n6006_));
INVX1 INVX1_1259 ( .A(core__abc_22172_new_n6010_), .Y(core__abc_22172_new_n6012_));
INVX1 INVX1_126 ( .A(_abc_19873_new_n2571_), .Y(_abc_19873_new_n2572_));
INVX1 INVX1_1260 ( .A(core__abc_22172_new_n6018_), .Y(core__abc_22172_new_n6019_));
INVX1 INVX1_1261 ( .A(core__abc_22172_new_n6029_), .Y(core__abc_22172_new_n6030_));
INVX1 INVX1_1262 ( .A(core__abc_22172_new_n6033_), .Y(core__abc_22172_new_n6034_));
INVX1 INVX1_1263 ( .A(core__abc_22172_new_n6037_), .Y(core__abc_22172_new_n6038_));
INVX1 INVX1_1264 ( .A(core__abc_22172_new_n6028_), .Y(core__abc_22172_new_n6040_));
INVX1 INVX1_1265 ( .A(core__abc_22172_new_n6042_), .Y(core__abc_22172_new_n6043_));
INVX1 INVX1_1266 ( .A(core_key_117_), .Y(core__abc_22172_new_n6048_));
INVX1 INVX1_1267 ( .A(core__abc_22172_new_n6051_), .Y(core__abc_22172_new_n6052_));
INVX1 INVX1_1268 ( .A(core__abc_22172_new_n6036_), .Y(core__abc_22172_new_n6063_));
INVX1 INVX1_1269 ( .A(core__abc_22172_new_n6068_), .Y(core__abc_22172_new_n6070_));
INVX1 INVX1_127 ( .A(_abc_19873_new_n2576_), .Y(_abc_19873_new_n2577_));
INVX1 INVX1_1270 ( .A(core__abc_22172_new_n6072_), .Y(core__abc_22172_new_n6073_));
INVX1 INVX1_1271 ( .A(core__abc_22172_new_n6076_), .Y(core__abc_22172_new_n6077_));
INVX1 INVX1_1272 ( .A(core__abc_22172_new_n6061_), .Y(core__abc_22172_new_n6079_));
INVX1 INVX1_1273 ( .A(core__abc_22172_new_n6065_), .Y(core__abc_22172_new_n6081_));
INVX1 INVX1_1274 ( .A(core__abc_22172_new_n6084_), .Y(core__abc_22172_new_n6086_));
INVX1 INVX1_1275 ( .A(core_key_118_), .Y(core__abc_22172_new_n6090_));
INVX1 INVX1_1276 ( .A(core__abc_22172_new_n6093_), .Y(core__abc_22172_new_n6094_));
INVX1 INVX1_1277 ( .A(core__abc_22172_new_n6104_), .Y(core__abc_22172_new_n6105_));
INVX1 INVX1_1278 ( .A(core__abc_22172_new_n6108_), .Y(core__abc_22172_new_n6109_));
INVX1 INVX1_1279 ( .A(core__abc_22172_new_n6074_), .Y(core__abc_22172_new_n6114_));
INVX1 INVX1_128 ( .A(_abc_19873_new_n2581_), .Y(_abc_19873_new_n2582_));
INVX1 INVX1_1280 ( .A(core__abc_22172_new_n6111_), .Y(core__abc_22172_new_n6118_));
INVX1 INVX1_1281 ( .A(core__abc_22172_new_n6131_), .Y(core__abc_22172_new_n6132_));
INVX1 INVX1_1282 ( .A(core__abc_22172_new_n5264_), .Y(core__abc_22172_new_n6141_));
INVX1 INVX1_1283 ( .A(core__abc_22172_new_n6149_), .Y(core__abc_22172_new_n6150_));
INVX1 INVX1_1284 ( .A(core__abc_22172_new_n6155_), .Y(core__abc_22172_new_n6157_));
INVX1 INVX1_1285 ( .A(core__abc_22172_new_n6159_), .Y(core__abc_22172_new_n6160_));
INVX1 INVX1_1286 ( .A(core__abc_22172_new_n6163_), .Y(core__abc_22172_new_n6164_));
INVX1 INVX1_1287 ( .A(core__abc_22172_new_n6176_), .Y(core__abc_22172_new_n6178_));
INVX1 INVX1_1288 ( .A(core__abc_22172_new_n6184_), .Y(core__abc_22172_new_n6185_));
INVX1 INVX1_1289 ( .A(core__abc_22172_new_n6195_), .Y(core__abc_22172_new_n6196_));
INVX1 INVX1_129 ( .A(_abc_19873_new_n2586_), .Y(_abc_19873_new_n2587_));
INVX1 INVX1_1290 ( .A(core__abc_22172_new_n6199_), .Y(core__abc_22172_new_n6200_));
INVX1 INVX1_1291 ( .A(core__abc_22172_new_n6203_), .Y(core__abc_22172_new_n6204_));
INVX1 INVX1_1292 ( .A(core__abc_22172_new_n6194_), .Y(core__abc_22172_new_n6206_));
INVX1 INVX1_1293 ( .A(core__abc_22172_new_n6208_), .Y(core__abc_22172_new_n6209_));
INVX1 INVX1_1294 ( .A(core__abc_22172_new_n6216_), .Y(core__abc_22172_new_n6217_));
INVX1 INVX1_1295 ( .A(core__abc_22172_new_n5357_), .Y(core__abc_22172_new_n6226_));
INVX1 INVX1_1296 ( .A(core__abc_22172_new_n6201_), .Y(core__abc_22172_new_n6227_));
INVX1 INVX1_1297 ( .A(core__abc_22172_new_n6161_), .Y(core__abc_22172_new_n6228_));
INVX1 INVX1_1298 ( .A(core__abc_22172_new_n6230_), .Y(core__abc_22172_new_n6231_));
INVX1 INVX1_1299 ( .A(core__abc_22172_new_n2964_), .Y(core__abc_22172_new_n6235_));
INVX1 INVX1_13 ( .A(\write_data[1] ), .Y(_abc_19873_new_n2128_));
INVX1 INVX1_130 ( .A(_abc_19873_new_n2591_), .Y(_abc_19873_new_n2592_));
INVX1 INVX1_1300 ( .A(core__abc_22172_new_n6238_), .Y(core__abc_22172_new_n6239_));
INVX1 INVX1_1301 ( .A(core__abc_22172_new_n6241_), .Y(core__abc_22172_new_n6242_));
INVX1 INVX1_1302 ( .A(core__abc_22172_new_n6245_), .Y(core__abc_22172_new_n6246_));
INVX1 INVX1_1303 ( .A(core__abc_22172_new_n6247_), .Y(core__abc_22172_new_n6248_));
INVX1 INVX1_1304 ( .A(core__abc_22172_new_n6250_), .Y(core__abc_22172_new_n6251_));
INVX1 INVX1_1305 ( .A(core_key_122_), .Y(core__abc_22172_new_n6256_));
INVX1 INVX1_1306 ( .A(core__abc_22172_new_n6259_), .Y(core__abc_22172_new_n6260_));
INVX1 INVX1_1307 ( .A(core__abc_22172_new_n6243_), .Y(core__abc_22172_new_n6268_));
INVX1 INVX1_1308 ( .A(core__abc_22172_new_n6269_), .Y(core__abc_22172_new_n6270_));
INVX1 INVX1_1309 ( .A(core__abc_22172_new_n6272_), .Y(core__abc_22172_new_n6273_));
INVX1 INVX1_131 ( .A(_abc_19873_new_n2596_), .Y(_abc_19873_new_n2597_));
INVX1 INVX1_1310 ( .A(core__abc_22172_new_n6275_), .Y(core__abc_22172_new_n6276_));
INVX1 INVX1_1311 ( .A(core__abc_22172_new_n6285_), .Y(core__abc_22172_new_n6286_));
INVX1 INVX1_1312 ( .A(core__abc_22172_new_n6292_), .Y(core__abc_22172_new_n6293_));
INVX1 INVX1_1313 ( .A(core__abc_22172_new_n6309_), .Y(core__abc_22172_new_n6310_));
INVX1 INVX1_1314 ( .A(core__abc_22172_new_n6314_), .Y(core__abc_22172_new_n6316_));
INVX1 INVX1_1315 ( .A(core__abc_22172_new_n6318_), .Y(core__abc_22172_new_n6319_));
INVX1 INVX1_1316 ( .A(core__abc_22172_new_n6322_), .Y(core__abc_22172_new_n6323_));
INVX1 INVX1_1317 ( .A(core__abc_22172_new_n6232_), .Y(core__abc_22172_new_n6325_));
INVX1 INVX1_1318 ( .A(core__abc_22172_new_n6307_), .Y(core__abc_22172_new_n6329_));
INVX1 INVX1_1319 ( .A(core__abc_22172_new_n6333_), .Y(core__abc_22172_new_n6335_));
INVX1 INVX1_132 ( .A(_abc_19873_new_n2601_), .Y(_abc_19873_new_n2602_));
INVX1 INVX1_1320 ( .A(core_key_124_), .Y(core__abc_22172_new_n6339_));
INVX1 INVX1_1321 ( .A(core__abc_22172_new_n6342_), .Y(core__abc_22172_new_n6343_));
INVX1 INVX1_1322 ( .A(core__abc_22172_new_n6353_), .Y(core__abc_22172_new_n6354_));
INVX1 INVX1_1323 ( .A(core__abc_22172_new_n6357_), .Y(core__abc_22172_new_n6358_));
INVX1 INVX1_1324 ( .A(core__abc_22172_new_n6320_), .Y(core__abc_22172_new_n6363_));
INVX1 INVX1_1325 ( .A(core__abc_22172_new_n6360_), .Y(core__abc_22172_new_n6367_));
INVX1 INVX1_1326 ( .A(core_key_125_), .Y(core__abc_22172_new_n6378_));
INVX1 INVX1_1327 ( .A(core__abc_22172_new_n6381_), .Y(core__abc_22172_new_n6382_));
INVX1 INVX1_1328 ( .A(core__abc_22172_new_n6394_), .Y(core__abc_22172_new_n6395_));
INVX1 INVX1_1329 ( .A(core__abc_22172_new_n6398_), .Y(core__abc_22172_new_n6400_));
INVX1 INVX1_133 ( .A(_abc_19873_new_n2606_), .Y(_abc_19873_new_n2607_));
INVX1 INVX1_1330 ( .A(core__abc_22172_new_n6402_), .Y(core__abc_22172_new_n6403_));
INVX1 INVX1_1331 ( .A(core__abc_22172_new_n6406_), .Y(core__abc_22172_new_n6411_));
INVX1 INVX1_1332 ( .A(core_key_126_), .Y(core__abc_22172_new_n6421_));
INVX1 INVX1_1333 ( .A(core__abc_22172_new_n6424_), .Y(core__abc_22172_new_n6425_));
INVX1 INVX1_1334 ( .A(core__abc_22172_new_n6434_), .Y(core__abc_22172_new_n6435_));
INVX1 INVX1_1335 ( .A(core__abc_22172_new_n6438_), .Y(core__abc_22172_new_n6439_));
INVX1 INVX1_1336 ( .A(core__abc_22172_new_n6404_), .Y(core__abc_22172_new_n6444_));
INVX1 INVX1_1337 ( .A(core__abc_22172_new_n6442_), .Y(core__abc_22172_new_n6446_));
INVX1 INVX1_1338 ( .A(core__abc_22172_new_n6457_), .Y(core__abc_22172_new_n6458_));
INVX1 INVX1_1339 ( .A(core_v1_reg_18_), .Y(core__abc_22172_new_n6468_));
INVX1 INVX1_134 ( .A(_abc_19873_new_n2611_), .Y(_abc_19873_new_n2612_));
INVX1 INVX1_1340 ( .A(core__abc_22172_new_n6473_), .Y(core__abc_22172_new_n6474_));
INVX1 INVX1_1341 ( .A(core_v1_reg_17_), .Y(core__abc_22172_new_n6476_));
INVX1 INVX1_1342 ( .A(core__abc_22172_new_n6479_), .Y(core__abc_22172_new_n6481_));
INVX1 INVX1_1343 ( .A(core__abc_22172_new_n4951_), .Y(core__abc_22172_new_n6485_));
INVX1 INVX1_1344 ( .A(core_v1_reg_16_), .Y(core__abc_22172_new_n6486_));
INVX1 INVX1_1345 ( .A(core__abc_22172_new_n6489_), .Y(core__abc_22172_new_n6490_));
INVX1 INVX1_1346 ( .A(core__abc_22172_new_n6491_), .Y(core__abc_22172_new_n6492_));
INVX1 INVX1_1347 ( .A(core__abc_22172_new_n6493_), .Y(core__abc_22172_new_n6494_));
INVX1 INVX1_1348 ( .A(core_v1_reg_15_), .Y(core__abc_22172_new_n6496_));
INVX1 INVX1_1349 ( .A(core__abc_22172_new_n6499_), .Y(core__abc_22172_new_n6500_));
INVX1 INVX1_135 ( .A(_abc_19873_new_n2616_), .Y(_abc_19873_new_n2617_));
INVX1 INVX1_1350 ( .A(core__abc_22172_new_n6503_), .Y(core__abc_22172_new_n6504_));
INVX1 INVX1_1351 ( .A(core__abc_22172_new_n6508_), .Y(core__abc_22172_new_n6509_));
INVX1 INVX1_1352 ( .A(core__abc_22172_new_n6510_), .Y(core__abc_22172_new_n6511_));
INVX1 INVX1_1353 ( .A(core__abc_22172_new_n4842_), .Y(core__abc_22172_new_n6513_));
INVX1 INVX1_1354 ( .A(core_v1_reg_13_), .Y(core__abc_22172_new_n6516_));
INVX1 INVX1_1355 ( .A(core__abc_22172_new_n6519_), .Y(core__abc_22172_new_n6520_));
INVX1 INVX1_1356 ( .A(core__abc_22172_new_n6523_), .Y(core__abc_22172_new_n6524_));
INVX1 INVX1_1357 ( .A(core__abc_22172_new_n4743_), .Y(core__abc_22172_new_n6526_));
INVX1 INVX1_1358 ( .A(core_v1_reg_12_), .Y(core__abc_22172_new_n6527_));
INVX1 INVX1_1359 ( .A(core__abc_22172_new_n6530_), .Y(core__abc_22172_new_n6531_));
INVX1 INVX1_136 ( .A(_abc_19873_new_n2621_), .Y(_abc_19873_new_n2622_));
INVX1 INVX1_1360 ( .A(core__abc_22172_new_n6532_), .Y(core__abc_22172_new_n6533_));
INVX1 INVX1_1361 ( .A(core_v1_reg_11_), .Y(core__abc_22172_new_n6534_));
INVX1 INVX1_1362 ( .A(core__abc_22172_new_n6537_), .Y(core__abc_22172_new_n6538_));
INVX1 INVX1_1363 ( .A(core__abc_22172_new_n6539_), .Y(core__abc_22172_new_n6540_));
INVX1 INVX1_1364 ( .A(core__abc_22172_new_n6543_), .Y(core__abc_22172_new_n6544_));
INVX1 INVX1_1365 ( .A(core__abc_22172_new_n6514_), .Y(core__abc_22172_new_n6546_));
INVX1 INVX1_1366 ( .A(core__abc_22172_new_n6521_), .Y(core__abc_22172_new_n6547_));
INVX1 INVX1_1367 ( .A(core__abc_22172_new_n6549_), .Y(core__abc_22172_new_n6550_));
INVX1 INVX1_1368 ( .A(core__abc_22172_new_n6472_), .Y(core__abc_22172_new_n6556_));
INVX1 INVX1_1369 ( .A(core__abc_22172_new_n6480_), .Y(core__abc_22172_new_n6557_));
INVX1 INVX1_137 ( .A(_abc_19873_new_n2626_), .Y(_abc_19873_new_n2627_));
INVX1 INVX1_1370 ( .A(core__abc_22172_new_n6541_), .Y(core__abc_22172_new_n6562_));
INVX1 INVX1_1371 ( .A(core__abc_22172_new_n6565_), .Y(core__abc_22172_new_n6566_));
INVX1 INVX1_1372 ( .A(core_v1_reg_10_), .Y(core__abc_22172_new_n6570_));
INVX1 INVX1_1373 ( .A(core__abc_22172_new_n6571_), .Y(core__abc_22172_new_n6572_));
INVX1 INVX1_1374 ( .A(core__abc_22172_new_n6574_), .Y(core__abc_22172_new_n6575_));
INVX1 INVX1_1375 ( .A(core_v1_reg_9_), .Y(core__abc_22172_new_n6579_));
INVX1 INVX1_1376 ( .A(core__abc_22172_new_n6582_), .Y(core__abc_22172_new_n6583_));
INVX1 INVX1_1377 ( .A(core__abc_22172_new_n6586_), .Y(core__abc_22172_new_n6587_));
INVX1 INVX1_1378 ( .A(core_v1_reg_8_), .Y(core__abc_22172_new_n6589_));
INVX1 INVX1_1379 ( .A(core__abc_22172_new_n6594_), .Y(core__abc_22172_new_n6595_));
INVX1 INVX1_138 ( .A(_abc_19873_new_n2631_), .Y(_abc_19873_new_n2632_));
INVX1 INVX1_1380 ( .A(core_v1_reg_7_), .Y(core__abc_22172_new_n6597_));
INVX1 INVX1_1381 ( .A(core__abc_22172_new_n6600_), .Y(core__abc_22172_new_n6601_));
INVX1 INVX1_1382 ( .A(core__abc_22172_new_n6604_), .Y(core__abc_22172_new_n6605_));
INVX1 INVX1_1383 ( .A(core_v1_reg_5_), .Y(core__abc_22172_new_n6608_));
INVX1 INVX1_1384 ( .A(core__abc_22172_new_n6611_), .Y(core__abc_22172_new_n6612_));
INVX1 INVX1_1385 ( .A(core__abc_22172_new_n6615_), .Y(core__abc_22172_new_n6616_));
INVX1 INVX1_1386 ( .A(core_v1_reg_6_), .Y(core__abc_22172_new_n6617_));
INVX1 INVX1_1387 ( .A(core__abc_22172_new_n6620_), .Y(core__abc_22172_new_n6622_));
INVX1 INVX1_1388 ( .A(core_v1_reg_4_), .Y(core__abc_22172_new_n6626_));
INVX1 INVX1_1389 ( .A(core__abc_22172_new_n6627_), .Y(core__abc_22172_new_n6628_));
INVX1 INVX1_139 ( .A(_abc_19873_new_n2637_), .Y(_abc_19873_new_n2638_));
INVX1 INVX1_1390 ( .A(core__abc_22172_new_n6631_), .Y(core__abc_22172_new_n6632_));
INVX1 INVX1_1391 ( .A(core_v1_reg_3_), .Y(core__abc_22172_new_n6633_));
INVX1 INVX1_1392 ( .A(core__abc_22172_new_n6636_), .Y(core__abc_22172_new_n6637_));
INVX1 INVX1_1393 ( .A(core__abc_22172_new_n6638_), .Y(core__abc_22172_new_n6639_));
INVX1 INVX1_1394 ( .A(core__abc_22172_new_n6630_), .Y(core__abc_22172_new_n6640_));
INVX1 INVX1_1395 ( .A(core__abc_22172_new_n6643_), .Y(core__abc_22172_new_n6644_));
INVX1 INVX1_1396 ( .A(core__abc_22172_new_n6613_), .Y(core__abc_22172_new_n6646_));
INVX1 INVX1_1397 ( .A(core__abc_22172_new_n6647_), .Y(core__abc_22172_new_n6648_));
INVX1 INVX1_1398 ( .A(core__abc_22172_new_n6602_), .Y(core__abc_22172_new_n6652_));
INVX1 INVX1_1399 ( .A(core__abc_22172_new_n6654_), .Y(core__abc_22172_new_n6655_));
INVX1 INVX1_14 ( .A(_abc_19873_new_n2129_), .Y(_abc_19873_new_n2130_));
INVX1 INVX1_140 ( .A(_abc_19873_new_n2642_), .Y(_abc_19873_new_n2643_));
INVX1 INVX1_1400 ( .A(core__abc_22172_new_n6576_), .Y(core__abc_22172_new_n6657_));
INVX1 INVX1_1401 ( .A(core_v1_reg_2_), .Y(core__abc_22172_new_n6662_));
INVX1 INVX1_1402 ( .A(core__abc_22172_new_n4139_), .Y(core__abc_22172_new_n6667_));
INVX1 INVX1_1403 ( .A(core__abc_22172_new_n6665_), .Y(core__abc_22172_new_n6668_));
INVX1 INVX1_1404 ( .A(core__abc_22172_new_n6673_), .Y(core__abc_22172_new_n6674_));
INVX1 INVX1_1405 ( .A(core__abc_22172_new_n6677_), .Y(core__abc_22172_new_n6678_));
INVX1 INVX1_1406 ( .A(core_v1_reg_0_), .Y(core__abc_22172_new_n6680_));
INVX1 INVX1_1407 ( .A(core__abc_22172_new_n6684_), .Y(core__abc_22172_new_n6685_));
INVX1 INVX1_1408 ( .A(core__abc_22172_new_n6683_), .Y(core__abc_22172_new_n6686_));
INVX1 INVX1_1409 ( .A(core__abc_22172_new_n6687_), .Y(core__abc_22172_new_n6688_));
INVX1 INVX1_141 ( .A(_abc_19873_new_n2647_), .Y(_abc_19873_new_n2648_));
INVX1 INVX1_1410 ( .A(core__abc_22172_new_n6691_), .Y(core__abc_22172_new_n6692_));
INVX1 INVX1_1411 ( .A(core__abc_22172_new_n6693_), .Y(core__abc_22172_new_n6694_));
INVX1 INVX1_1412 ( .A(core__abc_22172_new_n6695_), .Y(core__abc_22172_new_n6696_));
INVX1 INVX1_1413 ( .A(core__abc_22172_new_n6666_), .Y(core__abc_22172_new_n6699_));
INVX1 INVX1_1414 ( .A(core__abc_22172_new_n6705_), .Y(core__abc_22172_new_n6706_));
INVX1 INVX1_1415 ( .A(core__abc_22172_new_n6710_), .Y(core__abc_22172_new_n6711_));
INVX1 INVX1_1416 ( .A(core__abc_22172_new_n6712_), .Y(core__abc_22172_new_n6713_));
INVX1 INVX1_1417 ( .A(core__abc_22172_new_n6714_), .Y(core__abc_22172_new_n6715_));
INVX1 INVX1_1418 ( .A(core_v1_reg_61_), .Y(core__abc_22172_new_n6717_));
INVX1 INVX1_1419 ( .A(core__abc_22172_new_n6720_), .Y(core__abc_22172_new_n6721_));
INVX1 INVX1_142 ( .A(_abc_19873_new_n2652_), .Y(_abc_19873_new_n2653_));
INVX1 INVX1_1420 ( .A(core__abc_22172_new_n6727_), .Y(core__abc_22172_new_n6728_));
INVX1 INVX1_1421 ( .A(core_v1_reg_60_), .Y(core__abc_22172_new_n6730_));
INVX1 INVX1_1422 ( .A(core__abc_22172_new_n6734_), .Y(core__abc_22172_new_n6735_));
INVX1 INVX1_1423 ( .A(core__abc_22172_new_n6736_), .Y(core__abc_22172_new_n6737_));
INVX1 INVX1_1424 ( .A(core_v1_reg_59_), .Y(core__abc_22172_new_n6738_));
INVX1 INVX1_1425 ( .A(core__abc_22172_new_n6741_), .Y(core__abc_22172_new_n6742_));
INVX1 INVX1_1426 ( .A(core__abc_22172_new_n6749_), .Y(core__abc_22172_new_n6750_));
INVX1 INVX1_1427 ( .A(core_v1_reg_57_), .Y(core__abc_22172_new_n6754_));
INVX1 INVX1_1428 ( .A(core__abc_22172_new_n6757_), .Y(core__abc_22172_new_n6758_));
INVX1 INVX1_1429 ( .A(core__abc_22172_new_n6752_), .Y(core__abc_22172_new_n6762_));
INVX1 INVX1_143 ( .A(_abc_19873_new_n2657_), .Y(_abc_19873_new_n2658_));
INVX1 INVX1_1430 ( .A(core__abc_22172_new_n6765_), .Y(core__abc_22172_new_n6766_));
INVX1 INVX1_1431 ( .A(core_v1_reg_56_), .Y(core__abc_22172_new_n6768_));
INVX1 INVX1_1432 ( .A(core__abc_22172_new_n5348_), .Y(core__abc_22172_new_n6770_));
INVX1 INVX1_1433 ( .A(core__abc_22172_new_n6772_), .Y(core__abc_22172_new_n6773_));
INVX1 INVX1_1434 ( .A(core__abc_22172_new_n6775_), .Y(core__abc_22172_new_n6776_));
INVX1 INVX1_1435 ( .A(core_v1_reg_55_), .Y(core__abc_22172_new_n6777_));
INVX1 INVX1_1436 ( .A(core__abc_22172_new_n6780_), .Y(core__abc_22172_new_n6781_));
INVX1 INVX1_1437 ( .A(core_v1_reg_54_), .Y(core__abc_22172_new_n6783_));
INVX1 INVX1_1438 ( .A(core__abc_22172_new_n5254_), .Y(core__abc_22172_new_n6785_));
INVX1 INVX1_1439 ( .A(core__abc_22172_new_n6787_), .Y(core__abc_22172_new_n6788_));
INVX1 INVX1_144 ( .A(_abc_19873_new_n2662_), .Y(_abc_19873_new_n2663_));
INVX1 INVX1_1440 ( .A(core_v1_reg_53_), .Y(core__abc_22172_new_n6791_));
INVX1 INVX1_1441 ( .A(core__abc_22172_new_n6795_), .Y(core__abc_22172_new_n6796_));
INVX1 INVX1_1442 ( .A(core_v1_reg_52_), .Y(core__abc_22172_new_n6797_));
INVX1 INVX1_1443 ( .A(core__abc_22172_new_n6801_), .Y(core__abc_22172_new_n6802_));
INVX1 INVX1_1444 ( .A(core__abc_22172_new_n6803_), .Y(core__abc_22172_new_n6804_));
INVX1 INVX1_1445 ( .A(core__abc_22172_new_n6806_), .Y(core__abc_22172_new_n6807_));
INVX1 INVX1_1446 ( .A(core__abc_22172_new_n6800_), .Y(core__abc_22172_new_n6809_));
INVX1 INVX1_1447 ( .A(core__abc_22172_new_n6794_), .Y(core__abc_22172_new_n6814_));
INVX1 INVX1_1448 ( .A(core__abc_22172_new_n6822_), .Y(core__abc_22172_new_n6823_));
INVX1 INVX1_1449 ( .A(core__abc_22172_new_n6832_), .Y(core__abc_22172_new_n6833_));
INVX1 INVX1_145 ( .A(_abc_19873_new_n2667_), .Y(_abc_19873_new_n2668_));
INVX1 INVX1_1450 ( .A(core__abc_22172_new_n6641_), .Y(core__abc_22172_new_n6840_));
INVX1 INVX1_1451 ( .A(core__abc_22172_new_n6843_), .Y(core__abc_22172_new_n6844_));
INVX1 INVX1_1452 ( .A(core_v1_reg_19_), .Y(core__abc_22172_new_n6852_));
INVX1 INVX1_1453 ( .A(core__abc_22172_new_n6855_), .Y(core__abc_22172_new_n6856_));
INVX1 INVX1_1454 ( .A(core__abc_22172_new_n6859_), .Y(core__abc_22172_new_n6860_));
INVX1 INVX1_1455 ( .A(core__abc_22172_new_n6851_), .Y(core__abc_22172_new_n6862_));
INVX1 INVX1_1456 ( .A(core__abc_22172_new_n6864_), .Y(core__abc_22172_new_n6865_));
INVX1 INVX1_1457 ( .A(core_key_0_), .Y(core__abc_22172_new_n6867_));
INVX1 INVX1_1458 ( .A(core_long), .Y(core__abc_22172_new_n6870_));
INVX1 INVX1_1459 ( .A(core__abc_22172_new_n6877_), .Y(core__abc_22172_new_n6878_));
INVX1 INVX1_146 ( .A(_abc_19873_new_n2672_), .Y(_abc_19873_new_n2673_));
INVX1 INVX1_1460 ( .A(core__abc_22172_new_n5168_), .Y(core__abc_22172_new_n6884_));
INVX1 INVX1_1461 ( .A(core_v1_reg_20_), .Y(core__abc_22172_new_n6885_));
INVX1 INVX1_1462 ( .A(core__abc_22172_new_n6886_), .Y(core__abc_22172_new_n6887_));
INVX1 INVX1_1463 ( .A(core__abc_22172_new_n6889_), .Y(core__abc_22172_new_n6891_));
INVX1 INVX1_1464 ( .A(core__abc_22172_new_n6857_), .Y(core__abc_22172_new_n6894_));
INVX1 INVX1_1465 ( .A(core__abc_22172_new_n6861_), .Y(core__abc_22172_new_n6895_));
INVX1 INVX1_1466 ( .A(core__abc_22172_new_n6898_), .Y(core__abc_22172_new_n6899_));
INVX1 INVX1_1467 ( .A(core__abc_22172_new_n6900_), .Y(core__abc_22172_new_n6901_));
INVX1 INVX1_1468 ( .A(core__abc_22172_new_n6893_), .Y(core__abc_22172_new_n6911_));
INVX1 INVX1_1469 ( .A(core_v1_reg_21_), .Y(core__abc_22172_new_n6917_));
INVX1 INVX1_147 ( .A(_abc_19873_new_n2677_), .Y(_abc_19873_new_n2678_));
INVX1 INVX1_1470 ( .A(core__abc_22172_new_n6920_), .Y(core__abc_22172_new_n6922_));
INVX1 INVX1_1471 ( .A(core__abc_22172_new_n6924_), .Y(core__abc_22172_new_n6925_));
INVX1 INVX1_1472 ( .A(core__abc_22172_new_n6926_), .Y(core__abc_22172_new_n6927_));
INVX1 INVX1_1473 ( .A(core__abc_22172_new_n6923_), .Y(core__abc_22172_new_n6939_));
INVX1 INVX1_1474 ( .A(core__abc_22172_new_n6942_), .Y(core__abc_22172_new_n6943_));
INVX1 INVX1_1475 ( .A(core__abc_22172_new_n6944_), .Y(core__abc_22172_new_n6946_));
INVX1 INVX1_1476 ( .A(core__abc_22172_new_n6949_), .Y(core__abc_22172_new_n6950_));
INVX1 INVX1_1477 ( .A(core_v1_reg_23_), .Y(core__abc_22172_new_n6962_));
INVX1 INVX1_1478 ( .A(core__abc_22172_new_n6965_), .Y(core__abc_22172_new_n6967_));
INVX1 INVX1_1479 ( .A(core__abc_22172_new_n6969_), .Y(core__abc_22172_new_n6970_));
INVX1 INVX1_148 ( .A(_abc_19873_new_n2682_), .Y(_abc_19873_new_n2683_));
INVX1 INVX1_1480 ( .A(core__abc_22172_new_n6945_), .Y(core__abc_22172_new_n6971_));
INVX1 INVX1_1481 ( .A(core__abc_22172_new_n6974_), .Y(core__abc_22172_new_n6975_));
INVX1 INVX1_1482 ( .A(core__abc_22172_new_n6978_), .Y(core__abc_22172_new_n6979_));
INVX1 INVX1_1483 ( .A(core_v1_reg_24_), .Y(core__abc_22172_new_n6993_));
INVX1 INVX1_1484 ( .A(core__abc_22172_new_n3480_), .Y(core__abc_22172_new_n6994_));
INVX1 INVX1_1485 ( .A(core__abc_22172_new_n6998_), .Y(core__abc_22172_new_n6999_));
INVX1 INVX1_1486 ( .A(core__abc_22172_new_n7001_), .Y(core__abc_22172_new_n7002_));
INVX1 INVX1_1487 ( .A(core__abc_22172_new_n7003_), .Y(core__abc_22172_new_n7004_));
INVX1 INVX1_1488 ( .A(core__abc_22172_new_n7006_), .Y(core__abc_22172_new_n7007_));
INVX1 INVX1_1489 ( .A(core_key_5_), .Y(core__abc_22172_new_n7009_));
INVX1 INVX1_149 ( .A(_abc_19873_new_n2687_), .Y(_abc_19873_new_n2688_));
INVX1 INVX1_1490 ( .A(core_v1_reg_25_), .Y(core__abc_22172_new_n7018_));
INVX1 INVX1_1491 ( .A(core__abc_22172_new_n7021_), .Y(core__abc_22172_new_n7023_));
INVX1 INVX1_1492 ( .A(core__abc_22172_new_n6968_), .Y(core__abc_22172_new_n7026_));
INVX1 INVX1_1493 ( .A(core__abc_22172_new_n7029_), .Y(core__abc_22172_new_n7030_));
INVX1 INVX1_1494 ( .A(core__abc_22172_new_n7033_), .Y(core__abc_22172_new_n7034_));
INVX1 INVX1_1495 ( .A(core__abc_22172_new_n7036_), .Y(core__abc_22172_new_n7037_));
INVX1 INVX1_1496 ( .A(core_key_6_), .Y(core__abc_22172_new_n7039_));
INVX1 INVX1_1497 ( .A(core__abc_22172_new_n7024_), .Y(core__abc_22172_new_n7048_));
INVX1 INVX1_1498 ( .A(core__abc_22172_new_n5449_), .Y(core__abc_22172_new_n7050_));
INVX1 INVX1_1499 ( .A(core_v1_reg_26_), .Y(core__abc_22172_new_n7051_));
INVX1 INVX1_15 ( .A(\write_data[2] ), .Y(_abc_19873_new_n2134_));
INVX1 INVX1_150 ( .A(_abc_19873_new_n2692_), .Y(_abc_19873_new_n2693_));
INVX1 INVX1_1500 ( .A(core__abc_22172_new_n7054_), .Y(core__abc_22172_new_n7055_));
INVX1 INVX1_1501 ( .A(core__abc_22172_new_n7059_), .Y(core__abc_22172_new_n7060_));
INVX1 INVX1_1502 ( .A(core__abc_22172_new_n7072_), .Y(core__abc_22172_new_n7073_));
INVX1 INVX1_1503 ( .A(core__abc_22172_new_n7076_), .Y(core__abc_22172_new_n7077_));
INVX1 INVX1_1504 ( .A(core__abc_22172_new_n7081_), .Y(core__abc_22172_new_n7082_));
INVX1 INVX1_1505 ( .A(core__abc_22172_new_n7057_), .Y(core__abc_22172_new_n7085_));
INVX1 INVX1_1506 ( .A(core__abc_22172_new_n7087_), .Y(core__abc_22172_new_n7088_));
INVX1 INVX1_1507 ( .A(core__abc_22172_new_n7091_), .Y(core__abc_22172_new_n7092_));
INVX1 INVX1_1508 ( .A(core_v1_reg_27_), .Y(core__abc_22172_new_n7094_));
INVX1 INVX1_1509 ( .A(core__abc_22172_new_n7097_), .Y(core__abc_22172_new_n7099_));
INVX1 INVX1_151 ( .A(_abc_19873_new_n2697_), .Y(_abc_19873_new_n2698_));
INVX1 INVX1_1510 ( .A(core__abc_22172_new_n7101_), .Y(core__abc_22172_new_n7102_));
INVX1 INVX1_1511 ( .A(core__abc_22172_new_n7093_), .Y(core__abc_22172_new_n7104_));
INVX1 INVX1_1512 ( .A(core__abc_22172_new_n7106_), .Y(core__abc_22172_new_n7107_));
INVX1 INVX1_1513 ( .A(core__abc_22172_new_n6880_), .Y(core__abc_22172_new_n7114_));
INVX1 INVX1_1514 ( .A(core_v1_reg_28_), .Y(core__abc_22172_new_n7118_));
INVX1 INVX1_1515 ( .A(core__abc_22172_new_n3742_), .Y(core__abc_22172_new_n7119_));
INVX1 INVX1_1516 ( .A(core__abc_22172_new_n7124_), .Y(core__abc_22172_new_n7125_));
INVX1 INVX1_1517 ( .A(core__abc_22172_new_n7126_), .Y(core__abc_22172_new_n7127_));
INVX1 INVX1_1518 ( .A(core__abc_22172_new_n7100_), .Y(core__abc_22172_new_n7128_));
INVX1 INVX1_1519 ( .A(core__abc_22172_new_n7103_), .Y(core__abc_22172_new_n7129_));
INVX1 INVX1_152 ( .A(_abc_19873_new_n2702_), .Y(_abc_19873_new_n2703_));
INVX1 INVX1_1520 ( .A(core__abc_22172_new_n7132_), .Y(core__abc_22172_new_n7133_));
INVX1 INVX1_1521 ( .A(core__abc_22172_new_n7134_), .Y(core__abc_22172_new_n7135_));
INVX1 INVX1_1522 ( .A(core_key_9_), .Y(core__abc_22172_new_n7137_));
INVX1 INVX1_1523 ( .A(core__abc_22172_new_n7149_), .Y(core__abc_22172_new_n7150_));
INVX1 INVX1_1524 ( .A(core_v1_reg_29_), .Y(core__abc_22172_new_n7152_));
INVX1 INVX1_1525 ( .A(core__abc_22172_new_n7155_), .Y(core__abc_22172_new_n7156_));
INVX1 INVX1_1526 ( .A(core__abc_22172_new_n7159_), .Y(core__abc_22172_new_n7160_));
INVX1 INVX1_1527 ( .A(core__abc_22172_new_n7161_), .Y(core__abc_22172_new_n7162_));
INVX1 INVX1_1528 ( .A(core__abc_22172_new_n7157_), .Y(core__abc_22172_new_n7174_));
INVX1 INVX1_1529 ( .A(core_v1_reg_30_), .Y(core__abc_22172_new_n7176_));
INVX1 INVX1_153 ( .A(_abc_19873_new_n2707_), .Y(_abc_19873_new_n2708_));
INVX1 INVX1_1530 ( .A(core__abc_22172_new_n7181_), .Y(core__abc_22172_new_n7182_));
INVX1 INVX1_1531 ( .A(core__abc_22172_new_n7183_), .Y(core__abc_22172_new_n7184_));
INVX1 INVX1_1532 ( .A(core__abc_22172_new_n7185_), .Y(core__abc_22172_new_n7186_));
INVX1 INVX1_1533 ( .A(core__abc_22172_new_n7180_), .Y(core__abc_22172_new_n7200_));
INVX1 INVX1_1534 ( .A(core_v1_reg_31_), .Y(core__abc_22172_new_n7207_));
INVX1 INVX1_1535 ( .A(core__abc_22172_new_n7210_), .Y(core__abc_22172_new_n7211_));
INVX1 INVX1_1536 ( .A(core__abc_22172_new_n7214_), .Y(core__abc_22172_new_n7215_));
INVX1 INVX1_1537 ( .A(core__abc_22172_new_n7206_), .Y(core__abc_22172_new_n7217_));
INVX1 INVX1_1538 ( .A(core__abc_22172_new_n7219_), .Y(core__abc_22172_new_n7220_));
INVX1 INVX1_1539 ( .A(core_key_12_), .Y(core__abc_22172_new_n7222_));
INVX1 INVX1_154 ( .A(_abc_19873_new_n2712_), .Y(_abc_19873_new_n2713_));
INVX1 INVX1_1540 ( .A(core__abc_22172_new_n3325_), .Y(core__abc_22172_new_n7232_));
INVX1 INVX1_1541 ( .A(core_v1_reg_32_), .Y(core__abc_22172_new_n7233_));
INVX1 INVX1_1542 ( .A(core__abc_22172_new_n7236_), .Y(core__abc_22172_new_n7237_));
INVX1 INVX1_1543 ( .A(core__abc_22172_new_n7231_), .Y(core__abc_22172_new_n7242_));
INVX1 INVX1_1544 ( .A(core__abc_22172_new_n7240_), .Y(core__abc_22172_new_n7243_));
INVX1 INVX1_1545 ( .A(core_key_13_), .Y(core__abc_22172_new_n7247_));
INVX1 INVX1_1546 ( .A(core__abc_22172_new_n7239_), .Y(core__abc_22172_new_n7256_));
INVX1 INVX1_1547 ( .A(core__abc_22172_new_n7258_), .Y(core__abc_22172_new_n7259_));
INVX1 INVX1_1548 ( .A(core__abc_22172_new_n7260_), .Y(core__abc_22172_new_n7261_));
INVX1 INVX1_1549 ( .A(core__abc_22172_new_n7263_), .Y(core__abc_22172_new_n7264_));
INVX1 INVX1_155 ( .A(_abc_19873_new_n2717_), .Y(_abc_19873_new_n2718_));
INVX1 INVX1_1550 ( .A(core_v1_reg_33_), .Y(core__abc_22172_new_n7265_));
INVX1 INVX1_1551 ( .A(core__abc_22172_new_n4078_), .Y(core__abc_22172_new_n7266_));
INVX1 INVX1_1552 ( .A(core__abc_22172_new_n7269_), .Y(core__abc_22172_new_n7271_));
INVX1 INVX1_1553 ( .A(core__abc_22172_new_n7273_), .Y(core__abc_22172_new_n7274_));
INVX1 INVX1_1554 ( .A(core__abc_22172_new_n7277_), .Y(core__abc_22172_new_n7278_));
INVX1 INVX1_1555 ( .A(core_key_14_), .Y(core__abc_22172_new_n7280_));
INVX1 INVX1_1556 ( .A(core__abc_22172_new_n7289_), .Y(core__abc_22172_new_n7290_));
INVX1 INVX1_1557 ( .A(core__abc_22172_new_n7292_), .Y(core__abc_22172_new_n7293_));
INVX1 INVX1_1558 ( .A(core__abc_22172_new_n7291_), .Y(core__abc_22172_new_n7296_));
INVX1 INVX1_1559 ( .A(core__abc_22172_new_n7305_), .Y(core__abc_22172_new_n7306_));
INVX1 INVX1_156 ( .A(_abc_19873_new_n2722_), .Y(_abc_19873_new_n2723_));
INVX1 INVX1_1560 ( .A(core__abc_22172_new_n7203_), .Y(core__abc_22172_new_n7316_));
INVX1 INVX1_1561 ( .A(core__abc_22172_new_n7322_), .Y(core__abc_22172_new_n7323_));
INVX1 INVX1_1562 ( .A(core__abc_22172_new_n7204_), .Y(core__abc_22172_new_n7326_));
INVX1 INVX1_1563 ( .A(core__abc_22172_new_n7334_), .Y(core__abc_22172_new_n7335_));
INVX1 INVX1_1564 ( .A(core__abc_22172_new_n7336_), .Y(core__abc_22172_new_n7337_));
INVX1 INVX1_1565 ( .A(core_v1_reg_35_), .Y(core__abc_22172_new_n7338_));
INVX1 INVX1_1566 ( .A(core__abc_22172_new_n7341_), .Y(core__abc_22172_new_n7342_));
INVX1 INVX1_1567 ( .A(core__abc_22172_new_n7345_), .Y(core__abc_22172_new_n7346_));
INVX1 INVX1_1568 ( .A(core__abc_22172_new_n7349_), .Y(core__abc_22172_new_n7350_));
INVX1 INVX1_1569 ( .A(core_key_16_), .Y(core__abc_22172_new_n7352_));
INVX1 INVX1_157 ( .A(_abc_19873_new_n2727_), .Y(_abc_19873_new_n2728_));
INVX1 INVX1_1570 ( .A(core__abc_22172_new_n7343_), .Y(core__abc_22172_new_n7361_));
INVX1 INVX1_1571 ( .A(core__abc_22172_new_n7347_), .Y(core__abc_22172_new_n7362_));
INVX1 INVX1_1572 ( .A(core_v1_reg_36_), .Y(core__abc_22172_new_n7364_));
INVX1 INVX1_1573 ( .A(core__abc_22172_new_n4282_), .Y(core__abc_22172_new_n7365_));
INVX1 INVX1_1574 ( .A(core__abc_22172_new_n7368_), .Y(core__abc_22172_new_n7369_));
INVX1 INVX1_1575 ( .A(core__abc_22172_new_n7370_), .Y(core__abc_22172_new_n7371_));
INVX1 INVX1_1576 ( .A(core__abc_22172_new_n7372_), .Y(core__abc_22172_new_n7373_));
INVX1 INVX1_1577 ( .A(core__abc_22172_new_n7363_), .Y(core__abc_22172_new_n7376_));
INVX1 INVX1_1578 ( .A(core__abc_22172_new_n7374_), .Y(core__abc_22172_new_n7377_));
INVX1 INVX1_1579 ( .A(core__abc_22172_new_n7379_), .Y(core__abc_22172_new_n7380_));
INVX1 INVX1_158 ( .A(_abc_19873_new_n2732_), .Y(_abc_19873_new_n2733_));
INVX1 INVX1_1580 ( .A(core_v1_reg_37_), .Y(core__abc_22172_new_n7390_));
INVX1 INVX1_1581 ( .A(core__abc_22172_new_n7393_), .Y(core__abc_22172_new_n7394_));
INVX1 INVX1_1582 ( .A(core__abc_22172_new_n7397_), .Y(core__abc_22172_new_n7398_));
INVX1 INVX1_1583 ( .A(core__abc_22172_new_n7401_), .Y(core__abc_22172_new_n7402_));
INVX1 INVX1_1584 ( .A(core__abc_22172_new_n7405_), .Y(core__abc_22172_new_n7406_));
INVX1 INVX1_1585 ( .A(core_key_18_), .Y(core__abc_22172_new_n7408_));
INVX1 INVX1_1586 ( .A(core_v1_reg_38_), .Y(core__abc_22172_new_n7418_));
INVX1 INVX1_1587 ( .A(core__abc_22172_new_n4403_), .Y(core__abc_22172_new_n7419_));
INVX1 INVX1_1588 ( .A(core__abc_22172_new_n7422_), .Y(core__abc_22172_new_n7423_));
INVX1 INVX1_1589 ( .A(core__abc_22172_new_n7424_), .Y(core__abc_22172_new_n7425_));
INVX1 INVX1_159 ( .A(_abc_19873_new_n2737_), .Y(_abc_19873_new_n2738_));
INVX1 INVX1_1590 ( .A(core__abc_22172_new_n7426_), .Y(core__abc_22172_new_n7427_));
INVX1 INVX1_1591 ( .A(core__abc_22172_new_n7417_), .Y(core__abc_22172_new_n7430_));
INVX1 INVX1_1592 ( .A(core__abc_22172_new_n7428_), .Y(core__abc_22172_new_n7431_));
INVX1 INVX1_1593 ( .A(core__abc_22172_new_n7444_), .Y(core__abc_22172_new_n7445_));
INVX1 INVX1_1594 ( .A(core__abc_22172_new_n7447_), .Y(core__abc_22172_new_n7448_));
INVX1 INVX1_1595 ( .A(core__abc_22172_new_n7452_), .Y(core__abc_22172_new_n7453_));
INVX1 INVX1_1596 ( .A(core_v1_reg_39_), .Y(core__abc_22172_new_n7456_));
INVX1 INVX1_1597 ( .A(core__abc_22172_new_n7459_), .Y(core__abc_22172_new_n7460_));
INVX1 INVX1_1598 ( .A(core__abc_22172_new_n7464_), .Y(core__abc_22172_new_n7465_));
INVX1 INVX1_1599 ( .A(core__abc_22172_new_n7467_), .Y(core__abc_22172_new_n7468_));
INVX1 INVX1_16 ( .A(_abc_19873_new_n2135_), .Y(_abc_19873_new_n2136_));
INVX1 INVX1_160 ( .A(_abc_19873_new_n2742_), .Y(_abc_19873_new_n2743_));
INVX1 INVX1_1600 ( .A(core__abc_22172_new_n7461_), .Y(core__abc_22172_new_n7478_));
INVX1 INVX1_1601 ( .A(core__abc_22172_new_n7479_), .Y(core__abc_22172_new_n7480_));
INVX1 INVX1_1602 ( .A(core__abc_22172_new_n3845_), .Y(core__abc_22172_new_n7481_));
INVX1 INVX1_1603 ( .A(core_v1_reg_40_), .Y(core__abc_22172_new_n7482_));
INVX1 INVX1_1604 ( .A(core__abc_22172_new_n7485_), .Y(core__abc_22172_new_n7486_));
INVX1 INVX1_1605 ( .A(core__abc_22172_new_n7487_), .Y(core__abc_22172_new_n7488_));
INVX1 INVX1_1606 ( .A(core__abc_22172_new_n7489_), .Y(core__abc_22172_new_n7490_));
INVX1 INVX1_1607 ( .A(core__abc_22172_new_n7491_), .Y(core__abc_22172_new_n7493_));
INVX1 INVX1_1608 ( .A(core_key_21_), .Y(core__abc_22172_new_n7497_));
INVX1 INVX1_1609 ( .A(core_v1_reg_41_), .Y(core__abc_22172_new_n7506_));
INVX1 INVX1_161 ( .A(_abc_19873_new_n2747_), .Y(_abc_19873_new_n2748_));
INVX1 INVX1_1610 ( .A(core__abc_22172_new_n4583_), .Y(core__abc_22172_new_n7507_));
INVX1 INVX1_1611 ( .A(core__abc_22172_new_n7510_), .Y(core__abc_22172_new_n7511_));
INVX1 INVX1_1612 ( .A(core__abc_22172_new_n7520_), .Y(core__abc_22172_new_n7521_));
INVX1 INVX1_1613 ( .A(core__abc_22172_new_n7523_), .Y(core__abc_22172_new_n7524_));
INVX1 INVX1_1614 ( .A(core_key_22_), .Y(core__abc_22172_new_n7526_));
INVX1 INVX1_1615 ( .A(core__abc_22172_new_n7512_), .Y(core__abc_22172_new_n7535_));
INVX1 INVX1_1616 ( .A(core__abc_22172_new_n3972_), .Y(core__abc_22172_new_n7537_));
INVX1 INVX1_1617 ( .A(core_v1_reg_42_), .Y(core__abc_22172_new_n7538_));
INVX1 INVX1_1618 ( .A(core__abc_22172_new_n7541_), .Y(core__abc_22172_new_n7542_));
INVX1 INVX1_1619 ( .A(core__abc_22172_new_n7543_), .Y(core__abc_22172_new_n7544_));
INVX1 INVX1_162 ( .A(_abc_19873_new_n2752_), .Y(_abc_19873_new_n2753_));
INVX1 INVX1_1620 ( .A(core__abc_22172_new_n7545_), .Y(core__abc_22172_new_n7546_));
INVX1 INVX1_1621 ( .A(core__abc_22172_new_n7547_), .Y(core__abc_22172_new_n7548_));
INVX1 INVX1_1622 ( .A(core__abc_22172_new_n7536_), .Y(core__abc_22172_new_n7550_));
INVX1 INVX1_1623 ( .A(core__abc_22172_new_n7552_), .Y(core__abc_22172_new_n7553_));
INVX1 INVX1_1624 ( .A(core__abc_22172_new_n7450_), .Y(core__abc_22172_new_n7563_));
INVX1 INVX1_1625 ( .A(core__abc_22172_new_n7515_), .Y(core__abc_22172_new_n7564_));
INVX1 INVX1_1626 ( .A(core__abc_22172_new_n7514_), .Y(core__abc_22172_new_n7565_));
INVX1 INVX1_1627 ( .A(core__abc_22172_new_n7518_), .Y(core__abc_22172_new_n7569_));
INVX1 INVX1_1628 ( .A(core_v1_reg_43_), .Y(core__abc_22172_new_n7578_));
INVX1 INVX1_1629 ( .A(core__abc_22172_new_n7581_), .Y(core__abc_22172_new_n7582_));
INVX1 INVX1_163 ( .A(_abc_19873_new_n2757_), .Y(_abc_19873_new_n2758_));
INVX1 INVX1_1630 ( .A(core__abc_22172_new_n7585_), .Y(core__abc_22172_new_n7586_));
INVX1 INVX1_1631 ( .A(core__abc_22172_new_n7577_), .Y(core__abc_22172_new_n7588_));
INVX1 INVX1_1632 ( .A(core__abc_22172_new_n7590_), .Y(core__abc_22172_new_n7591_));
INVX1 INVX1_1633 ( .A(core__abc_22172_new_n7602_), .Y(core__abc_22172_new_n7603_));
INVX1 INVX1_1634 ( .A(core__abc_22172_new_n7606_), .Y(core__abc_22172_new_n7607_));
INVX1 INVX1_1635 ( .A(core__abc_22172_new_n7605_), .Y(core__abc_22172_new_n7608_));
INVX1 INVX1_1636 ( .A(core__abc_22172_new_n7609_), .Y(core__abc_22172_new_n7610_));
INVX1 INVX1_1637 ( .A(core__abc_22172_new_n7601_), .Y(core__abc_22172_new_n7613_));
INVX1 INVX1_1638 ( .A(core__abc_22172_new_n7611_), .Y(core__abc_22172_new_n7614_));
INVX1 INVX1_1639 ( .A(core_key_25_), .Y(core__abc_22172_new_n7618_));
INVX1 INVX1_164 ( .A(_abc_19873_new_n2762_), .Y(_abc_19873_new_n2763_));
INVX1 INVX1_1640 ( .A(core_v1_reg_45_), .Y(core__abc_22172_new_n7627_));
INVX1 INVX1_1641 ( .A(core__abc_22172_new_n7630_), .Y(core__abc_22172_new_n7631_));
INVX1 INVX1_1642 ( .A(core__abc_22172_new_n7634_), .Y(core__abc_22172_new_n7635_));
INVX1 INVX1_1643 ( .A(core__abc_22172_new_n7583_), .Y(core__abc_22172_new_n7638_));
INVX1 INVX1_1644 ( .A(core__abc_22172_new_n7640_), .Y(core__abc_22172_new_n7641_));
INVX1 INVX1_1645 ( .A(core__abc_22172_new_n7643_), .Y(core__abc_22172_new_n7644_));
INVX1 INVX1_1646 ( .A(core_key_26_), .Y(core__abc_22172_new_n7648_));
INVX1 INVX1_1647 ( .A(core__abc_22172_new_n7632_), .Y(core__abc_22172_new_n7657_));
INVX1 INVX1_1648 ( .A(core__abc_22172_new_n7658_), .Y(core__abc_22172_new_n7659_));
INVX1 INVX1_1649 ( .A(core_v1_reg_46_), .Y(core__abc_22172_new_n7660_));
INVX1 INVX1_165 ( .A(_abc_19873_new_n2767_), .Y(_abc_19873_new_n2768_));
INVX1 INVX1_1650 ( .A(core__abc_22172_new_n7663_), .Y(core__abc_22172_new_n7664_));
INVX1 INVX1_1651 ( .A(core__abc_22172_new_n7667_), .Y(core__abc_22172_new_n7668_));
INVX1 INVX1_1652 ( .A(core_key_27_), .Y(core__abc_22172_new_n7673_));
INVX1 INVX1_1653 ( .A(core__abc_22172_new_n7689_), .Y(core__abc_22172_new_n7690_));
INVX1 INVX1_1654 ( .A(core_v1_reg_47_), .Y(core__abc_22172_new_n7691_));
INVX1 INVX1_1655 ( .A(core__abc_22172_new_n7694_), .Y(core__abc_22172_new_n7695_));
INVX1 INVX1_1656 ( .A(core__abc_22172_new_n7698_), .Y(core__abc_22172_new_n7700_));
INVX1 INVX1_1657 ( .A(core__abc_22172_new_n7702_), .Y(core__abc_22172_new_n7703_));
INVX1 INVX1_1658 ( .A(core_v1_reg_48_), .Y(core__abc_22172_new_n7713_));
INVX1 INVX1_1659 ( .A(core__abc_22172_new_n7716_), .Y(core__abc_22172_new_n7718_));
INVX1 INVX1_166 ( .A(_abc_19873_new_n2772_), .Y(_abc_19873_new_n2773_));
INVX1 INVX1_1660 ( .A(core__abc_22172_new_n7721_), .Y(core__abc_22172_new_n7722_));
INVX1 INVX1_1661 ( .A(core__abc_22172_new_n7720_), .Y(core__abc_22172_new_n7724_));
INVX1 INVX1_1662 ( .A(core__abc_22172_new_n7726_), .Y(core__abc_22172_new_n7727_));
INVX1 INVX1_1663 ( .A(core_key_29_), .Y(core__abc_22172_new_n7729_));
INVX1 INVX1_1664 ( .A(core__abc_22172_new_n7742_), .Y(core__abc_22172_new_n7743_));
INVX1 INVX1_1665 ( .A(core_v1_reg_49_), .Y(core__abc_22172_new_n7744_));
INVX1 INVX1_1666 ( .A(core__abc_22172_new_n7747_), .Y(core__abc_22172_new_n7748_));
INVX1 INVX1_1667 ( .A(core__abc_22172_new_n7751_), .Y(core__abc_22172_new_n7753_));
INVX1 INVX1_1668 ( .A(core__abc_22172_new_n7755_), .Y(core__abc_22172_new_n7756_));
INVX1 INVX1_1669 ( .A(core_key_30_), .Y(core__abc_22172_new_n7758_));
INVX1 INVX1_167 ( .A(_abc_19873_new_n2777_), .Y(_abc_19873_new_n2778_));
INVX1 INVX1_1670 ( .A(core_v1_reg_50_), .Y(core__abc_22172_new_n7768_));
INVX1 INVX1_1671 ( .A(core__abc_22172_new_n7771_), .Y(core__abc_22172_new_n7772_));
INVX1 INVX1_1672 ( .A(core__abc_22172_new_n7767_), .Y(core__abc_22172_new_n7777_));
INVX1 INVX1_1673 ( .A(core__abc_22172_new_n7775_), .Y(core__abc_22172_new_n7778_));
INVX1 INVX1_1674 ( .A(core_key_32_), .Y(core__abc_22172_new_n7790_));
INVX1 INVX1_1675 ( .A(core__abc_22172_new_n7793_), .Y(core__abc_22172_new_n7794_));
INVX1 INVX1_1676 ( .A(core__abc_22172_new_n6812_), .Y(core__abc_22172_new_n7804_));
INVX1 INVX1_1677 ( .A(core__abc_22172_new_n6817_), .Y(core__abc_22172_new_n7812_));
INVX1 INVX1_1678 ( .A(core_key_34_), .Y(core__abc_22172_new_n7816_));
INVX1 INVX1_1679 ( .A(core__abc_22172_new_n6818_), .Y(core__abc_22172_new_n7825_));
INVX1 INVX1_168 ( .A(_abc_19873_new_n2782_), .Y(_abc_19873_new_n2783_));
INVX1 INVX1_1680 ( .A(core__abc_22172_new_n6789_), .Y(core__abc_22172_new_n7826_));
INVX1 INVX1_1681 ( .A(core__abc_22172_new_n7827_), .Y(core__abc_22172_new_n7828_));
INVX1 INVX1_1682 ( .A(core__abc_22172_new_n7831_), .Y(core__abc_22172_new_n7832_));
INVX1 INVX1_1683 ( .A(core__abc_22172_new_n6824_), .Y(core__abc_22172_new_n7842_));
INVX1 INVX1_1684 ( .A(core__abc_22172_new_n6825_), .Y(core__abc_22172_new_n7854_));
INVX1 INVX1_1685 ( .A(core__abc_22172_new_n6774_), .Y(core__abc_22172_new_n7855_));
INVX1 INVX1_1686 ( .A(core__abc_22172_new_n7857_), .Y(core__abc_22172_new_n7858_));
INVX1 INVX1_1687 ( .A(core__abc_22172_new_n7860_), .Y(core__abc_22172_new_n7861_));
INVX1 INVX1_1688 ( .A(core_key_37_), .Y(core__abc_22172_new_n7863_));
INVX1 INVX1_1689 ( .A(core__abc_22172_new_n7872_), .Y(core__abc_22172_new_n7873_));
INVX1 INVX1_169 ( .A(_abc_19873_new_n2787_), .Y(_abc_19873_new_n2788_));
INVX1 INVX1_1690 ( .A(core_key_38_), .Y(core__abc_22172_new_n7877_));
INVX1 INVX1_1691 ( .A(core__abc_22172_new_n6763_), .Y(core__abc_22172_new_n7888_));
INVX1 INVX1_1692 ( .A(core__abc_22172_new_n7886_), .Y(core__abc_22172_new_n7889_));
INVX1 INVX1_1693 ( .A(core__abc_22172_new_n7901_), .Y(core__abc_22172_new_n7902_));
INVX1 INVX1_1694 ( .A(core_key_40_), .Y(core__abc_22172_new_n7906_));
INVX1 INVX1_1695 ( .A(core__abc_22172_new_n6830_), .Y(core__abc_22172_new_n7915_));
INVX1 INVX1_1696 ( .A(core__abc_22172_new_n7916_), .Y(core__abc_22172_new_n7917_));
INVX1 INVX1_1697 ( .A(core__abc_22172_new_n7920_), .Y(core__abc_22172_new_n7921_));
INVX1 INVX1_1698 ( .A(core_key_41_), .Y(core__abc_22172_new_n7923_));
INVX1 INVX1_1699 ( .A(core__abc_22172_new_n7934_), .Y(core__abc_22172_new_n7935_));
INVX1 INVX1_17 ( .A(\write_data[3] ), .Y(_abc_19873_new_n2140_));
INVX1 INVX1_170 ( .A(_abc_19873_new_n2792_), .Y(_abc_19873_new_n2793_));
INVX1 INVX1_1700 ( .A(core_key_42_), .Y(core__abc_22172_new_n7939_));
INVX1 INVX1_1701 ( .A(core__abc_22172_new_n6725_), .Y(core__abc_22172_new_n7948_));
INVX1 INVX1_1702 ( .A(core__abc_22172_new_n7949_), .Y(core__abc_22172_new_n7950_));
INVX1 INVX1_1703 ( .A(core__abc_22172_new_n7953_), .Y(core__abc_22172_new_n7954_));
INVX1 INVX1_1704 ( .A(core__abc_22172_new_n7964_), .Y(core__abc_22172_new_n7965_));
INVX1 INVX1_1705 ( .A(core__abc_22172_new_n6703_), .Y(core__abc_22172_new_n7977_));
INVX1 INVX1_1706 ( .A(core__abc_22172_new_n7978_), .Y(core__abc_22172_new_n7979_));
INVX1 INVX1_1707 ( .A(core_key_45_), .Y(core__abc_22172_new_n7984_));
INVX1 INVX1_1708 ( .A(core__abc_22172_new_n7996_), .Y(core__abc_22172_new_n7997_));
INVX1 INVX1_1709 ( .A(core__abc_22172_new_n7998_), .Y(core__abc_22172_new_n7999_));
INVX1 INVX1_171 ( .A(_abc_19873_new_n2798_), .Y(_abc_19873_new_n2799_));
INVX1 INVX1_1710 ( .A(core_key_46_), .Y(core__abc_22172_new_n8001_));
INVX1 INVX1_1711 ( .A(core__abc_22172_new_n6670_), .Y(core__abc_22172_new_n8010_));
INVX1 INVX1_1712 ( .A(core__abc_22172_new_n8011_), .Y(core__abc_22172_new_n8012_));
INVX1 INVX1_1713 ( .A(core__abc_22172_new_n8015_), .Y(core__abc_22172_new_n8016_));
INVX1 INVX1_1714 ( .A(core__abc_22172_new_n6839_), .Y(core__abc_22172_new_n8026_));
INVX1 INVX1_1715 ( .A(core__abc_22172_new_n8029_), .Y(core__abc_22172_new_n8030_));
INVX1 INVX1_1716 ( .A(core_key_48_), .Y(core__abc_22172_new_n8032_));
INVX1 INVX1_1717 ( .A(core__abc_22172_new_n6841_), .Y(core__abc_22172_new_n8041_));
INVX1 INVX1_1718 ( .A(core__abc_22172_new_n8042_), .Y(core__abc_22172_new_n8044_));
INVX1 INVX1_1719 ( .A(core__abc_22172_new_n8058_), .Y(core__abc_22172_new_n8059_));
INVX1 INVX1_172 ( .A(_abc_19873_new_n2803_), .Y(_abc_19873_new_n2804_));
INVX1 INVX1_1720 ( .A(core__abc_22172_new_n6624_), .Y(core__abc_22172_new_n8071_));
INVX1 INVX1_1721 ( .A(core__abc_22172_new_n8073_), .Y(core__abc_22172_new_n8074_));
INVX1 INVX1_1722 ( .A(core_key_51_), .Y(core__abc_22172_new_n8078_));
INVX1 INVX1_1723 ( .A(core__abc_22172_new_n8087_), .Y(core__abc_22172_new_n8088_));
INVX1 INVX1_1724 ( .A(core__abc_22172_new_n8089_), .Y(core__abc_22172_new_n8091_));
INVX1 INVX1_1725 ( .A(core__abc_22172_new_n8093_), .Y(core__abc_22172_new_n8094_));
INVX1 INVX1_1726 ( .A(core_key_52_), .Y(core__abc_22172_new_n8096_));
INVX1 INVX1_1727 ( .A(core__abc_22172_new_n6596_), .Y(core__abc_22172_new_n8105_));
INVX1 INVX1_1728 ( .A(core__abc_22172_new_n8107_), .Y(core__abc_22172_new_n8108_));
INVX1 INVX1_1729 ( .A(core__abc_22172_new_n8110_), .Y(core__abc_22172_new_n8111_));
INVX1 INVX1_173 ( .A(_abc_19873_new_n2808_), .Y(_abc_19873_new_n2809_));
INVX1 INVX1_1730 ( .A(core_key_53_), .Y(core__abc_22172_new_n8113_));
INVX1 INVX1_1731 ( .A(core__abc_22172_new_n8124_), .Y(core__abc_22172_new_n8125_));
INVX1 INVX1_1732 ( .A(core_key_54_), .Y(core__abc_22172_new_n8129_));
INVX1 INVX1_1733 ( .A(core__abc_22172_new_n6578_), .Y(core__abc_22172_new_n8138_));
INVX1 INVX1_1734 ( .A(core__abc_22172_new_n8139_), .Y(core__abc_22172_new_n8140_));
INVX1 INVX1_1735 ( .A(core__abc_22172_new_n8143_), .Y(core__abc_22172_new_n8144_));
INVX1 INVX1_1736 ( .A(core__abc_22172_new_n6849_), .Y(core__abc_22172_new_n8154_));
INVX1 INVX1_1737 ( .A(core__abc_22172_new_n8157_), .Y(core__abc_22172_new_n8158_));
INVX1 INVX1_1738 ( .A(core__abc_22172_new_n6563_), .Y(core__abc_22172_new_n8168_));
INVX1 INVX1_1739 ( .A(core__abc_22172_new_n8156_), .Y(core__abc_22172_new_n8169_));
INVX1 INVX1_174 ( .A(_abc_19873_new_n2813_), .Y(_abc_19873_new_n2814_));
INVX1 INVX1_1740 ( .A(core__abc_22172_new_n8171_), .Y(core__abc_22172_new_n8172_));
INVX1 INVX1_1741 ( .A(core__abc_22172_new_n8186_), .Y(core__abc_22172_new_n8187_));
INVX1 INVX1_1742 ( .A(core_key_58_), .Y(core__abc_22172_new_n8191_));
INVX1 INVX1_1743 ( .A(core__abc_22172_new_n6515_), .Y(core__abc_22172_new_n8200_));
INVX1 INVX1_1744 ( .A(core__abc_22172_new_n8201_), .Y(core__abc_22172_new_n8202_));
INVX1 INVX1_1745 ( .A(core_key_59_), .Y(core__abc_22172_new_n8207_));
INVX1 INVX1_1746 ( .A(core__abc_22172_new_n8216_), .Y(core__abc_22172_new_n8217_));
INVX1 INVX1_1747 ( .A(core__abc_22172_new_n8218_), .Y(core__abc_22172_new_n8219_));
INVX1 INVX1_1748 ( .A(core__abc_22172_new_n8222_), .Y(core__abc_22172_new_n8223_));
INVX1 INVX1_1749 ( .A(core__abc_22172_new_n6495_), .Y(core__abc_22172_new_n8233_));
INVX1 INVX1_175 ( .A(_abc_19873_new_n2818_), .Y(_abc_19873_new_n2819_));
INVX1 INVX1_1750 ( .A(core__abc_22172_new_n8235_), .Y(core__abc_22172_new_n8236_));
INVX1 INVX1_1751 ( .A(core__abc_22172_new_n8238_), .Y(core__abc_22172_new_n8239_));
INVX1 INVX1_1752 ( .A(core_key_61_), .Y(core__abc_22172_new_n8241_));
INVX1 INVX1_1753 ( .A(core__abc_22172_new_n8252_), .Y(core__abc_22172_new_n8253_));
INVX1 INVX1_1754 ( .A(core_key_62_), .Y(core__abc_22172_new_n8257_));
INVX1 INVX1_1755 ( .A(core__abc_22172_new_n6475_), .Y(core__abc_22172_new_n8266_));
INVX1 INVX1_1756 ( .A(core__abc_22172_new_n8269_), .Y(core__abc_22172_new_n8270_));
INVX1 INVX1_1757 ( .A(core__abc_22172_new_n8271_), .Y(core__abc_22172_new_n8272_));
INVX1 INVX1_1758 ( .A(core__abc_22172_new_n8282_), .Y(core__abc_22172_new_n8283_));
INVX1 INVX1_1759 ( .A(core__abc_22172_new_n7806_), .Y(core__abc_22172_new_n8298_));
INVX1 INVX1_176 ( .A(_abc_19873_new_n2823_), .Y(_abc_19873_new_n2824_));
INVX1 INVX1_1760 ( .A(core__abc_22172_new_n8303_), .Y(core__abc_22172_new_n8304_));
INVX1 INVX1_1761 ( .A(core__abc_22172_new_n7814_), .Y(core__abc_22172_new_n8315_));
INVX1 INVX1_1762 ( .A(core_key_66_), .Y(core__abc_22172_new_n8319_));
INVX1 INVX1_1763 ( .A(core_key_67_), .Y(core__abc_22172_new_n8337_));
INVX1 INVX1_1764 ( .A(core__abc_22172_new_n7844_), .Y(core__abc_22172_new_n8348_));
INVX1 INVX1_1765 ( .A(core__abc_22172_new_n7875_), .Y(core__abc_22172_new_n8377_));
INVX1 INVX1_1766 ( .A(core__abc_22172_new_n7891_), .Y(core__abc_22172_new_n8392_));
INVX1 INVX1_1767 ( .A(core__abc_22172_new_n8397_), .Y(core__abc_22172_new_n8398_));
INVX1 INVX1_1768 ( .A(core__abc_22172_new_n7904_), .Y(core__abc_22172_new_n8408_));
INVX1 INVX1_1769 ( .A(core_key_73_), .Y(core__abc_22172_new_n8424_));
INVX1 INVX1_177 ( .A(_abc_19873_new_n2828_), .Y(_abc_19873_new_n2829_));
INVX1 INVX1_1770 ( .A(core__abc_22172_new_n7937_), .Y(core__abc_22172_new_n8433_));
INVX1 INVX1_1771 ( .A(core_key_75_), .Y(core__abc_22172_new_n8449_));
INVX1 INVX1_1772 ( .A(core__abc_22172_new_n7967_), .Y(core__abc_22172_new_n8458_));
INVX1 INVX1_1773 ( .A(core__abc_22172_new_n7982_), .Y(core__abc_22172_new_n8471_));
INVX1 INVX1_1774 ( .A(core__abc_22172_new_n8046_), .Y(core__abc_22172_new_n8515_));
INVX1 INVX1_1775 ( .A(core__abc_22172_new_n8061_), .Y(core__abc_22172_new_n8527_));
INVX1 INVX1_1776 ( .A(core__abc_22172_new_n8076_), .Y(core__abc_22172_new_n8539_));
INVX1 INVX1_1777 ( .A(core__abc_22172_new_n8127_), .Y(core__abc_22172_new_n8574_));
INVX1 INVX1_1778 ( .A(core__abc_22172_new_n6751_), .Y(core__abc_22172_new_n8597_));
INVX1 INVX1_1779 ( .A(core__abc_22172_new_n8174_), .Y(core__abc_22172_new_n8610_));
INVX1 INVX1_178 ( .A(_abc_19873_new_n2833_), .Y(_abc_19873_new_n2834_));
INVX1 INVX1_1780 ( .A(core_key_89_), .Y(core__abc_22172_new_n8615_));
INVX1 INVX1_1781 ( .A(core__abc_22172_new_n8189_), .Y(core__abc_22172_new_n8624_));
INVX1 INVX1_1782 ( .A(core__abc_22172_new_n6733_), .Y(core__abc_22172_new_n8626_));
INVX1 INVX1_1783 ( .A(core_key_90_), .Y(core__abc_22172_new_n8630_));
INVX1 INVX1_1784 ( .A(core__abc_22172_new_n8205_), .Y(core__abc_22172_new_n8639_));
INVX1 INVX1_1785 ( .A(core__abc_22172_new_n8255_), .Y(core__abc_22172_new_n8674_));
INVX1 INVX1_1786 ( .A(core_key_96_), .Y(core__abc_22172_new_n8701_));
INVX1 INVX1_1787 ( .A(core__abc_22172_new_n6929_), .Y(core__abc_22172_new_n8722_));
INVX1 INVX1_1788 ( .A(core__abc_22172_new_n6952_), .Y(core__abc_22172_new_n8734_));
INVX1 INVX1_1789 ( .A(core__abc_22172_new_n6592_), .Y(core__abc_22172_new_n8769_));
INVX1 INVX1_179 ( .A(_abc_19873_new_n2838_), .Y(_abc_19873_new_n2839_));
INVX1 INVX1_1790 ( .A(core__abc_22172_new_n7062_), .Y(core__abc_22172_new_n8780_));
INVX1 INVX1_1791 ( .A(core_key_105_), .Y(core__abc_22172_new_n8807_));
INVX1 INVX1_1792 ( .A(core__abc_22172_new_n7164_), .Y(core__abc_22172_new_n8816_));
INVX1 INVX1_1793 ( .A(core__abc_22172_new_n7188_), .Y(core__abc_22172_new_n8829_));
INVX1 INVX1_1794 ( .A(core_key_108_), .Y(core__abc_22172_new_n8845_));
INVX1 INVX1_1795 ( .A(core__abc_22172_new_n7245_), .Y(core__abc_22172_new_n8854_));
INVX1 INVX1_1796 ( .A(core__abc_22172_new_n6471_), .Y(core__abc_22172_new_n8889_));
INVX1 INVX1_1797 ( .A(core_key_113_), .Y(core__abc_22172_new_n8904_));
INVX1 INVX1_1798 ( .A(core__abc_22172_new_n7433_), .Y(core__abc_22172_new_n8924_));
INVX1 INVX1_1799 ( .A(core_key_115_), .Y(core__abc_22172_new_n8929_));
INVX1 INVX1_18 ( .A(_abc_19873_new_n2141_), .Y(_abc_19873_new_n2142_));
INVX1 INVX1_180 ( .A(_abc_19873_new_n2843_), .Y(_abc_19873_new_n2844_));
INVX1 INVX1_1800 ( .A(core__abc_22172_new_n7495_), .Y(core__abc_22172_new_n8949_));
INVX1 INVX1_1801 ( .A(core__abc_22172_new_n6997_), .Y(core__abc_22172_new_n8962_));
INVX1 INVX1_1802 ( .A(core__abc_22172_new_n7616_), .Y(core__abc_22172_new_n8995_));
INVX1 INVX1_1803 ( .A(core__abc_22172_new_n7646_), .Y(core__abc_22172_new_n9007_));
INVX1 INVX1_1804 ( .A(core__abc_22172_new_n7122_), .Y(core__abc_22172_new_n9009_));
INVX1 INVX1_1805 ( .A(core__abc_22172_new_n7671_), .Y(core__abc_22172_new_n9020_));
INVX1 INVX1_1806 ( .A(core__abc_22172_new_n7179_), .Y(core__abc_22172_new_n9033_));
INVX1 INVX1_1807 ( .A(core__abc_22172_new_n7780_), .Y(core__abc_22172_new_n9067_));
INVX1 INVX1_1808 ( .A(core__abc_22172_new_n9080_), .Y(core__abc_22172_new_n9081_));
INVX1 INVX1_1809 ( .A(core__abc_22172_new_n9087_), .Y(core__abc_22172_new_n9088_));
INVX1 INVX1_181 ( .A(_abc_19873_new_n2848_), .Y(_abc_19873_new_n2849_));
INVX1 INVX1_1810 ( .A(core__abc_22172_new_n9098_), .Y(core__abc_22172_new_n9099_));
INVX1 INVX1_1811 ( .A(core_key_2_), .Y(core__abc_22172_new_n9109_));
INVX1 INVX1_1812 ( .A(core__abc_22172_new_n9112_), .Y(core__abc_22172_new_n9113_));
INVX1 INVX1_1813 ( .A(core__abc_22172_new_n9125_), .Y(core__abc_22172_new_n9126_));
INVX1 INVX1_1814 ( .A(core_key_4_), .Y(core__abc_22172_new_n9135_));
INVX1 INVX1_1815 ( .A(core__abc_22172_new_n9138_), .Y(core__abc_22172_new_n9139_));
INVX1 INVX1_1816 ( .A(core__abc_22172_new_n9150_), .Y(core__abc_22172_new_n9151_));
INVX1 INVX1_1817 ( .A(core__abc_22172_new_n9162_), .Y(core__abc_22172_new_n9163_));
INVX1 INVX1_1818 ( .A(core__abc_22172_new_n9174_), .Y(core__abc_22172_new_n9175_));
INVX1 INVX1_1819 ( .A(core_key_8_), .Y(core__abc_22172_new_n9185_));
INVX1 INVX1_182 ( .A(_abc_19873_new_n2853_), .Y(_abc_19873_new_n2854_));
INVX1 INVX1_1820 ( .A(core__abc_22172_new_n9188_), .Y(core__abc_22172_new_n9189_));
INVX1 INVX1_1821 ( .A(core__abc_22172_new_n9201_), .Y(core__abc_22172_new_n9202_));
INVX1 INVX1_1822 ( .A(core_key_10_), .Y(core__abc_22172_new_n9212_));
INVX1 INVX1_1823 ( .A(core__abc_22172_new_n9215_), .Y(core__abc_22172_new_n9216_));
INVX1 INVX1_1824 ( .A(core__abc_22172_new_n9227_), .Y(core__abc_22172_new_n9228_));
INVX1 INVX1_1825 ( .A(core__abc_22172_new_n9240_), .Y(core__abc_22172_new_n9241_));
INVX1 INVX1_1826 ( .A(core__abc_22172_new_n9252_), .Y(core__abc_22172_new_n9253_));
INVX1 INVX1_1827 ( .A(core__abc_22172_new_n9264_), .Y(core__abc_22172_new_n9265_));
INVX1 INVX1_1828 ( .A(core__abc_22172_new_n9276_), .Y(core__abc_22172_new_n9277_));
INVX1 INVX1_1829 ( .A(core__abc_22172_new_n9288_), .Y(core__abc_22172_new_n9289_));
INVX1 INVX1_183 ( .A(_abc_19873_new_n2858_), .Y(_abc_19873_new_n2859_));
INVX1 INVX1_1830 ( .A(core_key_17_), .Y(core__abc_22172_new_n9299_));
INVX1 INVX1_1831 ( .A(core__abc_22172_new_n9302_), .Y(core__abc_22172_new_n9303_));
INVX1 INVX1_1832 ( .A(core__abc_22172_new_n9315_), .Y(core__abc_22172_new_n9316_));
INVX1 INVX1_1833 ( .A(core__abc_22172_new_n9327_), .Y(core__abc_22172_new_n9328_));
INVX1 INVX1_1834 ( .A(core_key_20_), .Y(core__abc_22172_new_n9338_));
INVX1 INVX1_1835 ( .A(core__abc_22172_new_n9341_), .Y(core__abc_22172_new_n9342_));
INVX1 INVX1_1836 ( .A(core__abc_22172_new_n9353_), .Y(core__abc_22172_new_n9354_));
INVX1 INVX1_1837 ( .A(core__abc_22172_new_n9365_), .Y(core__abc_22172_new_n9366_));
INVX1 INVX1_1838 ( .A(core__abc_22172_new_n9377_), .Y(core__abc_22172_new_n9378_));
INVX1 INVX1_1839 ( .A(core__abc_22172_new_n9389_), .Y(core__abc_22172_new_n9390_));
INVX1 INVX1_184 ( .A(_abc_19873_new_n2863_), .Y(_abc_19873_new_n2864_));
INVX1 INVX1_1840 ( .A(core__abc_22172_new_n9402_), .Y(core__abc_22172_new_n9403_));
INVX1 INVX1_1841 ( .A(core__abc_22172_new_n9415_), .Y(core__abc_22172_new_n9416_));
INVX1 INVX1_1842 ( .A(core__abc_22172_new_n9428_), .Y(core__abc_22172_new_n9429_));
INVX1 INVX1_1843 ( .A(core_key_28_), .Y(core__abc_22172_new_n9439_));
INVX1 INVX1_1844 ( .A(core__abc_22172_new_n9442_), .Y(core__abc_22172_new_n9443_));
INVX1 INVX1_1845 ( .A(core__abc_22172_new_n9454_), .Y(core__abc_22172_new_n9455_));
INVX1 INVX1_1846 ( .A(core__abc_22172_new_n9466_), .Y(core__abc_22172_new_n9467_));
INVX1 INVX1_1847 ( .A(core__abc_22172_new_n9478_), .Y(core__abc_22172_new_n9479_));
INVX1 INVX1_1848 ( .A(core__abc_22172_new_n9490_), .Y(core__abc_22172_new_n9491_));
INVX1 INVX1_1849 ( .A(core__abc_22172_new_n9502_), .Y(core__abc_22172_new_n9503_));
INVX1 INVX1_185 ( .A(_abc_19873_new_n2868_), .Y(_abc_19873_new_n2869_));
INVX1 INVX1_1850 ( .A(core__abc_22172_new_n9514_), .Y(core__abc_22172_new_n9515_));
INVX1 INVX1_1851 ( .A(core__abc_22172_new_n9526_), .Y(core__abc_22172_new_n9527_));
INVX1 INVX1_1852 ( .A(core__abc_22172_new_n9538_), .Y(core__abc_22172_new_n9539_));
INVX1 INVX1_1853 ( .A(core__abc_22172_new_n9550_), .Y(core__abc_22172_new_n9551_));
INVX1 INVX1_1854 ( .A(core__abc_22172_new_n9562_), .Y(core__abc_22172_new_n9563_));
INVX1 INVX1_1855 ( .A(core__abc_22172_new_n9574_), .Y(core__abc_22172_new_n9575_));
INVX1 INVX1_1856 ( .A(core__abc_22172_new_n9586_), .Y(core__abc_22172_new_n9587_));
INVX1 INVX1_1857 ( .A(core__abc_22172_new_n9599_), .Y(core__abc_22172_new_n9600_));
INVX1 INVX1_1858 ( .A(core__abc_22172_new_n9611_), .Y(core__abc_22172_new_n9612_));
INVX1 INVX1_1859 ( .A(core_key_43_), .Y(core__abc_22172_new_n9622_));
INVX1 INVX1_186 ( .A(_abc_19873_new_n2873_), .Y(_abc_19873_new_n2874_));
INVX1 INVX1_1860 ( .A(core__abc_22172_new_n9625_), .Y(core__abc_22172_new_n9626_));
INVX1 INVX1_1861 ( .A(core__abc_22172_new_n9637_), .Y(core__abc_22172_new_n9638_));
INVX1 INVX1_1862 ( .A(core__abc_22172_new_n9649_), .Y(core__abc_22172_new_n9650_));
INVX1 INVX1_1863 ( .A(core__abc_22172_new_n9661_), .Y(core__abc_22172_new_n9662_));
INVX1 INVX1_1864 ( .A(core__abc_22172_new_n9673_), .Y(core__abc_22172_new_n9674_));
INVX1 INVX1_1865 ( .A(core__abc_22172_new_n9685_), .Y(core__abc_22172_new_n9686_));
INVX1 INVX1_1866 ( .A(core_key_49_), .Y(core__abc_22172_new_n9696_));
INVX1 INVX1_1867 ( .A(core__abc_22172_new_n9699_), .Y(core__abc_22172_new_n9700_));
INVX1 INVX1_1868 ( .A(core_key_50_), .Y(core__abc_22172_new_n9710_));
INVX1 INVX1_1869 ( .A(core__abc_22172_new_n9713_), .Y(core__abc_22172_new_n9714_));
INVX1 INVX1_187 ( .A(_abc_19873_new_n2878_), .Y(_abc_19873_new_n2879_));
INVX1 INVX1_1870 ( .A(core__abc_22172_new_n9725_), .Y(core__abc_22172_new_n9726_));
INVX1 INVX1_1871 ( .A(core__abc_22172_new_n9738_), .Y(core__abc_22172_new_n9739_));
INVX1 INVX1_1872 ( .A(core__abc_22172_new_n9750_), .Y(core__abc_22172_new_n9751_));
INVX1 INVX1_1873 ( .A(core__abc_22172_new_n9762_), .Y(core__abc_22172_new_n9763_));
INVX1 INVX1_1874 ( .A(core__abc_22172_new_n9774_), .Y(core__abc_22172_new_n9775_));
INVX1 INVX1_1875 ( .A(core_key_56_), .Y(core__abc_22172_new_n9785_));
INVX1 INVX1_1876 ( .A(core__abc_22172_new_n9788_), .Y(core__abc_22172_new_n9789_));
INVX1 INVX1_1877 ( .A(core_key_57_), .Y(core__abc_22172_new_n9799_));
INVX1 INVX1_1878 ( .A(core__abc_22172_new_n9802_), .Y(core__abc_22172_new_n9803_));
INVX1 INVX1_1879 ( .A(core__abc_22172_new_n9815_), .Y(core__abc_22172_new_n9816_));
INVX1 INVX1_188 ( .A(_abc_19873_new_n2883_), .Y(_abc_19873_new_n2884_));
INVX1 INVX1_1880 ( .A(core__abc_22172_new_n9828_), .Y(core__abc_22172_new_n9829_));
INVX1 INVX1_1881 ( .A(core_key_60_), .Y(core__abc_22172_new_n9839_));
INVX1 INVX1_1882 ( .A(core__abc_22172_new_n9842_), .Y(core__abc_22172_new_n9843_));
INVX1 INVX1_1883 ( .A(core__abc_22172_new_n9854_), .Y(core__abc_22172_new_n9855_));
INVX1 INVX1_1884 ( .A(core__abc_22172_new_n9866_), .Y(core__abc_22172_new_n9867_));
INVX1 INVX1_1885 ( .A(core__abc_22172_new_n9878_), .Y(core__abc_22172_new_n9879_));
INVX1 INVX1_1886 ( .A(core__abc_22172_new_n2659_), .Y(core__abc_22172_new_n9895_));
INVX1 INVX1_189 ( .A(_abc_19873_new_n2888_), .Y(_abc_19873_new_n2889_));
INVX1 INVX1_19 ( .A(\write_data[4] ), .Y(_abc_19873_new_n2146_));
INVX1 INVX1_190 ( .A(_abc_19873_new_n2893_), .Y(_abc_19873_new_n2894_));
INVX1 INVX1_191 ( .A(_abc_19873_new_n2898_), .Y(_abc_19873_new_n2899_));
INVX1 INVX1_192 ( .A(_abc_19873_new_n2903_), .Y(_abc_19873_new_n2904_));
INVX1 INVX1_193 ( .A(_abc_19873_new_n2908_), .Y(_abc_19873_new_n2909_));
INVX1 INVX1_194 ( .A(_abc_19873_new_n2913_), .Y(_abc_19873_new_n2914_));
INVX1 INVX1_195 ( .A(_abc_19873_new_n2918_), .Y(_abc_19873_new_n2919_));
INVX1 INVX1_196 ( .A(_abc_19873_new_n2923_), .Y(_abc_19873_new_n2924_));
INVX1 INVX1_197 ( .A(_abc_19873_new_n2928_), .Y(_abc_19873_new_n2929_));
INVX1 INVX1_198 ( .A(_abc_19873_new_n2933_), .Y(_abc_19873_new_n2934_));
INVX1 INVX1_199 ( .A(_abc_19873_new_n2938_), .Y(_abc_19873_new_n2939_));
INVX1 INVX1_2 ( .A(\addr[6] ), .Y(_abc_19873_new_n871_));
INVX1 INVX1_20 ( .A(_abc_19873_new_n2147_), .Y(_abc_19873_new_n2148_));
INVX1 INVX1_200 ( .A(_abc_19873_new_n2943_), .Y(_abc_19873_new_n2944_));
INVX1 INVX1_201 ( .A(_abc_19873_new_n2948_), .Y(_abc_19873_new_n2949_));
INVX1 INVX1_202 ( .A(_abc_19873_new_n2953_), .Y(_abc_19873_new_n2954_));
INVX1 INVX1_203 ( .A(_abc_19873_new_n2959_), .Y(_abc_19873_new_n2960_));
INVX1 INVX1_204 ( .A(_abc_19873_new_n2964_), .Y(_abc_19873_new_n2965_));
INVX1 INVX1_205 ( .A(_abc_19873_new_n2969_), .Y(_abc_19873_new_n2970_));
INVX1 INVX1_206 ( .A(_abc_19873_new_n2974_), .Y(_abc_19873_new_n2975_));
INVX1 INVX1_207 ( .A(_abc_19873_new_n2979_), .Y(_abc_19873_new_n2980_));
INVX1 INVX1_208 ( .A(_abc_19873_new_n2984_), .Y(_abc_19873_new_n2985_));
INVX1 INVX1_209 ( .A(_abc_19873_new_n2989_), .Y(_abc_19873_new_n2990_));
INVX1 INVX1_21 ( .A(\write_data[5] ), .Y(_abc_19873_new_n2152_));
INVX1 INVX1_210 ( .A(_abc_19873_new_n2994_), .Y(_abc_19873_new_n2995_));
INVX1 INVX1_211 ( .A(_abc_19873_new_n2999_), .Y(_abc_19873_new_n3000_));
INVX1 INVX1_212 ( .A(_abc_19873_new_n3004_), .Y(_abc_19873_new_n3005_));
INVX1 INVX1_213 ( .A(_abc_19873_new_n3009_), .Y(_abc_19873_new_n3010_));
INVX1 INVX1_214 ( .A(_abc_19873_new_n3014_), .Y(_abc_19873_new_n3015_));
INVX1 INVX1_215 ( .A(_abc_19873_new_n3019_), .Y(_abc_19873_new_n3020_));
INVX1 INVX1_216 ( .A(_abc_19873_new_n3024_), .Y(_abc_19873_new_n3025_));
INVX1 INVX1_217 ( .A(_abc_19873_new_n3029_), .Y(_abc_19873_new_n3030_));
INVX1 INVX1_218 ( .A(_abc_19873_new_n3034_), .Y(_abc_19873_new_n3035_));
INVX1 INVX1_219 ( .A(_abc_19873_new_n3039_), .Y(_abc_19873_new_n3040_));
INVX1 INVX1_22 ( .A(_abc_19873_new_n2153_), .Y(_abc_19873_new_n2154_));
INVX1 INVX1_220 ( .A(_abc_19873_new_n3044_), .Y(_abc_19873_new_n3045_));
INVX1 INVX1_221 ( .A(_abc_19873_new_n3049_), .Y(_abc_19873_new_n3050_));
INVX1 INVX1_222 ( .A(_abc_19873_new_n3054_), .Y(_abc_19873_new_n3055_));
INVX1 INVX1_223 ( .A(_abc_19873_new_n3059_), .Y(_abc_19873_new_n3060_));
INVX1 INVX1_224 ( .A(_abc_19873_new_n3064_), .Y(_abc_19873_new_n3065_));
INVX1 INVX1_225 ( .A(_abc_19873_new_n3069_), .Y(_abc_19873_new_n3070_));
INVX1 INVX1_226 ( .A(_abc_19873_new_n3074_), .Y(_abc_19873_new_n3075_));
INVX1 INVX1_227 ( .A(_abc_19873_new_n3079_), .Y(_abc_19873_new_n3080_));
INVX1 INVX1_228 ( .A(_abc_19873_new_n3084_), .Y(_abc_19873_new_n3085_));
INVX1 INVX1_229 ( .A(_abc_19873_new_n3089_), .Y(_abc_19873_new_n3090_));
INVX1 INVX1_23 ( .A(\write_data[6] ), .Y(_abc_19873_new_n2158_));
INVX1 INVX1_230 ( .A(_abc_19873_new_n3094_), .Y(_abc_19873_new_n3095_));
INVX1 INVX1_231 ( .A(_abc_19873_new_n3099_), .Y(_abc_19873_new_n3100_));
INVX1 INVX1_232 ( .A(_abc_19873_new_n3104_), .Y(_abc_19873_new_n3105_));
INVX1 INVX1_233 ( .A(_abc_19873_new_n3109_), .Y(_abc_19873_new_n3110_));
INVX1 INVX1_234 ( .A(_abc_19873_new_n3114_), .Y(_abc_19873_new_n3115_));
INVX1 INVX1_235 ( .A(_abc_19873_new_n3118_), .Y(_abc_19873_new_n3120_));
INVX1 INVX1_236 ( .A(reset_n), .Y(_abc_19873_new_n3125_));
INVX1 INVX1_237 ( .A(_abc_19873_new_n3163_), .Y(_abc_19873_new_n3164_));
INVX1 INVX1_238 ( .A(core_final_rounds_3_), .Y(core__abc_22172_new_n1130_));
INVX1 INVX1_239 ( .A(core_final_rounds_2_), .Y(core__abc_22172_new_n1131_));
INVX1 INVX1_24 ( .A(_abc_19873_new_n2159_), .Y(_abc_19873_new_n2160_));
INVX1 INVX1_240 ( .A(core_final_rounds_1_), .Y(core__abc_22172_new_n1132_));
INVX1 INVX1_241 ( .A(core_final_rounds_0_), .Y(core__abc_22172_new_n1133_));
INVX1 INVX1_242 ( .A(core__abc_22172_new_n1135_), .Y(core__abc_22172_new_n1137_));
INVX1 INVX1_243 ( .A(core__abc_22172_new_n1139_), .Y(core__abc_22172_new_n1140_));
INVX1 INVX1_244 ( .A(core_loop_ctr_reg_3_), .Y(core__abc_22172_new_n1142_));
INVX1 INVX1_245 ( .A(core__abc_22172_new_n1144_), .Y(core__abc_22172_new_n1145_));
INVX1 INVX1_246 ( .A(core__abc_22172_new_n1148_), .Y(core__abc_22172_new_n1149_));
INVX1 INVX1_247 ( .A(core__abc_22172_new_n1153_), .Y(core__abc_22172_new_n1154_));
INVX1 INVX1_248 ( .A(core_loop_ctr_reg_1_), .Y(core__abc_22172_new_n1155_));
INVX1 INVX1_249 ( .A(core__abc_22172_new_n1159_), .Y(core__abc_22172_new_n1160_));
INVX1 INVX1_25 ( .A(\write_data[7] ), .Y(_abc_19873_new_n2164_));
INVX1 INVX1_250 ( .A(core_siphash_ctrl_reg_5_), .Y(core__abc_22172_new_n1168_));
INVX1 INVX1_251 ( .A(core_siphash_ctrl_reg_2_), .Y(core__abc_22172_new_n1169_));
INVX1 INVX1_252 ( .A(core__abc_22172_new_n1170_), .Y(core__abc_22172_new_n1171_));
INVX1 INVX1_253 ( .A(core__abc_22172_new_n1173_), .Y(core__abc_22172_new_n1174_));
INVX1 INVX1_254 ( .A(core_compression_rounds_3_), .Y(core__abc_22172_new_n1176_));
INVX1 INVX1_255 ( .A(core_compression_rounds_2_), .Y(core__abc_22172_new_n1177_));
INVX1 INVX1_256 ( .A(core_compression_rounds_1_), .Y(core__abc_22172_new_n1178_));
INVX1 INVX1_257 ( .A(core_compression_rounds_0_), .Y(core__abc_22172_new_n1179_));
INVX1 INVX1_258 ( .A(core__abc_22172_new_n1181_), .Y(core__abc_22172_new_n1183_));
INVX1 INVX1_259 ( .A(core__abc_22172_new_n1185_), .Y(core__abc_22172_new_n1186_));
INVX1 INVX1_26 ( .A(_abc_19873_new_n2165_), .Y(_abc_19873_new_n2166_));
INVX1 INVX1_260 ( .A(core__abc_22172_new_n1187_), .Y(core__abc_22172_new_n1188_));
INVX1 INVX1_261 ( .A(core__abc_22172_new_n1190_), .Y(core__abc_22172_new_n1191_));
INVX1 INVX1_262 ( .A(core__abc_22172_new_n1195_), .Y(core__abc_22172_new_n1196_));
INVX1 INVX1_263 ( .A(core__abc_22172_new_n1202_), .Y(core__abc_22172_new_n1203_));
INVX1 INVX1_264 ( .A(core_loop_ctr_reg_2_), .Y(core__abc_22172_new_n1205_));
INVX1 INVX1_265 ( .A(core__abc_22172_new_n1209_), .Y(core__abc_22172_new_n1210_));
INVX1 INVX1_266 ( .A(core_initalize), .Y(core__abc_22172_new_n1213_));
INVX1 INVX1_267 ( .A(core__abc_22172_new_n1217_), .Y(core__abc_22172_new_n1218_));
INVX1 INVX1_268 ( .A(core__abc_22172_new_n1222_), .Y(core__abc_22172_new_n1223_));
INVX1 INVX1_269 ( .A(core__abc_22172_new_n1225_), .Y(core__abc_22172_new_n1226_));
INVX1 INVX1_27 ( .A(\write_data[8] ), .Y(_abc_19873_new_n2170_));
INVX1 INVX1_270 ( .A(core__abc_22172_new_n1211_), .Y(core__abc_22172_new_n1230_));
INVX1 INVX1_271 ( .A(core__abc_22172_new_n1165_), .Y(core__abc_22172_new_n1232_));
INVX1 INVX1_272 ( .A(reset_n), .Y(core__abc_22172_new_n1238_));
INVX1 INVX1_273 ( .A(core__abc_22172_new_n1172_), .Y(core__abc_22172_new_n1239_));
INVX1 INVX1_274 ( .A(core_compress), .Y(core__abc_22172_new_n1252_));
INVX1 INVX1_275 ( .A(core_siphash_word1_we), .Y(core__abc_22172_new_n1256_));
INVX1 INVX1_276 ( .A(core__abc_22172_new_n1258_), .Y(core__abc_22172_new_n1259_));
INVX1 INVX1_277 ( .A(core_v2_reg_0_), .Y(core__abc_22172_new_n1261_));
INVX1 INVX1_278 ( .A(core_v3_reg_0_), .Y(core__abc_22172_new_n1262_));
INVX1 INVX1_279 ( .A(core__abc_22172_new_n1265_), .Y(core__abc_22172_new_n1266_));
INVX1 INVX1_28 ( .A(_abc_19873_new_n2171_), .Y(_abc_19873_new_n2172_));
INVX1 INVX1_280 ( .A(core__abc_22172_new_n1260_), .Y(core__abc_22172_new_n1268_));
INVX1 INVX1_281 ( .A(core__abc_22172_new_n1276_), .Y(core__abc_22172_new_n1277_));
INVX1 INVX1_282 ( .A(core_v2_reg_1_), .Y(core__abc_22172_new_n1280_));
INVX1 INVX1_283 ( .A(core_v3_reg_1_), .Y(core__abc_22172_new_n1281_));
INVX1 INVX1_284 ( .A(core__abc_22172_new_n1283_), .Y(core__abc_22172_new_n1284_));
INVX1 INVX1_285 ( .A(core_v1_reg_1_), .Y(core__abc_22172_new_n1286_));
INVX1 INVX1_286 ( .A(core_v0_reg_1_), .Y(core__abc_22172_new_n1287_));
INVX1 INVX1_287 ( .A(core__abc_22172_new_n1296_), .Y(core__abc_22172_new_n1297_));
INVX1 INVX1_288 ( .A(core__abc_22172_new_n1299_), .Y(core__abc_22172_new_n1300_));
INVX1 INVX1_289 ( .A(core_v2_reg_2_), .Y(core__abc_22172_new_n1302_));
INVX1 INVX1_29 ( .A(\write_data[9] ), .Y(_abc_19873_new_n2176_));
INVX1 INVX1_290 ( .A(core_v3_reg_2_), .Y(core__abc_22172_new_n1303_));
INVX1 INVX1_291 ( .A(core__abc_22172_new_n1305_), .Y(core__abc_22172_new_n1306_));
INVX1 INVX1_292 ( .A(core__abc_22172_new_n1315_), .Y(core__abc_22172_new_n1316_));
INVX1 INVX1_293 ( .A(core_v2_reg_3_), .Y(core__abc_22172_new_n1319_));
INVX1 INVX1_294 ( .A(core_v3_reg_3_), .Y(core__abc_22172_new_n1320_));
INVX1 INVX1_295 ( .A(core__abc_22172_new_n1322_), .Y(core__abc_22172_new_n1323_));
INVX1 INVX1_296 ( .A(core__abc_22172_new_n1317_), .Y(core__abc_22172_new_n1325_));
INVX1 INVX1_297 ( .A(core__abc_22172_new_n1333_), .Y(core__abc_22172_new_n1334_));
INVX1 INVX1_298 ( .A(core_v2_reg_4_), .Y(core__abc_22172_new_n1337_));
INVX1 INVX1_299 ( .A(core_v3_reg_4_), .Y(core__abc_22172_new_n1338_));
INVX1 INVX1_3 ( .A(\addr[5] ), .Y(_abc_19873_new_n873_));
INVX1 INVX1_30 ( .A(_abc_19873_new_n2177_), .Y(_abc_19873_new_n2178_));
INVX1 INVX1_300 ( .A(core__abc_22172_new_n1340_), .Y(core__abc_22172_new_n1341_));
INVX1 INVX1_301 ( .A(core__abc_22172_new_n1335_), .Y(core__abc_22172_new_n1343_));
INVX1 INVX1_302 ( .A(core__abc_22172_new_n1351_), .Y(core__abc_22172_new_n1352_));
INVX1 INVX1_303 ( .A(core__abc_22172_new_n1354_), .Y(core__abc_22172_new_n1355_));
INVX1 INVX1_304 ( .A(core_v2_reg_5_), .Y(core__abc_22172_new_n1356_));
INVX1 INVX1_305 ( .A(core_v3_reg_5_), .Y(core__abc_22172_new_n1357_));
INVX1 INVX1_306 ( .A(core__abc_22172_new_n1358_), .Y(core__abc_22172_new_n1359_));
INVX1 INVX1_307 ( .A(core__abc_22172_new_n1353_), .Y(core__abc_22172_new_n1362_));
INVX1 INVX1_308 ( .A(core__abc_22172_new_n1360_), .Y(core__abc_22172_new_n1363_));
INVX1 INVX1_309 ( .A(core__abc_22172_new_n1371_), .Y(core__abc_22172_new_n1372_));
INVX1 INVX1_31 ( .A(\write_data[10] ), .Y(_abc_19873_new_n2182_));
INVX1 INVX1_310 ( .A(core_v2_reg_6_), .Y(core__abc_22172_new_n1375_));
INVX1 INVX1_311 ( .A(core_v3_reg_6_), .Y(core__abc_22172_new_n1376_));
INVX1 INVX1_312 ( .A(core__abc_22172_new_n1378_), .Y(core__abc_22172_new_n1379_));
INVX1 INVX1_313 ( .A(core__abc_22172_new_n1373_), .Y(core__abc_22172_new_n1381_));
INVX1 INVX1_314 ( .A(core__abc_22172_new_n1389_), .Y(core__abc_22172_new_n1390_));
INVX1 INVX1_315 ( .A(core__abc_22172_new_n1392_), .Y(core__abc_22172_new_n1393_));
INVX1 INVX1_316 ( .A(core_v2_reg_7_), .Y(core__abc_22172_new_n1394_));
INVX1 INVX1_317 ( .A(core_v3_reg_7_), .Y(core__abc_22172_new_n1395_));
INVX1 INVX1_318 ( .A(core__abc_22172_new_n1396_), .Y(core__abc_22172_new_n1397_));
INVX1 INVX1_319 ( .A(core__abc_22172_new_n1391_), .Y(core__abc_22172_new_n1400_));
INVX1 INVX1_32 ( .A(_abc_19873_new_n2183_), .Y(_abc_19873_new_n2184_));
INVX1 INVX1_320 ( .A(core__abc_22172_new_n1398_), .Y(core__abc_22172_new_n1401_));
INVX1 INVX1_321 ( .A(core__abc_22172_new_n1409_), .Y(core__abc_22172_new_n1410_));
INVX1 INVX1_322 ( .A(core__abc_22172_new_n1412_), .Y(core__abc_22172_new_n1413_));
INVX1 INVX1_323 ( .A(core__abc_22172_new_n1411_), .Y(core__abc_22172_new_n1417_));
INVX1 INVX1_324 ( .A(core__abc_22172_new_n1415_), .Y(core__abc_22172_new_n1418_));
INVX1 INVX1_325 ( .A(core__abc_22172_new_n1426_), .Y(core__abc_22172_new_n1427_));
INVX1 INVX1_326 ( .A(core__abc_22172_new_n1429_), .Y(core__abc_22172_new_n1430_));
INVX1 INVX1_327 ( .A(core__abc_22172_new_n1428_), .Y(core__abc_22172_new_n1434_));
INVX1 INVX1_328 ( .A(core__abc_22172_new_n1432_), .Y(core__abc_22172_new_n1435_));
INVX1 INVX1_329 ( .A(core__abc_22172_new_n1443_), .Y(core__abc_22172_new_n1444_));
INVX1 INVX1_33 ( .A(\write_data[11] ), .Y(_abc_19873_new_n2188_));
INVX1 INVX1_330 ( .A(core__abc_22172_new_n1446_), .Y(core__abc_22172_new_n1447_));
INVX1 INVX1_331 ( .A(core__abc_22172_new_n1445_), .Y(core__abc_22172_new_n1451_));
INVX1 INVX1_332 ( .A(core__abc_22172_new_n1449_), .Y(core__abc_22172_new_n1452_));
INVX1 INVX1_333 ( .A(core__abc_22172_new_n1460_), .Y(core__abc_22172_new_n1461_));
INVX1 INVX1_334 ( .A(core__abc_22172_new_n1463_), .Y(core__abc_22172_new_n1464_));
INVX1 INVX1_335 ( .A(core__abc_22172_new_n1462_), .Y(core__abc_22172_new_n1468_));
INVX1 INVX1_336 ( .A(core__abc_22172_new_n1466_), .Y(core__abc_22172_new_n1469_));
INVX1 INVX1_337 ( .A(core__abc_22172_new_n1477_), .Y(core__abc_22172_new_n1478_));
INVX1 INVX1_338 ( .A(core__abc_22172_new_n1480_), .Y(core__abc_22172_new_n1481_));
INVX1 INVX1_339 ( .A(core__abc_22172_new_n1479_), .Y(core__abc_22172_new_n1485_));
INVX1 INVX1_34 ( .A(_abc_19873_new_n2189_), .Y(_abc_19873_new_n2190_));
INVX1 INVX1_340 ( .A(core__abc_22172_new_n1483_), .Y(core__abc_22172_new_n1486_));
INVX1 INVX1_341 ( .A(core__abc_22172_new_n1494_), .Y(core__abc_22172_new_n1495_));
INVX1 INVX1_342 ( .A(core__abc_22172_new_n1497_), .Y(core__abc_22172_new_n1498_));
INVX1 INVX1_343 ( .A(core__abc_22172_new_n1496_), .Y(core__abc_22172_new_n1502_));
INVX1 INVX1_344 ( .A(core__abc_22172_new_n1500_), .Y(core__abc_22172_new_n1503_));
INVX1 INVX1_345 ( .A(core__abc_22172_new_n1511_), .Y(core__abc_22172_new_n1512_));
INVX1 INVX1_346 ( .A(core__abc_22172_new_n1514_), .Y(core__abc_22172_new_n1515_));
INVX1 INVX1_347 ( .A(core__abc_22172_new_n1513_), .Y(core__abc_22172_new_n1519_));
INVX1 INVX1_348 ( .A(core__abc_22172_new_n1517_), .Y(core__abc_22172_new_n1520_));
INVX1 INVX1_349 ( .A(core__abc_22172_new_n1528_), .Y(core__abc_22172_new_n1529_));
INVX1 INVX1_35 ( .A(\write_data[12] ), .Y(_abc_19873_new_n2194_));
INVX1 INVX1_350 ( .A(core__abc_22172_new_n1531_), .Y(core__abc_22172_new_n1532_));
INVX1 INVX1_351 ( .A(core__abc_22172_new_n1530_), .Y(core__abc_22172_new_n1536_));
INVX1 INVX1_352 ( .A(core__abc_22172_new_n1534_), .Y(core__abc_22172_new_n1537_));
INVX1 INVX1_353 ( .A(core__abc_22172_new_n1545_), .Y(core__abc_22172_new_n1546_));
INVX1 INVX1_354 ( .A(core__abc_22172_new_n1548_), .Y(core__abc_22172_new_n1549_));
INVX1 INVX1_355 ( .A(core__abc_22172_new_n1547_), .Y(core__abc_22172_new_n1553_));
INVX1 INVX1_356 ( .A(core__abc_22172_new_n1551_), .Y(core__abc_22172_new_n1554_));
INVX1 INVX1_357 ( .A(core__abc_22172_new_n1562_), .Y(core__abc_22172_new_n1563_));
INVX1 INVX1_358 ( .A(core__abc_22172_new_n1565_), .Y(core__abc_22172_new_n1566_));
INVX1 INVX1_359 ( .A(core__abc_22172_new_n1564_), .Y(core__abc_22172_new_n1570_));
INVX1 INVX1_36 ( .A(_abc_19873_new_n2195_), .Y(_abc_19873_new_n2196_));
INVX1 INVX1_360 ( .A(core__abc_22172_new_n1568_), .Y(core__abc_22172_new_n1571_));
INVX1 INVX1_361 ( .A(core__abc_22172_new_n1579_), .Y(core__abc_22172_new_n1580_));
INVX1 INVX1_362 ( .A(core__abc_22172_new_n1582_), .Y(core__abc_22172_new_n1583_));
INVX1 INVX1_363 ( .A(core__abc_22172_new_n1581_), .Y(core__abc_22172_new_n1587_));
INVX1 INVX1_364 ( .A(core__abc_22172_new_n1585_), .Y(core__abc_22172_new_n1588_));
INVX1 INVX1_365 ( .A(core__abc_22172_new_n1596_), .Y(core__abc_22172_new_n1597_));
INVX1 INVX1_366 ( .A(core__abc_22172_new_n1599_), .Y(core__abc_22172_new_n1600_));
INVX1 INVX1_367 ( .A(core__abc_22172_new_n1598_), .Y(core__abc_22172_new_n1604_));
INVX1 INVX1_368 ( .A(core__abc_22172_new_n1602_), .Y(core__abc_22172_new_n1605_));
INVX1 INVX1_369 ( .A(core__abc_22172_new_n1613_), .Y(core__abc_22172_new_n1614_));
INVX1 INVX1_37 ( .A(\write_data[13] ), .Y(_abc_19873_new_n2200_));
INVX1 INVX1_370 ( .A(core__abc_22172_new_n1616_), .Y(core__abc_22172_new_n1617_));
INVX1 INVX1_371 ( .A(core__abc_22172_new_n1615_), .Y(core__abc_22172_new_n1621_));
INVX1 INVX1_372 ( .A(core__abc_22172_new_n1619_), .Y(core__abc_22172_new_n1622_));
INVX1 INVX1_373 ( .A(core__abc_22172_new_n1630_), .Y(core__abc_22172_new_n1631_));
INVX1 INVX1_374 ( .A(core__abc_22172_new_n1633_), .Y(core__abc_22172_new_n1634_));
INVX1 INVX1_375 ( .A(core__abc_22172_new_n1632_), .Y(core__abc_22172_new_n1638_));
INVX1 INVX1_376 ( .A(core__abc_22172_new_n1636_), .Y(core__abc_22172_new_n1639_));
INVX1 INVX1_377 ( .A(core__abc_22172_new_n1647_), .Y(core__abc_22172_new_n1648_));
INVX1 INVX1_378 ( .A(core__abc_22172_new_n1650_), .Y(core__abc_22172_new_n1651_));
INVX1 INVX1_379 ( .A(core__abc_22172_new_n1649_), .Y(core__abc_22172_new_n1655_));
INVX1 INVX1_38 ( .A(_abc_19873_new_n2201_), .Y(_abc_19873_new_n2202_));
INVX1 INVX1_380 ( .A(core__abc_22172_new_n1653_), .Y(core__abc_22172_new_n1656_));
INVX1 INVX1_381 ( .A(core__abc_22172_new_n1664_), .Y(core__abc_22172_new_n1665_));
INVX1 INVX1_382 ( .A(core__abc_22172_new_n1667_), .Y(core__abc_22172_new_n1668_));
INVX1 INVX1_383 ( .A(core__abc_22172_new_n1666_), .Y(core__abc_22172_new_n1672_));
INVX1 INVX1_384 ( .A(core__abc_22172_new_n1670_), .Y(core__abc_22172_new_n1673_));
INVX1 INVX1_385 ( .A(core__abc_22172_new_n1681_), .Y(core__abc_22172_new_n1682_));
INVX1 INVX1_386 ( .A(core__abc_22172_new_n1684_), .Y(core__abc_22172_new_n1685_));
INVX1 INVX1_387 ( .A(core__abc_22172_new_n1683_), .Y(core__abc_22172_new_n1689_));
INVX1 INVX1_388 ( .A(core__abc_22172_new_n1687_), .Y(core__abc_22172_new_n1690_));
INVX1 INVX1_389 ( .A(core__abc_22172_new_n1698_), .Y(core__abc_22172_new_n1699_));
INVX1 INVX1_39 ( .A(\write_data[14] ), .Y(_abc_19873_new_n2206_));
INVX1 INVX1_390 ( .A(core__abc_22172_new_n1701_), .Y(core__abc_22172_new_n1702_));
INVX1 INVX1_391 ( .A(core__abc_22172_new_n1700_), .Y(core__abc_22172_new_n1706_));
INVX1 INVX1_392 ( .A(core__abc_22172_new_n1704_), .Y(core__abc_22172_new_n1707_));
INVX1 INVX1_393 ( .A(core__abc_22172_new_n1715_), .Y(core__abc_22172_new_n1716_));
INVX1 INVX1_394 ( .A(core__abc_22172_new_n1718_), .Y(core__abc_22172_new_n1719_));
INVX1 INVX1_395 ( .A(core__abc_22172_new_n1717_), .Y(core__abc_22172_new_n1723_));
INVX1 INVX1_396 ( .A(core__abc_22172_new_n1721_), .Y(core__abc_22172_new_n1724_));
INVX1 INVX1_397 ( .A(core__abc_22172_new_n1732_), .Y(core__abc_22172_new_n1733_));
INVX1 INVX1_398 ( .A(core__abc_22172_new_n1735_), .Y(core__abc_22172_new_n1736_));
INVX1 INVX1_399 ( .A(core__abc_22172_new_n1734_), .Y(core__abc_22172_new_n1740_));
INVX1 INVX1_4 ( .A(\addr[3] ), .Y(_abc_19873_new_n877_));
INVX1 INVX1_40 ( .A(_abc_19873_new_n2207_), .Y(_abc_19873_new_n2208_));
INVX1 INVX1_400 ( .A(core__abc_22172_new_n1738_), .Y(core__abc_22172_new_n1741_));
INVX1 INVX1_401 ( .A(core__abc_22172_new_n1749_), .Y(core__abc_22172_new_n1750_));
INVX1 INVX1_402 ( .A(core__abc_22172_new_n1752_), .Y(core__abc_22172_new_n1753_));
INVX1 INVX1_403 ( .A(core__abc_22172_new_n1751_), .Y(core__abc_22172_new_n1757_));
INVX1 INVX1_404 ( .A(core__abc_22172_new_n1755_), .Y(core__abc_22172_new_n1758_));
INVX1 INVX1_405 ( .A(core__abc_22172_new_n1766_), .Y(core__abc_22172_new_n1767_));
INVX1 INVX1_406 ( .A(core__abc_22172_new_n1769_), .Y(core__abc_22172_new_n1770_));
INVX1 INVX1_407 ( .A(core__abc_22172_new_n1768_), .Y(core__abc_22172_new_n1774_));
INVX1 INVX1_408 ( .A(core__abc_22172_new_n1772_), .Y(core__abc_22172_new_n1775_));
INVX1 INVX1_409 ( .A(core__abc_22172_new_n1783_), .Y(core__abc_22172_new_n1784_));
INVX1 INVX1_41 ( .A(\write_data[15] ), .Y(_abc_19873_new_n2212_));
INVX1 INVX1_410 ( .A(core__abc_22172_new_n1786_), .Y(core__abc_22172_new_n1787_));
INVX1 INVX1_411 ( .A(core__abc_22172_new_n1785_), .Y(core__abc_22172_new_n1791_));
INVX1 INVX1_412 ( .A(core__abc_22172_new_n1789_), .Y(core__abc_22172_new_n1792_));
INVX1 INVX1_413 ( .A(core__abc_22172_new_n1800_), .Y(core__abc_22172_new_n1801_));
INVX1 INVX1_414 ( .A(core__abc_22172_new_n1803_), .Y(core__abc_22172_new_n1804_));
INVX1 INVX1_415 ( .A(core__abc_22172_new_n1802_), .Y(core__abc_22172_new_n1808_));
INVX1 INVX1_416 ( .A(core__abc_22172_new_n1806_), .Y(core__abc_22172_new_n1809_));
INVX1 INVX1_417 ( .A(core__abc_22172_new_n1817_), .Y(core__abc_22172_new_n1818_));
INVX1 INVX1_418 ( .A(core__abc_22172_new_n1820_), .Y(core__abc_22172_new_n1821_));
INVX1 INVX1_419 ( .A(core__abc_22172_new_n1819_), .Y(core__abc_22172_new_n1825_));
INVX1 INVX1_42 ( .A(_abc_19873_new_n2213_), .Y(_abc_19873_new_n2214_));
INVX1 INVX1_420 ( .A(core__abc_22172_new_n1823_), .Y(core__abc_22172_new_n1826_));
INVX1 INVX1_421 ( .A(core__abc_22172_new_n1834_), .Y(core__abc_22172_new_n1835_));
INVX1 INVX1_422 ( .A(core__abc_22172_new_n1837_), .Y(core__abc_22172_new_n1838_));
INVX1 INVX1_423 ( .A(core__abc_22172_new_n1836_), .Y(core__abc_22172_new_n1842_));
INVX1 INVX1_424 ( .A(core__abc_22172_new_n1840_), .Y(core__abc_22172_new_n1843_));
INVX1 INVX1_425 ( .A(core__abc_22172_new_n1851_), .Y(core__abc_22172_new_n1852_));
INVX1 INVX1_426 ( .A(core__abc_22172_new_n1855_), .Y(core__abc_22172_new_n1856_));
INVX1 INVX1_427 ( .A(core__abc_22172_new_n1853_), .Y(core__abc_22172_new_n1859_));
INVX1 INVX1_428 ( .A(core__abc_22172_new_n1857_), .Y(core__abc_22172_new_n1860_));
INVX1 INVX1_429 ( .A(core__abc_22172_new_n1868_), .Y(core__abc_22172_new_n1869_));
INVX1 INVX1_43 ( .A(\write_data[16] ), .Y(_abc_19873_new_n2218_));
INVX1 INVX1_430 ( .A(core__abc_22172_new_n1871_), .Y(core__abc_22172_new_n1872_));
INVX1 INVX1_431 ( .A(core__abc_22172_new_n1870_), .Y(core__abc_22172_new_n1876_));
INVX1 INVX1_432 ( .A(core__abc_22172_new_n1874_), .Y(core__abc_22172_new_n1877_));
INVX1 INVX1_433 ( .A(core__abc_22172_new_n1885_), .Y(core__abc_22172_new_n1886_));
INVX1 INVX1_434 ( .A(core__abc_22172_new_n1889_), .Y(core__abc_22172_new_n1890_));
INVX1 INVX1_435 ( .A(core__abc_22172_new_n1887_), .Y(core__abc_22172_new_n1893_));
INVX1 INVX1_436 ( .A(core__abc_22172_new_n1891_), .Y(core__abc_22172_new_n1894_));
INVX1 INVX1_437 ( .A(core__abc_22172_new_n1902_), .Y(core__abc_22172_new_n1903_));
INVX1 INVX1_438 ( .A(core__abc_22172_new_n1905_), .Y(core__abc_22172_new_n1906_));
INVX1 INVX1_439 ( .A(core__abc_22172_new_n1904_), .Y(core__abc_22172_new_n1910_));
INVX1 INVX1_44 ( .A(_abc_19873_new_n2219_), .Y(_abc_19873_new_n2220_));
INVX1 INVX1_440 ( .A(core__abc_22172_new_n1908_), .Y(core__abc_22172_new_n1911_));
INVX1 INVX1_441 ( .A(core__abc_22172_new_n1919_), .Y(core__abc_22172_new_n1920_));
INVX1 INVX1_442 ( .A(core__abc_22172_new_n1923_), .Y(core__abc_22172_new_n1924_));
INVX1 INVX1_443 ( .A(core__abc_22172_new_n1921_), .Y(core__abc_22172_new_n1927_));
INVX1 INVX1_444 ( .A(core__abc_22172_new_n1925_), .Y(core__abc_22172_new_n1928_));
INVX1 INVX1_445 ( .A(core__abc_22172_new_n1936_), .Y(core__abc_22172_new_n1937_));
INVX1 INVX1_446 ( .A(core__abc_22172_new_n1939_), .Y(core__abc_22172_new_n1940_));
INVX1 INVX1_447 ( .A(core__abc_22172_new_n1938_), .Y(core__abc_22172_new_n1944_));
INVX1 INVX1_448 ( .A(core__abc_22172_new_n1942_), .Y(core__abc_22172_new_n1945_));
INVX1 INVX1_449 ( .A(core__abc_22172_new_n1953_), .Y(core__abc_22172_new_n1954_));
INVX1 INVX1_45 ( .A(\write_data[17] ), .Y(_abc_19873_new_n2224_));
INVX1 INVX1_450 ( .A(core__abc_22172_new_n1956_), .Y(core__abc_22172_new_n1957_));
INVX1 INVX1_451 ( .A(core__abc_22172_new_n1955_), .Y(core__abc_22172_new_n1961_));
INVX1 INVX1_452 ( .A(core__abc_22172_new_n1959_), .Y(core__abc_22172_new_n1962_));
INVX1 INVX1_453 ( .A(core__abc_22172_new_n1970_), .Y(core__abc_22172_new_n1971_));
INVX1 INVX1_454 ( .A(core__abc_22172_new_n1973_), .Y(core__abc_22172_new_n1974_));
INVX1 INVX1_455 ( .A(core__abc_22172_new_n1972_), .Y(core__abc_22172_new_n1978_));
INVX1 INVX1_456 ( .A(core__abc_22172_new_n1976_), .Y(core__abc_22172_new_n1979_));
INVX1 INVX1_457 ( .A(core__abc_22172_new_n1987_), .Y(core__abc_22172_new_n1988_));
INVX1 INVX1_458 ( .A(core__abc_22172_new_n1990_), .Y(core__abc_22172_new_n1991_));
INVX1 INVX1_459 ( .A(core__abc_22172_new_n1989_), .Y(core__abc_22172_new_n1995_));
INVX1 INVX1_46 ( .A(_abc_19873_new_n2225_), .Y(_abc_19873_new_n2226_));
INVX1 INVX1_460 ( .A(core__abc_22172_new_n1993_), .Y(core__abc_22172_new_n1996_));
INVX1 INVX1_461 ( .A(core__abc_22172_new_n2004_), .Y(core__abc_22172_new_n2005_));
INVX1 INVX1_462 ( .A(core__abc_22172_new_n2008_), .Y(core__abc_22172_new_n2009_));
INVX1 INVX1_463 ( .A(core__abc_22172_new_n2006_), .Y(core__abc_22172_new_n2012_));
INVX1 INVX1_464 ( .A(core__abc_22172_new_n2010_), .Y(core__abc_22172_new_n2013_));
INVX1 INVX1_465 ( .A(core__abc_22172_new_n2021_), .Y(core__abc_22172_new_n2022_));
INVX1 INVX1_466 ( .A(core__abc_22172_new_n2025_), .Y(core__abc_22172_new_n2026_));
INVX1 INVX1_467 ( .A(core__abc_22172_new_n2023_), .Y(core__abc_22172_new_n2029_));
INVX1 INVX1_468 ( .A(core__abc_22172_new_n2027_), .Y(core__abc_22172_new_n2030_));
INVX1 INVX1_469 ( .A(core__abc_22172_new_n2038_), .Y(core__abc_22172_new_n2039_));
INVX1 INVX1_47 ( .A(\write_data[18] ), .Y(_abc_19873_new_n2230_));
INVX1 INVX1_470 ( .A(core__abc_22172_new_n2042_), .Y(core__abc_22172_new_n2043_));
INVX1 INVX1_471 ( .A(core__abc_22172_new_n2040_), .Y(core__abc_22172_new_n2046_));
INVX1 INVX1_472 ( .A(core__abc_22172_new_n2044_), .Y(core__abc_22172_new_n2047_));
INVX1 INVX1_473 ( .A(core__abc_22172_new_n2055_), .Y(core__abc_22172_new_n2056_));
INVX1 INVX1_474 ( .A(core__abc_22172_new_n2059_), .Y(core__abc_22172_new_n2060_));
INVX1 INVX1_475 ( .A(core__abc_22172_new_n2057_), .Y(core__abc_22172_new_n2063_));
INVX1 INVX1_476 ( .A(core__abc_22172_new_n2061_), .Y(core__abc_22172_new_n2064_));
INVX1 INVX1_477 ( .A(core__abc_22172_new_n2072_), .Y(core__abc_22172_new_n2073_));
INVX1 INVX1_478 ( .A(core__abc_22172_new_n2076_), .Y(core__abc_22172_new_n2077_));
INVX1 INVX1_479 ( .A(core__abc_22172_new_n2074_), .Y(core__abc_22172_new_n2080_));
INVX1 INVX1_48 ( .A(_abc_19873_new_n2231_), .Y(_abc_19873_new_n2232_));
INVX1 INVX1_480 ( .A(core__abc_22172_new_n2078_), .Y(core__abc_22172_new_n2081_));
INVX1 INVX1_481 ( .A(core__abc_22172_new_n2089_), .Y(core__abc_22172_new_n2090_));
INVX1 INVX1_482 ( .A(core__abc_22172_new_n2093_), .Y(core__abc_22172_new_n2094_));
INVX1 INVX1_483 ( .A(core__abc_22172_new_n2091_), .Y(core__abc_22172_new_n2097_));
INVX1 INVX1_484 ( .A(core__abc_22172_new_n2095_), .Y(core__abc_22172_new_n2098_));
INVX1 INVX1_485 ( .A(core__abc_22172_new_n2105_), .Y(core__abc_22172_new_n2106_));
INVX1 INVX1_486 ( .A(core__abc_22172_new_n2108_), .Y(core__abc_22172_new_n2109_));
INVX1 INVX1_487 ( .A(core__abc_22172_new_n2111_), .Y(core__abc_22172_new_n2112_));
INVX1 INVX1_488 ( .A(core__abc_22172_new_n2113_), .Y(core__abc_22172_new_n2115_));
INVX1 INVX1_489 ( .A(core__abc_22172_new_n2123_), .Y(core__abc_22172_new_n2124_));
INVX1 INVX1_49 ( .A(\write_data[19] ), .Y(_abc_19873_new_n2236_));
INVX1 INVX1_490 ( .A(core__abc_22172_new_n2127_), .Y(core__abc_22172_new_n2128_));
INVX1 INVX1_491 ( .A(core__abc_22172_new_n2125_), .Y(core__abc_22172_new_n2131_));
INVX1 INVX1_492 ( .A(core__abc_22172_new_n2129_), .Y(core__abc_22172_new_n2132_));
INVX1 INVX1_493 ( .A(core__abc_22172_new_n2140_), .Y(core__abc_22172_new_n2141_));
INVX1 INVX1_494 ( .A(core__abc_22172_new_n2144_), .Y(core__abc_22172_new_n2145_));
INVX1 INVX1_495 ( .A(core__abc_22172_new_n2142_), .Y(core__abc_22172_new_n2148_));
INVX1 INVX1_496 ( .A(core__abc_22172_new_n2146_), .Y(core__abc_22172_new_n2149_));
INVX1 INVX1_497 ( .A(core__abc_22172_new_n2157_), .Y(core__abc_22172_new_n2158_));
INVX1 INVX1_498 ( .A(core__abc_22172_new_n2161_), .Y(core__abc_22172_new_n2162_));
INVX1 INVX1_499 ( .A(core__abc_22172_new_n2159_), .Y(core__abc_22172_new_n2165_));
INVX1 INVX1_5 ( .A(\addr[2] ), .Y(_abc_19873_new_n878_));
INVX1 INVX1_50 ( .A(_abc_19873_new_n2237_), .Y(_abc_19873_new_n2238_));
INVX1 INVX1_500 ( .A(core__abc_22172_new_n2163_), .Y(core__abc_22172_new_n2166_));
INVX1 INVX1_501 ( .A(core__abc_22172_new_n2173_), .Y(core__abc_22172_new_n2174_));
INVX1 INVX1_502 ( .A(core__abc_22172_new_n2176_), .Y(core__abc_22172_new_n2177_));
INVX1 INVX1_503 ( .A(core__abc_22172_new_n2179_), .Y(core__abc_22172_new_n2180_));
INVX1 INVX1_504 ( .A(core__abc_22172_new_n2181_), .Y(core__abc_22172_new_n2183_));
INVX1 INVX1_505 ( .A(core__abc_22172_new_n2191_), .Y(core__abc_22172_new_n2192_));
INVX1 INVX1_506 ( .A(core__abc_22172_new_n2195_), .Y(core__abc_22172_new_n2196_));
INVX1 INVX1_507 ( .A(core__abc_22172_new_n2193_), .Y(core__abc_22172_new_n2199_));
INVX1 INVX1_508 ( .A(core__abc_22172_new_n2197_), .Y(core__abc_22172_new_n2200_));
INVX1 INVX1_509 ( .A(core__abc_22172_new_n2208_), .Y(core__abc_22172_new_n2209_));
INVX1 INVX1_51 ( .A(\write_data[20] ), .Y(_abc_19873_new_n2242_));
INVX1 INVX1_510 ( .A(core__abc_22172_new_n2212_), .Y(core__abc_22172_new_n2213_));
INVX1 INVX1_511 ( .A(core__abc_22172_new_n2210_), .Y(core__abc_22172_new_n2216_));
INVX1 INVX1_512 ( .A(core__abc_22172_new_n2214_), .Y(core__abc_22172_new_n2217_));
INVX1 INVX1_513 ( .A(core__abc_22172_new_n2225_), .Y(core__abc_22172_new_n2226_));
INVX1 INVX1_514 ( .A(core__abc_22172_new_n2229_), .Y(core__abc_22172_new_n2230_));
INVX1 INVX1_515 ( .A(core__abc_22172_new_n2227_), .Y(core__abc_22172_new_n2233_));
INVX1 INVX1_516 ( .A(core__abc_22172_new_n2231_), .Y(core__abc_22172_new_n2234_));
INVX1 INVX1_517 ( .A(core__abc_22172_new_n2242_), .Y(core__abc_22172_new_n2243_));
INVX1 INVX1_518 ( .A(core__abc_22172_new_n2246_), .Y(core__abc_22172_new_n2247_));
INVX1 INVX1_519 ( .A(core__abc_22172_new_n2244_), .Y(core__abc_22172_new_n2250_));
INVX1 INVX1_52 ( .A(_abc_19873_new_n2243_), .Y(_abc_19873_new_n2244_));
INVX1 INVX1_520 ( .A(core__abc_22172_new_n2248_), .Y(core__abc_22172_new_n2251_));
INVX1 INVX1_521 ( .A(core__abc_22172_new_n2259_), .Y(core__abc_22172_new_n2260_));
INVX1 INVX1_522 ( .A(core__abc_22172_new_n2263_), .Y(core__abc_22172_new_n2264_));
INVX1 INVX1_523 ( .A(core__abc_22172_new_n2261_), .Y(core__abc_22172_new_n2267_));
INVX1 INVX1_524 ( .A(core__abc_22172_new_n2265_), .Y(core__abc_22172_new_n2268_));
INVX1 INVX1_525 ( .A(core__abc_22172_new_n2276_), .Y(core__abc_22172_new_n2277_));
INVX1 INVX1_526 ( .A(core__abc_22172_new_n2280_), .Y(core__abc_22172_new_n2281_));
INVX1 INVX1_527 ( .A(core__abc_22172_new_n2278_), .Y(core__abc_22172_new_n2284_));
INVX1 INVX1_528 ( .A(core__abc_22172_new_n2282_), .Y(core__abc_22172_new_n2285_));
INVX1 INVX1_529 ( .A(core__abc_22172_new_n2293_), .Y(core__abc_22172_new_n2294_));
INVX1 INVX1_53 ( .A(\write_data[21] ), .Y(_abc_19873_new_n2248_));
INVX1 INVX1_530 ( .A(core__abc_22172_new_n2297_), .Y(core__abc_22172_new_n2298_));
INVX1 INVX1_531 ( .A(core__abc_22172_new_n2295_), .Y(core__abc_22172_new_n2301_));
INVX1 INVX1_532 ( .A(core__abc_22172_new_n2299_), .Y(core__abc_22172_new_n2302_));
INVX1 INVX1_533 ( .A(core__abc_22172_new_n2310_), .Y(core__abc_22172_new_n2311_));
INVX1 INVX1_534 ( .A(core__abc_22172_new_n2314_), .Y(core__abc_22172_new_n2315_));
INVX1 INVX1_535 ( .A(core__abc_22172_new_n2312_), .Y(core__abc_22172_new_n2318_));
INVX1 INVX1_536 ( .A(core__abc_22172_new_n2316_), .Y(core__abc_22172_new_n2319_));
INVX1 INVX1_537 ( .A(core__abc_22172_new_n2327_), .Y(core__abc_22172_new_n2328_));
INVX1 INVX1_538 ( .A(core__abc_22172_new_n2331_), .Y(core__abc_22172_new_n2332_));
INVX1 INVX1_539 ( .A(core__abc_22172_new_n2329_), .Y(core__abc_22172_new_n2335_));
INVX1 INVX1_54 ( .A(_abc_19873_new_n2249_), .Y(_abc_19873_new_n2250_));
INVX1 INVX1_540 ( .A(core__abc_22172_new_n2333_), .Y(core__abc_22172_new_n2336_));
INVX1 INVX1_541 ( .A(core_v1_reg_63_), .Y(core__abc_22172_new_n2343_));
INVX1 INVX1_542 ( .A(core_v0_reg_63_), .Y(core__abc_22172_new_n2345_));
INVX1 INVX1_543 ( .A(core__abc_22172_new_n2347_), .Y(core__abc_22172_new_n2348_));
INVX1 INVX1_544 ( .A(core__abc_22172_new_n2350_), .Y(core__abc_22172_new_n2351_));
INVX1 INVX1_545 ( .A(core__abc_22172_new_n2352_), .Y(core__abc_22172_new_n2354_));
INVX1 INVX1_546 ( .A(core_siphash_ctrl_reg_0_), .Y(core__abc_22172_new_n2361_));
INVX1 INVX1_547 ( .A(core__abc_22172_new_n2364_), .Y(core__abc_22172_new_n2366_));
INVX1 INVX1_548 ( .A(core__abc_22172_new_n1216_), .Y(core__abc_22172_new_n2622_));
INVX1 INVX1_549 ( .A(core__abc_22172_new_n2623_), .Y(core__abc_22172_new_n2624_));
INVX1 INVX1_55 ( .A(\write_data[22] ), .Y(_abc_19873_new_n2254_));
INVX1 INVX1_550 ( .A(core__abc_22172_new_n2628_), .Y(core__abc_22172_new_n2629_));
INVX1 INVX1_551 ( .A(core__abc_22172_new_n1220_), .Y(core__abc_22172_new_n2630_));
INVX1 INVX1_552 ( .A(core__abc_22172_new_n2632_), .Y(core__abc_22172_new_n2633_));
INVX1 INVX1_553 ( .A(core__abc_22172_new_n2634_), .Y(core__abc_22172_new_n2635_));
INVX1 INVX1_554 ( .A(core__abc_22172_new_n2640_), .Y(core__abc_22172_new_n2641_));
INVX1 INVX1_555 ( .A(core__abc_22172_new_n2648_), .Y(core__abc_22172_new_n2649_));
INVX1 INVX1_556 ( .A(core__abc_22172_new_n2660_), .Y(core__abc_22172_new_n2662_));
INVX1 INVX1_557 ( .A(core__abc_22172_new_n2948_), .Y(core__abc_22172_new_n2949_));
INVX1 INVX1_558 ( .A(core__abc_22172_new_n2953_), .Y(core__abc_22172_new_n2954_));
INVX1 INVX1_559 ( .A(core__abc_22172_new_n1629_), .Y(core__abc_22172_new_n2984_));
INVX1 INVX1_56 ( .A(_abc_19873_new_n2255_), .Y(_abc_19873_new_n2256_));
INVX1 INVX1_560 ( .A(core__abc_22172_new_n2986_), .Y(core__abc_22172_new_n2987_));
INVX1 INVX1_561 ( .A(core__abc_22172_new_n1697_), .Y(core__abc_22172_new_n2994_));
INVX1 INVX1_562 ( .A(core__abc_22172_new_n2996_), .Y(core__abc_22172_new_n2997_));
INVX1 INVX1_563 ( .A(core__abc_22172_new_n1765_), .Y(core__abc_22172_new_n3005_));
INVX1 INVX1_564 ( .A(core__abc_22172_new_n3007_), .Y(core__abc_22172_new_n3008_));
INVX1 INVX1_565 ( .A(core__abc_22172_new_n2920_), .Y(core__abc_22172_new_n3017_));
INVX1 INVX1_566 ( .A(core__abc_22172_new_n2923_), .Y(core__abc_22172_new_n3019_));
INVX1 INVX1_567 ( .A(core__abc_22172_new_n2927_), .Y(core__abc_22172_new_n3021_));
INVX1 INVX1_568 ( .A(core__abc_22172_new_n2934_), .Y(core__abc_22172_new_n3023_));
INVX1 INVX1_569 ( .A(core__abc_22172_new_n2942_), .Y(core__abc_22172_new_n3025_));
INVX1 INVX1_57 ( .A(\write_data[23] ), .Y(_abc_19873_new_n2260_));
INVX1 INVX1_570 ( .A(core__abc_22172_new_n2959_), .Y(core__abc_22172_new_n3027_));
INVX1 INVX1_571 ( .A(core__abc_22172_new_n2975_), .Y(core__abc_22172_new_n3029_));
INVX1 INVX1_572 ( .A(core__abc_22172_new_n3012_), .Y(core__abc_22172_new_n3031_));
INVX1 INVX1_573 ( .A(core__abc_22172_new_n3035_), .Y(core__abc_22172_new_n3036_));
INVX1 INVX1_574 ( .A(core__abc_22172_new_n3034_), .Y(core__abc_22172_new_n3040_));
INVX1 INVX1_575 ( .A(core__abc_22172_new_n3038_), .Y(core__abc_22172_new_n3041_));
INVX1 INVX1_576 ( .A(core__abc_22172_new_n3043_), .Y(core__abc_22172_new_n3044_));
INVX1 INVX1_577 ( .A(core__abc_22172_new_n1975_), .Y(core__abc_22172_new_n3045_));
INVX1 INVX1_578 ( .A(core__abc_22172_new_n3047_), .Y(core__abc_22172_new_n3048_));
INVX1 INVX1_579 ( .A(core__abc_22172_new_n3050_), .Y(core__abc_22172_new_n3051_));
INVX1 INVX1_58 ( .A(_abc_19873_new_n2261_), .Y(_abc_19873_new_n2262_));
INVX1 INVX1_580 ( .A(core__abc_22172_new_n1279_), .Y(core__abc_22172_new_n3052_));
INVX1 INVX1_581 ( .A(core__abc_22172_new_n1264_), .Y(core__abc_22172_new_n3053_));
INVX1 INVX1_582 ( .A(core__abc_22172_new_n3056_), .Y(core__abc_22172_new_n3057_));
INVX1 INVX1_583 ( .A(core__abc_22172_new_n3059_), .Y(core__abc_22172_new_n3060_));
INVX1 INVX1_584 ( .A(core__abc_22172_new_n1336_), .Y(core__abc_22172_new_n3065_));
INVX1 INVX1_585 ( .A(core__abc_22172_new_n3067_), .Y(core__abc_22172_new_n3068_));
INVX1 INVX1_586 ( .A(core__abc_22172_new_n1431_), .Y(core__abc_22172_new_n3082_));
INVX1 INVX1_587 ( .A(core__abc_22172_new_n3084_), .Y(core__abc_22172_new_n3085_));
INVX1 INVX1_588 ( .A(core__abc_22172_new_n3092_), .Y(core__abc_22172_new_n3093_));
INVX1 INVX1_589 ( .A(core__abc_22172_new_n3117_), .Y(core__abc_22172_new_n3118_));
INVX1 INVX1_59 ( .A(\write_data[24] ), .Y(_abc_19873_new_n2266_));
INVX1 INVX1_590 ( .A(core__abc_22172_new_n1635_), .Y(core__abc_22172_new_n3124_));
INVX1 INVX1_591 ( .A(core__abc_22172_new_n3126_), .Y(core__abc_22172_new_n3127_));
INVX1 INVX1_592 ( .A(core__abc_22172_new_n1703_), .Y(core__abc_22172_new_n3134_));
INVX1 INVX1_593 ( .A(core__abc_22172_new_n3136_), .Y(core__abc_22172_new_n3137_));
INVX1 INVX1_594 ( .A(core__abc_22172_new_n1771_), .Y(core__abc_22172_new_n3145_));
INVX1 INVX1_595 ( .A(core__abc_22172_new_n3147_), .Y(core__abc_22172_new_n3148_));
INVX1 INVX1_596 ( .A(core__abc_22172_new_n1839_), .Y(core__abc_22172_new_n3162_));
INVX1 INVX1_597 ( .A(core__abc_22172_new_n3164_), .Y(core__abc_22172_new_n3165_));
INVX1 INVX1_598 ( .A(core__abc_22172_new_n1907_), .Y(core__abc_22172_new_n3173_));
INVX1 INVX1_599 ( .A(core__abc_22172_new_n3175_), .Y(core__abc_22172_new_n3176_));
INVX1 INVX1_6 ( .A(\addr[0] ), .Y(_abc_19873_new_n883_));
INVX1 INVX1_60 ( .A(_abc_19873_new_n2267_), .Y(_abc_19873_new_n2268_));
INVX1 INVX1_600 ( .A(core__abc_22172_new_n3185_), .Y(core__abc_22172_new_n3186_));
INVX1 INVX1_601 ( .A(core__abc_22172_new_n3190_), .Y(core__abc_22172_new_n3191_));
INVX1 INVX1_602 ( .A(core__abc_22172_new_n3193_), .Y(core__abc_22172_new_n3194_));
INVX1 INVX1_603 ( .A(core__abc_22172_new_n3196_), .Y(core__abc_22172_new_n3197_));
INVX1 INVX1_604 ( .A(core__abc_22172_new_n3198_), .Y(core__abc_22172_new_n3199_));
INVX1 INVX1_605 ( .A(core__abc_22172_new_n3200_), .Y(core__abc_22172_new_n3201_));
INVX1 INVX1_606 ( .A(core__abc_22172_new_n3203_), .Y(core__abc_22172_new_n3204_));
INVX1 INVX1_607 ( .A(core__abc_22172_new_n3214_), .Y(core__abc_22172_new_n3215_));
INVX1 INVX1_608 ( .A(core_key_64_), .Y(core__abc_22172_new_n3218_));
INVX1 INVX1_609 ( .A(core__abc_22172_new_n3220_), .Y(core__abc_22172_new_n3221_));
INVX1 INVX1_61 ( .A(\write_data[25] ), .Y(_abc_19873_new_n2272_));
INVX1 INVX1_610 ( .A(core__abc_22172_new_n3217_), .Y(core__abc_22172_new_n3228_));
INVX1 INVX1_611 ( .A(core__abc_22172_new_n3014_), .Y(core__abc_22172_new_n3232_));
INVX1 INVX1_612 ( .A(core_v3_reg_49_), .Y(core__abc_22172_new_n3240_));
INVX1 INVX1_613 ( .A(core__abc_22172_new_n3054_), .Y(core__abc_22172_new_n3241_));
INVX1 INVX1_614 ( .A(core__abc_22172_new_n3243_), .Y(core__abc_22172_new_n3244_));
INVX1 INVX1_615 ( .A(core__abc_22172_new_n3248_), .Y(core__abc_22172_new_n3249_));
INVX1 INVX1_616 ( .A(core__abc_22172_new_n3252_), .Y(core__abc_22172_new_n3253_));
INVX1 INVX1_617 ( .A(core_v3_reg_28_), .Y(core__abc_22172_new_n3256_));
INVX1 INVX1_618 ( .A(core__abc_22172_new_n3264_), .Y(core__abc_22172_new_n3265_));
INVX1 INVX1_619 ( .A(core__abc_22172_new_n3268_), .Y(core__abc_22172_new_n3269_));
INVX1 INVX1_62 ( .A(_abc_19873_new_n2273_), .Y(_abc_19873_new_n2274_));
INVX1 INVX1_620 ( .A(core__abc_22172_new_n3272_), .Y(core__abc_22172_new_n3273_));
INVX1 INVX1_621 ( .A(core__abc_22172_new_n3255_), .Y(core__abc_22172_new_n3275_));
INVX1 INVX1_622 ( .A(core_key_65_), .Y(core__abc_22172_new_n3279_));
INVX1 INVX1_623 ( .A(core__abc_22172_new_n3281_), .Y(core__abc_22172_new_n3282_));
INVX1 INVX1_624 ( .A(core__abc_22172_new_n3250_), .Y(core__abc_22172_new_n3292_));
INVX1 INVX1_625 ( .A(core__abc_22172_new_n3235_), .Y(core__abc_22172_new_n3294_));
INVX1 INVX1_626 ( .A(core__abc_22172_new_n3295_), .Y(core__abc_22172_new_n3296_));
INVX1 INVX1_627 ( .A(core__abc_22172_new_n3298_), .Y(core__abc_22172_new_n3299_));
INVX1 INVX1_628 ( .A(core__abc_22172_new_n3301_), .Y(core__abc_22172_new_n3302_));
INVX1 INVX1_629 ( .A(core_v3_reg_50_), .Y(core__abc_22172_new_n3303_));
INVX1 INVX1_63 ( .A(\write_data[26] ), .Y(_abc_19873_new_n2278_));
INVX1 INVX1_630 ( .A(core__abc_22172_new_n3055_), .Y(core__abc_22172_new_n3304_));
INVX1 INVX1_631 ( .A(core__abc_22172_new_n3307_), .Y(core__abc_22172_new_n3308_));
INVX1 INVX1_632 ( .A(core__abc_22172_new_n3311_), .Y(core__abc_22172_new_n3313_));
INVX1 INVX1_633 ( .A(core__abc_22172_new_n3315_), .Y(core__abc_22172_new_n3316_));
INVX1 INVX1_634 ( .A(core__abc_22172_new_n3317_), .Y(core__abc_22172_new_n3318_));
INVX1 INVX1_635 ( .A(core__abc_22172_new_n3321_), .Y(core__abc_22172_new_n3322_));
INVX1 INVX1_636 ( .A(core__abc_22172_new_n3326_), .Y(core__abc_22172_new_n3327_));
INVX1 INVX1_637 ( .A(core__abc_22172_new_n3329_), .Y(core__abc_22172_new_n3330_));
INVX1 INVX1_638 ( .A(core__abc_22172_new_n3320_), .Y(core__abc_22172_new_n3332_));
INVX1 INVX1_639 ( .A(core__abc_22172_new_n3337_), .Y(core__abc_22172_new_n3338_));
INVX1 INVX1_64 ( .A(_abc_19873_new_n2279_), .Y(_abc_19873_new_n2280_));
INVX1 INVX1_640 ( .A(core__abc_22172_new_n2041_), .Y(core__abc_22172_new_n3350_));
INVX1 INVX1_641 ( .A(core__abc_22172_new_n3352_), .Y(core__abc_22172_new_n3353_));
INVX1 INVX1_642 ( .A(core__abc_22172_new_n3354_), .Y(core__abc_22172_new_n3356_));
INVX1 INVX1_643 ( .A(core__abc_22172_new_n3358_), .Y(core__abc_22172_new_n3359_));
INVX1 INVX1_644 ( .A(core_v3_reg_30_), .Y(core__abc_22172_new_n3361_));
INVX1 INVX1_645 ( .A(core__abc_22172_new_n3366_), .Y(core__abc_22172_new_n3367_));
INVX1 INVX1_646 ( .A(core__abc_22172_new_n1301_), .Y(core__abc_22172_new_n3370_));
INVX1 INVX1_647 ( .A(core__abc_22172_new_n3305_), .Y(core__abc_22172_new_n3371_));
INVX1 INVX1_648 ( .A(core__abc_22172_new_n3372_), .Y(core__abc_22172_new_n3373_));
INVX1 INVX1_649 ( .A(core__abc_22172_new_n3377_), .Y(core__abc_22172_new_n3378_));
INVX1 INVX1_65 ( .A(\write_data[27] ), .Y(_abc_19873_new_n2284_));
INVX1 INVX1_650 ( .A(core__abc_22172_new_n3381_), .Y(core__abc_22172_new_n3382_));
INVX1 INVX1_651 ( .A(core__abc_22172_new_n3369_), .Y(core__abc_22172_new_n3383_));
INVX1 INVX1_652 ( .A(core__abc_22172_new_n3380_), .Y(core__abc_22172_new_n3384_));
INVX1 INVX1_653 ( .A(core__abc_22172_new_n3385_), .Y(core__abc_22172_new_n3386_));
INVX1 INVX1_654 ( .A(core__abc_22172_new_n3387_), .Y(core__abc_22172_new_n3388_));
INVX1 INVX1_655 ( .A(core__abc_22172_new_n3364_), .Y(core__abc_22172_new_n3390_));
INVX1 INVX1_656 ( .A(core__abc_22172_new_n3392_), .Y(core__abc_22172_new_n3393_));
INVX1 INVX1_657 ( .A(core__abc_22172_new_n3363_), .Y(core__abc_22172_new_n3395_));
INVX1 INVX1_658 ( .A(core__abc_22172_new_n3400_), .Y(core__abc_22172_new_n3401_));
INVX1 INVX1_659 ( .A(core__abc_22172_new_n3418_), .Y(core__abc_22172_new_n3420_));
INVX1 INVX1_66 ( .A(_abc_19873_new_n2285_), .Y(_abc_19873_new_n2286_));
INVX1 INVX1_660 ( .A(core_v3_reg_52_), .Y(core__abc_22172_new_n3423_));
INVX1 INVX1_661 ( .A(core__abc_22172_new_n3426_), .Y(core__abc_22172_new_n3428_));
INVX1 INVX1_662 ( .A(core__abc_22172_new_n3422_), .Y(core__abc_22172_new_n3432_));
INVX1 INVX1_663 ( .A(core__abc_22172_new_n3430_), .Y(core__abc_22172_new_n3433_));
INVX1 INVX1_664 ( .A(core__abc_22172_new_n3435_), .Y(core__abc_22172_new_n3436_));
INVX1 INVX1_665 ( .A(core__abc_22172_new_n3439_), .Y(core__abc_22172_new_n3440_));
INVX1 INVX1_666 ( .A(core__abc_22172_new_n3443_), .Y(core__abc_22172_new_n3444_));
INVX1 INVX1_667 ( .A(core_v3_reg_31_), .Y(core__abc_22172_new_n3449_));
INVX1 INVX1_668 ( .A(core__abc_22172_new_n3447_), .Y(core__abc_22172_new_n3450_));
INVX1 INVX1_669 ( .A(core__abc_22172_new_n3442_), .Y(core__abc_22172_new_n3454_));
INVX1 INVX1_67 ( .A(\write_data[28] ), .Y(_abc_19873_new_n2290_));
INVX1 INVX1_670 ( .A(core__abc_22172_new_n3448_), .Y(core__abc_22172_new_n3455_));
INVX1 INVX1_671 ( .A(core_key_68_), .Y(core__abc_22172_new_n3461_));
INVX1 INVX1_672 ( .A(core__abc_22172_new_n3463_), .Y(core__abc_22172_new_n3464_));
INVX1 INVX1_673 ( .A(core__abc_22172_new_n3474_), .Y(core__abc_22172_new_n3475_));
INVX1 INVX1_674 ( .A(core__abc_22172_new_n3478_), .Y(core__abc_22172_new_n3479_));
INVX1 INVX1_675 ( .A(core_v3_reg_53_), .Y(core__abc_22172_new_n3481_));
INVX1 INVX1_676 ( .A(core__abc_22172_new_n3482_), .Y(core__abc_22172_new_n3483_));
INVX1 INVX1_677 ( .A(core__abc_22172_new_n3486_), .Y(core__abc_22172_new_n3488_));
INVX1 INVX1_678 ( .A(core__abc_22172_new_n3490_), .Y(core__abc_22172_new_n3491_));
INVX1 INVX1_679 ( .A(core__abc_22172_new_n3492_), .Y(core__abc_22172_new_n3493_));
INVX1 INVX1_68 ( .A(_abc_19873_new_n2291_), .Y(_abc_19873_new_n2292_));
INVX1 INVX1_680 ( .A(core__abc_22172_new_n3495_), .Y(core__abc_22172_new_n3497_));
INVX1 INVX1_681 ( .A(core__abc_22172_new_n3499_), .Y(core__abc_22172_new_n3500_));
INVX1 INVX1_682 ( .A(core_v3_reg_32_), .Y(core__abc_22172_new_n3501_));
INVX1 INVX1_683 ( .A(core__abc_22172_new_n3511_), .Y(core__abc_22172_new_n3512_));
INVX1 INVX1_684 ( .A(core__abc_22172_new_n3515_), .Y(core__abc_22172_new_n3516_));
INVX1 INVX1_685 ( .A(core__abc_22172_new_n3519_), .Y(core__abc_22172_new_n3520_));
INVX1 INVX1_686 ( .A(core_key_69_), .Y(core__abc_22172_new_n3525_));
INVX1 INVX1_687 ( .A(core__abc_22172_new_n3527_), .Y(core__abc_22172_new_n3528_));
INVX1 INVX1_688 ( .A(core__abc_22172_new_n1901_), .Y(core__abc_22172_new_n3538_));
INVX1 INVX1_689 ( .A(core__abc_22172_new_n3540_), .Y(core__abc_22172_new_n3541_));
INVX1 INVX1_69 ( .A(\write_data[29] ), .Y(_abc_19873_new_n2296_));
INVX1 INVX1_690 ( .A(core__abc_22172_new_n3544_), .Y(core__abc_22172_new_n3546_));
INVX1 INVX1_691 ( .A(core_v3_reg_54_), .Y(core__abc_22172_new_n3549_));
INVX1 INVX1_692 ( .A(core__abc_22172_new_n3062_), .Y(core__abc_22172_new_n3550_));
INVX1 INVX1_693 ( .A(core__abc_22172_new_n3552_), .Y(core__abc_22172_new_n3553_));
INVX1 INVX1_694 ( .A(core__abc_22172_new_n3556_), .Y(core__abc_22172_new_n3557_));
INVX1 INVX1_695 ( .A(core__abc_22172_new_n3548_), .Y(core__abc_22172_new_n3562_));
INVX1 INVX1_696 ( .A(core__abc_22172_new_n3560_), .Y(core__abc_22172_new_n3563_));
INVX1 INVX1_697 ( .A(core__abc_22172_new_n3565_), .Y(core__abc_22172_new_n3566_));
INVX1 INVX1_698 ( .A(core__abc_22172_new_n3568_), .Y(core__abc_22172_new_n3570_));
INVX1 INVX1_699 ( .A(core__abc_22172_new_n3572_), .Y(core__abc_22172_new_n3573_));
INVX1 INVX1_7 ( .A(\addr[1] ), .Y(_abc_19873_new_n884_));
INVX1 INVX1_70 ( .A(_abc_19873_new_n2297_), .Y(_abc_19873_new_n2298_));
INVX1 INVX1_700 ( .A(core_v3_reg_33_), .Y(core__abc_22172_new_n3574_));
INVX1 INVX1_701 ( .A(core__abc_22172_new_n3514_), .Y(core__abc_22172_new_n3575_));
INVX1 INVX1_702 ( .A(core__abc_22172_new_n3582_), .Y(core__abc_22172_new_n3584_));
INVX1 INVX1_703 ( .A(core__abc_22172_new_n3586_), .Y(core__abc_22172_new_n3587_));
INVX1 INVX1_704 ( .A(core_key_70_), .Y(core__abc_22172_new_n3592_));
INVX1 INVX1_705 ( .A(core__abc_22172_new_n3594_), .Y(core__abc_22172_new_n3595_));
INVX1 INVX1_706 ( .A(core__abc_22172_new_n3605_), .Y(core__abc_22172_new_n3606_));
INVX1 INVX1_707 ( .A(core__abc_22172_new_n3609_), .Y(core__abc_22172_new_n3610_));
INVX1 INVX1_708 ( .A(core_v3_reg_55_), .Y(core__abc_22172_new_n3611_));
INVX1 INVX1_709 ( .A(core__abc_22172_new_n3612_), .Y(core__abc_22172_new_n3613_));
INVX1 INVX1_71 ( .A(\write_data[30] ), .Y(_abc_19873_new_n2302_));
INVX1 INVX1_710 ( .A(core__abc_22172_new_n3616_), .Y(core__abc_22172_new_n3618_));
INVX1 INVX1_711 ( .A(core__abc_22172_new_n3620_), .Y(core__abc_22172_new_n3621_));
INVX1 INVX1_712 ( .A(core__abc_22172_new_n3624_), .Y(core__abc_22172_new_n3625_));
INVX1 INVX1_713 ( .A(core__abc_22172_new_n3626_), .Y(core__abc_22172_new_n3627_));
INVX1 INVX1_714 ( .A(core__abc_22172_new_n3630_), .Y(core__abc_22172_new_n3631_));
INVX1 INVX1_715 ( .A(core_v3_reg_34_), .Y(core__abc_22172_new_n3632_));
INVX1 INVX1_716 ( .A(core__abc_22172_new_n3634_), .Y(core__abc_22172_new_n3635_));
INVX1 INVX1_717 ( .A(core__abc_22172_new_n3638_), .Y(core__abc_22172_new_n3639_));
INVX1 INVX1_718 ( .A(core__abc_22172_new_n3642_), .Y(core__abc_22172_new_n3643_));
INVX1 INVX1_719 ( .A(core__abc_22172_new_n3649_), .Y(core__abc_22172_new_n3650_));
INVX1 INVX1_72 ( .A(_abc_19873_new_n2303_), .Y(_abc_19873_new_n2304_));
INVX1 INVX1_720 ( .A(core__abc_22172_new_n3623_), .Y(core__abc_22172_new_n3664_));
INVX1 INVX1_721 ( .A(core__abc_22172_new_n3671_), .Y(core__abc_22172_new_n3672_));
INVX1 INVX1_722 ( .A(core__abc_22172_new_n3683_), .Y(core__abc_22172_new_n3685_));
INVX1 INVX1_723 ( .A(core__abc_22172_new_n3687_), .Y(core__abc_22172_new_n3688_));
INVX1 INVX1_724 ( .A(core_v3_reg_56_), .Y(core__abc_22172_new_n3689_));
INVX1 INVX1_725 ( .A(core__abc_22172_new_n3073_), .Y(core__abc_22172_new_n3690_));
INVX1 INVX1_726 ( .A(core__abc_22172_new_n3693_), .Y(core__abc_22172_new_n3694_));
INVX1 INVX1_727 ( .A(core__abc_22172_new_n3697_), .Y(core__abc_22172_new_n3698_));
INVX1 INVX1_728 ( .A(core__abc_22172_new_n3701_), .Y(core__abc_22172_new_n3703_));
INVX1 INVX1_729 ( .A(core__abc_22172_new_n3705_), .Y(core__abc_22172_new_n3706_));
INVX1 INVX1_73 ( .A(\write_data[31] ), .Y(_abc_19873_new_n2308_));
INVX1 INVX1_730 ( .A(core__abc_22172_new_n3709_), .Y(core__abc_22172_new_n3710_));
INVX1 INVX1_731 ( .A(core__abc_22172_new_n3711_), .Y(core__abc_22172_new_n3712_));
INVX1 INVX1_732 ( .A(core__abc_22172_new_n3713_), .Y(core__abc_22172_new_n3714_));
INVX1 INVX1_733 ( .A(core__abc_22172_new_n3716_), .Y(core__abc_22172_new_n3717_));
INVX1 INVX1_734 ( .A(core_key_72_), .Y(core__abc_22172_new_n3722_));
INVX1 INVX1_735 ( .A(core__abc_22172_new_n3724_), .Y(core__abc_22172_new_n3725_));
INVX1 INVX1_736 ( .A(core__abc_22172_new_n3704_), .Y(core__abc_22172_new_n3735_));
INVX1 INVX1_737 ( .A(core__abc_22172_new_n3699_), .Y(core__abc_22172_new_n3736_));
INVX1 INVX1_738 ( .A(core__abc_22172_new_n3684_), .Y(core__abc_22172_new_n3737_));
INVX1 INVX1_739 ( .A(core__abc_22172_new_n3739_), .Y(core__abc_22172_new_n3740_));
INVX1 INVX1_74 ( .A(_abc_19873_new_n2309_), .Y(_abc_19873_new_n2310_));
INVX1 INVX1_740 ( .A(core_v3_reg_57_), .Y(core__abc_22172_new_n3743_));
INVX1 INVX1_741 ( .A(core__abc_22172_new_n3744_), .Y(core__abc_22172_new_n3745_));
INVX1 INVX1_742 ( .A(core__abc_22172_new_n3748_), .Y(core__abc_22172_new_n3750_));
INVX1 INVX1_743 ( .A(core__abc_22172_new_n3752_), .Y(core__abc_22172_new_n3753_));
INVX1 INVX1_744 ( .A(core__abc_22172_new_n3754_), .Y(core__abc_22172_new_n3755_));
INVX1 INVX1_745 ( .A(core__abc_22172_new_n3757_), .Y(core__abc_22172_new_n3758_));
INVX1 INVX1_746 ( .A(core__abc_22172_new_n3760_), .Y(core__abc_22172_new_n3761_));
INVX1 INVX1_747 ( .A(core__abc_22172_new_n3762_), .Y(core__abc_22172_new_n3763_));
INVX1 INVX1_748 ( .A(core__abc_22172_new_n3765_), .Y(core__abc_22172_new_n3766_));
INVX1 INVX1_749 ( .A(core_v3_reg_36_), .Y(core__abc_22172_new_n3769_));
INVX1 INVX1_75 ( .A(_abc_19873_new_n2315_), .Y(_abc_19873_new_n2316_));
INVX1 INVX1_750 ( .A(core__abc_22172_new_n3777_), .Y(core__abc_22172_new_n3778_));
INVX1 INVX1_751 ( .A(core__abc_22172_new_n3781_), .Y(core__abc_22172_new_n3782_));
INVX1 INVX1_752 ( .A(core__abc_22172_new_n3785_), .Y(core__abc_22172_new_n3786_));
INVX1 INVX1_753 ( .A(core__abc_22172_new_n3768_), .Y(core__abc_22172_new_n3788_));
INVX1 INVX1_754 ( .A(core__abc_22172_new_n3793_), .Y(core__abc_22172_new_n3794_));
INVX1 INVX1_755 ( .A(core__abc_22172_new_n3804_), .Y(core__abc_22172_new_n3805_));
INVX1 INVX1_756 ( .A(core__abc_22172_new_n3806_), .Y(core__abc_22172_new_n3807_));
INVX1 INVX1_757 ( .A(core__abc_22172_new_n1969_), .Y(core__abc_22172_new_n3810_));
INVX1 INVX1_758 ( .A(core__abc_22172_new_n3812_), .Y(core__abc_22172_new_n3813_));
INVX1 INVX1_759 ( .A(core__abc_22172_new_n3814_), .Y(core__abc_22172_new_n3816_));
INVX1 INVX1_76 ( .A(_abc_19873_new_n2320_), .Y(_abc_19873_new_n2321_));
INVX1 INVX1_760 ( .A(core_v3_reg_58_), .Y(core__abc_22172_new_n3819_));
INVX1 INVX1_761 ( .A(core__abc_22172_new_n3820_), .Y(core__abc_22172_new_n3821_));
INVX1 INVX1_762 ( .A(core__abc_22172_new_n3824_), .Y(core__abc_22172_new_n3825_));
INVX1 INVX1_763 ( .A(core__abc_22172_new_n3826_), .Y(core__abc_22172_new_n3827_));
INVX1 INVX1_764 ( .A(core__abc_22172_new_n3818_), .Y(core__abc_22172_new_n3832_));
INVX1 INVX1_765 ( .A(core__abc_22172_new_n3830_), .Y(core__abc_22172_new_n3833_));
INVX1 INVX1_766 ( .A(core__abc_22172_new_n3835_), .Y(core__abc_22172_new_n3836_));
INVX1 INVX1_767 ( .A(core__abc_22172_new_n3839_), .Y(core__abc_22172_new_n3840_));
INVX1 INVX1_768 ( .A(core__abc_22172_new_n3841_), .Y(core__abc_22172_new_n3842_));
INVX1 INVX1_769 ( .A(core__abc_22172_new_n3847_), .Y(core__abc_22172_new_n3848_));
INVX1 INVX1_77 ( .A(_abc_19873_new_n2325_), .Y(_abc_19873_new_n2326_));
INVX1 INVX1_770 ( .A(core__abc_22172_new_n3849_), .Y(core__abc_22172_new_n3850_));
INVX1 INVX1_771 ( .A(core_key_74_), .Y(core__abc_22172_new_n3855_));
INVX1 INVX1_772 ( .A(core__abc_22172_new_n3857_), .Y(core__abc_22172_new_n3858_));
INVX1 INVX1_773 ( .A(core__abc_22172_new_n3868_), .Y(core__abc_22172_new_n3869_));
INVX1 INVX1_774 ( .A(core__abc_22172_new_n3870_), .Y(core__abc_22172_new_n3871_));
INVX1 INVX1_775 ( .A(core__abc_22172_new_n3874_), .Y(core__abc_22172_new_n3875_));
INVX1 INVX1_776 ( .A(core__abc_22172_new_n3877_), .Y(core__abc_22172_new_n3878_));
INVX1 INVX1_777 ( .A(core__abc_22172_new_n3880_), .Y(core__abc_22172_new_n3881_));
INVX1 INVX1_778 ( .A(core__abc_22172_new_n3882_), .Y(core__abc_22172_new_n3883_));
INVX1 INVX1_779 ( .A(core__abc_22172_new_n3885_), .Y(core__abc_22172_new_n3886_));
INVX1 INVX1_78 ( .A(_abc_19873_new_n2330_), .Y(_abc_19873_new_n2331_));
INVX1 INVX1_780 ( .A(core__abc_22172_new_n3889_), .Y(core__abc_22172_new_n3890_));
INVX1 INVX1_781 ( .A(core__abc_22172_new_n3893_), .Y(core__abc_22172_new_n3894_));
INVX1 INVX1_782 ( .A(core_v3_reg_38_), .Y(core__abc_22172_new_n3895_));
INVX1 INVX1_783 ( .A(core__abc_22172_new_n3900_), .Y(core__abc_22172_new_n3902_));
INVX1 INVX1_784 ( .A(core__abc_22172_new_n3904_), .Y(core__abc_22172_new_n3905_));
INVX1 INVX1_785 ( .A(core__abc_22172_new_n3908_), .Y(core__abc_22172_new_n3909_));
INVX1 INVX1_786 ( .A(core__abc_22172_new_n3915_), .Y(core__abc_22172_new_n3916_));
INVX1 INVX1_787 ( .A(core__abc_22172_new_n3888_), .Y(core__abc_22172_new_n3928_));
INVX1 INVX1_788 ( .A(core__abc_22172_new_n3942_), .Y(core__abc_22172_new_n3944_));
INVX1 INVX1_789 ( .A(core_v3_reg_60_), .Y(core__abc_22172_new_n3947_));
INVX1 INVX1_79 ( .A(_abc_19873_new_n2335_), .Y(_abc_19873_new_n2336_));
INVX1 INVX1_790 ( .A(core__abc_22172_new_n3949_), .Y(core__abc_22172_new_n3951_));
INVX1 INVX1_791 ( .A(core__abc_22172_new_n3953_), .Y(core__abc_22172_new_n3954_));
INVX1 INVX1_792 ( .A(core__abc_22172_new_n3946_), .Y(core__abc_22172_new_n3959_));
INVX1 INVX1_793 ( .A(core__abc_22172_new_n3957_), .Y(core__abc_22172_new_n3960_));
INVX1 INVX1_794 ( .A(core__abc_22172_new_n3962_), .Y(core__abc_22172_new_n3963_));
INVX1 INVX1_795 ( .A(core__abc_22172_new_n3964_), .Y(core__abc_22172_new_n3965_));
INVX1 INVX1_796 ( .A(core__abc_22172_new_n3968_), .Y(core__abc_22172_new_n3969_));
INVX1 INVX1_797 ( .A(core__abc_22172_new_n3974_), .Y(core__abc_22172_new_n3975_));
INVX1 INVX1_798 ( .A(core__abc_22172_new_n3967_), .Y(core__abc_22172_new_n3978_));
INVX1 INVX1_799 ( .A(core__abc_22172_new_n3973_), .Y(core__abc_22172_new_n3979_));
INVX1 INVX1_8 ( .A(\addr[4] ), .Y(_abc_19873_new_n891_));
INVX1 INVX1_80 ( .A(_abc_19873_new_n2340_), .Y(_abc_19873_new_n2341_));
INVX1 INVX1_800 ( .A(core__abc_22172_new_n3985_), .Y(core__abc_22172_new_n3986_));
INVX1 INVX1_801 ( .A(core__abc_22172_new_n3961_), .Y(core__abc_22172_new_n3996_));
INVX1 INVX1_802 ( .A(core__abc_22172_new_n3997_), .Y(core__abc_22172_new_n3998_));
INVX1 INVX1_803 ( .A(core__abc_22172_new_n4001_), .Y(core__abc_22172_new_n4002_));
INVX1 INVX1_804 ( .A(core_v3_reg_61_), .Y(core__abc_22172_new_n4003_));
INVX1 INVX1_805 ( .A(core__abc_22172_new_n4004_), .Y(core__abc_22172_new_n4005_));
INVX1 INVX1_806 ( .A(core__abc_22172_new_n4008_), .Y(core__abc_22172_new_n4010_));
INVX1 INVX1_807 ( .A(core__abc_22172_new_n4012_), .Y(core__abc_22172_new_n4013_));
INVX1 INVX1_808 ( .A(core__abc_22172_new_n4016_), .Y(core__abc_22172_new_n4017_));
INVX1 INVX1_809 ( .A(core__abc_22172_new_n4019_), .Y(core__abc_22172_new_n4020_));
INVX1 INVX1_81 ( .A(_abc_19873_new_n2345_), .Y(_abc_19873_new_n2346_));
INVX1 INVX1_810 ( .A(core__abc_22172_new_n4021_), .Y(core__abc_22172_new_n4022_));
INVX1 INVX1_811 ( .A(core__abc_22172_new_n4024_), .Y(core__abc_22172_new_n4025_));
INVX1 INVX1_812 ( .A(core__abc_22172_new_n4027_), .Y(core__abc_22172_new_n4028_));
INVX1 INVX1_813 ( .A(core__abc_22172_new_n4035_), .Y(core__abc_22172_new_n4037_));
INVX1 INVX1_814 ( .A(core__abc_22172_new_n4039_), .Y(core__abc_22172_new_n4040_));
INVX1 INVX1_815 ( .A(core_v3_reg_40_), .Y(core__abc_22172_new_n4042_));
INVX1 INVX1_816 ( .A(core__abc_22172_new_n4044_), .Y(core__abc_22172_new_n4045_));
INVX1 INVX1_817 ( .A(core_key_77_), .Y(core__abc_22172_new_n4050_));
INVX1 INVX1_818 ( .A(core__abc_22172_new_n4052_), .Y(core__abc_22172_new_n4053_));
INVX1 INVX1_819 ( .A(core__abc_22172_new_n4015_), .Y(core__abc_22172_new_n4063_));
INVX1 INVX1_82 ( .A(_abc_19873_new_n2350_), .Y(_abc_19873_new_n2351_));
INVX1 INVX1_820 ( .A(core__abc_22172_new_n4064_), .Y(core__abc_22172_new_n4065_));
INVX1 INVX1_821 ( .A(core__abc_22172_new_n4066_), .Y(core__abc_22172_new_n4067_));
INVX1 INVX1_822 ( .A(core__abc_22172_new_n2037_), .Y(core__abc_22172_new_n4068_));
INVX1 INVX1_823 ( .A(core__abc_22172_new_n4070_), .Y(core__abc_22172_new_n4071_));
INVX1 INVX1_824 ( .A(core__abc_22172_new_n4074_), .Y(core__abc_22172_new_n4076_));
INVX1 INVX1_825 ( .A(core_v3_reg_62_), .Y(core__abc_22172_new_n4079_));
INVX1 INVX1_826 ( .A(core__abc_22172_new_n4081_), .Y(core__abc_22172_new_n4082_));
INVX1 INVX1_827 ( .A(core__abc_22172_new_n4085_), .Y(core__abc_22172_new_n4086_));
INVX1 INVX1_828 ( .A(core__abc_22172_new_n4090_), .Y(core__abc_22172_new_n4091_));
INVX1 INVX1_829 ( .A(core__abc_22172_new_n4093_), .Y(core__abc_22172_new_n4095_));
INVX1 INVX1_83 ( .A(_abc_19873_new_n2355_), .Y(_abc_19873_new_n2356_));
INVX1 INVX1_830 ( .A(core__abc_22172_new_n4097_), .Y(core__abc_22172_new_n4098_));
INVX1 INVX1_831 ( .A(core__abc_22172_new_n4099_), .Y(core__abc_22172_new_n4100_));
INVX1 INVX1_832 ( .A(core__abc_22172_new_n4103_), .Y(core__abc_22172_new_n4104_));
INVX1 INVX1_833 ( .A(core_v3_reg_41_), .Y(core__abc_22172_new_n4106_));
INVX1 INVX1_834 ( .A(core__abc_22172_new_n4108_), .Y(core__abc_22172_new_n4109_));
INVX1 INVX1_835 ( .A(core_key_78_), .Y(core__abc_22172_new_n4114_));
INVX1 INVX1_836 ( .A(core__abc_22172_new_n4116_), .Y(core__abc_22172_new_n4117_));
INVX1 INVX1_837 ( .A(core__abc_22172_new_n4092_), .Y(core__abc_22172_new_n4127_));
INVX1 INVX1_838 ( .A(core__abc_22172_new_n4128_), .Y(core__abc_22172_new_n4129_));
INVX1 INVX1_839 ( .A(core__abc_22172_new_n4132_), .Y(core__abc_22172_new_n4133_));
INVX1 INVX1_84 ( .A(_abc_19873_new_n2360_), .Y(_abc_19873_new_n2361_));
INVX1 INVX1_840 ( .A(core__abc_22172_new_n4135_), .Y(core__abc_22172_new_n4136_));
INVX1 INVX1_841 ( .A(core__abc_22172_new_n4140_), .Y(core__abc_22172_new_n4141_));
INVX1 INVX1_842 ( .A(core__abc_22172_new_n4143_), .Y(core__abc_22172_new_n4144_));
INVX1 INVX1_843 ( .A(core__abc_22172_new_n4131_), .Y(core__abc_22172_new_n4146_));
INVX1 INVX1_844 ( .A(core__abc_22172_new_n4149_), .Y(core__abc_22172_new_n4150_));
INVX1 INVX1_845 ( .A(core__abc_22172_new_n4153_), .Y(core__abc_22172_new_n4154_));
INVX1 INVX1_846 ( .A(core_v3_reg_42_), .Y(core__abc_22172_new_n4155_));
INVX1 INVX1_847 ( .A(core__abc_22172_new_n4160_), .Y(core__abc_22172_new_n4161_));
INVX1 INVX1_848 ( .A(core__abc_22172_new_n4164_), .Y(core__abc_22172_new_n4165_));
INVX1 INVX1_849 ( .A(core__abc_22172_new_n4168_), .Y(core__abc_22172_new_n4169_));
INVX1 INVX1_85 ( .A(_abc_19873_new_n2365_), .Y(_abc_19873_new_n2366_));
INVX1 INVX1_850 ( .A(core__abc_22172_new_n4175_), .Y(core__abc_22172_new_n4176_));
INVX1 INVX1_851 ( .A(core__abc_22172_new_n3212_), .Y(core__abc_22172_new_n4187_));
INVX1 INVX1_852 ( .A(core__abc_22172_new_n4148_), .Y(core__abc_22172_new_n4194_));
INVX1 INVX1_853 ( .A(core__abc_22172_new_n4210_), .Y(core__abc_22172_new_n4215_));
INVX1 INVX1_854 ( .A(core__abc_22172_new_n4211_), .Y(core__abc_22172_new_n4216_));
INVX1 INVX1_855 ( .A(core__abc_22172_new_n3099_), .Y(core__abc_22172_new_n4221_));
INVX1 INVX1_856 ( .A(core__abc_22172_new_n4224_), .Y(core__abc_22172_new_n4225_));
INVX1 INVX1_857 ( .A(core__abc_22172_new_n4228_), .Y(core__abc_22172_new_n4229_));
INVX1 INVX1_858 ( .A(core__abc_22172_new_n4220_), .Y(core__abc_22172_new_n4231_));
INVX1 INVX1_859 ( .A(core__abc_22172_new_n4233_), .Y(core__abc_22172_new_n4234_));
INVX1 INVX1_86 ( .A(_abc_19873_new_n2370_), .Y(_abc_19873_new_n2371_));
INVX1 INVX1_860 ( .A(core__abc_22172_new_n4199_), .Y(core__abc_22172_new_n4236_));
INVX1 INVX1_861 ( .A(core__abc_22172_new_n4238_), .Y(core__abc_22172_new_n4239_));
INVX1 INVX1_862 ( .A(core__abc_22172_new_n4163_), .Y(core__abc_22172_new_n4240_));
INVX1 INVX1_863 ( .A(core__abc_22172_new_n4243_), .Y(core__abc_22172_new_n4244_));
INVX1 INVX1_864 ( .A(core_v3_reg_43_), .Y(core__abc_22172_new_n4247_));
INVX1 INVX1_865 ( .A(core__abc_22172_new_n4242_), .Y(core__abc_22172_new_n4248_));
INVX1 INVX1_866 ( .A(core__abc_22172_new_n4250_), .Y(core__abc_22172_new_n4254_));
INVX1 INVX1_867 ( .A(core__abc_22172_new_n4261_), .Y(core__abc_22172_new_n4262_));
INVX1 INVX1_868 ( .A(core__abc_22172_new_n4235_), .Y(core__abc_22172_new_n4270_));
INVX1 INVX1_869 ( .A(core__abc_22172_new_n4232_), .Y(core__abc_22172_new_n4271_));
INVX1 INVX1_87 ( .A(_abc_19873_new_n2375_), .Y(_abc_19873_new_n2376_));
INVX1 INVX1_870 ( .A(core__abc_22172_new_n4214_), .Y(core__abc_22172_new_n4272_));
INVX1 INVX1_871 ( .A(core__abc_22172_new_n4274_), .Y(core__abc_22172_new_n4275_));
INVX1 INVX1_872 ( .A(core__abc_22172_new_n4276_), .Y(core__abc_22172_new_n4277_));
INVX1 INVX1_873 ( .A(core__abc_22172_new_n4278_), .Y(core__abc_22172_new_n4279_));
INVX1 INVX1_874 ( .A(core__abc_22172_new_n4283_), .Y(core__abc_22172_new_n4284_));
INVX1 INVX1_875 ( .A(core__abc_22172_new_n4287_), .Y(core__abc_22172_new_n4289_));
INVX1 INVX1_876 ( .A(core__abc_22172_new_n4292_), .Y(core__abc_22172_new_n4293_));
INVX1 INVX1_877 ( .A(core__abc_22172_new_n4295_), .Y(core__abc_22172_new_n4296_));
INVX1 INVX1_878 ( .A(core__abc_22172_new_n4298_), .Y(core__abc_22172_new_n4299_));
INVX1 INVX1_879 ( .A(core__abc_22172_new_n4300_), .Y(core__abc_22172_new_n4301_));
INVX1 INVX1_88 ( .A(_abc_19873_new_n2380_), .Y(_abc_19873_new_n2381_));
INVX1 INVX1_880 ( .A(core__abc_22172_new_n4303_), .Y(core__abc_22172_new_n4304_));
INVX1 INVX1_881 ( .A(core__abc_22172_new_n4306_), .Y(core__abc_22172_new_n4307_));
INVX1 INVX1_882 ( .A(core__abc_22172_new_n4311_), .Y(core__abc_22172_new_n4313_));
INVX1 INVX1_883 ( .A(core__abc_22172_new_n4315_), .Y(core__abc_22172_new_n4316_));
INVX1 INVX1_884 ( .A(core_v3_reg_44_), .Y(core__abc_22172_new_n4318_));
INVX1 INVX1_885 ( .A(core__abc_22172_new_n4320_), .Y(core__abc_22172_new_n4321_));
INVX1 INVX1_886 ( .A(core__abc_22172_new_n4327_), .Y(core__abc_22172_new_n4328_));
INVX1 INVX1_887 ( .A(core__abc_22172_new_n4338_), .Y(core__abc_22172_new_n4339_));
INVX1 INVX1_888 ( .A(core__abc_22172_new_n4340_), .Y(core__abc_22172_new_n4341_));
INVX1 INVX1_889 ( .A(core__abc_22172_new_n4345_), .Y(core__abc_22172_new_n4346_));
INVX1 INVX1_89 ( .A(_abc_19873_new_n2385_), .Y(_abc_19873_new_n2386_));
INVX1 INVX1_890 ( .A(core__abc_22172_new_n4350_), .Y(core__abc_22172_new_n4351_));
INVX1 INVX1_891 ( .A(core__abc_22172_new_n4353_), .Y(core__abc_22172_new_n4355_));
INVX1 INVX1_892 ( .A(core__abc_22172_new_n4357_), .Y(core__abc_22172_new_n4358_));
INVX1 INVX1_893 ( .A(core__abc_22172_new_n4347_), .Y(core__abc_22172_new_n4360_));
INVX1 INVX1_894 ( .A(core__abc_22172_new_n4362_), .Y(core__abc_22172_new_n4363_));
INVX1 INVX1_895 ( .A(core__abc_22172_new_n4368_), .Y(core__abc_22172_new_n4369_));
INVX1 INVX1_896 ( .A(core__abc_22172_new_n4371_), .Y(core__abc_22172_new_n4372_));
INVX1 INVX1_897 ( .A(core_v3_reg_45_), .Y(core__abc_22172_new_n4374_));
INVX1 INVX1_898 ( .A(core__abc_22172_new_n4366_), .Y(core__abc_22172_new_n4378_));
INVX1 INVX1_899 ( .A(core__abc_22172_new_n4373_), .Y(core__abc_22172_new_n4379_));
INVX1 INVX1_9 ( .A(we), .Y(_abc_19873_new_n936_));
INVX1 INVX1_90 ( .A(_abc_19873_new_n2390_), .Y(_abc_19873_new_n2391_));
INVX1 INVX1_900 ( .A(core__abc_22172_new_n4375_), .Y(core__abc_22172_new_n4380_));
INVX1 INVX1_901 ( .A(core_key_82_), .Y(core__abc_22172_new_n4385_));
INVX1 INVX1_902 ( .A(core__abc_22172_new_n4387_), .Y(core__abc_22172_new_n4388_));
INVX1 INVX1_903 ( .A(core__abc_22172_new_n4400_), .Y(core__abc_22172_new_n4401_));
INVX1 INVX1_904 ( .A(core__abc_22172_new_n4405_), .Y(core__abc_22172_new_n4406_));
INVX1 INVX1_905 ( .A(core__abc_22172_new_n4408_), .Y(core__abc_22172_new_n4409_));
INVX1 INVX1_906 ( .A(core__abc_22172_new_n4413_), .Y(core__abc_22172_new_n4414_));
INVX1 INVX1_907 ( .A(core__abc_22172_new_n4417_), .Y(core__abc_22172_new_n4418_));
INVX1 INVX1_908 ( .A(core__abc_22172_new_n4420_), .Y(core__abc_22172_new_n4421_));
INVX1 INVX1_909 ( .A(core_v3_reg_46_), .Y(core__abc_22172_new_n4422_));
INVX1 INVX1_91 ( .A(_abc_19873_new_n2395_), .Y(_abc_19873_new_n2396_));
INVX1 INVX1_910 ( .A(core__abc_22172_new_n4426_), .Y(core__abc_22172_new_n4427_));
INVX1 INVX1_911 ( .A(core__abc_22172_new_n4428_), .Y(core__abc_22172_new_n4429_));
INVX1 INVX1_912 ( .A(core__abc_22172_new_n4432_), .Y(core__abc_22172_new_n4434_));
INVX1 INVX1_913 ( .A(core__abc_22172_new_n4439_), .Y(core__abc_22172_new_n4440_));
INVX1 INVX1_914 ( .A(core__abc_22172_new_n4458_), .Y(core__abc_22172_new_n4459_));
INVX1 INVX1_915 ( .A(core__abc_22172_new_n4462_), .Y(core__abc_22172_new_n4463_));
INVX1 INVX1_916 ( .A(core__abc_22172_new_n4464_), .Y(core__abc_22172_new_n4465_));
INVX1 INVX1_917 ( .A(core__abc_22172_new_n4468_), .Y(core__abc_22172_new_n4470_));
INVX1 INVX1_918 ( .A(core__abc_22172_new_n4472_), .Y(core__abc_22172_new_n4473_));
INVX1 INVX1_919 ( .A(core__abc_22172_new_n4475_), .Y(core__abc_22172_new_n4477_));
INVX1 INVX1_92 ( .A(_abc_19873_new_n2400_), .Y(_abc_19873_new_n2401_));
INVX1 INVX1_920 ( .A(core__abc_22172_new_n4479_), .Y(core__abc_22172_new_n4480_));
INVX1 INVX1_921 ( .A(core__abc_22172_new_n4483_), .Y(core__abc_22172_new_n4484_));
INVX1 INVX1_922 ( .A(core__abc_22172_new_n4487_), .Y(core__abc_22172_new_n4488_));
INVX1 INVX1_923 ( .A(core__abc_22172_new_n4489_), .Y(core__abc_22172_new_n4490_));
INVX1 INVX1_924 ( .A(core__abc_22172_new_n4492_), .Y(core__abc_22172_new_n4493_));
INVX1 INVX1_925 ( .A(core__abc_22172_new_n4496_), .Y(core__abc_22172_new_n4497_));
INVX1 INVX1_926 ( .A(core_v3_reg_47_), .Y(core__abc_22172_new_n4500_));
INVX1 INVX1_927 ( .A(core__abc_22172_new_n4498_), .Y(core__abc_22172_new_n4501_));
INVX1 INVX1_928 ( .A(core__abc_22172_new_n4503_), .Y(core__abc_22172_new_n4504_));
INVX1 INVX1_929 ( .A(core_key_84_), .Y(core__abc_22172_new_n4509_));
INVX1 INVX1_93 ( .A(_abc_19873_new_n2405_), .Y(_abc_19873_new_n2406_));
INVX1 INVX1_930 ( .A(core__abc_22172_new_n4511_), .Y(core__abc_22172_new_n4512_));
INVX1 INVX1_931 ( .A(core__abc_22172_new_n4522_), .Y(core__abc_22172_new_n4523_));
INVX1 INVX1_932 ( .A(core__abc_22172_new_n4526_), .Y(core__abc_22172_new_n4527_));
INVX1 INVX1_933 ( .A(core__abc_22172_new_n4530_), .Y(core__abc_22172_new_n4531_));
INVX1 INVX1_934 ( .A(core__abc_22172_new_n4532_), .Y(core__abc_22172_new_n4533_));
INVX1 INVX1_935 ( .A(core__abc_22172_new_n4536_), .Y(core__abc_22172_new_n4538_));
INVX1 INVX1_936 ( .A(core__abc_22172_new_n4540_), .Y(core__abc_22172_new_n4541_));
INVX1 INVX1_937 ( .A(core__abc_22172_new_n4485_), .Y(core__abc_22172_new_n4542_));
INVX1 INVX1_938 ( .A(core__abc_22172_new_n4545_), .Y(core__abc_22172_new_n4546_));
INVX1 INVX1_939 ( .A(core__abc_22172_new_n4547_), .Y(core__abc_22172_new_n4548_));
INVX1 INVX1_94 ( .A(_abc_19873_new_n2410_), .Y(_abc_19873_new_n2411_));
INVX1 INVX1_940 ( .A(core_key_85_), .Y(core__abc_22172_new_n4553_));
INVX1 INVX1_941 ( .A(core__abc_22172_new_n4555_), .Y(core__abc_22172_new_n4556_));
INVX1 INVX1_942 ( .A(core__abc_22172_new_n3247_), .Y(core__abc_22172_new_n4566_));
INVX1 INVX1_943 ( .A(core__abc_22172_new_n4539_), .Y(core__abc_22172_new_n4569_));
INVX1 INVX1_944 ( .A(core__abc_22172_new_n2175_), .Y(core__abc_22172_new_n4575_));
INVX1 INVX1_945 ( .A(core__abc_22172_new_n4577_), .Y(core__abc_22172_new_n4578_));
INVX1 INVX1_946 ( .A(core__abc_22172_new_n4579_), .Y(core__abc_22172_new_n4581_));
INVX1 INVX1_947 ( .A(core__abc_22172_new_n4585_), .Y(core__abc_22172_new_n4587_));
INVX1 INVX1_948 ( .A(core__abc_22172_new_n4589_), .Y(core__abc_22172_new_n4590_));
INVX1 INVX1_949 ( .A(core__abc_22172_new_n4593_), .Y(core__abc_22172_new_n4594_));
INVX1 INVX1_95 ( .A(_abc_19873_new_n2415_), .Y(_abc_19873_new_n2416_));
INVX1 INVX1_950 ( .A(core__abc_22172_new_n4595_), .Y(core__abc_22172_new_n4596_));
INVX1 INVX1_951 ( .A(core__abc_22172_new_n4599_), .Y(core__abc_22172_new_n4600_));
INVX1 INVX1_952 ( .A(core__abc_22172_new_n4602_), .Y(core__abc_22172_new_n4604_));
INVX1 INVX1_953 ( .A(core_key_86_), .Y(core__abc_22172_new_n4608_));
INVX1 INVX1_954 ( .A(core__abc_22172_new_n4610_), .Y(core__abc_22172_new_n4611_));
INVX1 INVX1_955 ( .A(core__abc_22172_new_n4624_), .Y(core__abc_22172_new_n4625_));
INVX1 INVX1_956 ( .A(core__abc_22172_new_n4627_), .Y(core__abc_22172_new_n4628_));
INVX1 INVX1_957 ( .A(core__abc_22172_new_n4631_), .Y(core__abc_22172_new_n4633_));
INVX1 INVX1_958 ( .A(core__abc_22172_new_n4623_), .Y(core__abc_22172_new_n4637_));
INVX1 INVX1_959 ( .A(core__abc_22172_new_n4635_), .Y(core__abc_22172_new_n4639_));
INVX1 INVX1_96 ( .A(_abc_19873_new_n2420_), .Y(_abc_19873_new_n2421_));
INVX1 INVX1_960 ( .A(core__abc_22172_new_n4641_), .Y(core__abc_22172_new_n4642_));
INVX1 INVX1_961 ( .A(core__abc_22172_new_n4643_), .Y(core__abc_22172_new_n4644_));
INVX1 INVX1_962 ( .A(core__abc_22172_new_n4646_), .Y(core__abc_22172_new_n4648_));
INVX1 INVX1_963 ( .A(core__abc_22172_new_n4653_), .Y(core__abc_22172_new_n4654_));
INVX1 INVX1_964 ( .A(core__abc_22172_new_n4640_), .Y(core__abc_22172_new_n4668_));
INVX1 INVX1_965 ( .A(core__abc_22172_new_n4597_), .Y(core__abc_22172_new_n4669_));
INVX1 INVX1_966 ( .A(core__abc_22172_new_n4679_), .Y(core__abc_22172_new_n4689_));
INVX1 INVX1_967 ( .A(core__abc_22172_new_n4686_), .Y(core__abc_22172_new_n4691_));
INVX1 INVX1_968 ( .A(core__abc_22172_new_n4696_), .Y(core__abc_22172_new_n4698_));
INVX1 INVX1_969 ( .A(core__abc_22172_new_n4700_), .Y(core__abc_22172_new_n4701_));
INVX1 INVX1_97 ( .A(_abc_19873_new_n2425_), .Y(_abc_19873_new_n2426_));
INVX1 INVX1_970 ( .A(core_v3_reg_8_), .Y(core__abc_22172_new_n4703_));
INVX1 INVX1_971 ( .A(core__abc_22172_new_n4705_), .Y(core__abc_22172_new_n4706_));
INVX1 INVX1_972 ( .A(core__abc_22172_new_n4694_), .Y(core__abc_22172_new_n4708_));
INVX1 INVX1_973 ( .A(core__abc_22172_new_n4710_), .Y(core__abc_22172_new_n4711_));
INVX1 INVX1_974 ( .A(core__abc_22172_new_n4676_), .Y(core__abc_22172_new_n4713_));
INVX1 INVX1_975 ( .A(core__abc_22172_new_n4715_), .Y(core__abc_22172_new_n4717_));
INVX1 INVX1_976 ( .A(core_key_88_), .Y(core__abc_22172_new_n4721_));
INVX1 INVX1_977 ( .A(core__abc_22172_new_n4723_), .Y(core__abc_22172_new_n4724_));
INVX1 INVX1_978 ( .A(core__abc_22172_new_n4734_), .Y(core__abc_22172_new_n4735_));
INVX1 INVX1_979 ( .A(core__abc_22172_new_n4739_), .Y(core__abc_22172_new_n4740_));
INVX1 INVX1_98 ( .A(_abc_19873_new_n2430_), .Y(_abc_19873_new_n2431_));
INVX1 INVX1_980 ( .A(core__abc_22172_new_n4744_), .Y(core__abc_22172_new_n4745_));
INVX1 INVX1_981 ( .A(core__abc_22172_new_n4738_), .Y(core__abc_22172_new_n4749_));
INVX1 INVX1_982 ( .A(core__abc_22172_new_n4747_), .Y(core__abc_22172_new_n4750_));
INVX1 INVX1_983 ( .A(core__abc_22172_new_n4709_), .Y(core__abc_22172_new_n4753_));
INVX1 INVX1_984 ( .A(core__abc_22172_new_n4712_), .Y(core__abc_22172_new_n4754_));
INVX1 INVX1_985 ( .A(core__abc_22172_new_n4757_), .Y(core__abc_22172_new_n4758_));
INVX1 INVX1_986 ( .A(core__abc_22172_new_n4759_), .Y(core__abc_22172_new_n4760_));
INVX1 INVX1_987 ( .A(core__abc_22172_new_n4766_), .Y(core__abc_22172_new_n4767_));
INVX1 INVX1_988 ( .A(core__abc_22172_new_n4752_), .Y(core__abc_22172_new_n4777_));
INVX1 INVX1_989 ( .A(core__abc_22172_new_n4748_), .Y(core__abc_22172_new_n4780_));
INVX1 INVX1_99 ( .A(_abc_19873_new_n2435_), .Y(_abc_19873_new_n2436_));
INVX1 INVX1_990 ( .A(core__abc_22172_new_n4788_), .Y(core__abc_22172_new_n4790_));
INVX1 INVX1_991 ( .A(core__abc_22172_new_n4792_), .Y(core__abc_22172_new_n4793_));
INVX1 INVX1_992 ( .A(core_v3_reg_10_), .Y(core__abc_22172_new_n4794_));
INVX1 INVX1_993 ( .A(core__abc_22172_new_n4796_), .Y(core__abc_22172_new_n4797_));
INVX1 INVX1_994 ( .A(core__abc_22172_new_n4800_), .Y(core__abc_22172_new_n4801_));
INVX1 INVX1_995 ( .A(core__abc_22172_new_n4804_), .Y(core__abc_22172_new_n4805_));
INVX1 INVX1_996 ( .A(core__abc_22172_new_n4808_), .Y(core__abc_22172_new_n4809_));
INVX1 INVX1_997 ( .A(core__abc_22172_new_n4810_), .Y(core__abc_22172_new_n4811_));
INVX1 INVX1_998 ( .A(core__abc_22172_new_n4813_), .Y(core__abc_22172_new_n4814_));
INVX1 INVX1_999 ( .A(core__abc_22172_new_n4820_), .Y(core__abc_22172_new_n4821_));
OR2X2 OR2X2_1 ( .A(_abc_19873_new_n882_), .B(_abc_19873_new_n889_), .Y(_abc_19873_new_n890_));
OR2X2 OR2X2_10 ( .A(_abc_19873_new_n927_), .B(_abc_19873_new_n932_), .Y(_abc_19873_new_n933_));
OR2X2 OR2X2_100 ( .A(_abc_19873_new_n1125_), .B(_abc_19873_new_n1116_), .Y(_abc_19873_new_n1126_));
OR2X2 OR2X2_1000 ( .A(core_v2_reg_52_), .B(core_v3_reg_52_), .Y(core__abc_22172_new_n2160_));
OR2X2 OR2X2_1001 ( .A(core__abc_22172_new_n2159_), .B(core__abc_22172_new_n2163_), .Y(core__abc_22172_new_n2164_));
OR2X2 OR2X2_1002 ( .A(core__abc_22172_new_n2165_), .B(core__abc_22172_new_n2166_), .Y(core__abc_22172_new_n2167_));
OR2X2 OR2X2_1003 ( .A(core__abc_22172_new_n2168_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n2169_));
OR2X2 OR2X2_1004 ( .A(core_siphash_word1_we), .B(core_siphash_word_116_), .Y(core__abc_22172_new_n2170_));
OR2X2 OR2X2_1005 ( .A(core_v1_reg_53_), .B(core_v0_reg_53_), .Y(core__abc_22172_new_n2175_));
OR2X2 OR2X2_1006 ( .A(core_v2_reg_53_), .B(core_v3_reg_53_), .Y(core__abc_22172_new_n2178_));
OR2X2 OR2X2_1007 ( .A(core__abc_22172_new_n2182_), .B(core__abc_22172_new_n2184_), .Y(core__abc_22172_new_n2185_));
OR2X2 OR2X2_1008 ( .A(core__abc_22172_new_n2185_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n2186_));
OR2X2 OR2X2_1009 ( .A(core_siphash_word1_we), .B(core_siphash_word_117_), .Y(core__abc_22172_new_n2187_));
OR2X2 OR2X2_101 ( .A(_abc_19873_new_n1128_), .B(_abc_19873_new_n1129_), .Y(_abc_19873_new_n1130_));
OR2X2 OR2X2_1010 ( .A(core_v1_reg_54_), .B(core_v0_reg_54_), .Y(core__abc_22172_new_n2190_));
OR2X2 OR2X2_1011 ( .A(core_v2_reg_54_), .B(core_v3_reg_54_), .Y(core__abc_22172_new_n2194_));
OR2X2 OR2X2_1012 ( .A(core__abc_22172_new_n2193_), .B(core__abc_22172_new_n2197_), .Y(core__abc_22172_new_n2198_));
OR2X2 OR2X2_1013 ( .A(core__abc_22172_new_n2199_), .B(core__abc_22172_new_n2200_), .Y(core__abc_22172_new_n2201_));
OR2X2 OR2X2_1014 ( .A(core__abc_22172_new_n2202_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n2203_));
OR2X2 OR2X2_1015 ( .A(core_siphash_word1_we), .B(core_siphash_word_118_), .Y(core__abc_22172_new_n2204_));
OR2X2 OR2X2_1016 ( .A(core_v1_reg_55_), .B(core_v0_reg_55_), .Y(core__abc_22172_new_n2207_));
OR2X2 OR2X2_1017 ( .A(core_v2_reg_55_), .B(core_v3_reg_55_), .Y(core__abc_22172_new_n2211_));
OR2X2 OR2X2_1018 ( .A(core__abc_22172_new_n2210_), .B(core__abc_22172_new_n2214_), .Y(core__abc_22172_new_n2215_));
OR2X2 OR2X2_1019 ( .A(core__abc_22172_new_n2216_), .B(core__abc_22172_new_n2217_), .Y(core__abc_22172_new_n2218_));
OR2X2 OR2X2_102 ( .A(_abc_19873_new_n1132_), .B(_abc_19873_new_n1133_), .Y(_abc_19873_new_n1134_));
OR2X2 OR2X2_1020 ( .A(core__abc_22172_new_n2219_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n2220_));
OR2X2 OR2X2_1021 ( .A(core_siphash_word1_we), .B(core_siphash_word_119_), .Y(core__abc_22172_new_n2221_));
OR2X2 OR2X2_1022 ( .A(core_v1_reg_56_), .B(core_v0_reg_56_), .Y(core__abc_22172_new_n2224_));
OR2X2 OR2X2_1023 ( .A(core_v2_reg_56_), .B(core_v3_reg_56_), .Y(core__abc_22172_new_n2228_));
OR2X2 OR2X2_1024 ( .A(core__abc_22172_new_n2227_), .B(core__abc_22172_new_n2231_), .Y(core__abc_22172_new_n2232_));
OR2X2 OR2X2_1025 ( .A(core__abc_22172_new_n2233_), .B(core__abc_22172_new_n2234_), .Y(core__abc_22172_new_n2235_));
OR2X2 OR2X2_1026 ( .A(core__abc_22172_new_n2236_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n2237_));
OR2X2 OR2X2_1027 ( .A(core_siphash_word1_we), .B(core_siphash_word_120_), .Y(core__abc_22172_new_n2238_));
OR2X2 OR2X2_1028 ( .A(core_v1_reg_57_), .B(core_v0_reg_57_), .Y(core__abc_22172_new_n2241_));
OR2X2 OR2X2_1029 ( .A(core_v2_reg_57_), .B(core_v3_reg_57_), .Y(core__abc_22172_new_n2245_));
OR2X2 OR2X2_103 ( .A(_abc_19873_new_n1134_), .B(_abc_19873_new_n1131_), .Y(_abc_19873_new_n1135_));
OR2X2 OR2X2_1030 ( .A(core__abc_22172_new_n2244_), .B(core__abc_22172_new_n2248_), .Y(core__abc_22172_new_n2249_));
OR2X2 OR2X2_1031 ( .A(core__abc_22172_new_n2250_), .B(core__abc_22172_new_n2251_), .Y(core__abc_22172_new_n2252_));
OR2X2 OR2X2_1032 ( .A(core__abc_22172_new_n2253_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n2254_));
OR2X2 OR2X2_1033 ( .A(core_siphash_word1_we), .B(core_siphash_word_121_), .Y(core__abc_22172_new_n2255_));
OR2X2 OR2X2_1034 ( .A(core_v1_reg_58_), .B(core_v0_reg_58_), .Y(core__abc_22172_new_n2258_));
OR2X2 OR2X2_1035 ( .A(core_v2_reg_58_), .B(core_v3_reg_58_), .Y(core__abc_22172_new_n2262_));
OR2X2 OR2X2_1036 ( .A(core__abc_22172_new_n2261_), .B(core__abc_22172_new_n2265_), .Y(core__abc_22172_new_n2266_));
OR2X2 OR2X2_1037 ( .A(core__abc_22172_new_n2267_), .B(core__abc_22172_new_n2268_), .Y(core__abc_22172_new_n2269_));
OR2X2 OR2X2_1038 ( .A(core__abc_22172_new_n2270_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n2271_));
OR2X2 OR2X2_1039 ( .A(core_siphash_word1_we), .B(core_siphash_word_122_), .Y(core__abc_22172_new_n2272_));
OR2X2 OR2X2_104 ( .A(_abc_19873_new_n1135_), .B(_abc_19873_new_n1130_), .Y(_abc_19873_new_n1136_));
OR2X2 OR2X2_1040 ( .A(core_v1_reg_59_), .B(core_v0_reg_59_), .Y(core__abc_22172_new_n2275_));
OR2X2 OR2X2_1041 ( .A(core_v2_reg_59_), .B(core_v3_reg_59_), .Y(core__abc_22172_new_n2279_));
OR2X2 OR2X2_1042 ( .A(core__abc_22172_new_n2278_), .B(core__abc_22172_new_n2282_), .Y(core__abc_22172_new_n2283_));
OR2X2 OR2X2_1043 ( .A(core__abc_22172_new_n2284_), .B(core__abc_22172_new_n2285_), .Y(core__abc_22172_new_n2286_));
OR2X2 OR2X2_1044 ( .A(core__abc_22172_new_n2287_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n2288_));
OR2X2 OR2X2_1045 ( .A(core_siphash_word1_we), .B(core_siphash_word_123_), .Y(core__abc_22172_new_n2289_));
OR2X2 OR2X2_1046 ( .A(core_v1_reg_60_), .B(core_v0_reg_60_), .Y(core__abc_22172_new_n2292_));
OR2X2 OR2X2_1047 ( .A(core_v2_reg_60_), .B(core_v3_reg_60_), .Y(core__abc_22172_new_n2296_));
OR2X2 OR2X2_1048 ( .A(core__abc_22172_new_n2295_), .B(core__abc_22172_new_n2299_), .Y(core__abc_22172_new_n2300_));
OR2X2 OR2X2_1049 ( .A(core__abc_22172_new_n2301_), .B(core__abc_22172_new_n2302_), .Y(core__abc_22172_new_n2303_));
OR2X2 OR2X2_105 ( .A(_abc_19873_new_n1138_), .B(_abc_19873_new_n1139_), .Y(_abc_19873_new_n1140_));
OR2X2 OR2X2_1050 ( .A(core__abc_22172_new_n2304_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n2305_));
OR2X2 OR2X2_1051 ( .A(core_siphash_word1_we), .B(core_siphash_word_124_), .Y(core__abc_22172_new_n2306_));
OR2X2 OR2X2_1052 ( .A(core_v1_reg_61_), .B(core_v0_reg_61_), .Y(core__abc_22172_new_n2309_));
OR2X2 OR2X2_1053 ( .A(core_v2_reg_61_), .B(core_v3_reg_61_), .Y(core__abc_22172_new_n2313_));
OR2X2 OR2X2_1054 ( .A(core__abc_22172_new_n2312_), .B(core__abc_22172_new_n2316_), .Y(core__abc_22172_new_n2317_));
OR2X2 OR2X2_1055 ( .A(core__abc_22172_new_n2318_), .B(core__abc_22172_new_n2319_), .Y(core__abc_22172_new_n2320_));
OR2X2 OR2X2_1056 ( .A(core__abc_22172_new_n2321_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n2322_));
OR2X2 OR2X2_1057 ( .A(core_siphash_word1_we), .B(core_siphash_word_125_), .Y(core__abc_22172_new_n2323_));
OR2X2 OR2X2_1058 ( .A(core_v1_reg_62_), .B(core_v0_reg_62_), .Y(core__abc_22172_new_n2326_));
OR2X2 OR2X2_1059 ( .A(core_v2_reg_62_), .B(core_v3_reg_62_), .Y(core__abc_22172_new_n2330_));
OR2X2 OR2X2_106 ( .A(_abc_19873_new_n1141_), .B(_abc_19873_new_n1142_), .Y(_abc_19873_new_n1143_));
OR2X2 OR2X2_1060 ( .A(core__abc_22172_new_n2329_), .B(core__abc_22172_new_n2333_), .Y(core__abc_22172_new_n2334_));
OR2X2 OR2X2_1061 ( .A(core__abc_22172_new_n2335_), .B(core__abc_22172_new_n2336_), .Y(core__abc_22172_new_n2337_));
OR2X2 OR2X2_1062 ( .A(core__abc_22172_new_n2338_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n2339_));
OR2X2 OR2X2_1063 ( .A(core_siphash_word1_we), .B(core_siphash_word_126_), .Y(core__abc_22172_new_n2340_));
OR2X2 OR2X2_1064 ( .A(core__abc_22172_new_n2343_), .B(core_v0_reg_63_), .Y(core__abc_22172_new_n2344_));
OR2X2 OR2X2_1065 ( .A(core__abc_22172_new_n2345_), .B(core_v1_reg_63_), .Y(core__abc_22172_new_n2346_));
OR2X2 OR2X2_1066 ( .A(core_v2_reg_63_), .B(core_v3_reg_63_), .Y(core__abc_22172_new_n2349_));
OR2X2 OR2X2_1067 ( .A(core__abc_22172_new_n2348_), .B(core__abc_22172_new_n2352_), .Y(core__abc_22172_new_n2353_));
OR2X2 OR2X2_1068 ( .A(core__abc_22172_new_n2354_), .B(core__abc_22172_new_n2347_), .Y(core__abc_22172_new_n2355_));
OR2X2 OR2X2_1069 ( .A(core__abc_22172_new_n2356_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n2357_));
OR2X2 OR2X2_107 ( .A(_abc_19873_new_n1140_), .B(_abc_19873_new_n1143_), .Y(_abc_19873_new_n1144_));
OR2X2 OR2X2_1070 ( .A(core_siphash_word1_we), .B(core_siphash_word_127_), .Y(core__abc_22172_new_n2358_));
OR2X2 OR2X2_1071 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_0_), .Y(core__abc_22172_new_n2365_));
OR2X2 OR2X2_1072 ( .A(core__abc_22172_new_n1270_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2367_));
OR2X2 OR2X2_1073 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_1_), .Y(core__abc_22172_new_n2370_));
OR2X2 OR2X2_1074 ( .A(core__abc_22172_new_n1291_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2371_));
OR2X2 OR2X2_1075 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_2_), .Y(core__abc_22172_new_n2374_));
OR2X2 OR2X2_1076 ( .A(core__abc_22172_new_n1309_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2375_));
OR2X2 OR2X2_1077 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_3_), .Y(core__abc_22172_new_n2378_));
OR2X2 OR2X2_1078 ( .A(core__abc_22172_new_n1327_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2379_));
OR2X2 OR2X2_1079 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_4_), .Y(core__abc_22172_new_n2382_));
OR2X2 OR2X2_108 ( .A(_abc_19873_new_n1144_), .B(_abc_19873_new_n1137_), .Y(_abc_19873_new_n1145_));
OR2X2 OR2X2_1080 ( .A(core__abc_22172_new_n1345_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2383_));
OR2X2 OR2X2_1081 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_5_), .Y(core__abc_22172_new_n2386_));
OR2X2 OR2X2_1082 ( .A(core__abc_22172_new_n1365_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2387_));
OR2X2 OR2X2_1083 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_6_), .Y(core__abc_22172_new_n2390_));
OR2X2 OR2X2_1084 ( .A(core__abc_22172_new_n1383_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2391_));
OR2X2 OR2X2_1085 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_7_), .Y(core__abc_22172_new_n2394_));
OR2X2 OR2X2_1086 ( .A(core__abc_22172_new_n1403_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2395_));
OR2X2 OR2X2_1087 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_8_), .Y(core__abc_22172_new_n2398_));
OR2X2 OR2X2_1088 ( .A(core__abc_22172_new_n1420_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2399_));
OR2X2 OR2X2_1089 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_9_), .Y(core__abc_22172_new_n2402_));
OR2X2 OR2X2_109 ( .A(_abc_19873_new_n1145_), .B(_abc_19873_new_n1136_), .Y(_abc_19873_new_n1146_));
OR2X2 OR2X2_1090 ( .A(core__abc_22172_new_n1437_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2403_));
OR2X2 OR2X2_1091 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_10_), .Y(core__abc_22172_new_n2406_));
OR2X2 OR2X2_1092 ( .A(core__abc_22172_new_n1454_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2407_));
OR2X2 OR2X2_1093 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_11_), .Y(core__abc_22172_new_n2410_));
OR2X2 OR2X2_1094 ( .A(core__abc_22172_new_n1471_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2411_));
OR2X2 OR2X2_1095 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_12_), .Y(core__abc_22172_new_n2414_));
OR2X2 OR2X2_1096 ( .A(core__abc_22172_new_n1488_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2415_));
OR2X2 OR2X2_1097 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_13_), .Y(core__abc_22172_new_n2418_));
OR2X2 OR2X2_1098 ( .A(core__abc_22172_new_n1505_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2419_));
OR2X2 OR2X2_1099 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_14_), .Y(core__abc_22172_new_n2422_));
OR2X2 OR2X2_11 ( .A(_abc_19873_new_n933_), .B(_abc_19873_new_n922_), .Y(_abc_19873_new_n934_));
OR2X2 OR2X2_110 ( .A(_abc_19873_new_n1148_), .B(_abc_19873_new_n1149_), .Y(_abc_19873_new_n1150_));
OR2X2 OR2X2_1100 ( .A(core__abc_22172_new_n1522_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2423_));
OR2X2 OR2X2_1101 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_15_), .Y(core__abc_22172_new_n2426_));
OR2X2 OR2X2_1102 ( .A(core__abc_22172_new_n1539_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2427_));
OR2X2 OR2X2_1103 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_16_), .Y(core__abc_22172_new_n2430_));
OR2X2 OR2X2_1104 ( .A(core__abc_22172_new_n1556_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2431_));
OR2X2 OR2X2_1105 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_17_), .Y(core__abc_22172_new_n2434_));
OR2X2 OR2X2_1106 ( .A(core__abc_22172_new_n1573_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2435_));
OR2X2 OR2X2_1107 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_18_), .Y(core__abc_22172_new_n2438_));
OR2X2 OR2X2_1108 ( .A(core__abc_22172_new_n1590_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2439_));
OR2X2 OR2X2_1109 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_19_), .Y(core__abc_22172_new_n2442_));
OR2X2 OR2X2_111 ( .A(_abc_19873_new_n1152_), .B(_abc_19873_new_n1153_), .Y(_abc_19873_new_n1154_));
OR2X2 OR2X2_1110 ( .A(core__abc_22172_new_n1607_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2443_));
OR2X2 OR2X2_1111 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_20_), .Y(core__abc_22172_new_n2446_));
OR2X2 OR2X2_1112 ( .A(core__abc_22172_new_n1624_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2447_));
OR2X2 OR2X2_1113 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_21_), .Y(core__abc_22172_new_n2450_));
OR2X2 OR2X2_1114 ( .A(core__abc_22172_new_n1641_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2451_));
OR2X2 OR2X2_1115 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_22_), .Y(core__abc_22172_new_n2454_));
OR2X2 OR2X2_1116 ( .A(core__abc_22172_new_n1658_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2455_));
OR2X2 OR2X2_1117 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_23_), .Y(core__abc_22172_new_n2458_));
OR2X2 OR2X2_1118 ( .A(core__abc_22172_new_n1675_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2459_));
OR2X2 OR2X2_1119 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_24_), .Y(core__abc_22172_new_n2462_));
OR2X2 OR2X2_112 ( .A(_abc_19873_new_n1154_), .B(_abc_19873_new_n1151_), .Y(_abc_19873_new_n1155_));
OR2X2 OR2X2_1120 ( .A(core__abc_22172_new_n1692_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2463_));
OR2X2 OR2X2_1121 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_25_), .Y(core__abc_22172_new_n2466_));
OR2X2 OR2X2_1122 ( .A(core__abc_22172_new_n1709_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2467_));
OR2X2 OR2X2_1123 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_26_), .Y(core__abc_22172_new_n2470_));
OR2X2 OR2X2_1124 ( .A(core__abc_22172_new_n1726_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2471_));
OR2X2 OR2X2_1125 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_27_), .Y(core__abc_22172_new_n2474_));
OR2X2 OR2X2_1126 ( .A(core__abc_22172_new_n1743_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2475_));
OR2X2 OR2X2_1127 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_28_), .Y(core__abc_22172_new_n2478_));
OR2X2 OR2X2_1128 ( .A(core__abc_22172_new_n1760_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2479_));
OR2X2 OR2X2_1129 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_29_), .Y(core__abc_22172_new_n2482_));
OR2X2 OR2X2_113 ( .A(_abc_19873_new_n1155_), .B(_abc_19873_new_n1150_), .Y(_abc_19873_new_n1156_));
OR2X2 OR2X2_1130 ( .A(core__abc_22172_new_n1777_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2483_));
OR2X2 OR2X2_1131 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_30_), .Y(core__abc_22172_new_n2486_));
OR2X2 OR2X2_1132 ( .A(core__abc_22172_new_n1794_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2487_));
OR2X2 OR2X2_1133 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_31_), .Y(core__abc_22172_new_n2490_));
OR2X2 OR2X2_1134 ( .A(core__abc_22172_new_n1811_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2491_));
OR2X2 OR2X2_1135 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_32_), .Y(core__abc_22172_new_n2494_));
OR2X2 OR2X2_1136 ( .A(core__abc_22172_new_n1828_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2495_));
OR2X2 OR2X2_1137 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_33_), .Y(core__abc_22172_new_n2498_));
OR2X2 OR2X2_1138 ( .A(core__abc_22172_new_n1845_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2499_));
OR2X2 OR2X2_1139 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_34_), .Y(core__abc_22172_new_n2502_));
OR2X2 OR2X2_114 ( .A(_abc_19873_new_n1158_), .B(_abc_19873_new_n1159_), .Y(_abc_19873_new_n1160_));
OR2X2 OR2X2_1140 ( .A(core__abc_22172_new_n1862_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2503_));
OR2X2 OR2X2_1141 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_35_), .Y(core__abc_22172_new_n2506_));
OR2X2 OR2X2_1142 ( .A(core__abc_22172_new_n1879_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2507_));
OR2X2 OR2X2_1143 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_36_), .Y(core__abc_22172_new_n2510_));
OR2X2 OR2X2_1144 ( .A(core__abc_22172_new_n1896_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2511_));
OR2X2 OR2X2_1145 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_37_), .Y(core__abc_22172_new_n2514_));
OR2X2 OR2X2_1146 ( .A(core__abc_22172_new_n1913_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2515_));
OR2X2 OR2X2_1147 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_38_), .Y(core__abc_22172_new_n2518_));
OR2X2 OR2X2_1148 ( .A(core__abc_22172_new_n1930_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2519_));
OR2X2 OR2X2_1149 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_39_), .Y(core__abc_22172_new_n2522_));
OR2X2 OR2X2_115 ( .A(_abc_19873_new_n1161_), .B(_abc_19873_new_n1162_), .Y(_abc_19873_new_n1163_));
OR2X2 OR2X2_1150 ( .A(core__abc_22172_new_n1947_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2523_));
OR2X2 OR2X2_1151 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_40_), .Y(core__abc_22172_new_n2526_));
OR2X2 OR2X2_1152 ( .A(core__abc_22172_new_n1964_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2527_));
OR2X2 OR2X2_1153 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_41_), .Y(core__abc_22172_new_n2530_));
OR2X2 OR2X2_1154 ( .A(core__abc_22172_new_n1981_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2531_));
OR2X2 OR2X2_1155 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_42_), .Y(core__abc_22172_new_n2534_));
OR2X2 OR2X2_1156 ( .A(core__abc_22172_new_n1998_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2535_));
OR2X2 OR2X2_1157 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_43_), .Y(core__abc_22172_new_n2538_));
OR2X2 OR2X2_1158 ( .A(core__abc_22172_new_n2015_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2539_));
OR2X2 OR2X2_1159 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_44_), .Y(core__abc_22172_new_n2542_));
OR2X2 OR2X2_116 ( .A(_abc_19873_new_n1160_), .B(_abc_19873_new_n1163_), .Y(_abc_19873_new_n1164_));
OR2X2 OR2X2_1160 ( .A(core__abc_22172_new_n2032_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2543_));
OR2X2 OR2X2_1161 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_45_), .Y(core__abc_22172_new_n2546_));
OR2X2 OR2X2_1162 ( .A(core__abc_22172_new_n2049_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2547_));
OR2X2 OR2X2_1163 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_46_), .Y(core__abc_22172_new_n2550_));
OR2X2 OR2X2_1164 ( .A(core__abc_22172_new_n2066_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2551_));
OR2X2 OR2X2_1165 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_47_), .Y(core__abc_22172_new_n2554_));
OR2X2 OR2X2_1166 ( .A(core__abc_22172_new_n2083_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2555_));
OR2X2 OR2X2_1167 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_48_), .Y(core__abc_22172_new_n2558_));
OR2X2 OR2X2_1168 ( .A(core__abc_22172_new_n2100_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2559_));
OR2X2 OR2X2_1169 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_49_), .Y(core__abc_22172_new_n2562_));
OR2X2 OR2X2_117 ( .A(_abc_19873_new_n1164_), .B(_abc_19873_new_n1157_), .Y(_abc_19873_new_n1165_));
OR2X2 OR2X2_1170 ( .A(core__abc_22172_new_n2117_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2563_));
OR2X2 OR2X2_1171 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_50_), .Y(core__abc_22172_new_n2566_));
OR2X2 OR2X2_1172 ( .A(core__abc_22172_new_n2134_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2567_));
OR2X2 OR2X2_1173 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_51_), .Y(core__abc_22172_new_n2570_));
OR2X2 OR2X2_1174 ( .A(core__abc_22172_new_n2151_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2571_));
OR2X2 OR2X2_1175 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_52_), .Y(core__abc_22172_new_n2574_));
OR2X2 OR2X2_1176 ( .A(core__abc_22172_new_n2168_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2575_));
OR2X2 OR2X2_1177 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_53_), .Y(core__abc_22172_new_n2578_));
OR2X2 OR2X2_1178 ( .A(core__abc_22172_new_n2185_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2579_));
OR2X2 OR2X2_1179 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_54_), .Y(core__abc_22172_new_n2582_));
OR2X2 OR2X2_118 ( .A(_abc_19873_new_n1165_), .B(_abc_19873_new_n1156_), .Y(_abc_19873_new_n1166_));
OR2X2 OR2X2_1180 ( .A(core__abc_22172_new_n2202_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2583_));
OR2X2 OR2X2_1181 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_55_), .Y(core__abc_22172_new_n2586_));
OR2X2 OR2X2_1182 ( .A(core__abc_22172_new_n2219_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2587_));
OR2X2 OR2X2_1183 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_56_), .Y(core__abc_22172_new_n2590_));
OR2X2 OR2X2_1184 ( .A(core__abc_22172_new_n2236_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2591_));
OR2X2 OR2X2_1185 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_57_), .Y(core__abc_22172_new_n2594_));
OR2X2 OR2X2_1186 ( .A(core__abc_22172_new_n2253_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2595_));
OR2X2 OR2X2_1187 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_58_), .Y(core__abc_22172_new_n2598_));
OR2X2 OR2X2_1188 ( .A(core__abc_22172_new_n2270_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2599_));
OR2X2 OR2X2_1189 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_59_), .Y(core__abc_22172_new_n2602_));
OR2X2 OR2X2_119 ( .A(_abc_19873_new_n1169_), .B(_abc_19873_new_n1170_), .Y(_abc_19873_new_n1171_));
OR2X2 OR2X2_1190 ( .A(core__abc_22172_new_n2287_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2603_));
OR2X2 OR2X2_1191 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_60_), .Y(core__abc_22172_new_n2606_));
OR2X2 OR2X2_1192 ( .A(core__abc_22172_new_n2304_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2607_));
OR2X2 OR2X2_1193 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_61_), .Y(core__abc_22172_new_n2610_));
OR2X2 OR2X2_1194 ( .A(core__abc_22172_new_n2321_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2611_));
OR2X2 OR2X2_1195 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_62_), .Y(core__abc_22172_new_n2614_));
OR2X2 OR2X2_1196 ( .A(core__abc_22172_new_n2338_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2615_));
OR2X2 OR2X2_1197 ( .A(core__abc_22172_new_n2364_), .B(core_siphash_word_63_), .Y(core__abc_22172_new_n2618_));
OR2X2 OR2X2_1198 ( .A(core__abc_22172_new_n2356_), .B(core__abc_22172_new_n2366_), .Y(core__abc_22172_new_n2619_));
OR2X2 OR2X2_1199 ( .A(core__abc_22172_new_n2624_), .B(core__abc_22172_new_n2622_), .Y(core__abc_22172_new_n2625_));
OR2X2 OR2X2_12 ( .A(_abc_19873_new_n911_), .B(_abc_19873_new_n934_), .Y(_abc_19873_new_n935_));
OR2X2 OR2X2_120 ( .A(_abc_19873_new_n1171_), .B(_abc_19873_new_n1168_), .Y(_abc_19873_new_n1172_));
OR2X2 OR2X2_1200 ( .A(core__abc_22172_new_n2626_), .B(core__abc_22172_new_n1240_), .Y(core__0ready_reg_0_0_));
OR2X2 OR2X2_1201 ( .A(core__abc_22172_new_n2628_), .B(core_loop_ctr_reg_0_), .Y(core__abc_22172_new_n2636_));
OR2X2 OR2X2_1202 ( .A(core__abc_22172_new_n2634_), .B(core_loop_ctr_reg_1_), .Y(core__abc_22172_new_n2639_));
OR2X2 OR2X2_1203 ( .A(core__abc_22172_new_n2632_), .B(core__abc_22172_new_n2642_), .Y(core__abc_22172_new_n2643_));
OR2X2 OR2X2_1204 ( .A(core__abc_22172_new_n2646_), .B(core_loop_ctr_reg_2_), .Y(core__abc_22172_new_n2647_));
OR2X2 OR2X2_1205 ( .A(core__abc_22172_new_n2632_), .B(core__abc_22172_new_n2650_), .Y(core__abc_22172_new_n2651_));
OR2X2 OR2X2_1206 ( .A(core__abc_22172_new_n2651_), .B(core__abc_22172_new_n1142_), .Y(core__abc_22172_new_n2654_));
OR2X2 OR2X2_1207 ( .A(core__abc_22172_new_n2655_), .B(core_loop_ctr_reg_3_), .Y(core__abc_22172_new_n2656_));
OR2X2 OR2X2_1208 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_0_), .Y(core__abc_22172_new_n2661_));
OR2X2 OR2X2_1209 ( .A(core__abc_22172_new_n2662_), .B(core_mi_0_), .Y(core__abc_22172_new_n2663_));
OR2X2 OR2X2_121 ( .A(_abc_19873_new_n1173_), .B(_abc_19873_new_n1174_), .Y(_abc_19873_new_n1175_));
OR2X2 OR2X2_1210 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_1_), .Y(core__abc_22172_new_n2666_));
OR2X2 OR2X2_1211 ( .A(core__abc_22172_new_n2662_), .B(core_mi_1_), .Y(core__abc_22172_new_n2667_));
OR2X2 OR2X2_1212 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_2_), .Y(core__abc_22172_new_n2670_));
OR2X2 OR2X2_1213 ( .A(core__abc_22172_new_n2662_), .B(core_mi_2_), .Y(core__abc_22172_new_n2671_));
OR2X2 OR2X2_1214 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_3_), .Y(core__abc_22172_new_n2674_));
OR2X2 OR2X2_1215 ( .A(core__abc_22172_new_n2662_), .B(core_mi_3_), .Y(core__abc_22172_new_n2675_));
OR2X2 OR2X2_1216 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_4_), .Y(core__abc_22172_new_n2678_));
OR2X2 OR2X2_1217 ( .A(core__abc_22172_new_n2662_), .B(core_mi_4_), .Y(core__abc_22172_new_n2679_));
OR2X2 OR2X2_1218 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_5_), .Y(core__abc_22172_new_n2682_));
OR2X2 OR2X2_1219 ( .A(core__abc_22172_new_n2662_), .B(core_mi_5_), .Y(core__abc_22172_new_n2683_));
OR2X2 OR2X2_122 ( .A(_abc_19873_new_n1176_), .B(_abc_19873_new_n1177_), .Y(_abc_19873_new_n1178_));
OR2X2 OR2X2_1220 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_6_), .Y(core__abc_22172_new_n2686_));
OR2X2 OR2X2_1221 ( .A(core__abc_22172_new_n2662_), .B(core_mi_6_), .Y(core__abc_22172_new_n2687_));
OR2X2 OR2X2_1222 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_7_), .Y(core__abc_22172_new_n2690_));
OR2X2 OR2X2_1223 ( .A(core__abc_22172_new_n2662_), .B(core_mi_7_), .Y(core__abc_22172_new_n2691_));
OR2X2 OR2X2_1224 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_8_), .Y(core__abc_22172_new_n2694_));
OR2X2 OR2X2_1225 ( .A(core__abc_22172_new_n2662_), .B(core_mi_8_), .Y(core__abc_22172_new_n2695_));
OR2X2 OR2X2_1226 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_9_), .Y(core__abc_22172_new_n2698_));
OR2X2 OR2X2_1227 ( .A(core__abc_22172_new_n2662_), .B(core_mi_9_), .Y(core__abc_22172_new_n2699_));
OR2X2 OR2X2_1228 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_10_), .Y(core__abc_22172_new_n2702_));
OR2X2 OR2X2_1229 ( .A(core__abc_22172_new_n2662_), .B(core_mi_10_), .Y(core__abc_22172_new_n2703_));
OR2X2 OR2X2_123 ( .A(_abc_19873_new_n1175_), .B(_abc_19873_new_n1178_), .Y(_abc_19873_new_n1179_));
OR2X2 OR2X2_1230 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_11_), .Y(core__abc_22172_new_n2706_));
OR2X2 OR2X2_1231 ( .A(core__abc_22172_new_n2662_), .B(core_mi_11_), .Y(core__abc_22172_new_n2707_));
OR2X2 OR2X2_1232 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_12_), .Y(core__abc_22172_new_n2710_));
OR2X2 OR2X2_1233 ( .A(core__abc_22172_new_n2662_), .B(core_mi_12_), .Y(core__abc_22172_new_n2711_));
OR2X2 OR2X2_1234 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_13_), .Y(core__abc_22172_new_n2714_));
OR2X2 OR2X2_1235 ( .A(core__abc_22172_new_n2662_), .B(core_mi_13_), .Y(core__abc_22172_new_n2715_));
OR2X2 OR2X2_1236 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_14_), .Y(core__abc_22172_new_n2718_));
OR2X2 OR2X2_1237 ( .A(core__abc_22172_new_n2662_), .B(core_mi_14_), .Y(core__abc_22172_new_n2719_));
OR2X2 OR2X2_1238 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_15_), .Y(core__abc_22172_new_n2722_));
OR2X2 OR2X2_1239 ( .A(core__abc_22172_new_n2662_), .B(core_mi_15_), .Y(core__abc_22172_new_n2723_));
OR2X2 OR2X2_124 ( .A(_abc_19873_new_n1180_), .B(_abc_19873_new_n1181_), .Y(_abc_19873_new_n1182_));
OR2X2 OR2X2_1240 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_16_), .Y(core__abc_22172_new_n2726_));
OR2X2 OR2X2_1241 ( .A(core__abc_22172_new_n2662_), .B(core_mi_16_), .Y(core__abc_22172_new_n2727_));
OR2X2 OR2X2_1242 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_17_), .Y(core__abc_22172_new_n2730_));
OR2X2 OR2X2_1243 ( .A(core__abc_22172_new_n2662_), .B(core_mi_17_), .Y(core__abc_22172_new_n2731_));
OR2X2 OR2X2_1244 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_18_), .Y(core__abc_22172_new_n2734_));
OR2X2 OR2X2_1245 ( .A(core__abc_22172_new_n2662_), .B(core_mi_18_), .Y(core__abc_22172_new_n2735_));
OR2X2 OR2X2_1246 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_19_), .Y(core__abc_22172_new_n2738_));
OR2X2 OR2X2_1247 ( .A(core__abc_22172_new_n2662_), .B(core_mi_19_), .Y(core__abc_22172_new_n2739_));
OR2X2 OR2X2_1248 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_20_), .Y(core__abc_22172_new_n2742_));
OR2X2 OR2X2_1249 ( .A(core__abc_22172_new_n2662_), .B(core_mi_20_), .Y(core__abc_22172_new_n2743_));
OR2X2 OR2X2_125 ( .A(_abc_19873_new_n1183_), .B(_abc_19873_new_n1037_), .Y(_abc_19873_new_n1184_));
OR2X2 OR2X2_1250 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_21_), .Y(core__abc_22172_new_n2746_));
OR2X2 OR2X2_1251 ( .A(core__abc_22172_new_n2662_), .B(core_mi_21_), .Y(core__abc_22172_new_n2747_));
OR2X2 OR2X2_1252 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_22_), .Y(core__abc_22172_new_n2750_));
OR2X2 OR2X2_1253 ( .A(core__abc_22172_new_n2662_), .B(core_mi_22_), .Y(core__abc_22172_new_n2751_));
OR2X2 OR2X2_1254 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_23_), .Y(core__abc_22172_new_n2754_));
OR2X2 OR2X2_1255 ( .A(core__abc_22172_new_n2662_), .B(core_mi_23_), .Y(core__abc_22172_new_n2755_));
OR2X2 OR2X2_1256 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_24_), .Y(core__abc_22172_new_n2758_));
OR2X2 OR2X2_1257 ( .A(core__abc_22172_new_n2662_), .B(core_mi_24_), .Y(core__abc_22172_new_n2759_));
OR2X2 OR2X2_1258 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_25_), .Y(core__abc_22172_new_n2762_));
OR2X2 OR2X2_1259 ( .A(core__abc_22172_new_n2662_), .B(core_mi_25_), .Y(core__abc_22172_new_n2763_));
OR2X2 OR2X2_126 ( .A(_abc_19873_new_n1182_), .B(_abc_19873_new_n1184_), .Y(_abc_19873_new_n1185_));
OR2X2 OR2X2_1260 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_26_), .Y(core__abc_22172_new_n2766_));
OR2X2 OR2X2_1261 ( .A(core__abc_22172_new_n2662_), .B(core_mi_26_), .Y(core__abc_22172_new_n2767_));
OR2X2 OR2X2_1262 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_27_), .Y(core__abc_22172_new_n2770_));
OR2X2 OR2X2_1263 ( .A(core__abc_22172_new_n2662_), .B(core_mi_27_), .Y(core__abc_22172_new_n2771_));
OR2X2 OR2X2_1264 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_28_), .Y(core__abc_22172_new_n2774_));
OR2X2 OR2X2_1265 ( .A(core__abc_22172_new_n2662_), .B(core_mi_28_), .Y(core__abc_22172_new_n2775_));
OR2X2 OR2X2_1266 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_29_), .Y(core__abc_22172_new_n2778_));
OR2X2 OR2X2_1267 ( .A(core__abc_22172_new_n2662_), .B(core_mi_29_), .Y(core__abc_22172_new_n2779_));
OR2X2 OR2X2_1268 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_30_), .Y(core__abc_22172_new_n2782_));
OR2X2 OR2X2_1269 ( .A(core__abc_22172_new_n2662_), .B(core_mi_30_), .Y(core__abc_22172_new_n2783_));
OR2X2 OR2X2_127 ( .A(_abc_19873_new_n1179_), .B(_abc_19873_new_n1185_), .Y(_abc_19873_new_n1186_));
OR2X2 OR2X2_1270 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_31_), .Y(core__abc_22172_new_n2786_));
OR2X2 OR2X2_1271 ( .A(core__abc_22172_new_n2662_), .B(core_mi_31_), .Y(core__abc_22172_new_n2787_));
OR2X2 OR2X2_1272 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_32_), .Y(core__abc_22172_new_n2790_));
OR2X2 OR2X2_1273 ( .A(core__abc_22172_new_n2662_), .B(core_mi_32_), .Y(core__abc_22172_new_n2791_));
OR2X2 OR2X2_1274 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_33_), .Y(core__abc_22172_new_n2794_));
OR2X2 OR2X2_1275 ( .A(core__abc_22172_new_n2662_), .B(core_mi_33_), .Y(core__abc_22172_new_n2795_));
OR2X2 OR2X2_1276 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_34_), .Y(core__abc_22172_new_n2798_));
OR2X2 OR2X2_1277 ( .A(core__abc_22172_new_n2662_), .B(core_mi_34_), .Y(core__abc_22172_new_n2799_));
OR2X2 OR2X2_1278 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_35_), .Y(core__abc_22172_new_n2802_));
OR2X2 OR2X2_1279 ( .A(core__abc_22172_new_n2662_), .B(core_mi_35_), .Y(core__abc_22172_new_n2803_));
OR2X2 OR2X2_128 ( .A(_abc_19873_new_n1186_), .B(_abc_19873_new_n1172_), .Y(_abc_19873_new_n1187_));
OR2X2 OR2X2_1280 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_36_), .Y(core__abc_22172_new_n2806_));
OR2X2 OR2X2_1281 ( .A(core__abc_22172_new_n2662_), .B(core_mi_36_), .Y(core__abc_22172_new_n2807_));
OR2X2 OR2X2_1282 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_37_), .Y(core__abc_22172_new_n2810_));
OR2X2 OR2X2_1283 ( .A(core__abc_22172_new_n2662_), .B(core_mi_37_), .Y(core__abc_22172_new_n2811_));
OR2X2 OR2X2_1284 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_38_), .Y(core__abc_22172_new_n2814_));
OR2X2 OR2X2_1285 ( .A(core__abc_22172_new_n2662_), .B(core_mi_38_), .Y(core__abc_22172_new_n2815_));
OR2X2 OR2X2_1286 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_39_), .Y(core__abc_22172_new_n2818_));
OR2X2 OR2X2_1287 ( .A(core__abc_22172_new_n2662_), .B(core_mi_39_), .Y(core__abc_22172_new_n2819_));
OR2X2 OR2X2_1288 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_40_), .Y(core__abc_22172_new_n2822_));
OR2X2 OR2X2_1289 ( .A(core__abc_22172_new_n2662_), .B(core_mi_40_), .Y(core__abc_22172_new_n2823_));
OR2X2 OR2X2_129 ( .A(_abc_19873_new_n1189_), .B(_abc_19873_new_n1190_), .Y(_abc_19873_new_n1191_));
OR2X2 OR2X2_1290 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_41_), .Y(core__abc_22172_new_n2826_));
OR2X2 OR2X2_1291 ( .A(core__abc_22172_new_n2662_), .B(core_mi_41_), .Y(core__abc_22172_new_n2827_));
OR2X2 OR2X2_1292 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_42_), .Y(core__abc_22172_new_n2830_));
OR2X2 OR2X2_1293 ( .A(core__abc_22172_new_n2662_), .B(core_mi_42_), .Y(core__abc_22172_new_n2831_));
OR2X2 OR2X2_1294 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_43_), .Y(core__abc_22172_new_n2834_));
OR2X2 OR2X2_1295 ( .A(core__abc_22172_new_n2662_), .B(core_mi_43_), .Y(core__abc_22172_new_n2835_));
OR2X2 OR2X2_1296 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_44_), .Y(core__abc_22172_new_n2838_));
OR2X2 OR2X2_1297 ( .A(core__abc_22172_new_n2662_), .B(core_mi_44_), .Y(core__abc_22172_new_n2839_));
OR2X2 OR2X2_1298 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_45_), .Y(core__abc_22172_new_n2842_));
OR2X2 OR2X2_1299 ( .A(core__abc_22172_new_n2662_), .B(core_mi_45_), .Y(core__abc_22172_new_n2843_));
OR2X2 OR2X2_13 ( .A(_abc_19873_new_n939_), .B(_abc_19873_new_n940_), .Y(_abc_19873_new_n941_));
OR2X2 OR2X2_130 ( .A(_abc_19873_new_n994_), .B(_abc_19873_new_n1018_), .Y(_abc_19873_new_n1192_));
OR2X2 OR2X2_1300 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_46_), .Y(core__abc_22172_new_n2846_));
OR2X2 OR2X2_1301 ( .A(core__abc_22172_new_n2662_), .B(core_mi_46_), .Y(core__abc_22172_new_n2847_));
OR2X2 OR2X2_1302 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_47_), .Y(core__abc_22172_new_n2850_));
OR2X2 OR2X2_1303 ( .A(core__abc_22172_new_n2662_), .B(core_mi_47_), .Y(core__abc_22172_new_n2851_));
OR2X2 OR2X2_1304 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_48_), .Y(core__abc_22172_new_n2854_));
OR2X2 OR2X2_1305 ( .A(core__abc_22172_new_n2662_), .B(core_mi_48_), .Y(core__abc_22172_new_n2855_));
OR2X2 OR2X2_1306 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_49_), .Y(core__abc_22172_new_n2858_));
OR2X2 OR2X2_1307 ( .A(core__abc_22172_new_n2662_), .B(core_mi_49_), .Y(core__abc_22172_new_n2859_));
OR2X2 OR2X2_1308 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_50_), .Y(core__abc_22172_new_n2862_));
OR2X2 OR2X2_1309 ( .A(core__abc_22172_new_n2662_), .B(core_mi_50_), .Y(core__abc_22172_new_n2863_));
OR2X2 OR2X2_131 ( .A(_abc_19873_new_n1192_), .B(_abc_19873_new_n1193_), .Y(_abc_19873_new_n1194_));
OR2X2 OR2X2_1310 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_51_), .Y(core__abc_22172_new_n2866_));
OR2X2 OR2X2_1311 ( .A(core__abc_22172_new_n2662_), .B(core_mi_51_), .Y(core__abc_22172_new_n2867_));
OR2X2 OR2X2_1312 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_52_), .Y(core__abc_22172_new_n2870_));
OR2X2 OR2X2_1313 ( .A(core__abc_22172_new_n2662_), .B(core_mi_52_), .Y(core__abc_22172_new_n2871_));
OR2X2 OR2X2_1314 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_53_), .Y(core__abc_22172_new_n2874_));
OR2X2 OR2X2_1315 ( .A(core__abc_22172_new_n2662_), .B(core_mi_53_), .Y(core__abc_22172_new_n2875_));
OR2X2 OR2X2_1316 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_54_), .Y(core__abc_22172_new_n2878_));
OR2X2 OR2X2_1317 ( .A(core__abc_22172_new_n2662_), .B(core_mi_54_), .Y(core__abc_22172_new_n2879_));
OR2X2 OR2X2_1318 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_55_), .Y(core__abc_22172_new_n2882_));
OR2X2 OR2X2_1319 ( .A(core__abc_22172_new_n2662_), .B(core_mi_55_), .Y(core__abc_22172_new_n2883_));
OR2X2 OR2X2_132 ( .A(_abc_19873_new_n1194_), .B(_abc_19873_new_n1191_), .Y(_abc_19873_new_n1195_));
OR2X2 OR2X2_1320 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_56_), .Y(core__abc_22172_new_n2886_));
OR2X2 OR2X2_1321 ( .A(core__abc_22172_new_n2662_), .B(core_mi_56_), .Y(core__abc_22172_new_n2887_));
OR2X2 OR2X2_1322 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_57_), .Y(core__abc_22172_new_n2890_));
OR2X2 OR2X2_1323 ( .A(core__abc_22172_new_n2662_), .B(core_mi_57_), .Y(core__abc_22172_new_n2891_));
OR2X2 OR2X2_1324 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_58_), .Y(core__abc_22172_new_n2894_));
OR2X2 OR2X2_1325 ( .A(core__abc_22172_new_n2662_), .B(core_mi_58_), .Y(core__abc_22172_new_n2895_));
OR2X2 OR2X2_1326 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_59_), .Y(core__abc_22172_new_n2898_));
OR2X2 OR2X2_1327 ( .A(core__abc_22172_new_n2662_), .B(core_mi_59_), .Y(core__abc_22172_new_n2899_));
OR2X2 OR2X2_1328 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_60_), .Y(core__abc_22172_new_n2902_));
OR2X2 OR2X2_1329 ( .A(core__abc_22172_new_n2662_), .B(core_mi_60_), .Y(core__abc_22172_new_n2903_));
OR2X2 OR2X2_133 ( .A(_abc_19873_new_n1197_), .B(_abc_19873_new_n1198_), .Y(_abc_19873_new_n1199_));
OR2X2 OR2X2_1330 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_61_), .Y(core__abc_22172_new_n2906_));
OR2X2 OR2X2_1331 ( .A(core__abc_22172_new_n2662_), .B(core_mi_61_), .Y(core__abc_22172_new_n2907_));
OR2X2 OR2X2_1332 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_62_), .Y(core__abc_22172_new_n2910_));
OR2X2 OR2X2_1333 ( .A(core__abc_22172_new_n2662_), .B(core_mi_62_), .Y(core__abc_22172_new_n2911_));
OR2X2 OR2X2_1334 ( .A(core__abc_22172_new_n2660_), .B(core_mi_reg_63_), .Y(core__abc_22172_new_n2914_));
OR2X2 OR2X2_1335 ( .A(core__abc_22172_new_n2662_), .B(core_mi_63_), .Y(core__abc_22172_new_n2915_));
OR2X2 OR2X2_1336 ( .A(core__abc_22172_new_n2918_), .B(core__abc_22172_new_n1276_), .Y(core__abc_22172_new_n2919_));
OR2X2 OR2X2_1337 ( .A(core__abc_22172_new_n2922_), .B(core__abc_22172_new_n1315_), .Y(core__abc_22172_new_n2923_));
OR2X2 OR2X2_1338 ( .A(core__abc_22172_new_n2921_), .B(core__abc_22172_new_n2923_), .Y(core__abc_22172_new_n2924_));
OR2X2 OR2X2_1339 ( .A(core__abc_22172_new_n1333_), .B(core__abc_22172_new_n1351_), .Y(core__abc_22172_new_n2929_));
OR2X2 OR2X2_134 ( .A(_abc_19873_new_n1199_), .B(_abc_19873_new_n1196_), .Y(_abc_19873_new_n1200_));
OR2X2 OR2X2_1340 ( .A(core__abc_22172_new_n2932_), .B(core__abc_22172_new_n1389_), .Y(core__abc_22172_new_n2933_));
OR2X2 OR2X2_1341 ( .A(core__abc_22172_new_n2931_), .B(core__abc_22172_new_n2933_), .Y(core__abc_22172_new_n2934_));
OR2X2 OR2X2_1342 ( .A(core__abc_22172_new_n2928_), .B(core__abc_22172_new_n2934_), .Y(core__abc_22172_new_n2935_));
OR2X2 OR2X2_1343 ( .A(core__abc_22172_new_n1409_), .B(core__abc_22172_new_n1426_), .Y(core__abc_22172_new_n2944_));
OR2X2 OR2X2_1344 ( .A(core__abc_22172_new_n1468_), .B(core__abc_22172_new_n1444_), .Y(core__abc_22172_new_n2947_));
OR2X2 OR2X2_1345 ( .A(core__abc_22172_new_n2949_), .B(core__abc_22172_new_n2946_), .Y(core__abc_22172_new_n2950_));
OR2X2 OR2X2_1346 ( .A(core__abc_22172_new_n1502_), .B(core__abc_22172_new_n1478_), .Y(core__abc_22172_new_n2952_));
OR2X2 OR2X2_1347 ( .A(core__abc_22172_new_n2956_), .B(core__abc_22172_new_n1528_), .Y(core__abc_22172_new_n2957_));
OR2X2 OR2X2_1348 ( .A(core__abc_22172_new_n2955_), .B(core__abc_22172_new_n2957_), .Y(core__abc_22172_new_n2958_));
OR2X2 OR2X2_1349 ( .A(core__abc_22172_new_n2951_), .B(core__abc_22172_new_n2958_), .Y(core__abc_22172_new_n2959_));
OR2X2 OR2X2_135 ( .A(_abc_19873_new_n1201_), .B(_abc_19873_new_n1202_), .Y(_abc_19873_new_n1203_));
OR2X2 OR2X2_1350 ( .A(core__abc_22172_new_n2943_), .B(core__abc_22172_new_n2959_), .Y(core__abc_22172_new_n2960_));
OR2X2 OR2X2_1351 ( .A(core__abc_22172_new_n1545_), .B(core__abc_22172_new_n1562_), .Y(core__abc_22172_new_n2977_));
OR2X2 OR2X2_1352 ( .A(core__abc_22172_new_n2980_), .B(core__abc_22172_new_n1596_), .Y(core__abc_22172_new_n2981_));
OR2X2 OR2X2_1353 ( .A(core__abc_22172_new_n2979_), .B(core__abc_22172_new_n2981_), .Y(core__abc_22172_new_n2982_));
OR2X2 OR2X2_1354 ( .A(core__abc_22172_new_n2985_), .B(core__abc_22172_new_n2984_), .Y(core__abc_22172_new_n2986_));
OR2X2 OR2X2_1355 ( .A(core__abc_22172_new_n2989_), .B(core__abc_22172_new_n1664_), .Y(core__abc_22172_new_n2990_));
OR2X2 OR2X2_1356 ( .A(core__abc_22172_new_n2988_), .B(core__abc_22172_new_n2990_), .Y(core__abc_22172_new_n2991_));
OR2X2 OR2X2_1357 ( .A(core__abc_22172_new_n2983_), .B(core__abc_22172_new_n2991_), .Y(core__abc_22172_new_n2992_));
OR2X2 OR2X2_1358 ( .A(core__abc_22172_new_n2995_), .B(core__abc_22172_new_n2994_), .Y(core__abc_22172_new_n2996_));
OR2X2 OR2X2_1359 ( .A(core__abc_22172_new_n2999_), .B(core__abc_22172_new_n1732_), .Y(core__abc_22172_new_n3000_));
OR2X2 OR2X2_136 ( .A(_abc_19873_new_n1204_), .B(_abc_19873_new_n1205_), .Y(_abc_19873_new_n1206_));
OR2X2 OR2X2_1360 ( .A(core__abc_22172_new_n2998_), .B(core__abc_22172_new_n3000_), .Y(core__abc_22172_new_n3001_));
OR2X2 OR2X2_1361 ( .A(core__abc_22172_new_n3003_), .B(core__abc_22172_new_n1800_), .Y(core__abc_22172_new_n3004_));
OR2X2 OR2X2_1362 ( .A(core__abc_22172_new_n3006_), .B(core__abc_22172_new_n3005_), .Y(core__abc_22172_new_n3007_));
OR2X2 OR2X2_1363 ( .A(core__abc_22172_new_n3009_), .B(core__abc_22172_new_n3004_), .Y(core__abc_22172_new_n3010_));
OR2X2 OR2X2_1364 ( .A(core__abc_22172_new_n3002_), .B(core__abc_22172_new_n3010_), .Y(core__abc_22172_new_n3011_));
OR2X2 OR2X2_1365 ( .A(core__abc_22172_new_n2993_), .B(core__abc_22172_new_n3011_), .Y(core__abc_22172_new_n3012_));
OR2X2 OR2X2_1366 ( .A(core__abc_22172_new_n2976_), .B(core__abc_22172_new_n3012_), .Y(core__abc_22172_new_n3013_));
OR2X2 OR2X2_1367 ( .A(core__abc_22172_new_n1289_), .B(core__abc_22172_new_n1259_), .Y(core__abc_22172_new_n3015_));
OR2X2 OR2X2_1368 ( .A(core__abc_22172_new_n3016_), .B(core__abc_22172_new_n3017_), .Y(core__abc_22172_new_n3018_));
OR2X2 OR2X2_1369 ( .A(core__abc_22172_new_n3020_), .B(core__abc_22172_new_n3021_), .Y(core__abc_22172_new_n3022_));
OR2X2 OR2X2_137 ( .A(_abc_19873_new_n1203_), .B(_abc_19873_new_n1206_), .Y(_abc_19873_new_n1207_));
OR2X2 OR2X2_1370 ( .A(core__abc_22172_new_n3024_), .B(core__abc_22172_new_n3025_), .Y(core__abc_22172_new_n3026_));
OR2X2 OR2X2_1371 ( .A(core__abc_22172_new_n3028_), .B(core__abc_22172_new_n3029_), .Y(core__abc_22172_new_n3030_));
OR2X2 OR2X2_1372 ( .A(core__abc_22172_new_n3033_), .B(core__abc_22172_new_n3014_), .Y(core__abc_22172_new_n3034_));
OR2X2 OR2X2_1373 ( .A(core__abc_22172_new_n1265_), .B(core_v3_reg_48_), .Y(core__abc_22172_new_n3037_));
OR2X2 OR2X2_1374 ( .A(core__abc_22172_new_n3042_), .B(core__abc_22172_new_n3039_), .Y(core__abc_22172_new_n3043_));
OR2X2 OR2X2_1375 ( .A(core__abc_22172_new_n3046_), .B(core__abc_22172_new_n3045_), .Y(core__abc_22172_new_n3047_));
OR2X2 OR2X2_1376 ( .A(core__abc_22172_new_n3049_), .B(core__abc_22172_new_n1318_), .Y(core__abc_22172_new_n3050_));
OR2X2 OR2X2_1377 ( .A(core__abc_22172_new_n1283_), .B(core__abc_22172_new_n3053_), .Y(core__abc_22172_new_n3054_));
OR2X2 OR2X2_1378 ( .A(core__abc_22172_new_n3057_), .B(core__abc_22172_new_n3055_), .Y(core__abc_22172_new_n3058_));
OR2X2 OR2X2_1379 ( .A(core__abc_22172_new_n3066_), .B(core__abc_22172_new_n1358_), .Y(core__abc_22172_new_n3067_));
OR2X2 OR2X2_138 ( .A(_abc_19873_new_n1207_), .B(_abc_19873_new_n1200_), .Y(_abc_19873_new_n1208_));
OR2X2 OR2X2_1380 ( .A(core__abc_22172_new_n3070_), .B(core__abc_22172_new_n1392_), .Y(core__abc_22172_new_n3071_));
OR2X2 OR2X2_1381 ( .A(core__abc_22172_new_n3069_), .B(core__abc_22172_new_n3071_), .Y(core__abc_22172_new_n3072_));
OR2X2 OR2X2_1382 ( .A(core__abc_22172_new_n3064_), .B(core__abc_22172_new_n3072_), .Y(core__abc_22172_new_n3073_));
OR2X2 OR2X2_1383 ( .A(core__abc_22172_new_n3083_), .B(core__abc_22172_new_n3082_), .Y(core__abc_22172_new_n3084_));
OR2X2 OR2X2_1384 ( .A(core__abc_22172_new_n3087_), .B(core__abc_22172_new_n1463_), .Y(core__abc_22172_new_n3088_));
OR2X2 OR2X2_1385 ( .A(core__abc_22172_new_n3086_), .B(core__abc_22172_new_n3088_), .Y(core__abc_22172_new_n3089_));
OR2X2 OR2X2_1386 ( .A(core__abc_22172_new_n1503_), .B(core__abc_22172_new_n1481_), .Y(core__abc_22172_new_n3091_));
OR2X2 OR2X2_1387 ( .A(core__abc_22172_new_n3095_), .B(core__abc_22172_new_n1531_), .Y(core__abc_22172_new_n3096_));
OR2X2 OR2X2_1388 ( .A(core__abc_22172_new_n3094_), .B(core__abc_22172_new_n3096_), .Y(core__abc_22172_new_n3097_));
OR2X2 OR2X2_1389 ( .A(core__abc_22172_new_n3097_), .B(core__abc_22172_new_n3090_), .Y(core__abc_22172_new_n3098_));
OR2X2 OR2X2_139 ( .A(_abc_19873_new_n1208_), .B(_abc_19873_new_n1195_), .Y(_abc_19873_new_n1209_));
OR2X2 OR2X2_1390 ( .A(core__abc_22172_new_n3081_), .B(core__abc_22172_new_n3098_), .Y(core__abc_22172_new_n3099_));
OR2X2 OR2X2_1391 ( .A(core__abc_22172_new_n1571_), .B(core__abc_22172_new_n1549_), .Y(core__abc_22172_new_n3116_));
OR2X2 OR2X2_1392 ( .A(core__abc_22172_new_n3120_), .B(core__abc_22172_new_n1599_), .Y(core__abc_22172_new_n3121_));
OR2X2 OR2X2_1393 ( .A(core__abc_22172_new_n3119_), .B(core__abc_22172_new_n3121_), .Y(core__abc_22172_new_n3122_));
OR2X2 OR2X2_1394 ( .A(core__abc_22172_new_n3125_), .B(core__abc_22172_new_n3124_), .Y(core__abc_22172_new_n3126_));
OR2X2 OR2X2_1395 ( .A(core__abc_22172_new_n3129_), .B(core__abc_22172_new_n1667_), .Y(core__abc_22172_new_n3130_));
OR2X2 OR2X2_1396 ( .A(core__abc_22172_new_n3128_), .B(core__abc_22172_new_n3130_), .Y(core__abc_22172_new_n3131_));
OR2X2 OR2X2_1397 ( .A(core__abc_22172_new_n3123_), .B(core__abc_22172_new_n3131_), .Y(core__abc_22172_new_n3132_));
OR2X2 OR2X2_1398 ( .A(core__abc_22172_new_n3135_), .B(core__abc_22172_new_n3134_), .Y(core__abc_22172_new_n3136_));
OR2X2 OR2X2_1399 ( .A(core__abc_22172_new_n3139_), .B(core__abc_22172_new_n1735_), .Y(core__abc_22172_new_n3140_));
OR2X2 OR2X2_14 ( .A(_abc_19873_new_n942_), .B(_abc_19873_new_n943_), .Y(_abc_19873_new_n944_));
OR2X2 OR2X2_140 ( .A(_abc_19873_new_n1212_), .B(_abc_19873_new_n1213_), .Y(_abc_19873_new_n1214_));
OR2X2 OR2X2_1400 ( .A(core__abc_22172_new_n3138_), .B(core__abc_22172_new_n3140_), .Y(core__abc_22172_new_n3141_));
OR2X2 OR2X2_1401 ( .A(core__abc_22172_new_n3143_), .B(core__abc_22172_new_n1803_), .Y(core__abc_22172_new_n3144_));
OR2X2 OR2X2_1402 ( .A(core__abc_22172_new_n3146_), .B(core__abc_22172_new_n3145_), .Y(core__abc_22172_new_n3147_));
OR2X2 OR2X2_1403 ( .A(core__abc_22172_new_n3149_), .B(core__abc_22172_new_n3144_), .Y(core__abc_22172_new_n3150_));
OR2X2 OR2X2_1404 ( .A(core__abc_22172_new_n3142_), .B(core__abc_22172_new_n3150_), .Y(core__abc_22172_new_n3151_));
OR2X2 OR2X2_1405 ( .A(core__abc_22172_new_n3133_), .B(core__abc_22172_new_n3151_), .Y(core__abc_22172_new_n3152_));
OR2X2 OR2X2_1406 ( .A(core__abc_22172_new_n3115_), .B(core__abc_22172_new_n3152_), .Y(core__abc_22172_new_n3153_));
OR2X2 OR2X2_1407 ( .A(core__abc_22172_new_n3163_), .B(core__abc_22172_new_n3162_), .Y(core__abc_22172_new_n3164_));
OR2X2 OR2X2_1408 ( .A(core__abc_22172_new_n3167_), .B(core__abc_22172_new_n1871_), .Y(core__abc_22172_new_n3168_));
OR2X2 OR2X2_1409 ( .A(core__abc_22172_new_n3166_), .B(core__abc_22172_new_n3168_), .Y(core__abc_22172_new_n3169_));
OR2X2 OR2X2_141 ( .A(_abc_19873_new_n1215_), .B(_abc_19873_new_n1216_), .Y(_abc_19873_new_n1217_));
OR2X2 OR2X2_1410 ( .A(core__abc_22172_new_n3171_), .B(core__abc_22172_new_n1939_), .Y(core__abc_22172_new_n3172_));
OR2X2 OR2X2_1411 ( .A(core__abc_22172_new_n3174_), .B(core__abc_22172_new_n3173_), .Y(core__abc_22172_new_n3175_));
OR2X2 OR2X2_1412 ( .A(core__abc_22172_new_n3177_), .B(core__abc_22172_new_n3172_), .Y(core__abc_22172_new_n3178_));
OR2X2 OR2X2_1413 ( .A(core__abc_22172_new_n3170_), .B(core__abc_22172_new_n3178_), .Y(core__abc_22172_new_n3179_));
OR2X2 OR2X2_1414 ( .A(core__abc_22172_new_n3161_), .B(core__abc_22172_new_n3179_), .Y(core__abc_22172_new_n3180_));
OR2X2 OR2X2_1415 ( .A(core__abc_22172_new_n3182_), .B(core__abc_22172_new_n3048_), .Y(core__abc_22172_new_n3183_));
OR2X2 OR2X2_1416 ( .A(core__abc_22172_new_n3184_), .B(core__abc_22172_new_n1990_), .Y(core__abc_22172_new_n3185_));
OR2X2 OR2X2_1417 ( .A(core__abc_22172_new_n3187_), .B(core__abc_22172_new_n3188_), .Y(core__abc_22172_new_n3189_));
OR2X2 OR2X2_1418 ( .A(core__abc_22172_new_n3189_), .B(core_v3_reg_27_), .Y(core__abc_22172_new_n3192_));
OR2X2 OR2X2_1419 ( .A(core__abc_22172_new_n3194_), .B(core__abc_22172_new_n3044_), .Y(core__abc_22172_new_n3195_));
OR2X2 OR2X2_142 ( .A(_abc_19873_new_n1214_), .B(_abc_19873_new_n1217_), .Y(_abc_19873_new_n1218_));
OR2X2 OR2X2_1420 ( .A(core__abc_22172_new_n3199_), .B(core__abc_22172_new_n3202_), .Y(core__abc_22172_new_n3203_));
OR2X2 OR2X2_1421 ( .A(core__abc_22172_new_n3193_), .B(core__abc_22172_new_n3043_), .Y(core__abc_22172_new_n3206_));
OR2X2 OR2X2_1422 ( .A(core__abc_22172_new_n3209_), .B(core__abc_22172_new_n3211_), .Y(core__abc_22172_new_n3212_));
OR2X2 OR2X2_1423 ( .A(core__abc_22172_new_n3216_), .B(core__abc_22172_new_n3212_), .Y(core__abc_22172_new_n3217_));
OR2X2 OR2X2_1424 ( .A(core_v3_reg_0_), .B(core_mi_0_), .Y(core__abc_22172_new_n3222_));
OR2X2 OR2X2_1425 ( .A(core__abc_22172_new_n3219_), .B(core__abc_22172_new_n3224_), .Y(core__abc_22172_new_n3225_));
OR2X2 OR2X2_1426 ( .A(core__abc_22172_new_n3217_), .B(core__abc_22172_new_n3225_), .Y(core__abc_22172_new_n3226_));
OR2X2 OR2X2_1427 ( .A(core__abc_22172_new_n3208_), .B(core__abc_22172_new_n3226_), .Y(core__abc_22172_new_n3227_));
OR2X2 OR2X2_1428 ( .A(core__abc_22172_new_n3228_), .B(core_v3_reg_0_), .Y(core__abc_22172_new_n3229_));
OR2X2 OR2X2_1429 ( .A(core__abc_22172_new_n3237_), .B(core__abc_22172_new_n3235_), .Y(core__abc_22172_new_n3238_));
OR2X2 OR2X2_143 ( .A(_abc_19873_new_n1218_), .B(_abc_19873_new_n1211_), .Y(_abc_19873_new_n1219_));
OR2X2 OR2X2_1430 ( .A(core__abc_22172_new_n3234_), .B(core__abc_22172_new_n3238_), .Y(core__abc_22172_new_n3239_));
OR2X2 OR2X2_1431 ( .A(core__abc_22172_new_n3241_), .B(core__abc_22172_new_n3242_), .Y(core__abc_22172_new_n3243_));
OR2X2 OR2X2_1432 ( .A(core__abc_22172_new_n3244_), .B(core__abc_22172_new_n3240_), .Y(core__abc_22172_new_n3245_));
OR2X2 OR2X2_1433 ( .A(core__abc_22172_new_n3243_), .B(core_v3_reg_49_), .Y(core__abc_22172_new_n3246_));
OR2X2 OR2X2_1434 ( .A(core__abc_22172_new_n3239_), .B(core__abc_22172_new_n3247_), .Y(core__abc_22172_new_n3250_));
OR2X2 OR2X2_1435 ( .A(core__abc_22172_new_n3251_), .B(core__abc_22172_new_n3042_), .Y(core__abc_22172_new_n3254_));
OR2X2 OR2X2_1436 ( .A(core__abc_22172_new_n3259_), .B(core__abc_22172_new_n2008_), .Y(core__abc_22172_new_n3260_));
OR2X2 OR2X2_1437 ( .A(core__abc_22172_new_n3258_), .B(core__abc_22172_new_n3260_), .Y(core__abc_22172_new_n3261_));
OR2X2 OR2X2_1438 ( .A(core__abc_22172_new_n3263_), .B(core__abc_22172_new_n3261_), .Y(core__abc_22172_new_n3264_));
OR2X2 OR2X2_1439 ( .A(core__abc_22172_new_n3266_), .B(core__abc_22172_new_n3267_), .Y(core__abc_22172_new_n3268_));
OR2X2 OR2X2_144 ( .A(_abc_19873_new_n1220_), .B(_abc_19873_new_n1221_), .Y(_abc_19873_new_n1222_));
OR2X2 OR2X2_1440 ( .A(core__abc_22172_new_n3269_), .B(core__abc_22172_new_n3256_), .Y(core__abc_22172_new_n3270_));
OR2X2 OR2X2_1441 ( .A(core__abc_22172_new_n3268_), .B(core_v3_reg_28_), .Y(core__abc_22172_new_n3271_));
OR2X2 OR2X2_1442 ( .A(core__abc_22172_new_n3273_), .B(core__abc_22172_new_n3255_), .Y(core__abc_22172_new_n3274_));
OR2X2 OR2X2_1443 ( .A(core__abc_22172_new_n3272_), .B(core__abc_22172_new_n3275_), .Y(core__abc_22172_new_n3276_));
OR2X2 OR2X2_1444 ( .A(core_v3_reg_1_), .B(core_mi_1_), .Y(core__abc_22172_new_n3283_));
OR2X2 OR2X2_1445 ( .A(core__abc_22172_new_n3280_), .B(core__abc_22172_new_n3285_), .Y(core__abc_22172_new_n3286_));
OR2X2 OR2X2_1446 ( .A(core__abc_22172_new_n3217_), .B(core__abc_22172_new_n3286_), .Y(core__abc_22172_new_n3287_));
OR2X2 OR2X2_1447 ( .A(core__abc_22172_new_n3278_), .B(core__abc_22172_new_n3287_), .Y(core__abc_22172_new_n3288_));
OR2X2 OR2X2_1448 ( .A(core__abc_22172_new_n3228_), .B(core_v3_reg_1_), .Y(core__abc_22172_new_n3289_));
OR2X2 OR2X2_1449 ( .A(core__abc_22172_new_n3252_), .B(core__abc_22172_new_n3292_), .Y(core__abc_22172_new_n3293_));
OR2X2 OR2X2_145 ( .A(_abc_19873_new_n1222_), .B(_abc_19873_new_n1223_), .Y(_abc_19873_new_n1224_));
OR2X2 OR2X2_1450 ( .A(core__abc_22172_new_n3237_), .B(core__abc_22172_new_n3296_), .Y(core__abc_22172_new_n3297_));
OR2X2 OR2X2_1451 ( .A(core__abc_22172_new_n3297_), .B(core__abc_22172_new_n1853_), .Y(core__abc_22172_new_n3300_));
OR2X2 OR2X2_1452 ( .A(core__abc_22172_new_n3305_), .B(core__abc_22172_new_n3306_), .Y(core__abc_22172_new_n3307_));
OR2X2 OR2X2_1453 ( .A(core__abc_22172_new_n3308_), .B(core__abc_22172_new_n3303_), .Y(core__abc_22172_new_n3309_));
OR2X2 OR2X2_1454 ( .A(core__abc_22172_new_n3307_), .B(core_v3_reg_50_), .Y(core__abc_22172_new_n3310_));
OR2X2 OR2X2_1455 ( .A(core__abc_22172_new_n3312_), .B(core__abc_22172_new_n3314_), .Y(core__abc_22172_new_n3315_));
OR2X2 OR2X2_1456 ( .A(core__abc_22172_new_n3293_), .B(core__abc_22172_new_n3316_), .Y(core__abc_22172_new_n3319_));
OR2X2 OR2X2_1457 ( .A(core__abc_22172_new_n3267_), .B(core__abc_22172_new_n2025_), .Y(core__abc_22172_new_n3321_));
OR2X2 OR2X2_1458 ( .A(core__abc_22172_new_n3323_), .B(core__abc_22172_new_n3324_), .Y(core__abc_22172_new_n3325_));
OR2X2 OR2X2_1459 ( .A(core__abc_22172_new_n3325_), .B(core_v3_reg_29_), .Y(core__abc_22172_new_n3328_));
OR2X2 OR2X2_146 ( .A(_abc_19873_new_n1225_), .B(_abc_19873_new_n1226_), .Y(_abc_19873_new_n1227_));
OR2X2 OR2X2_1460 ( .A(core__abc_22172_new_n3330_), .B(core__abc_22172_new_n3320_), .Y(core__abc_22172_new_n3331_));
OR2X2 OR2X2_1461 ( .A(core__abc_22172_new_n3329_), .B(core__abc_22172_new_n3332_), .Y(core__abc_22172_new_n3333_));
OR2X2 OR2X2_1462 ( .A(core_v3_reg_2_), .B(core_mi_2_), .Y(core__abc_22172_new_n3339_));
OR2X2 OR2X2_1463 ( .A(core__abc_22172_new_n3336_), .B(core__abc_22172_new_n3341_), .Y(core__abc_22172_new_n3342_));
OR2X2 OR2X2_1464 ( .A(core__abc_22172_new_n3217_), .B(core__abc_22172_new_n3342_), .Y(core__abc_22172_new_n3343_));
OR2X2 OR2X2_1465 ( .A(core__abc_22172_new_n3335_), .B(core__abc_22172_new_n3343_), .Y(core__abc_22172_new_n3344_));
OR2X2 OR2X2_1466 ( .A(core__abc_22172_new_n3228_), .B(core_v3_reg_2_), .Y(core__abc_22172_new_n3345_));
OR2X2 OR2X2_1467 ( .A(core__abc_22172_new_n3351_), .B(core__abc_22172_new_n3350_), .Y(core__abc_22172_new_n3352_));
OR2X2 OR2X2_1468 ( .A(core__abc_22172_new_n3349_), .B(core__abc_22172_new_n3353_), .Y(core__abc_22172_new_n3354_));
OR2X2 OR2X2_1469 ( .A(core__abc_22172_new_n3357_), .B(core__abc_22172_new_n3355_), .Y(core__abc_22172_new_n3358_));
OR2X2 OR2X2_147 ( .A(_abc_19873_new_n1039_), .B(_abc_19873_new_n1227_), .Y(_abc_19873_new_n1228_));
OR2X2 OR2X2_1470 ( .A(core__abc_22172_new_n3359_), .B(core_v3_reg_30_), .Y(core__abc_22172_new_n3360_));
OR2X2 OR2X2_1471 ( .A(core__abc_22172_new_n3358_), .B(core__abc_22172_new_n3361_), .Y(core__abc_22172_new_n3362_));
OR2X2 OR2X2_1472 ( .A(core__abc_22172_new_n3317_), .B(core__abc_22172_new_n3314_), .Y(core__abc_22172_new_n3364_));
OR2X2 OR2X2_1473 ( .A(core__abc_22172_new_n3365_), .B(core__abc_22172_new_n1876_), .Y(core__abc_22172_new_n3368_));
OR2X2 OR2X2_1474 ( .A(core__abc_22172_new_n3374_), .B(core__abc_22172_new_n3375_), .Y(core__abc_22172_new_n3376_));
OR2X2 OR2X2_1475 ( .A(core__abc_22172_new_n3376_), .B(core_v3_reg_51_), .Y(core__abc_22172_new_n3379_));
OR2X2 OR2X2_1476 ( .A(core__abc_22172_new_n3388_), .B(core__abc_22172_new_n3364_), .Y(core__abc_22172_new_n3389_));
OR2X2 OR2X2_1477 ( .A(core__abc_22172_new_n3390_), .B(core__abc_22172_new_n3387_), .Y(core__abc_22172_new_n3391_));
OR2X2 OR2X2_1478 ( .A(core__abc_22172_new_n3393_), .B(core__abc_22172_new_n3363_), .Y(core__abc_22172_new_n3394_));
OR2X2 OR2X2_1479 ( .A(core__abc_22172_new_n3392_), .B(core__abc_22172_new_n3395_), .Y(core__abc_22172_new_n3396_));
OR2X2 OR2X2_148 ( .A(_abc_19873_new_n1228_), .B(_abc_19873_new_n1224_), .Y(_abc_19873_new_n1229_));
OR2X2 OR2X2_1480 ( .A(core_v3_reg_3_), .B(core_mi_3_), .Y(core__abc_22172_new_n3402_));
OR2X2 OR2X2_1481 ( .A(core__abc_22172_new_n3399_), .B(core__abc_22172_new_n3404_), .Y(core__abc_22172_new_n3405_));
OR2X2 OR2X2_1482 ( .A(core__abc_22172_new_n3217_), .B(core__abc_22172_new_n3405_), .Y(core__abc_22172_new_n3406_));
OR2X2 OR2X2_1483 ( .A(core__abc_22172_new_n3398_), .B(core__abc_22172_new_n3406_), .Y(core__abc_22172_new_n3407_));
OR2X2 OR2X2_1484 ( .A(core__abc_22172_new_n3228_), .B(core_v3_reg_3_), .Y(core__abc_22172_new_n3408_));
OR2X2 OR2X2_1485 ( .A(core__abc_22172_new_n3413_), .B(core__abc_22172_new_n1868_), .Y(core__abc_22172_new_n3414_));
OR2X2 OR2X2_1486 ( .A(core__abc_22172_new_n3412_), .B(core__abc_22172_new_n3414_), .Y(core__abc_22172_new_n3415_));
OR2X2 OR2X2_1487 ( .A(core__abc_22172_new_n3417_), .B(core__abc_22172_new_n3415_), .Y(core__abc_22172_new_n3418_));
OR2X2 OR2X2_1488 ( .A(core__abc_22172_new_n3421_), .B(core__abc_22172_new_n3419_), .Y(core__abc_22172_new_n3422_));
OR2X2 OR2X2_1489 ( .A(core__abc_22172_new_n3425_), .B(core__abc_22172_new_n3424_), .Y(core__abc_22172_new_n3426_));
OR2X2 OR2X2_149 ( .A(_abc_19873_new_n1229_), .B(_abc_19873_new_n1219_), .Y(_abc_19873_new_n1230_));
OR2X2 OR2X2_1490 ( .A(core__abc_22172_new_n3429_), .B(core__abc_22172_new_n3427_), .Y(core__abc_22172_new_n3430_));
OR2X2 OR2X2_1491 ( .A(core__abc_22172_new_n3434_), .B(core__abc_22172_new_n3431_), .Y(core__abc_22172_new_n3435_));
OR2X2 OR2X2_1492 ( .A(core__abc_22172_new_n3437_), .B(core__abc_22172_new_n3381_), .Y(core__abc_22172_new_n3438_));
OR2X2 OR2X2_1493 ( .A(core__abc_22172_new_n3438_), .B(core__abc_22172_new_n3436_), .Y(core__abc_22172_new_n3441_));
OR2X2 OR2X2_1494 ( .A(core__abc_22172_new_n3355_), .B(core__abc_22172_new_n2059_), .Y(core__abc_22172_new_n3443_));
OR2X2 OR2X2_1495 ( .A(core__abc_22172_new_n3445_), .B(core__abc_22172_new_n3446_), .Y(core__abc_22172_new_n3447_));
OR2X2 OR2X2_1496 ( .A(core__abc_22172_new_n3451_), .B(core__abc_22172_new_n3448_), .Y(core__abc_22172_new_n3452_));
OR2X2 OR2X2_1497 ( .A(core__abc_22172_new_n3442_), .B(core__abc_22172_new_n3452_), .Y(core__abc_22172_new_n3453_));
OR2X2 OR2X2_1498 ( .A(core__abc_22172_new_n3447_), .B(core_v3_reg_31_), .Y(core__abc_22172_new_n3456_));
OR2X2 OR2X2_1499 ( .A(core__abc_22172_new_n3454_), .B(core__abc_22172_new_n3457_), .Y(core__abc_22172_new_n3458_));
OR2X2 OR2X2_15 ( .A(_abc_19873_new_n945_), .B(_abc_19873_new_n946_), .Y(_abc_19873_new_n947_));
OR2X2 OR2X2_150 ( .A(_abc_19873_new_n1232_), .B(_abc_19873_new_n1233_), .Y(_abc_19873_new_n1234_));
OR2X2 OR2X2_1500 ( .A(core_v3_reg_4_), .B(core_mi_4_), .Y(core__abc_22172_new_n3465_));
OR2X2 OR2X2_1501 ( .A(core__abc_22172_new_n3462_), .B(core__abc_22172_new_n3467_), .Y(core__abc_22172_new_n3468_));
OR2X2 OR2X2_1502 ( .A(core__abc_22172_new_n3217_), .B(core__abc_22172_new_n3468_), .Y(core__abc_22172_new_n3469_));
OR2X2 OR2X2_1503 ( .A(core__abc_22172_new_n3460_), .B(core__abc_22172_new_n3469_), .Y(core__abc_22172_new_n3470_));
OR2X2 OR2X2_1504 ( .A(core__abc_22172_new_n3228_), .B(core_v3_reg_4_), .Y(core__abc_22172_new_n3471_));
OR2X2 OR2X2_1505 ( .A(core__abc_22172_new_n3439_), .B(core__abc_22172_new_n3434_), .Y(core__abc_22172_new_n3474_));
OR2X2 OR2X2_1506 ( .A(core__abc_22172_new_n3419_), .B(core__abc_22172_new_n1885_), .Y(core__abc_22172_new_n3476_));
OR2X2 OR2X2_1507 ( .A(core__abc_22172_new_n3476_), .B(core__abc_22172_new_n1904_), .Y(core__abc_22172_new_n3477_));
OR2X2 OR2X2_1508 ( .A(core__abc_22172_new_n3425_), .B(core__abc_22172_new_n1336_), .Y(core__abc_22172_new_n3482_));
OR2X2 OR2X2_1509 ( .A(core__abc_22172_new_n3484_), .B(core__abc_22172_new_n3485_), .Y(core__abc_22172_new_n3486_));
OR2X2 OR2X2_151 ( .A(_abc_19873_new_n1038_), .B(_abc_19873_new_n1235_), .Y(_abc_19873_new_n1236_));
OR2X2 OR2X2_1510 ( .A(core__abc_22172_new_n3489_), .B(core__abc_22172_new_n3487_), .Y(core__abc_22172_new_n3490_));
OR2X2 OR2X2_1511 ( .A(core__abc_22172_new_n3480_), .B(core__abc_22172_new_n3491_), .Y(core__abc_22172_new_n3494_));
OR2X2 OR2X2_1512 ( .A(core__abc_22172_new_n3475_), .B(core__abc_22172_new_n3495_), .Y(core__abc_22172_new_n3496_));
OR2X2 OR2X2_1513 ( .A(core__abc_22172_new_n3474_), .B(core__abc_22172_new_n3497_), .Y(core__abc_22172_new_n3498_));
OR2X2 OR2X2_1514 ( .A(core__abc_22172_new_n3506_), .B(core__abc_22172_new_n2076_), .Y(core__abc_22172_new_n3507_));
OR2X2 OR2X2_1515 ( .A(core__abc_22172_new_n3505_), .B(core__abc_22172_new_n3507_), .Y(core__abc_22172_new_n3508_));
OR2X2 OR2X2_1516 ( .A(core__abc_22172_new_n3504_), .B(core__abc_22172_new_n3508_), .Y(core__abc_22172_new_n3509_));
OR2X2 OR2X2_1517 ( .A(core__abc_22172_new_n3510_), .B(core__abc_22172_new_n3509_), .Y(core__abc_22172_new_n3511_));
OR2X2 OR2X2_1518 ( .A(core__abc_22172_new_n3513_), .B(core__abc_22172_new_n3514_), .Y(core__abc_22172_new_n3515_));
OR2X2 OR2X2_1519 ( .A(core__abc_22172_new_n3516_), .B(core__abc_22172_new_n3501_), .Y(core__abc_22172_new_n3517_));
OR2X2 OR2X2_152 ( .A(_abc_19873_new_n1236_), .B(_abc_19873_new_n1234_), .Y(_abc_19873_new_n1237_));
OR2X2 OR2X2_1520 ( .A(core__abc_22172_new_n3515_), .B(core_v3_reg_32_), .Y(core__abc_22172_new_n3518_));
OR2X2 OR2X2_1521 ( .A(core__abc_22172_new_n3500_), .B(core__abc_22172_new_n3520_), .Y(core__abc_22172_new_n3521_));
OR2X2 OR2X2_1522 ( .A(core__abc_22172_new_n3499_), .B(core__abc_22172_new_n3519_), .Y(core__abc_22172_new_n3522_));
OR2X2 OR2X2_1523 ( .A(core_v3_reg_5_), .B(core_mi_5_), .Y(core__abc_22172_new_n3529_));
OR2X2 OR2X2_1524 ( .A(core__abc_22172_new_n3526_), .B(core__abc_22172_new_n3531_), .Y(core__abc_22172_new_n3532_));
OR2X2 OR2X2_1525 ( .A(core__abc_22172_new_n3217_), .B(core__abc_22172_new_n3532_), .Y(core__abc_22172_new_n3533_));
OR2X2 OR2X2_1526 ( .A(core__abc_22172_new_n3524_), .B(core__abc_22172_new_n3533_), .Y(core__abc_22172_new_n3534_));
OR2X2 OR2X2_1527 ( .A(core__abc_22172_new_n3228_), .B(core_v3_reg_5_), .Y(core__abc_22172_new_n3535_));
OR2X2 OR2X2_1528 ( .A(core__abc_22172_new_n3539_), .B(core__abc_22172_new_n3538_), .Y(core__abc_22172_new_n3540_));
OR2X2 OR2X2_1529 ( .A(core__abc_22172_new_n3543_), .B(core__abc_22172_new_n3541_), .Y(core__abc_22172_new_n3544_));
OR2X2 OR2X2_153 ( .A(_abc_19873_new_n1239_), .B(_abc_19873_new_n1240_), .Y(_abc_19873_new_n1241_));
OR2X2 OR2X2_1530 ( .A(core__abc_22172_new_n3547_), .B(core__abc_22172_new_n3545_), .Y(core__abc_22172_new_n3548_));
OR2X2 OR2X2_1531 ( .A(core__abc_22172_new_n3059_), .B(core__abc_22172_new_n3550_), .Y(core__abc_22172_new_n3551_));
OR2X2 OR2X2_1532 ( .A(core__abc_22172_new_n3554_), .B(core__abc_22172_new_n3555_), .Y(core__abc_22172_new_n3556_));
OR2X2 OR2X2_1533 ( .A(core__abc_22172_new_n3557_), .B(core__abc_22172_new_n3549_), .Y(core__abc_22172_new_n3558_));
OR2X2 OR2X2_1534 ( .A(core__abc_22172_new_n3556_), .B(core_v3_reg_54_), .Y(core__abc_22172_new_n3559_));
OR2X2 OR2X2_1535 ( .A(core__abc_22172_new_n3564_), .B(core__abc_22172_new_n3561_), .Y(core__abc_22172_new_n3565_));
OR2X2 OR2X2_1536 ( .A(core__abc_22172_new_n3567_), .B(core__abc_22172_new_n3492_), .Y(core__abc_22172_new_n3568_));
OR2X2 OR2X2_1537 ( .A(core__abc_22172_new_n3571_), .B(core__abc_22172_new_n3569_), .Y(core__abc_22172_new_n3572_));
OR2X2 OR2X2_1538 ( .A(core__abc_22172_new_n3580_), .B(core__abc_22172_new_n3578_), .Y(core__abc_22172_new_n3581_));
OR2X2 OR2X2_1539 ( .A(core__abc_22172_new_n3577_), .B(core__abc_22172_new_n3581_), .Y(core__abc_22172_new_n3582_));
OR2X2 OR2X2_154 ( .A(_abc_19873_new_n1241_), .B(_abc_19873_new_n1238_), .Y(_abc_19873_new_n1242_));
OR2X2 OR2X2_1540 ( .A(core__abc_22172_new_n3585_), .B(core__abc_22172_new_n3583_), .Y(core__abc_22172_new_n3586_));
OR2X2 OR2X2_1541 ( .A(core__abc_22172_new_n3573_), .B(core__abc_22172_new_n3587_), .Y(core__abc_22172_new_n3588_));
OR2X2 OR2X2_1542 ( .A(core__abc_22172_new_n3572_), .B(core__abc_22172_new_n3586_), .Y(core__abc_22172_new_n3589_));
OR2X2 OR2X2_1543 ( .A(core_v3_reg_6_), .B(core_mi_6_), .Y(core__abc_22172_new_n3596_));
OR2X2 OR2X2_1544 ( .A(core__abc_22172_new_n3593_), .B(core__abc_22172_new_n3598_), .Y(core__abc_22172_new_n3599_));
OR2X2 OR2X2_1545 ( .A(core__abc_22172_new_n3217_), .B(core__abc_22172_new_n3599_), .Y(core__abc_22172_new_n3600_));
OR2X2 OR2X2_1546 ( .A(core__abc_22172_new_n3591_), .B(core__abc_22172_new_n3600_), .Y(core__abc_22172_new_n3601_));
OR2X2 OR2X2_1547 ( .A(core__abc_22172_new_n3228_), .B(core_v3_reg_6_), .Y(core__abc_22172_new_n3602_));
OR2X2 OR2X2_1548 ( .A(core__abc_22172_new_n3545_), .B(core__abc_22172_new_n1919_), .Y(core__abc_22172_new_n3605_));
OR2X2 OR2X2_1549 ( .A(core__abc_22172_new_n3607_), .B(core__abc_22172_new_n3608_), .Y(core__abc_22172_new_n3609_));
OR2X2 OR2X2_155 ( .A(_abc_19873_new_n1243_), .B(_abc_19873_new_n1244_), .Y(_abc_19873_new_n1245_));
OR2X2 OR2X2_1550 ( .A(core__abc_22172_new_n3554_), .B(core__abc_22172_new_n1374_), .Y(core__abc_22172_new_n3612_));
OR2X2 OR2X2_1551 ( .A(core__abc_22172_new_n3614_), .B(core__abc_22172_new_n3615_), .Y(core__abc_22172_new_n3616_));
OR2X2 OR2X2_1552 ( .A(core__abc_22172_new_n3619_), .B(core__abc_22172_new_n3617_), .Y(core__abc_22172_new_n3620_));
OR2X2 OR2X2_1553 ( .A(core__abc_22172_new_n3610_), .B(core__abc_22172_new_n3621_), .Y(core__abc_22172_new_n3622_));
OR2X2 OR2X2_1554 ( .A(core__abc_22172_new_n3609_), .B(core__abc_22172_new_n3620_), .Y(core__abc_22172_new_n3623_));
OR2X2 OR2X2_1555 ( .A(core__abc_22172_new_n3569_), .B(core__abc_22172_new_n3564_), .Y(core__abc_22172_new_n3626_));
OR2X2 OR2X2_1556 ( .A(core__abc_22172_new_n3628_), .B(core__abc_22172_new_n3629_), .Y(core__abc_22172_new_n3630_));
OR2X2 OR2X2_1557 ( .A(core__abc_22172_new_n3578_), .B(core__abc_22172_new_n2111_), .Y(core__abc_22172_new_n3633_));
OR2X2 OR2X2_1558 ( .A(core__abc_22172_new_n3580_), .B(core__abc_22172_new_n3633_), .Y(core__abc_22172_new_n3634_));
OR2X2 OR2X2_1559 ( .A(core__abc_22172_new_n3636_), .B(core__abc_22172_new_n3637_), .Y(core__abc_22172_new_n3638_));
OR2X2 OR2X2_156 ( .A(_abc_19873_new_n1246_), .B(_abc_19873_new_n1247_), .Y(_abc_19873_new_n1248_));
OR2X2 OR2X2_1560 ( .A(core__abc_22172_new_n3639_), .B(core__abc_22172_new_n3632_), .Y(core__abc_22172_new_n3640_));
OR2X2 OR2X2_1561 ( .A(core__abc_22172_new_n3638_), .B(core_v3_reg_34_), .Y(core__abc_22172_new_n3641_));
OR2X2 OR2X2_1562 ( .A(core__abc_22172_new_n3631_), .B(core__abc_22172_new_n3643_), .Y(core__abc_22172_new_n3644_));
OR2X2 OR2X2_1563 ( .A(core__abc_22172_new_n3630_), .B(core__abc_22172_new_n3642_), .Y(core__abc_22172_new_n3645_));
OR2X2 OR2X2_1564 ( .A(core_v3_reg_7_), .B(core_mi_7_), .Y(core__abc_22172_new_n3651_));
OR2X2 OR2X2_1565 ( .A(core__abc_22172_new_n3648_), .B(core__abc_22172_new_n3653_), .Y(core__abc_22172_new_n3654_));
OR2X2 OR2X2_1566 ( .A(core__abc_22172_new_n3217_), .B(core__abc_22172_new_n3654_), .Y(core__abc_22172_new_n3655_));
OR2X2 OR2X2_1567 ( .A(core__abc_22172_new_n3647_), .B(core__abc_22172_new_n3655_), .Y(core__abc_22172_new_n3656_));
OR2X2 OR2X2_1568 ( .A(core__abc_22172_new_n3228_), .B(core_v3_reg_7_), .Y(core__abc_22172_new_n3657_));
OR2X2 OR2X2_1569 ( .A(core__abc_22172_new_n3665_), .B(core__abc_22172_new_n3664_), .Y(core__abc_22172_new_n3666_));
OR2X2 OR2X2_157 ( .A(_abc_19873_new_n1245_), .B(_abc_19873_new_n1248_), .Y(_abc_19873_new_n1249_));
OR2X2 OR2X2_1570 ( .A(core__abc_22172_new_n3667_), .B(core__abc_22172_new_n3492_), .Y(core__abc_22172_new_n3668_));
OR2X2 OR2X2_1571 ( .A(core__abc_22172_new_n3669_), .B(core__abc_22172_new_n3666_), .Y(core__abc_22172_new_n3670_));
OR2X2 OR2X2_1572 ( .A(core__abc_22172_new_n3670_), .B(core__abc_22172_new_n3663_), .Y(core__abc_22172_new_n3671_));
OR2X2 OR2X2_1573 ( .A(core__abc_22172_new_n3677_), .B(core__abc_22172_new_n1936_), .Y(core__abc_22172_new_n3678_));
OR2X2 OR2X2_1574 ( .A(core__abc_22172_new_n3676_), .B(core__abc_22172_new_n3678_), .Y(core__abc_22172_new_n3679_));
OR2X2 OR2X2_1575 ( .A(core__abc_22172_new_n3675_), .B(core__abc_22172_new_n3679_), .Y(core__abc_22172_new_n3680_));
OR2X2 OR2X2_1576 ( .A(core__abc_22172_new_n3682_), .B(core__abc_22172_new_n3680_), .Y(core__abc_22172_new_n3683_));
OR2X2 OR2X2_1577 ( .A(core__abc_22172_new_n3686_), .B(core__abc_22172_new_n3684_), .Y(core__abc_22172_new_n3687_));
OR2X2 OR2X2_1578 ( .A(core__abc_22172_new_n3691_), .B(core__abc_22172_new_n3692_), .Y(core__abc_22172_new_n3693_));
OR2X2 OR2X2_1579 ( .A(core__abc_22172_new_n3694_), .B(core__abc_22172_new_n3689_), .Y(core__abc_22172_new_n3695_));
OR2X2 OR2X2_158 ( .A(_abc_19873_new_n1249_), .B(_abc_19873_new_n1242_), .Y(_abc_19873_new_n1250_));
OR2X2 OR2X2_1580 ( .A(core__abc_22172_new_n3693_), .B(core_v3_reg_56_), .Y(core__abc_22172_new_n3696_));
OR2X2 OR2X2_1581 ( .A(core__abc_22172_new_n3699_), .B(core__abc_22172_new_n3700_), .Y(core__abc_22172_new_n3701_));
OR2X2 OR2X2_1582 ( .A(core__abc_22172_new_n3702_), .B(core__abc_22172_new_n3704_), .Y(core__abc_22172_new_n3705_));
OR2X2 OR2X2_1583 ( .A(core__abc_22172_new_n3637_), .B(core__abc_22172_new_n2127_), .Y(core__abc_22172_new_n3707_));
OR2X2 OR2X2_1584 ( .A(core__abc_22172_new_n3707_), .B(core__abc_22172_new_n2146_), .Y(core__abc_22172_new_n3708_));
OR2X2 OR2X2_1585 ( .A(core__abc_22172_new_n3712_), .B(core_v3_reg_35_), .Y(core__abc_22172_new_n3715_));
OR2X2 OR2X2_1586 ( .A(core__abc_22172_new_n3706_), .B(core__abc_22172_new_n3717_), .Y(core__abc_22172_new_n3718_));
OR2X2 OR2X2_1587 ( .A(core__abc_22172_new_n3705_), .B(core__abc_22172_new_n3716_), .Y(core__abc_22172_new_n3719_));
OR2X2 OR2X2_1588 ( .A(core_v3_reg_8_), .B(core_mi_8_), .Y(core__abc_22172_new_n3726_));
OR2X2 OR2X2_1589 ( .A(core__abc_22172_new_n3723_), .B(core__abc_22172_new_n3728_), .Y(core__abc_22172_new_n3729_));
OR2X2 OR2X2_159 ( .A(_abc_19873_new_n1250_), .B(_abc_19873_new_n1237_), .Y(_abc_19873_new_n1251_));
OR2X2 OR2X2_1590 ( .A(core__abc_22172_new_n3217_), .B(core__abc_22172_new_n3729_), .Y(core__abc_22172_new_n3730_));
OR2X2 OR2X2_1591 ( .A(core__abc_22172_new_n3721_), .B(core__abc_22172_new_n3730_), .Y(core__abc_22172_new_n3731_));
OR2X2 OR2X2_1592 ( .A(core__abc_22172_new_n3228_), .B(core_v3_reg_8_), .Y(core__abc_22172_new_n3732_));
OR2X2 OR2X2_1593 ( .A(core__abc_22172_new_n3738_), .B(core__abc_22172_new_n1978_), .Y(core__abc_22172_new_n3741_));
OR2X2 OR2X2_1594 ( .A(core__abc_22172_new_n3692_), .B(core__abc_22172_new_n1412_), .Y(core__abc_22172_new_n3744_));
OR2X2 OR2X2_1595 ( .A(core__abc_22172_new_n3746_), .B(core__abc_22172_new_n3747_), .Y(core__abc_22172_new_n3748_));
OR2X2 OR2X2_1596 ( .A(core__abc_22172_new_n3751_), .B(core__abc_22172_new_n3749_), .Y(core__abc_22172_new_n3752_));
OR2X2 OR2X2_1597 ( .A(core__abc_22172_new_n3742_), .B(core__abc_22172_new_n3753_), .Y(core__abc_22172_new_n3756_));
OR2X2 OR2X2_1598 ( .A(core__abc_22172_new_n3774_), .B(core__abc_22172_new_n2144_), .Y(core__abc_22172_new_n3775_));
OR2X2 OR2X2_1599 ( .A(core__abc_22172_new_n3773_), .B(core__abc_22172_new_n3775_), .Y(core__abc_22172_new_n3776_));
OR2X2 OR2X2_16 ( .A(_abc_19873_new_n944_), .B(_abc_19873_new_n947_), .Y(_abc_19873_new_n948_));
OR2X2 OR2X2_160 ( .A(_abc_19873_new_n1253_), .B(_abc_19873_new_n1254_), .Y(_abc_19873_new_n1255_));
OR2X2 OR2X2_1600 ( .A(core__abc_22172_new_n3772_), .B(core__abc_22172_new_n3776_), .Y(core__abc_22172_new_n3777_));
OR2X2 OR2X2_1601 ( .A(core__abc_22172_new_n3779_), .B(core__abc_22172_new_n3780_), .Y(core__abc_22172_new_n3781_));
OR2X2 OR2X2_1602 ( .A(core__abc_22172_new_n3782_), .B(core__abc_22172_new_n3769_), .Y(core__abc_22172_new_n3783_));
OR2X2 OR2X2_1603 ( .A(core__abc_22172_new_n3781_), .B(core_v3_reg_36_), .Y(core__abc_22172_new_n3784_));
OR2X2 OR2X2_1604 ( .A(core__abc_22172_new_n3768_), .B(core__abc_22172_new_n3786_), .Y(core__abc_22172_new_n3787_));
OR2X2 OR2X2_1605 ( .A(core__abc_22172_new_n3788_), .B(core__abc_22172_new_n3785_), .Y(core__abc_22172_new_n3789_));
OR2X2 OR2X2_1606 ( .A(core_v3_reg_9_), .B(core_mi_9_), .Y(core__abc_22172_new_n3795_));
OR2X2 OR2X2_1607 ( .A(core__abc_22172_new_n3792_), .B(core__abc_22172_new_n3797_), .Y(core__abc_22172_new_n3798_));
OR2X2 OR2X2_1608 ( .A(core__abc_22172_new_n3217_), .B(core__abc_22172_new_n3798_), .Y(core__abc_22172_new_n3799_));
OR2X2 OR2X2_1609 ( .A(core__abc_22172_new_n3791_), .B(core__abc_22172_new_n3799_), .Y(core__abc_22172_new_n3800_));
OR2X2 OR2X2_161 ( .A(_abc_19873_new_n1257_), .B(_abc_19873_new_n1258_), .Y(_abc_19873_new_n1259_));
OR2X2 OR2X2_1610 ( .A(core__abc_22172_new_n3228_), .B(core_v3_reg_9_), .Y(core__abc_22172_new_n3801_));
OR2X2 OR2X2_1611 ( .A(core__abc_22172_new_n3762_), .B(core__abc_22172_new_n3754_), .Y(core__abc_22172_new_n3804_));
OR2X2 OR2X2_1612 ( .A(core__abc_22172_new_n3811_), .B(core__abc_22172_new_n3810_), .Y(core__abc_22172_new_n3812_));
OR2X2 OR2X2_1613 ( .A(core__abc_22172_new_n3809_), .B(core__abc_22172_new_n3813_), .Y(core__abc_22172_new_n3814_));
OR2X2 OR2X2_1614 ( .A(core__abc_22172_new_n3817_), .B(core__abc_22172_new_n3815_), .Y(core__abc_22172_new_n3818_));
OR2X2 OR2X2_1615 ( .A(core__abc_22172_new_n3822_), .B(core__abc_22172_new_n1452_), .Y(core__abc_22172_new_n3824_));
OR2X2 OR2X2_1616 ( .A(core__abc_22172_new_n3825_), .B(core__abc_22172_new_n3823_), .Y(core__abc_22172_new_n3826_));
OR2X2 OR2X2_1617 ( .A(core__abc_22172_new_n3827_), .B(core__abc_22172_new_n3819_), .Y(core__abc_22172_new_n3828_));
OR2X2 OR2X2_1618 ( .A(core__abc_22172_new_n3826_), .B(core_v3_reg_58_), .Y(core__abc_22172_new_n3829_));
OR2X2 OR2X2_1619 ( .A(core__abc_22172_new_n3834_), .B(core__abc_22172_new_n3831_), .Y(core__abc_22172_new_n3835_));
OR2X2 OR2X2_162 ( .A(_abc_19873_new_n1259_), .B(_abc_19873_new_n1256_), .Y(_abc_19873_new_n1260_));
OR2X2 OR2X2_1620 ( .A(core__abc_22172_new_n3837_), .B(core__abc_22172_new_n3838_), .Y(core__abc_22172_new_n3839_));
OR2X2 OR2X2_1621 ( .A(core__abc_22172_new_n3780_), .B(core__abc_22172_new_n2161_), .Y(core__abc_22172_new_n3841_));
OR2X2 OR2X2_1622 ( .A(core__abc_22172_new_n3843_), .B(core__abc_22172_new_n3844_), .Y(core__abc_22172_new_n3845_));
OR2X2 OR2X2_1623 ( .A(core__abc_22172_new_n3845_), .B(core_v3_reg_37_), .Y(core__abc_22172_new_n3846_));
OR2X2 OR2X2_1624 ( .A(core__abc_22172_new_n3840_), .B(core__abc_22172_new_n3850_), .Y(core__abc_22172_new_n3851_));
OR2X2 OR2X2_1625 ( .A(core__abc_22172_new_n3839_), .B(core__abc_22172_new_n3849_), .Y(core__abc_22172_new_n3852_));
OR2X2 OR2X2_1626 ( .A(core_v3_reg_10_), .B(core_mi_10_), .Y(core__abc_22172_new_n3859_));
OR2X2 OR2X2_1627 ( .A(core__abc_22172_new_n3856_), .B(core__abc_22172_new_n3861_), .Y(core__abc_22172_new_n3862_));
OR2X2 OR2X2_1628 ( .A(core__abc_22172_new_n3217_), .B(core__abc_22172_new_n3862_), .Y(core__abc_22172_new_n3863_));
OR2X2 OR2X2_1629 ( .A(core__abc_22172_new_n3854_), .B(core__abc_22172_new_n3863_), .Y(core__abc_22172_new_n3864_));
OR2X2 OR2X2_163 ( .A(_abc_19873_new_n1260_), .B(_abc_19873_new_n1255_), .Y(_abc_19873_new_n1261_));
OR2X2 OR2X2_1630 ( .A(core__abc_22172_new_n3228_), .B(core_v3_reg_10_), .Y(core__abc_22172_new_n3865_));
OR2X2 OR2X2_1631 ( .A(core__abc_22172_new_n3837_), .B(core__abc_22172_new_n3834_), .Y(core__abc_22172_new_n3868_));
OR2X2 OR2X2_1632 ( .A(core__abc_22172_new_n3815_), .B(core__abc_22172_new_n1987_), .Y(core__abc_22172_new_n3870_));
OR2X2 OR2X2_1633 ( .A(core__abc_22172_new_n3872_), .B(core__abc_22172_new_n3873_), .Y(core__abc_22172_new_n3874_));
OR2X2 OR2X2_1634 ( .A(core__abc_22172_new_n3876_), .B(core__abc_22172_new_n1469_), .Y(core__abc_22172_new_n3879_));
OR2X2 OR2X2_1635 ( .A(core__abc_22172_new_n3881_), .B(core_v3_reg_59_), .Y(core__abc_22172_new_n3884_));
OR2X2 OR2X2_1636 ( .A(core__abc_22172_new_n3875_), .B(core__abc_22172_new_n3886_), .Y(core__abc_22172_new_n3887_));
OR2X2 OR2X2_1637 ( .A(core__abc_22172_new_n3874_), .B(core__abc_22172_new_n3885_), .Y(core__abc_22172_new_n3888_));
OR2X2 OR2X2_1638 ( .A(core__abc_22172_new_n3891_), .B(core__abc_22172_new_n3892_), .Y(core__abc_22172_new_n3893_));
OR2X2 OR2X2_1639 ( .A(core__abc_22172_new_n3898_), .B(core__abc_22172_new_n2179_), .Y(core__abc_22172_new_n3899_));
OR2X2 OR2X2_164 ( .A(_abc_19873_new_n1263_), .B(_abc_19873_new_n1264_), .Y(_abc_19873_new_n1265_));
OR2X2 OR2X2_1640 ( .A(core__abc_22172_new_n3897_), .B(core__abc_22172_new_n3899_), .Y(core__abc_22172_new_n3900_));
OR2X2 OR2X2_1641 ( .A(core__abc_22172_new_n3903_), .B(core__abc_22172_new_n3901_), .Y(core__abc_22172_new_n3904_));
OR2X2 OR2X2_1642 ( .A(core__abc_22172_new_n3905_), .B(core__abc_22172_new_n3895_), .Y(core__abc_22172_new_n3906_));
OR2X2 OR2X2_1643 ( .A(core__abc_22172_new_n3904_), .B(core_v3_reg_38_), .Y(core__abc_22172_new_n3907_));
OR2X2 OR2X2_1644 ( .A(core__abc_22172_new_n3894_), .B(core__abc_22172_new_n3909_), .Y(core__abc_22172_new_n3910_));
OR2X2 OR2X2_1645 ( .A(core__abc_22172_new_n3893_), .B(core__abc_22172_new_n3908_), .Y(core__abc_22172_new_n3911_));
OR2X2 OR2X2_1646 ( .A(core_v3_reg_11_), .B(core_mi_11_), .Y(core__abc_22172_new_n3917_));
OR2X2 OR2X2_1647 ( .A(core__abc_22172_new_n3914_), .B(core__abc_22172_new_n3919_), .Y(core__abc_22172_new_n3920_));
OR2X2 OR2X2_1648 ( .A(core__abc_22172_new_n3217_), .B(core__abc_22172_new_n3920_), .Y(core__abc_22172_new_n3921_));
OR2X2 OR2X2_1649 ( .A(core__abc_22172_new_n3913_), .B(core__abc_22172_new_n3921_), .Y(core__abc_22172_new_n3922_));
OR2X2 OR2X2_165 ( .A(_abc_19873_new_n1266_), .B(_abc_19873_new_n1267_), .Y(_abc_19873_new_n1268_));
OR2X2 OR2X2_1650 ( .A(core__abc_22172_new_n3228_), .B(core_v3_reg_11_), .Y(core__abc_22172_new_n3923_));
OR2X2 OR2X2_1651 ( .A(core__abc_22172_new_n3929_), .B(core__abc_22172_new_n3928_), .Y(core__abc_22172_new_n3930_));
OR2X2 OR2X2_1652 ( .A(core__abc_22172_new_n3927_), .B(core__abc_22172_new_n3930_), .Y(core__abc_22172_new_n3931_));
OR2X2 OR2X2_1653 ( .A(core__abc_22172_new_n3933_), .B(core__abc_22172_new_n3931_), .Y(core__abc_22172_new_n3934_));
OR2X2 OR2X2_1654 ( .A(core__abc_22172_new_n3937_), .B(core__abc_22172_new_n2004_), .Y(core__abc_22172_new_n3938_));
OR2X2 OR2X2_1655 ( .A(core__abc_22172_new_n3936_), .B(core__abc_22172_new_n3938_), .Y(core__abc_22172_new_n3939_));
OR2X2 OR2X2_1656 ( .A(core__abc_22172_new_n3941_), .B(core__abc_22172_new_n3939_), .Y(core__abc_22172_new_n3942_));
OR2X2 OR2X2_1657 ( .A(core__abc_22172_new_n3945_), .B(core__abc_22172_new_n3943_), .Y(core__abc_22172_new_n3946_));
OR2X2 OR2X2_1658 ( .A(core__abc_22172_new_n3948_), .B(core__abc_22172_new_n3089_), .Y(core__abc_22172_new_n3949_));
OR2X2 OR2X2_1659 ( .A(core__abc_22172_new_n3952_), .B(core__abc_22172_new_n3950_), .Y(core__abc_22172_new_n3953_));
OR2X2 OR2X2_166 ( .A(_abc_19873_new_n1265_), .B(_abc_19873_new_n1268_), .Y(_abc_19873_new_n1269_));
OR2X2 OR2X2_1660 ( .A(core__abc_22172_new_n3954_), .B(core__abc_22172_new_n3947_), .Y(core__abc_22172_new_n3955_));
OR2X2 OR2X2_1661 ( .A(core__abc_22172_new_n3953_), .B(core_v3_reg_60_), .Y(core__abc_22172_new_n3956_));
OR2X2 OR2X2_1662 ( .A(core__abc_22172_new_n3961_), .B(core__abc_22172_new_n3958_), .Y(core__abc_22172_new_n3962_));
OR2X2 OR2X2_1663 ( .A(core__abc_22172_new_n3934_), .B(core__abc_22172_new_n3963_), .Y(core__abc_22172_new_n3966_));
OR2X2 OR2X2_1664 ( .A(core__abc_22172_new_n3901_), .B(core__abc_22172_new_n2195_), .Y(core__abc_22172_new_n3968_));
OR2X2 OR2X2_1665 ( .A(core__abc_22172_new_n3970_), .B(core__abc_22172_new_n3971_), .Y(core__abc_22172_new_n3972_));
OR2X2 OR2X2_1666 ( .A(core__abc_22172_new_n3972_), .B(core_v3_reg_39_), .Y(core__abc_22172_new_n3974_));
OR2X2 OR2X2_1667 ( .A(core__abc_22172_new_n3975_), .B(core__abc_22172_new_n3973_), .Y(core__abc_22172_new_n3976_));
OR2X2 OR2X2_1668 ( .A(core__abc_22172_new_n3967_), .B(core__abc_22172_new_n3976_), .Y(core__abc_22172_new_n3977_));
OR2X2 OR2X2_1669 ( .A(core__abc_22172_new_n3978_), .B(core__abc_22172_new_n3980_), .Y(core__abc_22172_new_n3981_));
OR2X2 OR2X2_167 ( .A(_abc_19873_new_n1269_), .B(_abc_19873_new_n1262_), .Y(_abc_19873_new_n1270_));
OR2X2 OR2X2_1670 ( .A(core_v3_reg_12_), .B(core_mi_12_), .Y(core__abc_22172_new_n3987_));
OR2X2 OR2X2_1671 ( .A(core__abc_22172_new_n3984_), .B(core__abc_22172_new_n3989_), .Y(core__abc_22172_new_n3990_));
OR2X2 OR2X2_1672 ( .A(core__abc_22172_new_n3217_), .B(core__abc_22172_new_n3990_), .Y(core__abc_22172_new_n3991_));
OR2X2 OR2X2_1673 ( .A(core__abc_22172_new_n3983_), .B(core__abc_22172_new_n3991_), .Y(core__abc_22172_new_n3992_));
OR2X2 OR2X2_1674 ( .A(core__abc_22172_new_n3228_), .B(core_v3_reg_12_), .Y(core__abc_22172_new_n3993_));
OR2X2 OR2X2_1675 ( .A(core__abc_22172_new_n3943_), .B(core__abc_22172_new_n2021_), .Y(core__abc_22172_new_n3997_));
OR2X2 OR2X2_1676 ( .A(core__abc_22172_new_n3999_), .B(core__abc_22172_new_n4000_), .Y(core__abc_22172_new_n4001_));
OR2X2 OR2X2_1677 ( .A(core__abc_22172_new_n3950_), .B(core__abc_22172_new_n1480_), .Y(core__abc_22172_new_n4004_));
OR2X2 OR2X2_1678 ( .A(core__abc_22172_new_n4006_), .B(core__abc_22172_new_n4007_), .Y(core__abc_22172_new_n4008_));
OR2X2 OR2X2_1679 ( .A(core__abc_22172_new_n4011_), .B(core__abc_22172_new_n4009_), .Y(core__abc_22172_new_n4012_));
OR2X2 OR2X2_168 ( .A(_abc_19873_new_n1270_), .B(_abc_19873_new_n1261_), .Y(_abc_19873_new_n1271_));
OR2X2 OR2X2_1680 ( .A(core__abc_22172_new_n4002_), .B(core__abc_22172_new_n4013_), .Y(core__abc_22172_new_n4014_));
OR2X2 OR2X2_1681 ( .A(core__abc_22172_new_n4001_), .B(core__abc_22172_new_n4012_), .Y(core__abc_22172_new_n4015_));
OR2X2 OR2X2_1682 ( .A(core__abc_22172_new_n4029_), .B(core__abc_22172_new_n2212_), .Y(core__abc_22172_new_n4030_));
OR2X2 OR2X2_1683 ( .A(core__abc_22172_new_n4032_), .B(core__abc_22172_new_n4030_), .Y(core__abc_22172_new_n4033_));
OR2X2 OR2X2_1684 ( .A(core__abc_22172_new_n4034_), .B(core__abc_22172_new_n4033_), .Y(core__abc_22172_new_n4035_));
OR2X2 OR2X2_1685 ( .A(core__abc_22172_new_n4038_), .B(core__abc_22172_new_n4036_), .Y(core__abc_22172_new_n4039_));
OR2X2 OR2X2_1686 ( .A(core__abc_22172_new_n4040_), .B(core_v3_reg_40_), .Y(core__abc_22172_new_n4041_));
OR2X2 OR2X2_1687 ( .A(core__abc_22172_new_n4039_), .B(core__abc_22172_new_n4042_), .Y(core__abc_22172_new_n4043_));
OR2X2 OR2X2_1688 ( .A(core__abc_22172_new_n4028_), .B(core__abc_22172_new_n4045_), .Y(core__abc_22172_new_n4046_));
OR2X2 OR2X2_1689 ( .A(core__abc_22172_new_n4027_), .B(core__abc_22172_new_n4044_), .Y(core__abc_22172_new_n4047_));
OR2X2 OR2X2_169 ( .A(_abc_19873_new_n1273_), .B(_abc_19873_new_n1274_), .Y(_abc_19873_new_n1275_));
OR2X2 OR2X2_1690 ( .A(core_v3_reg_13_), .B(core_mi_13_), .Y(core__abc_22172_new_n4054_));
OR2X2 OR2X2_1691 ( .A(core__abc_22172_new_n4051_), .B(core__abc_22172_new_n4056_), .Y(core__abc_22172_new_n4057_));
OR2X2 OR2X2_1692 ( .A(core__abc_22172_new_n3217_), .B(core__abc_22172_new_n4057_), .Y(core__abc_22172_new_n4058_));
OR2X2 OR2X2_1693 ( .A(core__abc_22172_new_n4049_), .B(core__abc_22172_new_n4058_), .Y(core__abc_22172_new_n4059_));
OR2X2 OR2X2_1694 ( .A(core__abc_22172_new_n3228_), .B(core_v3_reg_13_), .Y(core__abc_22172_new_n4060_));
OR2X2 OR2X2_1695 ( .A(core__abc_22172_new_n4021_), .B(core__abc_22172_new_n4063_), .Y(core__abc_22172_new_n4064_));
OR2X2 OR2X2_1696 ( .A(core__abc_22172_new_n4069_), .B(core__abc_22172_new_n4068_), .Y(core__abc_22172_new_n4070_));
OR2X2 OR2X2_1697 ( .A(core__abc_22172_new_n4073_), .B(core__abc_22172_new_n4071_), .Y(core__abc_22172_new_n4074_));
OR2X2 OR2X2_1698 ( .A(core__abc_22172_new_n4077_), .B(core__abc_22172_new_n4075_), .Y(core__abc_22172_new_n4078_));
OR2X2 OR2X2_1699 ( .A(core__abc_22172_new_n4080_), .B(core__abc_22172_new_n3093_), .Y(core__abc_22172_new_n4081_));
OR2X2 OR2X2_17 ( .A(_abc_19873_new_n948_), .B(_abc_19873_new_n941_), .Y(_abc_19873_new_n949_));
OR2X2 OR2X2_170 ( .A(_abc_19873_new_n1038_), .B(_abc_19873_new_n1276_), .Y(_abc_19873_new_n1277_));
OR2X2 OR2X2_1700 ( .A(core__abc_22172_new_n4083_), .B(core__abc_22172_new_n4084_), .Y(core__abc_22172_new_n4085_));
OR2X2 OR2X2_1701 ( .A(core__abc_22172_new_n4086_), .B(core__abc_22172_new_n4079_), .Y(core__abc_22172_new_n4087_));
OR2X2 OR2X2_1702 ( .A(core__abc_22172_new_n4085_), .B(core_v3_reg_62_), .Y(core__abc_22172_new_n4088_));
OR2X2 OR2X2_1703 ( .A(core__abc_22172_new_n4078_), .B(core__abc_22172_new_n4089_), .Y(core__abc_22172_new_n4092_));
OR2X2 OR2X2_1704 ( .A(core__abc_22172_new_n4094_), .B(core__abc_22172_new_n4096_), .Y(core__abc_22172_new_n4097_));
OR2X2 OR2X2_1705 ( .A(core__abc_22172_new_n4036_), .B(core__abc_22172_new_n2229_), .Y(core__abc_22172_new_n4099_));
OR2X2 OR2X2_1706 ( .A(core__abc_22172_new_n4101_), .B(core__abc_22172_new_n4102_), .Y(core__abc_22172_new_n4103_));
OR2X2 OR2X2_1707 ( .A(core__abc_22172_new_n4105_), .B(core__abc_22172_new_n4107_), .Y(core__abc_22172_new_n4108_));
OR2X2 OR2X2_1708 ( .A(core__abc_22172_new_n4098_), .B(core__abc_22172_new_n4109_), .Y(core__abc_22172_new_n4110_));
OR2X2 OR2X2_1709 ( .A(core__abc_22172_new_n4097_), .B(core__abc_22172_new_n4108_), .Y(core__abc_22172_new_n4111_));
OR2X2 OR2X2_171 ( .A(_abc_19873_new_n1277_), .B(_abc_19873_new_n1275_), .Y(_abc_19873_new_n1278_));
OR2X2 OR2X2_1710 ( .A(core_v3_reg_14_), .B(core_mi_14_), .Y(core__abc_22172_new_n4118_));
OR2X2 OR2X2_1711 ( .A(core__abc_22172_new_n4115_), .B(core__abc_22172_new_n4120_), .Y(core__abc_22172_new_n4121_));
OR2X2 OR2X2_1712 ( .A(core__abc_22172_new_n3217_), .B(core__abc_22172_new_n4121_), .Y(core__abc_22172_new_n4122_));
OR2X2 OR2X2_1713 ( .A(core__abc_22172_new_n4113_), .B(core__abc_22172_new_n4122_), .Y(core__abc_22172_new_n4123_));
OR2X2 OR2X2_1714 ( .A(core__abc_22172_new_n3228_), .B(core_v3_reg_14_), .Y(core__abc_22172_new_n4124_));
OR2X2 OR2X2_1715 ( .A(core__abc_22172_new_n4094_), .B(core__abc_22172_new_n4127_), .Y(core__abc_22172_new_n4128_));
OR2X2 OR2X2_1716 ( .A(core__abc_22172_new_n4075_), .B(core__abc_22172_new_n2055_), .Y(core__abc_22172_new_n4130_));
OR2X2 OR2X2_1717 ( .A(core__abc_22172_new_n4130_), .B(core__abc_22172_new_n2074_), .Y(core__abc_22172_new_n4131_));
OR2X2 OR2X2_1718 ( .A(core__abc_22172_new_n4084_), .B(core__abc_22172_new_n1514_), .Y(core__abc_22172_new_n4135_));
OR2X2 OR2X2_1719 ( .A(core__abc_22172_new_n4137_), .B(core__abc_22172_new_n4138_), .Y(core__abc_22172_new_n4139_));
OR2X2 OR2X2_172 ( .A(_abc_19873_new_n1280_), .B(_abc_19873_new_n1281_), .Y(_abc_19873_new_n1282_));
OR2X2 OR2X2_1720 ( .A(core__abc_22172_new_n4139_), .B(core_v3_reg_63_), .Y(core__abc_22172_new_n4142_));
OR2X2 OR2X2_1721 ( .A(core__abc_22172_new_n4134_), .B(core__abc_22172_new_n4144_), .Y(core__abc_22172_new_n4145_));
OR2X2 OR2X2_1722 ( .A(core__abc_22172_new_n4146_), .B(core__abc_22172_new_n4132_), .Y(core__abc_22172_new_n4147_));
OR2X2 OR2X2_1723 ( .A(core__abc_22172_new_n4147_), .B(core__abc_22172_new_n4143_), .Y(core__abc_22172_new_n4148_));
OR2X2 OR2X2_1724 ( .A(core__abc_22172_new_n4151_), .B(core__abc_22172_new_n4152_), .Y(core__abc_22172_new_n4153_));
OR2X2 OR2X2_1725 ( .A(core__abc_22172_new_n4158_), .B(core__abc_22172_new_n2246_), .Y(core__abc_22172_new_n4159_));
OR2X2 OR2X2_1726 ( .A(core__abc_22172_new_n4157_), .B(core__abc_22172_new_n4159_), .Y(core__abc_22172_new_n4160_));
OR2X2 OR2X2_1727 ( .A(core__abc_22172_new_n4162_), .B(core__abc_22172_new_n4163_), .Y(core__abc_22172_new_n4164_));
OR2X2 OR2X2_1728 ( .A(core__abc_22172_new_n4165_), .B(core__abc_22172_new_n4155_), .Y(core__abc_22172_new_n4166_));
OR2X2 OR2X2_1729 ( .A(core__abc_22172_new_n4164_), .B(core_v3_reg_42_), .Y(core__abc_22172_new_n4167_));
OR2X2 OR2X2_173 ( .A(_abc_19873_new_n1282_), .B(_abc_19873_new_n1279_), .Y(_abc_19873_new_n1283_));
OR2X2 OR2X2_1730 ( .A(core__abc_22172_new_n4154_), .B(core__abc_22172_new_n4169_), .Y(core__abc_22172_new_n4170_));
OR2X2 OR2X2_1731 ( .A(core__abc_22172_new_n4153_), .B(core__abc_22172_new_n4168_), .Y(core__abc_22172_new_n4171_));
OR2X2 OR2X2_1732 ( .A(core_v3_reg_15_), .B(core_mi_15_), .Y(core__abc_22172_new_n4177_));
OR2X2 OR2X2_1733 ( .A(core__abc_22172_new_n4174_), .B(core__abc_22172_new_n4179_), .Y(core__abc_22172_new_n4180_));
OR2X2 OR2X2_1734 ( .A(core__abc_22172_new_n3217_), .B(core__abc_22172_new_n4180_), .Y(core__abc_22172_new_n4181_));
OR2X2 OR2X2_1735 ( .A(core__abc_22172_new_n4173_), .B(core__abc_22172_new_n4181_), .Y(core__abc_22172_new_n4182_));
OR2X2 OR2X2_1736 ( .A(core__abc_22172_new_n3228_), .B(core_v3_reg_15_), .Y(core__abc_22172_new_n4183_));
OR2X2 OR2X2_1737 ( .A(core__abc_22172_new_n4195_), .B(core__abc_22172_new_n4194_), .Y(core__abc_22172_new_n4196_));
OR2X2 OR2X2_1738 ( .A(core__abc_22172_new_n4193_), .B(core__abc_22172_new_n4196_), .Y(core__abc_22172_new_n4197_));
OR2X2 OR2X2_1739 ( .A(core__abc_22172_new_n4197_), .B(core__abc_22172_new_n4192_), .Y(core__abc_22172_new_n4198_));
OR2X2 OR2X2_174 ( .A(_abc_19873_new_n1284_), .B(_abc_19873_new_n1285_), .Y(_abc_19873_new_n1286_));
OR2X2 OR2X2_1740 ( .A(core__abc_22172_new_n4198_), .B(core__abc_22172_new_n4191_), .Y(core__abc_22172_new_n4199_));
OR2X2 OR2X2_1741 ( .A(core__abc_22172_new_n4206_), .B(core__abc_22172_new_n2072_), .Y(core__abc_22172_new_n4207_));
OR2X2 OR2X2_1742 ( .A(core__abc_22172_new_n4205_), .B(core__abc_22172_new_n4207_), .Y(core__abc_22172_new_n4208_));
OR2X2 OR2X2_1743 ( .A(core__abc_22172_new_n4204_), .B(core__abc_22172_new_n4208_), .Y(core__abc_22172_new_n4209_));
OR2X2 OR2X2_1744 ( .A(core__abc_22172_new_n4203_), .B(core__abc_22172_new_n4209_), .Y(core__abc_22172_new_n4210_));
OR2X2 OR2X2_1745 ( .A(core__abc_22172_new_n4212_), .B(core__abc_22172_new_n4210_), .Y(core__abc_22172_new_n4213_));
OR2X2 OR2X2_1746 ( .A(core__abc_22172_new_n3032_), .B(core__abc_22172_new_n4216_), .Y(core__abc_22172_new_n4217_));
OR2X2 OR2X2_1747 ( .A(core__abc_22172_new_n4219_), .B(core__abc_22172_new_n4214_), .Y(core__abc_22172_new_n4220_));
OR2X2 OR2X2_1748 ( .A(core__abc_22172_new_n4222_), .B(core__abc_22172_new_n4223_), .Y(core__abc_22172_new_n4224_));
OR2X2 OR2X2_1749 ( .A(core__abc_22172_new_n4225_), .B(core_v3_reg_0_), .Y(core__abc_22172_new_n4226_));
OR2X2 OR2X2_175 ( .A(_abc_19873_new_n1287_), .B(_abc_19873_new_n1288_), .Y(_abc_19873_new_n1289_));
OR2X2 OR2X2_1750 ( .A(core__abc_22172_new_n4224_), .B(core__abc_22172_new_n1262_), .Y(core__abc_22172_new_n4227_));
OR2X2 OR2X2_1751 ( .A(core__abc_22172_new_n4232_), .B(core__abc_22172_new_n4230_), .Y(core__abc_22172_new_n4233_));
OR2X2 OR2X2_1752 ( .A(core__abc_22172_new_n4237_), .B(core__abc_22172_new_n4235_), .Y(core__abc_22172_new_n4238_));
OR2X2 OR2X2_1753 ( .A(core__abc_22172_new_n4241_), .B(core__abc_22172_new_n2285_), .Y(core__abc_22172_new_n4243_));
OR2X2 OR2X2_1754 ( .A(core__abc_22172_new_n4244_), .B(core__abc_22172_new_n4242_), .Y(core__abc_22172_new_n4245_));
OR2X2 OR2X2_1755 ( .A(core__abc_22172_new_n4246_), .B(core__abc_22172_new_n4250_), .Y(core__abc_22172_new_n4251_));
OR2X2 OR2X2_1756 ( .A(core__abc_22172_new_n4239_), .B(core__abc_22172_new_n4251_), .Y(core__abc_22172_new_n4252_));
OR2X2 OR2X2_1757 ( .A(core__abc_22172_new_n4249_), .B(core__abc_22172_new_n4247_), .Y(core__abc_22172_new_n4253_));
OR2X2 OR2X2_1758 ( .A(core__abc_22172_new_n4238_), .B(core__abc_22172_new_n4255_), .Y(core__abc_22172_new_n4256_));
OR2X2 OR2X2_1759 ( .A(core_v3_reg_16_), .B(core_mi_16_), .Y(core__abc_22172_new_n4260_));
OR2X2 OR2X2_176 ( .A(_abc_19873_new_n1286_), .B(_abc_19873_new_n1289_), .Y(_abc_19873_new_n1290_));
OR2X2 OR2X2_1760 ( .A(core__abc_22172_new_n4259_), .B(core__abc_22172_new_n4264_), .Y(core__abc_22172_new_n4265_));
OR2X2 OR2X2_1761 ( .A(core__abc_22172_new_n4258_), .B(core__abc_22172_new_n4265_), .Y(core__abc_22172_new_n4266_));
OR2X2 OR2X2_1762 ( .A(core__abc_22172_new_n4267_), .B(core__abc_22172_new_n4186_), .Y(core__abc_22172_new_n4268_));
OR2X2 OR2X2_1763 ( .A(core__abc_22172_new_n4218_), .B(core__abc_22172_new_n4279_), .Y(core__abc_22172_new_n4280_));
OR2X2 OR2X2_1764 ( .A(core__abc_22172_new_n4223_), .B(core__abc_22172_new_n1548_), .Y(core__abc_22172_new_n4283_));
OR2X2 OR2X2_1765 ( .A(core__abc_22172_new_n4285_), .B(core__abc_22172_new_n4286_), .Y(core__abc_22172_new_n4287_));
OR2X2 OR2X2_1766 ( .A(core__abc_22172_new_n4290_), .B(core__abc_22172_new_n4288_), .Y(core__abc_22172_new_n4291_));
OR2X2 OR2X2_1767 ( .A(core__abc_22172_new_n4282_), .B(core__abc_22172_new_n4291_), .Y(core__abc_22172_new_n4294_));
OR2X2 OR2X2_1768 ( .A(core__abc_22172_new_n4309_), .B(core__abc_22172_new_n2280_), .Y(core__abc_22172_new_n4310_));
OR2X2 OR2X2_1769 ( .A(core__abc_22172_new_n4308_), .B(core__abc_22172_new_n4310_), .Y(core__abc_22172_new_n4311_));
OR2X2 OR2X2_177 ( .A(_abc_19873_new_n1290_), .B(_abc_19873_new_n1283_), .Y(_abc_19873_new_n1291_));
OR2X2 OR2X2_1770 ( .A(core__abc_22172_new_n4314_), .B(core__abc_22172_new_n4312_), .Y(core__abc_22172_new_n4315_));
OR2X2 OR2X2_1771 ( .A(core__abc_22172_new_n4316_), .B(core_v3_reg_44_), .Y(core__abc_22172_new_n4317_));
OR2X2 OR2X2_1772 ( .A(core__abc_22172_new_n4315_), .B(core__abc_22172_new_n4318_), .Y(core__abc_22172_new_n4319_));
OR2X2 OR2X2_1773 ( .A(core__abc_22172_new_n4307_), .B(core__abc_22172_new_n4321_), .Y(core__abc_22172_new_n4322_));
OR2X2 OR2X2_1774 ( .A(core__abc_22172_new_n4306_), .B(core__abc_22172_new_n4320_), .Y(core__abc_22172_new_n4323_));
OR2X2 OR2X2_1775 ( .A(core_v3_reg_17_), .B(core_mi_17_), .Y(core__abc_22172_new_n4329_));
OR2X2 OR2X2_1776 ( .A(core__abc_22172_new_n4326_), .B(core__abc_22172_new_n4331_), .Y(core__abc_22172_new_n4332_));
OR2X2 OR2X2_1777 ( .A(core__abc_22172_new_n3217_), .B(core__abc_22172_new_n4332_), .Y(core__abc_22172_new_n4333_));
OR2X2 OR2X2_1778 ( .A(core__abc_22172_new_n4325_), .B(core__abc_22172_new_n4333_), .Y(core__abc_22172_new_n4334_));
OR2X2 OR2X2_1779 ( .A(core__abc_22172_new_n3228_), .B(core_v3_reg_17_), .Y(core__abc_22172_new_n4335_));
OR2X2 OR2X2_178 ( .A(_abc_19873_new_n1291_), .B(_abc_19873_new_n1278_), .Y(_abc_19873_new_n1292_));
OR2X2 OR2X2_1780 ( .A(core__abc_22172_new_n4300_), .B(core__abc_22172_new_n4292_), .Y(core__abc_22172_new_n4338_));
OR2X2 OR2X2_1781 ( .A(core__abc_22172_new_n4343_), .B(core__abc_22172_new_n2131_), .Y(core__abc_22172_new_n4344_));
OR2X2 OR2X2_1782 ( .A(core__abc_22172_new_n4348_), .B(core__abc_22172_new_n3118_), .Y(core__abc_22172_new_n4349_));
OR2X2 OR2X2_1783 ( .A(core__abc_22172_new_n4349_), .B(core__abc_22172_new_n1585_), .Y(core__abc_22172_new_n4352_));
OR2X2 OR2X2_1784 ( .A(core__abc_22172_new_n4353_), .B(core__abc_22172_new_n1303_), .Y(core__abc_22172_new_n4354_));
OR2X2 OR2X2_1785 ( .A(core__abc_22172_new_n4355_), .B(core_v3_reg_2_), .Y(core__abc_22172_new_n4356_));
OR2X2 OR2X2_1786 ( .A(core__abc_22172_new_n4361_), .B(core__abc_22172_new_n4359_), .Y(core__abc_22172_new_n4362_));
OR2X2 OR2X2_1787 ( .A(core__abc_22172_new_n4364_), .B(core__abc_22172_new_n4365_), .Y(core__abc_22172_new_n4366_));
OR2X2 OR2X2_1788 ( .A(core__abc_22172_new_n4312_), .B(core__abc_22172_new_n2297_), .Y(core__abc_22172_new_n4367_));
OR2X2 OR2X2_1789 ( .A(core__abc_22172_new_n4367_), .B(core__abc_22172_new_n2319_), .Y(core__abc_22172_new_n4370_));
OR2X2 OR2X2_179 ( .A(_abc_19873_new_n1018_), .B(_abc_19873_new_n1037_), .Y(_abc_19873_new_n1295_));
OR2X2 OR2X2_1790 ( .A(core__abc_22172_new_n4373_), .B(core__abc_22172_new_n4375_), .Y(core__abc_22172_new_n4376_));
OR2X2 OR2X2_1791 ( .A(core__abc_22172_new_n4366_), .B(core__abc_22172_new_n4376_), .Y(core__abc_22172_new_n4377_));
OR2X2 OR2X2_1792 ( .A(core__abc_22172_new_n4378_), .B(core__abc_22172_new_n4381_), .Y(core__abc_22172_new_n4382_));
OR2X2 OR2X2_1793 ( .A(core_v3_reg_18_), .B(core_mi_18_), .Y(core__abc_22172_new_n4389_));
OR2X2 OR2X2_1794 ( .A(core__abc_22172_new_n4386_), .B(core__abc_22172_new_n4391_), .Y(core__abc_22172_new_n4392_));
OR2X2 OR2X2_1795 ( .A(core__abc_22172_new_n3217_), .B(core__abc_22172_new_n4392_), .Y(core__abc_22172_new_n4393_));
OR2X2 OR2X2_1796 ( .A(core__abc_22172_new_n4384_), .B(core__abc_22172_new_n4393_), .Y(core__abc_22172_new_n4394_));
OR2X2 OR2X2_1797 ( .A(core__abc_22172_new_n3228_), .B(core_v3_reg_18_), .Y(core__abc_22172_new_n4395_));
OR2X2 OR2X2_1798 ( .A(core__abc_22172_new_n4364_), .B(core__abc_22172_new_n4359_), .Y(core__abc_22172_new_n4398_));
OR2X2 OR2X2_1799 ( .A(core__abc_22172_new_n4399_), .B(core__abc_22172_new_n2148_), .Y(core__abc_22172_new_n4402_));
OR2X2 OR2X2_18 ( .A(_abc_19873_new_n951_), .B(_abc_19873_new_n952_), .Y(_abc_19873_new_n953_));
OR2X2 OR2X2_180 ( .A(_abc_19873_new_n1295_), .B(_abc_19873_new_n1294_), .Y(_abc_19873_new_n1296_));
OR2X2 OR2X2_1800 ( .A(core__abc_22172_new_n4404_), .B(core__abc_22172_new_n1605_), .Y(core__abc_22172_new_n4407_));
OR2X2 OR2X2_1801 ( .A(core__abc_22172_new_n4410_), .B(core__abc_22172_new_n4411_), .Y(core__abc_22172_new_n4412_));
OR2X2 OR2X2_1802 ( .A(core__abc_22172_new_n4403_), .B(core__abc_22172_new_n4412_), .Y(core__abc_22172_new_n4415_));
OR2X2 OR2X2_1803 ( .A(core__abc_22172_new_n4398_), .B(core__abc_22172_new_n4416_), .Y(core__abc_22172_new_n4419_));
OR2X2 OR2X2_1804 ( .A(core__abc_22172_new_n4367_), .B(core__abc_22172_new_n2314_), .Y(core__abc_22172_new_n4423_));
OR2X2 OR2X2_1805 ( .A(core__abc_22172_new_n4424_), .B(core__abc_22172_new_n2333_), .Y(core__abc_22172_new_n4425_));
OR2X2 OR2X2_1806 ( .A(core__abc_22172_new_n4430_), .B(core__abc_22172_new_n4431_), .Y(core__abc_22172_new_n4432_));
OR2X2 OR2X2_1807 ( .A(core__abc_22172_new_n4421_), .B(core__abc_22172_new_n4432_), .Y(core__abc_22172_new_n4433_));
OR2X2 OR2X2_1808 ( .A(core__abc_22172_new_n4420_), .B(core__abc_22172_new_n4434_), .Y(core__abc_22172_new_n4435_));
OR2X2 OR2X2_1809 ( .A(core_v3_reg_19_), .B(core_mi_19_), .Y(core__abc_22172_new_n4441_));
OR2X2 OR2X2_181 ( .A(_abc_19873_new_n1297_), .B(_abc_19873_new_n1298_), .Y(_abc_19873_new_n1299_));
OR2X2 OR2X2_1810 ( .A(core__abc_22172_new_n4438_), .B(core__abc_22172_new_n4443_), .Y(core__abc_22172_new_n4444_));
OR2X2 OR2X2_1811 ( .A(core__abc_22172_new_n3217_), .B(core__abc_22172_new_n4444_), .Y(core__abc_22172_new_n4445_));
OR2X2 OR2X2_1812 ( .A(core__abc_22172_new_n4437_), .B(core__abc_22172_new_n4445_), .Y(core__abc_22172_new_n4446_));
OR2X2 OR2X2_1813 ( .A(core__abc_22172_new_n3228_), .B(core_v3_reg_19_), .Y(core__abc_22172_new_n4447_));
OR2X2 OR2X2_1814 ( .A(core__abc_22172_new_n4413_), .B(core__abc_22172_new_n4359_), .Y(core__abc_22172_new_n4452_));
OR2X2 OR2X2_1815 ( .A(core__abc_22172_new_n4451_), .B(core__abc_22172_new_n4453_), .Y(core__abc_22172_new_n4454_));
OR2X2 OR2X2_1816 ( .A(core__abc_22172_new_n4456_), .B(core__abc_22172_new_n4454_), .Y(core__abc_22172_new_n4457_));
OR2X2 OR2X2_1817 ( .A(core__abc_22172_new_n4342_), .B(core__abc_22172_new_n4459_), .Y(core__abc_22172_new_n4460_));
OR2X2 OR2X2_1818 ( .A(core__abc_22172_new_n4461_), .B(core__abc_22172_new_n2140_), .Y(core__abc_22172_new_n4462_));
OR2X2 OR2X2_1819 ( .A(core__abc_22172_new_n4467_), .B(core__abc_22172_new_n4465_), .Y(core__abc_22172_new_n4468_));
OR2X2 OR2X2_182 ( .A(_abc_19873_new_n1296_), .B(_abc_19873_new_n1299_), .Y(_abc_19873_new_n1300_));
OR2X2 OR2X2_1820 ( .A(core__abc_22172_new_n4471_), .B(core__abc_22172_new_n4469_), .Y(core__abc_22172_new_n4472_));
OR2X2 OR2X2_1821 ( .A(core__abc_22172_new_n4474_), .B(core__abc_22172_new_n3122_), .Y(core__abc_22172_new_n4475_));
OR2X2 OR2X2_1822 ( .A(core__abc_22172_new_n4478_), .B(core__abc_22172_new_n4476_), .Y(core__abc_22172_new_n4479_));
OR2X2 OR2X2_1823 ( .A(core__abc_22172_new_n4480_), .B(core__abc_22172_new_n1338_), .Y(core__abc_22172_new_n4481_));
OR2X2 OR2X2_1824 ( .A(core__abc_22172_new_n4479_), .B(core_v3_reg_4_), .Y(core__abc_22172_new_n4482_));
OR2X2 OR2X2_1825 ( .A(core__abc_22172_new_n4485_), .B(core__abc_22172_new_n4486_), .Y(core__abc_22172_new_n4487_));
OR2X2 OR2X2_1826 ( .A(core__abc_22172_new_n4457_), .B(core__abc_22172_new_n4488_), .Y(core__abc_22172_new_n4491_));
OR2X2 OR2X2_1827 ( .A(core__abc_22172_new_n4426_), .B(core__abc_22172_new_n2331_), .Y(core__abc_22172_new_n4494_));
OR2X2 OR2X2_1828 ( .A(core__abc_22172_new_n4494_), .B(core__abc_22172_new_n2352_), .Y(core__abc_22172_new_n4495_));
OR2X2 OR2X2_1829 ( .A(core__abc_22172_new_n4498_), .B(core_v3_reg_47_), .Y(core__abc_22172_new_n4499_));
OR2X2 OR2X2_183 ( .A(_abc_19873_new_n1302_), .B(_abc_19873_new_n1303_), .Y(_abc_19873_new_n1304_));
OR2X2 OR2X2_1830 ( .A(core__abc_22172_new_n4501_), .B(core__abc_22172_new_n4500_), .Y(core__abc_22172_new_n4502_));
OR2X2 OR2X2_1831 ( .A(core__abc_22172_new_n4504_), .B(core__abc_22172_new_n4493_), .Y(core__abc_22172_new_n4505_));
OR2X2 OR2X2_1832 ( .A(core__abc_22172_new_n4503_), .B(core__abc_22172_new_n4492_), .Y(core__abc_22172_new_n4506_));
OR2X2 OR2X2_1833 ( .A(core_v3_reg_20_), .B(core_mi_20_), .Y(core__abc_22172_new_n4513_));
OR2X2 OR2X2_1834 ( .A(core__abc_22172_new_n4510_), .B(core__abc_22172_new_n4515_), .Y(core__abc_22172_new_n4516_));
OR2X2 OR2X2_1835 ( .A(core__abc_22172_new_n3217_), .B(core__abc_22172_new_n4516_), .Y(core__abc_22172_new_n4517_));
OR2X2 OR2X2_1836 ( .A(core__abc_22172_new_n4508_), .B(core__abc_22172_new_n4517_), .Y(core__abc_22172_new_n4518_));
OR2X2 OR2X2_1837 ( .A(core__abc_22172_new_n3228_), .B(core_v3_reg_20_), .Y(core__abc_22172_new_n4519_));
OR2X2 OR2X2_1838 ( .A(core__abc_22172_new_n4469_), .B(core__abc_22172_new_n2157_), .Y(core__abc_22172_new_n4522_));
OR2X2 OR2X2_1839 ( .A(core__abc_22172_new_n4524_), .B(core__abc_22172_new_n4525_), .Y(core__abc_22172_new_n4526_));
OR2X2 OR2X2_184 ( .A(_abc_19873_new_n1304_), .B(_abc_19873_new_n1301_), .Y(_abc_19873_new_n1305_));
OR2X2 OR2X2_1840 ( .A(core__abc_22172_new_n4476_), .B(core__abc_22172_new_n1616_), .Y(core__abc_22172_new_n4528_));
OR2X2 OR2X2_1841 ( .A(core__abc_22172_new_n4528_), .B(core__abc_22172_new_n1636_), .Y(core__abc_22172_new_n4529_));
OR2X2 OR2X2_1842 ( .A(core__abc_22172_new_n4534_), .B(core__abc_22172_new_n4535_), .Y(core__abc_22172_new_n4536_));
OR2X2 OR2X2_1843 ( .A(core__abc_22172_new_n4527_), .B(core__abc_22172_new_n4536_), .Y(core__abc_22172_new_n4537_));
OR2X2 OR2X2_1844 ( .A(core__abc_22172_new_n4526_), .B(core__abc_22172_new_n4538_), .Y(core__abc_22172_new_n4539_));
OR2X2 OR2X2_1845 ( .A(core__abc_22172_new_n4543_), .B(core__abc_22172_new_n4541_), .Y(core__abc_22172_new_n4545_));
OR2X2 OR2X2_1846 ( .A(core__abc_22172_new_n4546_), .B(core__abc_22172_new_n4544_), .Y(core__abc_22172_new_n4547_));
OR2X2 OR2X2_1847 ( .A(core__abc_22172_new_n4548_), .B(core__abc_22172_new_n3041_), .Y(core__abc_22172_new_n4549_));
OR2X2 OR2X2_1848 ( .A(core__abc_22172_new_n4547_), .B(core__abc_22172_new_n3038_), .Y(core__abc_22172_new_n4550_));
OR2X2 OR2X2_1849 ( .A(core_v3_reg_21_), .B(core_mi_21_), .Y(core__abc_22172_new_n4557_));
OR2X2 OR2X2_185 ( .A(_abc_19873_new_n1306_), .B(_abc_19873_new_n1307_), .Y(_abc_19873_new_n1308_));
OR2X2 OR2X2_1850 ( .A(core__abc_22172_new_n4554_), .B(core__abc_22172_new_n4559_), .Y(core__abc_22172_new_n4560_));
OR2X2 OR2X2_1851 ( .A(core__abc_22172_new_n3217_), .B(core__abc_22172_new_n4560_), .Y(core__abc_22172_new_n4561_));
OR2X2 OR2X2_1852 ( .A(core__abc_22172_new_n4552_), .B(core__abc_22172_new_n4561_), .Y(core__abc_22172_new_n4562_));
OR2X2 OR2X2_1853 ( .A(core__abc_22172_new_n3228_), .B(core_v3_reg_21_), .Y(core__abc_22172_new_n4563_));
OR2X2 OR2X2_1854 ( .A(core__abc_22172_new_n4569_), .B(core__abc_22172_new_n4485_), .Y(core__abc_22172_new_n4570_));
OR2X2 OR2X2_1855 ( .A(core__abc_22172_new_n4568_), .B(core__abc_22172_new_n4571_), .Y(core__abc_22172_new_n4572_));
OR2X2 OR2X2_1856 ( .A(core__abc_22172_new_n4576_), .B(core__abc_22172_new_n4575_), .Y(core__abc_22172_new_n4577_));
OR2X2 OR2X2_1857 ( .A(core__abc_22172_new_n4574_), .B(core__abc_22172_new_n4578_), .Y(core__abc_22172_new_n4579_));
OR2X2 OR2X2_1858 ( .A(core__abc_22172_new_n4582_), .B(core__abc_22172_new_n4580_), .Y(core__abc_22172_new_n4583_));
OR2X2 OR2X2_1859 ( .A(core__abc_22172_new_n4584_), .B(core__abc_22172_new_n3127_), .Y(core__abc_22172_new_n4585_));
OR2X2 OR2X2_186 ( .A(_abc_19873_new_n1309_), .B(_abc_19873_new_n1310_), .Y(_abc_19873_new_n1311_));
OR2X2 OR2X2_1860 ( .A(core__abc_22172_new_n4588_), .B(core__abc_22172_new_n4586_), .Y(core__abc_22172_new_n4589_));
OR2X2 OR2X2_1861 ( .A(core__abc_22172_new_n4590_), .B(core_v3_reg_6_), .Y(core__abc_22172_new_n4591_));
OR2X2 OR2X2_1862 ( .A(core__abc_22172_new_n4589_), .B(core__abc_22172_new_n1376_), .Y(core__abc_22172_new_n4592_));
OR2X2 OR2X2_1863 ( .A(core__abc_22172_new_n4583_), .B(core__abc_22172_new_n4594_), .Y(core__abc_22172_new_n4597_));
OR2X2 OR2X2_1864 ( .A(core__abc_22172_new_n4572_), .B(core__abc_22172_new_n4598_), .Y(core__abc_22172_new_n4601_));
OR2X2 OR2X2_1865 ( .A(core__abc_22172_new_n4602_), .B(core__abc_22172_new_n4566_), .Y(core__abc_22172_new_n4603_));
OR2X2 OR2X2_1866 ( .A(core__abc_22172_new_n4604_), .B(core__abc_22172_new_n3247_), .Y(core__abc_22172_new_n4605_));
OR2X2 OR2X2_1867 ( .A(core_v3_reg_22_), .B(core_mi_22_), .Y(core__abc_22172_new_n4612_));
OR2X2 OR2X2_1868 ( .A(core__abc_22172_new_n4609_), .B(core__abc_22172_new_n4614_), .Y(core__abc_22172_new_n4615_));
OR2X2 OR2X2_1869 ( .A(core__abc_22172_new_n3217_), .B(core__abc_22172_new_n4615_), .Y(core__abc_22172_new_n4616_));
OR2X2 OR2X2_187 ( .A(_abc_19873_new_n1308_), .B(_abc_19873_new_n1311_), .Y(_abc_19873_new_n1312_));
OR2X2 OR2X2_1870 ( .A(core__abc_22172_new_n4607_), .B(core__abc_22172_new_n4616_), .Y(core__abc_22172_new_n4617_));
OR2X2 OR2X2_1871 ( .A(core__abc_22172_new_n3228_), .B(core_v3_reg_22_), .Y(core__abc_22172_new_n4618_));
OR2X2 OR2X2_1872 ( .A(core__abc_22172_new_n4580_), .B(core__abc_22172_new_n2191_), .Y(core__abc_22172_new_n4622_));
OR2X2 OR2X2_1873 ( .A(core__abc_22172_new_n4622_), .B(core__abc_22172_new_n2210_), .Y(core__abc_22172_new_n4623_));
OR2X2 OR2X2_1874 ( .A(core__abc_22172_new_n4586_), .B(core__abc_22172_new_n1650_), .Y(core__abc_22172_new_n4627_));
OR2X2 OR2X2_1875 ( .A(core__abc_22172_new_n4629_), .B(core__abc_22172_new_n4630_), .Y(core__abc_22172_new_n4631_));
OR2X2 OR2X2_1876 ( .A(core__abc_22172_new_n4634_), .B(core__abc_22172_new_n4632_), .Y(core__abc_22172_new_n4635_));
OR2X2 OR2X2_1877 ( .A(core__abc_22172_new_n4626_), .B(core__abc_22172_new_n4635_), .Y(core__abc_22172_new_n4636_));
OR2X2 OR2X2_1878 ( .A(core__abc_22172_new_n4637_), .B(core__abc_22172_new_n4624_), .Y(core__abc_22172_new_n4638_));
OR2X2 OR2X2_1879 ( .A(core__abc_22172_new_n4638_), .B(core__abc_22172_new_n4639_), .Y(core__abc_22172_new_n4640_));
OR2X2 OR2X2_188 ( .A(_abc_19873_new_n1312_), .B(_abc_19873_new_n1305_), .Y(_abc_19873_new_n1313_));
OR2X2 OR2X2_1880 ( .A(core__abc_22172_new_n4621_), .B(core__abc_22172_new_n4642_), .Y(core__abc_22172_new_n4645_));
OR2X2 OR2X2_1881 ( .A(core__abc_22172_new_n4646_), .B(core__abc_22172_new_n3313_), .Y(core__abc_22172_new_n4647_));
OR2X2 OR2X2_1882 ( .A(core__abc_22172_new_n4648_), .B(core__abc_22172_new_n3311_), .Y(core__abc_22172_new_n4649_));
OR2X2 OR2X2_1883 ( .A(core_v3_reg_23_), .B(core_mi_23_), .Y(core__abc_22172_new_n4655_));
OR2X2 OR2X2_1884 ( .A(core__abc_22172_new_n4652_), .B(core__abc_22172_new_n4657_), .Y(core__abc_22172_new_n4658_));
OR2X2 OR2X2_1885 ( .A(core__abc_22172_new_n3217_), .B(core__abc_22172_new_n4658_), .Y(core__abc_22172_new_n4659_));
OR2X2 OR2X2_1886 ( .A(core__abc_22172_new_n4651_), .B(core__abc_22172_new_n4659_), .Y(core__abc_22172_new_n4660_));
OR2X2 OR2X2_1887 ( .A(core__abc_22172_new_n3228_), .B(core_v3_reg_23_), .Y(core__abc_22172_new_n4661_));
OR2X2 OR2X2_1888 ( .A(core__abc_22172_new_n4670_), .B(core__abc_22172_new_n4668_), .Y(core__abc_22172_new_n4671_));
OR2X2 OR2X2_1889 ( .A(core__abc_22172_new_n4667_), .B(core__abc_22172_new_n4671_), .Y(core__abc_22172_new_n4672_));
OR2X2 OR2X2_189 ( .A(_abc_19873_new_n1313_), .B(_abc_19873_new_n1300_), .Y(_abc_19873_new_n1314_));
OR2X2 OR2X2_1890 ( .A(core__abc_22172_new_n4672_), .B(core__abc_22172_new_n4666_), .Y(core__abc_22172_new_n4673_));
OR2X2 OR2X2_1891 ( .A(core__abc_22172_new_n4675_), .B(core__abc_22172_new_n4673_), .Y(core__abc_22172_new_n4676_));
OR2X2 OR2X2_1892 ( .A(core__abc_22172_new_n4683_), .B(core__abc_22172_new_n2208_), .Y(core__abc_22172_new_n4684_));
OR2X2 OR2X2_1893 ( .A(core__abc_22172_new_n4682_), .B(core__abc_22172_new_n4684_), .Y(core__abc_22172_new_n4685_));
OR2X2 OR2X2_1894 ( .A(core__abc_22172_new_n4681_), .B(core__abc_22172_new_n4685_), .Y(core__abc_22172_new_n4686_));
OR2X2 OR2X2_1895 ( .A(core__abc_22172_new_n4680_), .B(core__abc_22172_new_n4686_), .Y(core__abc_22172_new_n4687_));
OR2X2 OR2X2_1896 ( .A(core__abc_22172_new_n4218_), .B(core__abc_22172_new_n4689_), .Y(core__abc_22172_new_n4690_));
OR2X2 OR2X2_1897 ( .A(core__abc_22172_new_n4693_), .B(core__abc_22172_new_n4688_), .Y(core__abc_22172_new_n4694_));
OR2X2 OR2X2_1898 ( .A(core__abc_22172_new_n4695_), .B(core__abc_22172_new_n3132_), .Y(core__abc_22172_new_n4696_));
OR2X2 OR2X2_1899 ( .A(core__abc_22172_new_n4699_), .B(core__abc_22172_new_n4697_), .Y(core__abc_22172_new_n4700_));
OR2X2 OR2X2_19 ( .A(_abc_19873_new_n953_), .B(_abc_19873_new_n950_), .Y(_abc_19873_new_n954_));
OR2X2 OR2X2_190 ( .A(_abc_19873_new_n1317_), .B(_abc_19873_new_n1318_), .Y(_abc_19873_new_n1319_));
OR2X2 OR2X2_1900 ( .A(core__abc_22172_new_n4701_), .B(core_v3_reg_8_), .Y(core__abc_22172_new_n4702_));
OR2X2 OR2X2_1901 ( .A(core__abc_22172_new_n4700_), .B(core__abc_22172_new_n4703_), .Y(core__abc_22172_new_n4704_));
OR2X2 OR2X2_1902 ( .A(core__abc_22172_new_n4709_), .B(core__abc_22172_new_n4707_), .Y(core__abc_22172_new_n4710_));
OR2X2 OR2X2_1903 ( .A(core__abc_22172_new_n4714_), .B(core__abc_22172_new_n4712_), .Y(core__abc_22172_new_n4715_));
OR2X2 OR2X2_1904 ( .A(core__abc_22172_new_n4715_), .B(core__abc_22172_new_n3384_), .Y(core__abc_22172_new_n4716_));
OR2X2 OR2X2_1905 ( .A(core__abc_22172_new_n4717_), .B(core__abc_22172_new_n3380_), .Y(core__abc_22172_new_n4718_));
OR2X2 OR2X2_1906 ( .A(core_v3_reg_24_), .B(core_mi_24_), .Y(core__abc_22172_new_n4725_));
OR2X2 OR2X2_1907 ( .A(core__abc_22172_new_n4722_), .B(core__abc_22172_new_n4727_), .Y(core__abc_22172_new_n4728_));
OR2X2 OR2X2_1908 ( .A(core__abc_22172_new_n3217_), .B(core__abc_22172_new_n4728_), .Y(core__abc_22172_new_n4729_));
OR2X2 OR2X2_1909 ( .A(core__abc_22172_new_n4720_), .B(core__abc_22172_new_n4729_), .Y(core__abc_22172_new_n4730_));
OR2X2 OR2X2_191 ( .A(_abc_19873_new_n1319_), .B(_abc_19873_new_n1316_), .Y(_abc_19873_new_n1320_));
OR2X2 OR2X2_1910 ( .A(core__abc_22172_new_n3228_), .B(core_v3_reg_24_), .Y(core__abc_22172_new_n4731_));
OR2X2 OR2X2_1911 ( .A(core__abc_22172_new_n4688_), .B(core__abc_22172_new_n2225_), .Y(core__abc_22172_new_n4734_));
OR2X2 OR2X2_1912 ( .A(core__abc_22172_new_n4736_), .B(core__abc_22172_new_n4737_), .Y(core__abc_22172_new_n4738_));
OR2X2 OR2X2_1913 ( .A(core__abc_22172_new_n4697_), .B(core__abc_22172_new_n1684_), .Y(core__abc_22172_new_n4739_));
OR2X2 OR2X2_1914 ( .A(core__abc_22172_new_n4741_), .B(core__abc_22172_new_n4742_), .Y(core__abc_22172_new_n4743_));
OR2X2 OR2X2_1915 ( .A(core__abc_22172_new_n4743_), .B(core_v3_reg_9_), .Y(core__abc_22172_new_n4746_));
OR2X2 OR2X2_1916 ( .A(core__abc_22172_new_n4751_), .B(core__abc_22172_new_n4748_), .Y(core__abc_22172_new_n4752_));
OR2X2 OR2X2_1917 ( .A(core__abc_22172_new_n4755_), .B(core__abc_22172_new_n4752_), .Y(core__abc_22172_new_n4757_));
OR2X2 OR2X2_1918 ( .A(core__abc_22172_new_n4758_), .B(core__abc_22172_new_n4756_), .Y(core__abc_22172_new_n4759_));
OR2X2 OR2X2_1919 ( .A(core__abc_22172_new_n4760_), .B(core__abc_22172_new_n3433_), .Y(core__abc_22172_new_n4761_));
OR2X2 OR2X2_192 ( .A(_abc_19873_new_n1321_), .B(_abc_19873_new_n1322_), .Y(_abc_19873_new_n1323_));
OR2X2 OR2X2_1920 ( .A(core__abc_22172_new_n4759_), .B(core__abc_22172_new_n3430_), .Y(core__abc_22172_new_n4762_));
OR2X2 OR2X2_1921 ( .A(core_v3_reg_25_), .B(core_mi_25_), .Y(core__abc_22172_new_n4768_));
OR2X2 OR2X2_1922 ( .A(core__abc_22172_new_n4765_), .B(core__abc_22172_new_n4770_), .Y(core__abc_22172_new_n4771_));
OR2X2 OR2X2_1923 ( .A(core__abc_22172_new_n3217_), .B(core__abc_22172_new_n4771_), .Y(core__abc_22172_new_n4772_));
OR2X2 OR2X2_1924 ( .A(core__abc_22172_new_n4764_), .B(core__abc_22172_new_n4772_), .Y(core__abc_22172_new_n4773_));
OR2X2 OR2X2_1925 ( .A(core__abc_22172_new_n3228_), .B(core_v3_reg_25_), .Y(core__abc_22172_new_n4774_));
OR2X2 OR2X2_1926 ( .A(core__abc_22172_new_n4751_), .B(core__abc_22172_new_n4709_), .Y(core__abc_22172_new_n4781_));
OR2X2 OR2X2_1927 ( .A(core__abc_22172_new_n4779_), .B(core__abc_22172_new_n4782_), .Y(core__abc_22172_new_n4783_));
OR2X2 OR2X2_1928 ( .A(core__abc_22172_new_n4786_), .B(core__abc_22172_new_n2242_), .Y(core__abc_22172_new_n4787_));
OR2X2 OR2X2_1929 ( .A(core__abc_22172_new_n4785_), .B(core__abc_22172_new_n4787_), .Y(core__abc_22172_new_n4788_));
OR2X2 OR2X2_193 ( .A(_abc_19873_new_n1324_), .B(_abc_19873_new_n1325_), .Y(_abc_19873_new_n1326_));
OR2X2 OR2X2_1930 ( .A(core__abc_22172_new_n4791_), .B(core__abc_22172_new_n4789_), .Y(core__abc_22172_new_n4792_));
OR2X2 OR2X2_1931 ( .A(core__abc_22172_new_n4795_), .B(core__abc_22172_new_n3137_), .Y(core__abc_22172_new_n4796_));
OR2X2 OR2X2_1932 ( .A(core__abc_22172_new_n4798_), .B(core__abc_22172_new_n4799_), .Y(core__abc_22172_new_n4800_));
OR2X2 OR2X2_1933 ( .A(core__abc_22172_new_n4801_), .B(core__abc_22172_new_n4794_), .Y(core__abc_22172_new_n4802_));
OR2X2 OR2X2_1934 ( .A(core__abc_22172_new_n4800_), .B(core_v3_reg_10_), .Y(core__abc_22172_new_n4803_));
OR2X2 OR2X2_1935 ( .A(core__abc_22172_new_n4806_), .B(core__abc_22172_new_n4807_), .Y(core__abc_22172_new_n4808_));
OR2X2 OR2X2_1936 ( .A(core__abc_22172_new_n4783_), .B(core__abc_22172_new_n4809_), .Y(core__abc_22172_new_n4812_));
OR2X2 OR2X2_1937 ( .A(core__abc_22172_new_n4814_), .B(core__abc_22172_new_n3490_), .Y(core__abc_22172_new_n4815_));
OR2X2 OR2X2_1938 ( .A(core__abc_22172_new_n4813_), .B(core__abc_22172_new_n3491_), .Y(core__abc_22172_new_n4816_));
OR2X2 OR2X2_1939 ( .A(core_v3_reg_26_), .B(core_mi_26_), .Y(core__abc_22172_new_n4822_));
OR2X2 OR2X2_194 ( .A(_abc_19873_new_n1323_), .B(_abc_19873_new_n1326_), .Y(_abc_19873_new_n1327_));
OR2X2 OR2X2_1940 ( .A(core__abc_22172_new_n4819_), .B(core__abc_22172_new_n4824_), .Y(core__abc_22172_new_n4825_));
OR2X2 OR2X2_1941 ( .A(core__abc_22172_new_n3217_), .B(core__abc_22172_new_n4825_), .Y(core__abc_22172_new_n4826_));
OR2X2 OR2X2_1942 ( .A(core__abc_22172_new_n4818_), .B(core__abc_22172_new_n4826_), .Y(core__abc_22172_new_n4827_));
OR2X2 OR2X2_1943 ( .A(core__abc_22172_new_n3228_), .B(core_v3_reg_26_), .Y(core__abc_22172_new_n4828_));
OR2X2 OR2X2_1944 ( .A(core__abc_22172_new_n4789_), .B(core__abc_22172_new_n2259_), .Y(core__abc_22172_new_n4833_));
OR2X2 OR2X2_1945 ( .A(core__abc_22172_new_n4835_), .B(core__abc_22172_new_n4836_), .Y(core__abc_22172_new_n4837_));
OR2X2 OR2X2_1946 ( .A(core__abc_22172_new_n4799_), .B(core__abc_22172_new_n1718_), .Y(core__abc_22172_new_n4838_));
OR2X2 OR2X2_1947 ( .A(core__abc_22172_new_n4840_), .B(core__abc_22172_new_n4841_), .Y(core__abc_22172_new_n4842_));
OR2X2 OR2X2_1948 ( .A(core__abc_22172_new_n4842_), .B(core_v3_reg_11_), .Y(core__abc_22172_new_n4845_));
OR2X2 OR2X2_1949 ( .A(core__abc_22172_new_n4850_), .B(core__abc_22172_new_n4847_), .Y(core__abc_22172_new_n4851_));
OR2X2 OR2X2_195 ( .A(_abc_19873_new_n1328_), .B(_abc_19873_new_n1329_), .Y(_abc_19873_new_n1330_));
OR2X2 OR2X2_1950 ( .A(core__abc_22172_new_n4832_), .B(core__abc_22172_new_n4851_), .Y(core__abc_22172_new_n4854_));
OR2X2 OR2X2_1951 ( .A(core__abc_22172_new_n4855_), .B(core__abc_22172_new_n3563_), .Y(core__abc_22172_new_n4856_));
OR2X2 OR2X2_1952 ( .A(core__abc_22172_new_n4857_), .B(core__abc_22172_new_n3560_), .Y(core__abc_22172_new_n4858_));
OR2X2 OR2X2_1953 ( .A(core_v3_reg_27_), .B(core_mi_27_), .Y(core__abc_22172_new_n4865_));
OR2X2 OR2X2_1954 ( .A(core__abc_22172_new_n4862_), .B(core__abc_22172_new_n4867_), .Y(core__abc_22172_new_n4868_));
OR2X2 OR2X2_1955 ( .A(core__abc_22172_new_n3217_), .B(core__abc_22172_new_n4868_), .Y(core__abc_22172_new_n4869_));
OR2X2 OR2X2_1956 ( .A(core__abc_22172_new_n4860_), .B(core__abc_22172_new_n4869_), .Y(core__abc_22172_new_n4870_));
OR2X2 OR2X2_1957 ( .A(core__abc_22172_new_n3228_), .B(core_v3_reg_27_), .Y(core__abc_22172_new_n4871_));
OR2X2 OR2X2_1958 ( .A(core__abc_22172_new_n4837_), .B(core__abc_22172_new_n4846_), .Y(core__abc_22172_new_n4876_));
OR2X2 OR2X2_1959 ( .A(core__abc_22172_new_n4880_), .B(core__abc_22172_new_n4850_), .Y(core__abc_22172_new_n4881_));
OR2X2 OR2X2_196 ( .A(_abc_19873_new_n1331_), .B(_abc_19873_new_n1018_), .Y(_abc_19873_new_n1332_));
OR2X2 OR2X2_1960 ( .A(core__abc_22172_new_n4879_), .B(core__abc_22172_new_n4881_), .Y(core__abc_22172_new_n4882_));
OR2X2 OR2X2_1961 ( .A(core__abc_22172_new_n4884_), .B(core__abc_22172_new_n4882_), .Y(core__abc_22172_new_n4885_));
OR2X2 OR2X2_1962 ( .A(core__abc_22172_new_n4890_), .B(core__abc_22172_new_n2276_), .Y(core__abc_22172_new_n4891_));
OR2X2 OR2X2_1963 ( .A(core__abc_22172_new_n4889_), .B(core__abc_22172_new_n4891_), .Y(core__abc_22172_new_n4892_));
OR2X2 OR2X2_1964 ( .A(core__abc_22172_new_n4888_), .B(core__abc_22172_new_n4892_), .Y(core__abc_22172_new_n4893_));
OR2X2 OR2X2_1965 ( .A(core__abc_22172_new_n4692_), .B(core__abc_22172_new_n4895_), .Y(core__abc_22172_new_n4896_));
OR2X2 OR2X2_1966 ( .A(core__abc_22172_new_n4899_), .B(core__abc_22172_new_n4894_), .Y(core__abc_22172_new_n4900_));
OR2X2 OR2X2_1967 ( .A(core__abc_22172_new_n4903_), .B(core__abc_22172_new_n3141_), .Y(core__abc_22172_new_n4904_));
OR2X2 OR2X2_1968 ( .A(core__abc_22172_new_n4907_), .B(core__abc_22172_new_n4905_), .Y(core__abc_22172_new_n4908_));
OR2X2 OR2X2_1969 ( .A(core__abc_22172_new_n4909_), .B(core__abc_22172_new_n4902_), .Y(core__abc_22172_new_n4910_));
OR2X2 OR2X2_197 ( .A(_abc_19873_new_n1330_), .B(_abc_19873_new_n1332_), .Y(_abc_19873_new_n1333_));
OR2X2 OR2X2_1970 ( .A(core__abc_22172_new_n4908_), .B(core_v3_reg_12_), .Y(core__abc_22172_new_n4911_));
OR2X2 OR2X2_1971 ( .A(core__abc_22172_new_n4914_), .B(core__abc_22172_new_n4915_), .Y(core__abc_22172_new_n4916_));
OR2X2 OR2X2_1972 ( .A(core__abc_22172_new_n4885_), .B(core__abc_22172_new_n4917_), .Y(core__abc_22172_new_n4920_));
OR2X2 OR2X2_1973 ( .A(core__abc_22172_new_n4922_), .B(core__abc_22172_new_n3620_), .Y(core__abc_22172_new_n4923_));
OR2X2 OR2X2_1974 ( .A(core__abc_22172_new_n4921_), .B(core__abc_22172_new_n3621_), .Y(core__abc_22172_new_n4924_));
OR2X2 OR2X2_1975 ( .A(core_v3_reg_28_), .B(core_mi_28_), .Y(core__abc_22172_new_n4929_));
OR2X2 OR2X2_1976 ( .A(core__abc_22172_new_n4928_), .B(core__abc_22172_new_n4933_), .Y(core__abc_22172_new_n4934_));
OR2X2 OR2X2_1977 ( .A(core__abc_22172_new_n4926_), .B(core__abc_22172_new_n4934_), .Y(core__abc_22172_new_n4935_));
OR2X2 OR2X2_1978 ( .A(core__abc_22172_new_n4936_), .B(core__abc_22172_new_n4874_), .Y(core__abc_22172_new_n4937_));
OR2X2 OR2X2_1979 ( .A(core__abc_22172_new_n4894_), .B(core__abc_22172_new_n2293_), .Y(core__abc_22172_new_n4942_));
OR2X2 OR2X2_198 ( .A(_abc_19873_new_n1327_), .B(_abc_19873_new_n1333_), .Y(_abc_19873_new_n1334_));
OR2X2 OR2X2_1980 ( .A(core__abc_22172_new_n4944_), .B(core__abc_22172_new_n4945_), .Y(core__abc_22172_new_n4946_));
OR2X2 OR2X2_1981 ( .A(core__abc_22172_new_n4905_), .B(core__abc_22172_new_n1752_), .Y(core__abc_22172_new_n4947_));
OR2X2 OR2X2_1982 ( .A(core__abc_22172_new_n4949_), .B(core__abc_22172_new_n4950_), .Y(core__abc_22172_new_n4951_));
OR2X2 OR2X2_1983 ( .A(core__abc_22172_new_n4951_), .B(core_v3_reg_13_), .Y(core__abc_22172_new_n4954_));
OR2X2 OR2X2_1984 ( .A(core__abc_22172_new_n4964_), .B(core__abc_22172_new_n4965_), .Y(core__abc_22172_new_n4966_));
OR2X2 OR2X2_1985 ( .A(core__abc_22172_new_n4966_), .B(core__abc_22172_new_n3698_), .Y(core__abc_22172_new_n4967_));
OR2X2 OR2X2_1986 ( .A(core__abc_22172_new_n4968_), .B(core__abc_22172_new_n3697_), .Y(core__abc_22172_new_n4969_));
OR2X2 OR2X2_1987 ( .A(core_v3_reg_29_), .B(core_mi_29_), .Y(core__abc_22172_new_n4976_));
OR2X2 OR2X2_1988 ( .A(core__abc_22172_new_n4973_), .B(core__abc_22172_new_n4978_), .Y(core__abc_22172_new_n4979_));
OR2X2 OR2X2_1989 ( .A(core__abc_22172_new_n3217_), .B(core__abc_22172_new_n4979_), .Y(core__abc_22172_new_n4980_));
OR2X2 OR2X2_199 ( .A(_abc_19873_new_n1334_), .B(_abc_19873_new_n1320_), .Y(_abc_19873_new_n1335_));
OR2X2 OR2X2_1990 ( .A(core__abc_22172_new_n4971_), .B(core__abc_22172_new_n4980_), .Y(core__abc_22172_new_n4981_));
OR2X2 OR2X2_1991 ( .A(core__abc_22172_new_n3228_), .B(core_v3_reg_29_), .Y(core__abc_22172_new_n4982_));
OR2X2 OR2X2_1992 ( .A(core__abc_22172_new_n4987_), .B(core__abc_22172_new_n2310_), .Y(core__abc_22172_new_n4988_));
OR2X2 OR2X2_1993 ( .A(core__abc_22172_new_n4986_), .B(core__abc_22172_new_n4988_), .Y(core__abc_22172_new_n4989_));
OR2X2 OR2X2_1994 ( .A(core__abc_22172_new_n4898_), .B(core__abc_22172_new_n4991_), .Y(core__abc_22172_new_n4992_));
OR2X2 OR2X2_1995 ( .A(core__abc_22172_new_n4995_), .B(core__abc_22172_new_n4990_), .Y(core__abc_22172_new_n4996_));
OR2X2 OR2X2_1996 ( .A(core__abc_22172_new_n4998_), .B(core__abc_22172_new_n3148_), .Y(core__abc_22172_new_n4999_));
OR2X2 OR2X2_1997 ( .A(core__abc_22172_new_n5002_), .B(core__abc_22172_new_n5000_), .Y(core__abc_22172_new_n5003_));
OR2X2 OR2X2_1998 ( .A(core__abc_22172_new_n5004_), .B(core__abc_22172_new_n4997_), .Y(core__abc_22172_new_n5005_));
OR2X2 OR2X2_1999 ( .A(core__abc_22172_new_n5003_), .B(core_v3_reg_14_), .Y(core__abc_22172_new_n5006_));
OR2X2 OR2X2_2 ( .A(_abc_19873_new_n895_), .B(_abc_19873_new_n898_), .Y(_abc_19873_new_n899_));
OR2X2 OR2X2_20 ( .A(_abc_19873_new_n955_), .B(_abc_19873_new_n956_), .Y(_abc_19873_new_n957_));
OR2X2 OR2X2_200 ( .A(_abc_19873_new_n1337_), .B(_abc_19873_new_n1338_), .Y(_abc_19873_new_n1339_));
OR2X2 OR2X2_2000 ( .A(core__abc_22172_new_n5011_), .B(core__abc_22172_new_n5008_), .Y(core__abc_22172_new_n5012_));
OR2X2 OR2X2_2001 ( .A(core__abc_22172_new_n5015_), .B(core__abc_22172_new_n4956_), .Y(core__abc_22172_new_n5016_));
OR2X2 OR2X2_2002 ( .A(core__abc_22172_new_n5018_), .B(core__abc_22172_new_n5019_), .Y(core__abc_22172_new_n5020_));
OR2X2 OR2X2_2003 ( .A(core__abc_22172_new_n5020_), .B(core__abc_22172_new_n3752_), .Y(core__abc_22172_new_n5021_));
OR2X2 OR2X2_2004 ( .A(core__abc_22172_new_n5022_), .B(core__abc_22172_new_n3753_), .Y(core__abc_22172_new_n5023_));
OR2X2 OR2X2_2005 ( .A(core_v3_reg_30_), .B(core_mi_30_), .Y(core__abc_22172_new_n5030_));
OR2X2 OR2X2_2006 ( .A(core__abc_22172_new_n5027_), .B(core__abc_22172_new_n5032_), .Y(core__abc_22172_new_n5033_));
OR2X2 OR2X2_2007 ( .A(core__abc_22172_new_n3217_), .B(core__abc_22172_new_n5033_), .Y(core__abc_22172_new_n5034_));
OR2X2 OR2X2_2008 ( .A(core__abc_22172_new_n5025_), .B(core__abc_22172_new_n5034_), .Y(core__abc_22172_new_n5035_));
OR2X2 OR2X2_2009 ( .A(core__abc_22172_new_n3228_), .B(core_v3_reg_30_), .Y(core__abc_22172_new_n5036_));
OR2X2 OR2X2_201 ( .A(_abc_19873_new_n1192_), .B(_abc_19873_new_n1340_), .Y(_abc_19873_new_n1341_));
OR2X2 OR2X2_2010 ( .A(core__abc_22172_new_n5018_), .B(core__abc_22172_new_n5011_), .Y(core__abc_22172_new_n5039_));
OR2X2 OR2X2_2011 ( .A(core__abc_22172_new_n4990_), .B(core__abc_22172_new_n2327_), .Y(core__abc_22172_new_n5040_));
OR2X2 OR2X2_2012 ( .A(core__abc_22172_new_n5040_), .B(core__abc_22172_new_n2348_), .Y(core__abc_22172_new_n5041_));
OR2X2 OR2X2_2013 ( .A(core__abc_22172_new_n4994_), .B(core__abc_22172_new_n2335_), .Y(core__abc_22172_new_n5042_));
OR2X2 OR2X2_2014 ( .A(core__abc_22172_new_n5043_), .B(core__abc_22172_new_n2347_), .Y(core__abc_22172_new_n5044_));
OR2X2 OR2X2_2015 ( .A(core__abc_22172_new_n5000_), .B(core__abc_22172_new_n1786_), .Y(core__abc_22172_new_n5046_));
OR2X2 OR2X2_2016 ( .A(core__abc_22172_new_n5048_), .B(core__abc_22172_new_n5049_), .Y(core__abc_22172_new_n5050_));
OR2X2 OR2X2_2017 ( .A(core__abc_22172_new_n5054_), .B(core__abc_22172_new_n5051_), .Y(core__abc_22172_new_n5055_));
OR2X2 OR2X2_2018 ( .A(core__abc_22172_new_n5045_), .B(core__abc_22172_new_n5055_), .Y(core__abc_22172_new_n5056_));
OR2X2 OR2X2_2019 ( .A(core__abc_22172_new_n5057_), .B(core__abc_22172_new_n5058_), .Y(core__abc_22172_new_n5059_));
OR2X2 OR2X2_202 ( .A(_abc_19873_new_n1341_), .B(_abc_19873_new_n1339_), .Y(_abc_19873_new_n1342_));
OR2X2 OR2X2_2020 ( .A(core__abc_22172_new_n5050_), .B(core_v3_reg_15_), .Y(core__abc_22172_new_n5061_));
OR2X2 OR2X2_2021 ( .A(core__abc_22172_new_n5059_), .B(core__abc_22172_new_n5062_), .Y(core__abc_22172_new_n5063_));
OR2X2 OR2X2_2022 ( .A(core__abc_22172_new_n5039_), .B(core__abc_22172_new_n5064_), .Y(core__abc_22172_new_n5067_));
OR2X2 OR2X2_2023 ( .A(core__abc_22172_new_n5068_), .B(core__abc_22172_new_n3833_), .Y(core__abc_22172_new_n5069_));
OR2X2 OR2X2_2024 ( .A(core__abc_22172_new_n5070_), .B(core__abc_22172_new_n3830_), .Y(core__abc_22172_new_n5071_));
OR2X2 OR2X2_2025 ( .A(core_v3_reg_31_), .B(core_mi_31_), .Y(core__abc_22172_new_n5077_));
OR2X2 OR2X2_2026 ( .A(core__abc_22172_new_n5074_), .B(core__abc_22172_new_n5079_), .Y(core__abc_22172_new_n5080_));
OR2X2 OR2X2_2027 ( .A(core__abc_22172_new_n3217_), .B(core__abc_22172_new_n5080_), .Y(core__abc_22172_new_n5081_));
OR2X2 OR2X2_2028 ( .A(core__abc_22172_new_n5073_), .B(core__abc_22172_new_n5081_), .Y(core__abc_22172_new_n5082_));
OR2X2 OR2X2_2029 ( .A(core__abc_22172_new_n3228_), .B(core_v3_reg_31_), .Y(core__abc_22172_new_n5083_));
OR2X2 OR2X2_203 ( .A(_abc_19873_new_n1344_), .B(_abc_19873_new_n1345_), .Y(_abc_19873_new_n1346_));
OR2X2 OR2X2_2030 ( .A(core__abc_22172_new_n5098_), .B(core__abc_22172_new_n5011_), .Y(core__abc_22172_new_n5099_));
OR2X2 OR2X2_2031 ( .A(core__abc_22172_new_n5097_), .B(core__abc_22172_new_n5100_), .Y(core__abc_22172_new_n5101_));
OR2X2 OR2X2_2032 ( .A(core__abc_22172_new_n5101_), .B(core__abc_22172_new_n5094_), .Y(core__abc_22172_new_n5102_));
OR2X2 OR2X2_2033 ( .A(core__abc_22172_new_n5102_), .B(core__abc_22172_new_n5093_), .Y(core__abc_22172_new_n5103_));
OR2X2 OR2X2_2034 ( .A(core__abc_22172_new_n5103_), .B(core__abc_22172_new_n5092_), .Y(core__abc_22172_new_n5104_));
OR2X2 OR2X2_2035 ( .A(core__abc_22172_new_n5107_), .B(core__abc_22172_new_n5108_), .Y(core__abc_22172_new_n5109_));
OR2X2 OR2X2_2036 ( .A(core__abc_22172_new_n5110_), .B(core__abc_22172_new_n5105_), .Y(core__abc_22172_new_n5111_));
OR2X2 OR2X2_2037 ( .A(core__abc_22172_new_n5109_), .B(core_v3_reg_16_), .Y(core__abc_22172_new_n5112_));
OR2X2 OR2X2_2038 ( .A(core__abc_22172_new_n5115_), .B(core__abc_22172_new_n5116_), .Y(core__abc_22172_new_n5117_));
OR2X2 OR2X2_2039 ( .A(core__abc_22172_new_n4851_), .B(core__abc_22172_new_n4808_), .Y(core__abc_22172_new_n5123_));
OR2X2 OR2X2_204 ( .A(_abc_19873_new_n1346_), .B(_abc_19873_new_n1343_), .Y(_abc_19873_new_n1347_));
OR2X2 OR2X2_2040 ( .A(core__abc_22172_new_n5123_), .B(core__abc_22172_new_n5122_), .Y(core__abc_22172_new_n5124_));
OR2X2 OR2X2_2041 ( .A(core__abc_22172_new_n5128_), .B(core__abc_22172_new_n5098_), .Y(core__abc_22172_new_n5129_));
OR2X2 OR2X2_2042 ( .A(core__abc_22172_new_n5129_), .B(core__abc_22172_new_n5012_), .Y(core__abc_22172_new_n5130_));
OR2X2 OR2X2_2043 ( .A(core__abc_22172_new_n5130_), .B(core__abc_22172_new_n5127_), .Y(core__abc_22172_new_n5131_));
OR2X2 OR2X2_2044 ( .A(core__abc_22172_new_n5131_), .B(core__abc_22172_new_n5126_), .Y(core__abc_22172_new_n5132_));
OR2X2 OR2X2_2045 ( .A(core__abc_22172_new_n5014_), .B(core__abc_22172_new_n4956_), .Y(core__abc_22172_new_n5133_));
OR2X2 OR2X2_2046 ( .A(core__abc_22172_new_n5130_), .B(core__abc_22172_new_n5133_), .Y(core__abc_22172_new_n5134_));
OR2X2 OR2X2_2047 ( .A(core__abc_22172_new_n5140_), .B(core__abc_22172_new_n5119_), .Y(core__abc_22172_new_n5141_));
OR2X2 OR2X2_2048 ( .A(core__abc_22172_new_n5144_), .B(core__abc_22172_new_n5142_), .Y(core__abc_22172_new_n5145_));
OR2X2 OR2X2_2049 ( .A(core_v3_reg_32_), .B(core_mi_32_), .Y(core__abc_22172_new_n5148_));
OR2X2 OR2X2_205 ( .A(_abc_19873_new_n1348_), .B(_abc_19873_new_n1349_), .Y(_abc_19873_new_n1350_));
OR2X2 OR2X2_2050 ( .A(core__abc_22172_new_n5147_), .B(core__abc_22172_new_n5152_), .Y(core__abc_22172_new_n5153_));
OR2X2 OR2X2_2051 ( .A(core__abc_22172_new_n5146_), .B(core__abc_22172_new_n5153_), .Y(core__abc_22172_new_n5154_));
OR2X2 OR2X2_2052 ( .A(core__abc_22172_new_n5155_), .B(core__abc_22172_new_n5086_), .Y(core__abc_22172_new_n5156_));
OR2X2 OR2X2_2053 ( .A(core__abc_22172_new_n5119_), .B(core__abc_22172_new_n5115_), .Y(core__abc_22172_new_n5159_));
OR2X2 OR2X2_2054 ( .A(core__abc_22172_new_n5161_), .B(core__abc_22172_new_n2918_), .Y(core__abc_22172_new_n5162_));
OR2X2 OR2X2_2055 ( .A(core__abc_22172_new_n5108_), .B(core__abc_22172_new_n1820_), .Y(core__abc_22172_new_n5164_));
OR2X2 OR2X2_2056 ( .A(core__abc_22172_new_n5166_), .B(core__abc_22172_new_n5167_), .Y(core__abc_22172_new_n5168_));
OR2X2 OR2X2_2057 ( .A(core__abc_22172_new_n5168_), .B(core_v3_reg_17_), .Y(core__abc_22172_new_n5171_));
OR2X2 OR2X2_2058 ( .A(core__abc_22172_new_n5160_), .B(core__abc_22172_new_n5179_), .Y(core__abc_22172_new_n5180_));
OR2X2 OR2X2_2059 ( .A(core__abc_22172_new_n5159_), .B(core__abc_22172_new_n5178_), .Y(core__abc_22172_new_n5181_));
OR2X2 OR2X2_206 ( .A(_abc_19873_new_n1351_), .B(_abc_19873_new_n1352_), .Y(_abc_19873_new_n1353_));
OR2X2 OR2X2_2060 ( .A(core__abc_22172_new_n5184_), .B(core__abc_22172_new_n5185_), .Y(core__abc_22172_new_n5186_));
OR2X2 OR2X2_2061 ( .A(core_v3_reg_33_), .B(core_mi_33_), .Y(core__abc_22172_new_n5190_));
OR2X2 OR2X2_2062 ( .A(core__abc_22172_new_n5189_), .B(core__abc_22172_new_n5194_), .Y(core__abc_22172_new_n5195_));
OR2X2 OR2X2_2063 ( .A(core__abc_22172_new_n5187_), .B(core__abc_22172_new_n5195_), .Y(core__abc_22172_new_n5196_));
OR2X2 OR2X2_2064 ( .A(core__abc_22172_new_n5197_), .B(core__abc_22172_new_n5158_), .Y(core__abc_22172_new_n5198_));
OR2X2 OR2X2_2065 ( .A(core__abc_22172_new_n5174_), .B(core__abc_22172_new_n5115_), .Y(core__abc_22172_new_n5201_));
OR2X2 OR2X2_2066 ( .A(core__abc_22172_new_n5204_), .B(core__abc_22172_new_n5202_), .Y(core__abc_22172_new_n5205_));
OR2X2 OR2X2_2067 ( .A(core__abc_22172_new_n5207_), .B(core__abc_22172_new_n5206_), .Y(core__abc_22172_new_n5208_));
OR2X2 OR2X2_2068 ( .A(core__abc_22172_new_n5106_), .B(core__abc_22172_new_n5211_), .Y(core__abc_22172_new_n5212_));
OR2X2 OR2X2_2069 ( .A(core__abc_22172_new_n5215_), .B(core__abc_22172_new_n5216_), .Y(core__abc_22172_new_n5217_));
OR2X2 OR2X2_207 ( .A(_abc_19873_new_n1350_), .B(_abc_19873_new_n1353_), .Y(_abc_19873_new_n1354_));
OR2X2 OR2X2_2070 ( .A(core__abc_22172_new_n5218_), .B(core__abc_22172_new_n5210_), .Y(core__abc_22172_new_n5219_));
OR2X2 OR2X2_2071 ( .A(core__abc_22172_new_n5217_), .B(core_v3_reg_18_), .Y(core__abc_22172_new_n5220_));
OR2X2 OR2X2_2072 ( .A(core__abc_22172_new_n5223_), .B(core__abc_22172_new_n5224_), .Y(core__abc_22172_new_n5225_));
OR2X2 OR2X2_2073 ( .A(core__abc_22172_new_n5205_), .B(core__abc_22172_new_n5226_), .Y(core__abc_22172_new_n5229_));
OR2X2 OR2X2_2074 ( .A(core__abc_22172_new_n5231_), .B(core__abc_22172_new_n4012_), .Y(core__abc_22172_new_n5232_));
OR2X2 OR2X2_2075 ( .A(core__abc_22172_new_n5230_), .B(core__abc_22172_new_n4013_), .Y(core__abc_22172_new_n5233_));
OR2X2 OR2X2_2076 ( .A(core_v3_reg_34_), .B(core_mi_34_), .Y(core__abc_22172_new_n5237_));
OR2X2 OR2X2_2077 ( .A(core__abc_22172_new_n5236_), .B(core__abc_22172_new_n5241_), .Y(core__abc_22172_new_n5242_));
OR2X2 OR2X2_2078 ( .A(core__abc_22172_new_n5235_), .B(core__abc_22172_new_n5242_), .Y(core__abc_22172_new_n5243_));
OR2X2 OR2X2_2079 ( .A(core__abc_22172_new_n5244_), .B(core__abc_22172_new_n5200_), .Y(core__abc_22172_new_n5245_));
OR2X2 OR2X2_208 ( .A(_abc_19873_new_n1354_), .B(_abc_19873_new_n1347_), .Y(_abc_19873_new_n1355_));
OR2X2 OR2X2_2080 ( .A(core__abc_22172_new_n5206_), .B(core__abc_22172_new_n1296_), .Y(core__abc_22172_new_n5250_));
OR2X2 OR2X2_2081 ( .A(core__abc_22172_new_n5252_), .B(core__abc_22172_new_n5253_), .Y(core__abc_22172_new_n5254_));
OR2X2 OR2X2_2082 ( .A(core__abc_22172_new_n5215_), .B(core__abc_22172_new_n1855_), .Y(core__abc_22172_new_n5255_));
OR2X2 OR2X2_2083 ( .A(core__abc_22172_new_n5255_), .B(core__abc_22172_new_n1874_), .Y(core__abc_22172_new_n5256_));
OR2X2 OR2X2_2084 ( .A(core__abc_22172_new_n5260_), .B(core_v3_reg_19_), .Y(core__abc_22172_new_n5263_));
OR2X2 OR2X2_2085 ( .A(core__abc_22172_new_n5264_), .B(core__abc_22172_new_n5254_), .Y(core__abc_22172_new_n5265_));
OR2X2 OR2X2_2086 ( .A(core__abc_22172_new_n5266_), .B(core__abc_22172_new_n5267_), .Y(core__abc_22172_new_n5268_));
OR2X2 OR2X2_2087 ( .A(core__abc_22172_new_n5249_), .B(core__abc_22172_new_n5268_), .Y(core__abc_22172_new_n5269_));
OR2X2 OR2X2_2088 ( .A(core__abc_22172_new_n5270_), .B(core__abc_22172_new_n5272_), .Y(core__abc_22172_new_n5273_));
OR2X2 OR2X2_2089 ( .A(core__abc_22172_new_n5274_), .B(core__abc_22172_new_n5247_), .Y(core__abc_22172_new_n5275_));
OR2X2 OR2X2_209 ( .A(_abc_19873_new_n1355_), .B(_abc_19873_new_n1342_), .Y(_abc_19873_new_n1356_));
OR2X2 OR2X2_2090 ( .A(core__abc_22172_new_n5276_), .B(core__abc_22172_new_n4089_), .Y(core__abc_22172_new_n5277_));
OR2X2 OR2X2_2091 ( .A(core_v3_reg_35_), .B(core_mi_35_), .Y(core__abc_22172_new_n5283_));
OR2X2 OR2X2_2092 ( .A(core__abc_22172_new_n5280_), .B(core__abc_22172_new_n5285_), .Y(core__abc_22172_new_n5286_));
OR2X2 OR2X2_2093 ( .A(core__abc_22172_new_n3217_), .B(core__abc_22172_new_n5286_), .Y(core__abc_22172_new_n5287_));
OR2X2 OR2X2_2094 ( .A(core__abc_22172_new_n5279_), .B(core__abc_22172_new_n5287_), .Y(core__abc_22172_new_n5288_));
OR2X2 OR2X2_2095 ( .A(core__abc_22172_new_n3228_), .B(core_v3_reg_35_), .Y(core__abc_22172_new_n5289_));
OR2X2 OR2X2_2096 ( .A(core__abc_22172_new_n5267_), .B(core__abc_22172_new_n5248_), .Y(core__abc_22172_new_n5295_));
OR2X2 OR2X2_2097 ( .A(core__abc_22172_new_n5294_), .B(core__abc_22172_new_n5297_), .Y(core__abc_22172_new_n5298_));
OR2X2 OR2X2_2098 ( .A(core__abc_22172_new_n5300_), .B(core__abc_22172_new_n5298_), .Y(core__abc_22172_new_n5301_));
OR2X2 OR2X2_2099 ( .A(core__abc_22172_new_n5303_), .B(core__abc_22172_new_n5302_), .Y(core__abc_22172_new_n5304_));
OR2X2 OR2X2_21 ( .A(_abc_19873_new_n958_), .B(_abc_19873_new_n959_), .Y(_abc_19873_new_n960_));
OR2X2 OR2X2_210 ( .A(_abc_19873_new_n1359_), .B(_abc_19873_new_n1360_), .Y(_abc_19873_new_n1361_));
OR2X2 OR2X2_2100 ( .A(core__abc_22172_new_n5307_), .B(core__abc_22172_new_n3169_), .Y(core__abc_22172_new_n5308_));
OR2X2 OR2X2_2101 ( .A(core__abc_22172_new_n5311_), .B(core__abc_22172_new_n5309_), .Y(core__abc_22172_new_n5312_));
OR2X2 OR2X2_2102 ( .A(core__abc_22172_new_n5313_), .B(core__abc_22172_new_n5306_), .Y(core__abc_22172_new_n5314_));
OR2X2 OR2X2_2103 ( .A(core__abc_22172_new_n5312_), .B(core_v3_reg_20_), .Y(core__abc_22172_new_n5315_));
OR2X2 OR2X2_2104 ( .A(core__abc_22172_new_n5318_), .B(core__abc_22172_new_n5319_), .Y(core__abc_22172_new_n5320_));
OR2X2 OR2X2_2105 ( .A(core__abc_22172_new_n5301_), .B(core__abc_22172_new_n5321_), .Y(core__abc_22172_new_n5324_));
OR2X2 OR2X2_2106 ( .A(core__abc_22172_new_n5325_), .B(core__abc_22172_new_n4144_), .Y(core__abc_22172_new_n5326_));
OR2X2 OR2X2_2107 ( .A(core__abc_22172_new_n5327_), .B(core__abc_22172_new_n4143_), .Y(core__abc_22172_new_n5328_));
OR2X2 OR2X2_2108 ( .A(core_v3_reg_36_), .B(core_mi_36_), .Y(core__abc_22172_new_n5332_));
OR2X2 OR2X2_2109 ( .A(core__abc_22172_new_n5331_), .B(core__abc_22172_new_n5336_), .Y(core__abc_22172_new_n5337_));
OR2X2 OR2X2_211 ( .A(_abc_19873_new_n1361_), .B(_abc_19873_new_n1358_), .Y(_abc_19873_new_n1362_));
OR2X2 OR2X2_2110 ( .A(core__abc_22172_new_n5330_), .B(core__abc_22172_new_n5337_), .Y(core__abc_22172_new_n5338_));
OR2X2 OR2X2_2111 ( .A(core__abc_22172_new_n5339_), .B(core__abc_22172_new_n5292_), .Y(core__abc_22172_new_n5340_));
OR2X2 OR2X2_2112 ( .A(core__abc_22172_new_n5302_), .B(core__abc_22172_new_n1333_), .Y(core__abc_22172_new_n5344_));
OR2X2 OR2X2_2113 ( .A(core__abc_22172_new_n5346_), .B(core__abc_22172_new_n5347_), .Y(core__abc_22172_new_n5348_));
OR2X2 OR2X2_2114 ( .A(core__abc_22172_new_n5309_), .B(core__abc_22172_new_n1889_), .Y(core__abc_22172_new_n5349_));
OR2X2 OR2X2_2115 ( .A(core__abc_22172_new_n5351_), .B(core__abc_22172_new_n5352_), .Y(core__abc_22172_new_n5353_));
OR2X2 OR2X2_2116 ( .A(core__abc_22172_new_n5353_), .B(core_v3_reg_21_), .Y(core__abc_22172_new_n5356_));
OR2X2 OR2X2_2117 ( .A(core__abc_22172_new_n5357_), .B(core__abc_22172_new_n5348_), .Y(core__abc_22172_new_n5359_));
OR2X2 OR2X2_2118 ( .A(core__abc_22172_new_n5360_), .B(core__abc_22172_new_n5358_), .Y(core__abc_22172_new_n5361_));
OR2X2 OR2X2_2119 ( .A(core__abc_22172_new_n5375_), .B(core__abc_22172_new_n5373_), .Y(core__abc_22172_new_n5376_));
OR2X2 OR2X2_212 ( .A(_abc_19873_new_n1363_), .B(_abc_19873_new_n1364_), .Y(_abc_19873_new_n1365_));
OR2X2 OR2X2_2120 ( .A(core_v3_reg_37_), .B(core_mi_37_), .Y(core__abc_22172_new_n5380_));
OR2X2 OR2X2_2121 ( .A(core__abc_22172_new_n5379_), .B(core__abc_22172_new_n5384_), .Y(core__abc_22172_new_n5385_));
OR2X2 OR2X2_2122 ( .A(core__abc_22172_new_n5377_), .B(core__abc_22172_new_n5385_), .Y(core__abc_22172_new_n5386_));
OR2X2 OR2X2_2123 ( .A(core__abc_22172_new_n5387_), .B(core__abc_22172_new_n5342_), .Y(core__abc_22172_new_n5388_));
OR2X2 OR2X2_2124 ( .A(core__abc_22172_new_n5366_), .B(core__abc_22172_new_n5360_), .Y(core__abc_22172_new_n5391_));
OR2X2 OR2X2_2125 ( .A(core__abc_22172_new_n5395_), .B(core__abc_22172_new_n2930_), .Y(core__abc_22172_new_n5396_));
OR2X2 OR2X2_2126 ( .A(core__abc_22172_new_n5396_), .B(core__abc_22172_new_n1373_), .Y(core__abc_22172_new_n5399_));
OR2X2 OR2X2_2127 ( .A(core__abc_22172_new_n5402_), .B(core__abc_22172_new_n3176_), .Y(core__abc_22172_new_n5403_));
OR2X2 OR2X2_2128 ( .A(core__abc_22172_new_n5405_), .B(core__abc_22172_new_n5406_), .Y(core__abc_22172_new_n5407_));
OR2X2 OR2X2_2129 ( .A(core__abc_22172_new_n5408_), .B(core_v3_reg_22_), .Y(core__abc_22172_new_n5409_));
OR2X2 OR2X2_213 ( .A(_abc_19873_new_n1366_), .B(_abc_19873_new_n1367_), .Y(_abc_19873_new_n1368_));
OR2X2 OR2X2_2130 ( .A(core__abc_22172_new_n5407_), .B(core__abc_22172_new_n5410_), .Y(core__abc_22172_new_n5411_));
OR2X2 OR2X2_2131 ( .A(core__abc_22172_new_n5414_), .B(core__abc_22172_new_n5415_), .Y(core__abc_22172_new_n5416_));
OR2X2 OR2X2_2132 ( .A(core__abc_22172_new_n5418_), .B(core__abc_22172_new_n5419_), .Y(core__abc_22172_new_n5420_));
OR2X2 OR2X2_2133 ( .A(core__abc_22172_new_n5424_), .B(core__abc_22172_new_n5421_), .Y(core__abc_22172_new_n5425_));
OR2X2 OR2X2_2134 ( .A(core_v3_reg_38_), .B(core_mi_38_), .Y(core__abc_22172_new_n5429_));
OR2X2 OR2X2_2135 ( .A(core__abc_22172_new_n5428_), .B(core__abc_22172_new_n5433_), .Y(core__abc_22172_new_n5434_));
OR2X2 OR2X2_2136 ( .A(core__abc_22172_new_n5426_), .B(core__abc_22172_new_n5434_), .Y(core__abc_22172_new_n5435_));
OR2X2 OR2X2_2137 ( .A(core__abc_22172_new_n5436_), .B(core__abc_22172_new_n5390_), .Y(core__abc_22172_new_n5437_));
OR2X2 OR2X2_2138 ( .A(core__abc_22172_new_n5418_), .B(core__abc_22172_new_n5415_), .Y(core__abc_22172_new_n5439_));
OR2X2 OR2X2_2139 ( .A(core__abc_22172_new_n5440_), .B(core__abc_22172_new_n1400_), .Y(core__abc_22172_new_n5443_));
OR2X2 OR2X2_214 ( .A(_abc_19873_new_n1365_), .B(_abc_19873_new_n1368_), .Y(_abc_19873_new_n1369_));
OR2X2 OR2X2_2140 ( .A(core__abc_22172_new_n5406_), .B(core__abc_22172_new_n1923_), .Y(core__abc_22172_new_n5445_));
OR2X2 OR2X2_2141 ( .A(core__abc_22172_new_n5447_), .B(core__abc_22172_new_n5448_), .Y(core__abc_22172_new_n5449_));
OR2X2 OR2X2_2142 ( .A(core__abc_22172_new_n5449_), .B(core_v3_reg_23_), .Y(core__abc_22172_new_n5452_));
OR2X2 OR2X2_2143 ( .A(core__abc_22172_new_n5454_), .B(core__abc_22172_new_n5444_), .Y(core__abc_22172_new_n5457_));
OR2X2 OR2X2_2144 ( .A(core__abc_22172_new_n5439_), .B(core__abc_22172_new_n5458_), .Y(core__abc_22172_new_n5459_));
OR2X2 OR2X2_2145 ( .A(core__abc_22172_new_n5461_), .B(core__abc_22172_new_n5455_), .Y(core__abc_22172_new_n5462_));
OR2X2 OR2X2_2146 ( .A(core__abc_22172_new_n5460_), .B(core__abc_22172_new_n5462_), .Y(core__abc_22172_new_n5463_));
OR2X2 OR2X2_2147 ( .A(core__abc_22172_new_n5465_), .B(core__abc_22172_new_n4357_), .Y(core__abc_22172_new_n5466_));
OR2X2 OR2X2_2148 ( .A(core__abc_22172_new_n5464_), .B(core__abc_22172_new_n4358_), .Y(core__abc_22172_new_n5467_));
OR2X2 OR2X2_2149 ( .A(core_v3_reg_39_), .B(core_mi_39_), .Y(core__abc_22172_new_n5473_));
OR2X2 OR2X2_215 ( .A(_abc_19873_new_n1370_), .B(_abc_19873_new_n1371_), .Y(_abc_19873_new_n1372_));
OR2X2 OR2X2_2150 ( .A(core__abc_22172_new_n5470_), .B(core__abc_22172_new_n5475_), .Y(core__abc_22172_new_n5476_));
OR2X2 OR2X2_2151 ( .A(core__abc_22172_new_n3217_), .B(core__abc_22172_new_n5476_), .Y(core__abc_22172_new_n5477_));
OR2X2 OR2X2_2152 ( .A(core__abc_22172_new_n5469_), .B(core__abc_22172_new_n5477_), .Y(core__abc_22172_new_n5478_));
OR2X2 OR2X2_2153 ( .A(core__abc_22172_new_n3228_), .B(core_v3_reg_39_), .Y(core__abc_22172_new_n5479_));
OR2X2 OR2X2_2154 ( .A(core__abc_22172_new_n5455_), .B(core__abc_22172_new_n5415_), .Y(core__abc_22172_new_n5487_));
OR2X2 OR2X2_2155 ( .A(core__abc_22172_new_n5486_), .B(core__abc_22172_new_n5488_), .Y(core__abc_22172_new_n5489_));
OR2X2 OR2X2_2156 ( .A(core__abc_22172_new_n5489_), .B(core__abc_22172_new_n5485_), .Y(core__abc_22172_new_n5490_));
OR2X2 OR2X2_2157 ( .A(core__abc_22172_new_n5492_), .B(core__abc_22172_new_n5490_), .Y(core__abc_22172_new_n5493_));
OR2X2 OR2X2_2158 ( .A(core__abc_22172_new_n5495_), .B(core__abc_22172_new_n5494_), .Y(core__abc_22172_new_n5496_));
OR2X2 OR2X2_2159 ( .A(core__abc_22172_new_n5501_), .B(core__abc_22172_new_n5499_), .Y(core__abc_22172_new_n5502_));
OR2X2 OR2X2_216 ( .A(_abc_19873_new_n1373_), .B(_abc_19873_new_n1037_), .Y(_abc_19873_new_n1374_));
OR2X2 OR2X2_2160 ( .A(core__abc_22172_new_n5503_), .B(core__abc_22172_new_n5498_), .Y(core__abc_22172_new_n5504_));
OR2X2 OR2X2_2161 ( .A(core__abc_22172_new_n5502_), .B(core_v3_reg_24_), .Y(core__abc_22172_new_n5505_));
OR2X2 OR2X2_2162 ( .A(core__abc_22172_new_n5508_), .B(core__abc_22172_new_n5509_), .Y(core__abc_22172_new_n5510_));
OR2X2 OR2X2_2163 ( .A(core__abc_22172_new_n5139_), .B(core__abc_22172_new_n5514_), .Y(core__abc_22172_new_n5515_));
OR2X2 OR2X2_2164 ( .A(core__abc_22172_new_n5517_), .B(core__abc_22172_new_n5512_), .Y(core__abc_22172_new_n5518_));
OR2X2 OR2X2_2165 ( .A(core__abc_22172_new_n5522_), .B(core__abc_22172_new_n5519_), .Y(core__abc_22172_new_n5523_));
OR2X2 OR2X2_2166 ( .A(core_v3_reg_40_), .B(core_mi_40_), .Y(core__abc_22172_new_n5526_));
OR2X2 OR2X2_2167 ( .A(core__abc_22172_new_n5525_), .B(core__abc_22172_new_n5530_), .Y(core__abc_22172_new_n5531_));
OR2X2 OR2X2_2168 ( .A(core__abc_22172_new_n5524_), .B(core__abc_22172_new_n5531_), .Y(core__abc_22172_new_n5532_));
OR2X2 OR2X2_2169 ( .A(core__abc_22172_new_n5533_), .B(core__abc_22172_new_n5482_), .Y(core__abc_22172_new_n5534_));
OR2X2 OR2X2_217 ( .A(_abc_19873_new_n1372_), .B(_abc_19873_new_n1374_), .Y(_abc_19873_new_n1375_));
OR2X2 OR2X2_2170 ( .A(core__abc_22172_new_n5494_), .B(core__abc_22172_new_n1409_), .Y(core__abc_22172_new_n5541_));
OR2X2 OR2X2_2171 ( .A(core__abc_22172_new_n5543_), .B(core__abc_22172_new_n5544_), .Y(core__abc_22172_new_n5545_));
OR2X2 OR2X2_2172 ( .A(core__abc_22172_new_n5499_), .B(core__abc_22172_new_n1956_), .Y(core__abc_22172_new_n5548_));
OR2X2 OR2X2_2173 ( .A(core__abc_22172_new_n5550_), .B(core__abc_22172_new_n5551_), .Y(core__abc_22172_new_n5552_));
OR2X2 OR2X2_2174 ( .A(core__abc_22172_new_n5555_), .B(core__abc_22172_new_n5553_), .Y(core__abc_22172_new_n5556_));
OR2X2 OR2X2_2175 ( .A(core__abc_22172_new_n5540_), .B(core__abc_22172_new_n5562_), .Y(core__abc_22172_new_n5563_));
OR2X2 OR2X2_2176 ( .A(core__abc_22172_new_n5539_), .B(core__abc_22172_new_n5564_), .Y(core__abc_22172_new_n5565_));
OR2X2 OR2X2_2177 ( .A(core__abc_22172_new_n5567_), .B(core__abc_22172_new_n4483_), .Y(core__abc_22172_new_n5568_));
OR2X2 OR2X2_2178 ( .A(core__abc_22172_new_n5566_), .B(core__abc_22172_new_n4484_), .Y(core__abc_22172_new_n5569_));
OR2X2 OR2X2_2179 ( .A(core_v3_reg_41_), .B(core_mi_41_), .Y(core__abc_22172_new_n5573_));
OR2X2 OR2X2_218 ( .A(_abc_19873_new_n1369_), .B(_abc_19873_new_n1375_), .Y(_abc_19873_new_n1376_));
OR2X2 OR2X2_2180 ( .A(core__abc_22172_new_n5572_), .B(core__abc_22172_new_n5577_), .Y(core__abc_22172_new_n5578_));
OR2X2 OR2X2_2181 ( .A(core__abc_22172_new_n5571_), .B(core__abc_22172_new_n5578_), .Y(core__abc_22172_new_n5579_));
OR2X2 OR2X2_2182 ( .A(core__abc_22172_new_n5580_), .B(core__abc_22172_new_n5536_), .Y(core__abc_22172_new_n5581_));
OR2X2 OR2X2_2183 ( .A(core__abc_22172_new_n5584_), .B(core__abc_22172_new_n2945_), .Y(core__abc_22172_new_n5585_));
OR2X2 OR2X2_2184 ( .A(core__abc_22172_new_n5588_), .B(core__abc_22172_new_n5586_), .Y(core__abc_22172_new_n5589_));
OR2X2 OR2X2_2185 ( .A(core__abc_22172_new_n5593_), .B(core__abc_22172_new_n3184_), .Y(core__abc_22172_new_n5594_));
OR2X2 OR2X2_2186 ( .A(core__abc_22172_new_n5595_), .B(core__abc_22172_new_n5591_), .Y(core__abc_22172_new_n5596_));
OR2X2 OR2X2_2187 ( .A(core__abc_22172_new_n5594_), .B(core_v3_reg_26_), .Y(core__abc_22172_new_n5597_));
OR2X2 OR2X2_2188 ( .A(core__abc_22172_new_n5600_), .B(core__abc_22172_new_n5601_), .Y(core__abc_22172_new_n5602_));
OR2X2 OR2X2_2189 ( .A(core__abc_22172_new_n5558_), .B(core__abc_22172_new_n5508_), .Y(core__abc_22172_new_n5603_));
OR2X2 OR2X2_219 ( .A(_abc_19873_new_n1376_), .B(_abc_19873_new_n1362_), .Y(_abc_19873_new_n1377_));
OR2X2 OR2X2_2190 ( .A(core__abc_22172_new_n5605_), .B(core__abc_22172_new_n5560_), .Y(core__abc_22172_new_n5606_));
OR2X2 OR2X2_2191 ( .A(core__abc_22172_new_n5606_), .B(core__abc_22172_new_n5602_), .Y(core__abc_22172_new_n5607_));
OR2X2 OR2X2_2192 ( .A(core__abc_22172_new_n5610_), .B(core__abc_22172_new_n4536_), .Y(core__abc_22172_new_n5611_));
OR2X2 OR2X2_2193 ( .A(core__abc_22172_new_n5612_), .B(core__abc_22172_new_n4538_), .Y(core__abc_22172_new_n5613_));
OR2X2 OR2X2_2194 ( .A(core_v3_reg_42_), .B(core_mi_42_), .Y(core__abc_22172_new_n5618_));
OR2X2 OR2X2_2195 ( .A(core__abc_22172_new_n5617_), .B(core__abc_22172_new_n5622_), .Y(core__abc_22172_new_n5623_));
OR2X2 OR2X2_2196 ( .A(core__abc_22172_new_n5615_), .B(core__abc_22172_new_n5623_), .Y(core__abc_22172_new_n5624_));
OR2X2 OR2X2_2197 ( .A(core__abc_22172_new_n5625_), .B(core__abc_22172_new_n5583_), .Y(core__abc_22172_new_n5626_));
OR2X2 OR2X2_2198 ( .A(core__abc_22172_new_n5586_), .B(core__abc_22172_new_n1443_), .Y(core__abc_22172_new_n5630_));
OR2X2 OR2X2_2199 ( .A(core__abc_22172_new_n5630_), .B(core__abc_22172_new_n1462_), .Y(core__abc_22172_new_n5631_));
OR2X2 OR2X2_22 ( .A(_abc_19873_new_n957_), .B(_abc_19873_new_n960_), .Y(_abc_19873_new_n961_));
OR2X2 OR2X2_220 ( .A(_abc_19873_new_n1380_), .B(_abc_19873_new_n1381_), .Y(_abc_19873_new_n1382_));
OR2X2 OR2X2_2200 ( .A(core__abc_22172_new_n5635_), .B(core__abc_22172_new_n5637_), .Y(core__abc_22172_new_n5638_));
OR2X2 OR2X2_2201 ( .A(core__abc_22172_new_n5629_), .B(core__abc_22172_new_n5638_), .Y(core__abc_22172_new_n5639_));
OR2X2 OR2X2_2202 ( .A(core__abc_22172_new_n5640_), .B(core__abc_22172_new_n5641_), .Y(core__abc_22172_new_n5642_));
OR2X2 OR2X2_2203 ( .A(core__abc_22172_new_n5644_), .B(core__abc_22172_new_n4594_), .Y(core__abc_22172_new_n5645_));
OR2X2 OR2X2_2204 ( .A(core__abc_22172_new_n5643_), .B(core__abc_22172_new_n4593_), .Y(core__abc_22172_new_n5646_));
OR2X2 OR2X2_2205 ( .A(core_v3_reg_43_), .B(core_mi_43_), .Y(core__abc_22172_new_n5652_));
OR2X2 OR2X2_2206 ( .A(core__abc_22172_new_n5649_), .B(core__abc_22172_new_n5654_), .Y(core__abc_22172_new_n5655_));
OR2X2 OR2X2_2207 ( .A(core__abc_22172_new_n3217_), .B(core__abc_22172_new_n5655_), .Y(core__abc_22172_new_n5656_));
OR2X2 OR2X2_2208 ( .A(core__abc_22172_new_n5648_), .B(core__abc_22172_new_n5656_), .Y(core__abc_22172_new_n5657_));
OR2X2 OR2X2_2209 ( .A(core__abc_22172_new_n3228_), .B(core_v3_reg_43_), .Y(core__abc_22172_new_n5658_));
OR2X2 OR2X2_221 ( .A(_abc_19873_new_n1383_), .B(_abc_19873_new_n1384_), .Y(_abc_19873_new_n1385_));
OR2X2 OR2X2_2210 ( .A(core__abc_22172_new_n5637_), .B(core__abc_22172_new_n5628_), .Y(core__abc_22172_new_n5667_));
OR2X2 OR2X2_2211 ( .A(core__abc_22172_new_n5665_), .B(core__abc_22172_new_n5669_), .Y(core__abc_22172_new_n5670_));
OR2X2 OR2X2_2212 ( .A(core__abc_22172_new_n5673_), .B(core__abc_22172_new_n5670_), .Y(core__abc_22172_new_n5674_));
OR2X2 OR2X2_2213 ( .A(core__abc_22172_new_n5675_), .B(core__abc_22172_new_n2950_), .Y(core__abc_22172_new_n5676_));
OR2X2 OR2X2_2214 ( .A(core__abc_22172_new_n5679_), .B(core__abc_22172_new_n5677_), .Y(core__abc_22172_new_n5680_));
OR2X2 OR2X2_2215 ( .A(core__abc_22172_new_n5682_), .B(core__abc_22172_new_n5683_), .Y(core__abc_22172_new_n5684_));
OR2X2 OR2X2_2216 ( .A(core__abc_22172_new_n5516_), .B(core__abc_22172_new_n5689_), .Y(core__abc_22172_new_n5690_));
OR2X2 OR2X2_2217 ( .A(core__abc_22172_new_n5692_), .B(core__abc_22172_new_n5686_), .Y(core__abc_22172_new_n5693_));
OR2X2 OR2X2_2218 ( .A(core__abc_22172_new_n5696_), .B(core__abc_22172_new_n5694_), .Y(core__abc_22172_new_n5697_));
OR2X2 OR2X2_2219 ( .A(core_v3_reg_44_), .B(core_mi_44_), .Y(core__abc_22172_new_n5700_));
OR2X2 OR2X2_222 ( .A(_abc_19873_new_n1382_), .B(_abc_19873_new_n1385_), .Y(_abc_19873_new_n1386_));
OR2X2 OR2X2_2220 ( .A(core__abc_22172_new_n5699_), .B(core__abc_22172_new_n5704_), .Y(core__abc_22172_new_n5705_));
OR2X2 OR2X2_2221 ( .A(core__abc_22172_new_n5698_), .B(core__abc_22172_new_n5705_), .Y(core__abc_22172_new_n5706_));
OR2X2 OR2X2_2222 ( .A(core__abc_22172_new_n5707_), .B(core__abc_22172_new_n5661_), .Y(core__abc_22172_new_n5708_));
OR2X2 OR2X2_2223 ( .A(core__abc_22172_new_n5686_), .B(core__abc_22172_new_n5682_), .Y(core__abc_22172_new_n5711_));
OR2X2 OR2X2_2224 ( .A(core__abc_22172_new_n5677_), .B(core__abc_22172_new_n1477_), .Y(core__abc_22172_new_n5712_));
OR2X2 OR2X2_2225 ( .A(core__abc_22172_new_n5714_), .B(core__abc_22172_new_n5715_), .Y(core__abc_22172_new_n5716_));
OR2X2 OR2X2_2226 ( .A(core__abc_22172_new_n5718_), .B(core__abc_22172_new_n5719_), .Y(core__abc_22172_new_n5720_));
OR2X2 OR2X2_2227 ( .A(core__abc_22172_new_n5711_), .B(core__abc_22172_new_n5721_), .Y(core__abc_22172_new_n5722_));
OR2X2 OR2X2_2228 ( .A(core__abc_22172_new_n5723_), .B(core__abc_22172_new_n5720_), .Y(core__abc_22172_new_n5724_));
OR2X2 OR2X2_2229 ( .A(core__abc_22172_new_n5728_), .B(core__abc_22172_new_n5726_), .Y(core__abc_22172_new_n5729_));
OR2X2 OR2X2_223 ( .A(_abc_19873_new_n1386_), .B(_abc_19873_new_n1379_), .Y(_abc_19873_new_n1387_));
OR2X2 OR2X2_2230 ( .A(core_v3_reg_45_), .B(core_mi_45_), .Y(core__abc_22172_new_n5733_));
OR2X2 OR2X2_2231 ( .A(core__abc_22172_new_n5732_), .B(core__abc_22172_new_n5737_), .Y(core__abc_22172_new_n5738_));
OR2X2 OR2X2_2232 ( .A(core__abc_22172_new_n5730_), .B(core__abc_22172_new_n5738_), .Y(core__abc_22172_new_n5739_));
OR2X2 OR2X2_2233 ( .A(core__abc_22172_new_n5740_), .B(core__abc_22172_new_n5710_), .Y(core__abc_22172_new_n5741_));
OR2X2 OR2X2_2234 ( .A(core__abc_22172_new_n5718_), .B(core__abc_22172_new_n5682_), .Y(core__abc_22172_new_n5747_));
OR2X2 OR2X2_2235 ( .A(core__abc_22172_new_n5745_), .B(core__abc_22172_new_n5748_), .Y(core__abc_22172_new_n5749_));
OR2X2 OR2X2_2236 ( .A(core__abc_22172_new_n5750_), .B(core__abc_22172_new_n2954_), .Y(core__abc_22172_new_n5751_));
OR2X2 OR2X2_2237 ( .A(core__abc_22172_new_n5751_), .B(core__abc_22172_new_n1513_), .Y(core__abc_22172_new_n5754_));
OR2X2 OR2X2_2238 ( .A(core__abc_22172_new_n5757_), .B(core__abc_22172_new_n5758_), .Y(core__abc_22172_new_n5759_));
OR2X2 OR2X2_2239 ( .A(core__abc_22172_new_n5691_), .B(core__abc_22172_new_n5762_), .Y(core__abc_22172_new_n5763_));
OR2X2 OR2X2_224 ( .A(_abc_19873_new_n1389_), .B(_abc_19873_new_n1390_), .Y(_abc_19873_new_n1391_));
OR2X2 OR2X2_2240 ( .A(core__abc_22172_new_n5766_), .B(core__abc_22172_new_n5761_), .Y(core__abc_22172_new_n5767_));
OR2X2 OR2X2_2241 ( .A(core__abc_22172_new_n5770_), .B(core__abc_22172_new_n5768_), .Y(core__abc_22172_new_n5771_));
OR2X2 OR2X2_2242 ( .A(core_v3_reg_46_), .B(core_mi_46_), .Y(core__abc_22172_new_n5775_));
OR2X2 OR2X2_2243 ( .A(core__abc_22172_new_n5774_), .B(core__abc_22172_new_n5779_), .Y(core__abc_22172_new_n5780_));
OR2X2 OR2X2_2244 ( .A(core__abc_22172_new_n5772_), .B(core__abc_22172_new_n5780_), .Y(core__abc_22172_new_n5781_));
OR2X2 OR2X2_2245 ( .A(core__abc_22172_new_n5782_), .B(core__abc_22172_new_n5743_), .Y(core__abc_22172_new_n5783_));
OR2X2 OR2X2_2246 ( .A(core__abc_22172_new_n5761_), .B(core__abc_22172_new_n5758_), .Y(core__abc_22172_new_n5786_));
OR2X2 OR2X2_2247 ( .A(core__abc_22172_new_n5752_), .B(core__abc_22172_new_n1511_), .Y(core__abc_22172_new_n5787_));
OR2X2 OR2X2_2248 ( .A(core__abc_22172_new_n5787_), .B(core__abc_22172_new_n1530_), .Y(core__abc_22172_new_n5788_));
OR2X2 OR2X2_2249 ( .A(core__abc_22172_new_n5792_), .B(core__abc_22172_new_n5794_), .Y(core__abc_22172_new_n5795_));
OR2X2 OR2X2_225 ( .A(_abc_19873_new_n1391_), .B(_abc_19873_new_n1388_), .Y(_abc_19873_new_n1392_));
OR2X2 OR2X2_2250 ( .A(core__abc_22172_new_n5786_), .B(core__abc_22172_new_n5795_), .Y(core__abc_22172_new_n5796_));
OR2X2 OR2X2_2251 ( .A(core__abc_22172_new_n5765_), .B(core__abc_22172_new_n5759_), .Y(core__abc_22172_new_n5798_));
OR2X2 OR2X2_2252 ( .A(core__abc_22172_new_n3457_), .B(core__abc_22172_new_n5793_), .Y(core__abc_22172_new_n5800_));
OR2X2 OR2X2_2253 ( .A(core__abc_22172_new_n3452_), .B(core__abc_22172_new_n5791_), .Y(core__abc_22172_new_n5801_));
OR2X2 OR2X2_2254 ( .A(core__abc_22172_new_n5799_), .B(core__abc_22172_new_n5802_), .Y(core__abc_22172_new_n5803_));
OR2X2 OR2X2_2255 ( .A(core__abc_22172_new_n5804_), .B(core__abc_22172_new_n4804_), .Y(core__abc_22172_new_n5805_));
OR2X2 OR2X2_2256 ( .A(core__abc_22172_new_n5786_), .B(core__abc_22172_new_n5802_), .Y(core__abc_22172_new_n5806_));
OR2X2 OR2X2_2257 ( .A(core__abc_22172_new_n5799_), .B(core__abc_22172_new_n5795_), .Y(core__abc_22172_new_n5807_));
OR2X2 OR2X2_2258 ( .A(core__abc_22172_new_n5808_), .B(core__abc_22172_new_n4805_), .Y(core__abc_22172_new_n5809_));
OR2X2 OR2X2_2259 ( .A(core_v3_reg_47_), .B(core_mi_47_), .Y(core__abc_22172_new_n5813_));
OR2X2 OR2X2_226 ( .A(_abc_19873_new_n1393_), .B(_abc_19873_new_n1394_), .Y(_abc_19873_new_n1395_));
OR2X2 OR2X2_2260 ( .A(core__abc_22172_new_n5812_), .B(core__abc_22172_new_n5817_), .Y(core__abc_22172_new_n5818_));
OR2X2 OR2X2_2261 ( .A(core__abc_22172_new_n5811_), .B(core__abc_22172_new_n5818_), .Y(core__abc_22172_new_n5819_));
OR2X2 OR2X2_2262 ( .A(core__abc_22172_new_n5820_), .B(core__abc_22172_new_n5785_), .Y(core__abc_22172_new_n5821_));
OR2X2 OR2X2_2263 ( .A(core__abc_22172_new_n5792_), .B(core__abc_22172_new_n5758_), .Y(core__abc_22172_new_n5832_));
OR2X2 OR2X2_2264 ( .A(core__abc_22172_new_n5831_), .B(core__abc_22172_new_n5833_), .Y(core__abc_22172_new_n5834_));
OR2X2 OR2X2_2265 ( .A(core__abc_22172_new_n5834_), .B(core__abc_22172_new_n5830_), .Y(core__abc_22172_new_n5835_));
OR2X2 OR2X2_2266 ( .A(core__abc_22172_new_n5835_), .B(core__abc_22172_new_n5829_), .Y(core__abc_22172_new_n5836_));
OR2X2 OR2X2_2267 ( .A(core__abc_22172_new_n5828_), .B(core__abc_22172_new_n5836_), .Y(core__abc_22172_new_n5837_));
OR2X2 OR2X2_2268 ( .A(core__abc_22172_new_n5839_), .B(core__abc_22172_new_n5838_), .Y(core__abc_22172_new_n5840_));
OR2X2 OR2X2_2269 ( .A(core__abc_22172_new_n5842_), .B(core__abc_22172_new_n5843_), .Y(core__abc_22172_new_n5844_));
OR2X2 OR2X2_227 ( .A(_abc_19873_new_n1039_), .B(_abc_19873_new_n1395_), .Y(_abc_19873_new_n1396_));
OR2X2 OR2X2_2270 ( .A(core__abc_22172_new_n5139_), .B(core__abc_22172_new_n5847_), .Y(core__abc_22172_new_n5848_));
OR2X2 OR2X2_2271 ( .A(core__abc_22172_new_n5855_), .B(core__abc_22172_new_n5846_), .Y(core__abc_22172_new_n5856_));
OR2X2 OR2X2_2272 ( .A(core__abc_22172_new_n5859_), .B(core__abc_22172_new_n5857_), .Y(core__abc_22172_new_n5860_));
OR2X2 OR2X2_2273 ( .A(core_v3_reg_48_), .B(core_mi_48_), .Y(core__abc_22172_new_n5864_));
OR2X2 OR2X2_2274 ( .A(core__abc_22172_new_n5863_), .B(core__abc_22172_new_n5868_), .Y(core__abc_22172_new_n5869_));
OR2X2 OR2X2_2275 ( .A(core__abc_22172_new_n5861_), .B(core__abc_22172_new_n5869_), .Y(core__abc_22172_new_n5870_));
OR2X2 OR2X2_2276 ( .A(core__abc_22172_new_n5871_), .B(core__abc_22172_new_n5823_), .Y(core__abc_22172_new_n5872_));
OR2X2 OR2X2_2277 ( .A(core__abc_22172_new_n5838_), .B(core__abc_22172_new_n1545_), .Y(core__abc_22172_new_n5877_));
OR2X2 OR2X2_2278 ( .A(core__abc_22172_new_n5879_), .B(core__abc_22172_new_n5880_), .Y(core__abc_22172_new_n5881_));
OR2X2 OR2X2_2279 ( .A(core__abc_22172_new_n3586_), .B(core__abc_22172_new_n5881_), .Y(core__abc_22172_new_n5882_));
OR2X2 OR2X2_228 ( .A(_abc_19873_new_n1396_), .B(_abc_19873_new_n1392_), .Y(_abc_19873_new_n1397_));
OR2X2 OR2X2_2280 ( .A(core__abc_22172_new_n5883_), .B(core__abc_22172_new_n5884_), .Y(core__abc_22172_new_n5885_));
OR2X2 OR2X2_2281 ( .A(core__abc_22172_new_n5854_), .B(core__abc_22172_new_n5893_), .Y(core__abc_22172_new_n5894_));
OR2X2 OR2X2_2282 ( .A(core__abc_22172_new_n5898_), .B(core__abc_22172_new_n5899_), .Y(core__abc_22172_new_n5900_));
OR2X2 OR2X2_2283 ( .A(core_v3_reg_49_), .B(core_mi_49_), .Y(core__abc_22172_new_n5903_));
OR2X2 OR2X2_2284 ( .A(core__abc_22172_new_n5902_), .B(core__abc_22172_new_n5907_), .Y(core__abc_22172_new_n5908_));
OR2X2 OR2X2_2285 ( .A(core__abc_22172_new_n5901_), .B(core__abc_22172_new_n5908_), .Y(core__abc_22172_new_n5909_));
OR2X2 OR2X2_2286 ( .A(core__abc_22172_new_n5910_), .B(core__abc_22172_new_n5874_), .Y(core__abc_22172_new_n5911_));
OR2X2 OR2X2_2287 ( .A(core__abc_22172_new_n5916_), .B(core__abc_22172_new_n2978_), .Y(core__abc_22172_new_n5917_));
OR2X2 OR2X2_2288 ( .A(core__abc_22172_new_n5917_), .B(core__abc_22172_new_n1581_), .Y(core__abc_22172_new_n5920_));
OR2X2 OR2X2_2289 ( .A(core__abc_22172_new_n5922_), .B(core__abc_22172_new_n5924_), .Y(core__abc_22172_new_n5925_));
OR2X2 OR2X2_229 ( .A(_abc_19873_new_n1397_), .B(_abc_19873_new_n1387_), .Y(_abc_19873_new_n1398_));
OR2X2 OR2X2_2290 ( .A(core__abc_22172_new_n5915_), .B(core__abc_22172_new_n5925_), .Y(core__abc_22172_new_n5926_));
OR2X2 OR2X2_2291 ( .A(core__abc_22172_new_n5927_), .B(core__abc_22172_new_n5928_), .Y(core__abc_22172_new_n5929_));
OR2X2 OR2X2_2292 ( .A(core__abc_22172_new_n5932_), .B(core__abc_22172_new_n5930_), .Y(core__abc_22172_new_n5933_));
OR2X2 OR2X2_2293 ( .A(core_v3_reg_50_), .B(core_mi_50_), .Y(core__abc_22172_new_n5937_));
OR2X2 OR2X2_2294 ( .A(core__abc_22172_new_n5936_), .B(core__abc_22172_new_n5941_), .Y(core__abc_22172_new_n5942_));
OR2X2 OR2X2_2295 ( .A(core__abc_22172_new_n5934_), .B(core__abc_22172_new_n5942_), .Y(core__abc_22172_new_n5943_));
OR2X2 OR2X2_2296 ( .A(core__abc_22172_new_n5944_), .B(core__abc_22172_new_n5913_), .Y(core__abc_22172_new_n5945_));
OR2X2 OR2X2_2297 ( .A(core__abc_22172_new_n5918_), .B(core__abc_22172_new_n1579_), .Y(core__abc_22172_new_n5950_));
OR2X2 OR2X2_2298 ( .A(core__abc_22172_new_n5950_), .B(core__abc_22172_new_n1598_), .Y(core__abc_22172_new_n5951_));
OR2X2 OR2X2_2299 ( .A(core__abc_22172_new_n3716_), .B(core__abc_22172_new_n5955_), .Y(core__abc_22172_new_n5956_));
OR2X2 OR2X2_23 ( .A(_abc_19873_new_n961_), .B(_abc_19873_new_n954_), .Y(_abc_19873_new_n962_));
OR2X2 OR2X2_230 ( .A(_abc_19873_new_n1400_), .B(_abc_19873_new_n1401_), .Y(_abc_19873_new_n1402_));
OR2X2 OR2X2_2300 ( .A(core__abc_22172_new_n5949_), .B(core__abc_22172_new_n5960_), .Y(core__abc_22172_new_n5963_));
OR2X2 OR2X2_2301 ( .A(core__abc_22172_new_n5967_), .B(core__abc_22172_new_n5965_), .Y(core__abc_22172_new_n5968_));
OR2X2 OR2X2_2302 ( .A(core_v3_reg_51_), .B(core_mi_51_), .Y(core__abc_22172_new_n5971_));
OR2X2 OR2X2_2303 ( .A(core__abc_22172_new_n5970_), .B(core__abc_22172_new_n5975_), .Y(core__abc_22172_new_n5976_));
OR2X2 OR2X2_2304 ( .A(core__abc_22172_new_n5969_), .B(core__abc_22172_new_n5976_), .Y(core__abc_22172_new_n5977_));
OR2X2 OR2X2_2305 ( .A(core__abc_22172_new_n5978_), .B(core__abc_22172_new_n5947_), .Y(core__abc_22172_new_n5979_));
OR2X2 OR2X2_2306 ( .A(core__abc_22172_new_n5957_), .B(core__abc_22172_new_n5948_), .Y(core__abc_22172_new_n5986_));
OR2X2 OR2X2_2307 ( .A(core__abc_22172_new_n5985_), .B(core__abc_22172_new_n5988_), .Y(core__abc_22172_new_n5989_));
OR2X2 OR2X2_2308 ( .A(core__abc_22172_new_n5991_), .B(core__abc_22172_new_n5989_), .Y(core__abc_22172_new_n5992_));
OR2X2 OR2X2_2309 ( .A(core__abc_22172_new_n5993_), .B(core__abc_22172_new_n2982_), .Y(core__abc_22172_new_n5994_));
OR2X2 OR2X2_231 ( .A(_abc_19873_new_n1038_), .B(_abc_19873_new_n1403_), .Y(_abc_19873_new_n1404_));
OR2X2 OR2X2_2310 ( .A(core__abc_22172_new_n5997_), .B(core__abc_22172_new_n5995_), .Y(core__abc_22172_new_n5998_));
OR2X2 OR2X2_2311 ( .A(core__abc_22172_new_n6000_), .B(core__abc_22172_new_n6001_), .Y(core__abc_22172_new_n6002_));
OR2X2 OR2X2_2312 ( .A(core__abc_22172_new_n5854_), .B(core__abc_22172_new_n6006_), .Y(core__abc_22172_new_n6007_));
OR2X2 OR2X2_2313 ( .A(core__abc_22172_new_n6009_), .B(core__abc_22172_new_n6004_), .Y(core__abc_22172_new_n6010_));
OR2X2 OR2X2_2314 ( .A(core__abc_22172_new_n6013_), .B(core__abc_22172_new_n6011_), .Y(core__abc_22172_new_n6014_));
OR2X2 OR2X2_2315 ( .A(core_v3_reg_52_), .B(core_mi_52_), .Y(core__abc_22172_new_n6017_));
OR2X2 OR2X2_2316 ( .A(core__abc_22172_new_n6016_), .B(core__abc_22172_new_n6021_), .Y(core__abc_22172_new_n6022_));
OR2X2 OR2X2_2317 ( .A(core__abc_22172_new_n6015_), .B(core__abc_22172_new_n6022_), .Y(core__abc_22172_new_n6023_));
OR2X2 OR2X2_2318 ( .A(core__abc_22172_new_n6024_), .B(core__abc_22172_new_n5981_), .Y(core__abc_22172_new_n6025_));
OR2X2 OR2X2_2319 ( .A(core__abc_22172_new_n6004_), .B(core__abc_22172_new_n6000_), .Y(core__abc_22172_new_n6028_));
OR2X2 OR2X2_232 ( .A(_abc_19873_new_n1404_), .B(_abc_19873_new_n1402_), .Y(_abc_19873_new_n1405_));
OR2X2 OR2X2_2320 ( .A(core__abc_22172_new_n5995_), .B(core__abc_22172_new_n1613_), .Y(core__abc_22172_new_n6029_));
OR2X2 OR2X2_2321 ( .A(core__abc_22172_new_n6031_), .B(core__abc_22172_new_n6032_), .Y(core__abc_22172_new_n6033_));
OR2X2 OR2X2_2322 ( .A(core__abc_22172_new_n6035_), .B(core__abc_22172_new_n6036_), .Y(core__abc_22172_new_n6037_));
OR2X2 OR2X2_2323 ( .A(core__abc_22172_new_n6028_), .B(core__abc_22172_new_n6038_), .Y(core__abc_22172_new_n6039_));
OR2X2 OR2X2_2324 ( .A(core__abc_22172_new_n6040_), .B(core__abc_22172_new_n6037_), .Y(core__abc_22172_new_n6041_));
OR2X2 OR2X2_2325 ( .A(core__abc_22172_new_n6043_), .B(core__abc_22172_new_n5113_), .Y(core__abc_22172_new_n6044_));
OR2X2 OR2X2_2326 ( .A(core__abc_22172_new_n6042_), .B(core__abc_22172_new_n5114_), .Y(core__abc_22172_new_n6045_));
OR2X2 OR2X2_2327 ( .A(core_v3_reg_53_), .B(core_mi_53_), .Y(core__abc_22172_new_n6050_));
OR2X2 OR2X2_2328 ( .A(core__abc_22172_new_n6049_), .B(core__abc_22172_new_n6054_), .Y(core__abc_22172_new_n6055_));
OR2X2 OR2X2_2329 ( .A(core__abc_22172_new_n6047_), .B(core__abc_22172_new_n6055_), .Y(core__abc_22172_new_n6056_));
OR2X2 OR2X2_233 ( .A(_abc_19873_new_n1407_), .B(_abc_19873_new_n1408_), .Y(_abc_19873_new_n1409_));
OR2X2 OR2X2_2330 ( .A(core__abc_22172_new_n6057_), .B(core__abc_22172_new_n6027_), .Y(core__abc_22172_new_n6058_));
OR2X2 OR2X2_2331 ( .A(core__abc_22172_new_n6035_), .B(core__abc_22172_new_n6000_), .Y(core__abc_22172_new_n6064_));
OR2X2 OR2X2_2332 ( .A(core__abc_22172_new_n6062_), .B(core__abc_22172_new_n6065_), .Y(core__abc_22172_new_n6066_));
OR2X2 OR2X2_2333 ( .A(core__abc_22172_new_n6067_), .B(core__abc_22172_new_n2987_), .Y(core__abc_22172_new_n6068_));
OR2X2 OR2X2_2334 ( .A(core__abc_22172_new_n6071_), .B(core__abc_22172_new_n6069_), .Y(core__abc_22172_new_n6072_));
OR2X2 OR2X2_2335 ( .A(core__abc_22172_new_n6074_), .B(core__abc_22172_new_n6075_), .Y(core__abc_22172_new_n6076_));
OR2X2 OR2X2_2336 ( .A(core__abc_22172_new_n6008_), .B(core__abc_22172_new_n6079_), .Y(core__abc_22172_new_n6080_));
OR2X2 OR2X2_2337 ( .A(core__abc_22172_new_n6083_), .B(core__abc_22172_new_n6078_), .Y(core__abc_22172_new_n6084_));
OR2X2 OR2X2_2338 ( .A(core__abc_22172_new_n6087_), .B(core__abc_22172_new_n6085_), .Y(core__abc_22172_new_n6088_));
OR2X2 OR2X2_2339 ( .A(core_v3_reg_54_), .B(core_mi_54_), .Y(core__abc_22172_new_n6092_));
OR2X2 OR2X2_234 ( .A(_abc_19873_new_n1409_), .B(_abc_19873_new_n1406_), .Y(_abc_19873_new_n1410_));
OR2X2 OR2X2_2340 ( .A(core__abc_22172_new_n6091_), .B(core__abc_22172_new_n6096_), .Y(core__abc_22172_new_n6097_));
OR2X2 OR2X2_2341 ( .A(core__abc_22172_new_n6089_), .B(core__abc_22172_new_n6097_), .Y(core__abc_22172_new_n6098_));
OR2X2 OR2X2_2342 ( .A(core__abc_22172_new_n6099_), .B(core__abc_22172_new_n6060_), .Y(core__abc_22172_new_n6100_));
OR2X2 OR2X2_2343 ( .A(core__abc_22172_new_n6078_), .B(core__abc_22172_new_n6074_), .Y(core__abc_22172_new_n6103_));
OR2X2 OR2X2_2344 ( .A(core__abc_22172_new_n6069_), .B(core__abc_22172_new_n1647_), .Y(core__abc_22172_new_n6104_));
OR2X2 OR2X2_2345 ( .A(core__abc_22172_new_n6106_), .B(core__abc_22172_new_n6107_), .Y(core__abc_22172_new_n6108_));
OR2X2 OR2X2_2346 ( .A(core__abc_22172_new_n6110_), .B(core__abc_22172_new_n6111_), .Y(core__abc_22172_new_n6112_));
OR2X2 OR2X2_2347 ( .A(core__abc_22172_new_n6103_), .B(core__abc_22172_new_n6112_), .Y(core__abc_22172_new_n6113_));
OR2X2 OR2X2_2348 ( .A(core__abc_22172_new_n6082_), .B(core__abc_22172_new_n6076_), .Y(core__abc_22172_new_n6115_));
OR2X2 OR2X2_2349 ( .A(core__abc_22172_new_n3980_), .B(core__abc_22172_new_n6108_), .Y(core__abc_22172_new_n6117_));
OR2X2 OR2X2_235 ( .A(_abc_19873_new_n1411_), .B(_abc_19873_new_n1412_), .Y(_abc_19873_new_n1413_));
OR2X2 OR2X2_2350 ( .A(core__abc_22172_new_n6116_), .B(core__abc_22172_new_n6119_), .Y(core__abc_22172_new_n6120_));
OR2X2 OR2X2_2351 ( .A(core__abc_22172_new_n6121_), .B(core__abc_22172_new_n5221_), .Y(core__abc_22172_new_n6122_));
OR2X2 OR2X2_2352 ( .A(core__abc_22172_new_n6103_), .B(core__abc_22172_new_n6119_), .Y(core__abc_22172_new_n6123_));
OR2X2 OR2X2_2353 ( .A(core__abc_22172_new_n6116_), .B(core__abc_22172_new_n6112_), .Y(core__abc_22172_new_n6124_));
OR2X2 OR2X2_2354 ( .A(core__abc_22172_new_n6125_), .B(core__abc_22172_new_n5222_), .Y(core__abc_22172_new_n6126_));
OR2X2 OR2X2_2355 ( .A(core_v3_reg_55_), .B(core_mi_55_), .Y(core__abc_22172_new_n6130_));
OR2X2 OR2X2_2356 ( .A(core__abc_22172_new_n6129_), .B(core__abc_22172_new_n6134_), .Y(core__abc_22172_new_n6135_));
OR2X2 OR2X2_2357 ( .A(core__abc_22172_new_n6128_), .B(core__abc_22172_new_n6135_), .Y(core__abc_22172_new_n6136_));
OR2X2 OR2X2_2358 ( .A(core__abc_22172_new_n6137_), .B(core__abc_22172_new_n6102_), .Y(core__abc_22172_new_n6138_));
OR2X2 OR2X2_2359 ( .A(core__abc_22172_new_n6111_), .B(core__abc_22172_new_n6114_), .Y(core__abc_22172_new_n6148_));
OR2X2 OR2X2_236 ( .A(_abc_19873_new_n1414_), .B(_abc_19873_new_n1415_), .Y(_abc_19873_new_n1416_));
OR2X2 OR2X2_2360 ( .A(core__abc_22172_new_n6147_), .B(core__abc_22172_new_n6150_), .Y(core__abc_22172_new_n6151_));
OR2X2 OR2X2_2361 ( .A(core__abc_22172_new_n6151_), .B(core__abc_22172_new_n6146_), .Y(core__abc_22172_new_n6152_));
OR2X2 OR2X2_2362 ( .A(core__abc_22172_new_n6145_), .B(core__abc_22172_new_n6152_), .Y(core__abc_22172_new_n6153_));
OR2X2 OR2X2_2363 ( .A(core__abc_22172_new_n6154_), .B(core__abc_22172_new_n2992_), .Y(core__abc_22172_new_n6155_));
OR2X2 OR2X2_2364 ( .A(core__abc_22172_new_n6158_), .B(core__abc_22172_new_n6156_), .Y(core__abc_22172_new_n6159_));
OR2X2 OR2X2_2365 ( .A(core__abc_22172_new_n6162_), .B(core__abc_22172_new_n6161_), .Y(core__abc_22172_new_n6163_));
OR2X2 OR2X2_2366 ( .A(core__abc_22172_new_n6112_), .B(core__abc_22172_new_n6076_), .Y(core__abc_22172_new_n6166_));
OR2X2 OR2X2_2367 ( .A(core__abc_22172_new_n6166_), .B(core__abc_22172_new_n6079_), .Y(core__abc_22172_new_n6167_));
OR2X2 OR2X2_2368 ( .A(core__abc_22172_new_n6167_), .B(core__abc_22172_new_n6006_), .Y(core__abc_22172_new_n6168_));
OR2X2 OR2X2_2369 ( .A(core__abc_22172_new_n5854_), .B(core__abc_22172_new_n6168_), .Y(core__abc_22172_new_n6169_));
OR2X2 OR2X2_237 ( .A(_abc_19873_new_n1413_), .B(_abc_19873_new_n1416_), .Y(_abc_19873_new_n1417_));
OR2X2 OR2X2_2370 ( .A(core__abc_22172_new_n6167_), .B(core__abc_22172_new_n6005_), .Y(core__abc_22172_new_n6170_));
OR2X2 OR2X2_2371 ( .A(core__abc_22172_new_n6166_), .B(core__abc_22172_new_n6081_), .Y(core__abc_22172_new_n6171_));
OR2X2 OR2X2_2372 ( .A(core__abc_22172_new_n6175_), .B(core__abc_22172_new_n6165_), .Y(core__abc_22172_new_n6176_));
OR2X2 OR2X2_2373 ( .A(core__abc_22172_new_n6179_), .B(core__abc_22172_new_n6177_), .Y(core__abc_22172_new_n6180_));
OR2X2 OR2X2_2374 ( .A(core_v3_reg_56_), .B(core_mi_56_), .Y(core__abc_22172_new_n6183_));
OR2X2 OR2X2_2375 ( .A(core__abc_22172_new_n6182_), .B(core__abc_22172_new_n6187_), .Y(core__abc_22172_new_n6188_));
OR2X2 OR2X2_2376 ( .A(core__abc_22172_new_n6181_), .B(core__abc_22172_new_n6188_), .Y(core__abc_22172_new_n6189_));
OR2X2 OR2X2_2377 ( .A(core__abc_22172_new_n6190_), .B(core__abc_22172_new_n6140_), .Y(core__abc_22172_new_n6191_));
OR2X2 OR2X2_2378 ( .A(core__abc_22172_new_n6165_), .B(core__abc_22172_new_n6161_), .Y(core__abc_22172_new_n6194_));
OR2X2 OR2X2_2379 ( .A(core__abc_22172_new_n6156_), .B(core__abc_22172_new_n1681_), .Y(core__abc_22172_new_n6195_));
OR2X2 OR2X2_238 ( .A(_abc_19873_new_n1417_), .B(_abc_19873_new_n1410_), .Y(_abc_19873_new_n1418_));
OR2X2 OR2X2_2380 ( .A(core__abc_22172_new_n6197_), .B(core__abc_22172_new_n6198_), .Y(core__abc_22172_new_n6199_));
OR2X2 OR2X2_2381 ( .A(core__abc_22172_new_n6201_), .B(core__abc_22172_new_n6202_), .Y(core__abc_22172_new_n6203_));
OR2X2 OR2X2_2382 ( .A(core__abc_22172_new_n6194_), .B(core__abc_22172_new_n6204_), .Y(core__abc_22172_new_n6205_));
OR2X2 OR2X2_2383 ( .A(core__abc_22172_new_n6206_), .B(core__abc_22172_new_n6203_), .Y(core__abc_22172_new_n6207_));
OR2X2 OR2X2_2384 ( .A(core__abc_22172_new_n6209_), .B(core__abc_22172_new_n5316_), .Y(core__abc_22172_new_n6210_));
OR2X2 OR2X2_2385 ( .A(core__abc_22172_new_n6208_), .B(core__abc_22172_new_n5317_), .Y(core__abc_22172_new_n6211_));
OR2X2 OR2X2_2386 ( .A(core_v3_reg_57_), .B(core_mi_57_), .Y(core__abc_22172_new_n6215_));
OR2X2 OR2X2_2387 ( .A(core__abc_22172_new_n6214_), .B(core__abc_22172_new_n6219_), .Y(core__abc_22172_new_n6220_));
OR2X2 OR2X2_2388 ( .A(core__abc_22172_new_n6213_), .B(core__abc_22172_new_n6220_), .Y(core__abc_22172_new_n6221_));
OR2X2 OR2X2_2389 ( .A(core__abc_22172_new_n6222_), .B(core__abc_22172_new_n6193_), .Y(core__abc_22172_new_n6223_));
OR2X2 OR2X2_239 ( .A(_abc_19873_new_n1418_), .B(_abc_19873_new_n1405_), .Y(_abc_19873_new_n1419_));
OR2X2 OR2X2_2390 ( .A(core__abc_22172_new_n6202_), .B(core__abc_22172_new_n6228_), .Y(core__abc_22172_new_n6229_));
OR2X2 OR2X2_2391 ( .A(core__abc_22172_new_n6233_), .B(core__abc_22172_new_n6231_), .Y(core__abc_22172_new_n6234_));
OR2X2 OR2X2_2392 ( .A(core__abc_22172_new_n6157_), .B(core__abc_22172_new_n6235_), .Y(core__abc_22172_new_n6236_));
OR2X2 OR2X2_2393 ( .A(core__abc_22172_new_n6237_), .B(core__abc_22172_new_n1723_), .Y(core__abc_22172_new_n6238_));
OR2X2 OR2X2_2394 ( .A(core__abc_22172_new_n6239_), .B(core__abc_22172_new_n6240_), .Y(core__abc_22172_new_n6241_));
OR2X2 OR2X2_2395 ( .A(core__abc_22172_new_n6243_), .B(core__abc_22172_new_n6244_), .Y(core__abc_22172_new_n6245_));
OR2X2 OR2X2_2396 ( .A(core__abc_22172_new_n6234_), .B(core__abc_22172_new_n6246_), .Y(core__abc_22172_new_n6249_));
OR2X2 OR2X2_2397 ( .A(core__abc_22172_new_n6252_), .B(core__abc_22172_new_n6253_), .Y(core__abc_22172_new_n6254_));
OR2X2 OR2X2_2398 ( .A(core_v3_reg_58_), .B(core_mi_58_), .Y(core__abc_22172_new_n6258_));
OR2X2 OR2X2_2399 ( .A(core__abc_22172_new_n6257_), .B(core__abc_22172_new_n6262_), .Y(core__abc_22172_new_n6263_));
OR2X2 OR2X2_24 ( .A(_abc_19873_new_n949_), .B(_abc_19873_new_n962_), .Y(_abc_19873_new_n963_));
OR2X2 OR2X2_240 ( .A(_abc_19873_new_n1421_), .B(_abc_19873_new_n1422_), .Y(_abc_19873_new_n1423_));
OR2X2 OR2X2_2400 ( .A(core__abc_22172_new_n6255_), .B(core__abc_22172_new_n6263_), .Y(core__abc_22172_new_n6264_));
OR2X2 OR2X2_2401 ( .A(core__abc_22172_new_n6265_), .B(core__abc_22172_new_n6225_), .Y(core__abc_22172_new_n6266_));
OR2X2 OR2X2_2402 ( .A(core__abc_22172_new_n6271_), .B(core__abc_22172_new_n1740_), .Y(core__abc_22172_new_n6274_));
OR2X2 OR2X2_2403 ( .A(core__abc_22172_new_n4255_), .B(core__abc_22172_new_n6276_), .Y(core__abc_22172_new_n6277_));
OR2X2 OR2X2_2404 ( .A(core__abc_22172_new_n4251_), .B(core__abc_22172_new_n6275_), .Y(core__abc_22172_new_n6278_));
OR2X2 OR2X2_2405 ( .A(core__abc_22172_new_n6270_), .B(core__abc_22172_new_n6279_), .Y(core__abc_22172_new_n6280_));
OR2X2 OR2X2_2406 ( .A(core__abc_22172_new_n6282_), .B(core__abc_22172_new_n6281_), .Y(core__abc_22172_new_n6283_));
OR2X2 OR2X2_2407 ( .A(core__abc_22172_new_n6269_), .B(core__abc_22172_new_n6283_), .Y(core__abc_22172_new_n6284_));
OR2X2 OR2X2_2408 ( .A(core__abc_22172_new_n6286_), .B(core__abc_22172_new_n5413_), .Y(core__abc_22172_new_n6287_));
OR2X2 OR2X2_2409 ( .A(core__abc_22172_new_n6285_), .B(core__abc_22172_new_n5412_), .Y(core__abc_22172_new_n6288_));
OR2X2 OR2X2_241 ( .A(_abc_19873_new_n1425_), .B(_abc_19873_new_n1426_), .Y(_abc_19873_new_n1427_));
OR2X2 OR2X2_2410 ( .A(core_v3_reg_59_), .B(core_mi_59_), .Y(core__abc_22172_new_n6294_));
OR2X2 OR2X2_2411 ( .A(core__abc_22172_new_n6291_), .B(core__abc_22172_new_n6296_), .Y(core__abc_22172_new_n6297_));
OR2X2 OR2X2_2412 ( .A(core__abc_22172_new_n3217_), .B(core__abc_22172_new_n6297_), .Y(core__abc_22172_new_n6298_));
OR2X2 OR2X2_2413 ( .A(core__abc_22172_new_n6290_), .B(core__abc_22172_new_n6298_), .Y(core__abc_22172_new_n6299_));
OR2X2 OR2X2_2414 ( .A(core__abc_22172_new_n3228_), .B(core_v3_reg_59_), .Y(core__abc_22172_new_n6300_));
OR2X2 OR2X2_2415 ( .A(core__abc_22172_new_n6282_), .B(core__abc_22172_new_n6268_), .Y(core__abc_22172_new_n6308_));
OR2X2 OR2X2_2416 ( .A(core__abc_22172_new_n6307_), .B(core__abc_22172_new_n6310_), .Y(core__abc_22172_new_n6311_));
OR2X2 OR2X2_2417 ( .A(core__abc_22172_new_n6306_), .B(core__abc_22172_new_n6311_), .Y(core__abc_22172_new_n6312_));
OR2X2 OR2X2_2418 ( .A(core__abc_22172_new_n6313_), .B(core__abc_22172_new_n3001_), .Y(core__abc_22172_new_n6314_));
OR2X2 OR2X2_2419 ( .A(core__abc_22172_new_n6317_), .B(core__abc_22172_new_n6315_), .Y(core__abc_22172_new_n6318_));
OR2X2 OR2X2_242 ( .A(_abc_19873_new_n1427_), .B(_abc_19873_new_n1424_), .Y(_abc_19873_new_n1428_));
OR2X2 OR2X2_2420 ( .A(core__abc_22172_new_n6321_), .B(core__abc_22172_new_n6320_), .Y(core__abc_22172_new_n6322_));
OR2X2 OR2X2_2421 ( .A(core__abc_22172_new_n6283_), .B(core__abc_22172_new_n6245_), .Y(core__abc_22172_new_n6326_));
OR2X2 OR2X2_2422 ( .A(core__abc_22172_new_n6326_), .B(core__abc_22172_new_n6325_), .Y(core__abc_22172_new_n6327_));
OR2X2 OR2X2_2423 ( .A(core__abc_22172_new_n6174_), .B(core__abc_22172_new_n6327_), .Y(core__abc_22172_new_n6328_));
OR2X2 OR2X2_2424 ( .A(core__abc_22172_new_n6332_), .B(core__abc_22172_new_n6324_), .Y(core__abc_22172_new_n6333_));
OR2X2 OR2X2_2425 ( .A(core__abc_22172_new_n6336_), .B(core__abc_22172_new_n6334_), .Y(core__abc_22172_new_n6337_));
OR2X2 OR2X2_2426 ( .A(core_v3_reg_60_), .B(core_mi_60_), .Y(core__abc_22172_new_n6341_));
OR2X2 OR2X2_2427 ( .A(core__abc_22172_new_n6340_), .B(core__abc_22172_new_n6345_), .Y(core__abc_22172_new_n6346_));
OR2X2 OR2X2_2428 ( .A(core__abc_22172_new_n6338_), .B(core__abc_22172_new_n6346_), .Y(core__abc_22172_new_n6347_));
OR2X2 OR2X2_2429 ( .A(core__abc_22172_new_n6348_), .B(core__abc_22172_new_n6303_), .Y(core__abc_22172_new_n6349_));
OR2X2 OR2X2_243 ( .A(_abc_19873_new_n1428_), .B(_abc_19873_new_n1423_), .Y(_abc_19873_new_n1429_));
OR2X2 OR2X2_2430 ( .A(core__abc_22172_new_n6324_), .B(core__abc_22172_new_n6320_), .Y(core__abc_22172_new_n6352_));
OR2X2 OR2X2_2431 ( .A(core__abc_22172_new_n6315_), .B(core__abc_22172_new_n1749_), .Y(core__abc_22172_new_n6353_));
OR2X2 OR2X2_2432 ( .A(core__abc_22172_new_n6355_), .B(core__abc_22172_new_n6356_), .Y(core__abc_22172_new_n6357_));
OR2X2 OR2X2_2433 ( .A(core__abc_22172_new_n6359_), .B(core__abc_22172_new_n6360_), .Y(core__abc_22172_new_n6361_));
OR2X2 OR2X2_2434 ( .A(core__abc_22172_new_n6352_), .B(core__abc_22172_new_n6361_), .Y(core__abc_22172_new_n6362_));
OR2X2 OR2X2_2435 ( .A(core__abc_22172_new_n6331_), .B(core__abc_22172_new_n6322_), .Y(core__abc_22172_new_n6364_));
OR2X2 OR2X2_2436 ( .A(core__abc_22172_new_n4376_), .B(core__abc_22172_new_n6357_), .Y(core__abc_22172_new_n6366_));
OR2X2 OR2X2_2437 ( .A(core__abc_22172_new_n6365_), .B(core__abc_22172_new_n6368_), .Y(core__abc_22172_new_n6369_));
OR2X2 OR2X2_2438 ( .A(core__abc_22172_new_n6370_), .B(core__abc_22172_new_n5506_), .Y(core__abc_22172_new_n6371_));
OR2X2 OR2X2_2439 ( .A(core__abc_22172_new_n6352_), .B(core__abc_22172_new_n6368_), .Y(core__abc_22172_new_n6372_));
OR2X2 OR2X2_244 ( .A(_abc_19873_new_n1431_), .B(_abc_19873_new_n1432_), .Y(_abc_19873_new_n1433_));
OR2X2 OR2X2_2440 ( .A(core__abc_22172_new_n6365_), .B(core__abc_22172_new_n6361_), .Y(core__abc_22172_new_n6373_));
OR2X2 OR2X2_2441 ( .A(core__abc_22172_new_n6374_), .B(core__abc_22172_new_n5507_), .Y(core__abc_22172_new_n6375_));
OR2X2 OR2X2_2442 ( .A(core_v3_reg_61_), .B(core_mi_61_), .Y(core__abc_22172_new_n6380_));
OR2X2 OR2X2_2443 ( .A(core__abc_22172_new_n6379_), .B(core__abc_22172_new_n6384_), .Y(core__abc_22172_new_n6385_));
OR2X2 OR2X2_2444 ( .A(core__abc_22172_new_n6377_), .B(core__abc_22172_new_n6385_), .Y(core__abc_22172_new_n6386_));
OR2X2 OR2X2_2445 ( .A(core__abc_22172_new_n6387_), .B(core__abc_22172_new_n6351_), .Y(core__abc_22172_new_n6388_));
OR2X2 OR2X2_2446 ( .A(core__abc_22172_new_n6361_), .B(core__abc_22172_new_n6322_), .Y(core__abc_22172_new_n6391_));
OR2X2 OR2X2_2447 ( .A(core__abc_22172_new_n6331_), .B(core__abc_22172_new_n6391_), .Y(core__abc_22172_new_n6392_));
OR2X2 OR2X2_2448 ( .A(core__abc_22172_new_n6393_), .B(core__abc_22172_new_n6359_), .Y(core__abc_22172_new_n6394_));
OR2X2 OR2X2_2449 ( .A(core__abc_22172_new_n6397_), .B(core__abc_22172_new_n3008_), .Y(core__abc_22172_new_n6398_));
OR2X2 OR2X2_245 ( .A(_abc_19873_new_n1434_), .B(_abc_19873_new_n1435_), .Y(_abc_19873_new_n1436_));
OR2X2 OR2X2_2450 ( .A(core__abc_22172_new_n6401_), .B(core__abc_22172_new_n6399_), .Y(core__abc_22172_new_n6402_));
OR2X2 OR2X2_2451 ( .A(core__abc_22172_new_n6404_), .B(core__abc_22172_new_n6405_), .Y(core__abc_22172_new_n6406_));
OR2X2 OR2X2_2452 ( .A(core__abc_22172_new_n6409_), .B(core__abc_22172_new_n6394_), .Y(core__abc_22172_new_n6410_));
OR2X2 OR2X2_2453 ( .A(core__abc_22172_new_n6407_), .B(core__abc_22172_new_n6412_), .Y(core__abc_22172_new_n6413_));
OR2X2 OR2X2_2454 ( .A(core__abc_22172_new_n6413_), .B(core__abc_22172_new_n5556_), .Y(core__abc_22172_new_n6414_));
OR2X2 OR2X2_2455 ( .A(core__abc_22172_new_n6410_), .B(core__abc_22172_new_n6411_), .Y(core__abc_22172_new_n6415_));
OR2X2 OR2X2_2456 ( .A(core__abc_22172_new_n6396_), .B(core__abc_22172_new_n6406_), .Y(core__abc_22172_new_n6416_));
OR2X2 OR2X2_2457 ( .A(core__abc_22172_new_n6417_), .B(core__abc_22172_new_n5557_), .Y(core__abc_22172_new_n6418_));
OR2X2 OR2X2_2458 ( .A(core_v3_reg_62_), .B(core_mi_62_), .Y(core__abc_22172_new_n6423_));
OR2X2 OR2X2_2459 ( .A(core__abc_22172_new_n6422_), .B(core__abc_22172_new_n6427_), .Y(core__abc_22172_new_n6428_));
OR2X2 OR2X2_246 ( .A(_abc_19873_new_n1433_), .B(_abc_19873_new_n1436_), .Y(_abc_19873_new_n1437_));
OR2X2 OR2X2_2460 ( .A(core__abc_22172_new_n6420_), .B(core__abc_22172_new_n6428_), .Y(core__abc_22172_new_n6429_));
OR2X2 OR2X2_2461 ( .A(core__abc_22172_new_n6430_), .B(core__abc_22172_new_n6390_), .Y(core__abc_22172_new_n6431_));
OR2X2 OR2X2_2462 ( .A(core__abc_22172_new_n6412_), .B(core__abc_22172_new_n6404_), .Y(core__abc_22172_new_n6433_));
OR2X2 OR2X2_2463 ( .A(core__abc_22172_new_n6399_), .B(core__abc_22172_new_n1783_), .Y(core__abc_22172_new_n6434_));
OR2X2 OR2X2_2464 ( .A(core__abc_22172_new_n6436_), .B(core__abc_22172_new_n6437_), .Y(core__abc_22172_new_n6438_));
OR2X2 OR2X2_2465 ( .A(core__abc_22172_new_n6440_), .B(core__abc_22172_new_n6441_), .Y(core__abc_22172_new_n6442_));
OR2X2 OR2X2_2466 ( .A(core__abc_22172_new_n6433_), .B(core__abc_22172_new_n6442_), .Y(core__abc_22172_new_n6443_));
OR2X2 OR2X2_2467 ( .A(core__abc_22172_new_n6445_), .B(core__abc_22172_new_n6446_), .Y(core__abc_22172_new_n6447_));
OR2X2 OR2X2_2468 ( .A(core__abc_22172_new_n6448_), .B(core__abc_22172_new_n5599_), .Y(core__abc_22172_new_n6449_));
OR2X2 OR2X2_2469 ( .A(core__abc_22172_new_n6433_), .B(core__abc_22172_new_n6446_), .Y(core__abc_22172_new_n6450_));
OR2X2 OR2X2_247 ( .A(_abc_19873_new_n1437_), .B(_abc_19873_new_n1430_), .Y(_abc_19873_new_n1438_));
OR2X2 OR2X2_2470 ( .A(core__abc_22172_new_n6445_), .B(core__abc_22172_new_n6442_), .Y(core__abc_22172_new_n6451_));
OR2X2 OR2X2_2471 ( .A(core__abc_22172_new_n6452_), .B(core__abc_22172_new_n5598_), .Y(core__abc_22172_new_n6453_));
OR2X2 OR2X2_2472 ( .A(core_v3_reg_63_), .B(core_mi_63_), .Y(core__abc_22172_new_n6459_));
OR2X2 OR2X2_2473 ( .A(core__abc_22172_new_n6456_), .B(core__abc_22172_new_n6461_), .Y(core__abc_22172_new_n6462_));
OR2X2 OR2X2_2474 ( .A(core__abc_22172_new_n3217_), .B(core__abc_22172_new_n6462_), .Y(core__abc_22172_new_n6463_));
OR2X2 OR2X2_2475 ( .A(core__abc_22172_new_n6455_), .B(core__abc_22172_new_n6463_), .Y(core__abc_22172_new_n6464_));
OR2X2 OR2X2_2476 ( .A(core__abc_22172_new_n3228_), .B(core_v3_reg_63_), .Y(core__abc_22172_new_n6465_));
OR2X2 OR2X2_2477 ( .A(core__abc_22172_new_n6470_), .B(core__abc_22172_new_n6469_), .Y(core__abc_22172_new_n6471_));
OR2X2 OR2X2_2478 ( .A(core__abc_22172_new_n6471_), .B(core__abc_22172_new_n5050_), .Y(core__abc_22172_new_n6472_));
OR2X2 OR2X2_2479 ( .A(core__abc_22172_new_n6403_), .B(core__abc_22172_new_n6476_), .Y(core__abc_22172_new_n6477_));
OR2X2 OR2X2_248 ( .A(_abc_19873_new_n1438_), .B(_abc_19873_new_n1429_), .Y(_abc_19873_new_n1439_));
OR2X2 OR2X2_2480 ( .A(core__abc_22172_new_n6402_), .B(core_v1_reg_17_), .Y(core__abc_22172_new_n6478_));
OR2X2 OR2X2_2481 ( .A(core__abc_22172_new_n6479_), .B(core__abc_22172_new_n5003_), .Y(core__abc_22172_new_n6480_));
OR2X2 OR2X2_2482 ( .A(core__abc_22172_new_n6481_), .B(core__abc_22172_new_n5004_), .Y(core__abc_22172_new_n6482_));
OR2X2 OR2X2_2483 ( .A(core__abc_22172_new_n6488_), .B(core__abc_22172_new_n6487_), .Y(core__abc_22172_new_n6489_));
OR2X2 OR2X2_2484 ( .A(core__abc_22172_new_n6319_), .B(core__abc_22172_new_n6496_), .Y(core__abc_22172_new_n6497_));
OR2X2 OR2X2_2485 ( .A(core__abc_22172_new_n6318_), .B(core_v1_reg_15_), .Y(core__abc_22172_new_n6498_));
OR2X2 OR2X2_2486 ( .A(core__abc_22172_new_n6501_), .B(core__abc_22172_new_n6502_), .Y(core__abc_22172_new_n6503_));
OR2X2 OR2X2_2487 ( .A(core__abc_22172_new_n6275_), .B(core_v1_reg_14_), .Y(core__abc_22172_new_n6507_));
OR2X2 OR2X2_2488 ( .A(core__abc_22172_new_n6511_), .B(core__abc_22172_new_n4842_), .Y(core__abc_22172_new_n6512_));
OR2X2 OR2X2_2489 ( .A(core__abc_22172_new_n6510_), .B(core__abc_22172_new_n6513_), .Y(core__abc_22172_new_n6514_));
OR2X2 OR2X2_249 ( .A(_abc_19873_new_n1441_), .B(_abc_19873_new_n1442_), .Y(_abc_19873_new_n1443_));
OR2X2 OR2X2_2490 ( .A(core__abc_22172_new_n6242_), .B(core__abc_22172_new_n6516_), .Y(core__abc_22172_new_n6517_));
OR2X2 OR2X2_2491 ( .A(core__abc_22172_new_n6241_), .B(core_v1_reg_13_), .Y(core__abc_22172_new_n6518_));
OR2X2 OR2X2_2492 ( .A(core__abc_22172_new_n6521_), .B(core__abc_22172_new_n6522_), .Y(core__abc_22172_new_n6523_));
OR2X2 OR2X2_2493 ( .A(core__abc_22172_new_n6529_), .B(core__abc_22172_new_n6528_), .Y(core__abc_22172_new_n6530_));
OR2X2 OR2X2_2494 ( .A(core__abc_22172_new_n6160_), .B(core__abc_22172_new_n6534_), .Y(core__abc_22172_new_n6535_));
OR2X2 OR2X2_2495 ( .A(core__abc_22172_new_n6159_), .B(core_v1_reg_11_), .Y(core__abc_22172_new_n6536_));
OR2X2 OR2X2_2496 ( .A(core__abc_22172_new_n6541_), .B(core__abc_22172_new_n6540_), .Y(core__abc_22172_new_n6542_));
OR2X2 OR2X2_2497 ( .A(core__abc_22172_new_n6548_), .B(core__abc_22172_new_n6546_), .Y(core__abc_22172_new_n6549_));
OR2X2 OR2X2_2498 ( .A(core__abc_22172_new_n6545_), .B(core__abc_22172_new_n6550_), .Y(core__abc_22172_new_n6551_));
OR2X2 OR2X2_2499 ( .A(core__abc_22172_new_n6491_), .B(core__abc_22172_new_n6501_), .Y(core__abc_22172_new_n6553_));
OR2X2 OR2X2_25 ( .A(_abc_19873_new_n966_), .B(_abc_19873_new_n967_), .Y(_abc_19873_new_n968_));
OR2X2 OR2X2_250 ( .A(_abc_19873_new_n1038_), .B(_abc_19873_new_n1444_), .Y(_abc_19873_new_n1445_));
OR2X2 OR2X2_2500 ( .A(core__abc_22172_new_n6558_), .B(core__abc_22172_new_n6556_), .Y(core__abc_22172_new_n6559_));
OR2X2 OR2X2_2501 ( .A(core__abc_22172_new_n6555_), .B(core__abc_22172_new_n6559_), .Y(core__abc_22172_new_n6560_));
OR2X2 OR2X2_2502 ( .A(core__abc_22172_new_n6560_), .B(core__abc_22172_new_n6552_), .Y(core__abc_22172_new_n6561_));
OR2X2 OR2X2_2503 ( .A(core__abc_22172_new_n6539_), .B(core__abc_22172_new_n6564_), .Y(core__abc_22172_new_n6565_));
OR2X2 OR2X2_2504 ( .A(core__abc_22172_new_n6108_), .B(core__abc_22172_new_n6570_), .Y(core__abc_22172_new_n6573_));
OR2X2 OR2X2_2505 ( .A(core__abc_22172_new_n6575_), .B(core__abc_22172_new_n4631_), .Y(core__abc_22172_new_n6576_));
OR2X2 OR2X2_2506 ( .A(core__abc_22172_new_n6574_), .B(core__abc_22172_new_n4633_), .Y(core__abc_22172_new_n6577_));
OR2X2 OR2X2_2507 ( .A(core__abc_22172_new_n6073_), .B(core__abc_22172_new_n6579_), .Y(core__abc_22172_new_n6580_));
OR2X2 OR2X2_2508 ( .A(core__abc_22172_new_n6072_), .B(core_v1_reg_9_), .Y(core__abc_22172_new_n6581_));
OR2X2 OR2X2_2509 ( .A(core__abc_22172_new_n6584_), .B(core__abc_22172_new_n6585_), .Y(core__abc_22172_new_n6586_));
OR2X2 OR2X2_251 ( .A(_abc_19873_new_n1445_), .B(_abc_19873_new_n1443_), .Y(_abc_19873_new_n1446_));
OR2X2 OR2X2_2510 ( .A(core__abc_22172_new_n6591_), .B(core__abc_22172_new_n6590_), .Y(core__abc_22172_new_n6592_));
OR2X2 OR2X2_2511 ( .A(core__abc_22172_new_n6592_), .B(core__abc_22172_new_n4533_), .Y(core__abc_22172_new_n6593_));
OR2X2 OR2X2_2512 ( .A(core__abc_22172_new_n5999_), .B(core__abc_22172_new_n6597_), .Y(core__abc_22172_new_n6598_));
OR2X2 OR2X2_2513 ( .A(core__abc_22172_new_n5998_), .B(core_v1_reg_7_), .Y(core__abc_22172_new_n6599_));
OR2X2 OR2X2_2514 ( .A(core__abc_22172_new_n6602_), .B(core__abc_22172_new_n6603_), .Y(core__abc_22172_new_n6604_));
OR2X2 OR2X2_2515 ( .A(core__abc_22172_new_n5921_), .B(core__abc_22172_new_n6608_), .Y(core__abc_22172_new_n6609_));
OR2X2 OR2X2_2516 ( .A(core__abc_22172_new_n5923_), .B(core_v1_reg_5_), .Y(core__abc_22172_new_n6610_));
OR2X2 OR2X2_2517 ( .A(core__abc_22172_new_n6613_), .B(core__abc_22172_new_n6614_), .Y(core__abc_22172_new_n6615_));
OR2X2 OR2X2_2518 ( .A(core__abc_22172_new_n6618_), .B(core__abc_22172_new_n6619_), .Y(core__abc_22172_new_n6620_));
OR2X2 OR2X2_2519 ( .A(core__abc_22172_new_n6620_), .B(core__abc_22172_new_n4409_), .Y(core__abc_22172_new_n6621_));
OR2X2 OR2X2_252 ( .A(_abc_19873_new_n1448_), .B(_abc_19873_new_n1449_), .Y(_abc_19873_new_n1450_));
OR2X2 OR2X2_2520 ( .A(core__abc_22172_new_n6622_), .B(core__abc_22172_new_n4408_), .Y(core__abc_22172_new_n6623_));
OR2X2 OR2X2_2521 ( .A(core__abc_22172_new_n5881_), .B(core__abc_22172_new_n6626_), .Y(core__abc_22172_new_n6629_));
OR2X2 OR2X2_2522 ( .A(core__abc_22172_new_n5841_), .B(core__abc_22172_new_n6633_), .Y(core__abc_22172_new_n6634_));
OR2X2 OR2X2_2523 ( .A(core__abc_22172_new_n5840_), .B(core_v1_reg_3_), .Y(core__abc_22172_new_n6635_));
OR2X2 OR2X2_2524 ( .A(core__abc_22172_new_n6641_), .B(core__abc_22172_new_n6639_), .Y(core__abc_22172_new_n6642_));
OR2X2 OR2X2_2525 ( .A(core__abc_22172_new_n6645_), .B(core__abc_22172_new_n6649_), .Y(core__abc_22172_new_n6650_));
OR2X2 OR2X2_2526 ( .A(core__abc_22172_new_n6653_), .B(core__abc_22172_new_n6594_), .Y(core__abc_22172_new_n6654_));
OR2X2 OR2X2_2527 ( .A(core__abc_22172_new_n6658_), .B(core__abc_22172_new_n6657_), .Y(core__abc_22172_new_n6659_));
OR2X2 OR2X2_2528 ( .A(core__abc_22172_new_n6656_), .B(core__abc_22172_new_n6659_), .Y(core__abc_22172_new_n6660_));
OR2X2 OR2X2_2529 ( .A(core__abc_22172_new_n6660_), .B(core__abc_22172_new_n6651_), .Y(core__abc_22172_new_n6661_));
OR2X2 OR2X2_253 ( .A(_abc_19873_new_n1450_), .B(_abc_19873_new_n1447_), .Y(_abc_19873_new_n1451_));
OR2X2 OR2X2_2530 ( .A(core__abc_22172_new_n6663_), .B(core__abc_22172_new_n6664_), .Y(core__abc_22172_new_n6665_));
OR2X2 OR2X2_2531 ( .A(core__abc_22172_new_n6665_), .B(core__abc_22172_new_n4139_), .Y(core__abc_22172_new_n6666_));
OR2X2 OR2X2_2532 ( .A(core__abc_22172_new_n6668_), .B(core__abc_22172_new_n6667_), .Y(core__abc_22172_new_n6669_));
OR2X2 OR2X2_2533 ( .A(core__abc_22172_new_n5755_), .B(core__abc_22172_new_n1286_), .Y(core__abc_22172_new_n6671_));
OR2X2 OR2X2_2534 ( .A(core__abc_22172_new_n5756_), .B(core_v1_reg_1_), .Y(core__abc_22172_new_n6672_));
OR2X2 OR2X2_2535 ( .A(core__abc_22172_new_n6675_), .B(core__abc_22172_new_n6676_), .Y(core__abc_22172_new_n6677_));
OR2X2 OR2X2_2536 ( .A(core__abc_22172_new_n6682_), .B(core__abc_22172_new_n6681_), .Y(core__abc_22172_new_n6683_));
OR2X2 OR2X2_2537 ( .A(core__abc_22172_new_n5681_), .B(core__abc_22172_new_n2343_), .Y(core__abc_22172_new_n6689_));
OR2X2 OR2X2_2538 ( .A(core__abc_22172_new_n5680_), .B(core_v1_reg_63_), .Y(core__abc_22172_new_n6690_));
OR2X2 OR2X2_2539 ( .A(core__abc_22172_new_n6700_), .B(core__abc_22172_new_n6699_), .Y(core__abc_22172_new_n6701_));
OR2X2 OR2X2_254 ( .A(_abc_19873_new_n1452_), .B(_abc_19873_new_n1453_), .Y(_abc_19873_new_n1454_));
OR2X2 OR2X2_2540 ( .A(core__abc_22172_new_n6698_), .B(core__abc_22172_new_n6701_), .Y(core__abc_22172_new_n6702_));
OR2X2 OR2X2_2541 ( .A(core__abc_22172_new_n6693_), .B(core__abc_22172_new_n6704_), .Y(core__abc_22172_new_n6705_));
OR2X2 OR2X2_2542 ( .A(core__abc_22172_new_n5634_), .B(core_v1_reg_62_), .Y(core__abc_22172_new_n6709_));
OR2X2 OR2X2_2543 ( .A(core__abc_22172_new_n6713_), .B(core__abc_22172_new_n3881_), .Y(core__abc_22172_new_n6714_));
OR2X2 OR2X2_2544 ( .A(core__abc_22172_new_n6712_), .B(core__abc_22172_new_n3880_), .Y(core__abc_22172_new_n6716_));
OR2X2 OR2X2_2545 ( .A(core__abc_22172_new_n5590_), .B(core__abc_22172_new_n6717_), .Y(core__abc_22172_new_n6718_));
OR2X2 OR2X2_2546 ( .A(core__abc_22172_new_n5589_), .B(core_v1_reg_61_), .Y(core__abc_22172_new_n6719_));
OR2X2 OR2X2_2547 ( .A(core__abc_22172_new_n6715_), .B(core__abc_22172_new_n6723_), .Y(core__abc_22172_new_n6724_));
OR2X2 OR2X2_2548 ( .A(core__abc_22172_new_n6722_), .B(core__abc_22172_new_n6726_), .Y(core__abc_22172_new_n6727_));
OR2X2 OR2X2_2549 ( .A(core__abc_22172_new_n6732_), .B(core__abc_22172_new_n6731_), .Y(core__abc_22172_new_n6733_));
OR2X2 OR2X2_255 ( .A(_abc_19873_new_n1455_), .B(_abc_19873_new_n1456_), .Y(_abc_19873_new_n1457_));
OR2X2 OR2X2_2550 ( .A(core__abc_22172_new_n6733_), .B(core__abc_22172_new_n3748_), .Y(core__abc_22172_new_n6734_));
OR2X2 OR2X2_2551 ( .A(core__abc_22172_new_n5497_), .B(core__abc_22172_new_n6738_), .Y(core__abc_22172_new_n6739_));
OR2X2 OR2X2_2552 ( .A(core__abc_22172_new_n5496_), .B(core_v1_reg_59_), .Y(core__abc_22172_new_n6740_));
OR2X2 OR2X2_2553 ( .A(core__abc_22172_new_n6744_), .B(core__abc_22172_new_n6735_), .Y(core__abc_22172_new_n6745_));
OR2X2 OR2X2_2554 ( .A(core__abc_22172_new_n6746_), .B(core__abc_22172_new_n6724_), .Y(core__abc_22172_new_n6747_));
OR2X2 OR2X2_2555 ( .A(core__abc_22172_new_n5444_), .B(core_v1_reg_58_), .Y(core__abc_22172_new_n6748_));
OR2X2 OR2X2_2556 ( .A(core__abc_22172_new_n6751_), .B(core__abc_22172_new_n3618_), .Y(core__abc_22172_new_n6753_));
OR2X2 OR2X2_2557 ( .A(core__abc_22172_new_n5400_), .B(core__abc_22172_new_n6754_), .Y(core__abc_22172_new_n6755_));
OR2X2 OR2X2_2558 ( .A(core__abc_22172_new_n5401_), .B(core_v1_reg_57_), .Y(core__abc_22172_new_n6756_));
OR2X2 OR2X2_2559 ( .A(core__abc_22172_new_n6760_), .B(core__abc_22172_new_n6752_), .Y(core__abc_22172_new_n6761_));
OR2X2 OR2X2_256 ( .A(_abc_19873_new_n1454_), .B(_abc_19873_new_n1457_), .Y(_abc_19873_new_n1458_));
OR2X2 OR2X2_2560 ( .A(core__abc_22172_new_n6759_), .B(core__abc_22172_new_n6764_), .Y(core__abc_22172_new_n6765_));
OR2X2 OR2X2_2561 ( .A(core__abc_22172_new_n6771_), .B(core__abc_22172_new_n6769_), .Y(core__abc_22172_new_n6772_));
OR2X2 OR2X2_2562 ( .A(core__abc_22172_new_n5305_), .B(core__abc_22172_new_n6777_), .Y(core__abc_22172_new_n6778_));
OR2X2 OR2X2_2563 ( .A(core__abc_22172_new_n5304_), .B(core_v1_reg_55_), .Y(core__abc_22172_new_n6779_));
OR2X2 OR2X2_2564 ( .A(core__abc_22172_new_n6786_), .B(core__abc_22172_new_n6784_), .Y(core__abc_22172_new_n6787_));
OR2X2 OR2X2_2565 ( .A(core__abc_22172_new_n6788_), .B(core__abc_22172_new_n3376_), .Y(core__abc_22172_new_n6790_));
OR2X2 OR2X2_2566 ( .A(core__abc_22172_new_n5209_), .B(core__abc_22172_new_n6791_), .Y(core__abc_22172_new_n6792_));
OR2X2 OR2X2_2567 ( .A(core__abc_22172_new_n5208_), .B(core_v1_reg_53_), .Y(core__abc_22172_new_n6793_));
OR2X2 OR2X2_2568 ( .A(core__abc_22172_new_n6794_), .B(core__abc_22172_new_n3307_), .Y(core__abc_22172_new_n6795_));
OR2X2 OR2X2_2569 ( .A(core__abc_22172_new_n5163_), .B(core__abc_22172_new_n6797_), .Y(core__abc_22172_new_n6798_));
OR2X2 OR2X2_257 ( .A(_abc_19873_new_n1458_), .B(_abc_19873_new_n1451_), .Y(_abc_19873_new_n1459_));
OR2X2 OR2X2_2570 ( .A(core__abc_22172_new_n5162_), .B(core_v1_reg_52_), .Y(core__abc_22172_new_n6799_));
OR2X2 OR2X2_2571 ( .A(core__abc_22172_new_n6800_), .B(core__abc_22172_new_n3243_), .Y(core__abc_22172_new_n6801_));
OR2X2 OR2X2_2572 ( .A(core__abc_22172_new_n1268_), .B(core_v1_reg_51_), .Y(core__abc_22172_new_n6805_));
OR2X2 OR2X2_2573 ( .A(core__abc_22172_new_n6809_), .B(core__abc_22172_new_n3244_), .Y(core__abc_22172_new_n6810_));
OR2X2 OR2X2_2574 ( .A(core__abc_22172_new_n6812_), .B(core__abc_22172_new_n6802_), .Y(core__abc_22172_new_n6813_));
OR2X2 OR2X2_2575 ( .A(core__abc_22172_new_n6814_), .B(core__abc_22172_new_n3308_), .Y(core__abc_22172_new_n6815_));
OR2X2 OR2X2_2576 ( .A(core__abc_22172_new_n6817_), .B(core__abc_22172_new_n6796_), .Y(core__abc_22172_new_n6818_));
OR2X2 OR2X2_2577 ( .A(core__abc_22172_new_n6819_), .B(core__abc_22172_new_n6789_), .Y(core__abc_22172_new_n6820_));
OR2X2 OR2X2_2578 ( .A(core__abc_22172_new_n6782_), .B(core__abc_22172_new_n6821_), .Y(core__abc_22172_new_n6822_));
OR2X2 OR2X2_2579 ( .A(core__abc_22172_new_n6824_), .B(core__abc_22172_new_n6782_), .Y(core__abc_22172_new_n6825_));
OR2X2 OR2X2_258 ( .A(_abc_19873_new_n1459_), .B(_abc_19873_new_n1446_), .Y(_abc_19873_new_n1460_));
OR2X2 OR2X2_2580 ( .A(core__abc_22172_new_n6826_), .B(core__abc_22172_new_n6774_), .Y(core__abc_22172_new_n6827_));
OR2X2 OR2X2_2581 ( .A(core__abc_22172_new_n6828_), .B(core__abc_22172_new_n6761_), .Y(core__abc_22172_new_n6829_));
OR2X2 OR2X2_2582 ( .A(core__abc_22172_new_n6743_), .B(core__abc_22172_new_n6831_), .Y(core__abc_22172_new_n6832_));
OR2X2 OR2X2_2583 ( .A(core__abc_22172_new_n6747_), .B(core__abc_22172_new_n6836_), .Y(core__abc_22172_new_n6837_));
OR2X2 OR2X2_2584 ( .A(core__abc_22172_new_n6702_), .B(core__abc_22172_new_n6838_), .Y(core__abc_22172_new_n6839_));
OR2X2 OR2X2_2585 ( .A(core__abc_22172_new_n6638_), .B(core__abc_22172_new_n6842_), .Y(core__abc_22172_new_n6843_));
OR2X2 OR2X2_2586 ( .A(core__abc_22172_new_n6661_), .B(core__abc_22172_new_n6848_), .Y(core__abc_22172_new_n6849_));
OR2X2 OR2X2_2587 ( .A(core__abc_22172_new_n6561_), .B(core__abc_22172_new_n6850_), .Y(core__abc_22172_new_n6851_));
OR2X2 OR2X2_2588 ( .A(core__abc_22172_new_n3040_), .B(core__abc_22172_new_n6852_), .Y(core__abc_22172_new_n6853_));
OR2X2 OR2X2_2589 ( .A(core__abc_22172_new_n3034_), .B(core_v1_reg_19_), .Y(core__abc_22172_new_n6854_));
OR2X2 OR2X2_259 ( .A(_abc_19873_new_n1462_), .B(_abc_19873_new_n1463_), .Y(_abc_19873_new_n1464_));
OR2X2 OR2X2_2590 ( .A(core__abc_22172_new_n6857_), .B(core__abc_22172_new_n6858_), .Y(core__abc_22172_new_n6859_));
OR2X2 OR2X2_2591 ( .A(core__abc_22172_new_n6863_), .B(core__abc_22172_new_n6861_), .Y(core__abc_22172_new_n6864_));
OR2X2 OR2X2_2592 ( .A(core__abc_22172_new_n1261_), .B(core_long), .Y(core__abc_22172_new_n6869_));
OR2X2 OR2X2_2593 ( .A(core__abc_22172_new_n6870_), .B(core_v2_reg_0_), .Y(core__abc_22172_new_n6871_));
OR2X2 OR2X2_2594 ( .A(core__abc_22172_new_n6868_), .B(core__abc_22172_new_n6873_), .Y(core__abc_22172_new_n6874_));
OR2X2 OR2X2_2595 ( .A(core__abc_22172_new_n6866_), .B(core__abc_22172_new_n6874_), .Y(core__abc_22172_new_n6875_));
OR2X2 OR2X2_2596 ( .A(core__abc_22172_new_n3205_), .B(core__abc_22172_new_n3214_), .Y(core__abc_22172_new_n6877_));
OR2X2 OR2X2_2597 ( .A(core__abc_22172_new_n6879_), .B(core__abc_22172_new_n3212_), .Y(core__abc_22172_new_n6880_));
OR2X2 OR2X2_2598 ( .A(core__abc_22172_new_n6876_), .B(core__abc_22172_new_n6881_), .Y(core__abc_22172_new_n6882_));
OR2X2 OR2X2_2599 ( .A(core__abc_22172_new_n3239_), .B(core__abc_22172_new_n6885_), .Y(core__abc_22172_new_n6888_));
OR2X2 OR2X2_26 ( .A(_abc_19873_new_n969_), .B(_abc_19873_new_n970_), .Y(_abc_19873_new_n971_));
OR2X2 OR2X2_260 ( .A(_abc_19873_new_n1192_), .B(_abc_19873_new_n1465_), .Y(_abc_19873_new_n1466_));
OR2X2 OR2X2_2600 ( .A(core__abc_22172_new_n6892_), .B(core__abc_22172_new_n6890_), .Y(core__abc_22172_new_n6893_));
OR2X2 OR2X2_2601 ( .A(core__abc_22172_new_n6896_), .B(core__abc_22172_new_n6893_), .Y(core__abc_22172_new_n6898_));
OR2X2 OR2X2_2602 ( .A(core__abc_22172_new_n6899_), .B(core__abc_22172_new_n6897_), .Y(core__abc_22172_new_n6900_));
OR2X2 OR2X2_2603 ( .A(core__abc_22172_new_n6903_), .B(core__abc_22172_new_n6904_), .Y(core__abc_22172_new_n6905_));
OR2X2 OR2X2_2604 ( .A(core__abc_22172_new_n6902_), .B(core__abc_22172_new_n6905_), .Y(core__abc_22172_new_n6906_));
OR2X2 OR2X2_2605 ( .A(core__abc_22172_new_n6907_), .B(core__abc_22172_new_n6908_), .Y(core__abc_22172_new_n6909_));
OR2X2 OR2X2_2606 ( .A(core__abc_22172_new_n6914_), .B(core__abc_22172_new_n6890_), .Y(core__abc_22172_new_n6915_));
OR2X2 OR2X2_2607 ( .A(core__abc_22172_new_n6913_), .B(core__abc_22172_new_n6915_), .Y(core__abc_22172_new_n6916_));
OR2X2 OR2X2_2608 ( .A(core__abc_22172_new_n3301_), .B(core__abc_22172_new_n6917_), .Y(core__abc_22172_new_n6918_));
OR2X2 OR2X2_2609 ( .A(core__abc_22172_new_n3302_), .B(core_v1_reg_21_), .Y(core__abc_22172_new_n6919_));
OR2X2 OR2X2_261 ( .A(_abc_19873_new_n1466_), .B(_abc_19873_new_n1464_), .Y(_abc_19873_new_n1467_));
OR2X2 OR2X2_2610 ( .A(core__abc_22172_new_n6923_), .B(core__abc_22172_new_n6921_), .Y(core__abc_22172_new_n6924_));
OR2X2 OR2X2_2611 ( .A(core__abc_22172_new_n6916_), .B(core__abc_22172_new_n6925_), .Y(core__abc_22172_new_n6928_));
OR2X2 OR2X2_2612 ( .A(core__abc_22172_new_n6931_), .B(core__abc_22172_new_n6932_), .Y(core__abc_22172_new_n6933_));
OR2X2 OR2X2_2613 ( .A(core__abc_22172_new_n6930_), .B(core__abc_22172_new_n6933_), .Y(core__abc_22172_new_n6934_));
OR2X2 OR2X2_2614 ( .A(core__abc_22172_new_n6935_), .B(core__abc_22172_new_n6936_), .Y(core__abc_22172_new_n6937_));
OR2X2 OR2X2_2615 ( .A(core__abc_22172_new_n3369_), .B(core_v1_reg_22_), .Y(core__abc_22172_new_n6941_));
OR2X2 OR2X2_2616 ( .A(core__abc_22172_new_n6947_), .B(core__abc_22172_new_n6945_), .Y(core__abc_22172_new_n6948_));
OR2X2 OR2X2_2617 ( .A(core__abc_22172_new_n6940_), .B(core__abc_22172_new_n6948_), .Y(core__abc_22172_new_n6951_));
OR2X2 OR2X2_2618 ( .A(core__abc_22172_new_n6954_), .B(core__abc_22172_new_n6955_), .Y(core__abc_22172_new_n6956_));
OR2X2 OR2X2_2619 ( .A(core__abc_22172_new_n6953_), .B(core__abc_22172_new_n6956_), .Y(core__abc_22172_new_n6957_));
OR2X2 OR2X2_262 ( .A(_abc_19873_new_n1469_), .B(_abc_19873_new_n1470_), .Y(_abc_19873_new_n1471_));
OR2X2 OR2X2_2620 ( .A(core__abc_22172_new_n6958_), .B(core__abc_22172_new_n6959_), .Y(core__abc_22172_new_n6960_));
OR2X2 OR2X2_2621 ( .A(core__abc_22172_new_n3432_), .B(core__abc_22172_new_n6962_), .Y(core__abc_22172_new_n6963_));
OR2X2 OR2X2_2622 ( .A(core__abc_22172_new_n3422_), .B(core_v1_reg_23_), .Y(core__abc_22172_new_n6964_));
OR2X2 OR2X2_2623 ( .A(core__abc_22172_new_n6968_), .B(core__abc_22172_new_n6966_), .Y(core__abc_22172_new_n6969_));
OR2X2 OR2X2_2624 ( .A(core__abc_22172_new_n6973_), .B(core__abc_22172_new_n6947_), .Y(core__abc_22172_new_n6974_));
OR2X2 OR2X2_2625 ( .A(core__abc_22172_new_n6976_), .B(core__abc_22172_new_n6977_), .Y(core__abc_22172_new_n6978_));
OR2X2 OR2X2_2626 ( .A(core__abc_22172_new_n1337_), .B(core_long), .Y(core__abc_22172_new_n6982_));
OR2X2 OR2X2_2627 ( .A(core__abc_22172_new_n6870_), .B(core_v2_reg_4_), .Y(core__abc_22172_new_n6983_));
OR2X2 OR2X2_2628 ( .A(core__abc_22172_new_n6981_), .B(core__abc_22172_new_n6985_), .Y(core__abc_22172_new_n6986_));
OR2X2 OR2X2_2629 ( .A(core__abc_22172_new_n6980_), .B(core__abc_22172_new_n6986_), .Y(core__abc_22172_new_n6987_));
OR2X2 OR2X2_263 ( .A(_abc_19873_new_n1471_), .B(_abc_19873_new_n1468_), .Y(_abc_19873_new_n1472_));
OR2X2 OR2X2_2630 ( .A(core__abc_22172_new_n6988_), .B(core__abc_22172_new_n6989_), .Y(core__abc_22172_new_n6990_));
OR2X2 OR2X2_2631 ( .A(core__abc_22172_new_n6976_), .B(core__abc_22172_new_n6968_), .Y(core__abc_22172_new_n6992_));
OR2X2 OR2X2_2632 ( .A(core__abc_22172_new_n6995_), .B(core__abc_22172_new_n6996_), .Y(core__abc_22172_new_n6997_));
OR2X2 OR2X2_2633 ( .A(core__abc_22172_new_n6997_), .B(core__abc_22172_new_n5353_), .Y(core__abc_22172_new_n7000_));
OR2X2 OR2X2_2634 ( .A(core__abc_22172_new_n6992_), .B(core__abc_22172_new_n7002_), .Y(core__abc_22172_new_n7005_));
OR2X2 OR2X2_2635 ( .A(core__abc_22172_new_n7010_), .B(core__abc_22172_new_n7011_), .Y(core__abc_22172_new_n7012_));
OR2X2 OR2X2_2636 ( .A(core__abc_22172_new_n7008_), .B(core__abc_22172_new_n7012_), .Y(core__abc_22172_new_n7013_));
OR2X2 OR2X2_2637 ( .A(core__abc_22172_new_n7014_), .B(core__abc_22172_new_n7015_), .Y(core__abc_22172_new_n7016_));
OR2X2 OR2X2_2638 ( .A(core__abc_22172_new_n3562_), .B(core__abc_22172_new_n7018_), .Y(core__abc_22172_new_n7019_));
OR2X2 OR2X2_2639 ( .A(core__abc_22172_new_n3548_), .B(core_v1_reg_25_), .Y(core__abc_22172_new_n7020_));
OR2X2 OR2X2_264 ( .A(_abc_19873_new_n1473_), .B(_abc_19873_new_n1474_), .Y(_abc_19873_new_n1475_));
OR2X2 OR2X2_2640 ( .A(core__abc_22172_new_n7024_), .B(core__abc_22172_new_n7022_), .Y(core__abc_22172_new_n7025_));
OR2X2 OR2X2_2641 ( .A(core__abc_22172_new_n7027_), .B(core__abc_22172_new_n6998_), .Y(core__abc_22172_new_n7028_));
OR2X2 OR2X2_2642 ( .A(core__abc_22172_new_n6974_), .B(core__abc_22172_new_n7030_), .Y(core__abc_22172_new_n7031_));
OR2X2 OR2X2_2643 ( .A(core__abc_22172_new_n7032_), .B(core__abc_22172_new_n7025_), .Y(core__abc_22172_new_n7033_));
OR2X2 OR2X2_2644 ( .A(core__abc_22172_new_n7034_), .B(core__abc_22172_new_n7035_), .Y(core__abc_22172_new_n7036_));
OR2X2 OR2X2_2645 ( .A(core__abc_22172_new_n7040_), .B(core__abc_22172_new_n7041_), .Y(core__abc_22172_new_n7042_));
OR2X2 OR2X2_2646 ( .A(core__abc_22172_new_n7038_), .B(core__abc_22172_new_n7042_), .Y(core__abc_22172_new_n7043_));
OR2X2 OR2X2_2647 ( .A(core__abc_22172_new_n7044_), .B(core__abc_22172_new_n7045_), .Y(core__abc_22172_new_n7046_));
OR2X2 OR2X2_2648 ( .A(core__abc_22172_new_n7053_), .B(core__abc_22172_new_n7052_), .Y(core__abc_22172_new_n7054_));
OR2X2 OR2X2_2649 ( .A(core__abc_22172_new_n7056_), .B(core__abc_22172_new_n7057_), .Y(core__abc_22172_new_n7058_));
OR2X2 OR2X2_265 ( .A(_abc_19873_new_n1476_), .B(_abc_19873_new_n1477_), .Y(_abc_19873_new_n1478_));
OR2X2 OR2X2_2650 ( .A(core__abc_22172_new_n7049_), .B(core__abc_22172_new_n7058_), .Y(core__abc_22172_new_n7061_));
OR2X2 OR2X2_2651 ( .A(core__abc_22172_new_n7064_), .B(core__abc_22172_new_n7065_), .Y(core__abc_22172_new_n7066_));
OR2X2 OR2X2_2652 ( .A(core__abc_22172_new_n7063_), .B(core__abc_22172_new_n7066_), .Y(core__abc_22172_new_n7067_));
OR2X2 OR2X2_2653 ( .A(core__abc_22172_new_n7068_), .B(core__abc_22172_new_n7069_), .Y(core__abc_22172_new_n7070_));
OR2X2 OR2X2_2654 ( .A(core__abc_22172_new_n6948_), .B(core__abc_22172_new_n6924_), .Y(core__abc_22172_new_n7072_));
OR2X2 OR2X2_2655 ( .A(core__abc_22172_new_n7058_), .B(core__abc_22172_new_n7025_), .Y(core__abc_22172_new_n7075_));
OR2X2 OR2X2_2656 ( .A(core__abc_22172_new_n7075_), .B(core__abc_22172_new_n7030_), .Y(core__abc_22172_new_n7076_));
OR2X2 OR2X2_2657 ( .A(core__abc_22172_new_n6972_), .B(core__abc_22172_new_n6947_), .Y(core__abc_22172_new_n7080_));
OR2X2 OR2X2_2658 ( .A(core__abc_22172_new_n7083_), .B(core__abc_22172_new_n7076_), .Y(core__abc_22172_new_n7084_));
OR2X2 OR2X2_2659 ( .A(core__abc_22172_new_n7056_), .B(core__abc_22172_new_n7024_), .Y(core__abc_22172_new_n7086_));
OR2X2 OR2X2_266 ( .A(_abc_19873_new_n1475_), .B(_abc_19873_new_n1478_), .Y(_abc_19873_new_n1479_));
OR2X2 OR2X2_2660 ( .A(core__abc_22172_new_n7075_), .B(core__abc_22172_new_n7028_), .Y(core__abc_22172_new_n7089_));
OR2X2 OR2X2_2661 ( .A(core__abc_22172_new_n7079_), .B(core__abc_22172_new_n7092_), .Y(core__abc_22172_new_n7093_));
OR2X2 OR2X2_2662 ( .A(core__abc_22172_new_n3688_), .B(core__abc_22172_new_n7094_), .Y(core__abc_22172_new_n7095_));
OR2X2 OR2X2_2663 ( .A(core__abc_22172_new_n3687_), .B(core_v1_reg_27_), .Y(core__abc_22172_new_n7096_));
OR2X2 OR2X2_2664 ( .A(core__abc_22172_new_n7100_), .B(core__abc_22172_new_n7098_), .Y(core__abc_22172_new_n7101_));
OR2X2 OR2X2_2665 ( .A(core__abc_22172_new_n7105_), .B(core__abc_22172_new_n7103_), .Y(core__abc_22172_new_n7106_));
OR2X2 OR2X2_2666 ( .A(core__abc_22172_new_n7109_), .B(core__abc_22172_new_n7110_), .Y(core__abc_22172_new_n7111_));
OR2X2 OR2X2_2667 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n7111_), .Y(core__abc_22172_new_n7112_));
OR2X2 OR2X2_2668 ( .A(core__abc_22172_new_n7108_), .B(core__abc_22172_new_n7112_), .Y(core__abc_22172_new_n7113_));
OR2X2 OR2X2_2669 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_8_), .Y(core__abc_22172_new_n7115_));
OR2X2 OR2X2_267 ( .A(_abc_19873_new_n1479_), .B(_abc_19873_new_n1472_), .Y(_abc_19873_new_n1480_));
OR2X2 OR2X2_2670 ( .A(core__abc_22172_new_n7120_), .B(core__abc_22172_new_n7121_), .Y(core__abc_22172_new_n7122_));
OR2X2 OR2X2_2671 ( .A(core__abc_22172_new_n7122_), .B(core__abc_22172_new_n5552_), .Y(core__abc_22172_new_n7123_));
OR2X2 OR2X2_2672 ( .A(core__abc_22172_new_n7130_), .B(core__abc_22172_new_n7127_), .Y(core__abc_22172_new_n7132_));
OR2X2 OR2X2_2673 ( .A(core__abc_22172_new_n7133_), .B(core__abc_22172_new_n7131_), .Y(core__abc_22172_new_n7134_));
OR2X2 OR2X2_2674 ( .A(core__abc_22172_new_n7138_), .B(core__abc_22172_new_n7139_), .Y(core__abc_22172_new_n7140_));
OR2X2 OR2X2_2675 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n7140_), .Y(core__abc_22172_new_n7141_));
OR2X2 OR2X2_2676 ( .A(core__abc_22172_new_n7136_), .B(core__abc_22172_new_n7141_), .Y(core__abc_22172_new_n7142_));
OR2X2 OR2X2_2677 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_9_), .Y(core__abc_22172_new_n7143_));
OR2X2 OR2X2_2678 ( .A(core__abc_22172_new_n7124_), .B(core__abc_22172_new_n7128_), .Y(core__abc_22172_new_n7148_));
OR2X2 OR2X2_2679 ( .A(core__abc_22172_new_n7147_), .B(core__abc_22172_new_n7150_), .Y(core__abc_22172_new_n7151_));
OR2X2 OR2X2_268 ( .A(_abc_19873_new_n1480_), .B(_abc_19873_new_n1467_), .Y(_abc_19873_new_n1481_));
OR2X2 OR2X2_2680 ( .A(core__abc_22172_new_n3832_), .B(core__abc_22172_new_n7152_), .Y(core__abc_22172_new_n7153_));
OR2X2 OR2X2_2681 ( .A(core__abc_22172_new_n3818_), .B(core_v1_reg_29_), .Y(core__abc_22172_new_n7154_));
OR2X2 OR2X2_2682 ( .A(core__abc_22172_new_n7157_), .B(core__abc_22172_new_n7158_), .Y(core__abc_22172_new_n7159_));
OR2X2 OR2X2_2683 ( .A(core__abc_22172_new_n7151_), .B(core__abc_22172_new_n7160_), .Y(core__abc_22172_new_n7163_));
OR2X2 OR2X2_2684 ( .A(core__abc_22172_new_n7166_), .B(core__abc_22172_new_n7167_), .Y(core__abc_22172_new_n7168_));
OR2X2 OR2X2_2685 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n7168_), .Y(core__abc_22172_new_n7169_));
OR2X2 OR2X2_2686 ( .A(core__abc_22172_new_n7165_), .B(core__abc_22172_new_n7169_), .Y(core__abc_22172_new_n7170_));
OR2X2 OR2X2_2687 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_10_), .Y(core__abc_22172_new_n7171_));
OR2X2 OR2X2_2688 ( .A(core__abc_22172_new_n7178_), .B(core__abc_22172_new_n7177_), .Y(core__abc_22172_new_n7179_));
OR2X2 OR2X2_2689 ( .A(core__abc_22172_new_n7179_), .B(core__abc_22172_new_n3189_), .Y(core__abc_22172_new_n7180_));
OR2X2 OR2X2_269 ( .A(_abc_19873_new_n1483_), .B(_abc_19873_new_n1484_), .Y(_abc_19873_new_n1485_));
OR2X2 OR2X2_2690 ( .A(core__abc_22172_new_n7175_), .B(core__abc_22172_new_n7184_), .Y(core__abc_22172_new_n7187_));
OR2X2 OR2X2_2691 ( .A(core__abc_22172_new_n7190_), .B(core__abc_22172_new_n7191_), .Y(core__abc_22172_new_n7192_));
OR2X2 OR2X2_2692 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n7192_), .Y(core__abc_22172_new_n7193_));
OR2X2 OR2X2_2693 ( .A(core__abc_22172_new_n7189_), .B(core__abc_22172_new_n7193_), .Y(core__abc_22172_new_n7194_));
OR2X2 OR2X2_2694 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_11_), .Y(core__abc_22172_new_n7195_));
OR2X2 OR2X2_2695 ( .A(core__abc_22172_new_n7201_), .B(core__abc_22172_new_n7200_), .Y(core__abc_22172_new_n7202_));
OR2X2 OR2X2_2696 ( .A(core__abc_22172_new_n7199_), .B(core__abc_22172_new_n7202_), .Y(core__abc_22172_new_n7203_));
OR2X2 OR2X2_2697 ( .A(core__abc_22172_new_n7205_), .B(core__abc_22172_new_n7203_), .Y(core__abc_22172_new_n7206_));
OR2X2 OR2X2_2698 ( .A(core__abc_22172_new_n3959_), .B(core__abc_22172_new_n7207_), .Y(core__abc_22172_new_n7208_));
OR2X2 OR2X2_2699 ( .A(core__abc_22172_new_n3946_), .B(core_v1_reg_31_), .Y(core__abc_22172_new_n7209_));
OR2X2 OR2X2_27 ( .A(_abc_19873_new_n968_), .B(_abc_19873_new_n971_), .Y(_abc_19873_new_n972_));
OR2X2 OR2X2_270 ( .A(_abc_19873_new_n1487_), .B(_abc_19873_new_n1488_), .Y(_abc_19873_new_n1489_));
OR2X2 OR2X2_2700 ( .A(core__abc_22172_new_n7212_), .B(core__abc_22172_new_n7213_), .Y(core__abc_22172_new_n7214_));
OR2X2 OR2X2_2701 ( .A(core__abc_22172_new_n7218_), .B(core__abc_22172_new_n7216_), .Y(core__abc_22172_new_n7219_));
OR2X2 OR2X2_2702 ( .A(core__abc_22172_new_n7223_), .B(core__abc_22172_new_n7224_), .Y(core__abc_22172_new_n7225_));
OR2X2 OR2X2_2703 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n7225_), .Y(core__abc_22172_new_n7226_));
OR2X2 OR2X2_2704 ( .A(core__abc_22172_new_n7221_), .B(core__abc_22172_new_n7226_), .Y(core__abc_22172_new_n7227_));
OR2X2 OR2X2_2705 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_12_), .Y(core__abc_22172_new_n7228_));
OR2X2 OR2X2_2706 ( .A(core__abc_22172_new_n7216_), .B(core__abc_22172_new_n7212_), .Y(core__abc_22172_new_n7231_));
OR2X2 OR2X2_2707 ( .A(core__abc_22172_new_n7235_), .B(core__abc_22172_new_n7234_), .Y(core__abc_22172_new_n7236_));
OR2X2 OR2X2_2708 ( .A(core__abc_22172_new_n7238_), .B(core__abc_22172_new_n7239_), .Y(core__abc_22172_new_n7240_));
OR2X2 OR2X2_2709 ( .A(core__abc_22172_new_n7244_), .B(core__abc_22172_new_n7241_), .Y(core__abc_22172_new_n7245_));
OR2X2 OR2X2_271 ( .A(_abc_19873_new_n1489_), .B(_abc_19873_new_n1486_), .Y(_abc_19873_new_n1490_));
OR2X2 OR2X2_2710 ( .A(core__abc_22172_new_n7248_), .B(core__abc_22172_new_n7249_), .Y(core__abc_22172_new_n7250_));
OR2X2 OR2X2_2711 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n7250_), .Y(core__abc_22172_new_n7251_));
OR2X2 OR2X2_2712 ( .A(core__abc_22172_new_n7246_), .B(core__abc_22172_new_n7251_), .Y(core__abc_22172_new_n7252_));
OR2X2 OR2X2_2713 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_13_), .Y(core__abc_22172_new_n7253_));
OR2X2 OR2X2_2714 ( .A(core__abc_22172_new_n7238_), .B(core__abc_22172_new_n7212_), .Y(core__abc_22172_new_n7257_));
OR2X2 OR2X2_2715 ( .A(core__abc_22172_new_n7217_), .B(core__abc_22172_new_n7261_), .Y(core__abc_22172_new_n7262_));
OR2X2 OR2X2_2716 ( .A(core__abc_22172_new_n7266_), .B(core__abc_22172_new_n7265_), .Y(core__abc_22172_new_n7267_));
OR2X2 OR2X2_2717 ( .A(core__abc_22172_new_n4078_), .B(core_v1_reg_33_), .Y(core__abc_22172_new_n7268_));
OR2X2 OR2X2_2718 ( .A(core__abc_22172_new_n7272_), .B(core__abc_22172_new_n7270_), .Y(core__abc_22172_new_n7273_));
OR2X2 OR2X2_2719 ( .A(core__abc_22172_new_n7275_), .B(core__abc_22172_new_n7276_), .Y(core__abc_22172_new_n7277_));
OR2X2 OR2X2_272 ( .A(_abc_19873_new_n1490_), .B(_abc_19873_new_n1485_), .Y(_abc_19873_new_n1491_));
OR2X2 OR2X2_2720 ( .A(core__abc_22172_new_n7281_), .B(core__abc_22172_new_n7282_), .Y(core__abc_22172_new_n7283_));
OR2X2 OR2X2_2721 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n7283_), .Y(core__abc_22172_new_n7284_));
OR2X2 OR2X2_2722 ( .A(core__abc_22172_new_n7279_), .B(core__abc_22172_new_n7284_), .Y(core__abc_22172_new_n7285_));
OR2X2 OR2X2_2723 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_14_), .Y(core__abc_22172_new_n7286_));
OR2X2 OR2X2_2724 ( .A(core__abc_22172_new_n7275_), .B(core__abc_22172_new_n7272_), .Y(core__abc_22172_new_n7289_));
OR2X2 OR2X2_2725 ( .A(core__abc_22172_new_n4134_), .B(core_v1_reg_34_), .Y(core__abc_22172_new_n7291_));
OR2X2 OR2X2_2726 ( .A(core__abc_22172_new_n7296_), .B(core__abc_22172_new_n7292_), .Y(core__abc_22172_new_n7297_));
OR2X2 OR2X2_2727 ( .A(core__abc_22172_new_n7298_), .B(core__abc_22172_new_n7295_), .Y(core__abc_22172_new_n7299_));
OR2X2 OR2X2_2728 ( .A(core__abc_22172_new_n7297_), .B(core__abc_22172_new_n3447_), .Y(core__abc_22172_new_n7301_));
OR2X2 OR2X2_2729 ( .A(core__abc_22172_new_n7294_), .B(core__abc_22172_new_n3450_), .Y(core__abc_22172_new_n7302_));
OR2X2 OR2X2_273 ( .A(_abc_19873_new_n1493_), .B(_abc_19873_new_n1494_), .Y(_abc_19873_new_n1495_));
OR2X2 OR2X2_2730 ( .A(core__abc_22172_new_n7300_), .B(core__abc_22172_new_n7304_), .Y(core__abc_22172_new_n7305_));
OR2X2 OR2X2_2731 ( .A(core__abc_22172_new_n7308_), .B(core__abc_22172_new_n7309_), .Y(core__abc_22172_new_n7310_));
OR2X2 OR2X2_2732 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n7310_), .Y(core__abc_22172_new_n7311_));
OR2X2 OR2X2_2733 ( .A(core__abc_22172_new_n7307_), .B(core__abc_22172_new_n7311_), .Y(core__abc_22172_new_n7312_));
OR2X2 OR2X2_2734 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_15_), .Y(core__abc_22172_new_n7313_));
OR2X2 OR2X2_2735 ( .A(core__abc_22172_new_n7299_), .B(core__abc_22172_new_n7273_), .Y(core__abc_22172_new_n7317_));
OR2X2 OR2X2_2736 ( .A(core__abc_22172_new_n7317_), .B(core__abc_22172_new_n7261_), .Y(core__abc_22172_new_n7318_));
OR2X2 OR2X2_2737 ( .A(core__abc_22172_new_n7318_), .B(core__abc_22172_new_n7316_), .Y(core__abc_22172_new_n7319_));
OR2X2 OR2X2_2738 ( .A(core__abc_22172_new_n7317_), .B(core__abc_22172_new_n7259_), .Y(core__abc_22172_new_n7320_));
OR2X2 OR2X2_2739 ( .A(core__abc_22172_new_n7321_), .B(core__abc_22172_new_n7295_), .Y(core__abc_22172_new_n7322_));
OR2X2 OR2X2_274 ( .A(_abc_19873_new_n1496_), .B(_abc_19873_new_n1497_), .Y(_abc_19873_new_n1498_));
OR2X2 OR2X2_2740 ( .A(core__abc_22172_new_n7318_), .B(core__abc_22172_new_n7326_), .Y(core__abc_22172_new_n7327_));
OR2X2 OR2X2_2741 ( .A(core__abc_22172_new_n7327_), .B(core__abc_22172_new_n7091_), .Y(core__abc_22172_new_n7328_));
OR2X2 OR2X2_2742 ( .A(core__abc_22172_new_n4231_), .B(core__abc_22172_new_n7338_), .Y(core__abc_22172_new_n7339_));
OR2X2 OR2X2_2743 ( .A(core__abc_22172_new_n4220_), .B(core_v1_reg_35_), .Y(core__abc_22172_new_n7340_));
OR2X2 OR2X2_2744 ( .A(core__abc_22172_new_n7343_), .B(core__abc_22172_new_n7344_), .Y(core__abc_22172_new_n7345_));
OR2X2 OR2X2_2745 ( .A(core__abc_22172_new_n7347_), .B(core__abc_22172_new_n7348_), .Y(core__abc_22172_new_n7349_));
OR2X2 OR2X2_2746 ( .A(core__abc_22172_new_n7353_), .B(core__abc_22172_new_n7354_), .Y(core__abc_22172_new_n7355_));
OR2X2 OR2X2_2747 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n7355_), .Y(core__abc_22172_new_n7356_));
OR2X2 OR2X2_2748 ( .A(core__abc_22172_new_n7351_), .B(core__abc_22172_new_n7356_), .Y(core__abc_22172_new_n7357_));
OR2X2 OR2X2_2749 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_16_), .Y(core__abc_22172_new_n7358_));
OR2X2 OR2X2_275 ( .A(_abc_19873_new_n1495_), .B(_abc_19873_new_n1498_), .Y(_abc_19873_new_n1499_));
OR2X2 OR2X2_2750 ( .A(core__abc_22172_new_n7366_), .B(core__abc_22172_new_n7367_), .Y(core__abc_22172_new_n7368_));
OR2X2 OR2X2_2751 ( .A(core__abc_22172_new_n7363_), .B(core__abc_22172_new_n7374_), .Y(core__abc_22172_new_n7375_));
OR2X2 OR2X2_2752 ( .A(core__abc_22172_new_n7376_), .B(core__abc_22172_new_n7377_), .Y(core__abc_22172_new_n7378_));
OR2X2 OR2X2_2753 ( .A(core__abc_22172_new_n7382_), .B(core__abc_22172_new_n7383_), .Y(core__abc_22172_new_n7384_));
OR2X2 OR2X2_2754 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n7384_), .Y(core__abc_22172_new_n7385_));
OR2X2 OR2X2_2755 ( .A(core__abc_22172_new_n7381_), .B(core__abc_22172_new_n7385_), .Y(core__abc_22172_new_n7386_));
OR2X2 OR2X2_2756 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_17_), .Y(core__abc_22172_new_n7387_));
OR2X2 OR2X2_2757 ( .A(core__abc_22172_new_n4347_), .B(core__abc_22172_new_n7390_), .Y(core__abc_22172_new_n7391_));
OR2X2 OR2X2_2758 ( .A(core__abc_22172_new_n4360_), .B(core_v1_reg_37_), .Y(core__abc_22172_new_n7392_));
OR2X2 OR2X2_2759 ( .A(core__abc_22172_new_n7395_), .B(core__abc_22172_new_n7396_), .Y(core__abc_22172_new_n7397_));
OR2X2 OR2X2_276 ( .A(_abc_19873_new_n1499_), .B(_abc_19873_new_n1492_), .Y(_abc_19873_new_n1500_));
OR2X2 OR2X2_2760 ( .A(core__abc_22172_new_n7400_), .B(core__abc_22172_new_n7372_), .Y(core__abc_22172_new_n7401_));
OR2X2 OR2X2_2761 ( .A(core__abc_22172_new_n7403_), .B(core__abc_22172_new_n7404_), .Y(core__abc_22172_new_n7405_));
OR2X2 OR2X2_2762 ( .A(core__abc_22172_new_n7409_), .B(core__abc_22172_new_n7410_), .Y(core__abc_22172_new_n7411_));
OR2X2 OR2X2_2763 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n7411_), .Y(core__abc_22172_new_n7412_));
OR2X2 OR2X2_2764 ( .A(core__abc_22172_new_n7407_), .B(core__abc_22172_new_n7412_), .Y(core__abc_22172_new_n7413_));
OR2X2 OR2X2_2765 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_18_), .Y(core__abc_22172_new_n7414_));
OR2X2 OR2X2_2766 ( .A(core__abc_22172_new_n7403_), .B(core__abc_22172_new_n7395_), .Y(core__abc_22172_new_n7417_));
OR2X2 OR2X2_2767 ( .A(core__abc_22172_new_n7420_), .B(core__abc_22172_new_n7421_), .Y(core__abc_22172_new_n7422_));
OR2X2 OR2X2_2768 ( .A(core__abc_22172_new_n7417_), .B(core__abc_22172_new_n7428_), .Y(core__abc_22172_new_n7429_));
OR2X2 OR2X2_2769 ( .A(core__abc_22172_new_n7430_), .B(core__abc_22172_new_n7431_), .Y(core__abc_22172_new_n7432_));
OR2X2 OR2X2_277 ( .A(_abc_19873_new_n1500_), .B(_abc_19873_new_n1491_), .Y(_abc_19873_new_n1501_));
OR2X2 OR2X2_2770 ( .A(core__abc_22172_new_n7435_), .B(core__abc_22172_new_n7436_), .Y(core__abc_22172_new_n7437_));
OR2X2 OR2X2_2771 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n7437_), .Y(core__abc_22172_new_n7438_));
OR2X2 OR2X2_2772 ( .A(core__abc_22172_new_n7434_), .B(core__abc_22172_new_n7438_), .Y(core__abc_22172_new_n7439_));
OR2X2 OR2X2_2773 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_19_), .Y(core__abc_22172_new_n7440_));
OR2X2 OR2X2_2774 ( .A(core__abc_22172_new_n7424_), .B(core__abc_22172_new_n7395_), .Y(core__abc_22172_new_n7443_));
OR2X2 OR2X2_2775 ( .A(core__abc_22172_new_n7399_), .B(core__abc_22172_new_n7372_), .Y(core__abc_22172_new_n7446_));
OR2X2 OR2X2_2776 ( .A(core__abc_22172_new_n7448_), .B(core__abc_22172_new_n7446_), .Y(core__abc_22172_new_n7449_));
OR2X2 OR2X2_2777 ( .A(core__abc_22172_new_n7336_), .B(core__abc_22172_new_n7453_), .Y(core__abc_22172_new_n7454_));
OR2X2 OR2X2_2778 ( .A(core__abc_22172_new_n4473_), .B(core__abc_22172_new_n7456_), .Y(core__abc_22172_new_n7457_));
OR2X2 OR2X2_2779 ( .A(core__abc_22172_new_n4472_), .B(core_v1_reg_39_), .Y(core__abc_22172_new_n7458_));
OR2X2 OR2X2_278 ( .A(_abc_19873_new_n1503_), .B(_abc_19873_new_n1504_), .Y(_abc_19873_new_n1505_));
OR2X2 OR2X2_2780 ( .A(core__abc_22172_new_n7461_), .B(core__abc_22172_new_n7462_), .Y(core__abc_22172_new_n7463_));
OR2X2 OR2X2_2781 ( .A(core__abc_22172_new_n7455_), .B(core__abc_22172_new_n7463_), .Y(core__abc_22172_new_n7464_));
OR2X2 OR2X2_2782 ( .A(core__abc_22172_new_n7465_), .B(core__abc_22172_new_n7466_), .Y(core__abc_22172_new_n7467_));
OR2X2 OR2X2_2783 ( .A(core__abc_22172_new_n7470_), .B(core__abc_22172_new_n7471_), .Y(core__abc_22172_new_n7472_));
OR2X2 OR2X2_2784 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n7472_), .Y(core__abc_22172_new_n7473_));
OR2X2 OR2X2_2785 ( .A(core__abc_22172_new_n7469_), .B(core__abc_22172_new_n7473_), .Y(core__abc_22172_new_n7474_));
OR2X2 OR2X2_2786 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_20_), .Y(core__abc_22172_new_n7475_));
OR2X2 OR2X2_2787 ( .A(core__abc_22172_new_n7484_), .B(core__abc_22172_new_n7483_), .Y(core__abc_22172_new_n7485_));
OR2X2 OR2X2_2788 ( .A(core__abc_22172_new_n7480_), .B(core__abc_22172_new_n7491_), .Y(core__abc_22172_new_n7492_));
OR2X2 OR2X2_2789 ( .A(core__abc_22172_new_n7479_), .B(core__abc_22172_new_n7493_), .Y(core__abc_22172_new_n7494_));
OR2X2 OR2X2_279 ( .A(_abc_19873_new_n1507_), .B(_abc_19873_new_n1508_), .Y(_abc_19873_new_n1509_));
OR2X2 OR2X2_2790 ( .A(core__abc_22172_new_n7498_), .B(core__abc_22172_new_n7499_), .Y(core__abc_22172_new_n7500_));
OR2X2 OR2X2_2791 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n7500_), .Y(core__abc_22172_new_n7501_));
OR2X2 OR2X2_2792 ( .A(core__abc_22172_new_n7496_), .B(core__abc_22172_new_n7501_), .Y(core__abc_22172_new_n7502_));
OR2X2 OR2X2_2793 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_21_), .Y(core__abc_22172_new_n7503_));
OR2X2 OR2X2_2794 ( .A(core__abc_22172_new_n7507_), .B(core__abc_22172_new_n7506_), .Y(core__abc_22172_new_n7508_));
OR2X2 OR2X2_2795 ( .A(core__abc_22172_new_n4583_), .B(core_v1_reg_41_), .Y(core__abc_22172_new_n7509_));
OR2X2 OR2X2_2796 ( .A(core__abc_22172_new_n7512_), .B(core__abc_22172_new_n7513_), .Y(core__abc_22172_new_n7514_));
OR2X2 OR2X2_2797 ( .A(core__abc_22172_new_n7493_), .B(core__abc_22172_new_n7463_), .Y(core__abc_22172_new_n7515_));
OR2X2 OR2X2_2798 ( .A(core__abc_22172_new_n7455_), .B(core__abc_22172_new_n7515_), .Y(core__abc_22172_new_n7516_));
OR2X2 OR2X2_2799 ( .A(core__abc_22172_new_n7517_), .B(core__abc_22172_new_n7489_), .Y(core__abc_22172_new_n7518_));
OR2X2 OR2X2_28 ( .A(_abc_19873_new_n972_), .B(_abc_19873_new_n965_), .Y(_abc_19873_new_n973_));
OR2X2 OR2X2_280 ( .A(_abc_19873_new_n1509_), .B(_abc_19873_new_n1506_), .Y(_abc_19873_new_n1510_));
OR2X2 OR2X2_2800 ( .A(core__abc_22172_new_n7519_), .B(core__abc_22172_new_n7514_), .Y(core__abc_22172_new_n7520_));
OR2X2 OR2X2_2801 ( .A(core__abc_22172_new_n7521_), .B(core__abc_22172_new_n7522_), .Y(core__abc_22172_new_n7523_));
OR2X2 OR2X2_2802 ( .A(core__abc_22172_new_n7527_), .B(core__abc_22172_new_n7528_), .Y(core__abc_22172_new_n7529_));
OR2X2 OR2X2_2803 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n7529_), .Y(core__abc_22172_new_n7530_));
OR2X2 OR2X2_2804 ( .A(core__abc_22172_new_n7525_), .B(core__abc_22172_new_n7530_), .Y(core__abc_22172_new_n7531_));
OR2X2 OR2X2_2805 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_22_), .Y(core__abc_22172_new_n7532_));
OR2X2 OR2X2_2806 ( .A(core__abc_22172_new_n7539_), .B(core__abc_22172_new_n7540_), .Y(core__abc_22172_new_n7541_));
OR2X2 OR2X2_2807 ( .A(core__abc_22172_new_n7551_), .B(core__abc_22172_new_n7549_), .Y(core__abc_22172_new_n7552_));
OR2X2 OR2X2_2808 ( .A(core__abc_22172_new_n7555_), .B(core__abc_22172_new_n7556_), .Y(core__abc_22172_new_n7557_));
OR2X2 OR2X2_2809 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n7557_), .Y(core__abc_22172_new_n7558_));
OR2X2 OR2X2_281 ( .A(_abc_19873_new_n1510_), .B(_abc_19873_new_n1505_), .Y(_abc_19873_new_n1511_));
OR2X2 OR2X2_2810 ( .A(core__abc_22172_new_n7554_), .B(core__abc_22172_new_n7558_), .Y(core__abc_22172_new_n7559_));
OR2X2 OR2X2_2811 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_23_), .Y(core__abc_22172_new_n7560_));
OR2X2 OR2X2_2812 ( .A(core__abc_22172_new_n7571_), .B(core__abc_22172_new_n7543_), .Y(core__abc_22172_new_n7572_));
OR2X2 OR2X2_2813 ( .A(core__abc_22172_new_n7570_), .B(core__abc_22172_new_n7572_), .Y(core__abc_22172_new_n7573_));
OR2X2 OR2X2_2814 ( .A(core__abc_22172_new_n7573_), .B(core__abc_22172_new_n7568_), .Y(core__abc_22172_new_n7574_));
OR2X2 OR2X2_2815 ( .A(core__abc_22172_new_n7576_), .B(core__abc_22172_new_n7574_), .Y(core__abc_22172_new_n7577_));
OR2X2 OR2X2_2816 ( .A(core__abc_22172_new_n4708_), .B(core__abc_22172_new_n7578_), .Y(core__abc_22172_new_n7579_));
OR2X2 OR2X2_2817 ( .A(core__abc_22172_new_n4694_), .B(core_v1_reg_43_), .Y(core__abc_22172_new_n7580_));
OR2X2 OR2X2_2818 ( .A(core__abc_22172_new_n7583_), .B(core__abc_22172_new_n7584_), .Y(core__abc_22172_new_n7585_));
OR2X2 OR2X2_2819 ( .A(core__abc_22172_new_n7589_), .B(core__abc_22172_new_n7587_), .Y(core__abc_22172_new_n7590_));
OR2X2 OR2X2_282 ( .A(_abc_19873_new_n1513_), .B(_abc_19873_new_n1514_), .Y(_abc_19873_new_n1515_));
OR2X2 OR2X2_2820 ( .A(core__abc_22172_new_n7593_), .B(core__abc_22172_new_n7594_), .Y(core__abc_22172_new_n7595_));
OR2X2 OR2X2_2821 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n7595_), .Y(core__abc_22172_new_n7596_));
OR2X2 OR2X2_2822 ( .A(core__abc_22172_new_n7592_), .B(core__abc_22172_new_n7596_), .Y(core__abc_22172_new_n7597_));
OR2X2 OR2X2_2823 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_24_), .Y(core__abc_22172_new_n7598_));
OR2X2 OR2X2_2824 ( .A(core__abc_22172_new_n7587_), .B(core__abc_22172_new_n7583_), .Y(core__abc_22172_new_n7601_));
OR2X2 OR2X2_2825 ( .A(core__abc_22172_new_n4749_), .B(core_v1_reg_44_), .Y(core__abc_22172_new_n7604_));
OR2X2 OR2X2_2826 ( .A(core__abc_22172_new_n7601_), .B(core__abc_22172_new_n7611_), .Y(core__abc_22172_new_n7612_));
OR2X2 OR2X2_2827 ( .A(core__abc_22172_new_n7613_), .B(core__abc_22172_new_n7614_), .Y(core__abc_22172_new_n7615_));
OR2X2 OR2X2_2828 ( .A(core__abc_22172_new_n7619_), .B(core__abc_22172_new_n7620_), .Y(core__abc_22172_new_n7621_));
OR2X2 OR2X2_2829 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n7621_), .Y(core__abc_22172_new_n7622_));
OR2X2 OR2X2_283 ( .A(_abc_19873_new_n1516_), .B(_abc_19873_new_n1517_), .Y(_abc_19873_new_n1518_));
OR2X2 OR2X2_2830 ( .A(core__abc_22172_new_n7617_), .B(core__abc_22172_new_n7622_), .Y(core__abc_22172_new_n7623_));
OR2X2 OR2X2_2831 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_25_), .Y(core__abc_22172_new_n7624_));
OR2X2 OR2X2_2832 ( .A(core__abc_22172_new_n4793_), .B(core__abc_22172_new_n7627_), .Y(core__abc_22172_new_n7628_));
OR2X2 OR2X2_2833 ( .A(core__abc_22172_new_n4792_), .B(core_v1_reg_45_), .Y(core__abc_22172_new_n7629_));
OR2X2 OR2X2_2834 ( .A(core__abc_22172_new_n7632_), .B(core__abc_22172_new_n7633_), .Y(core__abc_22172_new_n7634_));
OR2X2 OR2X2_2835 ( .A(core__abc_22172_new_n7639_), .B(core__abc_22172_new_n7609_), .Y(core__abc_22172_new_n7640_));
OR2X2 OR2X2_2836 ( .A(core__abc_22172_new_n7637_), .B(core__abc_22172_new_n7641_), .Y(core__abc_22172_new_n7642_));
OR2X2 OR2X2_2837 ( .A(core__abc_22172_new_n7642_), .B(core__abc_22172_new_n7635_), .Y(core__abc_22172_new_n7645_));
OR2X2 OR2X2_2838 ( .A(core__abc_22172_new_n7649_), .B(core__abc_22172_new_n7650_), .Y(core__abc_22172_new_n7651_));
OR2X2 OR2X2_2839 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n7651_), .Y(core__abc_22172_new_n7652_));
OR2X2 OR2X2_284 ( .A(_abc_19873_new_n1515_), .B(_abc_19873_new_n1518_), .Y(_abc_19873_new_n1519_));
OR2X2 OR2X2_2840 ( .A(core__abc_22172_new_n7647_), .B(core__abc_22172_new_n7652_), .Y(core__abc_22172_new_n7653_));
OR2X2 OR2X2_2841 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_26_), .Y(core__abc_22172_new_n7654_));
OR2X2 OR2X2_2842 ( .A(core__abc_22172_new_n7662_), .B(core__abc_22172_new_n7661_), .Y(core__abc_22172_new_n7663_));
OR2X2 OR2X2_2843 ( .A(core__abc_22172_new_n7666_), .B(core__abc_22172_new_n7665_), .Y(core__abc_22172_new_n7667_));
OR2X2 OR2X2_2844 ( .A(core__abc_22172_new_n7659_), .B(core__abc_22172_new_n7668_), .Y(core__abc_22172_new_n7669_));
OR2X2 OR2X2_2845 ( .A(core__abc_22172_new_n7658_), .B(core__abc_22172_new_n7667_), .Y(core__abc_22172_new_n7670_));
OR2X2 OR2X2_2846 ( .A(core__abc_22172_new_n7674_), .B(core__abc_22172_new_n7675_), .Y(core__abc_22172_new_n7676_));
OR2X2 OR2X2_2847 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n7676_), .Y(core__abc_22172_new_n7677_));
OR2X2 OR2X2_2848 ( .A(core__abc_22172_new_n7672_), .B(core__abc_22172_new_n7677_), .Y(core__abc_22172_new_n7678_));
OR2X2 OR2X2_2849 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_27_), .Y(core__abc_22172_new_n7679_));
OR2X2 OR2X2_285 ( .A(_abc_19873_new_n1519_), .B(_abc_19873_new_n1512_), .Y(_abc_19873_new_n1520_));
OR2X2 OR2X2_2850 ( .A(core__abc_22172_new_n7686_), .B(core__abc_22172_new_n7665_), .Y(core__abc_22172_new_n7687_));
OR2X2 OR2X2_2851 ( .A(core__abc_22172_new_n7687_), .B(core__abc_22172_new_n7685_), .Y(core__abc_22172_new_n7688_));
OR2X2 OR2X2_2852 ( .A(core__abc_22172_new_n7684_), .B(core__abc_22172_new_n7688_), .Y(core__abc_22172_new_n7689_));
OR2X2 OR2X2_2853 ( .A(core__abc_22172_new_n4901_), .B(core__abc_22172_new_n7691_), .Y(core__abc_22172_new_n7692_));
OR2X2 OR2X2_2854 ( .A(core__abc_22172_new_n4900_), .B(core_v1_reg_47_), .Y(core__abc_22172_new_n7693_));
OR2X2 OR2X2_2855 ( .A(core__abc_22172_new_n7696_), .B(core__abc_22172_new_n7697_), .Y(core__abc_22172_new_n7698_));
OR2X2 OR2X2_2856 ( .A(core__abc_22172_new_n7699_), .B(core__abc_22172_new_n7701_), .Y(core__abc_22172_new_n7702_));
OR2X2 OR2X2_2857 ( .A(core__abc_22172_new_n7705_), .B(core__abc_22172_new_n7706_), .Y(core__abc_22172_new_n7707_));
OR2X2 OR2X2_2858 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n7707_), .Y(core__abc_22172_new_n7708_));
OR2X2 OR2X2_2859 ( .A(core__abc_22172_new_n7704_), .B(core__abc_22172_new_n7708_), .Y(core__abc_22172_new_n7709_));
OR2X2 OR2X2_286 ( .A(_abc_19873_new_n1520_), .B(_abc_19873_new_n1511_), .Y(_abc_19873_new_n1521_));
OR2X2 OR2X2_2860 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_28_), .Y(core__abc_22172_new_n7710_));
OR2X2 OR2X2_2861 ( .A(core__abc_22172_new_n7714_), .B(core__abc_22172_new_n7715_), .Y(core__abc_22172_new_n7716_));
OR2X2 OR2X2_2862 ( .A(core__abc_22172_new_n7717_), .B(core__abc_22172_new_n7719_), .Y(core__abc_22172_new_n7720_));
OR2X2 OR2X2_2863 ( .A(core__abc_22172_new_n7701_), .B(core__abc_22172_new_n7696_), .Y(core__abc_22172_new_n7721_));
OR2X2 OR2X2_2864 ( .A(core__abc_22172_new_n7723_), .B(core__abc_22172_new_n7725_), .Y(core__abc_22172_new_n7726_));
OR2X2 OR2X2_2865 ( .A(core__abc_22172_new_n7730_), .B(core__abc_22172_new_n7731_), .Y(core__abc_22172_new_n7732_));
OR2X2 OR2X2_2866 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n7732_), .Y(core__abc_22172_new_n7733_));
OR2X2 OR2X2_2867 ( .A(core__abc_22172_new_n7728_), .B(core__abc_22172_new_n7733_), .Y(core__abc_22172_new_n7734_));
OR2X2 OR2X2_2868 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_29_), .Y(core__abc_22172_new_n7735_));
OR2X2 OR2X2_2869 ( .A(core__abc_22172_new_n7740_), .B(core__abc_22172_new_n7717_), .Y(core__abc_22172_new_n7741_));
OR2X2 OR2X2_287 ( .A(_abc_19873_new_n1523_), .B(_abc_19873_new_n1524_), .Y(_abc_19873_new_n1525_));
OR2X2 OR2X2_2870 ( .A(core__abc_22172_new_n7739_), .B(core__abc_22172_new_n7741_), .Y(core__abc_22172_new_n7742_));
OR2X2 OR2X2_2871 ( .A(core__abc_22172_new_n5009_), .B(core__abc_22172_new_n7744_), .Y(core__abc_22172_new_n7745_));
OR2X2 OR2X2_2872 ( .A(core__abc_22172_new_n4996_), .B(core_v1_reg_49_), .Y(core__abc_22172_new_n7746_));
OR2X2 OR2X2_2873 ( .A(core__abc_22172_new_n7750_), .B(core__abc_22172_new_n7749_), .Y(core__abc_22172_new_n7751_));
OR2X2 OR2X2_2874 ( .A(core__abc_22172_new_n7752_), .B(core__abc_22172_new_n7754_), .Y(core__abc_22172_new_n7755_));
OR2X2 OR2X2_2875 ( .A(core__abc_22172_new_n7759_), .B(core__abc_22172_new_n7760_), .Y(core__abc_22172_new_n7761_));
OR2X2 OR2X2_2876 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n7761_), .Y(core__abc_22172_new_n7762_));
OR2X2 OR2X2_2877 ( .A(core__abc_22172_new_n7757_), .B(core__abc_22172_new_n7762_), .Y(core__abc_22172_new_n7763_));
OR2X2 OR2X2_2878 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_30_), .Y(core__abc_22172_new_n7764_));
OR2X2 OR2X2_2879 ( .A(core__abc_22172_new_n7754_), .B(core__abc_22172_new_n7749_), .Y(core__abc_22172_new_n7767_));
OR2X2 OR2X2_288 ( .A(_abc_19873_new_n1192_), .B(_abc_19873_new_n1526_), .Y(_abc_19873_new_n1527_));
OR2X2 OR2X2_2880 ( .A(core__abc_22172_new_n7769_), .B(core__abc_22172_new_n7770_), .Y(core__abc_22172_new_n7771_));
OR2X2 OR2X2_2881 ( .A(core__abc_22172_new_n4498_), .B(core__abc_22172_new_n7772_), .Y(core__abc_22172_new_n7773_));
OR2X2 OR2X2_2882 ( .A(core__abc_22172_new_n4501_), .B(core__abc_22172_new_n7771_), .Y(core__abc_22172_new_n7774_));
OR2X2 OR2X2_2883 ( .A(core__abc_22172_new_n7767_), .B(core__abc_22172_new_n7775_), .Y(core__abc_22172_new_n7776_));
OR2X2 OR2X2_2884 ( .A(core__abc_22172_new_n7777_), .B(core__abc_22172_new_n7778_), .Y(core__abc_22172_new_n7779_));
OR2X2 OR2X2_2885 ( .A(core__abc_22172_new_n7782_), .B(core__abc_22172_new_n7783_), .Y(core__abc_22172_new_n7784_));
OR2X2 OR2X2_2886 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n7784_), .Y(core__abc_22172_new_n7785_));
OR2X2 OR2X2_2887 ( .A(core__abc_22172_new_n7781_), .B(core__abc_22172_new_n7785_), .Y(core__abc_22172_new_n7786_));
OR2X2 OR2X2_2888 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_31_), .Y(core__abc_22172_new_n7787_));
OR2X2 OR2X2_2889 ( .A(core__abc_22172_new_n6808_), .B(core__abc_22172_new_n7792_), .Y(core__abc_22172_new_n7793_));
OR2X2 OR2X2_289 ( .A(_abc_19873_new_n1527_), .B(_abc_19873_new_n1525_), .Y(_abc_19873_new_n1528_));
OR2X2 OR2X2_2890 ( .A(core__abc_22172_new_n7795_), .B(core__abc_22172_new_n7791_), .Y(core__abc_22172_new_n7796_));
OR2X2 OR2X2_2891 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n3196_), .Y(core__abc_22172_new_n7798_));
OR2X2 OR2X2_2892 ( .A(core__abc_22172_new_n7799_), .B(core__abc_22172_new_n7797_), .Y(core__abc_22172_new_n7800_));
OR2X2 OR2X2_2893 ( .A(core__abc_22172_new_n6811_), .B(core__abc_22172_new_n6808_), .Y(core__abc_22172_new_n7805_));
OR2X2 OR2X2_2894 ( .A(core__abc_22172_new_n7807_), .B(core__abc_22172_new_n7803_), .Y(core__abc_22172_new_n7808_));
OR2X2 OR2X2_2895 ( .A(core__abc_22172_new_n7802_), .B(core__abc_22172_new_n7809_), .Y(core__abc_22172_new_n7810_));
OR2X2 OR2X2_2896 ( .A(core__abc_22172_new_n6813_), .B(core__abc_22172_new_n6816_), .Y(core__abc_22172_new_n7813_));
OR2X2 OR2X2_2897 ( .A(core__abc_22172_new_n7817_), .B(core__abc_22172_new_n7818_), .Y(core__abc_22172_new_n7819_));
OR2X2 OR2X2_2898 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n7819_), .Y(core__abc_22172_new_n7820_));
OR2X2 OR2X2_2899 ( .A(core__abc_22172_new_n7815_), .B(core__abc_22172_new_n7820_), .Y(core__abc_22172_new_n7821_));
OR2X2 OR2X2_29 ( .A(_abc_19873_new_n974_), .B(_abc_19873_new_n975_), .Y(_abc_19873_new_n976_));
OR2X2 OR2X2_290 ( .A(_abc_19873_new_n1530_), .B(_abc_19873_new_n1531_), .Y(_abc_19873_new_n1532_));
OR2X2 OR2X2_2900 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_34_), .Y(core__abc_22172_new_n7822_));
OR2X2 OR2X2_2901 ( .A(core__abc_22172_new_n7829_), .B(core__abc_22172_new_n7830_), .Y(core__abc_22172_new_n7831_));
OR2X2 OR2X2_2902 ( .A(core__abc_22172_new_n7834_), .B(core__abc_22172_new_n7835_), .Y(core__abc_22172_new_n7836_));
OR2X2 OR2X2_2903 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n7836_), .Y(core__abc_22172_new_n7837_));
OR2X2 OR2X2_2904 ( .A(core__abc_22172_new_n7833_), .B(core__abc_22172_new_n7837_), .Y(core__abc_22172_new_n7838_));
OR2X2 OR2X2_2905 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_35_), .Y(core__abc_22172_new_n7839_));
OR2X2 OR2X2_2906 ( .A(core__abc_22172_new_n6820_), .B(core__abc_22172_new_n6823_), .Y(core__abc_22172_new_n7843_));
OR2X2 OR2X2_2907 ( .A(core__abc_22172_new_n7846_), .B(core__abc_22172_new_n7847_), .Y(core__abc_22172_new_n7848_));
OR2X2 OR2X2_2908 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n7848_), .Y(core__abc_22172_new_n7849_));
OR2X2 OR2X2_2909 ( .A(core__abc_22172_new_n7845_), .B(core__abc_22172_new_n7849_), .Y(core__abc_22172_new_n7850_));
OR2X2 OR2X2_291 ( .A(_abc_19873_new_n1532_), .B(_abc_19873_new_n1529_), .Y(_abc_19873_new_n1533_));
OR2X2 OR2X2_2910 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_36_), .Y(core__abc_22172_new_n7851_));
OR2X2 OR2X2_2911 ( .A(core__abc_22172_new_n7854_), .B(core__abc_22172_new_n7856_), .Y(core__abc_22172_new_n7859_));
OR2X2 OR2X2_2912 ( .A(core__abc_22172_new_n7864_), .B(core__abc_22172_new_n7865_), .Y(core__abc_22172_new_n7866_));
OR2X2 OR2X2_2913 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n7866_), .Y(core__abc_22172_new_n7867_));
OR2X2 OR2X2_2914 ( .A(core__abc_22172_new_n7862_), .B(core__abc_22172_new_n7867_), .Y(core__abc_22172_new_n7868_));
OR2X2 OR2X2_2915 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_37_), .Y(core__abc_22172_new_n7869_));
OR2X2 OR2X2_2916 ( .A(core__abc_22172_new_n6827_), .B(core__abc_22172_new_n6766_), .Y(core__abc_22172_new_n7874_));
OR2X2 OR2X2_2917 ( .A(core__abc_22172_new_n7878_), .B(core__abc_22172_new_n7879_), .Y(core__abc_22172_new_n7880_));
OR2X2 OR2X2_2918 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n7880_), .Y(core__abc_22172_new_n7881_));
OR2X2 OR2X2_2919 ( .A(core__abc_22172_new_n7876_), .B(core__abc_22172_new_n7881_), .Y(core__abc_22172_new_n7882_));
OR2X2 OR2X2_292 ( .A(_abc_19873_new_n1534_), .B(_abc_19873_new_n1535_), .Y(_abc_19873_new_n1536_));
OR2X2 OR2X2_2920 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_38_), .Y(core__abc_22172_new_n7883_));
OR2X2 OR2X2_2921 ( .A(core__abc_22172_new_n7872_), .B(core__abc_22172_new_n6759_), .Y(core__abc_22172_new_n7886_));
OR2X2 OR2X2_2922 ( .A(core__abc_22172_new_n7886_), .B(core__abc_22172_new_n6763_), .Y(core__abc_22172_new_n7887_));
OR2X2 OR2X2_2923 ( .A(core__abc_22172_new_n7889_), .B(core__abc_22172_new_n7888_), .Y(core__abc_22172_new_n7890_));
OR2X2 OR2X2_2924 ( .A(core__abc_22172_new_n7893_), .B(core__abc_22172_new_n7894_), .Y(core__abc_22172_new_n7895_));
OR2X2 OR2X2_2925 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n7895_), .Y(core__abc_22172_new_n7896_));
OR2X2 OR2X2_2926 ( .A(core__abc_22172_new_n7892_), .B(core__abc_22172_new_n7896_), .Y(core__abc_22172_new_n7897_));
OR2X2 OR2X2_2927 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_39_), .Y(core__abc_22172_new_n7898_));
OR2X2 OR2X2_2928 ( .A(core__abc_22172_new_n6829_), .B(core__abc_22172_new_n6833_), .Y(core__abc_22172_new_n7903_));
OR2X2 OR2X2_2929 ( .A(core__abc_22172_new_n7907_), .B(core__abc_22172_new_n7908_), .Y(core__abc_22172_new_n7909_));
OR2X2 OR2X2_293 ( .A(_abc_19873_new_n1537_), .B(_abc_19873_new_n1538_), .Y(_abc_19873_new_n1539_));
OR2X2 OR2X2_2930 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n7909_), .Y(core__abc_22172_new_n7910_));
OR2X2 OR2X2_2931 ( .A(core__abc_22172_new_n7905_), .B(core__abc_22172_new_n7910_), .Y(core__abc_22172_new_n7911_));
OR2X2 OR2X2_2932 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_40_), .Y(core__abc_22172_new_n7912_));
OR2X2 OR2X2_2933 ( .A(core__abc_22172_new_n7901_), .B(core__abc_22172_new_n6743_), .Y(core__abc_22172_new_n7916_));
OR2X2 OR2X2_2934 ( .A(core__abc_22172_new_n7918_), .B(core__abc_22172_new_n7919_), .Y(core__abc_22172_new_n7920_));
OR2X2 OR2X2_2935 ( .A(core__abc_22172_new_n7924_), .B(core__abc_22172_new_n7925_), .Y(core__abc_22172_new_n7926_));
OR2X2 OR2X2_2936 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n7926_), .Y(core__abc_22172_new_n7927_));
OR2X2 OR2X2_2937 ( .A(core__abc_22172_new_n7922_), .B(core__abc_22172_new_n7927_), .Y(core__abc_22172_new_n7928_));
OR2X2 OR2X2_2938 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_41_), .Y(core__abc_22172_new_n7929_));
OR2X2 OR2X2_2939 ( .A(core__abc_22172_new_n7932_), .B(core__abc_22172_new_n6745_), .Y(core__abc_22172_new_n7933_));
OR2X2 OR2X2_294 ( .A(_abc_19873_new_n1536_), .B(_abc_19873_new_n1539_), .Y(_abc_19873_new_n1540_));
OR2X2 OR2X2_2940 ( .A(core__abc_22172_new_n7933_), .B(core__abc_22172_new_n6728_), .Y(core__abc_22172_new_n7936_));
OR2X2 OR2X2_2941 ( .A(core__abc_22172_new_n7940_), .B(core__abc_22172_new_n7941_), .Y(core__abc_22172_new_n7942_));
OR2X2 OR2X2_2942 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n7942_), .Y(core__abc_22172_new_n7943_));
OR2X2 OR2X2_2943 ( .A(core__abc_22172_new_n7938_), .B(core__abc_22172_new_n7943_), .Y(core__abc_22172_new_n7944_));
OR2X2 OR2X2_2944 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_42_), .Y(core__abc_22172_new_n7945_));
OR2X2 OR2X2_2945 ( .A(core__abc_22172_new_n7934_), .B(core__abc_22172_new_n6722_), .Y(core__abc_22172_new_n7949_));
OR2X2 OR2X2_2946 ( .A(core__abc_22172_new_n7951_), .B(core__abc_22172_new_n7952_), .Y(core__abc_22172_new_n7953_));
OR2X2 OR2X2_2947 ( .A(core__abc_22172_new_n7956_), .B(core__abc_22172_new_n7957_), .Y(core__abc_22172_new_n7958_));
OR2X2 OR2X2_2948 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n7958_), .Y(core__abc_22172_new_n7959_));
OR2X2 OR2X2_2949 ( .A(core__abc_22172_new_n7955_), .B(core__abc_22172_new_n7959_), .Y(core__abc_22172_new_n7960_));
OR2X2 OR2X2_295 ( .A(_abc_19873_new_n1540_), .B(_abc_19873_new_n1533_), .Y(_abc_19873_new_n1541_));
OR2X2 OR2X2_2950 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_43_), .Y(core__abc_22172_new_n7961_));
OR2X2 OR2X2_2951 ( .A(core__abc_22172_new_n6837_), .B(core__abc_22172_new_n6706_), .Y(core__abc_22172_new_n7966_));
OR2X2 OR2X2_2952 ( .A(core__abc_22172_new_n7969_), .B(core__abc_22172_new_n7970_), .Y(core__abc_22172_new_n7971_));
OR2X2 OR2X2_2953 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n7971_), .Y(core__abc_22172_new_n7972_));
OR2X2 OR2X2_2954 ( .A(core__abc_22172_new_n7968_), .B(core__abc_22172_new_n7972_), .Y(core__abc_22172_new_n7973_));
OR2X2 OR2X2_2955 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_44_), .Y(core__abc_22172_new_n7974_));
OR2X2 OR2X2_2956 ( .A(core__abc_22172_new_n7980_), .B(core__abc_22172_new_n7981_), .Y(core__abc_22172_new_n7982_));
OR2X2 OR2X2_2957 ( .A(core__abc_22172_new_n7985_), .B(core__abc_22172_new_n7986_), .Y(core__abc_22172_new_n7987_));
OR2X2 OR2X2_2958 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n7987_), .Y(core__abc_22172_new_n7988_));
OR2X2 OR2X2_2959 ( .A(core__abc_22172_new_n7983_), .B(core__abc_22172_new_n7988_), .Y(core__abc_22172_new_n7989_));
OR2X2 OR2X2_296 ( .A(_abc_19873_new_n1541_), .B(_abc_19873_new_n1528_), .Y(_abc_19873_new_n1542_));
OR2X2 OR2X2_2960 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_45_), .Y(core__abc_22172_new_n7990_));
OR2X2 OR2X2_2961 ( .A(core__abc_22172_new_n7993_), .B(core__abc_22172_new_n6684_), .Y(core__abc_22172_new_n7994_));
OR2X2 OR2X2_2962 ( .A(core__abc_22172_new_n7994_), .B(core__abc_22172_new_n6677_), .Y(core__abc_22172_new_n7996_));
OR2X2 OR2X2_2963 ( .A(core__abc_22172_new_n7997_), .B(core__abc_22172_new_n7995_), .Y(core__abc_22172_new_n7998_));
OR2X2 OR2X2_2964 ( .A(core__abc_22172_new_n8002_), .B(core__abc_22172_new_n8003_), .Y(core__abc_22172_new_n8004_));
OR2X2 OR2X2_2965 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n8004_), .Y(core__abc_22172_new_n8005_));
OR2X2 OR2X2_2966 ( .A(core__abc_22172_new_n8000_), .B(core__abc_22172_new_n8005_), .Y(core__abc_22172_new_n8006_));
OR2X2 OR2X2_2967 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_46_), .Y(core__abc_22172_new_n8007_));
OR2X2 OR2X2_2968 ( .A(core__abc_22172_new_n7997_), .B(core__abc_22172_new_n6675_), .Y(core__abc_22172_new_n8011_));
OR2X2 OR2X2_2969 ( .A(core__abc_22172_new_n8013_), .B(core__abc_22172_new_n8014_), .Y(core__abc_22172_new_n8015_));
OR2X2 OR2X2_297 ( .A(_abc_19873_new_n1544_), .B(_abc_19873_new_n1545_), .Y(_abc_19873_new_n1546_));
OR2X2 OR2X2_2970 ( .A(core__abc_22172_new_n8018_), .B(core__abc_22172_new_n8019_), .Y(core__abc_22172_new_n8020_));
OR2X2 OR2X2_2971 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n8020_), .Y(core__abc_22172_new_n8021_));
OR2X2 OR2X2_2972 ( .A(core__abc_22172_new_n8017_), .B(core__abc_22172_new_n8021_), .Y(core__abc_22172_new_n8022_));
OR2X2 OR2X2_2973 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_47_), .Y(core__abc_22172_new_n8023_));
OR2X2 OR2X2_2974 ( .A(core__abc_22172_new_n8027_), .B(core__abc_22172_new_n8028_), .Y(core__abc_22172_new_n8029_));
OR2X2 OR2X2_2975 ( .A(core__abc_22172_new_n8033_), .B(core__abc_22172_new_n8034_), .Y(core__abc_22172_new_n8035_));
OR2X2 OR2X2_2976 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n8035_), .Y(core__abc_22172_new_n8036_));
OR2X2 OR2X2_2977 ( .A(core__abc_22172_new_n8031_), .B(core__abc_22172_new_n8036_), .Y(core__abc_22172_new_n8037_));
OR2X2 OR2X2_2978 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_48_), .Y(core__abc_22172_new_n8038_));
OR2X2 OR2X2_2979 ( .A(core__abc_22172_new_n8028_), .B(core__abc_22172_new_n6638_), .Y(core__abc_22172_new_n8042_));
OR2X2 OR2X2_298 ( .A(_abc_19873_new_n1547_), .B(_abc_19873_new_n1548_), .Y(_abc_19873_new_n1549_));
OR2X2 OR2X2_2980 ( .A(core__abc_22172_new_n8045_), .B(core__abc_22172_new_n8043_), .Y(core__abc_22172_new_n8046_));
OR2X2 OR2X2_2981 ( .A(core__abc_22172_new_n8048_), .B(core__abc_22172_new_n8049_), .Y(core__abc_22172_new_n8050_));
OR2X2 OR2X2_2982 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n8050_), .Y(core__abc_22172_new_n8051_));
OR2X2 OR2X2_2983 ( .A(core__abc_22172_new_n8047_), .B(core__abc_22172_new_n8051_), .Y(core__abc_22172_new_n8052_));
OR2X2 OR2X2_2984 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_49_), .Y(core__abc_22172_new_n8053_));
OR2X2 OR2X2_2985 ( .A(core__abc_22172_new_n8056_), .B(core__abc_22172_new_n6644_), .Y(core__abc_22172_new_n8057_));
OR2X2 OR2X2_2986 ( .A(core__abc_22172_new_n8057_), .B(core__abc_22172_new_n6616_), .Y(core__abc_22172_new_n8060_));
OR2X2 OR2X2_2987 ( .A(core__abc_22172_new_n8063_), .B(core__abc_22172_new_n8064_), .Y(core__abc_22172_new_n8065_));
OR2X2 OR2X2_2988 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n8065_), .Y(core__abc_22172_new_n8066_));
OR2X2 OR2X2_2989 ( .A(core__abc_22172_new_n8062_), .B(core__abc_22172_new_n8066_), .Y(core__abc_22172_new_n8067_));
OR2X2 OR2X2_299 ( .A(_abc_19873_new_n1546_), .B(_abc_19873_new_n1549_), .Y(_abc_19873_new_n1550_));
OR2X2 OR2X2_2990 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_50_), .Y(core__abc_22172_new_n8068_));
OR2X2 OR2X2_2991 ( .A(core__abc_22172_new_n8072_), .B(core__abc_22172_new_n8071_), .Y(core__abc_22172_new_n8075_));
OR2X2 OR2X2_2992 ( .A(core__abc_22172_new_n8079_), .B(core__abc_22172_new_n8080_), .Y(core__abc_22172_new_n8081_));
OR2X2 OR2X2_2993 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n8081_), .Y(core__abc_22172_new_n8082_));
OR2X2 OR2X2_2994 ( .A(core__abc_22172_new_n8077_), .B(core__abc_22172_new_n8082_), .Y(core__abc_22172_new_n8083_));
OR2X2 OR2X2_2995 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_51_), .Y(core__abc_22172_new_n8084_));
OR2X2 OR2X2_2996 ( .A(core__abc_22172_new_n8092_), .B(core__abc_22172_new_n8090_), .Y(core__abc_22172_new_n8093_));
OR2X2 OR2X2_2997 ( .A(core__abc_22172_new_n8097_), .B(core__abc_22172_new_n8098_), .Y(core__abc_22172_new_n8099_));
OR2X2 OR2X2_2998 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n8099_), .Y(core__abc_22172_new_n8100_));
OR2X2 OR2X2_2999 ( .A(core__abc_22172_new_n8095_), .B(core__abc_22172_new_n8100_), .Y(core__abc_22172_new_n8101_));
OR2X2 OR2X2_3 ( .A(_abc_19873_new_n902_), .B(_abc_19873_new_n908_), .Y(_abc_19873_new_n909_));
OR2X2 OR2X2_30 ( .A(_abc_19873_new_n976_), .B(_abc_19873_new_n977_), .Y(_abc_19873_new_n978_));
OR2X2 OR2X2_300 ( .A(_abc_19873_new_n1551_), .B(_abc_19873_new_n1552_), .Y(_abc_19873_new_n1553_));
OR2X2 OR2X2_3000 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_52_), .Y(core__abc_22172_new_n8102_));
OR2X2 OR2X2_3001 ( .A(core__abc_22172_new_n8090_), .B(core__abc_22172_new_n6602_), .Y(core__abc_22172_new_n8106_));
OR2X2 OR2X2_3002 ( .A(core__abc_22172_new_n8106_), .B(core__abc_22172_new_n8105_), .Y(core__abc_22172_new_n8109_));
OR2X2 OR2X2_3003 ( .A(core__abc_22172_new_n8114_), .B(core__abc_22172_new_n8115_), .Y(core__abc_22172_new_n8116_));
OR2X2 OR2X2_3004 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n8116_), .Y(core__abc_22172_new_n8117_));
OR2X2 OR2X2_3005 ( .A(core__abc_22172_new_n8112_), .B(core__abc_22172_new_n8117_), .Y(core__abc_22172_new_n8118_));
OR2X2 OR2X2_3006 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_53_), .Y(core__abc_22172_new_n8119_));
OR2X2 OR2X2_3007 ( .A(core__abc_22172_new_n8122_), .B(core__abc_22172_new_n6655_), .Y(core__abc_22172_new_n8123_));
OR2X2 OR2X2_3008 ( .A(core__abc_22172_new_n8123_), .B(core__abc_22172_new_n6587_), .Y(core__abc_22172_new_n8126_));
OR2X2 OR2X2_3009 ( .A(core__abc_22172_new_n8130_), .B(core__abc_22172_new_n8131_), .Y(core__abc_22172_new_n8132_));
OR2X2 OR2X2_301 ( .A(_abc_19873_new_n1554_), .B(_abc_19873_new_n1555_), .Y(_abc_19873_new_n1556_));
OR2X2 OR2X2_3010 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n8132_), .Y(core__abc_22172_new_n8133_));
OR2X2 OR2X2_3011 ( .A(core__abc_22172_new_n8128_), .B(core__abc_22172_new_n8133_), .Y(core__abc_22172_new_n8134_));
OR2X2 OR2X2_3012 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_54_), .Y(core__abc_22172_new_n8135_));
OR2X2 OR2X2_3013 ( .A(core__abc_22172_new_n8124_), .B(core__abc_22172_new_n6584_), .Y(core__abc_22172_new_n8139_));
OR2X2 OR2X2_3014 ( .A(core__abc_22172_new_n8141_), .B(core__abc_22172_new_n8142_), .Y(core__abc_22172_new_n8143_));
OR2X2 OR2X2_3015 ( .A(core__abc_22172_new_n8146_), .B(core__abc_22172_new_n8147_), .Y(core__abc_22172_new_n8148_));
OR2X2 OR2X2_3016 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n8148_), .Y(core__abc_22172_new_n8149_));
OR2X2 OR2X2_3017 ( .A(core__abc_22172_new_n8145_), .B(core__abc_22172_new_n8149_), .Y(core__abc_22172_new_n8150_));
OR2X2 OR2X2_3018 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_55_), .Y(core__abc_22172_new_n8151_));
OR2X2 OR2X2_3019 ( .A(core__abc_22172_new_n8155_), .B(core__abc_22172_new_n8156_), .Y(core__abc_22172_new_n8157_));
OR2X2 OR2X2_302 ( .A(_abc_19873_new_n1553_), .B(_abc_19873_new_n1556_), .Y(_abc_19873_new_n1557_));
OR2X2 OR2X2_3020 ( .A(core__abc_22172_new_n8160_), .B(core__abc_22172_new_n8161_), .Y(core__abc_22172_new_n8162_));
OR2X2 OR2X2_3021 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n8162_), .Y(core__abc_22172_new_n8163_));
OR2X2 OR2X2_3022 ( .A(core__abc_22172_new_n8159_), .B(core__abc_22172_new_n8163_), .Y(core__abc_22172_new_n8164_));
OR2X2 OR2X2_3023 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_56_), .Y(core__abc_22172_new_n8165_));
OR2X2 OR2X2_3024 ( .A(core__abc_22172_new_n8170_), .B(core__abc_22172_new_n8168_), .Y(core__abc_22172_new_n8173_));
OR2X2 OR2X2_3025 ( .A(core__abc_22172_new_n8176_), .B(core__abc_22172_new_n8177_), .Y(core__abc_22172_new_n8178_));
OR2X2 OR2X2_3026 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n8178_), .Y(core__abc_22172_new_n8179_));
OR2X2 OR2X2_3027 ( .A(core__abc_22172_new_n8175_), .B(core__abc_22172_new_n8179_), .Y(core__abc_22172_new_n8180_));
OR2X2 OR2X2_3028 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_57_), .Y(core__abc_22172_new_n8181_));
OR2X2 OR2X2_3029 ( .A(core__abc_22172_new_n8184_), .B(core__abc_22172_new_n6544_), .Y(core__abc_22172_new_n8185_));
OR2X2 OR2X2_303 ( .A(_abc_19873_new_n1558_), .B(_abc_19873_new_n1559_), .Y(_abc_19873_new_n1560_));
OR2X2 OR2X2_3030 ( .A(core__abc_22172_new_n8185_), .B(core__abc_22172_new_n6524_), .Y(core__abc_22172_new_n8188_));
OR2X2 OR2X2_3031 ( .A(core__abc_22172_new_n8192_), .B(core__abc_22172_new_n8193_), .Y(core__abc_22172_new_n8194_));
OR2X2 OR2X2_3032 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n8194_), .Y(core__abc_22172_new_n8195_));
OR2X2 OR2X2_3033 ( .A(core__abc_22172_new_n8190_), .B(core__abc_22172_new_n8195_), .Y(core__abc_22172_new_n8196_));
OR2X2 OR2X2_3034 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_58_), .Y(core__abc_22172_new_n8197_));
OR2X2 OR2X2_3035 ( .A(core__abc_22172_new_n8203_), .B(core__abc_22172_new_n8204_), .Y(core__abc_22172_new_n8205_));
OR2X2 OR2X2_3036 ( .A(core__abc_22172_new_n8208_), .B(core__abc_22172_new_n8209_), .Y(core__abc_22172_new_n8210_));
OR2X2 OR2X2_3037 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n8210_), .Y(core__abc_22172_new_n8211_));
OR2X2 OR2X2_3038 ( .A(core__abc_22172_new_n8206_), .B(core__abc_22172_new_n8211_), .Y(core__abc_22172_new_n8212_));
OR2X2 OR2X2_3039 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_59_), .Y(core__abc_22172_new_n8213_));
OR2X2 OR2X2_304 ( .A(_abc_19873_new_n1039_), .B(_abc_19873_new_n1560_), .Y(_abc_19873_new_n1561_));
OR2X2 OR2X2_3040 ( .A(core__abc_22172_new_n8220_), .B(core__abc_22172_new_n8221_), .Y(core__abc_22172_new_n8222_));
OR2X2 OR2X2_3041 ( .A(core__abc_22172_new_n8225_), .B(core__abc_22172_new_n8226_), .Y(core__abc_22172_new_n8227_));
OR2X2 OR2X2_3042 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n8227_), .Y(core__abc_22172_new_n8228_));
OR2X2 OR2X2_3043 ( .A(core__abc_22172_new_n8224_), .B(core__abc_22172_new_n8228_), .Y(core__abc_22172_new_n8229_));
OR2X2 OR2X2_3044 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_60_), .Y(core__abc_22172_new_n8230_));
OR2X2 OR2X2_3045 ( .A(core__abc_22172_new_n8220_), .B(core__abc_22172_new_n6501_), .Y(core__abc_22172_new_n8234_));
OR2X2 OR2X2_3046 ( .A(core__abc_22172_new_n8234_), .B(core__abc_22172_new_n8233_), .Y(core__abc_22172_new_n8237_));
OR2X2 OR2X2_3047 ( .A(core__abc_22172_new_n8242_), .B(core__abc_22172_new_n8243_), .Y(core__abc_22172_new_n8244_));
OR2X2 OR2X2_3048 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n8244_), .Y(core__abc_22172_new_n8245_));
OR2X2 OR2X2_3049 ( .A(core__abc_22172_new_n8240_), .B(core__abc_22172_new_n8245_), .Y(core__abc_22172_new_n8246_));
OR2X2 OR2X2_305 ( .A(_abc_19873_new_n1561_), .B(_abc_19873_new_n1557_), .Y(_abc_19873_new_n1562_));
OR2X2 OR2X2_3050 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_61_), .Y(core__abc_22172_new_n8247_));
OR2X2 OR2X2_3051 ( .A(core__abc_22172_new_n8250_), .B(core__abc_22172_new_n6554_), .Y(core__abc_22172_new_n8251_));
OR2X2 OR2X2_3052 ( .A(core__abc_22172_new_n8251_), .B(core__abc_22172_new_n6483_), .Y(core__abc_22172_new_n8254_));
OR2X2 OR2X2_3053 ( .A(core__abc_22172_new_n8258_), .B(core__abc_22172_new_n8259_), .Y(core__abc_22172_new_n8260_));
OR2X2 OR2X2_3054 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n8260_), .Y(core__abc_22172_new_n8261_));
OR2X2 OR2X2_3055 ( .A(core__abc_22172_new_n8256_), .B(core__abc_22172_new_n8261_), .Y(core__abc_22172_new_n8262_));
OR2X2 OR2X2_3056 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_62_), .Y(core__abc_22172_new_n8263_));
OR2X2 OR2X2_3057 ( .A(core__abc_22172_new_n8267_), .B(core__abc_22172_new_n8266_), .Y(core__abc_22172_new_n8269_));
OR2X2 OR2X2_3058 ( .A(core__abc_22172_new_n8270_), .B(core__abc_22172_new_n8268_), .Y(core__abc_22172_new_n8271_));
OR2X2 OR2X2_3059 ( .A(core__abc_22172_new_n8274_), .B(core__abc_22172_new_n8275_), .Y(core__abc_22172_new_n8276_));
OR2X2 OR2X2_306 ( .A(_abc_19873_new_n1562_), .B(_abc_19873_new_n1550_), .Y(_abc_19873_new_n1563_));
OR2X2 OR2X2_3060 ( .A(core__abc_22172_new_n6880_), .B(core__abc_22172_new_n8276_), .Y(core__abc_22172_new_n8277_));
OR2X2 OR2X2_3061 ( .A(core__abc_22172_new_n8273_), .B(core__abc_22172_new_n8277_), .Y(core__abc_22172_new_n8278_));
OR2X2 OR2X2_3062 ( .A(core__abc_22172_new_n7114_), .B(core_v2_reg_63_), .Y(core__abc_22172_new_n8279_));
OR2X2 OR2X2_3063 ( .A(core__abc_22172_new_n3219_), .B(core__abc_22172_new_n8290_), .Y(core__abc_22172_new_n8291_));
OR2X2 OR2X2_3064 ( .A(core__abc_22172_new_n8287_), .B(core__abc_22172_new_n8291_), .Y(core__abc_22172_new_n8292_));
OR2X2 OR2X2_3065 ( .A(core__abc_22172_new_n8292_), .B(core__abc_22172_new_n8285_), .Y(core__abc_22172_new_n8293_));
OR2X2 OR2X2_3066 ( .A(core__abc_22172_new_n8294_), .B(core__abc_22172_new_n8284_), .Y(core__abc_22172_new_n8295_));
OR2X2 OR2X2_3067 ( .A(core__abc_22172_new_n7342_), .B(core__abc_22172_new_n7806_), .Y(core__abc_22172_new_n8297_));
OR2X2 OR2X2_3068 ( .A(core__abc_22172_new_n7341_), .B(core__abc_22172_new_n8298_), .Y(core__abc_22172_new_n8299_));
OR2X2 OR2X2_3069 ( .A(core_key_65_), .B(core_long), .Y(core__abc_22172_new_n8302_));
OR2X2 OR2X2_307 ( .A(_abc_19873_new_n1565_), .B(_abc_19873_new_n1566_), .Y(_abc_19873_new_n1567_));
OR2X2 OR2X2_3070 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8307_), .Y(core__abc_22172_new_n8308_));
OR2X2 OR2X2_3071 ( .A(core__abc_22172_new_n8308_), .B(core__abc_22172_new_n8306_), .Y(core__abc_22172_new_n8309_));
OR2X2 OR2X2_3072 ( .A(core__abc_22172_new_n8301_), .B(core__abc_22172_new_n8309_), .Y(core__abc_22172_new_n8310_));
OR2X2 OR2X2_3073 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_1_), .Y(core__abc_22172_new_n8311_));
OR2X2 OR2X2_3074 ( .A(core__abc_22172_new_n8319_), .B(core_long), .Y(core__abc_22172_new_n8320_));
OR2X2 OR2X2_3075 ( .A(core__abc_22172_new_n6870_), .B(core_key_66_), .Y(core__abc_22172_new_n8321_));
OR2X2 OR2X2_3076 ( .A(core__abc_22172_new_n8323_), .B(core__abc_22172_new_n8324_), .Y(core__abc_22172_new_n8325_));
OR2X2 OR2X2_3077 ( .A(core__abc_22172_new_n8318_), .B(core__abc_22172_new_n8325_), .Y(core__abc_22172_new_n8326_));
OR2X2 OR2X2_3078 ( .A(core__abc_22172_new_n8326_), .B(core__abc_22172_new_n8317_), .Y(core__abc_22172_new_n8327_));
OR2X2 OR2X2_3079 ( .A(core__abc_22172_new_n8328_), .B(core__abc_22172_new_n8314_), .Y(core__abc_22172_new_n8329_));
OR2X2 OR2X2_308 ( .A(_abc_19873_new_n1038_), .B(_abc_19873_new_n1568_), .Y(_abc_19873_new_n1569_));
OR2X2 OR2X2_3080 ( .A(core__abc_22172_new_n7394_), .B(core__abc_22172_new_n7833_), .Y(core__abc_22172_new_n8332_));
OR2X2 OR2X2_3081 ( .A(core__abc_22172_new_n7393_), .B(core__abc_22172_new_n8333_), .Y(core__abc_22172_new_n8334_));
OR2X2 OR2X2_3082 ( .A(core__abc_22172_new_n6870_), .B(core_key_67_), .Y(core__abc_22172_new_n8336_));
OR2X2 OR2X2_3083 ( .A(core__abc_22172_new_n8337_), .B(core_long), .Y(core__abc_22172_new_n8338_));
OR2X2 OR2X2_3084 ( .A(core__abc_22172_new_n8340_), .B(core__abc_22172_new_n8341_), .Y(core__abc_22172_new_n8342_));
OR2X2 OR2X2_3085 ( .A(core__abc_22172_new_n8335_), .B(core__abc_22172_new_n8342_), .Y(core__abc_22172_new_n8343_));
OR2X2 OR2X2_3086 ( .A(core__abc_22172_new_n8344_), .B(core__abc_22172_new_n8331_), .Y(core__abc_22172_new_n8345_));
OR2X2 OR2X2_3087 ( .A(core__abc_22172_new_n8352_), .B(core__abc_22172_new_n8353_), .Y(core__abc_22172_new_n8354_));
OR2X2 OR2X2_3088 ( .A(core__abc_22172_new_n8351_), .B(core__abc_22172_new_n8354_), .Y(core__abc_22172_new_n8355_));
OR2X2 OR2X2_3089 ( .A(core__abc_22172_new_n8355_), .B(core__abc_22172_new_n8350_), .Y(core__abc_22172_new_n8356_));
OR2X2 OR2X2_309 ( .A(_abc_19873_new_n1569_), .B(_abc_19873_new_n1567_), .Y(_abc_19873_new_n1570_));
OR2X2 OR2X2_3090 ( .A(core__abc_22172_new_n8357_), .B(core__abc_22172_new_n8347_), .Y(core__abc_22172_new_n8358_));
OR2X2 OR2X2_3091 ( .A(core__abc_22172_new_n8360_), .B(core__abc_22172_new_n7459_), .Y(core__abc_22172_new_n8361_));
OR2X2 OR2X2_3092 ( .A(core__abc_22172_new_n7862_), .B(core__abc_22172_new_n7460_), .Y(core__abc_22172_new_n8362_));
OR2X2 OR2X2_3093 ( .A(core__abc_22172_new_n3525_), .B(core_long), .Y(core__abc_22172_new_n8364_));
OR2X2 OR2X2_3094 ( .A(core__abc_22172_new_n6870_), .B(core_key_69_), .Y(core__abc_22172_new_n8365_));
OR2X2 OR2X2_3095 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8368_), .Y(core__abc_22172_new_n8369_));
OR2X2 OR2X2_3096 ( .A(core__abc_22172_new_n8369_), .B(core__abc_22172_new_n8367_), .Y(core__abc_22172_new_n8370_));
OR2X2 OR2X2_3097 ( .A(core__abc_22172_new_n8363_), .B(core__abc_22172_new_n8370_), .Y(core__abc_22172_new_n8371_));
OR2X2 OR2X2_3098 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_5_), .Y(core__abc_22172_new_n8372_));
OR2X2 OR2X2_3099 ( .A(core__abc_22172_new_n3592_), .B(core_long), .Y(core__abc_22172_new_n8380_));
OR2X2 OR2X2_31 ( .A(_abc_19873_new_n979_), .B(_abc_19873_new_n980_), .Y(_abc_19873_new_n981_));
OR2X2 OR2X2_310 ( .A(_abc_19873_new_n1572_), .B(_abc_19873_new_n1573_), .Y(_abc_19873_new_n1574_));
OR2X2 OR2X2_3100 ( .A(core__abc_22172_new_n6870_), .B(core_key_70_), .Y(core__abc_22172_new_n8381_));
OR2X2 OR2X2_3101 ( .A(core__abc_22172_new_n8383_), .B(core__abc_22172_new_n8384_), .Y(core__abc_22172_new_n8385_));
OR2X2 OR2X2_3102 ( .A(core__abc_22172_new_n8379_), .B(core__abc_22172_new_n8385_), .Y(core__abc_22172_new_n8386_));
OR2X2 OR2X2_3103 ( .A(core__abc_22172_new_n8386_), .B(core__abc_22172_new_n8376_), .Y(core__abc_22172_new_n8387_));
OR2X2 OR2X2_3104 ( .A(core__abc_22172_new_n8388_), .B(core__abc_22172_new_n8375_), .Y(core__abc_22172_new_n8389_));
OR2X2 OR2X2_3105 ( .A(core__abc_22172_new_n8392_), .B(core__abc_22172_new_n7510_), .Y(core__abc_22172_new_n8393_));
OR2X2 OR2X2_3106 ( .A(core__abc_22172_new_n7891_), .B(core__abc_22172_new_n7511_), .Y(core__abc_22172_new_n8394_));
OR2X2 OR2X2_3107 ( .A(core_key_71_), .B(core_long), .Y(core__abc_22172_new_n8399_));
OR2X2 OR2X2_3108 ( .A(core__abc_22172_new_n8401_), .B(core__abc_22172_new_n8402_), .Y(core__abc_22172_new_n8403_));
OR2X2 OR2X2_3109 ( .A(core__abc_22172_new_n8396_), .B(core__abc_22172_new_n8403_), .Y(core__abc_22172_new_n8404_));
OR2X2 OR2X2_311 ( .A(_abc_19873_new_n1574_), .B(_abc_19873_new_n1571_), .Y(_abc_19873_new_n1575_));
OR2X2 OR2X2_3110 ( .A(core__abc_22172_new_n8405_), .B(core__abc_22172_new_n8391_), .Y(core__abc_22172_new_n8406_));
OR2X2 OR2X2_3111 ( .A(core__abc_22172_new_n8409_), .B(core__abc_22172_new_n7541_), .Y(core__abc_22172_new_n8410_));
OR2X2 OR2X2_3112 ( .A(core__abc_22172_new_n7542_), .B(core__abc_22172_new_n7905_), .Y(core__abc_22172_new_n8411_));
OR2X2 OR2X2_3113 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8413_), .Y(core__abc_22172_new_n8414_));
OR2X2 OR2X2_3114 ( .A(core__abc_22172_new_n8414_), .B(core__abc_22172_new_n3723_), .Y(core__abc_22172_new_n8415_));
OR2X2 OR2X2_3115 ( .A(core__abc_22172_new_n8412_), .B(core__abc_22172_new_n8415_), .Y(core__abc_22172_new_n8416_));
OR2X2 OR2X2_3116 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_8_), .Y(core__abc_22172_new_n8417_));
OR2X2 OR2X2_3117 ( .A(core__abc_22172_new_n7921_), .B(core__abc_22172_new_n7582_), .Y(core__abc_22172_new_n8420_));
OR2X2 OR2X2_3118 ( .A(core__abc_22172_new_n7920_), .B(core__abc_22172_new_n7581_), .Y(core__abc_22172_new_n8421_));
OR2X2 OR2X2_3119 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8426_), .Y(core__abc_22172_new_n8427_));
OR2X2 OR2X2_312 ( .A(_abc_19873_new_n1576_), .B(_abc_19873_new_n1577_), .Y(_abc_19873_new_n1578_));
OR2X2 OR2X2_3120 ( .A(core__abc_22172_new_n8427_), .B(core__abc_22172_new_n8425_), .Y(core__abc_22172_new_n8428_));
OR2X2 OR2X2_3121 ( .A(core__abc_22172_new_n8423_), .B(core__abc_22172_new_n8428_), .Y(core__abc_22172_new_n8429_));
OR2X2 OR2X2_3122 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_9_), .Y(core__abc_22172_new_n8430_));
OR2X2 OR2X2_3123 ( .A(core__abc_22172_new_n8433_), .B(core__abc_22172_new_n7608_), .Y(core__abc_22172_new_n8434_));
OR2X2 OR2X2_3124 ( .A(core__abc_22172_new_n7937_), .B(core__abc_22172_new_n7605_), .Y(core__abc_22172_new_n8435_));
OR2X2 OR2X2_3125 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8438_), .Y(core__abc_22172_new_n8439_));
OR2X2 OR2X2_3126 ( .A(core__abc_22172_new_n8439_), .B(core__abc_22172_new_n3856_), .Y(core__abc_22172_new_n8440_));
OR2X2 OR2X2_3127 ( .A(core__abc_22172_new_n8437_), .B(core__abc_22172_new_n8440_), .Y(core__abc_22172_new_n8441_));
OR2X2 OR2X2_3128 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_10_), .Y(core__abc_22172_new_n8442_));
OR2X2 OR2X2_3129 ( .A(core__abc_22172_new_n7954_), .B(core__abc_22172_new_n7631_), .Y(core__abc_22172_new_n8445_));
OR2X2 OR2X2_313 ( .A(_abc_19873_new_n1579_), .B(_abc_19873_new_n1580_), .Y(_abc_19873_new_n1581_));
OR2X2 OR2X2_3130 ( .A(core__abc_22172_new_n7953_), .B(core__abc_22172_new_n7630_), .Y(core__abc_22172_new_n8446_));
OR2X2 OR2X2_3131 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8451_), .Y(core__abc_22172_new_n8452_));
OR2X2 OR2X2_3132 ( .A(core__abc_22172_new_n8452_), .B(core__abc_22172_new_n8450_), .Y(core__abc_22172_new_n8453_));
OR2X2 OR2X2_3133 ( .A(core__abc_22172_new_n8448_), .B(core__abc_22172_new_n8453_), .Y(core__abc_22172_new_n8454_));
OR2X2 OR2X2_3134 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_11_), .Y(core__abc_22172_new_n8455_));
OR2X2 OR2X2_3135 ( .A(core__abc_22172_new_n8458_), .B(core__abc_22172_new_n7663_), .Y(core__abc_22172_new_n8459_));
OR2X2 OR2X2_3136 ( .A(core__abc_22172_new_n7967_), .B(core__abc_22172_new_n7664_), .Y(core__abc_22172_new_n8460_));
OR2X2 OR2X2_3137 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8463_), .Y(core__abc_22172_new_n8464_));
OR2X2 OR2X2_3138 ( .A(core__abc_22172_new_n8464_), .B(core__abc_22172_new_n3984_), .Y(core__abc_22172_new_n8465_));
OR2X2 OR2X2_3139 ( .A(core__abc_22172_new_n8462_), .B(core__abc_22172_new_n8465_), .Y(core__abc_22172_new_n8466_));
OR2X2 OR2X2_314 ( .A(_abc_19873_new_n1578_), .B(_abc_19873_new_n1581_), .Y(_abc_19873_new_n1582_));
OR2X2 OR2X2_3140 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_12_), .Y(core__abc_22172_new_n8467_));
OR2X2 OR2X2_3141 ( .A(core__abc_22172_new_n7982_), .B(core__abc_22172_new_n7695_), .Y(core__abc_22172_new_n8470_));
OR2X2 OR2X2_3142 ( .A(core__abc_22172_new_n8471_), .B(core__abc_22172_new_n7694_), .Y(core__abc_22172_new_n8472_));
OR2X2 OR2X2_3143 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8475_), .Y(core__abc_22172_new_n8476_));
OR2X2 OR2X2_3144 ( .A(core__abc_22172_new_n8476_), .B(core__abc_22172_new_n4051_), .Y(core__abc_22172_new_n8477_));
OR2X2 OR2X2_3145 ( .A(core__abc_22172_new_n8474_), .B(core__abc_22172_new_n8477_), .Y(core__abc_22172_new_n8478_));
OR2X2 OR2X2_3146 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_13_), .Y(core__abc_22172_new_n8479_));
OR2X2 OR2X2_3147 ( .A(core__abc_22172_new_n7999_), .B(core__abc_22172_new_n7716_), .Y(core__abc_22172_new_n8482_));
OR2X2 OR2X2_3148 ( .A(core__abc_22172_new_n7998_), .B(core__abc_22172_new_n7718_), .Y(core__abc_22172_new_n8483_));
OR2X2 OR2X2_3149 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8486_), .Y(core__abc_22172_new_n8487_));
OR2X2 OR2X2_315 ( .A(_abc_19873_new_n1582_), .B(_abc_19873_new_n1575_), .Y(_abc_19873_new_n1583_));
OR2X2 OR2X2_3150 ( .A(core__abc_22172_new_n8487_), .B(core__abc_22172_new_n4115_), .Y(core__abc_22172_new_n8488_));
OR2X2 OR2X2_3151 ( .A(core__abc_22172_new_n8485_), .B(core__abc_22172_new_n8488_), .Y(core__abc_22172_new_n8489_));
OR2X2 OR2X2_3152 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_14_), .Y(core__abc_22172_new_n8490_));
OR2X2 OR2X2_3153 ( .A(core__abc_22172_new_n8016_), .B(core__abc_22172_new_n7748_), .Y(core__abc_22172_new_n8493_));
OR2X2 OR2X2_3154 ( .A(core__abc_22172_new_n8015_), .B(core__abc_22172_new_n7747_), .Y(core__abc_22172_new_n8494_));
OR2X2 OR2X2_3155 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8497_), .Y(core__abc_22172_new_n8498_));
OR2X2 OR2X2_3156 ( .A(core__abc_22172_new_n8498_), .B(core__abc_22172_new_n4174_), .Y(core__abc_22172_new_n8499_));
OR2X2 OR2X2_3157 ( .A(core__abc_22172_new_n8496_), .B(core__abc_22172_new_n8499_), .Y(core__abc_22172_new_n8500_));
OR2X2 OR2X2_3158 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_15_), .Y(core__abc_22172_new_n8501_));
OR2X2 OR2X2_3159 ( .A(core__abc_22172_new_n8029_), .B(core__abc_22172_new_n7771_), .Y(core__abc_22172_new_n8504_));
OR2X2 OR2X2_316 ( .A(_abc_19873_new_n1583_), .B(_abc_19873_new_n1570_), .Y(_abc_19873_new_n1584_));
OR2X2 OR2X2_3160 ( .A(core__abc_22172_new_n8030_), .B(core__abc_22172_new_n7772_), .Y(core__abc_22172_new_n8505_));
OR2X2 OR2X2_3161 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8508_), .Y(core__abc_22172_new_n8509_));
OR2X2 OR2X2_3162 ( .A(core__abc_22172_new_n8509_), .B(core__abc_22172_new_n4259_), .Y(core__abc_22172_new_n8510_));
OR2X2 OR2X2_3163 ( .A(core__abc_22172_new_n8507_), .B(core__abc_22172_new_n8510_), .Y(core__abc_22172_new_n8511_));
OR2X2 OR2X2_3164 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_16_), .Y(core__abc_22172_new_n8512_));
OR2X2 OR2X2_3165 ( .A(core__abc_22172_new_n8515_), .B(core__abc_22172_new_n6806_), .Y(core__abc_22172_new_n8516_));
OR2X2 OR2X2_3166 ( .A(core__abc_22172_new_n8046_), .B(core__abc_22172_new_n6807_), .Y(core__abc_22172_new_n8517_));
OR2X2 OR2X2_3167 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8520_), .Y(core__abc_22172_new_n8521_));
OR2X2 OR2X2_3168 ( .A(core__abc_22172_new_n8521_), .B(core__abc_22172_new_n4326_), .Y(core__abc_22172_new_n8522_));
OR2X2 OR2X2_3169 ( .A(core__abc_22172_new_n8519_), .B(core__abc_22172_new_n8522_), .Y(core__abc_22172_new_n8523_));
OR2X2 OR2X2_317 ( .A(_abc_19873_new_n1586_), .B(_abc_19873_new_n1587_), .Y(_abc_19873_new_n1588_));
OR2X2 OR2X2_3170 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_17_), .Y(core__abc_22172_new_n8524_));
OR2X2 OR2X2_3171 ( .A(core__abc_22172_new_n8527_), .B(core__abc_22172_new_n6800_), .Y(core__abc_22172_new_n8528_));
OR2X2 OR2X2_3172 ( .A(core__abc_22172_new_n8061_), .B(core__abc_22172_new_n6809_), .Y(core__abc_22172_new_n8529_));
OR2X2 OR2X2_3173 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8532_), .Y(core__abc_22172_new_n8533_));
OR2X2 OR2X2_3174 ( .A(core__abc_22172_new_n8533_), .B(core__abc_22172_new_n4386_), .Y(core__abc_22172_new_n8534_));
OR2X2 OR2X2_3175 ( .A(core__abc_22172_new_n8531_), .B(core__abc_22172_new_n8534_), .Y(core__abc_22172_new_n8535_));
OR2X2 OR2X2_3176 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_18_), .Y(core__abc_22172_new_n8536_));
OR2X2 OR2X2_3177 ( .A(core__abc_22172_new_n8539_), .B(core__abc_22172_new_n6794_), .Y(core__abc_22172_new_n8540_));
OR2X2 OR2X2_3178 ( .A(core__abc_22172_new_n8076_), .B(core__abc_22172_new_n6814_), .Y(core__abc_22172_new_n8541_));
OR2X2 OR2X2_3179 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8544_), .Y(core__abc_22172_new_n8545_));
OR2X2 OR2X2_318 ( .A(_abc_19873_new_n1590_), .B(_abc_19873_new_n1591_), .Y(_abc_19873_new_n1592_));
OR2X2 OR2X2_3180 ( .A(core__abc_22172_new_n8545_), .B(core__abc_22172_new_n4438_), .Y(core__abc_22172_new_n8546_));
OR2X2 OR2X2_3181 ( .A(core__abc_22172_new_n8543_), .B(core__abc_22172_new_n8546_), .Y(core__abc_22172_new_n8547_));
OR2X2 OR2X2_3182 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_19_), .Y(core__abc_22172_new_n8548_));
OR2X2 OR2X2_3183 ( .A(core__abc_22172_new_n8093_), .B(core__abc_22172_new_n6787_), .Y(core__abc_22172_new_n8551_));
OR2X2 OR2X2_3184 ( .A(core__abc_22172_new_n8094_), .B(core__abc_22172_new_n6788_), .Y(core__abc_22172_new_n8552_));
OR2X2 OR2X2_3185 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8556_), .Y(core__abc_22172_new_n8557_));
OR2X2 OR2X2_3186 ( .A(core__abc_22172_new_n8557_), .B(core__abc_22172_new_n8555_), .Y(core__abc_22172_new_n8558_));
OR2X2 OR2X2_3187 ( .A(core__abc_22172_new_n8554_), .B(core__abc_22172_new_n8558_), .Y(core__abc_22172_new_n8559_));
OR2X2 OR2X2_3188 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_20_), .Y(core__abc_22172_new_n8560_));
OR2X2 OR2X2_3189 ( .A(core__abc_22172_new_n8111_), .B(core__abc_22172_new_n6781_), .Y(core__abc_22172_new_n8563_));
OR2X2 OR2X2_319 ( .A(_abc_19873_new_n1592_), .B(_abc_19873_new_n1589_), .Y(_abc_19873_new_n1593_));
OR2X2 OR2X2_3190 ( .A(core__abc_22172_new_n8110_), .B(core__abc_22172_new_n6780_), .Y(core__abc_22172_new_n8564_));
OR2X2 OR2X2_3191 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8567_), .Y(core__abc_22172_new_n8568_));
OR2X2 OR2X2_3192 ( .A(core__abc_22172_new_n8568_), .B(core__abc_22172_new_n4554_), .Y(core__abc_22172_new_n8569_));
OR2X2 OR2X2_3193 ( .A(core__abc_22172_new_n8566_), .B(core__abc_22172_new_n8569_), .Y(core__abc_22172_new_n8570_));
OR2X2 OR2X2_3194 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_21_), .Y(core__abc_22172_new_n8571_));
OR2X2 OR2X2_3195 ( .A(core__abc_22172_new_n8574_), .B(core__abc_22172_new_n6772_), .Y(core__abc_22172_new_n8575_));
OR2X2 OR2X2_3196 ( .A(core__abc_22172_new_n8127_), .B(core__abc_22172_new_n6773_), .Y(core__abc_22172_new_n8576_));
OR2X2 OR2X2_3197 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8579_), .Y(core__abc_22172_new_n8580_));
OR2X2 OR2X2_3198 ( .A(core__abc_22172_new_n8580_), .B(core__abc_22172_new_n4609_), .Y(core__abc_22172_new_n8581_));
OR2X2 OR2X2_3199 ( .A(core__abc_22172_new_n8578_), .B(core__abc_22172_new_n8581_), .Y(core__abc_22172_new_n8582_));
OR2X2 OR2X2_32 ( .A(_abc_19873_new_n982_), .B(_abc_19873_new_n983_), .Y(_abc_19873_new_n984_));
OR2X2 OR2X2_320 ( .A(_abc_19873_new_n1593_), .B(_abc_19873_new_n1588_), .Y(_abc_19873_new_n1594_));
OR2X2 OR2X2_3200 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_22_), .Y(core__abc_22172_new_n8583_));
OR2X2 OR2X2_3201 ( .A(core__abc_22172_new_n8144_), .B(core__abc_22172_new_n6758_), .Y(core__abc_22172_new_n8586_));
OR2X2 OR2X2_3202 ( .A(core__abc_22172_new_n8143_), .B(core__abc_22172_new_n6757_), .Y(core__abc_22172_new_n8587_));
OR2X2 OR2X2_3203 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8590_), .Y(core__abc_22172_new_n8591_));
OR2X2 OR2X2_3204 ( .A(core__abc_22172_new_n8591_), .B(core__abc_22172_new_n4652_), .Y(core__abc_22172_new_n8592_));
OR2X2 OR2X2_3205 ( .A(core__abc_22172_new_n8589_), .B(core__abc_22172_new_n8592_), .Y(core__abc_22172_new_n8593_));
OR2X2 OR2X2_3206 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_23_), .Y(core__abc_22172_new_n8594_));
OR2X2 OR2X2_3207 ( .A(core__abc_22172_new_n8157_), .B(core__abc_22172_new_n8597_), .Y(core__abc_22172_new_n8598_));
OR2X2 OR2X2_3208 ( .A(core__abc_22172_new_n8158_), .B(core__abc_22172_new_n6751_), .Y(core__abc_22172_new_n8599_));
OR2X2 OR2X2_3209 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8603_), .Y(core__abc_22172_new_n8604_));
OR2X2 OR2X2_321 ( .A(_abc_19873_new_n1596_), .B(_abc_19873_new_n1597_), .Y(_abc_19873_new_n1598_));
OR2X2 OR2X2_3210 ( .A(core__abc_22172_new_n8604_), .B(core__abc_22172_new_n8602_), .Y(core__abc_22172_new_n8605_));
OR2X2 OR2X2_3211 ( .A(core__abc_22172_new_n8601_), .B(core__abc_22172_new_n8605_), .Y(core__abc_22172_new_n8606_));
OR2X2 OR2X2_3212 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_24_), .Y(core__abc_22172_new_n8607_));
OR2X2 OR2X2_3213 ( .A(core__abc_22172_new_n8610_), .B(core__abc_22172_new_n6741_), .Y(core__abc_22172_new_n8611_));
OR2X2 OR2X2_3214 ( .A(core__abc_22172_new_n8174_), .B(core__abc_22172_new_n6742_), .Y(core__abc_22172_new_n8612_));
OR2X2 OR2X2_3215 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8617_), .Y(core__abc_22172_new_n8618_));
OR2X2 OR2X2_3216 ( .A(core__abc_22172_new_n8618_), .B(core__abc_22172_new_n8616_), .Y(core__abc_22172_new_n8619_));
OR2X2 OR2X2_3217 ( .A(core__abc_22172_new_n8614_), .B(core__abc_22172_new_n8619_), .Y(core__abc_22172_new_n8620_));
OR2X2 OR2X2_3218 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_25_), .Y(core__abc_22172_new_n8621_));
OR2X2 OR2X2_3219 ( .A(core__abc_22172_new_n8624_), .B(core__abc_22172_new_n6733_), .Y(core__abc_22172_new_n8625_));
OR2X2 OR2X2_322 ( .A(_abc_19873_new_n1599_), .B(_abc_19873_new_n1600_), .Y(_abc_19873_new_n1601_));
OR2X2 OR2X2_3220 ( .A(core__abc_22172_new_n8189_), .B(core__abc_22172_new_n8626_), .Y(core__abc_22172_new_n8627_));
OR2X2 OR2X2_3221 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8632_), .Y(core__abc_22172_new_n8633_));
OR2X2 OR2X2_3222 ( .A(core__abc_22172_new_n8633_), .B(core__abc_22172_new_n8631_), .Y(core__abc_22172_new_n8634_));
OR2X2 OR2X2_3223 ( .A(core__abc_22172_new_n8629_), .B(core__abc_22172_new_n8634_), .Y(core__abc_22172_new_n8635_));
OR2X2 OR2X2_3224 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_26_), .Y(core__abc_22172_new_n8636_));
OR2X2 OR2X2_3225 ( .A(core__abc_22172_new_n8639_), .B(core__abc_22172_new_n6720_), .Y(core__abc_22172_new_n8640_));
OR2X2 OR2X2_3226 ( .A(core__abc_22172_new_n8205_), .B(core__abc_22172_new_n6721_), .Y(core__abc_22172_new_n8641_));
OR2X2 OR2X2_3227 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8644_), .Y(core__abc_22172_new_n8645_));
OR2X2 OR2X2_3228 ( .A(core__abc_22172_new_n8645_), .B(core__abc_22172_new_n4862_), .Y(core__abc_22172_new_n8646_));
OR2X2 OR2X2_3229 ( .A(core__abc_22172_new_n8643_), .B(core__abc_22172_new_n8646_), .Y(core__abc_22172_new_n8647_));
OR2X2 OR2X2_323 ( .A(_abc_19873_new_n1598_), .B(_abc_19873_new_n1601_), .Y(_abc_19873_new_n1602_));
OR2X2 OR2X2_3230 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_27_), .Y(core__abc_22172_new_n8648_));
OR2X2 OR2X2_3231 ( .A(core__abc_22172_new_n8222_), .B(core__abc_22172_new_n6713_), .Y(core__abc_22172_new_n8651_));
OR2X2 OR2X2_3232 ( .A(core__abc_22172_new_n8223_), .B(core__abc_22172_new_n6712_), .Y(core__abc_22172_new_n8652_));
OR2X2 OR2X2_3233 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8656_), .Y(core__abc_22172_new_n8657_));
OR2X2 OR2X2_3234 ( .A(core__abc_22172_new_n8657_), .B(core__abc_22172_new_n8655_), .Y(core__abc_22172_new_n8658_));
OR2X2 OR2X2_3235 ( .A(core__abc_22172_new_n8654_), .B(core__abc_22172_new_n8658_), .Y(core__abc_22172_new_n8659_));
OR2X2 OR2X2_3236 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_28_), .Y(core__abc_22172_new_n8660_));
OR2X2 OR2X2_3237 ( .A(core__abc_22172_new_n8239_), .B(core__abc_22172_new_n6692_), .Y(core__abc_22172_new_n8663_));
OR2X2 OR2X2_3238 ( .A(core__abc_22172_new_n8238_), .B(core__abc_22172_new_n6691_), .Y(core__abc_22172_new_n8664_));
OR2X2 OR2X2_3239 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8667_), .Y(core__abc_22172_new_n8668_));
OR2X2 OR2X2_324 ( .A(_abc_19873_new_n1602_), .B(_abc_19873_new_n1595_), .Y(_abc_19873_new_n1603_));
OR2X2 OR2X2_3240 ( .A(core__abc_22172_new_n8668_), .B(core__abc_22172_new_n4973_), .Y(core__abc_22172_new_n8669_));
OR2X2 OR2X2_3241 ( .A(core__abc_22172_new_n8666_), .B(core__abc_22172_new_n8669_), .Y(core__abc_22172_new_n8670_));
OR2X2 OR2X2_3242 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_29_), .Y(core__abc_22172_new_n8671_));
OR2X2 OR2X2_3243 ( .A(core__abc_22172_new_n8674_), .B(core__abc_22172_new_n6683_), .Y(core__abc_22172_new_n8675_));
OR2X2 OR2X2_3244 ( .A(core__abc_22172_new_n8255_), .B(core__abc_22172_new_n6686_), .Y(core__abc_22172_new_n8676_));
OR2X2 OR2X2_3245 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8679_), .Y(core__abc_22172_new_n8680_));
OR2X2 OR2X2_3246 ( .A(core__abc_22172_new_n8680_), .B(core__abc_22172_new_n5027_), .Y(core__abc_22172_new_n8681_));
OR2X2 OR2X2_3247 ( .A(core__abc_22172_new_n8678_), .B(core__abc_22172_new_n8681_), .Y(core__abc_22172_new_n8682_));
OR2X2 OR2X2_3248 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_30_), .Y(core__abc_22172_new_n8683_));
OR2X2 OR2X2_3249 ( .A(core__abc_22172_new_n8272_), .B(core__abc_22172_new_n6674_), .Y(core__abc_22172_new_n8686_));
OR2X2 OR2X2_325 ( .A(_abc_19873_new_n1603_), .B(_abc_19873_new_n1594_), .Y(_abc_19873_new_n1604_));
OR2X2 OR2X2_3250 ( .A(core__abc_22172_new_n8271_), .B(core__abc_22172_new_n6673_), .Y(core__abc_22172_new_n8687_));
OR2X2 OR2X2_3251 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8690_), .Y(core__abc_22172_new_n8691_));
OR2X2 OR2X2_3252 ( .A(core__abc_22172_new_n8691_), .B(core__abc_22172_new_n5074_), .Y(core__abc_22172_new_n8692_));
OR2X2 OR2X2_3253 ( .A(core__abc_22172_new_n8689_), .B(core__abc_22172_new_n8692_), .Y(core__abc_22172_new_n8693_));
OR2X2 OR2X2_3254 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_31_), .Y(core__abc_22172_new_n8694_));
OR2X2 OR2X2_3255 ( .A(core__abc_22172_new_n6864_), .B(core__abc_22172_new_n6665_), .Y(core__abc_22172_new_n8697_));
OR2X2 OR2X2_3256 ( .A(core__abc_22172_new_n6865_), .B(core__abc_22172_new_n6668_), .Y(core__abc_22172_new_n8698_));
OR2X2 OR2X2_3257 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8703_), .Y(core__abc_22172_new_n8704_));
OR2X2 OR2X2_3258 ( .A(core__abc_22172_new_n8704_), .B(core__abc_22172_new_n8702_), .Y(core__abc_22172_new_n8705_));
OR2X2 OR2X2_3259 ( .A(core__abc_22172_new_n8700_), .B(core__abc_22172_new_n8705_), .Y(core__abc_22172_new_n8706_));
OR2X2 OR2X2_326 ( .A(_abc_19873_new_n1608_), .B(_abc_19873_new_n1606_), .Y(_abc_19873_new_n1609_));
OR2X2 OR2X2_3260 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_32_), .Y(core__abc_22172_new_n8707_));
OR2X2 OR2X2_3261 ( .A(core__abc_22172_new_n6901_), .B(core__abc_22172_new_n6637_), .Y(core__abc_22172_new_n8710_));
OR2X2 OR2X2_3262 ( .A(core__abc_22172_new_n6900_), .B(core__abc_22172_new_n6636_), .Y(core__abc_22172_new_n8711_));
OR2X2 OR2X2_3263 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8715_), .Y(core__abc_22172_new_n8716_));
OR2X2 OR2X2_3264 ( .A(core__abc_22172_new_n8716_), .B(core__abc_22172_new_n8714_), .Y(core__abc_22172_new_n8717_));
OR2X2 OR2X2_3265 ( .A(core__abc_22172_new_n8713_), .B(core__abc_22172_new_n8717_), .Y(core__abc_22172_new_n8718_));
OR2X2 OR2X2_3266 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_33_), .Y(core__abc_22172_new_n8719_));
OR2X2 OR2X2_3267 ( .A(core__abc_22172_new_n8722_), .B(core__abc_22172_new_n6640_), .Y(core__abc_22172_new_n8723_));
OR2X2 OR2X2_3268 ( .A(core__abc_22172_new_n6929_), .B(core__abc_22172_new_n6630_), .Y(core__abc_22172_new_n8724_));
OR2X2 OR2X2_3269 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8727_), .Y(core__abc_22172_new_n8728_));
OR2X2 OR2X2_327 ( .A(_abc_19873_new_n1612_), .B(_abc_19873_new_n1611_), .Y(_abc_19873_new_n1613_));
OR2X2 OR2X2_3270 ( .A(core__abc_22172_new_n8728_), .B(core__abc_22172_new_n5236_), .Y(core__abc_22172_new_n8729_));
OR2X2 OR2X2_3271 ( .A(core__abc_22172_new_n8726_), .B(core__abc_22172_new_n8729_), .Y(core__abc_22172_new_n8730_));
OR2X2 OR2X2_3272 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_34_), .Y(core__abc_22172_new_n8731_));
OR2X2 OR2X2_3273 ( .A(core__abc_22172_new_n8734_), .B(core__abc_22172_new_n6611_), .Y(core__abc_22172_new_n8735_));
OR2X2 OR2X2_3274 ( .A(core__abc_22172_new_n6952_), .B(core__abc_22172_new_n6612_), .Y(core__abc_22172_new_n8736_));
OR2X2 OR2X2_3275 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8739_), .Y(core__abc_22172_new_n8740_));
OR2X2 OR2X2_3276 ( .A(core__abc_22172_new_n8740_), .B(core__abc_22172_new_n5280_), .Y(core__abc_22172_new_n8741_));
OR2X2 OR2X2_3277 ( .A(core__abc_22172_new_n8738_), .B(core__abc_22172_new_n8741_), .Y(core__abc_22172_new_n8742_));
OR2X2 OR2X2_3278 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_35_), .Y(core__abc_22172_new_n8743_));
OR2X2 OR2X2_3279 ( .A(core__abc_22172_new_n6978_), .B(core__abc_22172_new_n6620_), .Y(core__abc_22172_new_n8746_));
OR2X2 OR2X2_328 ( .A(_abc_19873_new_n1616_), .B(_abc_19873_new_n1615_), .Y(_abc_19873_new_n1617_));
OR2X2 OR2X2_3280 ( .A(core__abc_22172_new_n6979_), .B(core__abc_22172_new_n6622_), .Y(core__abc_22172_new_n8747_));
OR2X2 OR2X2_3281 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8750_), .Y(core__abc_22172_new_n8751_));
OR2X2 OR2X2_3282 ( .A(core__abc_22172_new_n8751_), .B(core__abc_22172_new_n5331_), .Y(core__abc_22172_new_n8752_));
OR2X2 OR2X2_3283 ( .A(core__abc_22172_new_n8749_), .B(core__abc_22172_new_n8752_), .Y(core__abc_22172_new_n8753_));
OR2X2 OR2X2_3284 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_36_), .Y(core__abc_22172_new_n8754_));
OR2X2 OR2X2_3285 ( .A(core__abc_22172_new_n7007_), .B(core__abc_22172_new_n6601_), .Y(core__abc_22172_new_n8757_));
OR2X2 OR2X2_3286 ( .A(core__abc_22172_new_n7006_), .B(core__abc_22172_new_n6600_), .Y(core__abc_22172_new_n8758_));
OR2X2 OR2X2_3287 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8761_), .Y(core__abc_22172_new_n8762_));
OR2X2 OR2X2_3288 ( .A(core__abc_22172_new_n8762_), .B(core__abc_22172_new_n5379_), .Y(core__abc_22172_new_n8763_));
OR2X2 OR2X2_3289 ( .A(core__abc_22172_new_n8760_), .B(core__abc_22172_new_n8763_), .Y(core__abc_22172_new_n8764_));
OR2X2 OR2X2_329 ( .A(_abc_19873_new_n1620_), .B(_abc_19873_new_n1619_), .Y(_abc_19873_new_n1621_));
OR2X2 OR2X2_3290 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_37_), .Y(core__abc_22172_new_n8765_));
OR2X2 OR2X2_3291 ( .A(core__abc_22172_new_n7036_), .B(core__abc_22172_new_n6592_), .Y(core__abc_22172_new_n8768_));
OR2X2 OR2X2_3292 ( .A(core__abc_22172_new_n7037_), .B(core__abc_22172_new_n8769_), .Y(core__abc_22172_new_n8770_));
OR2X2 OR2X2_3293 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8773_), .Y(core__abc_22172_new_n8774_));
OR2X2 OR2X2_3294 ( .A(core__abc_22172_new_n8774_), .B(core__abc_22172_new_n5428_), .Y(core__abc_22172_new_n8775_));
OR2X2 OR2X2_3295 ( .A(core__abc_22172_new_n8772_), .B(core__abc_22172_new_n8775_), .Y(core__abc_22172_new_n8776_));
OR2X2 OR2X2_3296 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_38_), .Y(core__abc_22172_new_n8777_));
OR2X2 OR2X2_3297 ( .A(core__abc_22172_new_n8780_), .B(core__abc_22172_new_n6582_), .Y(core__abc_22172_new_n8781_));
OR2X2 OR2X2_3298 ( .A(core__abc_22172_new_n7062_), .B(core__abc_22172_new_n6583_), .Y(core__abc_22172_new_n8782_));
OR2X2 OR2X2_3299 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8785_), .Y(core__abc_22172_new_n8786_));
OR2X2 OR2X2_33 ( .A(_abc_19873_new_n981_), .B(_abc_19873_new_n984_), .Y(_abc_19873_new_n985_));
OR2X2 OR2X2_330 ( .A(_abc_19873_new_n1624_), .B(_abc_19873_new_n1623_), .Y(_abc_19873_new_n1625_));
OR2X2 OR2X2_3300 ( .A(core__abc_22172_new_n8786_), .B(core__abc_22172_new_n5470_), .Y(core__abc_22172_new_n8787_));
OR2X2 OR2X2_3301 ( .A(core__abc_22172_new_n8784_), .B(core__abc_22172_new_n8787_), .Y(core__abc_22172_new_n8788_));
OR2X2 OR2X2_3302 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_39_), .Y(core__abc_22172_new_n8789_));
OR2X2 OR2X2_3303 ( .A(core__abc_22172_new_n7106_), .B(core__abc_22172_new_n6575_), .Y(core__abc_22172_new_n8792_));
OR2X2 OR2X2_3304 ( .A(core__abc_22172_new_n7107_), .B(core__abc_22172_new_n6574_), .Y(core__abc_22172_new_n8793_));
OR2X2 OR2X2_3305 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8796_), .Y(core__abc_22172_new_n8797_));
OR2X2 OR2X2_3306 ( .A(core__abc_22172_new_n8797_), .B(core__abc_22172_new_n5525_), .Y(core__abc_22172_new_n8798_));
OR2X2 OR2X2_3307 ( .A(core__abc_22172_new_n8795_), .B(core__abc_22172_new_n8798_), .Y(core__abc_22172_new_n8799_));
OR2X2 OR2X2_3308 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_40_), .Y(core__abc_22172_new_n8800_));
OR2X2 OR2X2_3309 ( .A(core__abc_22172_new_n7135_), .B(core__abc_22172_new_n6538_), .Y(core__abc_22172_new_n8803_));
OR2X2 OR2X2_331 ( .A(_abc_19873_new_n1628_), .B(_abc_19873_new_n1627_), .Y(_abc_19873_new_n1629_));
OR2X2 OR2X2_3310 ( .A(core__abc_22172_new_n7134_), .B(core__abc_22172_new_n6537_), .Y(core__abc_22172_new_n8804_));
OR2X2 OR2X2_3311 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8809_), .Y(core__abc_22172_new_n8810_));
OR2X2 OR2X2_3312 ( .A(core__abc_22172_new_n8810_), .B(core__abc_22172_new_n8808_), .Y(core__abc_22172_new_n8811_));
OR2X2 OR2X2_3313 ( .A(core__abc_22172_new_n8806_), .B(core__abc_22172_new_n8811_), .Y(core__abc_22172_new_n8812_));
OR2X2 OR2X2_3314 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_41_), .Y(core__abc_22172_new_n8813_));
OR2X2 OR2X2_3315 ( .A(core__abc_22172_new_n8816_), .B(core__abc_22172_new_n6530_), .Y(core__abc_22172_new_n8817_));
OR2X2 OR2X2_3316 ( .A(core__abc_22172_new_n7164_), .B(core__abc_22172_new_n6531_), .Y(core__abc_22172_new_n8818_));
OR2X2 OR2X2_3317 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8822_), .Y(core__abc_22172_new_n8823_));
OR2X2 OR2X2_3318 ( .A(core__abc_22172_new_n8823_), .B(core__abc_22172_new_n8821_), .Y(core__abc_22172_new_n8824_));
OR2X2 OR2X2_3319 ( .A(core__abc_22172_new_n8820_), .B(core__abc_22172_new_n8824_), .Y(core__abc_22172_new_n8825_));
OR2X2 OR2X2_332 ( .A(_abc_19873_new_n1632_), .B(_abc_19873_new_n1631_), .Y(_abc_19873_new_n1633_));
OR2X2 OR2X2_3320 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_42_), .Y(core__abc_22172_new_n8826_));
OR2X2 OR2X2_3321 ( .A(core__abc_22172_new_n8829_), .B(core__abc_22172_new_n6519_), .Y(core__abc_22172_new_n8830_));
OR2X2 OR2X2_3322 ( .A(core__abc_22172_new_n7188_), .B(core__abc_22172_new_n6520_), .Y(core__abc_22172_new_n8831_));
OR2X2 OR2X2_3323 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8834_), .Y(core__abc_22172_new_n8835_));
OR2X2 OR2X2_3324 ( .A(core__abc_22172_new_n8835_), .B(core__abc_22172_new_n5649_), .Y(core__abc_22172_new_n8836_));
OR2X2 OR2X2_3325 ( .A(core__abc_22172_new_n8833_), .B(core__abc_22172_new_n8836_), .Y(core__abc_22172_new_n8837_));
OR2X2 OR2X2_3326 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_43_), .Y(core__abc_22172_new_n8838_));
OR2X2 OR2X2_3327 ( .A(core__abc_22172_new_n7219_), .B(core__abc_22172_new_n6511_), .Y(core__abc_22172_new_n8841_));
OR2X2 OR2X2_3328 ( .A(core__abc_22172_new_n7220_), .B(core__abc_22172_new_n6510_), .Y(core__abc_22172_new_n8842_));
OR2X2 OR2X2_3329 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8847_), .Y(core__abc_22172_new_n8848_));
OR2X2 OR2X2_333 ( .A(_abc_19873_new_n1636_), .B(_abc_19873_new_n1635_), .Y(_abc_19873_new_n1637_));
OR2X2 OR2X2_3330 ( .A(core__abc_22172_new_n8848_), .B(core__abc_22172_new_n8846_), .Y(core__abc_22172_new_n8849_));
OR2X2 OR2X2_3331 ( .A(core__abc_22172_new_n8844_), .B(core__abc_22172_new_n8849_), .Y(core__abc_22172_new_n8850_));
OR2X2 OR2X2_3332 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_44_), .Y(core__abc_22172_new_n8851_));
OR2X2 OR2X2_3333 ( .A(core__abc_22172_new_n8854_), .B(core__abc_22172_new_n6499_), .Y(core__abc_22172_new_n8855_));
OR2X2 OR2X2_3334 ( .A(core__abc_22172_new_n7245_), .B(core__abc_22172_new_n6500_), .Y(core__abc_22172_new_n8856_));
OR2X2 OR2X2_3335 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8859_), .Y(core__abc_22172_new_n8860_));
OR2X2 OR2X2_3336 ( .A(core__abc_22172_new_n8860_), .B(core__abc_22172_new_n5732_), .Y(core__abc_22172_new_n8861_));
OR2X2 OR2X2_3337 ( .A(core__abc_22172_new_n8858_), .B(core__abc_22172_new_n8861_), .Y(core__abc_22172_new_n8862_));
OR2X2 OR2X2_3338 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_45_), .Y(core__abc_22172_new_n8863_));
OR2X2 OR2X2_3339 ( .A(core__abc_22172_new_n7277_), .B(core__abc_22172_new_n6489_), .Y(core__abc_22172_new_n8866_));
OR2X2 OR2X2_334 ( .A(_abc_19873_new_n1640_), .B(_abc_19873_new_n1639_), .Y(_abc_19873_new_n1641_));
OR2X2 OR2X2_3340 ( .A(core__abc_22172_new_n7278_), .B(core__abc_22172_new_n6490_), .Y(core__abc_22172_new_n8867_));
OR2X2 OR2X2_3341 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8870_), .Y(core__abc_22172_new_n8871_));
OR2X2 OR2X2_3342 ( .A(core__abc_22172_new_n8871_), .B(core__abc_22172_new_n5774_), .Y(core__abc_22172_new_n8872_));
OR2X2 OR2X2_3343 ( .A(core__abc_22172_new_n8869_), .B(core__abc_22172_new_n8872_), .Y(core__abc_22172_new_n8873_));
OR2X2 OR2X2_3344 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_46_), .Y(core__abc_22172_new_n8874_));
OR2X2 OR2X2_3345 ( .A(core__abc_22172_new_n7306_), .B(core__abc_22172_new_n6481_), .Y(core__abc_22172_new_n8877_));
OR2X2 OR2X2_3346 ( .A(core__abc_22172_new_n7305_), .B(core__abc_22172_new_n6479_), .Y(core__abc_22172_new_n8878_));
OR2X2 OR2X2_3347 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8881_), .Y(core__abc_22172_new_n8882_));
OR2X2 OR2X2_3348 ( .A(core__abc_22172_new_n8882_), .B(core__abc_22172_new_n5812_), .Y(core__abc_22172_new_n8883_));
OR2X2 OR2X2_3349 ( .A(core__abc_22172_new_n8880_), .B(core__abc_22172_new_n8883_), .Y(core__abc_22172_new_n8884_));
OR2X2 OR2X2_335 ( .A(_abc_19873_new_n1644_), .B(_abc_19873_new_n1643_), .Y(_abc_19873_new_n1645_));
OR2X2 OR2X2_3350 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_47_), .Y(core__abc_22172_new_n8885_));
OR2X2 OR2X2_3351 ( .A(core__abc_22172_new_n7349_), .B(core__abc_22172_new_n6471_), .Y(core__abc_22172_new_n8888_));
OR2X2 OR2X2_3352 ( .A(core__abc_22172_new_n7350_), .B(core__abc_22172_new_n8889_), .Y(core__abc_22172_new_n8890_));
OR2X2 OR2X2_3353 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8893_), .Y(core__abc_22172_new_n8894_));
OR2X2 OR2X2_3354 ( .A(core__abc_22172_new_n8894_), .B(core__abc_22172_new_n5863_), .Y(core__abc_22172_new_n8895_));
OR2X2 OR2X2_3355 ( .A(core__abc_22172_new_n8892_), .B(core__abc_22172_new_n8895_), .Y(core__abc_22172_new_n8896_));
OR2X2 OR2X2_3356 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_48_), .Y(core__abc_22172_new_n8897_));
OR2X2 OR2X2_3357 ( .A(core__abc_22172_new_n7380_), .B(core__abc_22172_new_n6856_), .Y(core__abc_22172_new_n8900_));
OR2X2 OR2X2_3358 ( .A(core__abc_22172_new_n7379_), .B(core__abc_22172_new_n6855_), .Y(core__abc_22172_new_n8901_));
OR2X2 OR2X2_3359 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8906_), .Y(core__abc_22172_new_n8907_));
OR2X2 OR2X2_336 ( .A(_abc_19873_new_n1648_), .B(_abc_19873_new_n1647_), .Y(_abc_19873_new_n1649_));
OR2X2 OR2X2_3360 ( .A(core__abc_22172_new_n8907_), .B(core__abc_22172_new_n8905_), .Y(core__abc_22172_new_n8908_));
OR2X2 OR2X2_3361 ( .A(core__abc_22172_new_n8903_), .B(core__abc_22172_new_n8908_), .Y(core__abc_22172_new_n8909_));
OR2X2 OR2X2_3362 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_49_), .Y(core__abc_22172_new_n8910_));
OR2X2 OR2X2_3363 ( .A(core__abc_22172_new_n7405_), .B(core__abc_22172_new_n6891_), .Y(core__abc_22172_new_n8913_));
OR2X2 OR2X2_3364 ( .A(core__abc_22172_new_n7406_), .B(core__abc_22172_new_n6889_), .Y(core__abc_22172_new_n8914_));
OR2X2 OR2X2_3365 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8917_), .Y(core__abc_22172_new_n8918_));
OR2X2 OR2X2_3366 ( .A(core__abc_22172_new_n8918_), .B(core__abc_22172_new_n5936_), .Y(core__abc_22172_new_n8919_));
OR2X2 OR2X2_3367 ( .A(core__abc_22172_new_n8916_), .B(core__abc_22172_new_n8919_), .Y(core__abc_22172_new_n8920_));
OR2X2 OR2X2_3368 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_50_), .Y(core__abc_22172_new_n8921_));
OR2X2 OR2X2_3369 ( .A(core__abc_22172_new_n8924_), .B(core__abc_22172_new_n6920_), .Y(core__abc_22172_new_n8925_));
OR2X2 OR2X2_337 ( .A(_abc_19873_new_n1652_), .B(_abc_19873_new_n1651_), .Y(_abc_19873_new_n1653_));
OR2X2 OR2X2_3370 ( .A(core__abc_22172_new_n7433_), .B(core__abc_22172_new_n6922_), .Y(core__abc_22172_new_n8926_));
OR2X2 OR2X2_3371 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8931_), .Y(core__abc_22172_new_n8932_));
OR2X2 OR2X2_3372 ( .A(core__abc_22172_new_n8932_), .B(core__abc_22172_new_n8930_), .Y(core__abc_22172_new_n8933_));
OR2X2 OR2X2_3373 ( .A(core__abc_22172_new_n8928_), .B(core__abc_22172_new_n8933_), .Y(core__abc_22172_new_n8934_));
OR2X2 OR2X2_3374 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_51_), .Y(core__abc_22172_new_n8935_));
OR2X2 OR2X2_3375 ( .A(core__abc_22172_new_n7467_), .B(core__abc_22172_new_n6946_), .Y(core__abc_22172_new_n8938_));
OR2X2 OR2X2_3376 ( .A(core__abc_22172_new_n7468_), .B(core__abc_22172_new_n6944_), .Y(core__abc_22172_new_n8939_));
OR2X2 OR2X2_3377 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8942_), .Y(core__abc_22172_new_n8943_));
OR2X2 OR2X2_3378 ( .A(core__abc_22172_new_n8943_), .B(core__abc_22172_new_n6016_), .Y(core__abc_22172_new_n8944_));
OR2X2 OR2X2_3379 ( .A(core__abc_22172_new_n8941_), .B(core__abc_22172_new_n8944_), .Y(core__abc_22172_new_n8945_));
OR2X2 OR2X2_338 ( .A(_abc_19873_new_n1656_), .B(_abc_19873_new_n1655_), .Y(_abc_19873_new_n1657_));
OR2X2 OR2X2_3380 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_52_), .Y(core__abc_22172_new_n8946_));
OR2X2 OR2X2_3381 ( .A(core__abc_22172_new_n8949_), .B(core__abc_22172_new_n6965_), .Y(core__abc_22172_new_n8950_));
OR2X2 OR2X2_3382 ( .A(core__abc_22172_new_n7495_), .B(core__abc_22172_new_n6967_), .Y(core__abc_22172_new_n8951_));
OR2X2 OR2X2_3383 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8954_), .Y(core__abc_22172_new_n8955_));
OR2X2 OR2X2_3384 ( .A(core__abc_22172_new_n8955_), .B(core__abc_22172_new_n6049_), .Y(core__abc_22172_new_n8956_));
OR2X2 OR2X2_3385 ( .A(core__abc_22172_new_n8953_), .B(core__abc_22172_new_n8956_), .Y(core__abc_22172_new_n8957_));
OR2X2 OR2X2_3386 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_53_), .Y(core__abc_22172_new_n8958_));
OR2X2 OR2X2_3387 ( .A(core__abc_22172_new_n7523_), .B(core__abc_22172_new_n6997_), .Y(core__abc_22172_new_n8961_));
OR2X2 OR2X2_3388 ( .A(core__abc_22172_new_n7524_), .B(core__abc_22172_new_n8962_), .Y(core__abc_22172_new_n8963_));
OR2X2 OR2X2_3389 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8966_), .Y(core__abc_22172_new_n8967_));
OR2X2 OR2X2_339 ( .A(_abc_19873_new_n1660_), .B(_abc_19873_new_n1659_), .Y(_abc_19873_new_n1661_));
OR2X2 OR2X2_3390 ( .A(core__abc_22172_new_n8967_), .B(core__abc_22172_new_n6091_), .Y(core__abc_22172_new_n8968_));
OR2X2 OR2X2_3391 ( .A(core__abc_22172_new_n8965_), .B(core__abc_22172_new_n8968_), .Y(core__abc_22172_new_n8969_));
OR2X2 OR2X2_3392 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_54_), .Y(core__abc_22172_new_n8970_));
OR2X2 OR2X2_3393 ( .A(core__abc_22172_new_n7553_), .B(core__abc_22172_new_n7023_), .Y(core__abc_22172_new_n8973_));
OR2X2 OR2X2_3394 ( .A(core__abc_22172_new_n7552_), .B(core__abc_22172_new_n7021_), .Y(core__abc_22172_new_n8974_));
OR2X2 OR2X2_3395 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8977_), .Y(core__abc_22172_new_n8978_));
OR2X2 OR2X2_3396 ( .A(core__abc_22172_new_n8978_), .B(core__abc_22172_new_n6129_), .Y(core__abc_22172_new_n8979_));
OR2X2 OR2X2_3397 ( .A(core__abc_22172_new_n8976_), .B(core__abc_22172_new_n8979_), .Y(core__abc_22172_new_n8980_));
OR2X2 OR2X2_3398 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_55_), .Y(core__abc_22172_new_n8981_));
OR2X2 OR2X2_3399 ( .A(core__abc_22172_new_n7590_), .B(core__abc_22172_new_n7054_), .Y(core__abc_22172_new_n8984_));
OR2X2 OR2X2_34 ( .A(_abc_19873_new_n985_), .B(_abc_19873_new_n978_), .Y(_abc_19873_new_n986_));
OR2X2 OR2X2_340 ( .A(_abc_19873_new_n1664_), .B(_abc_19873_new_n1663_), .Y(_abc_19873_new_n1665_));
OR2X2 OR2X2_3400 ( .A(core__abc_22172_new_n7591_), .B(core__abc_22172_new_n7055_), .Y(core__abc_22172_new_n8985_));
OR2X2 OR2X2_3401 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n8988_), .Y(core__abc_22172_new_n8989_));
OR2X2 OR2X2_3402 ( .A(core__abc_22172_new_n8989_), .B(core__abc_22172_new_n6182_), .Y(core__abc_22172_new_n8990_));
OR2X2 OR2X2_3403 ( .A(core__abc_22172_new_n8987_), .B(core__abc_22172_new_n8990_), .Y(core__abc_22172_new_n8991_));
OR2X2 OR2X2_3404 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_56_), .Y(core__abc_22172_new_n8992_));
OR2X2 OR2X2_3405 ( .A(core__abc_22172_new_n8995_), .B(core__abc_22172_new_n7097_), .Y(core__abc_22172_new_n8996_));
OR2X2 OR2X2_3406 ( .A(core__abc_22172_new_n7616_), .B(core__abc_22172_new_n7099_), .Y(core__abc_22172_new_n8997_));
OR2X2 OR2X2_3407 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n9000_), .Y(core__abc_22172_new_n9001_));
OR2X2 OR2X2_3408 ( .A(core__abc_22172_new_n9001_), .B(core__abc_22172_new_n6214_), .Y(core__abc_22172_new_n9002_));
OR2X2 OR2X2_3409 ( .A(core__abc_22172_new_n8999_), .B(core__abc_22172_new_n9002_), .Y(core__abc_22172_new_n9003_));
OR2X2 OR2X2_341 ( .A(_abc_19873_new_n1668_), .B(_abc_19873_new_n1667_), .Y(_abc_19873_new_n1669_));
OR2X2 OR2X2_3410 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_57_), .Y(core__abc_22172_new_n9004_));
OR2X2 OR2X2_3411 ( .A(core__abc_22172_new_n9007_), .B(core__abc_22172_new_n7122_), .Y(core__abc_22172_new_n9008_));
OR2X2 OR2X2_3412 ( .A(core__abc_22172_new_n7646_), .B(core__abc_22172_new_n9009_), .Y(core__abc_22172_new_n9010_));
OR2X2 OR2X2_3413 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n9013_), .Y(core__abc_22172_new_n9014_));
OR2X2 OR2X2_3414 ( .A(core__abc_22172_new_n9014_), .B(core__abc_22172_new_n6257_), .Y(core__abc_22172_new_n9015_));
OR2X2 OR2X2_3415 ( .A(core__abc_22172_new_n9012_), .B(core__abc_22172_new_n9015_), .Y(core__abc_22172_new_n9016_));
OR2X2 OR2X2_3416 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_58_), .Y(core__abc_22172_new_n9017_));
OR2X2 OR2X2_3417 ( .A(core__abc_22172_new_n9020_), .B(core__abc_22172_new_n7155_), .Y(core__abc_22172_new_n9021_));
OR2X2 OR2X2_3418 ( .A(core__abc_22172_new_n7671_), .B(core__abc_22172_new_n7156_), .Y(core__abc_22172_new_n9022_));
OR2X2 OR2X2_3419 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n9025_), .Y(core__abc_22172_new_n9026_));
OR2X2 OR2X2_342 ( .A(_abc_19873_new_n1672_), .B(_abc_19873_new_n1671_), .Y(_abc_19873_new_n1673_));
OR2X2 OR2X2_3420 ( .A(core__abc_22172_new_n9026_), .B(core__abc_22172_new_n6291_), .Y(core__abc_22172_new_n9027_));
OR2X2 OR2X2_3421 ( .A(core__abc_22172_new_n9024_), .B(core__abc_22172_new_n9027_), .Y(core__abc_22172_new_n9028_));
OR2X2 OR2X2_3422 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_59_), .Y(core__abc_22172_new_n9029_));
OR2X2 OR2X2_3423 ( .A(core__abc_22172_new_n7702_), .B(core__abc_22172_new_n7179_), .Y(core__abc_22172_new_n9032_));
OR2X2 OR2X2_3424 ( .A(core__abc_22172_new_n7703_), .B(core__abc_22172_new_n9033_), .Y(core__abc_22172_new_n9034_));
OR2X2 OR2X2_3425 ( .A(core__abc_22172_new_n9037_), .B(core__abc_22172_new_n9038_), .Y(core__abc_22172_new_n9039_));
OR2X2 OR2X2_3426 ( .A(core__abc_22172_new_n9039_), .B(core__abc_22172_new_n8283_), .Y(core__abc_22172_new_n9040_));
OR2X2 OR2X2_3427 ( .A(core__abc_22172_new_n9036_), .B(core__abc_22172_new_n9040_), .Y(core__abc_22172_new_n9041_));
OR2X2 OR2X2_3428 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_60_), .Y(core__abc_22172_new_n9042_));
OR2X2 OR2X2_3429 ( .A(core__abc_22172_new_n7727_), .B(core__abc_22172_new_n7211_), .Y(core__abc_22172_new_n9045_));
OR2X2 OR2X2_343 ( .A(_abc_19873_new_n1676_), .B(_abc_19873_new_n1675_), .Y(_abc_19873_new_n1677_));
OR2X2 OR2X2_3430 ( .A(core__abc_22172_new_n7726_), .B(core__abc_22172_new_n7210_), .Y(core__abc_22172_new_n9046_));
OR2X2 OR2X2_3431 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n9049_), .Y(core__abc_22172_new_n9050_));
OR2X2 OR2X2_3432 ( .A(core__abc_22172_new_n9050_), .B(core__abc_22172_new_n6379_), .Y(core__abc_22172_new_n9051_));
OR2X2 OR2X2_3433 ( .A(core__abc_22172_new_n9048_), .B(core__abc_22172_new_n9051_), .Y(core__abc_22172_new_n9052_));
OR2X2 OR2X2_3434 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_61_), .Y(core__abc_22172_new_n9053_));
OR2X2 OR2X2_3435 ( .A(core__abc_22172_new_n7755_), .B(core__abc_22172_new_n7236_), .Y(core__abc_22172_new_n9056_));
OR2X2 OR2X2_3436 ( .A(core__abc_22172_new_n7756_), .B(core__abc_22172_new_n7237_), .Y(core__abc_22172_new_n9057_));
OR2X2 OR2X2_3437 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n9060_), .Y(core__abc_22172_new_n9061_));
OR2X2 OR2X2_3438 ( .A(core__abc_22172_new_n9061_), .B(core__abc_22172_new_n6422_), .Y(core__abc_22172_new_n9062_));
OR2X2 OR2X2_3439 ( .A(core__abc_22172_new_n9059_), .B(core__abc_22172_new_n9062_), .Y(core__abc_22172_new_n9063_));
OR2X2 OR2X2_344 ( .A(_abc_19873_new_n1680_), .B(_abc_19873_new_n1679_), .Y(_abc_19873_new_n1681_));
OR2X2 OR2X2_3440 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_62_), .Y(core__abc_22172_new_n9064_));
OR2X2 OR2X2_3441 ( .A(core__abc_22172_new_n9067_), .B(core__abc_22172_new_n7269_), .Y(core__abc_22172_new_n9068_));
OR2X2 OR2X2_3442 ( .A(core__abc_22172_new_n7780_), .B(core__abc_22172_new_n7271_), .Y(core__abc_22172_new_n9069_));
OR2X2 OR2X2_3443 ( .A(core__abc_22172_new_n8283_), .B(core__abc_22172_new_n9072_), .Y(core__abc_22172_new_n9073_));
OR2X2 OR2X2_3444 ( .A(core__abc_22172_new_n9073_), .B(core__abc_22172_new_n6456_), .Y(core__abc_22172_new_n9074_));
OR2X2 OR2X2_3445 ( .A(core__abc_22172_new_n9071_), .B(core__abc_22172_new_n9074_), .Y(core__abc_22172_new_n9075_));
OR2X2 OR2X2_3446 ( .A(core__abc_22172_new_n8282_), .B(core_v1_reg_63_), .Y(core__abc_22172_new_n9076_));
OR2X2 OR2X2_3447 ( .A(core__abc_22172_new_n9082_), .B(core__abc_22172_new_n3212_), .Y(core__abc_22172_new_n9083_));
OR2X2 OR2X2_3448 ( .A(core_v0_reg_0_), .B(core_mi_reg_0_), .Y(core__abc_22172_new_n9086_));
OR2X2 OR2X2_3449 ( .A(core__abc_22172_new_n6868_), .B(core__abc_22172_new_n9090_), .Y(core__abc_22172_new_n9091_));
OR2X2 OR2X2_345 ( .A(_abc_19873_new_n1684_), .B(_abc_19873_new_n1683_), .Y(_abc_19873_new_n1685_));
OR2X2 OR2X2_3450 ( .A(core__abc_22172_new_n9085_), .B(core__abc_22172_new_n9091_), .Y(core__abc_22172_new_n9092_));
OR2X2 OR2X2_3451 ( .A(core__abc_22172_new_n9093_), .B(core__abc_22172_new_n9084_), .Y(core__abc_22172_new_n9094_));
OR2X2 OR2X2_3452 ( .A(core_v0_reg_1_), .B(core_mi_reg_1_), .Y(core__abc_22172_new_n9097_));
OR2X2 OR2X2_3453 ( .A(core__abc_22172_new_n6903_), .B(core__abc_22172_new_n9101_), .Y(core__abc_22172_new_n9102_));
OR2X2 OR2X2_3454 ( .A(core__abc_22172_new_n9096_), .B(core__abc_22172_new_n9102_), .Y(core__abc_22172_new_n9103_));
OR2X2 OR2X2_3455 ( .A(core__abc_22172_new_n9104_), .B(core__abc_22172_new_n9105_), .Y(core__abc_22172_new_n9106_));
OR2X2 OR2X2_3456 ( .A(core_v0_reg_2_), .B(core_mi_reg_2_), .Y(core__abc_22172_new_n9111_));
OR2X2 OR2X2_3457 ( .A(core__abc_22172_new_n9110_), .B(core__abc_22172_new_n9115_), .Y(core__abc_22172_new_n9116_));
OR2X2 OR2X2_3458 ( .A(core__abc_22172_new_n9108_), .B(core__abc_22172_new_n9116_), .Y(core__abc_22172_new_n9117_));
OR2X2 OR2X2_3459 ( .A(core__abc_22172_new_n9118_), .B(core__abc_22172_new_n9119_), .Y(core__abc_22172_new_n9120_));
OR2X2 OR2X2_346 ( .A(_abc_19873_new_n1688_), .B(_abc_19873_new_n1687_), .Y(_abc_19873_new_n1689_));
OR2X2 OR2X2_3460 ( .A(core_v0_reg_3_), .B(core_mi_reg_3_), .Y(core__abc_22172_new_n9124_));
OR2X2 OR2X2_3461 ( .A(core__abc_22172_new_n6954_), .B(core__abc_22172_new_n9128_), .Y(core__abc_22172_new_n9129_));
OR2X2 OR2X2_3462 ( .A(core__abc_22172_new_n9123_), .B(core__abc_22172_new_n9129_), .Y(core__abc_22172_new_n9130_));
OR2X2 OR2X2_3463 ( .A(core__abc_22172_new_n9131_), .B(core__abc_22172_new_n9122_), .Y(core__abc_22172_new_n9132_));
OR2X2 OR2X2_3464 ( .A(core_v0_reg_4_), .B(core_mi_reg_4_), .Y(core__abc_22172_new_n9137_));
OR2X2 OR2X2_3465 ( .A(core__abc_22172_new_n9136_), .B(core__abc_22172_new_n9141_), .Y(core__abc_22172_new_n9142_));
OR2X2 OR2X2_3466 ( .A(core__abc_22172_new_n9134_), .B(core__abc_22172_new_n9142_), .Y(core__abc_22172_new_n9143_));
OR2X2 OR2X2_3467 ( .A(core__abc_22172_new_n9144_), .B(core__abc_22172_new_n9145_), .Y(core__abc_22172_new_n9146_));
OR2X2 OR2X2_3468 ( .A(core_v0_reg_5_), .B(core_mi_reg_5_), .Y(core__abc_22172_new_n9149_));
OR2X2 OR2X2_3469 ( .A(core__abc_22172_new_n7010_), .B(core__abc_22172_new_n9153_), .Y(core__abc_22172_new_n9154_));
OR2X2 OR2X2_347 ( .A(_abc_19873_new_n1692_), .B(_abc_19873_new_n1691_), .Y(_abc_19873_new_n1693_));
OR2X2 OR2X2_3470 ( .A(core__abc_22172_new_n9148_), .B(core__abc_22172_new_n9154_), .Y(core__abc_22172_new_n9155_));
OR2X2 OR2X2_3471 ( .A(core__abc_22172_new_n9156_), .B(core__abc_22172_new_n9157_), .Y(core__abc_22172_new_n9158_));
OR2X2 OR2X2_3472 ( .A(core_v0_reg_6_), .B(core_mi_reg_6_), .Y(core__abc_22172_new_n9161_));
OR2X2 OR2X2_3473 ( .A(core__abc_22172_new_n7040_), .B(core__abc_22172_new_n9165_), .Y(core__abc_22172_new_n9166_));
OR2X2 OR2X2_3474 ( .A(core__abc_22172_new_n9160_), .B(core__abc_22172_new_n9166_), .Y(core__abc_22172_new_n9167_));
OR2X2 OR2X2_3475 ( .A(core__abc_22172_new_n9168_), .B(core__abc_22172_new_n9169_), .Y(core__abc_22172_new_n9170_));
OR2X2 OR2X2_3476 ( .A(core_v0_reg_7_), .B(core_mi_reg_7_), .Y(core__abc_22172_new_n9173_));
OR2X2 OR2X2_3477 ( .A(core__abc_22172_new_n7064_), .B(core__abc_22172_new_n9177_), .Y(core__abc_22172_new_n9178_));
OR2X2 OR2X2_3478 ( .A(core__abc_22172_new_n9172_), .B(core__abc_22172_new_n9178_), .Y(core__abc_22172_new_n9179_));
OR2X2 OR2X2_3479 ( .A(core__abc_22172_new_n9180_), .B(core__abc_22172_new_n9181_), .Y(core__abc_22172_new_n9182_));
OR2X2 OR2X2_348 ( .A(_abc_19873_new_n1696_), .B(_abc_19873_new_n1695_), .Y(_abc_19873_new_n1697_));
OR2X2 OR2X2_3480 ( .A(core_v0_reg_8_), .B(core_mi_reg_8_), .Y(core__abc_22172_new_n9187_));
OR2X2 OR2X2_3481 ( .A(core__abc_22172_new_n9186_), .B(core__abc_22172_new_n9191_), .Y(core__abc_22172_new_n9192_));
OR2X2 OR2X2_3482 ( .A(core__abc_22172_new_n9184_), .B(core__abc_22172_new_n9192_), .Y(core__abc_22172_new_n9193_));
OR2X2 OR2X2_3483 ( .A(core__abc_22172_new_n9194_), .B(core__abc_22172_new_n9195_), .Y(core__abc_22172_new_n9196_));
OR2X2 OR2X2_3484 ( .A(core_v0_reg_9_), .B(core_mi_reg_9_), .Y(core__abc_22172_new_n9200_));
OR2X2 OR2X2_3485 ( .A(core__abc_22172_new_n9199_), .B(core__abc_22172_new_n9204_), .Y(core__abc_22172_new_n9205_));
OR2X2 OR2X2_3486 ( .A(core__abc_22172_new_n9198_), .B(core__abc_22172_new_n9205_), .Y(core__abc_22172_new_n9206_));
OR2X2 OR2X2_3487 ( .A(core__abc_22172_new_n9207_), .B(core__abc_22172_new_n9208_), .Y(core__abc_22172_new_n9209_));
OR2X2 OR2X2_3488 ( .A(core_v0_reg_10_), .B(core_mi_reg_10_), .Y(core__abc_22172_new_n9214_));
OR2X2 OR2X2_3489 ( .A(core__abc_22172_new_n9213_), .B(core__abc_22172_new_n9218_), .Y(core__abc_22172_new_n9219_));
OR2X2 OR2X2_349 ( .A(_abc_19873_new_n1700_), .B(_abc_19873_new_n1699_), .Y(_abc_19873_new_n1701_));
OR2X2 OR2X2_3490 ( .A(core__abc_22172_new_n9211_), .B(core__abc_22172_new_n9219_), .Y(core__abc_22172_new_n9220_));
OR2X2 OR2X2_3491 ( .A(core__abc_22172_new_n9221_), .B(core__abc_22172_new_n9222_), .Y(core__abc_22172_new_n9223_));
OR2X2 OR2X2_3492 ( .A(core_v0_reg_11_), .B(core_mi_reg_11_), .Y(core__abc_22172_new_n9226_));
OR2X2 OR2X2_3493 ( .A(core__abc_22172_new_n7190_), .B(core__abc_22172_new_n9230_), .Y(core__abc_22172_new_n9231_));
OR2X2 OR2X2_3494 ( .A(core__abc_22172_new_n9225_), .B(core__abc_22172_new_n9231_), .Y(core__abc_22172_new_n9232_));
OR2X2 OR2X2_3495 ( .A(core__abc_22172_new_n9233_), .B(core__abc_22172_new_n9234_), .Y(core__abc_22172_new_n9235_));
OR2X2 OR2X2_3496 ( .A(core_v0_reg_12_), .B(core_mi_reg_12_), .Y(core__abc_22172_new_n9239_));
OR2X2 OR2X2_3497 ( .A(core__abc_22172_new_n9238_), .B(core__abc_22172_new_n9243_), .Y(core__abc_22172_new_n9244_));
OR2X2 OR2X2_3498 ( .A(core__abc_22172_new_n9237_), .B(core__abc_22172_new_n9244_), .Y(core__abc_22172_new_n9245_));
OR2X2 OR2X2_3499 ( .A(core__abc_22172_new_n9246_), .B(core__abc_22172_new_n9247_), .Y(core__abc_22172_new_n9248_));
OR2X2 OR2X2_35 ( .A(_abc_19873_new_n973_), .B(_abc_19873_new_n986_), .Y(_abc_19873_new_n987_));
OR2X2 OR2X2_350 ( .A(_abc_19873_new_n1704_), .B(_abc_19873_new_n1703_), .Y(_abc_19873_new_n1705_));
OR2X2 OR2X2_3500 ( .A(core_v0_reg_13_), .B(core_mi_reg_13_), .Y(core__abc_22172_new_n9251_));
OR2X2 OR2X2_3501 ( .A(core__abc_22172_new_n7248_), .B(core__abc_22172_new_n9255_), .Y(core__abc_22172_new_n9256_));
OR2X2 OR2X2_3502 ( .A(core__abc_22172_new_n9250_), .B(core__abc_22172_new_n9256_), .Y(core__abc_22172_new_n9257_));
OR2X2 OR2X2_3503 ( .A(core__abc_22172_new_n9258_), .B(core__abc_22172_new_n9259_), .Y(core__abc_22172_new_n9260_));
OR2X2 OR2X2_3504 ( .A(core_v0_reg_14_), .B(core_mi_reg_14_), .Y(core__abc_22172_new_n9263_));
OR2X2 OR2X2_3505 ( .A(core__abc_22172_new_n7281_), .B(core__abc_22172_new_n9267_), .Y(core__abc_22172_new_n9268_));
OR2X2 OR2X2_3506 ( .A(core__abc_22172_new_n9262_), .B(core__abc_22172_new_n9268_), .Y(core__abc_22172_new_n9269_));
OR2X2 OR2X2_3507 ( .A(core__abc_22172_new_n9270_), .B(core__abc_22172_new_n9271_), .Y(core__abc_22172_new_n9272_));
OR2X2 OR2X2_3508 ( .A(core_v0_reg_15_), .B(core_mi_reg_15_), .Y(core__abc_22172_new_n9275_));
OR2X2 OR2X2_3509 ( .A(core__abc_22172_new_n7308_), .B(core__abc_22172_new_n9279_), .Y(core__abc_22172_new_n9280_));
OR2X2 OR2X2_351 ( .A(_abc_19873_new_n1708_), .B(_abc_19873_new_n1707_), .Y(_abc_19873_new_n1709_));
OR2X2 OR2X2_3510 ( .A(core__abc_22172_new_n9274_), .B(core__abc_22172_new_n9280_), .Y(core__abc_22172_new_n9281_));
OR2X2 OR2X2_3511 ( .A(core__abc_22172_new_n9282_), .B(core__abc_22172_new_n9283_), .Y(core__abc_22172_new_n9284_));
OR2X2 OR2X2_3512 ( .A(core_v0_reg_16_), .B(core_mi_reg_16_), .Y(core__abc_22172_new_n9287_));
OR2X2 OR2X2_3513 ( .A(core__abc_22172_new_n7353_), .B(core__abc_22172_new_n9291_), .Y(core__abc_22172_new_n9292_));
OR2X2 OR2X2_3514 ( .A(core__abc_22172_new_n9286_), .B(core__abc_22172_new_n9292_), .Y(core__abc_22172_new_n9293_));
OR2X2 OR2X2_3515 ( .A(core__abc_22172_new_n9294_), .B(core__abc_22172_new_n9295_), .Y(core__abc_22172_new_n9296_));
OR2X2 OR2X2_3516 ( .A(core_v0_reg_17_), .B(core_mi_reg_17_), .Y(core__abc_22172_new_n9301_));
OR2X2 OR2X2_3517 ( .A(core__abc_22172_new_n9300_), .B(core__abc_22172_new_n9305_), .Y(core__abc_22172_new_n9306_));
OR2X2 OR2X2_3518 ( .A(core__abc_22172_new_n9298_), .B(core__abc_22172_new_n9306_), .Y(core__abc_22172_new_n9307_));
OR2X2 OR2X2_3519 ( .A(core__abc_22172_new_n9308_), .B(core__abc_22172_new_n9309_), .Y(core__abc_22172_new_n9310_));
OR2X2 OR2X2_352 ( .A(_abc_19873_new_n1712_), .B(_abc_19873_new_n1711_), .Y(_abc_19873_new_n1713_));
OR2X2 OR2X2_3520 ( .A(core_v0_reg_18_), .B(core_mi_reg_18_), .Y(core__abc_22172_new_n9314_));
OR2X2 OR2X2_3521 ( .A(core__abc_22172_new_n9313_), .B(core__abc_22172_new_n9318_), .Y(core__abc_22172_new_n9319_));
OR2X2 OR2X2_3522 ( .A(core__abc_22172_new_n9312_), .B(core__abc_22172_new_n9319_), .Y(core__abc_22172_new_n9320_));
OR2X2 OR2X2_3523 ( .A(core__abc_22172_new_n9321_), .B(core__abc_22172_new_n9322_), .Y(core__abc_22172_new_n9323_));
OR2X2 OR2X2_3524 ( .A(core_v0_reg_19_), .B(core_mi_reg_19_), .Y(core__abc_22172_new_n9326_));
OR2X2 OR2X2_3525 ( .A(core__abc_22172_new_n7435_), .B(core__abc_22172_new_n9330_), .Y(core__abc_22172_new_n9331_));
OR2X2 OR2X2_3526 ( .A(core__abc_22172_new_n9325_), .B(core__abc_22172_new_n9331_), .Y(core__abc_22172_new_n9332_));
OR2X2 OR2X2_3527 ( .A(core__abc_22172_new_n9333_), .B(core__abc_22172_new_n9334_), .Y(core__abc_22172_new_n9335_));
OR2X2 OR2X2_3528 ( .A(core_v0_reg_20_), .B(core_mi_reg_20_), .Y(core__abc_22172_new_n9340_));
OR2X2 OR2X2_3529 ( .A(core__abc_22172_new_n9339_), .B(core__abc_22172_new_n9344_), .Y(core__abc_22172_new_n9345_));
OR2X2 OR2X2_353 ( .A(_abc_19873_new_n1716_), .B(_abc_19873_new_n1715_), .Y(_abc_19873_new_n1717_));
OR2X2 OR2X2_3530 ( .A(core__abc_22172_new_n9337_), .B(core__abc_22172_new_n9345_), .Y(core__abc_22172_new_n9346_));
OR2X2 OR2X2_3531 ( .A(core__abc_22172_new_n9347_), .B(core__abc_22172_new_n9348_), .Y(core__abc_22172_new_n9349_));
OR2X2 OR2X2_3532 ( .A(core_v0_reg_21_), .B(core_mi_reg_21_), .Y(core__abc_22172_new_n9352_));
OR2X2 OR2X2_3533 ( .A(core__abc_22172_new_n7498_), .B(core__abc_22172_new_n9356_), .Y(core__abc_22172_new_n9357_));
OR2X2 OR2X2_3534 ( .A(core__abc_22172_new_n9351_), .B(core__abc_22172_new_n9357_), .Y(core__abc_22172_new_n9358_));
OR2X2 OR2X2_3535 ( .A(core__abc_22172_new_n9359_), .B(core__abc_22172_new_n9360_), .Y(core__abc_22172_new_n9361_));
OR2X2 OR2X2_3536 ( .A(core_v0_reg_22_), .B(core_mi_reg_22_), .Y(core__abc_22172_new_n9364_));
OR2X2 OR2X2_3537 ( .A(core__abc_22172_new_n7527_), .B(core__abc_22172_new_n9368_), .Y(core__abc_22172_new_n9369_));
OR2X2 OR2X2_3538 ( .A(core__abc_22172_new_n9363_), .B(core__abc_22172_new_n9369_), .Y(core__abc_22172_new_n9370_));
OR2X2 OR2X2_3539 ( .A(core__abc_22172_new_n9371_), .B(core__abc_22172_new_n9372_), .Y(core__abc_22172_new_n9373_));
OR2X2 OR2X2_354 ( .A(_abc_19873_new_n1720_), .B(_abc_19873_new_n1719_), .Y(_abc_19873_new_n1721_));
OR2X2 OR2X2_3540 ( .A(core_v0_reg_23_), .B(core_mi_reg_23_), .Y(core__abc_22172_new_n9376_));
OR2X2 OR2X2_3541 ( .A(core__abc_22172_new_n7555_), .B(core__abc_22172_new_n9380_), .Y(core__abc_22172_new_n9381_));
OR2X2 OR2X2_3542 ( .A(core__abc_22172_new_n9375_), .B(core__abc_22172_new_n9381_), .Y(core__abc_22172_new_n9382_));
OR2X2 OR2X2_3543 ( .A(core__abc_22172_new_n9383_), .B(core__abc_22172_new_n9384_), .Y(core__abc_22172_new_n9385_));
OR2X2 OR2X2_3544 ( .A(core_v0_reg_24_), .B(core_mi_reg_24_), .Y(core__abc_22172_new_n9388_));
OR2X2 OR2X2_3545 ( .A(core__abc_22172_new_n7593_), .B(core__abc_22172_new_n9392_), .Y(core__abc_22172_new_n9393_));
OR2X2 OR2X2_3546 ( .A(core__abc_22172_new_n9387_), .B(core__abc_22172_new_n9393_), .Y(core__abc_22172_new_n9394_));
OR2X2 OR2X2_3547 ( .A(core__abc_22172_new_n9395_), .B(core__abc_22172_new_n9396_), .Y(core__abc_22172_new_n9397_));
OR2X2 OR2X2_3548 ( .A(core_v0_reg_25_), .B(core_mi_reg_25_), .Y(core__abc_22172_new_n9401_));
OR2X2 OR2X2_3549 ( .A(core__abc_22172_new_n9400_), .B(core__abc_22172_new_n9405_), .Y(core__abc_22172_new_n9406_));
OR2X2 OR2X2_355 ( .A(_abc_19873_new_n1724_), .B(_abc_19873_new_n1723_), .Y(_abc_19873_new_n1725_));
OR2X2 OR2X2_3550 ( .A(core__abc_22172_new_n9399_), .B(core__abc_22172_new_n9406_), .Y(core__abc_22172_new_n9407_));
OR2X2 OR2X2_3551 ( .A(core__abc_22172_new_n9408_), .B(core__abc_22172_new_n9409_), .Y(core__abc_22172_new_n9410_));
OR2X2 OR2X2_3552 ( .A(core_v0_reg_26_), .B(core_mi_reg_26_), .Y(core__abc_22172_new_n9414_));
OR2X2 OR2X2_3553 ( .A(core__abc_22172_new_n9413_), .B(core__abc_22172_new_n9418_), .Y(core__abc_22172_new_n9419_));
OR2X2 OR2X2_3554 ( .A(core__abc_22172_new_n9412_), .B(core__abc_22172_new_n9419_), .Y(core__abc_22172_new_n9420_));
OR2X2 OR2X2_3555 ( .A(core__abc_22172_new_n9421_), .B(core__abc_22172_new_n9422_), .Y(core__abc_22172_new_n9423_));
OR2X2 OR2X2_3556 ( .A(core_v0_reg_27_), .B(core_mi_reg_27_), .Y(core__abc_22172_new_n9427_));
OR2X2 OR2X2_3557 ( .A(core__abc_22172_new_n9426_), .B(core__abc_22172_new_n9431_), .Y(core__abc_22172_new_n9432_));
OR2X2 OR2X2_3558 ( .A(core__abc_22172_new_n9425_), .B(core__abc_22172_new_n9432_), .Y(core__abc_22172_new_n9433_));
OR2X2 OR2X2_3559 ( .A(core__abc_22172_new_n9434_), .B(core__abc_22172_new_n9435_), .Y(core__abc_22172_new_n9436_));
OR2X2 OR2X2_356 ( .A(_abc_19873_new_n1728_), .B(_abc_19873_new_n1727_), .Y(_abc_19873_new_n1729_));
OR2X2 OR2X2_3560 ( .A(core_v0_reg_28_), .B(core_mi_reg_28_), .Y(core__abc_22172_new_n9441_));
OR2X2 OR2X2_3561 ( .A(core__abc_22172_new_n9440_), .B(core__abc_22172_new_n9445_), .Y(core__abc_22172_new_n9446_));
OR2X2 OR2X2_3562 ( .A(core__abc_22172_new_n9438_), .B(core__abc_22172_new_n9446_), .Y(core__abc_22172_new_n9447_));
OR2X2 OR2X2_3563 ( .A(core__abc_22172_new_n9448_), .B(core__abc_22172_new_n9449_), .Y(core__abc_22172_new_n9450_));
OR2X2 OR2X2_3564 ( .A(core_v0_reg_29_), .B(core_mi_reg_29_), .Y(core__abc_22172_new_n9453_));
OR2X2 OR2X2_3565 ( .A(core__abc_22172_new_n7730_), .B(core__abc_22172_new_n9457_), .Y(core__abc_22172_new_n9458_));
OR2X2 OR2X2_3566 ( .A(core__abc_22172_new_n9452_), .B(core__abc_22172_new_n9458_), .Y(core__abc_22172_new_n9459_));
OR2X2 OR2X2_3567 ( .A(core__abc_22172_new_n9460_), .B(core__abc_22172_new_n9461_), .Y(core__abc_22172_new_n9462_));
OR2X2 OR2X2_3568 ( .A(core_v0_reg_30_), .B(core_mi_reg_30_), .Y(core__abc_22172_new_n9465_));
OR2X2 OR2X2_3569 ( .A(core__abc_22172_new_n7759_), .B(core__abc_22172_new_n9469_), .Y(core__abc_22172_new_n9470_));
OR2X2 OR2X2_357 ( .A(_abc_19873_new_n1732_), .B(_abc_19873_new_n1731_), .Y(_abc_19873_new_n1733_));
OR2X2 OR2X2_3570 ( .A(core__abc_22172_new_n9464_), .B(core__abc_22172_new_n9470_), .Y(core__abc_22172_new_n9471_));
OR2X2 OR2X2_3571 ( .A(core__abc_22172_new_n9472_), .B(core__abc_22172_new_n9473_), .Y(core__abc_22172_new_n9474_));
OR2X2 OR2X2_3572 ( .A(core_v0_reg_31_), .B(core_mi_reg_31_), .Y(core__abc_22172_new_n9477_));
OR2X2 OR2X2_3573 ( .A(core__abc_22172_new_n7782_), .B(core__abc_22172_new_n9481_), .Y(core__abc_22172_new_n9482_));
OR2X2 OR2X2_3574 ( .A(core__abc_22172_new_n9476_), .B(core__abc_22172_new_n9482_), .Y(core__abc_22172_new_n9483_));
OR2X2 OR2X2_3575 ( .A(core__abc_22172_new_n9484_), .B(core__abc_22172_new_n9485_), .Y(core__abc_22172_new_n9486_));
OR2X2 OR2X2_3576 ( .A(core_v0_reg_32_), .B(core_mi_reg_32_), .Y(core__abc_22172_new_n9489_));
OR2X2 OR2X2_3577 ( .A(core__abc_22172_new_n7791_), .B(core__abc_22172_new_n9493_), .Y(core__abc_22172_new_n9494_));
OR2X2 OR2X2_3578 ( .A(core__abc_22172_new_n9488_), .B(core__abc_22172_new_n9494_), .Y(core__abc_22172_new_n9495_));
OR2X2 OR2X2_3579 ( .A(core__abc_22172_new_n9496_), .B(core__abc_22172_new_n9497_), .Y(core__abc_22172_new_n9498_));
OR2X2 OR2X2_358 ( .A(_abc_19873_new_n1736_), .B(_abc_19873_new_n1735_), .Y(_abc_19873_new_n1737_));
OR2X2 OR2X2_3580 ( .A(core_v0_reg_33_), .B(core_mi_reg_33_), .Y(core__abc_22172_new_n9501_));
OR2X2 OR2X2_3581 ( .A(core__abc_22172_new_n7803_), .B(core__abc_22172_new_n9505_), .Y(core__abc_22172_new_n9506_));
OR2X2 OR2X2_3582 ( .A(core__abc_22172_new_n9500_), .B(core__abc_22172_new_n9506_), .Y(core__abc_22172_new_n9507_));
OR2X2 OR2X2_3583 ( .A(core__abc_22172_new_n9508_), .B(core__abc_22172_new_n9509_), .Y(core__abc_22172_new_n9510_));
OR2X2 OR2X2_3584 ( .A(core_v0_reg_34_), .B(core_mi_reg_34_), .Y(core__abc_22172_new_n9513_));
OR2X2 OR2X2_3585 ( .A(core__abc_22172_new_n7817_), .B(core__abc_22172_new_n9517_), .Y(core__abc_22172_new_n9518_));
OR2X2 OR2X2_3586 ( .A(core__abc_22172_new_n9512_), .B(core__abc_22172_new_n9518_), .Y(core__abc_22172_new_n9519_));
OR2X2 OR2X2_3587 ( .A(core__abc_22172_new_n9520_), .B(core__abc_22172_new_n9521_), .Y(core__abc_22172_new_n9522_));
OR2X2 OR2X2_3588 ( .A(core_v0_reg_35_), .B(core_mi_reg_35_), .Y(core__abc_22172_new_n9525_));
OR2X2 OR2X2_3589 ( .A(core__abc_22172_new_n7834_), .B(core__abc_22172_new_n9529_), .Y(core__abc_22172_new_n9530_));
OR2X2 OR2X2_359 ( .A(_abc_19873_new_n1740_), .B(_abc_19873_new_n1739_), .Y(_abc_19873_new_n1741_));
OR2X2 OR2X2_3590 ( .A(core__abc_22172_new_n9524_), .B(core__abc_22172_new_n9530_), .Y(core__abc_22172_new_n9531_));
OR2X2 OR2X2_3591 ( .A(core__abc_22172_new_n9532_), .B(core__abc_22172_new_n9533_), .Y(core__abc_22172_new_n9534_));
OR2X2 OR2X2_3592 ( .A(core_v0_reg_36_), .B(core_mi_reg_36_), .Y(core__abc_22172_new_n9537_));
OR2X2 OR2X2_3593 ( .A(core__abc_22172_new_n7846_), .B(core__abc_22172_new_n9541_), .Y(core__abc_22172_new_n9542_));
OR2X2 OR2X2_3594 ( .A(core__abc_22172_new_n9536_), .B(core__abc_22172_new_n9542_), .Y(core__abc_22172_new_n9543_));
OR2X2 OR2X2_3595 ( .A(core__abc_22172_new_n9544_), .B(core__abc_22172_new_n9545_), .Y(core__abc_22172_new_n9546_));
OR2X2 OR2X2_3596 ( .A(core_v0_reg_37_), .B(core_mi_reg_37_), .Y(core__abc_22172_new_n9549_));
OR2X2 OR2X2_3597 ( .A(core__abc_22172_new_n7864_), .B(core__abc_22172_new_n9553_), .Y(core__abc_22172_new_n9554_));
OR2X2 OR2X2_3598 ( .A(core__abc_22172_new_n9548_), .B(core__abc_22172_new_n9554_), .Y(core__abc_22172_new_n9555_));
OR2X2 OR2X2_3599 ( .A(core__abc_22172_new_n9556_), .B(core__abc_22172_new_n9557_), .Y(core__abc_22172_new_n9558_));
OR2X2 OR2X2_36 ( .A(_abc_19873_new_n990_), .B(_abc_19873_new_n991_), .Y(_abc_19873_new_n992_));
OR2X2 OR2X2_360 ( .A(_abc_19873_new_n1744_), .B(_abc_19873_new_n1743_), .Y(_abc_19873_new_n1745_));
OR2X2 OR2X2_3600 ( .A(core_v0_reg_38_), .B(core_mi_reg_38_), .Y(core__abc_22172_new_n9561_));
OR2X2 OR2X2_3601 ( .A(core__abc_22172_new_n7878_), .B(core__abc_22172_new_n9565_), .Y(core__abc_22172_new_n9566_));
OR2X2 OR2X2_3602 ( .A(core__abc_22172_new_n9560_), .B(core__abc_22172_new_n9566_), .Y(core__abc_22172_new_n9567_));
OR2X2 OR2X2_3603 ( .A(core__abc_22172_new_n9568_), .B(core__abc_22172_new_n9569_), .Y(core__abc_22172_new_n9570_));
OR2X2 OR2X2_3604 ( .A(core_v0_reg_39_), .B(core_mi_reg_39_), .Y(core__abc_22172_new_n9573_));
OR2X2 OR2X2_3605 ( .A(core__abc_22172_new_n7893_), .B(core__abc_22172_new_n9577_), .Y(core__abc_22172_new_n9578_));
OR2X2 OR2X2_3606 ( .A(core__abc_22172_new_n9572_), .B(core__abc_22172_new_n9578_), .Y(core__abc_22172_new_n9579_));
OR2X2 OR2X2_3607 ( .A(core__abc_22172_new_n9580_), .B(core__abc_22172_new_n9581_), .Y(core__abc_22172_new_n9582_));
OR2X2 OR2X2_3608 ( .A(core_v0_reg_40_), .B(core_mi_reg_40_), .Y(core__abc_22172_new_n9585_));
OR2X2 OR2X2_3609 ( .A(core__abc_22172_new_n7907_), .B(core__abc_22172_new_n9589_), .Y(core__abc_22172_new_n9590_));
OR2X2 OR2X2_361 ( .A(_abc_19873_new_n1748_), .B(_abc_19873_new_n1747_), .Y(_abc_19873_new_n1749_));
OR2X2 OR2X2_3610 ( .A(core__abc_22172_new_n9584_), .B(core__abc_22172_new_n9590_), .Y(core__abc_22172_new_n9591_));
OR2X2 OR2X2_3611 ( .A(core__abc_22172_new_n9592_), .B(core__abc_22172_new_n9593_), .Y(core__abc_22172_new_n9594_));
OR2X2 OR2X2_3612 ( .A(core_v0_reg_41_), .B(core_mi_reg_41_), .Y(core__abc_22172_new_n9598_));
OR2X2 OR2X2_3613 ( .A(core__abc_22172_new_n9597_), .B(core__abc_22172_new_n9602_), .Y(core__abc_22172_new_n9603_));
OR2X2 OR2X2_3614 ( .A(core__abc_22172_new_n9596_), .B(core__abc_22172_new_n9603_), .Y(core__abc_22172_new_n9604_));
OR2X2 OR2X2_3615 ( .A(core__abc_22172_new_n9605_), .B(core__abc_22172_new_n9606_), .Y(core__abc_22172_new_n9607_));
OR2X2 OR2X2_3616 ( .A(core_v0_reg_42_), .B(core_mi_reg_42_), .Y(core__abc_22172_new_n9610_));
OR2X2 OR2X2_3617 ( .A(core__abc_22172_new_n7940_), .B(core__abc_22172_new_n9614_), .Y(core__abc_22172_new_n9615_));
OR2X2 OR2X2_3618 ( .A(core__abc_22172_new_n9609_), .B(core__abc_22172_new_n9615_), .Y(core__abc_22172_new_n9616_));
OR2X2 OR2X2_3619 ( .A(core__abc_22172_new_n9617_), .B(core__abc_22172_new_n9618_), .Y(core__abc_22172_new_n9619_));
OR2X2 OR2X2_362 ( .A(_abc_19873_new_n1752_), .B(_abc_19873_new_n1751_), .Y(_abc_19873_new_n1753_));
OR2X2 OR2X2_3620 ( .A(core_v0_reg_43_), .B(core_mi_reg_43_), .Y(core__abc_22172_new_n9624_));
OR2X2 OR2X2_3621 ( .A(core__abc_22172_new_n9623_), .B(core__abc_22172_new_n9628_), .Y(core__abc_22172_new_n9629_));
OR2X2 OR2X2_3622 ( .A(core__abc_22172_new_n9621_), .B(core__abc_22172_new_n9629_), .Y(core__abc_22172_new_n9630_));
OR2X2 OR2X2_3623 ( .A(core__abc_22172_new_n9631_), .B(core__abc_22172_new_n9632_), .Y(core__abc_22172_new_n9633_));
OR2X2 OR2X2_3624 ( .A(core_v0_reg_44_), .B(core_mi_reg_44_), .Y(core__abc_22172_new_n9636_));
OR2X2 OR2X2_3625 ( .A(core__abc_22172_new_n7969_), .B(core__abc_22172_new_n9640_), .Y(core__abc_22172_new_n9641_));
OR2X2 OR2X2_3626 ( .A(core__abc_22172_new_n9635_), .B(core__abc_22172_new_n9641_), .Y(core__abc_22172_new_n9642_));
OR2X2 OR2X2_3627 ( .A(core__abc_22172_new_n9643_), .B(core__abc_22172_new_n9644_), .Y(core__abc_22172_new_n9645_));
OR2X2 OR2X2_3628 ( .A(core_v0_reg_45_), .B(core_mi_reg_45_), .Y(core__abc_22172_new_n9648_));
OR2X2 OR2X2_3629 ( .A(core__abc_22172_new_n7985_), .B(core__abc_22172_new_n9652_), .Y(core__abc_22172_new_n9653_));
OR2X2 OR2X2_363 ( .A(_abc_19873_new_n1756_), .B(_abc_19873_new_n1755_), .Y(_abc_19873_new_n1757_));
OR2X2 OR2X2_3630 ( .A(core__abc_22172_new_n9647_), .B(core__abc_22172_new_n9653_), .Y(core__abc_22172_new_n9654_));
OR2X2 OR2X2_3631 ( .A(core__abc_22172_new_n9655_), .B(core__abc_22172_new_n9656_), .Y(core__abc_22172_new_n9657_));
OR2X2 OR2X2_3632 ( .A(core_v0_reg_46_), .B(core_mi_reg_46_), .Y(core__abc_22172_new_n9660_));
OR2X2 OR2X2_3633 ( .A(core__abc_22172_new_n8002_), .B(core__abc_22172_new_n9664_), .Y(core__abc_22172_new_n9665_));
OR2X2 OR2X2_3634 ( .A(core__abc_22172_new_n9659_), .B(core__abc_22172_new_n9665_), .Y(core__abc_22172_new_n9666_));
OR2X2 OR2X2_3635 ( .A(core__abc_22172_new_n9667_), .B(core__abc_22172_new_n9668_), .Y(core__abc_22172_new_n9669_));
OR2X2 OR2X2_3636 ( .A(core_v0_reg_47_), .B(core_mi_reg_47_), .Y(core__abc_22172_new_n9672_));
OR2X2 OR2X2_3637 ( .A(core__abc_22172_new_n8018_), .B(core__abc_22172_new_n9676_), .Y(core__abc_22172_new_n9677_));
OR2X2 OR2X2_3638 ( .A(core__abc_22172_new_n9671_), .B(core__abc_22172_new_n9677_), .Y(core__abc_22172_new_n9678_));
OR2X2 OR2X2_3639 ( .A(core__abc_22172_new_n9679_), .B(core__abc_22172_new_n9680_), .Y(core__abc_22172_new_n9681_));
OR2X2 OR2X2_364 ( .A(_abc_19873_new_n1760_), .B(_abc_19873_new_n1759_), .Y(_abc_19873_new_n1761_));
OR2X2 OR2X2_3640 ( .A(core_v0_reg_48_), .B(core_mi_reg_48_), .Y(core__abc_22172_new_n9684_));
OR2X2 OR2X2_3641 ( .A(core__abc_22172_new_n8033_), .B(core__abc_22172_new_n9688_), .Y(core__abc_22172_new_n9689_));
OR2X2 OR2X2_3642 ( .A(core__abc_22172_new_n9683_), .B(core__abc_22172_new_n9689_), .Y(core__abc_22172_new_n9690_));
OR2X2 OR2X2_3643 ( .A(core__abc_22172_new_n9691_), .B(core__abc_22172_new_n9692_), .Y(core__abc_22172_new_n9693_));
OR2X2 OR2X2_3644 ( .A(core_v0_reg_49_), .B(core_mi_reg_49_), .Y(core__abc_22172_new_n9698_));
OR2X2 OR2X2_3645 ( .A(core__abc_22172_new_n9697_), .B(core__abc_22172_new_n9702_), .Y(core__abc_22172_new_n9703_));
OR2X2 OR2X2_3646 ( .A(core__abc_22172_new_n9695_), .B(core__abc_22172_new_n9703_), .Y(core__abc_22172_new_n9704_));
OR2X2 OR2X2_3647 ( .A(core__abc_22172_new_n9705_), .B(core__abc_22172_new_n9706_), .Y(core__abc_22172_new_n9707_));
OR2X2 OR2X2_3648 ( .A(core_v0_reg_50_), .B(core_mi_reg_50_), .Y(core__abc_22172_new_n9712_));
OR2X2 OR2X2_3649 ( .A(core__abc_22172_new_n9711_), .B(core__abc_22172_new_n9716_), .Y(core__abc_22172_new_n9717_));
OR2X2 OR2X2_365 ( .A(_abc_19873_new_n1764_), .B(_abc_19873_new_n1763_), .Y(_abc_19873_new_n1765_));
OR2X2 OR2X2_3650 ( .A(core__abc_22172_new_n9709_), .B(core__abc_22172_new_n9717_), .Y(core__abc_22172_new_n9718_));
OR2X2 OR2X2_3651 ( .A(core__abc_22172_new_n9719_), .B(core__abc_22172_new_n9720_), .Y(core__abc_22172_new_n9721_));
OR2X2 OR2X2_3652 ( .A(core_v0_reg_51_), .B(core_mi_reg_51_), .Y(core__abc_22172_new_n9724_));
OR2X2 OR2X2_3653 ( .A(core__abc_22172_new_n8079_), .B(core__abc_22172_new_n9728_), .Y(core__abc_22172_new_n9729_));
OR2X2 OR2X2_3654 ( .A(core__abc_22172_new_n9723_), .B(core__abc_22172_new_n9729_), .Y(core__abc_22172_new_n9730_));
OR2X2 OR2X2_3655 ( .A(core__abc_22172_new_n9731_), .B(core__abc_22172_new_n9732_), .Y(core__abc_22172_new_n9733_));
OR2X2 OR2X2_3656 ( .A(core_v0_reg_52_), .B(core_mi_reg_52_), .Y(core__abc_22172_new_n9737_));
OR2X2 OR2X2_3657 ( .A(core__abc_22172_new_n9736_), .B(core__abc_22172_new_n9741_), .Y(core__abc_22172_new_n9742_));
OR2X2 OR2X2_3658 ( .A(core__abc_22172_new_n9735_), .B(core__abc_22172_new_n9742_), .Y(core__abc_22172_new_n9743_));
OR2X2 OR2X2_3659 ( .A(core__abc_22172_new_n9744_), .B(core__abc_22172_new_n9745_), .Y(core__abc_22172_new_n9746_));
OR2X2 OR2X2_366 ( .A(_abc_19873_new_n1768_), .B(_abc_19873_new_n1767_), .Y(_abc_19873_new_n1769_));
OR2X2 OR2X2_3660 ( .A(core_v0_reg_53_), .B(core_mi_reg_53_), .Y(core__abc_22172_new_n9749_));
OR2X2 OR2X2_3661 ( .A(core__abc_22172_new_n8114_), .B(core__abc_22172_new_n9753_), .Y(core__abc_22172_new_n9754_));
OR2X2 OR2X2_3662 ( .A(core__abc_22172_new_n9748_), .B(core__abc_22172_new_n9754_), .Y(core__abc_22172_new_n9755_));
OR2X2 OR2X2_3663 ( .A(core__abc_22172_new_n9756_), .B(core__abc_22172_new_n9757_), .Y(core__abc_22172_new_n9758_));
OR2X2 OR2X2_3664 ( .A(core_v0_reg_54_), .B(core_mi_reg_54_), .Y(core__abc_22172_new_n9761_));
OR2X2 OR2X2_3665 ( .A(core__abc_22172_new_n8130_), .B(core__abc_22172_new_n9765_), .Y(core__abc_22172_new_n9766_));
OR2X2 OR2X2_3666 ( .A(core__abc_22172_new_n9760_), .B(core__abc_22172_new_n9766_), .Y(core__abc_22172_new_n9767_));
OR2X2 OR2X2_3667 ( .A(core__abc_22172_new_n9768_), .B(core__abc_22172_new_n9769_), .Y(core__abc_22172_new_n9770_));
OR2X2 OR2X2_3668 ( .A(core_v0_reg_55_), .B(core_mi_reg_55_), .Y(core__abc_22172_new_n9773_));
OR2X2 OR2X2_3669 ( .A(core__abc_22172_new_n8146_), .B(core__abc_22172_new_n9777_), .Y(core__abc_22172_new_n9778_));
OR2X2 OR2X2_367 ( .A(_abc_19873_new_n1772_), .B(_abc_19873_new_n1771_), .Y(_abc_19873_new_n1773_));
OR2X2 OR2X2_3670 ( .A(core__abc_22172_new_n9772_), .B(core__abc_22172_new_n9778_), .Y(core__abc_22172_new_n9779_));
OR2X2 OR2X2_3671 ( .A(core__abc_22172_new_n9780_), .B(core__abc_22172_new_n9781_), .Y(core__abc_22172_new_n9782_));
OR2X2 OR2X2_3672 ( .A(core_v0_reg_56_), .B(core_mi_reg_56_), .Y(core__abc_22172_new_n9787_));
OR2X2 OR2X2_3673 ( .A(core__abc_22172_new_n9786_), .B(core__abc_22172_new_n9791_), .Y(core__abc_22172_new_n9792_));
OR2X2 OR2X2_3674 ( .A(core__abc_22172_new_n9784_), .B(core__abc_22172_new_n9792_), .Y(core__abc_22172_new_n9793_));
OR2X2 OR2X2_3675 ( .A(core__abc_22172_new_n9794_), .B(core__abc_22172_new_n9795_), .Y(core__abc_22172_new_n9796_));
OR2X2 OR2X2_3676 ( .A(core_v0_reg_57_), .B(core_mi_reg_57_), .Y(core__abc_22172_new_n9801_));
OR2X2 OR2X2_3677 ( .A(core__abc_22172_new_n9800_), .B(core__abc_22172_new_n9805_), .Y(core__abc_22172_new_n9806_));
OR2X2 OR2X2_3678 ( .A(core__abc_22172_new_n9798_), .B(core__abc_22172_new_n9806_), .Y(core__abc_22172_new_n9807_));
OR2X2 OR2X2_3679 ( .A(core__abc_22172_new_n9808_), .B(core__abc_22172_new_n9809_), .Y(core__abc_22172_new_n9810_));
OR2X2 OR2X2_368 ( .A(_abc_19873_new_n1776_), .B(_abc_19873_new_n1775_), .Y(_abc_19873_new_n1777_));
OR2X2 OR2X2_3680 ( .A(core_v0_reg_58_), .B(core_mi_reg_58_), .Y(core__abc_22172_new_n9814_));
OR2X2 OR2X2_3681 ( .A(core__abc_22172_new_n9813_), .B(core__abc_22172_new_n9818_), .Y(core__abc_22172_new_n9819_));
OR2X2 OR2X2_3682 ( .A(core__abc_22172_new_n9812_), .B(core__abc_22172_new_n9819_), .Y(core__abc_22172_new_n9820_));
OR2X2 OR2X2_3683 ( .A(core__abc_22172_new_n9821_), .B(core__abc_22172_new_n9822_), .Y(core__abc_22172_new_n9823_));
OR2X2 OR2X2_3684 ( .A(core_v0_reg_59_), .B(core_mi_reg_59_), .Y(core__abc_22172_new_n9827_));
OR2X2 OR2X2_3685 ( .A(core__abc_22172_new_n9826_), .B(core__abc_22172_new_n9831_), .Y(core__abc_22172_new_n9832_));
OR2X2 OR2X2_3686 ( .A(core__abc_22172_new_n9825_), .B(core__abc_22172_new_n9832_), .Y(core__abc_22172_new_n9833_));
OR2X2 OR2X2_3687 ( .A(core__abc_22172_new_n9834_), .B(core__abc_22172_new_n9835_), .Y(core__abc_22172_new_n9836_));
OR2X2 OR2X2_3688 ( .A(core_v0_reg_60_), .B(core_mi_reg_60_), .Y(core__abc_22172_new_n9841_));
OR2X2 OR2X2_3689 ( .A(core__abc_22172_new_n9840_), .B(core__abc_22172_new_n9845_), .Y(core__abc_22172_new_n9846_));
OR2X2 OR2X2_369 ( .A(_abc_19873_new_n1780_), .B(_abc_19873_new_n1779_), .Y(_abc_19873_new_n1781_));
OR2X2 OR2X2_3690 ( .A(core__abc_22172_new_n9838_), .B(core__abc_22172_new_n9846_), .Y(core__abc_22172_new_n9847_));
OR2X2 OR2X2_3691 ( .A(core__abc_22172_new_n9848_), .B(core__abc_22172_new_n9849_), .Y(core__abc_22172_new_n9850_));
OR2X2 OR2X2_3692 ( .A(core_v0_reg_61_), .B(core_mi_reg_61_), .Y(core__abc_22172_new_n9853_));
OR2X2 OR2X2_3693 ( .A(core__abc_22172_new_n8242_), .B(core__abc_22172_new_n9857_), .Y(core__abc_22172_new_n9858_));
OR2X2 OR2X2_3694 ( .A(core__abc_22172_new_n9852_), .B(core__abc_22172_new_n9858_), .Y(core__abc_22172_new_n9859_));
OR2X2 OR2X2_3695 ( .A(core__abc_22172_new_n9860_), .B(core__abc_22172_new_n9861_), .Y(core__abc_22172_new_n9862_));
OR2X2 OR2X2_3696 ( .A(core_v0_reg_62_), .B(core_mi_reg_62_), .Y(core__abc_22172_new_n9865_));
OR2X2 OR2X2_3697 ( .A(core__abc_22172_new_n8258_), .B(core__abc_22172_new_n9869_), .Y(core__abc_22172_new_n9870_));
OR2X2 OR2X2_3698 ( .A(core__abc_22172_new_n9864_), .B(core__abc_22172_new_n9870_), .Y(core__abc_22172_new_n9871_));
OR2X2 OR2X2_3699 ( .A(core__abc_22172_new_n9872_), .B(core__abc_22172_new_n9873_), .Y(core__abc_22172_new_n9874_));
OR2X2 OR2X2_37 ( .A(_abc_19873_new_n993_), .B(_abc_19873_new_n994_), .Y(_abc_19873_new_n995_));
OR2X2 OR2X2_370 ( .A(_abc_19873_new_n1784_), .B(_abc_19873_new_n1783_), .Y(_abc_19873_new_n1785_));
OR2X2 OR2X2_3700 ( .A(core_v0_reg_63_), .B(core_mi_reg_63_), .Y(core__abc_22172_new_n9877_));
OR2X2 OR2X2_3701 ( .A(core__abc_22172_new_n8274_), .B(core__abc_22172_new_n9881_), .Y(core__abc_22172_new_n9882_));
OR2X2 OR2X2_3702 ( .A(core__abc_22172_new_n9876_), .B(core__abc_22172_new_n9882_), .Y(core__abc_22172_new_n9883_));
OR2X2 OR2X2_3703 ( .A(core__abc_22172_new_n9884_), .B(core__abc_22172_new_n9885_), .Y(core__abc_22172_new_n9886_));
OR2X2 OR2X2_3704 ( .A(core__abc_22172_new_n9895_), .B(core__abc_22172_new_n1213_), .Y(core__abc_22172_new_n9896_));
OR2X2 OR2X2_3705 ( .A(core__abc_22172_new_n9897_), .B(core__abc_22172_new_n1170_), .Y(core__abc_22172_new_n9898_));
OR2X2 OR2X2_371 ( .A(_abc_19873_new_n1788_), .B(_abc_19873_new_n1787_), .Y(_abc_19873_new_n1789_));
OR2X2 OR2X2_372 ( .A(_abc_19873_new_n1792_), .B(_abc_19873_new_n1791_), .Y(_abc_19873_new_n1793_));
OR2X2 OR2X2_373 ( .A(_abc_19873_new_n1796_), .B(_abc_19873_new_n1795_), .Y(_abc_19873_new_n1797_));
OR2X2 OR2X2_374 ( .A(_abc_19873_new_n1800_), .B(_abc_19873_new_n1799_), .Y(_abc_19873_new_n1801_));
OR2X2 OR2X2_375 ( .A(_abc_19873_new_n1804_), .B(_abc_19873_new_n1803_), .Y(_abc_19873_new_n1805_));
OR2X2 OR2X2_376 ( .A(_abc_19873_new_n1808_), .B(_abc_19873_new_n1807_), .Y(_abc_19873_new_n1809_));
OR2X2 OR2X2_377 ( .A(_abc_19873_new_n1812_), .B(_abc_19873_new_n1811_), .Y(_abc_19873_new_n1813_));
OR2X2 OR2X2_378 ( .A(_abc_19873_new_n1816_), .B(_abc_19873_new_n1815_), .Y(_abc_19873_new_n1817_));
OR2X2 OR2X2_379 ( .A(_abc_19873_new_n1820_), .B(_abc_19873_new_n1819_), .Y(_abc_19873_new_n1821_));
OR2X2 OR2X2_38 ( .A(_abc_19873_new_n992_), .B(_abc_19873_new_n995_), .Y(_abc_19873_new_n996_));
OR2X2 OR2X2_380 ( .A(_abc_19873_new_n1824_), .B(_abc_19873_new_n1823_), .Y(_abc_19873_new_n1825_));
OR2X2 OR2X2_381 ( .A(_abc_19873_new_n1828_), .B(_abc_19873_new_n1827_), .Y(_abc_19873_new_n1829_));
OR2X2 OR2X2_382 ( .A(_abc_19873_new_n1832_), .B(_abc_19873_new_n1831_), .Y(_abc_19873_new_n1833_));
OR2X2 OR2X2_383 ( .A(_abc_19873_new_n1836_), .B(_abc_19873_new_n1835_), .Y(_abc_19873_new_n1837_));
OR2X2 OR2X2_384 ( .A(_abc_19873_new_n1840_), .B(_abc_19873_new_n1839_), .Y(_abc_19873_new_n1841_));
OR2X2 OR2X2_385 ( .A(_abc_19873_new_n1844_), .B(_abc_19873_new_n1843_), .Y(_abc_19873_new_n1845_));
OR2X2 OR2X2_386 ( .A(_abc_19873_new_n1848_), .B(_abc_19873_new_n1847_), .Y(_abc_19873_new_n1849_));
OR2X2 OR2X2_387 ( .A(_abc_19873_new_n1852_), .B(_abc_19873_new_n1851_), .Y(_abc_19873_new_n1853_));
OR2X2 OR2X2_388 ( .A(_abc_19873_new_n1856_), .B(_abc_19873_new_n1855_), .Y(_abc_19873_new_n1857_));
OR2X2 OR2X2_389 ( .A(_abc_19873_new_n1860_), .B(_abc_19873_new_n1859_), .Y(_abc_19873_new_n1861_));
OR2X2 OR2X2_39 ( .A(_abc_19873_new_n996_), .B(_abc_19873_new_n989_), .Y(_abc_19873_new_n997_));
OR2X2 OR2X2_390 ( .A(_abc_19873_new_n1864_), .B(_abc_19873_new_n1863_), .Y(_abc_19873_new_n1865_));
OR2X2 OR2X2_391 ( .A(_abc_19873_new_n1868_), .B(_abc_19873_new_n1867_), .Y(_abc_19873_new_n1869_));
OR2X2 OR2X2_392 ( .A(_abc_19873_new_n1872_), .B(_abc_19873_new_n1871_), .Y(_abc_19873_new_n1873_));
OR2X2 OR2X2_393 ( .A(_abc_19873_new_n1876_), .B(_abc_19873_new_n1875_), .Y(_abc_19873_new_n1877_));
OR2X2 OR2X2_394 ( .A(_abc_19873_new_n1880_), .B(_abc_19873_new_n1879_), .Y(_abc_19873_new_n1881_));
OR2X2 OR2X2_395 ( .A(_abc_19873_new_n1884_), .B(_abc_19873_new_n1883_), .Y(_abc_19873_new_n1885_));
OR2X2 OR2X2_396 ( .A(_abc_19873_new_n1888_), .B(_abc_19873_new_n1887_), .Y(_abc_19873_new_n1889_));
OR2X2 OR2X2_397 ( .A(_abc_19873_new_n1892_), .B(_abc_19873_new_n1891_), .Y(_abc_19873_new_n1893_));
OR2X2 OR2X2_398 ( .A(_abc_19873_new_n1896_), .B(_abc_19873_new_n1895_), .Y(_abc_19873_new_n1897_));
OR2X2 OR2X2_399 ( .A(_abc_19873_new_n1900_), .B(_abc_19873_new_n1899_), .Y(_abc_19873_new_n1901_));
OR2X2 OR2X2_4 ( .A(_abc_19873_new_n899_), .B(_abc_19873_new_n909_), .Y(_abc_19873_new_n910_));
OR2X2 OR2X2_40 ( .A(_abc_19873_new_n999_), .B(_abc_19873_new_n1000_), .Y(_abc_19873_new_n1001_));
OR2X2 OR2X2_400 ( .A(_abc_19873_new_n1904_), .B(_abc_19873_new_n1903_), .Y(_abc_19873_new_n1905_));
OR2X2 OR2X2_401 ( .A(_abc_19873_new_n1908_), .B(_abc_19873_new_n1907_), .Y(_abc_19873_new_n1909_));
OR2X2 OR2X2_402 ( .A(_abc_19873_new_n1912_), .B(_abc_19873_new_n1911_), .Y(_abc_19873_new_n1913_));
OR2X2 OR2X2_403 ( .A(_abc_19873_new_n1916_), .B(_abc_19873_new_n1915_), .Y(_abc_19873_new_n1917_));
OR2X2 OR2X2_404 ( .A(_abc_19873_new_n1920_), .B(_abc_19873_new_n1919_), .Y(_abc_19873_new_n1921_));
OR2X2 OR2X2_405 ( .A(_abc_19873_new_n1924_), .B(_abc_19873_new_n1923_), .Y(_abc_19873_new_n1925_));
OR2X2 OR2X2_406 ( .A(_abc_19873_new_n1928_), .B(_abc_19873_new_n1927_), .Y(_abc_19873_new_n1929_));
OR2X2 OR2X2_407 ( .A(_abc_19873_new_n1932_), .B(_abc_19873_new_n1931_), .Y(_abc_19873_new_n1933_));
OR2X2 OR2X2_408 ( .A(_abc_19873_new_n1936_), .B(_abc_19873_new_n1935_), .Y(_abc_19873_new_n1937_));
OR2X2 OR2X2_409 ( .A(_abc_19873_new_n1940_), .B(_abc_19873_new_n1939_), .Y(_abc_19873_new_n1941_));
OR2X2 OR2X2_41 ( .A(_abc_19873_new_n1001_), .B(_abc_19873_new_n998_), .Y(_abc_19873_new_n1002_));
OR2X2 OR2X2_410 ( .A(_abc_19873_new_n1944_), .B(_abc_19873_new_n1943_), .Y(_abc_19873_new_n1945_));
OR2X2 OR2X2_411 ( .A(_abc_19873_new_n1948_), .B(_abc_19873_new_n1947_), .Y(_abc_19873_new_n1949_));
OR2X2 OR2X2_412 ( .A(_abc_19873_new_n1952_), .B(_abc_19873_new_n1951_), .Y(_abc_19873_new_n1953_));
OR2X2 OR2X2_413 ( .A(_abc_19873_new_n1956_), .B(_abc_19873_new_n1955_), .Y(_abc_19873_new_n1957_));
OR2X2 OR2X2_414 ( .A(_abc_19873_new_n1960_), .B(_abc_19873_new_n1959_), .Y(_abc_19873_new_n1961_));
OR2X2 OR2X2_415 ( .A(_abc_19873_new_n1964_), .B(_abc_19873_new_n1963_), .Y(_abc_19873_new_n1965_));
OR2X2 OR2X2_416 ( .A(_abc_19873_new_n1968_), .B(_abc_19873_new_n1967_), .Y(_abc_19873_new_n1969_));
OR2X2 OR2X2_417 ( .A(_abc_19873_new_n1972_), .B(_abc_19873_new_n1971_), .Y(_abc_19873_new_n1973_));
OR2X2 OR2X2_418 ( .A(_abc_19873_new_n1976_), .B(_abc_19873_new_n1975_), .Y(_abc_19873_new_n1977_));
OR2X2 OR2X2_419 ( .A(_abc_19873_new_n1980_), .B(_abc_19873_new_n1979_), .Y(_abc_19873_new_n1981_));
OR2X2 OR2X2_42 ( .A(_abc_19873_new_n1003_), .B(_abc_19873_new_n1004_), .Y(_abc_19873_new_n1005_));
OR2X2 OR2X2_420 ( .A(_abc_19873_new_n1984_), .B(_abc_19873_new_n1983_), .Y(_abc_19873_new_n1985_));
OR2X2 OR2X2_421 ( .A(_abc_19873_new_n1988_), .B(_abc_19873_new_n1987_), .Y(_abc_19873_new_n1989_));
OR2X2 OR2X2_422 ( .A(_abc_19873_new_n1992_), .B(_abc_19873_new_n1991_), .Y(_abc_19873_new_n1993_));
OR2X2 OR2X2_423 ( .A(_abc_19873_new_n1996_), .B(_abc_19873_new_n1995_), .Y(_abc_19873_new_n1997_));
OR2X2 OR2X2_424 ( .A(_abc_19873_new_n2000_), .B(_abc_19873_new_n1999_), .Y(_abc_19873_new_n2001_));
OR2X2 OR2X2_425 ( .A(_abc_19873_new_n2004_), .B(_abc_19873_new_n2003_), .Y(_abc_19873_new_n2005_));
OR2X2 OR2X2_426 ( .A(_abc_19873_new_n2008_), .B(_abc_19873_new_n2007_), .Y(_abc_19873_new_n2009_));
OR2X2 OR2X2_427 ( .A(_abc_19873_new_n2012_), .B(_abc_19873_new_n2011_), .Y(_abc_19873_new_n2013_));
OR2X2 OR2X2_428 ( .A(_abc_19873_new_n2016_), .B(_abc_19873_new_n2015_), .Y(_abc_19873_new_n2017_));
OR2X2 OR2X2_429 ( .A(_abc_19873_new_n2020_), .B(_abc_19873_new_n2019_), .Y(_abc_19873_new_n2021_));
OR2X2 OR2X2_43 ( .A(_abc_19873_new_n1006_), .B(_abc_19873_new_n1007_), .Y(_abc_19873_new_n1008_));
OR2X2 OR2X2_430 ( .A(_abc_19873_new_n2024_), .B(_abc_19873_new_n2023_), .Y(_abc_19873_new_n2025_));
OR2X2 OR2X2_431 ( .A(_abc_19873_new_n2028_), .B(_abc_19873_new_n2027_), .Y(_abc_19873_new_n2029_));
OR2X2 OR2X2_432 ( .A(_abc_19873_new_n2032_), .B(_abc_19873_new_n2031_), .Y(_abc_19873_new_n2033_));
OR2X2 OR2X2_433 ( .A(_abc_19873_new_n2036_), .B(_abc_19873_new_n2035_), .Y(_abc_19873_new_n2037_));
OR2X2 OR2X2_434 ( .A(_abc_19873_new_n2040_), .B(_abc_19873_new_n2039_), .Y(_abc_19873_new_n2041_));
OR2X2 OR2X2_435 ( .A(_abc_19873_new_n2044_), .B(_abc_19873_new_n2043_), .Y(_abc_19873_new_n2045_));
OR2X2 OR2X2_436 ( .A(_abc_19873_new_n2048_), .B(_abc_19873_new_n2047_), .Y(_abc_19873_new_n2049_));
OR2X2 OR2X2_437 ( .A(_abc_19873_new_n2052_), .B(_abc_19873_new_n2051_), .Y(_abc_19873_new_n2053_));
OR2X2 OR2X2_438 ( .A(_abc_19873_new_n2056_), .B(_abc_19873_new_n2055_), .Y(_abc_19873_new_n2057_));
OR2X2 OR2X2_439 ( .A(_abc_19873_new_n2060_), .B(_abc_19873_new_n2059_), .Y(_abc_19873_new_n2061_));
OR2X2 OR2X2_44 ( .A(_abc_19873_new_n1005_), .B(_abc_19873_new_n1008_), .Y(_abc_19873_new_n1009_));
OR2X2 OR2X2_440 ( .A(_abc_19873_new_n2064_), .B(_abc_19873_new_n2063_), .Y(_abc_19873_new_n2065_));
OR2X2 OR2X2_441 ( .A(_abc_19873_new_n2068_), .B(_abc_19873_new_n2067_), .Y(_abc_19873_new_n2069_));
OR2X2 OR2X2_442 ( .A(_abc_19873_new_n2072_), .B(_abc_19873_new_n2071_), .Y(_abc_19873_new_n2073_));
OR2X2 OR2X2_443 ( .A(_abc_19873_new_n2076_), .B(_abc_19873_new_n2075_), .Y(_abc_19873_new_n2077_));
OR2X2 OR2X2_444 ( .A(_abc_19873_new_n2080_), .B(_abc_19873_new_n2079_), .Y(_abc_19873_new_n2081_));
OR2X2 OR2X2_445 ( .A(_abc_19873_new_n2084_), .B(_abc_19873_new_n2083_), .Y(_abc_19873_new_n2085_));
OR2X2 OR2X2_446 ( .A(_abc_19873_new_n2088_), .B(_abc_19873_new_n2087_), .Y(_abc_19873_new_n2089_));
OR2X2 OR2X2_447 ( .A(_abc_19873_new_n2092_), .B(_abc_19873_new_n2091_), .Y(_abc_19873_new_n2093_));
OR2X2 OR2X2_448 ( .A(_abc_19873_new_n2096_), .B(_abc_19873_new_n2095_), .Y(_abc_19873_new_n2097_));
OR2X2 OR2X2_449 ( .A(_abc_19873_new_n2100_), .B(_abc_19873_new_n2099_), .Y(_abc_19873_new_n2101_));
OR2X2 OR2X2_45 ( .A(_abc_19873_new_n1009_), .B(_abc_19873_new_n1002_), .Y(_abc_19873_new_n1010_));
OR2X2 OR2X2_450 ( .A(_abc_19873_new_n2104_), .B(_abc_19873_new_n2103_), .Y(_abc_19873_new_n2105_));
OR2X2 OR2X2_451 ( .A(_abc_19873_new_n2108_), .B(_abc_19873_new_n2107_), .Y(_abc_19873_new_n2109_));
OR2X2 OR2X2_452 ( .A(_abc_19873_new_n2112_), .B(_abc_19873_new_n2111_), .Y(_abc_19873_new_n2113_));
OR2X2 OR2X2_453 ( .A(_abc_19873_new_n2116_), .B(_abc_19873_new_n2115_), .Y(_abc_19873_new_n2117_));
OR2X2 OR2X2_454 ( .A(_abc_19873_new_n2120_), .B(core_mi_32_), .Y(_abc_19873_new_n2121_));
OR2X2 OR2X2_455 ( .A(_abc_19873_new_n2120_), .B(core_mi_33_), .Y(_abc_19873_new_n2127_));
OR2X2 OR2X2_456 ( .A(_abc_19873_new_n2120_), .B(core_mi_34_), .Y(_abc_19873_new_n2133_));
OR2X2 OR2X2_457 ( .A(_abc_19873_new_n2120_), .B(core_mi_35_), .Y(_abc_19873_new_n2139_));
OR2X2 OR2X2_458 ( .A(_abc_19873_new_n2120_), .B(core_mi_36_), .Y(_abc_19873_new_n2145_));
OR2X2 OR2X2_459 ( .A(_abc_19873_new_n2120_), .B(core_mi_37_), .Y(_abc_19873_new_n2151_));
OR2X2 OR2X2_46 ( .A(_abc_19873_new_n1010_), .B(_abc_19873_new_n997_), .Y(_abc_19873_new_n1011_));
OR2X2 OR2X2_460 ( .A(_abc_19873_new_n2120_), .B(core_mi_38_), .Y(_abc_19873_new_n2157_));
OR2X2 OR2X2_461 ( .A(_abc_19873_new_n2120_), .B(core_mi_39_), .Y(_abc_19873_new_n2163_));
OR2X2 OR2X2_462 ( .A(_abc_19873_new_n2120_), .B(core_mi_40_), .Y(_abc_19873_new_n2169_));
OR2X2 OR2X2_463 ( .A(_abc_19873_new_n2120_), .B(core_mi_41_), .Y(_abc_19873_new_n2175_));
OR2X2 OR2X2_464 ( .A(_abc_19873_new_n2120_), .B(core_mi_42_), .Y(_abc_19873_new_n2181_));
OR2X2 OR2X2_465 ( .A(_abc_19873_new_n2120_), .B(core_mi_43_), .Y(_abc_19873_new_n2187_));
OR2X2 OR2X2_466 ( .A(_abc_19873_new_n2120_), .B(core_mi_44_), .Y(_abc_19873_new_n2193_));
OR2X2 OR2X2_467 ( .A(_abc_19873_new_n2120_), .B(core_mi_45_), .Y(_abc_19873_new_n2199_));
OR2X2 OR2X2_468 ( .A(_abc_19873_new_n2120_), .B(core_mi_46_), .Y(_abc_19873_new_n2205_));
OR2X2 OR2X2_469 ( .A(_abc_19873_new_n2120_), .B(core_mi_47_), .Y(_abc_19873_new_n2211_));
OR2X2 OR2X2_47 ( .A(_abc_19873_new_n1014_), .B(_abc_19873_new_n1015_), .Y(_abc_19873_new_n1016_));
OR2X2 OR2X2_470 ( .A(_abc_19873_new_n2120_), .B(core_mi_48_), .Y(_abc_19873_new_n2217_));
OR2X2 OR2X2_471 ( .A(_abc_19873_new_n2120_), .B(core_mi_49_), .Y(_abc_19873_new_n2223_));
OR2X2 OR2X2_472 ( .A(_abc_19873_new_n2120_), .B(core_mi_50_), .Y(_abc_19873_new_n2229_));
OR2X2 OR2X2_473 ( .A(_abc_19873_new_n2120_), .B(core_mi_51_), .Y(_abc_19873_new_n2235_));
OR2X2 OR2X2_474 ( .A(_abc_19873_new_n2120_), .B(core_mi_52_), .Y(_abc_19873_new_n2241_));
OR2X2 OR2X2_475 ( .A(_abc_19873_new_n2120_), .B(core_mi_53_), .Y(_abc_19873_new_n2247_));
OR2X2 OR2X2_476 ( .A(_abc_19873_new_n2120_), .B(core_mi_54_), .Y(_abc_19873_new_n2253_));
OR2X2 OR2X2_477 ( .A(_abc_19873_new_n2120_), .B(core_mi_55_), .Y(_abc_19873_new_n2259_));
OR2X2 OR2X2_478 ( .A(_abc_19873_new_n2120_), .B(core_mi_56_), .Y(_abc_19873_new_n2265_));
OR2X2 OR2X2_479 ( .A(_abc_19873_new_n2120_), .B(core_mi_57_), .Y(_abc_19873_new_n2271_));
OR2X2 OR2X2_48 ( .A(_abc_19873_new_n1017_), .B(_abc_19873_new_n1018_), .Y(_abc_19873_new_n1019_));
OR2X2 OR2X2_480 ( .A(_abc_19873_new_n2120_), .B(core_mi_58_), .Y(_abc_19873_new_n2277_));
OR2X2 OR2X2_481 ( .A(_abc_19873_new_n2120_), .B(core_mi_59_), .Y(_abc_19873_new_n2283_));
OR2X2 OR2X2_482 ( .A(_abc_19873_new_n2120_), .B(core_mi_60_), .Y(_abc_19873_new_n2289_));
OR2X2 OR2X2_483 ( .A(_abc_19873_new_n2120_), .B(core_mi_61_), .Y(_abc_19873_new_n2295_));
OR2X2 OR2X2_484 ( .A(_abc_19873_new_n2120_), .B(core_mi_62_), .Y(_abc_19873_new_n2301_));
OR2X2 OR2X2_485 ( .A(_abc_19873_new_n2120_), .B(core_mi_63_), .Y(_abc_19873_new_n2307_));
OR2X2 OR2X2_486 ( .A(_abc_19873_new_n2313_), .B(core_mi_0_), .Y(_abc_19873_new_n2314_));
OR2X2 OR2X2_487 ( .A(_abc_19873_new_n2313_), .B(core_mi_1_), .Y(_abc_19873_new_n2319_));
OR2X2 OR2X2_488 ( .A(_abc_19873_new_n2313_), .B(core_mi_2_), .Y(_abc_19873_new_n2324_));
OR2X2 OR2X2_489 ( .A(_abc_19873_new_n2313_), .B(core_mi_3_), .Y(_abc_19873_new_n2329_));
OR2X2 OR2X2_49 ( .A(_abc_19873_new_n1016_), .B(_abc_19873_new_n1019_), .Y(_abc_19873_new_n1020_));
OR2X2 OR2X2_490 ( .A(_abc_19873_new_n2313_), .B(core_mi_4_), .Y(_abc_19873_new_n2334_));
OR2X2 OR2X2_491 ( .A(_abc_19873_new_n2313_), .B(core_mi_5_), .Y(_abc_19873_new_n2339_));
OR2X2 OR2X2_492 ( .A(_abc_19873_new_n2313_), .B(core_mi_6_), .Y(_abc_19873_new_n2344_));
OR2X2 OR2X2_493 ( .A(_abc_19873_new_n2313_), .B(core_mi_7_), .Y(_abc_19873_new_n2349_));
OR2X2 OR2X2_494 ( .A(_abc_19873_new_n2313_), .B(core_mi_8_), .Y(_abc_19873_new_n2354_));
OR2X2 OR2X2_495 ( .A(_abc_19873_new_n2313_), .B(core_mi_9_), .Y(_abc_19873_new_n2359_));
OR2X2 OR2X2_496 ( .A(_abc_19873_new_n2313_), .B(core_mi_10_), .Y(_abc_19873_new_n2364_));
OR2X2 OR2X2_497 ( .A(_abc_19873_new_n2313_), .B(core_mi_11_), .Y(_abc_19873_new_n2369_));
OR2X2 OR2X2_498 ( .A(_abc_19873_new_n2313_), .B(core_mi_12_), .Y(_abc_19873_new_n2374_));
OR2X2 OR2X2_499 ( .A(_abc_19873_new_n2313_), .B(core_mi_13_), .Y(_abc_19873_new_n2379_));
OR2X2 OR2X2_5 ( .A(_abc_19873_new_n910_), .B(_abc_19873_new_n890_), .Y(_abc_19873_new_n911_));
OR2X2 OR2X2_50 ( .A(_abc_19873_new_n1020_), .B(_abc_19873_new_n1013_), .Y(_abc_19873_new_n1021_));
OR2X2 OR2X2_500 ( .A(_abc_19873_new_n2313_), .B(core_mi_14_), .Y(_abc_19873_new_n2384_));
OR2X2 OR2X2_501 ( .A(_abc_19873_new_n2313_), .B(core_mi_15_), .Y(_abc_19873_new_n2389_));
OR2X2 OR2X2_502 ( .A(_abc_19873_new_n2313_), .B(core_mi_16_), .Y(_abc_19873_new_n2394_));
OR2X2 OR2X2_503 ( .A(_abc_19873_new_n2313_), .B(core_mi_17_), .Y(_abc_19873_new_n2399_));
OR2X2 OR2X2_504 ( .A(_abc_19873_new_n2313_), .B(core_mi_18_), .Y(_abc_19873_new_n2404_));
OR2X2 OR2X2_505 ( .A(_abc_19873_new_n2313_), .B(core_mi_19_), .Y(_abc_19873_new_n2409_));
OR2X2 OR2X2_506 ( .A(_abc_19873_new_n2313_), .B(core_mi_20_), .Y(_abc_19873_new_n2414_));
OR2X2 OR2X2_507 ( .A(_abc_19873_new_n2313_), .B(core_mi_21_), .Y(_abc_19873_new_n2419_));
OR2X2 OR2X2_508 ( .A(_abc_19873_new_n2313_), .B(core_mi_22_), .Y(_abc_19873_new_n2424_));
OR2X2 OR2X2_509 ( .A(_abc_19873_new_n2313_), .B(core_mi_23_), .Y(_abc_19873_new_n2429_));
OR2X2 OR2X2_51 ( .A(_abc_19873_new_n1023_), .B(_abc_19873_new_n1024_), .Y(_abc_19873_new_n1025_));
OR2X2 OR2X2_510 ( .A(_abc_19873_new_n2313_), .B(core_mi_24_), .Y(_abc_19873_new_n2434_));
OR2X2 OR2X2_511 ( .A(_abc_19873_new_n2313_), .B(core_mi_25_), .Y(_abc_19873_new_n2439_));
OR2X2 OR2X2_512 ( .A(_abc_19873_new_n2313_), .B(core_mi_26_), .Y(_abc_19873_new_n2444_));
OR2X2 OR2X2_513 ( .A(_abc_19873_new_n2313_), .B(core_mi_27_), .Y(_abc_19873_new_n2449_));
OR2X2 OR2X2_514 ( .A(_abc_19873_new_n2313_), .B(core_mi_28_), .Y(_abc_19873_new_n2454_));
OR2X2 OR2X2_515 ( .A(_abc_19873_new_n2313_), .B(core_mi_29_), .Y(_abc_19873_new_n2459_));
OR2X2 OR2X2_516 ( .A(_abc_19873_new_n2313_), .B(core_mi_30_), .Y(_abc_19873_new_n2464_));
OR2X2 OR2X2_517 ( .A(_abc_19873_new_n2313_), .B(core_mi_31_), .Y(_abc_19873_new_n2469_));
OR2X2 OR2X2_518 ( .A(_abc_19873_new_n2474_), .B(core_key_96_), .Y(_abc_19873_new_n2475_));
OR2X2 OR2X2_519 ( .A(_abc_19873_new_n2474_), .B(core_key_97_), .Y(_abc_19873_new_n2480_));
OR2X2 OR2X2_52 ( .A(_abc_19873_new_n1025_), .B(_abc_19873_new_n1022_), .Y(_abc_19873_new_n1026_));
OR2X2 OR2X2_520 ( .A(_abc_19873_new_n2474_), .B(core_key_98_), .Y(_abc_19873_new_n2485_));
OR2X2 OR2X2_521 ( .A(_abc_19873_new_n2474_), .B(core_key_99_), .Y(_abc_19873_new_n2490_));
OR2X2 OR2X2_522 ( .A(_abc_19873_new_n2474_), .B(core_key_100_), .Y(_abc_19873_new_n2495_));
OR2X2 OR2X2_523 ( .A(_abc_19873_new_n2474_), .B(core_key_101_), .Y(_abc_19873_new_n2500_));
OR2X2 OR2X2_524 ( .A(_abc_19873_new_n2474_), .B(core_key_102_), .Y(_abc_19873_new_n2505_));
OR2X2 OR2X2_525 ( .A(_abc_19873_new_n2474_), .B(core_key_103_), .Y(_abc_19873_new_n2510_));
OR2X2 OR2X2_526 ( .A(_abc_19873_new_n2474_), .B(core_key_104_), .Y(_abc_19873_new_n2515_));
OR2X2 OR2X2_527 ( .A(_abc_19873_new_n2474_), .B(core_key_105_), .Y(_abc_19873_new_n2520_));
OR2X2 OR2X2_528 ( .A(_abc_19873_new_n2474_), .B(core_key_106_), .Y(_abc_19873_new_n2525_));
OR2X2 OR2X2_529 ( .A(_abc_19873_new_n2474_), .B(core_key_107_), .Y(_abc_19873_new_n2530_));
OR2X2 OR2X2_53 ( .A(_abc_19873_new_n1027_), .B(_abc_19873_new_n1028_), .Y(_abc_19873_new_n1029_));
OR2X2 OR2X2_530 ( .A(_abc_19873_new_n2474_), .B(core_key_108_), .Y(_abc_19873_new_n2535_));
OR2X2 OR2X2_531 ( .A(_abc_19873_new_n2474_), .B(core_key_109_), .Y(_abc_19873_new_n2540_));
OR2X2 OR2X2_532 ( .A(_abc_19873_new_n2474_), .B(core_key_110_), .Y(_abc_19873_new_n2545_));
OR2X2 OR2X2_533 ( .A(_abc_19873_new_n2474_), .B(core_key_111_), .Y(_abc_19873_new_n2550_));
OR2X2 OR2X2_534 ( .A(_abc_19873_new_n2474_), .B(core_key_112_), .Y(_abc_19873_new_n2555_));
OR2X2 OR2X2_535 ( .A(_abc_19873_new_n2474_), .B(core_key_113_), .Y(_abc_19873_new_n2560_));
OR2X2 OR2X2_536 ( .A(_abc_19873_new_n2474_), .B(core_key_114_), .Y(_abc_19873_new_n2565_));
OR2X2 OR2X2_537 ( .A(_abc_19873_new_n2474_), .B(core_key_115_), .Y(_abc_19873_new_n2570_));
OR2X2 OR2X2_538 ( .A(_abc_19873_new_n2474_), .B(core_key_116_), .Y(_abc_19873_new_n2575_));
OR2X2 OR2X2_539 ( .A(_abc_19873_new_n2474_), .B(core_key_117_), .Y(_abc_19873_new_n2580_));
OR2X2 OR2X2_54 ( .A(_abc_19873_new_n1030_), .B(_abc_19873_new_n1031_), .Y(_abc_19873_new_n1032_));
OR2X2 OR2X2_540 ( .A(_abc_19873_new_n2474_), .B(core_key_118_), .Y(_abc_19873_new_n2585_));
OR2X2 OR2X2_541 ( .A(_abc_19873_new_n2474_), .B(core_key_119_), .Y(_abc_19873_new_n2590_));
OR2X2 OR2X2_542 ( .A(_abc_19873_new_n2474_), .B(core_key_120_), .Y(_abc_19873_new_n2595_));
OR2X2 OR2X2_543 ( .A(_abc_19873_new_n2474_), .B(core_key_121_), .Y(_abc_19873_new_n2600_));
OR2X2 OR2X2_544 ( .A(_abc_19873_new_n2474_), .B(core_key_122_), .Y(_abc_19873_new_n2605_));
OR2X2 OR2X2_545 ( .A(_abc_19873_new_n2474_), .B(core_key_123_), .Y(_abc_19873_new_n2610_));
OR2X2 OR2X2_546 ( .A(_abc_19873_new_n2474_), .B(core_key_124_), .Y(_abc_19873_new_n2615_));
OR2X2 OR2X2_547 ( .A(_abc_19873_new_n2474_), .B(core_key_125_), .Y(_abc_19873_new_n2620_));
OR2X2 OR2X2_548 ( .A(_abc_19873_new_n2474_), .B(core_key_126_), .Y(_abc_19873_new_n2625_));
OR2X2 OR2X2_549 ( .A(_abc_19873_new_n2474_), .B(core_key_127_), .Y(_abc_19873_new_n2630_));
OR2X2 OR2X2_55 ( .A(_abc_19873_new_n1029_), .B(_abc_19873_new_n1032_), .Y(_abc_19873_new_n1033_));
OR2X2 OR2X2_550 ( .A(_abc_19873_new_n2635_), .B(core_key_64_), .Y(_abc_19873_new_n2636_));
OR2X2 OR2X2_551 ( .A(_abc_19873_new_n2635_), .B(core_key_65_), .Y(_abc_19873_new_n2641_));
OR2X2 OR2X2_552 ( .A(_abc_19873_new_n2635_), .B(core_key_66_), .Y(_abc_19873_new_n2646_));
OR2X2 OR2X2_553 ( .A(_abc_19873_new_n2635_), .B(core_key_67_), .Y(_abc_19873_new_n2651_));
OR2X2 OR2X2_554 ( .A(_abc_19873_new_n2635_), .B(core_key_68_), .Y(_abc_19873_new_n2656_));
OR2X2 OR2X2_555 ( .A(_abc_19873_new_n2635_), .B(core_key_69_), .Y(_abc_19873_new_n2661_));
OR2X2 OR2X2_556 ( .A(_abc_19873_new_n2635_), .B(core_key_70_), .Y(_abc_19873_new_n2666_));
OR2X2 OR2X2_557 ( .A(_abc_19873_new_n2635_), .B(core_key_71_), .Y(_abc_19873_new_n2671_));
OR2X2 OR2X2_558 ( .A(_abc_19873_new_n2635_), .B(core_key_72_), .Y(_abc_19873_new_n2676_));
OR2X2 OR2X2_559 ( .A(_abc_19873_new_n2635_), .B(core_key_73_), .Y(_abc_19873_new_n2681_));
OR2X2 OR2X2_56 ( .A(_abc_19873_new_n1033_), .B(_abc_19873_new_n1026_), .Y(_abc_19873_new_n1034_));
OR2X2 OR2X2_560 ( .A(_abc_19873_new_n2635_), .B(core_key_74_), .Y(_abc_19873_new_n2686_));
OR2X2 OR2X2_561 ( .A(_abc_19873_new_n2635_), .B(core_key_75_), .Y(_abc_19873_new_n2691_));
OR2X2 OR2X2_562 ( .A(_abc_19873_new_n2635_), .B(core_key_76_), .Y(_abc_19873_new_n2696_));
OR2X2 OR2X2_563 ( .A(_abc_19873_new_n2635_), .B(core_key_77_), .Y(_abc_19873_new_n2701_));
OR2X2 OR2X2_564 ( .A(_abc_19873_new_n2635_), .B(core_key_78_), .Y(_abc_19873_new_n2706_));
OR2X2 OR2X2_565 ( .A(_abc_19873_new_n2635_), .B(core_key_79_), .Y(_abc_19873_new_n2711_));
OR2X2 OR2X2_566 ( .A(_abc_19873_new_n2635_), .B(core_key_80_), .Y(_abc_19873_new_n2716_));
OR2X2 OR2X2_567 ( .A(_abc_19873_new_n2635_), .B(core_key_81_), .Y(_abc_19873_new_n2721_));
OR2X2 OR2X2_568 ( .A(_abc_19873_new_n2635_), .B(core_key_82_), .Y(_abc_19873_new_n2726_));
OR2X2 OR2X2_569 ( .A(_abc_19873_new_n2635_), .B(core_key_83_), .Y(_abc_19873_new_n2731_));
OR2X2 OR2X2_57 ( .A(_abc_19873_new_n1034_), .B(_abc_19873_new_n1021_), .Y(_abc_19873_new_n1035_));
OR2X2 OR2X2_570 ( .A(_abc_19873_new_n2635_), .B(core_key_84_), .Y(_abc_19873_new_n2736_));
OR2X2 OR2X2_571 ( .A(_abc_19873_new_n2635_), .B(core_key_85_), .Y(_abc_19873_new_n2741_));
OR2X2 OR2X2_572 ( .A(_abc_19873_new_n2635_), .B(core_key_86_), .Y(_abc_19873_new_n2746_));
OR2X2 OR2X2_573 ( .A(_abc_19873_new_n2635_), .B(core_key_87_), .Y(_abc_19873_new_n2751_));
OR2X2 OR2X2_574 ( .A(_abc_19873_new_n2635_), .B(core_key_88_), .Y(_abc_19873_new_n2756_));
OR2X2 OR2X2_575 ( .A(_abc_19873_new_n2635_), .B(core_key_89_), .Y(_abc_19873_new_n2761_));
OR2X2 OR2X2_576 ( .A(_abc_19873_new_n2635_), .B(core_key_90_), .Y(_abc_19873_new_n2766_));
OR2X2 OR2X2_577 ( .A(_abc_19873_new_n2635_), .B(core_key_91_), .Y(_abc_19873_new_n2771_));
OR2X2 OR2X2_578 ( .A(_abc_19873_new_n2635_), .B(core_key_92_), .Y(_abc_19873_new_n2776_));
OR2X2 OR2X2_579 ( .A(_abc_19873_new_n2635_), .B(core_key_93_), .Y(_abc_19873_new_n2781_));
OR2X2 OR2X2_58 ( .A(_abc_19873_new_n994_), .B(_abc_19873_new_n1037_), .Y(_abc_19873_new_n1038_));
OR2X2 OR2X2_580 ( .A(_abc_19873_new_n2635_), .B(core_key_94_), .Y(_abc_19873_new_n2786_));
OR2X2 OR2X2_581 ( .A(_abc_19873_new_n2635_), .B(core_key_95_), .Y(_abc_19873_new_n2791_));
OR2X2 OR2X2_582 ( .A(_abc_19873_new_n2796_), .B(core_key_32_), .Y(_abc_19873_new_n2797_));
OR2X2 OR2X2_583 ( .A(_abc_19873_new_n2796_), .B(core_key_33_), .Y(_abc_19873_new_n2802_));
OR2X2 OR2X2_584 ( .A(_abc_19873_new_n2796_), .B(core_key_34_), .Y(_abc_19873_new_n2807_));
OR2X2 OR2X2_585 ( .A(_abc_19873_new_n2796_), .B(core_key_35_), .Y(_abc_19873_new_n2812_));
OR2X2 OR2X2_586 ( .A(_abc_19873_new_n2796_), .B(core_key_36_), .Y(_abc_19873_new_n2817_));
OR2X2 OR2X2_587 ( .A(_abc_19873_new_n2796_), .B(core_key_37_), .Y(_abc_19873_new_n2822_));
OR2X2 OR2X2_588 ( .A(_abc_19873_new_n2796_), .B(core_key_38_), .Y(_abc_19873_new_n2827_));
OR2X2 OR2X2_589 ( .A(_abc_19873_new_n2796_), .B(core_key_39_), .Y(_abc_19873_new_n2832_));
OR2X2 OR2X2_59 ( .A(_abc_19873_new_n1038_), .B(_abc_19873_new_n1018_), .Y(_abc_19873_new_n1039_));
OR2X2 OR2X2_590 ( .A(_abc_19873_new_n2796_), .B(core_key_40_), .Y(_abc_19873_new_n2837_));
OR2X2 OR2X2_591 ( .A(_abc_19873_new_n2796_), .B(core_key_41_), .Y(_abc_19873_new_n2842_));
OR2X2 OR2X2_592 ( .A(_abc_19873_new_n2796_), .B(core_key_42_), .Y(_abc_19873_new_n2847_));
OR2X2 OR2X2_593 ( .A(_abc_19873_new_n2796_), .B(core_key_43_), .Y(_abc_19873_new_n2852_));
OR2X2 OR2X2_594 ( .A(_abc_19873_new_n2796_), .B(core_key_44_), .Y(_abc_19873_new_n2857_));
OR2X2 OR2X2_595 ( .A(_abc_19873_new_n2796_), .B(core_key_45_), .Y(_abc_19873_new_n2862_));
OR2X2 OR2X2_596 ( .A(_abc_19873_new_n2796_), .B(core_key_46_), .Y(_abc_19873_new_n2867_));
OR2X2 OR2X2_597 ( .A(_abc_19873_new_n2796_), .B(core_key_47_), .Y(_abc_19873_new_n2872_));
OR2X2 OR2X2_598 ( .A(_abc_19873_new_n2796_), .B(core_key_48_), .Y(_abc_19873_new_n2877_));
OR2X2 OR2X2_599 ( .A(_abc_19873_new_n2796_), .B(core_key_49_), .Y(_abc_19873_new_n2882_));
OR2X2 OR2X2_6 ( .A(_abc_19873_new_n917_), .B(_abc_19873_new_n920_), .Y(_abc_19873_new_n921_));
OR2X2 OR2X2_60 ( .A(_abc_19873_new_n1040_), .B(_abc_19873_new_n1041_), .Y(_abc_19873_new_n1042_));
OR2X2 OR2X2_600 ( .A(_abc_19873_new_n2796_), .B(core_key_50_), .Y(_abc_19873_new_n2887_));
OR2X2 OR2X2_601 ( .A(_abc_19873_new_n2796_), .B(core_key_51_), .Y(_abc_19873_new_n2892_));
OR2X2 OR2X2_602 ( .A(_abc_19873_new_n2796_), .B(core_key_52_), .Y(_abc_19873_new_n2897_));
OR2X2 OR2X2_603 ( .A(_abc_19873_new_n2796_), .B(core_key_53_), .Y(_abc_19873_new_n2902_));
OR2X2 OR2X2_604 ( .A(_abc_19873_new_n2796_), .B(core_key_54_), .Y(_abc_19873_new_n2907_));
OR2X2 OR2X2_605 ( .A(_abc_19873_new_n2796_), .B(core_key_55_), .Y(_abc_19873_new_n2912_));
OR2X2 OR2X2_606 ( .A(_abc_19873_new_n2796_), .B(core_key_56_), .Y(_abc_19873_new_n2917_));
OR2X2 OR2X2_607 ( .A(_abc_19873_new_n2796_), .B(core_key_57_), .Y(_abc_19873_new_n2922_));
OR2X2 OR2X2_608 ( .A(_abc_19873_new_n2796_), .B(core_key_58_), .Y(_abc_19873_new_n2927_));
OR2X2 OR2X2_609 ( .A(_abc_19873_new_n2796_), .B(core_key_59_), .Y(_abc_19873_new_n2932_));
OR2X2 OR2X2_61 ( .A(_abc_19873_new_n1039_), .B(_abc_19873_new_n1042_), .Y(_abc_19873_new_n1043_));
OR2X2 OR2X2_610 ( .A(_abc_19873_new_n2796_), .B(core_key_60_), .Y(_abc_19873_new_n2937_));
OR2X2 OR2X2_611 ( .A(_abc_19873_new_n2796_), .B(core_key_61_), .Y(_abc_19873_new_n2942_));
OR2X2 OR2X2_612 ( .A(_abc_19873_new_n2796_), .B(core_key_62_), .Y(_abc_19873_new_n2947_));
OR2X2 OR2X2_613 ( .A(_abc_19873_new_n2796_), .B(core_key_63_), .Y(_abc_19873_new_n2952_));
OR2X2 OR2X2_614 ( .A(_abc_19873_new_n2957_), .B(core_key_0_), .Y(_abc_19873_new_n2958_));
OR2X2 OR2X2_615 ( .A(_abc_19873_new_n2957_), .B(core_key_1_), .Y(_abc_19873_new_n2963_));
OR2X2 OR2X2_616 ( .A(_abc_19873_new_n2957_), .B(core_key_2_), .Y(_abc_19873_new_n2968_));
OR2X2 OR2X2_617 ( .A(_abc_19873_new_n2957_), .B(core_key_3_), .Y(_abc_19873_new_n2973_));
OR2X2 OR2X2_618 ( .A(_abc_19873_new_n2957_), .B(core_key_4_), .Y(_abc_19873_new_n2978_));
OR2X2 OR2X2_619 ( .A(_abc_19873_new_n2957_), .B(core_key_5_), .Y(_abc_19873_new_n2983_));
OR2X2 OR2X2_62 ( .A(_abc_19873_new_n1045_), .B(_abc_19873_new_n1046_), .Y(_abc_19873_new_n1047_));
OR2X2 OR2X2_620 ( .A(_abc_19873_new_n2957_), .B(core_key_6_), .Y(_abc_19873_new_n2988_));
OR2X2 OR2X2_621 ( .A(_abc_19873_new_n2957_), .B(core_key_7_), .Y(_abc_19873_new_n2993_));
OR2X2 OR2X2_622 ( .A(_abc_19873_new_n2957_), .B(core_key_8_), .Y(_abc_19873_new_n2998_));
OR2X2 OR2X2_623 ( .A(_abc_19873_new_n2957_), .B(core_key_9_), .Y(_abc_19873_new_n3003_));
OR2X2 OR2X2_624 ( .A(_abc_19873_new_n2957_), .B(core_key_10_), .Y(_abc_19873_new_n3008_));
OR2X2 OR2X2_625 ( .A(_abc_19873_new_n2957_), .B(core_key_11_), .Y(_abc_19873_new_n3013_));
OR2X2 OR2X2_626 ( .A(_abc_19873_new_n2957_), .B(core_key_12_), .Y(_abc_19873_new_n3018_));
OR2X2 OR2X2_627 ( .A(_abc_19873_new_n2957_), .B(core_key_13_), .Y(_abc_19873_new_n3023_));
OR2X2 OR2X2_628 ( .A(_abc_19873_new_n2957_), .B(core_key_14_), .Y(_abc_19873_new_n3028_));
OR2X2 OR2X2_629 ( .A(_abc_19873_new_n2957_), .B(core_key_15_), .Y(_abc_19873_new_n3033_));
OR2X2 OR2X2_63 ( .A(_abc_19873_new_n1047_), .B(_abc_19873_new_n1044_), .Y(_abc_19873_new_n1048_));
OR2X2 OR2X2_630 ( .A(_abc_19873_new_n2957_), .B(core_key_16_), .Y(_abc_19873_new_n3038_));
OR2X2 OR2X2_631 ( .A(_abc_19873_new_n2957_), .B(core_key_17_), .Y(_abc_19873_new_n3043_));
OR2X2 OR2X2_632 ( .A(_abc_19873_new_n2957_), .B(core_key_18_), .Y(_abc_19873_new_n3048_));
OR2X2 OR2X2_633 ( .A(_abc_19873_new_n2957_), .B(core_key_19_), .Y(_abc_19873_new_n3053_));
OR2X2 OR2X2_634 ( .A(_abc_19873_new_n2957_), .B(core_key_20_), .Y(_abc_19873_new_n3058_));
OR2X2 OR2X2_635 ( .A(_abc_19873_new_n2957_), .B(core_key_21_), .Y(_abc_19873_new_n3063_));
OR2X2 OR2X2_636 ( .A(_abc_19873_new_n2957_), .B(core_key_22_), .Y(_abc_19873_new_n3068_));
OR2X2 OR2X2_637 ( .A(_abc_19873_new_n2957_), .B(core_key_23_), .Y(_abc_19873_new_n3073_));
OR2X2 OR2X2_638 ( .A(_abc_19873_new_n2957_), .B(core_key_24_), .Y(_abc_19873_new_n3078_));
OR2X2 OR2X2_639 ( .A(_abc_19873_new_n2957_), .B(core_key_25_), .Y(_abc_19873_new_n3083_));
OR2X2 OR2X2_64 ( .A(_abc_19873_new_n1043_), .B(_abc_19873_new_n1048_), .Y(_abc_19873_new_n1049_));
OR2X2 OR2X2_640 ( .A(_abc_19873_new_n2957_), .B(core_key_26_), .Y(_abc_19873_new_n3088_));
OR2X2 OR2X2_641 ( .A(_abc_19873_new_n2957_), .B(core_key_27_), .Y(_abc_19873_new_n3093_));
OR2X2 OR2X2_642 ( .A(_abc_19873_new_n2957_), .B(core_key_28_), .Y(_abc_19873_new_n3098_));
OR2X2 OR2X2_643 ( .A(_abc_19873_new_n2957_), .B(core_key_29_), .Y(_abc_19873_new_n3103_));
OR2X2 OR2X2_644 ( .A(_abc_19873_new_n2957_), .B(core_key_30_), .Y(_abc_19873_new_n3108_));
OR2X2 OR2X2_645 ( .A(_abc_19873_new_n2957_), .B(core_key_31_), .Y(_abc_19873_new_n3113_));
OR2X2 OR2X2_646 ( .A(_abc_19873_new_n3121_), .B(_abc_19873_new_n3119_), .Y(_abc_19873_new_n3122_));
OR2X2 OR2X2_647 ( .A(_abc_19873_new_n3126_), .B(_abc_19873_new_n3125_), .Y(_abc_19873_new_n3127_));
OR2X2 OR2X2_648 ( .A(_abc_19873_new_n3127_), .B(_abc_19873_new_n3124_), .Y(_0param_reg_7_0__1_));
OR2X2 OR2X2_649 ( .A(_abc_19873_new_n3129_), .B(_abc_19873_new_n3130_), .Y(_abc_19873_new_n3131_));
OR2X2 OR2X2_65 ( .A(_abc_19873_new_n1050_), .B(_abc_19873_new_n1051_), .Y(_abc_19873_new_n1052_));
OR2X2 OR2X2_650 ( .A(_abc_19873_new_n3134_), .B(_abc_19873_new_n3133_), .Y(_abc_19873_new_n3135_));
OR2X2 OR2X2_651 ( .A(_abc_19873_new_n3138_), .B(_abc_19873_new_n3137_), .Y(_abc_19873_new_n3139_));
OR2X2 OR2X2_652 ( .A(_abc_19873_new_n3142_), .B(_abc_19873_new_n3141_), .Y(_abc_19873_new_n3143_));
OR2X2 OR2X2_653 ( .A(_abc_19873_new_n3146_), .B(_abc_19873_new_n3125_), .Y(_abc_19873_new_n3147_));
OR2X2 OR2X2_654 ( .A(_abc_19873_new_n3147_), .B(_abc_19873_new_n3145_), .Y(_0param_reg_7_0__6_));
OR2X2 OR2X2_655 ( .A(_abc_19873_new_n3150_), .B(_abc_19873_new_n3149_), .Y(_abc_19873_new_n3151_));
OR2X2 OR2X2_656 ( .A(_abc_19873_new_n3162_), .B(core_long), .Y(_abc_19873_new_n3165_));
OR2X2 OR2X2_657 ( .A(core__abc_22172_new_n1138_), .B(core__abc_22172_new_n1136_), .Y(core__abc_22172_new_n1139_));
OR2X2 OR2X2_658 ( .A(core__abc_22172_new_n1141_), .B(core__abc_22172_new_n1143_), .Y(core__abc_22172_new_n1144_));
OR2X2 OR2X2_659 ( .A(core__abc_22172_new_n1134_), .B(core__abc_22172_new_n1131_), .Y(core__abc_22172_new_n1146_));
OR2X2 OR2X2_66 ( .A(_abc_19873_new_n1053_), .B(_abc_19873_new_n1054_), .Y(_abc_19873_new_n1055_));
OR2X2 OR2X2_660 ( .A(core__abc_22172_new_n1147_), .B(core_loop_ctr_reg_2_), .Y(core__abc_22172_new_n1150_));
OR2X2 OR2X2_661 ( .A(core__abc_22172_new_n1136_), .B(core__abc_22172_new_n1152_), .Y(core__abc_22172_new_n1153_));
OR2X2 OR2X2_662 ( .A(core__abc_22172_new_n1156_), .B(core__abc_22172_new_n1157_), .Y(core__abc_22172_new_n1158_));
OR2X2 OR2X2_663 ( .A(core__abc_22172_new_n1158_), .B(core_loop_ctr_reg_0_), .Y(core__abc_22172_new_n1161_));
OR2X2 OR2X2_664 ( .A(core_siphash_ctrl_reg_3_), .B(core_siphash_ctrl_reg_6_), .Y(core__abc_22172_new_n1166_));
OR2X2 OR2X2_665 ( .A(core_siphash_word1_we), .B(core_siphash_ctrl_reg_1_), .Y(core__abc_22172_new_n1170_));
OR2X2 OR2X2_666 ( .A(core__abc_22172_new_n1167_), .B(core__abc_22172_new_n1174_), .Y(core__abc_22172_new_n1175_));
OR2X2 OR2X2_667 ( .A(core__abc_22172_new_n1184_), .B(core__abc_22172_new_n1182_), .Y(core__abc_22172_new_n1185_));
OR2X2 OR2X2_668 ( .A(core__abc_22172_new_n1182_), .B(core__abc_22172_new_n1189_), .Y(core__abc_22172_new_n1190_));
OR2X2 OR2X2_669 ( .A(core__abc_22172_new_n1192_), .B(core__abc_22172_new_n1193_), .Y(core__abc_22172_new_n1194_));
OR2X2 OR2X2_67 ( .A(_abc_19873_new_n1056_), .B(_abc_19873_new_n1057_), .Y(_abc_19873_new_n1058_));
OR2X2 OR2X2_670 ( .A(core__abc_22172_new_n1194_), .B(core_loop_ctr_reg_0_), .Y(core__abc_22172_new_n1197_));
OR2X2 OR2X2_671 ( .A(core__abc_22172_new_n1180_), .B(core__abc_22172_new_n1177_), .Y(core__abc_22172_new_n1201_));
OR2X2 OR2X2_672 ( .A(core__abc_22172_new_n1203_), .B(core_loop_ctr_reg_2_), .Y(core__abc_22172_new_n1204_));
OR2X2 OR2X2_673 ( .A(core__abc_22172_new_n1202_), .B(core__abc_22172_new_n1205_), .Y(core__abc_22172_new_n1206_));
OR2X2 OR2X2_674 ( .A(core__abc_22172_new_n1207_), .B(core__abc_22172_new_n1208_), .Y(core__abc_22172_new_n1209_));
OR2X2 OR2X2_675 ( .A(core__abc_22172_new_n1214_), .B(core__abc_22172_new_n1215_), .Y(core__abc_22172_new_n1216_));
OR2X2 OR2X2_676 ( .A(core__abc_22172_new_n1166_), .B(core_siphash_ctrl_reg_4_), .Y(core__abc_22172_new_n1217_));
OR2X2 OR2X2_677 ( .A(core__abc_22172_new_n1212_), .B(core__abc_22172_new_n1220_), .Y(core__abc_22172_new_n1221_));
OR2X2 OR2X2_678 ( .A(core__abc_22172_new_n1175_), .B(core__abc_22172_new_n1221_), .Y(core__abc_22172_new_n1222_));
OR2X2 OR2X2_679 ( .A(core_initalize), .B(core_compress), .Y(core__abc_22172_new_n1224_));
OR2X2 OR2X2_68 ( .A(_abc_19873_new_n1055_), .B(_abc_19873_new_n1058_), .Y(_abc_19873_new_n1059_));
OR2X2 OR2X2_680 ( .A(core__abc_22172_new_n1224_), .B(core_finalize), .Y(core__abc_22172_new_n1225_));
OR2X2 OR2X2_681 ( .A(core__abc_22172_new_n1223_), .B(core__abc_22172_new_n1226_), .Y(core__abc_22172_new_n1227_));
OR2X2 OR2X2_682 ( .A(core__abc_22172_new_n1233_), .B(core__abc_22172_new_n1234_), .Y(core__abc_22172_new_n1235_));
OR2X2 OR2X2_683 ( .A(core__abc_22172_new_n1235_), .B(core__abc_22172_new_n1231_), .Y(core__abc_22172_new_n1236_));
OR2X2 OR2X2_684 ( .A(core__abc_22172_new_n1239_), .B(core__abc_22172_new_n1238_), .Y(core__abc_22172_new_n1240_));
OR2X2 OR2X2_685 ( .A(core__abc_22172_new_n1237_), .B(core__abc_22172_new_n1240_), .Y(core__abc_22172_new_n1241_));
OR2X2 OR2X2_686 ( .A(core__abc_22172_new_n1229_), .B(core__abc_22172_new_n1241_), .Y(core__abc_15204_auto_fsm_map_cc_170_map_fsm_1439_0_));
OR2X2 OR2X2_687 ( .A(core__abc_22172_new_n1245_), .B(core__abc_22172_new_n1243_), .Y(core__abc_15204_auto_fsm_map_cc_170_map_fsm_1439_3_));
OR2X2 OR2X2_688 ( .A(core__abc_22172_new_n1247_), .B(core__abc_22172_new_n1249_), .Y(core__abc_15204_auto_fsm_map_cc_170_map_fsm_1439_4_));
OR2X2 OR2X2_689 ( .A(core__abc_22172_new_n1251_), .B(core__abc_22172_new_n1254_), .Y(core__abc_15204_auto_fsm_map_cc_170_map_fsm_1439_6_));
OR2X2 OR2X2_69 ( .A(_abc_19873_new_n1059_), .B(_abc_19873_new_n1052_), .Y(_abc_19873_new_n1060_));
OR2X2 OR2X2_690 ( .A(core_v1_reg_0_), .B(core_v0_reg_0_), .Y(core__abc_22172_new_n1257_));
OR2X2 OR2X2_691 ( .A(core__abc_22172_new_n1263_), .B(core__abc_22172_new_n1264_), .Y(core__abc_22172_new_n1265_));
OR2X2 OR2X2_692 ( .A(core__abc_22172_new_n1266_), .B(core__abc_22172_new_n1260_), .Y(core__abc_22172_new_n1267_));
OR2X2 OR2X2_693 ( .A(core__abc_22172_new_n1268_), .B(core__abc_22172_new_n1265_), .Y(core__abc_22172_new_n1269_));
OR2X2 OR2X2_694 ( .A(core__abc_22172_new_n1270_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n1271_));
OR2X2 OR2X2_695 ( .A(core_siphash_word1_we), .B(core_siphash_word_64_), .Y(core__abc_22172_new_n1272_));
OR2X2 OR2X2_696 ( .A(core_v1_reg_1_), .B(core_v0_reg_1_), .Y(core__abc_22172_new_n1275_));
OR2X2 OR2X2_697 ( .A(core__abc_22172_new_n1282_), .B(core__abc_22172_new_n1279_), .Y(core__abc_22172_new_n1283_));
OR2X2 OR2X2_698 ( .A(core__abc_22172_new_n1284_), .B(core__abc_22172_new_n1278_), .Y(core__abc_22172_new_n1285_));
OR2X2 OR2X2_699 ( .A(core__abc_22172_new_n1288_), .B(core__abc_22172_new_n1276_), .Y(core__abc_22172_new_n1289_));
OR2X2 OR2X2_7 ( .A(_abc_19873_new_n921_), .B(_abc_19873_new_n913_), .Y(_abc_19873_new_n922_));
OR2X2 OR2X2_70 ( .A(_abc_19873_new_n1049_), .B(_abc_19873_new_n1060_), .Y(_abc_19873_new_n1061_));
OR2X2 OR2X2_700 ( .A(core__abc_22172_new_n1289_), .B(core__abc_22172_new_n1283_), .Y(core__abc_22172_new_n1290_));
OR2X2 OR2X2_701 ( .A(core__abc_22172_new_n1291_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n1292_));
OR2X2 OR2X2_702 ( .A(core_siphash_word1_we), .B(core_siphash_word_65_), .Y(core__abc_22172_new_n1293_));
OR2X2 OR2X2_703 ( .A(core_v1_reg_2_), .B(core_v0_reg_2_), .Y(core__abc_22172_new_n1298_));
OR2X2 OR2X2_704 ( .A(core__abc_22172_new_n1304_), .B(core__abc_22172_new_n1301_), .Y(core__abc_22172_new_n1305_));
OR2X2 OR2X2_705 ( .A(core__abc_22172_new_n1307_), .B(core__abc_22172_new_n1308_), .Y(core__abc_22172_new_n1309_));
OR2X2 OR2X2_706 ( .A(core__abc_22172_new_n1309_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n1310_));
OR2X2 OR2X2_707 ( .A(core_siphash_word1_we), .B(core_siphash_word_66_), .Y(core__abc_22172_new_n1311_));
OR2X2 OR2X2_708 ( .A(core_v1_reg_3_), .B(core_v0_reg_3_), .Y(core__abc_22172_new_n1314_));
OR2X2 OR2X2_709 ( .A(core__abc_22172_new_n1321_), .B(core__abc_22172_new_n1318_), .Y(core__abc_22172_new_n1322_));
OR2X2 OR2X2_71 ( .A(_abc_19873_new_n1063_), .B(_abc_19873_new_n1064_), .Y(_abc_19873_new_n1065_));
OR2X2 OR2X2_710 ( .A(core__abc_22172_new_n1323_), .B(core__abc_22172_new_n1317_), .Y(core__abc_22172_new_n1324_));
OR2X2 OR2X2_711 ( .A(core__abc_22172_new_n1325_), .B(core__abc_22172_new_n1322_), .Y(core__abc_22172_new_n1326_));
OR2X2 OR2X2_712 ( .A(core__abc_22172_new_n1327_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n1328_));
OR2X2 OR2X2_713 ( .A(core_siphash_word1_we), .B(core_siphash_word_67_), .Y(core__abc_22172_new_n1329_));
OR2X2 OR2X2_714 ( .A(core_v1_reg_4_), .B(core_v0_reg_4_), .Y(core__abc_22172_new_n1332_));
OR2X2 OR2X2_715 ( .A(core__abc_22172_new_n1339_), .B(core__abc_22172_new_n1336_), .Y(core__abc_22172_new_n1340_));
OR2X2 OR2X2_716 ( .A(core__abc_22172_new_n1341_), .B(core__abc_22172_new_n1335_), .Y(core__abc_22172_new_n1342_));
OR2X2 OR2X2_717 ( .A(core__abc_22172_new_n1343_), .B(core__abc_22172_new_n1340_), .Y(core__abc_22172_new_n1344_));
OR2X2 OR2X2_718 ( .A(core__abc_22172_new_n1345_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n1346_));
OR2X2 OR2X2_719 ( .A(core_siphash_word1_we), .B(core_siphash_word_68_), .Y(core__abc_22172_new_n1347_));
OR2X2 OR2X2_72 ( .A(_abc_19873_new_n1066_), .B(_abc_19873_new_n1067_), .Y(_abc_19873_new_n1068_));
OR2X2 OR2X2_720 ( .A(core_v1_reg_5_), .B(core_v0_reg_5_), .Y(core__abc_22172_new_n1350_));
OR2X2 OR2X2_721 ( .A(core__abc_22172_new_n1360_), .B(core__abc_22172_new_n1353_), .Y(core__abc_22172_new_n1361_));
OR2X2 OR2X2_722 ( .A(core__abc_22172_new_n1363_), .B(core__abc_22172_new_n1362_), .Y(core__abc_22172_new_n1364_));
OR2X2 OR2X2_723 ( .A(core__abc_22172_new_n1365_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n1366_));
OR2X2 OR2X2_724 ( .A(core_siphash_word1_we), .B(core_siphash_word_69_), .Y(core__abc_22172_new_n1367_));
OR2X2 OR2X2_725 ( .A(core_v1_reg_6_), .B(core_v0_reg_6_), .Y(core__abc_22172_new_n1370_));
OR2X2 OR2X2_726 ( .A(core__abc_22172_new_n1377_), .B(core__abc_22172_new_n1374_), .Y(core__abc_22172_new_n1378_));
OR2X2 OR2X2_727 ( .A(core__abc_22172_new_n1379_), .B(core__abc_22172_new_n1373_), .Y(core__abc_22172_new_n1380_));
OR2X2 OR2X2_728 ( .A(core__abc_22172_new_n1381_), .B(core__abc_22172_new_n1378_), .Y(core__abc_22172_new_n1382_));
OR2X2 OR2X2_729 ( .A(core__abc_22172_new_n1383_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n1384_));
OR2X2 OR2X2_73 ( .A(_abc_19873_new_n1065_), .B(_abc_19873_new_n1068_), .Y(_abc_19873_new_n1069_));
OR2X2 OR2X2_730 ( .A(core_siphash_word1_we), .B(core_siphash_word_70_), .Y(core__abc_22172_new_n1385_));
OR2X2 OR2X2_731 ( .A(core_v1_reg_7_), .B(core_v0_reg_7_), .Y(core__abc_22172_new_n1388_));
OR2X2 OR2X2_732 ( .A(core__abc_22172_new_n1398_), .B(core__abc_22172_new_n1391_), .Y(core__abc_22172_new_n1399_));
OR2X2 OR2X2_733 ( .A(core__abc_22172_new_n1401_), .B(core__abc_22172_new_n1400_), .Y(core__abc_22172_new_n1402_));
OR2X2 OR2X2_734 ( .A(core__abc_22172_new_n1403_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n1404_));
OR2X2 OR2X2_735 ( .A(core_siphash_word1_we), .B(core_siphash_word_71_), .Y(core__abc_22172_new_n1405_));
OR2X2 OR2X2_736 ( .A(core_v1_reg_8_), .B(core_v0_reg_8_), .Y(core__abc_22172_new_n1408_));
OR2X2 OR2X2_737 ( .A(core_v2_reg_8_), .B(core_v3_reg_8_), .Y(core__abc_22172_new_n1414_));
OR2X2 OR2X2_738 ( .A(core__abc_22172_new_n1411_), .B(core__abc_22172_new_n1415_), .Y(core__abc_22172_new_n1416_));
OR2X2 OR2X2_739 ( .A(core__abc_22172_new_n1417_), .B(core__abc_22172_new_n1418_), .Y(core__abc_22172_new_n1419_));
OR2X2 OR2X2_74 ( .A(_abc_19873_new_n1070_), .B(_abc_19873_new_n1071_), .Y(_abc_19873_new_n1072_));
OR2X2 OR2X2_740 ( .A(core__abc_22172_new_n1420_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n1421_));
OR2X2 OR2X2_741 ( .A(core_siphash_word1_we), .B(core_siphash_word_72_), .Y(core__abc_22172_new_n1422_));
OR2X2 OR2X2_742 ( .A(core_v1_reg_9_), .B(core_v0_reg_9_), .Y(core__abc_22172_new_n1425_));
OR2X2 OR2X2_743 ( .A(core_v2_reg_9_), .B(core_v3_reg_9_), .Y(core__abc_22172_new_n1431_));
OR2X2 OR2X2_744 ( .A(core__abc_22172_new_n1428_), .B(core__abc_22172_new_n1432_), .Y(core__abc_22172_new_n1433_));
OR2X2 OR2X2_745 ( .A(core__abc_22172_new_n1434_), .B(core__abc_22172_new_n1435_), .Y(core__abc_22172_new_n1436_));
OR2X2 OR2X2_746 ( .A(core__abc_22172_new_n1437_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n1438_));
OR2X2 OR2X2_747 ( .A(core_siphash_word1_we), .B(core_siphash_word_73_), .Y(core__abc_22172_new_n1439_));
OR2X2 OR2X2_748 ( .A(core_v1_reg_10_), .B(core_v0_reg_10_), .Y(core__abc_22172_new_n1442_));
OR2X2 OR2X2_749 ( .A(core_v2_reg_10_), .B(core_v3_reg_10_), .Y(core__abc_22172_new_n1448_));
OR2X2 OR2X2_75 ( .A(_abc_19873_new_n1073_), .B(_abc_19873_new_n1074_), .Y(_abc_19873_new_n1075_));
OR2X2 OR2X2_750 ( .A(core__abc_22172_new_n1445_), .B(core__abc_22172_new_n1449_), .Y(core__abc_22172_new_n1450_));
OR2X2 OR2X2_751 ( .A(core__abc_22172_new_n1452_), .B(core__abc_22172_new_n1451_), .Y(core__abc_22172_new_n1453_));
OR2X2 OR2X2_752 ( .A(core__abc_22172_new_n1454_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n1455_));
OR2X2 OR2X2_753 ( .A(core_siphash_word1_we), .B(core_siphash_word_74_), .Y(core__abc_22172_new_n1456_));
OR2X2 OR2X2_754 ( .A(core_v1_reg_11_), .B(core_v0_reg_11_), .Y(core__abc_22172_new_n1459_));
OR2X2 OR2X2_755 ( .A(core_v2_reg_11_), .B(core_v3_reg_11_), .Y(core__abc_22172_new_n1465_));
OR2X2 OR2X2_756 ( .A(core__abc_22172_new_n1462_), .B(core__abc_22172_new_n1466_), .Y(core__abc_22172_new_n1467_));
OR2X2 OR2X2_757 ( .A(core__abc_22172_new_n1469_), .B(core__abc_22172_new_n1468_), .Y(core__abc_22172_new_n1470_));
OR2X2 OR2X2_758 ( .A(core__abc_22172_new_n1471_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n1472_));
OR2X2 OR2X2_759 ( .A(core_siphash_word1_we), .B(core_siphash_word_75_), .Y(core__abc_22172_new_n1473_));
OR2X2 OR2X2_76 ( .A(_abc_19873_new_n1072_), .B(_abc_19873_new_n1075_), .Y(_abc_19873_new_n1076_));
OR2X2 OR2X2_760 ( .A(core_v1_reg_12_), .B(core_v0_reg_12_), .Y(core__abc_22172_new_n1476_));
OR2X2 OR2X2_761 ( .A(core_v2_reg_12_), .B(core_v3_reg_12_), .Y(core__abc_22172_new_n1482_));
OR2X2 OR2X2_762 ( .A(core__abc_22172_new_n1479_), .B(core__abc_22172_new_n1483_), .Y(core__abc_22172_new_n1484_));
OR2X2 OR2X2_763 ( .A(core__abc_22172_new_n1485_), .B(core__abc_22172_new_n1486_), .Y(core__abc_22172_new_n1487_));
OR2X2 OR2X2_764 ( .A(core__abc_22172_new_n1488_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n1489_));
OR2X2 OR2X2_765 ( .A(core_siphash_word1_we), .B(core_siphash_word_76_), .Y(core__abc_22172_new_n1490_));
OR2X2 OR2X2_766 ( .A(core_v1_reg_13_), .B(core_v0_reg_13_), .Y(core__abc_22172_new_n1493_));
OR2X2 OR2X2_767 ( .A(core_v2_reg_13_), .B(core_v3_reg_13_), .Y(core__abc_22172_new_n1499_));
OR2X2 OR2X2_768 ( .A(core__abc_22172_new_n1496_), .B(core__abc_22172_new_n1500_), .Y(core__abc_22172_new_n1501_));
OR2X2 OR2X2_769 ( .A(core__abc_22172_new_n1502_), .B(core__abc_22172_new_n1503_), .Y(core__abc_22172_new_n1504_));
OR2X2 OR2X2_77 ( .A(_abc_19873_new_n1077_), .B(_abc_19873_new_n994_), .Y(_abc_19873_new_n1078_));
OR2X2 OR2X2_770 ( .A(core__abc_22172_new_n1505_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n1506_));
OR2X2 OR2X2_771 ( .A(core_siphash_word1_we), .B(core_siphash_word_77_), .Y(core__abc_22172_new_n1507_));
OR2X2 OR2X2_772 ( .A(core_v1_reg_14_), .B(core_v0_reg_14_), .Y(core__abc_22172_new_n1510_));
OR2X2 OR2X2_773 ( .A(core_v2_reg_14_), .B(core_v3_reg_14_), .Y(core__abc_22172_new_n1516_));
OR2X2 OR2X2_774 ( .A(core__abc_22172_new_n1513_), .B(core__abc_22172_new_n1517_), .Y(core__abc_22172_new_n1518_));
OR2X2 OR2X2_775 ( .A(core__abc_22172_new_n1519_), .B(core__abc_22172_new_n1520_), .Y(core__abc_22172_new_n1521_));
OR2X2 OR2X2_776 ( .A(core__abc_22172_new_n1522_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n1523_));
OR2X2 OR2X2_777 ( .A(core_siphash_word1_we), .B(core_siphash_word_78_), .Y(core__abc_22172_new_n1524_));
OR2X2 OR2X2_778 ( .A(core_v1_reg_15_), .B(core_v0_reg_15_), .Y(core__abc_22172_new_n1527_));
OR2X2 OR2X2_779 ( .A(core_v2_reg_15_), .B(core_v3_reg_15_), .Y(core__abc_22172_new_n1533_));
OR2X2 OR2X2_78 ( .A(_abc_19873_new_n1079_), .B(_abc_19873_new_n1080_), .Y(_abc_19873_new_n1081_));
OR2X2 OR2X2_780 ( .A(core__abc_22172_new_n1530_), .B(core__abc_22172_new_n1534_), .Y(core__abc_22172_new_n1535_));
OR2X2 OR2X2_781 ( .A(core__abc_22172_new_n1536_), .B(core__abc_22172_new_n1537_), .Y(core__abc_22172_new_n1538_));
OR2X2 OR2X2_782 ( .A(core__abc_22172_new_n1539_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n1540_));
OR2X2 OR2X2_783 ( .A(core_siphash_word1_we), .B(core_siphash_word_79_), .Y(core__abc_22172_new_n1541_));
OR2X2 OR2X2_784 ( .A(core_v1_reg_16_), .B(core_v0_reg_16_), .Y(core__abc_22172_new_n1544_));
OR2X2 OR2X2_785 ( .A(core_v2_reg_16_), .B(core_v3_reg_16_), .Y(core__abc_22172_new_n1550_));
OR2X2 OR2X2_786 ( .A(core__abc_22172_new_n1547_), .B(core__abc_22172_new_n1551_), .Y(core__abc_22172_new_n1552_));
OR2X2 OR2X2_787 ( .A(core__abc_22172_new_n1553_), .B(core__abc_22172_new_n1554_), .Y(core__abc_22172_new_n1555_));
OR2X2 OR2X2_788 ( .A(core__abc_22172_new_n1556_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n1557_));
OR2X2 OR2X2_789 ( .A(core_siphash_word1_we), .B(core_siphash_word_80_), .Y(core__abc_22172_new_n1558_));
OR2X2 OR2X2_79 ( .A(_abc_19873_new_n1081_), .B(_abc_19873_new_n1078_), .Y(_abc_19873_new_n1082_));
OR2X2 OR2X2_790 ( .A(core_v1_reg_17_), .B(core_v0_reg_17_), .Y(core__abc_22172_new_n1561_));
OR2X2 OR2X2_791 ( .A(core_v2_reg_17_), .B(core_v3_reg_17_), .Y(core__abc_22172_new_n1567_));
OR2X2 OR2X2_792 ( .A(core__abc_22172_new_n1564_), .B(core__abc_22172_new_n1568_), .Y(core__abc_22172_new_n1569_));
OR2X2 OR2X2_793 ( .A(core__abc_22172_new_n1570_), .B(core__abc_22172_new_n1571_), .Y(core__abc_22172_new_n1572_));
OR2X2 OR2X2_794 ( .A(core__abc_22172_new_n1573_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n1574_));
OR2X2 OR2X2_795 ( .A(core_siphash_word1_we), .B(core_siphash_word_81_), .Y(core__abc_22172_new_n1575_));
OR2X2 OR2X2_796 ( .A(core_v1_reg_18_), .B(core_v0_reg_18_), .Y(core__abc_22172_new_n1578_));
OR2X2 OR2X2_797 ( .A(core_v2_reg_18_), .B(core_v3_reg_18_), .Y(core__abc_22172_new_n1584_));
OR2X2 OR2X2_798 ( .A(core__abc_22172_new_n1581_), .B(core__abc_22172_new_n1585_), .Y(core__abc_22172_new_n1586_));
OR2X2 OR2X2_799 ( .A(core__abc_22172_new_n1588_), .B(core__abc_22172_new_n1587_), .Y(core__abc_22172_new_n1589_));
OR2X2 OR2X2_8 ( .A(_abc_19873_new_n924_), .B(_abc_19873_new_n926_), .Y(_abc_19873_new_n927_));
OR2X2 OR2X2_80 ( .A(_abc_19873_new_n1076_), .B(_abc_19873_new_n1082_), .Y(_abc_19873_new_n1083_));
OR2X2 OR2X2_800 ( .A(core__abc_22172_new_n1590_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n1591_));
OR2X2 OR2X2_801 ( .A(core_siphash_word1_we), .B(core_siphash_word_82_), .Y(core__abc_22172_new_n1592_));
OR2X2 OR2X2_802 ( .A(core_v1_reg_19_), .B(core_v0_reg_19_), .Y(core__abc_22172_new_n1595_));
OR2X2 OR2X2_803 ( .A(core_v2_reg_19_), .B(core_v3_reg_19_), .Y(core__abc_22172_new_n1601_));
OR2X2 OR2X2_804 ( .A(core__abc_22172_new_n1598_), .B(core__abc_22172_new_n1602_), .Y(core__abc_22172_new_n1603_));
OR2X2 OR2X2_805 ( .A(core__abc_22172_new_n1605_), .B(core__abc_22172_new_n1604_), .Y(core__abc_22172_new_n1606_));
OR2X2 OR2X2_806 ( .A(core__abc_22172_new_n1607_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n1608_));
OR2X2 OR2X2_807 ( .A(core_siphash_word1_we), .B(core_siphash_word_83_), .Y(core__abc_22172_new_n1609_));
OR2X2 OR2X2_808 ( .A(core_v1_reg_20_), .B(core_v0_reg_20_), .Y(core__abc_22172_new_n1612_));
OR2X2 OR2X2_809 ( .A(core_v2_reg_20_), .B(core_v3_reg_20_), .Y(core__abc_22172_new_n1618_));
OR2X2 OR2X2_81 ( .A(_abc_19873_new_n1083_), .B(_abc_19873_new_n1069_), .Y(_abc_19873_new_n1084_));
OR2X2 OR2X2_810 ( .A(core__abc_22172_new_n1615_), .B(core__abc_22172_new_n1619_), .Y(core__abc_22172_new_n1620_));
OR2X2 OR2X2_811 ( .A(core__abc_22172_new_n1621_), .B(core__abc_22172_new_n1622_), .Y(core__abc_22172_new_n1623_));
OR2X2 OR2X2_812 ( .A(core__abc_22172_new_n1624_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n1625_));
OR2X2 OR2X2_813 ( .A(core_siphash_word1_we), .B(core_siphash_word_84_), .Y(core__abc_22172_new_n1626_));
OR2X2 OR2X2_814 ( .A(core_v1_reg_21_), .B(core_v0_reg_21_), .Y(core__abc_22172_new_n1629_));
OR2X2 OR2X2_815 ( .A(core_v2_reg_21_), .B(core_v3_reg_21_), .Y(core__abc_22172_new_n1635_));
OR2X2 OR2X2_816 ( .A(core__abc_22172_new_n1632_), .B(core__abc_22172_new_n1636_), .Y(core__abc_22172_new_n1637_));
OR2X2 OR2X2_817 ( .A(core__abc_22172_new_n1638_), .B(core__abc_22172_new_n1639_), .Y(core__abc_22172_new_n1640_));
OR2X2 OR2X2_818 ( .A(core__abc_22172_new_n1641_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n1642_));
OR2X2 OR2X2_819 ( .A(core_siphash_word1_we), .B(core_siphash_word_85_), .Y(core__abc_22172_new_n1643_));
OR2X2 OR2X2_82 ( .A(_abc_19873_new_n1086_), .B(_abc_19873_new_n1087_), .Y(_abc_19873_new_n1088_));
OR2X2 OR2X2_820 ( .A(core_v1_reg_22_), .B(core_v0_reg_22_), .Y(core__abc_22172_new_n1646_));
OR2X2 OR2X2_821 ( .A(core_v2_reg_22_), .B(core_v3_reg_22_), .Y(core__abc_22172_new_n1652_));
OR2X2 OR2X2_822 ( .A(core__abc_22172_new_n1649_), .B(core__abc_22172_new_n1653_), .Y(core__abc_22172_new_n1654_));
OR2X2 OR2X2_823 ( .A(core__abc_22172_new_n1655_), .B(core__abc_22172_new_n1656_), .Y(core__abc_22172_new_n1657_));
OR2X2 OR2X2_824 ( .A(core__abc_22172_new_n1658_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n1659_));
OR2X2 OR2X2_825 ( .A(core_siphash_word1_we), .B(core_siphash_word_86_), .Y(core__abc_22172_new_n1660_));
OR2X2 OR2X2_826 ( .A(core_v1_reg_23_), .B(core_v0_reg_23_), .Y(core__abc_22172_new_n1663_));
OR2X2 OR2X2_827 ( .A(core_v2_reg_23_), .B(core_v3_reg_23_), .Y(core__abc_22172_new_n1669_));
OR2X2 OR2X2_828 ( .A(core__abc_22172_new_n1666_), .B(core__abc_22172_new_n1670_), .Y(core__abc_22172_new_n1671_));
OR2X2 OR2X2_829 ( .A(core__abc_22172_new_n1672_), .B(core__abc_22172_new_n1673_), .Y(core__abc_22172_new_n1674_));
OR2X2 OR2X2_83 ( .A(_abc_19873_new_n1089_), .B(_abc_19873_new_n1090_), .Y(_abc_19873_new_n1091_));
OR2X2 OR2X2_830 ( .A(core__abc_22172_new_n1675_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n1676_));
OR2X2 OR2X2_831 ( .A(core_siphash_word1_we), .B(core_siphash_word_87_), .Y(core__abc_22172_new_n1677_));
OR2X2 OR2X2_832 ( .A(core_v1_reg_24_), .B(core_v0_reg_24_), .Y(core__abc_22172_new_n1680_));
OR2X2 OR2X2_833 ( .A(core_v2_reg_24_), .B(core_v3_reg_24_), .Y(core__abc_22172_new_n1686_));
OR2X2 OR2X2_834 ( .A(core__abc_22172_new_n1683_), .B(core__abc_22172_new_n1687_), .Y(core__abc_22172_new_n1688_));
OR2X2 OR2X2_835 ( .A(core__abc_22172_new_n1689_), .B(core__abc_22172_new_n1690_), .Y(core__abc_22172_new_n1691_));
OR2X2 OR2X2_836 ( .A(core__abc_22172_new_n1692_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n1693_));
OR2X2 OR2X2_837 ( .A(core_siphash_word1_we), .B(core_siphash_word_88_), .Y(core__abc_22172_new_n1694_));
OR2X2 OR2X2_838 ( .A(core_v1_reg_25_), .B(core_v0_reg_25_), .Y(core__abc_22172_new_n1697_));
OR2X2 OR2X2_839 ( .A(core_v2_reg_25_), .B(core_v3_reg_25_), .Y(core__abc_22172_new_n1703_));
OR2X2 OR2X2_84 ( .A(_abc_19873_new_n1088_), .B(_abc_19873_new_n1091_), .Y(_abc_19873_new_n1092_));
OR2X2 OR2X2_840 ( .A(core__abc_22172_new_n1700_), .B(core__abc_22172_new_n1704_), .Y(core__abc_22172_new_n1705_));
OR2X2 OR2X2_841 ( .A(core__abc_22172_new_n1706_), .B(core__abc_22172_new_n1707_), .Y(core__abc_22172_new_n1708_));
OR2X2 OR2X2_842 ( .A(core__abc_22172_new_n1709_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n1710_));
OR2X2 OR2X2_843 ( .A(core_siphash_word1_we), .B(core_siphash_word_89_), .Y(core__abc_22172_new_n1711_));
OR2X2 OR2X2_844 ( .A(core_v1_reg_26_), .B(core_v0_reg_26_), .Y(core__abc_22172_new_n1714_));
OR2X2 OR2X2_845 ( .A(core_v2_reg_26_), .B(core_v3_reg_26_), .Y(core__abc_22172_new_n1720_));
OR2X2 OR2X2_846 ( .A(core__abc_22172_new_n1717_), .B(core__abc_22172_new_n1721_), .Y(core__abc_22172_new_n1722_));
OR2X2 OR2X2_847 ( .A(core__abc_22172_new_n1723_), .B(core__abc_22172_new_n1724_), .Y(core__abc_22172_new_n1725_));
OR2X2 OR2X2_848 ( .A(core__abc_22172_new_n1726_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n1727_));
OR2X2 OR2X2_849 ( .A(core_siphash_word1_we), .B(core_siphash_word_90_), .Y(core__abc_22172_new_n1728_));
OR2X2 OR2X2_85 ( .A(_abc_19873_new_n1094_), .B(_abc_19873_new_n1095_), .Y(_abc_19873_new_n1096_));
OR2X2 OR2X2_850 ( .A(core_v1_reg_27_), .B(core_v0_reg_27_), .Y(core__abc_22172_new_n1731_));
OR2X2 OR2X2_851 ( .A(core_v2_reg_27_), .B(core_v3_reg_27_), .Y(core__abc_22172_new_n1737_));
OR2X2 OR2X2_852 ( .A(core__abc_22172_new_n1734_), .B(core__abc_22172_new_n1738_), .Y(core__abc_22172_new_n1739_));
OR2X2 OR2X2_853 ( .A(core__abc_22172_new_n1740_), .B(core__abc_22172_new_n1741_), .Y(core__abc_22172_new_n1742_));
OR2X2 OR2X2_854 ( .A(core__abc_22172_new_n1743_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n1744_));
OR2X2 OR2X2_855 ( .A(core_siphash_word1_we), .B(core_siphash_word_91_), .Y(core__abc_22172_new_n1745_));
OR2X2 OR2X2_856 ( .A(core_v1_reg_28_), .B(core_v0_reg_28_), .Y(core__abc_22172_new_n1748_));
OR2X2 OR2X2_857 ( .A(core_v2_reg_28_), .B(core_v3_reg_28_), .Y(core__abc_22172_new_n1754_));
OR2X2 OR2X2_858 ( .A(core__abc_22172_new_n1751_), .B(core__abc_22172_new_n1755_), .Y(core__abc_22172_new_n1756_));
OR2X2 OR2X2_859 ( .A(core__abc_22172_new_n1757_), .B(core__abc_22172_new_n1758_), .Y(core__abc_22172_new_n1759_));
OR2X2 OR2X2_86 ( .A(_abc_19873_new_n1096_), .B(_abc_19873_new_n1093_), .Y(_abc_19873_new_n1097_));
OR2X2 OR2X2_860 ( .A(core__abc_22172_new_n1760_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n1761_));
OR2X2 OR2X2_861 ( .A(core_siphash_word1_we), .B(core_siphash_word_92_), .Y(core__abc_22172_new_n1762_));
OR2X2 OR2X2_862 ( .A(core_v1_reg_29_), .B(core_v0_reg_29_), .Y(core__abc_22172_new_n1765_));
OR2X2 OR2X2_863 ( .A(core_v2_reg_29_), .B(core_v3_reg_29_), .Y(core__abc_22172_new_n1771_));
OR2X2 OR2X2_864 ( .A(core__abc_22172_new_n1768_), .B(core__abc_22172_new_n1772_), .Y(core__abc_22172_new_n1773_));
OR2X2 OR2X2_865 ( .A(core__abc_22172_new_n1774_), .B(core__abc_22172_new_n1775_), .Y(core__abc_22172_new_n1776_));
OR2X2 OR2X2_866 ( .A(core__abc_22172_new_n1777_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n1778_));
OR2X2 OR2X2_867 ( .A(core_siphash_word1_we), .B(core_siphash_word_93_), .Y(core__abc_22172_new_n1779_));
OR2X2 OR2X2_868 ( .A(core_v1_reg_30_), .B(core_v0_reg_30_), .Y(core__abc_22172_new_n1782_));
OR2X2 OR2X2_869 ( .A(core_v2_reg_30_), .B(core_v3_reg_30_), .Y(core__abc_22172_new_n1788_));
OR2X2 OR2X2_87 ( .A(_abc_19873_new_n1098_), .B(_abc_19873_new_n1099_), .Y(_abc_19873_new_n1100_));
OR2X2 OR2X2_870 ( .A(core__abc_22172_new_n1785_), .B(core__abc_22172_new_n1789_), .Y(core__abc_22172_new_n1790_));
OR2X2 OR2X2_871 ( .A(core__abc_22172_new_n1791_), .B(core__abc_22172_new_n1792_), .Y(core__abc_22172_new_n1793_));
OR2X2 OR2X2_872 ( .A(core__abc_22172_new_n1794_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n1795_));
OR2X2 OR2X2_873 ( .A(core_siphash_word1_we), .B(core_siphash_word_94_), .Y(core__abc_22172_new_n1796_));
OR2X2 OR2X2_874 ( .A(core_v1_reg_31_), .B(core_v0_reg_31_), .Y(core__abc_22172_new_n1799_));
OR2X2 OR2X2_875 ( .A(core_v2_reg_31_), .B(core_v3_reg_31_), .Y(core__abc_22172_new_n1805_));
OR2X2 OR2X2_876 ( .A(core__abc_22172_new_n1802_), .B(core__abc_22172_new_n1806_), .Y(core__abc_22172_new_n1807_));
OR2X2 OR2X2_877 ( .A(core__abc_22172_new_n1808_), .B(core__abc_22172_new_n1809_), .Y(core__abc_22172_new_n1810_));
OR2X2 OR2X2_878 ( .A(core__abc_22172_new_n1811_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n1812_));
OR2X2 OR2X2_879 ( .A(core_siphash_word1_we), .B(core_siphash_word_95_), .Y(core__abc_22172_new_n1813_));
OR2X2 OR2X2_88 ( .A(_abc_19873_new_n1101_), .B(_abc_19873_new_n1102_), .Y(_abc_19873_new_n1103_));
OR2X2 OR2X2_880 ( .A(core_v1_reg_32_), .B(core_v0_reg_32_), .Y(core__abc_22172_new_n1816_));
OR2X2 OR2X2_881 ( .A(core_v2_reg_32_), .B(core_v3_reg_32_), .Y(core__abc_22172_new_n1822_));
OR2X2 OR2X2_882 ( .A(core__abc_22172_new_n1819_), .B(core__abc_22172_new_n1823_), .Y(core__abc_22172_new_n1824_));
OR2X2 OR2X2_883 ( .A(core__abc_22172_new_n1825_), .B(core__abc_22172_new_n1826_), .Y(core__abc_22172_new_n1827_));
OR2X2 OR2X2_884 ( .A(core__abc_22172_new_n1828_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n1829_));
OR2X2 OR2X2_885 ( .A(core_siphash_word1_we), .B(core_siphash_word_96_), .Y(core__abc_22172_new_n1830_));
OR2X2 OR2X2_886 ( .A(core_v1_reg_33_), .B(core_v0_reg_33_), .Y(core__abc_22172_new_n1833_));
OR2X2 OR2X2_887 ( .A(core_v2_reg_33_), .B(core_v3_reg_33_), .Y(core__abc_22172_new_n1839_));
OR2X2 OR2X2_888 ( .A(core__abc_22172_new_n1836_), .B(core__abc_22172_new_n1840_), .Y(core__abc_22172_new_n1841_));
OR2X2 OR2X2_889 ( .A(core__abc_22172_new_n1842_), .B(core__abc_22172_new_n1843_), .Y(core__abc_22172_new_n1844_));
OR2X2 OR2X2_89 ( .A(_abc_19873_new_n1100_), .B(_abc_19873_new_n1103_), .Y(_abc_19873_new_n1104_));
OR2X2 OR2X2_890 ( .A(core__abc_22172_new_n1845_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n1846_));
OR2X2 OR2X2_891 ( .A(core_siphash_word1_we), .B(core_siphash_word_97_), .Y(core__abc_22172_new_n1847_));
OR2X2 OR2X2_892 ( .A(core_v1_reg_34_), .B(core_v0_reg_34_), .Y(core__abc_22172_new_n1850_));
OR2X2 OR2X2_893 ( .A(core_v2_reg_34_), .B(core_v3_reg_34_), .Y(core__abc_22172_new_n1854_));
OR2X2 OR2X2_894 ( .A(core__abc_22172_new_n1853_), .B(core__abc_22172_new_n1857_), .Y(core__abc_22172_new_n1858_));
OR2X2 OR2X2_895 ( .A(core__abc_22172_new_n1859_), .B(core__abc_22172_new_n1860_), .Y(core__abc_22172_new_n1861_));
OR2X2 OR2X2_896 ( .A(core__abc_22172_new_n1862_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n1863_));
OR2X2 OR2X2_897 ( .A(core_siphash_word1_we), .B(core_siphash_word_98_), .Y(core__abc_22172_new_n1864_));
OR2X2 OR2X2_898 ( .A(core_v1_reg_35_), .B(core_v0_reg_35_), .Y(core__abc_22172_new_n1867_));
OR2X2 OR2X2_899 ( .A(core_v2_reg_35_), .B(core_v3_reg_35_), .Y(core__abc_22172_new_n1873_));
OR2X2 OR2X2_9 ( .A(_abc_19873_new_n929_), .B(_abc_19873_new_n931_), .Y(_abc_19873_new_n932_));
OR2X2 OR2X2_90 ( .A(_abc_19873_new_n1104_), .B(_abc_19873_new_n1097_), .Y(_abc_19873_new_n1105_));
OR2X2 OR2X2_900 ( .A(core__abc_22172_new_n1870_), .B(core__abc_22172_new_n1874_), .Y(core__abc_22172_new_n1875_));
OR2X2 OR2X2_901 ( .A(core__abc_22172_new_n1876_), .B(core__abc_22172_new_n1877_), .Y(core__abc_22172_new_n1878_));
OR2X2 OR2X2_902 ( .A(core__abc_22172_new_n1879_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n1880_));
OR2X2 OR2X2_903 ( .A(core_siphash_word1_we), .B(core_siphash_word_99_), .Y(core__abc_22172_new_n1881_));
OR2X2 OR2X2_904 ( .A(core_v1_reg_36_), .B(core_v0_reg_36_), .Y(core__abc_22172_new_n1884_));
OR2X2 OR2X2_905 ( .A(core_v2_reg_36_), .B(core_v3_reg_36_), .Y(core__abc_22172_new_n1888_));
OR2X2 OR2X2_906 ( .A(core__abc_22172_new_n1887_), .B(core__abc_22172_new_n1891_), .Y(core__abc_22172_new_n1892_));
OR2X2 OR2X2_907 ( .A(core__abc_22172_new_n1893_), .B(core__abc_22172_new_n1894_), .Y(core__abc_22172_new_n1895_));
OR2X2 OR2X2_908 ( .A(core__abc_22172_new_n1896_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n1897_));
OR2X2 OR2X2_909 ( .A(core_siphash_word1_we), .B(core_siphash_word_100_), .Y(core__abc_22172_new_n1898_));
OR2X2 OR2X2_91 ( .A(_abc_19873_new_n1105_), .B(_abc_19873_new_n1092_), .Y(_abc_19873_new_n1106_));
OR2X2 OR2X2_910 ( .A(core_v1_reg_37_), .B(core_v0_reg_37_), .Y(core__abc_22172_new_n1901_));
OR2X2 OR2X2_911 ( .A(core_v2_reg_37_), .B(core_v3_reg_37_), .Y(core__abc_22172_new_n1907_));
OR2X2 OR2X2_912 ( .A(core__abc_22172_new_n1904_), .B(core__abc_22172_new_n1908_), .Y(core__abc_22172_new_n1909_));
OR2X2 OR2X2_913 ( .A(core__abc_22172_new_n1910_), .B(core__abc_22172_new_n1911_), .Y(core__abc_22172_new_n1912_));
OR2X2 OR2X2_914 ( .A(core__abc_22172_new_n1913_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n1914_));
OR2X2 OR2X2_915 ( .A(core_siphash_word1_we), .B(core_siphash_word_101_), .Y(core__abc_22172_new_n1915_));
OR2X2 OR2X2_916 ( .A(core_v1_reg_38_), .B(core_v0_reg_38_), .Y(core__abc_22172_new_n1918_));
OR2X2 OR2X2_917 ( .A(core_v2_reg_38_), .B(core_v3_reg_38_), .Y(core__abc_22172_new_n1922_));
OR2X2 OR2X2_918 ( .A(core__abc_22172_new_n1921_), .B(core__abc_22172_new_n1925_), .Y(core__abc_22172_new_n1926_));
OR2X2 OR2X2_919 ( .A(core__abc_22172_new_n1927_), .B(core__abc_22172_new_n1928_), .Y(core__abc_22172_new_n1929_));
OR2X2 OR2X2_92 ( .A(_abc_19873_new_n1108_), .B(_abc_19873_new_n1109_), .Y(_abc_19873_new_n1110_));
OR2X2 OR2X2_920 ( .A(core__abc_22172_new_n1930_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n1931_));
OR2X2 OR2X2_921 ( .A(core_siphash_word1_we), .B(core_siphash_word_102_), .Y(core__abc_22172_new_n1932_));
OR2X2 OR2X2_922 ( .A(core_v1_reg_39_), .B(core_v0_reg_39_), .Y(core__abc_22172_new_n1935_));
OR2X2 OR2X2_923 ( .A(core_v2_reg_39_), .B(core_v3_reg_39_), .Y(core__abc_22172_new_n1941_));
OR2X2 OR2X2_924 ( .A(core__abc_22172_new_n1938_), .B(core__abc_22172_new_n1942_), .Y(core__abc_22172_new_n1943_));
OR2X2 OR2X2_925 ( .A(core__abc_22172_new_n1944_), .B(core__abc_22172_new_n1945_), .Y(core__abc_22172_new_n1946_));
OR2X2 OR2X2_926 ( .A(core__abc_22172_new_n1947_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n1948_));
OR2X2 OR2X2_927 ( .A(core_siphash_word1_we), .B(core_siphash_word_103_), .Y(core__abc_22172_new_n1949_));
OR2X2 OR2X2_928 ( .A(core_v1_reg_40_), .B(core_v0_reg_40_), .Y(core__abc_22172_new_n1952_));
OR2X2 OR2X2_929 ( .A(core_v2_reg_40_), .B(core_v3_reg_40_), .Y(core__abc_22172_new_n1958_));
OR2X2 OR2X2_93 ( .A(_abc_19873_new_n1112_), .B(_abc_19873_new_n1113_), .Y(_abc_19873_new_n1114_));
OR2X2 OR2X2_930 ( .A(core__abc_22172_new_n1955_), .B(core__abc_22172_new_n1959_), .Y(core__abc_22172_new_n1960_));
OR2X2 OR2X2_931 ( .A(core__abc_22172_new_n1961_), .B(core__abc_22172_new_n1962_), .Y(core__abc_22172_new_n1963_));
OR2X2 OR2X2_932 ( .A(core__abc_22172_new_n1964_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n1965_));
OR2X2 OR2X2_933 ( .A(core_siphash_word1_we), .B(core_siphash_word_104_), .Y(core__abc_22172_new_n1966_));
OR2X2 OR2X2_934 ( .A(core_v1_reg_41_), .B(core_v0_reg_41_), .Y(core__abc_22172_new_n1969_));
OR2X2 OR2X2_935 ( .A(core_v2_reg_41_), .B(core_v3_reg_41_), .Y(core__abc_22172_new_n1975_));
OR2X2 OR2X2_936 ( .A(core__abc_22172_new_n1972_), .B(core__abc_22172_new_n1976_), .Y(core__abc_22172_new_n1977_));
OR2X2 OR2X2_937 ( .A(core__abc_22172_new_n1978_), .B(core__abc_22172_new_n1979_), .Y(core__abc_22172_new_n1980_));
OR2X2 OR2X2_938 ( .A(core__abc_22172_new_n1981_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n1982_));
OR2X2 OR2X2_939 ( .A(core_siphash_word1_we), .B(core_siphash_word_105_), .Y(core__abc_22172_new_n1983_));
OR2X2 OR2X2_94 ( .A(_abc_19873_new_n1114_), .B(_abc_19873_new_n1111_), .Y(_abc_19873_new_n1115_));
OR2X2 OR2X2_940 ( .A(core_v1_reg_42_), .B(core_v0_reg_42_), .Y(core__abc_22172_new_n1986_));
OR2X2 OR2X2_941 ( .A(core_v2_reg_42_), .B(core_v3_reg_42_), .Y(core__abc_22172_new_n1992_));
OR2X2 OR2X2_942 ( .A(core__abc_22172_new_n1989_), .B(core__abc_22172_new_n1993_), .Y(core__abc_22172_new_n1994_));
OR2X2 OR2X2_943 ( .A(core__abc_22172_new_n1995_), .B(core__abc_22172_new_n1996_), .Y(core__abc_22172_new_n1997_));
OR2X2 OR2X2_944 ( .A(core__abc_22172_new_n1998_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n1999_));
OR2X2 OR2X2_945 ( .A(core_siphash_word1_we), .B(core_siphash_word_106_), .Y(core__abc_22172_new_n2000_));
OR2X2 OR2X2_946 ( .A(core_v1_reg_43_), .B(core_v0_reg_43_), .Y(core__abc_22172_new_n2003_));
OR2X2 OR2X2_947 ( .A(core_v2_reg_43_), .B(core_v3_reg_43_), .Y(core__abc_22172_new_n2007_));
OR2X2 OR2X2_948 ( .A(core__abc_22172_new_n2006_), .B(core__abc_22172_new_n2010_), .Y(core__abc_22172_new_n2011_));
OR2X2 OR2X2_949 ( .A(core__abc_22172_new_n2012_), .B(core__abc_22172_new_n2013_), .Y(core__abc_22172_new_n2014_));
OR2X2 OR2X2_95 ( .A(_abc_19873_new_n1115_), .B(_abc_19873_new_n1110_), .Y(_abc_19873_new_n1116_));
OR2X2 OR2X2_950 ( .A(core__abc_22172_new_n2015_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n2016_));
OR2X2 OR2X2_951 ( .A(core_siphash_word1_we), .B(core_siphash_word_107_), .Y(core__abc_22172_new_n2017_));
OR2X2 OR2X2_952 ( .A(core_v1_reg_44_), .B(core_v0_reg_44_), .Y(core__abc_22172_new_n2020_));
OR2X2 OR2X2_953 ( .A(core_v2_reg_44_), .B(core_v3_reg_44_), .Y(core__abc_22172_new_n2024_));
OR2X2 OR2X2_954 ( .A(core__abc_22172_new_n2023_), .B(core__abc_22172_new_n2027_), .Y(core__abc_22172_new_n2028_));
OR2X2 OR2X2_955 ( .A(core__abc_22172_new_n2029_), .B(core__abc_22172_new_n2030_), .Y(core__abc_22172_new_n2031_));
OR2X2 OR2X2_956 ( .A(core__abc_22172_new_n2032_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n2033_));
OR2X2 OR2X2_957 ( .A(core_siphash_word1_we), .B(core_siphash_word_108_), .Y(core__abc_22172_new_n2034_));
OR2X2 OR2X2_958 ( .A(core_v1_reg_45_), .B(core_v0_reg_45_), .Y(core__abc_22172_new_n2037_));
OR2X2 OR2X2_959 ( .A(core_v2_reg_45_), .B(core_v3_reg_45_), .Y(core__abc_22172_new_n2041_));
OR2X2 OR2X2_96 ( .A(_abc_19873_new_n1118_), .B(_abc_19873_new_n1119_), .Y(_abc_19873_new_n1120_));
OR2X2 OR2X2_960 ( .A(core__abc_22172_new_n2040_), .B(core__abc_22172_new_n2044_), .Y(core__abc_22172_new_n2045_));
OR2X2 OR2X2_961 ( .A(core__abc_22172_new_n2046_), .B(core__abc_22172_new_n2047_), .Y(core__abc_22172_new_n2048_));
OR2X2 OR2X2_962 ( .A(core__abc_22172_new_n2049_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n2050_));
OR2X2 OR2X2_963 ( .A(core_siphash_word1_we), .B(core_siphash_word_109_), .Y(core__abc_22172_new_n2051_));
OR2X2 OR2X2_964 ( .A(core_v1_reg_46_), .B(core_v0_reg_46_), .Y(core__abc_22172_new_n2054_));
OR2X2 OR2X2_965 ( .A(core_v2_reg_46_), .B(core_v3_reg_46_), .Y(core__abc_22172_new_n2058_));
OR2X2 OR2X2_966 ( .A(core__abc_22172_new_n2057_), .B(core__abc_22172_new_n2061_), .Y(core__abc_22172_new_n2062_));
OR2X2 OR2X2_967 ( .A(core__abc_22172_new_n2063_), .B(core__abc_22172_new_n2064_), .Y(core__abc_22172_new_n2065_));
OR2X2 OR2X2_968 ( .A(core__abc_22172_new_n2066_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n2067_));
OR2X2 OR2X2_969 ( .A(core_siphash_word1_we), .B(core_siphash_word_110_), .Y(core__abc_22172_new_n2068_));
OR2X2 OR2X2_97 ( .A(_abc_19873_new_n1121_), .B(_abc_19873_new_n1122_), .Y(_abc_19873_new_n1123_));
OR2X2 OR2X2_970 ( .A(core_v1_reg_47_), .B(core_v0_reg_47_), .Y(core__abc_22172_new_n2071_));
OR2X2 OR2X2_971 ( .A(core_v2_reg_47_), .B(core_v3_reg_47_), .Y(core__abc_22172_new_n2075_));
OR2X2 OR2X2_972 ( .A(core__abc_22172_new_n2074_), .B(core__abc_22172_new_n2078_), .Y(core__abc_22172_new_n2079_));
OR2X2 OR2X2_973 ( .A(core__abc_22172_new_n2080_), .B(core__abc_22172_new_n2081_), .Y(core__abc_22172_new_n2082_));
OR2X2 OR2X2_974 ( .A(core__abc_22172_new_n2083_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n2084_));
OR2X2 OR2X2_975 ( .A(core_siphash_word1_we), .B(core_siphash_word_111_), .Y(core__abc_22172_new_n2085_));
OR2X2 OR2X2_976 ( .A(core_v1_reg_48_), .B(core_v0_reg_48_), .Y(core__abc_22172_new_n2088_));
OR2X2 OR2X2_977 ( .A(core_v2_reg_48_), .B(core_v3_reg_48_), .Y(core__abc_22172_new_n2092_));
OR2X2 OR2X2_978 ( .A(core__abc_22172_new_n2091_), .B(core__abc_22172_new_n2095_), .Y(core__abc_22172_new_n2096_));
OR2X2 OR2X2_979 ( .A(core__abc_22172_new_n2097_), .B(core__abc_22172_new_n2098_), .Y(core__abc_22172_new_n2099_));
OR2X2 OR2X2_98 ( .A(_abc_19873_new_n1120_), .B(_abc_19873_new_n1123_), .Y(_abc_19873_new_n1124_));
OR2X2 OR2X2_980 ( .A(core__abc_22172_new_n2100_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n2101_));
OR2X2 OR2X2_981 ( .A(core_siphash_word1_we), .B(core_siphash_word_112_), .Y(core__abc_22172_new_n2102_));
OR2X2 OR2X2_982 ( .A(core_v1_reg_49_), .B(core_v0_reg_49_), .Y(core__abc_22172_new_n2107_));
OR2X2 OR2X2_983 ( .A(core_v2_reg_49_), .B(core_v3_reg_49_), .Y(core__abc_22172_new_n2110_));
OR2X2 OR2X2_984 ( .A(core__abc_22172_new_n2114_), .B(core__abc_22172_new_n2116_), .Y(core__abc_22172_new_n2117_));
OR2X2 OR2X2_985 ( .A(core__abc_22172_new_n2117_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n2118_));
OR2X2 OR2X2_986 ( .A(core_siphash_word1_we), .B(core_siphash_word_113_), .Y(core__abc_22172_new_n2119_));
OR2X2 OR2X2_987 ( .A(core_v1_reg_50_), .B(core_v0_reg_50_), .Y(core__abc_22172_new_n2122_));
OR2X2 OR2X2_988 ( .A(core_v2_reg_50_), .B(core_v3_reg_50_), .Y(core__abc_22172_new_n2126_));
OR2X2 OR2X2_989 ( .A(core__abc_22172_new_n2125_), .B(core__abc_22172_new_n2129_), .Y(core__abc_22172_new_n2130_));
OR2X2 OR2X2_99 ( .A(_abc_19873_new_n1124_), .B(_abc_19873_new_n1117_), .Y(_abc_19873_new_n1125_));
OR2X2 OR2X2_990 ( .A(core__abc_22172_new_n2131_), .B(core__abc_22172_new_n2132_), .Y(core__abc_22172_new_n2133_));
OR2X2 OR2X2_991 ( .A(core__abc_22172_new_n2134_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n2135_));
OR2X2 OR2X2_992 ( .A(core_siphash_word1_we), .B(core_siphash_word_114_), .Y(core__abc_22172_new_n2136_));
OR2X2 OR2X2_993 ( .A(core_v1_reg_51_), .B(core_v0_reg_51_), .Y(core__abc_22172_new_n2139_));
OR2X2 OR2X2_994 ( .A(core_v2_reg_51_), .B(core_v3_reg_51_), .Y(core__abc_22172_new_n2143_));
OR2X2 OR2X2_995 ( .A(core__abc_22172_new_n2142_), .B(core__abc_22172_new_n2146_), .Y(core__abc_22172_new_n2147_));
OR2X2 OR2X2_996 ( .A(core__abc_22172_new_n2148_), .B(core__abc_22172_new_n2149_), .Y(core__abc_22172_new_n2150_));
OR2X2 OR2X2_997 ( .A(core__abc_22172_new_n2151_), .B(core__abc_22172_new_n1256_), .Y(core__abc_22172_new_n2152_));
OR2X2 OR2X2_998 ( .A(core_siphash_word1_we), .B(core_siphash_word_115_), .Y(core__abc_22172_new_n2153_));
OR2X2 OR2X2_999 ( .A(core_v1_reg_52_), .B(core_v0_reg_52_), .Y(core__abc_22172_new_n2156_));


endmodule