module b06_reset(clock, RESET_G, nRESET_G, EQL, CONT_EQL, CC_MUX_REG_2_, CC_MUX_REG_1_, USCITE_REG_2_, USCITE_REG_1_, ENABLE_COUNT_REG, ACKOUT_REG);

output ACKOUT_REG;
output CC_MUX_REG_1_;
output CC_MUX_REG_2_;
input CONT_EQL;
output ENABLE_COUNT_REG;
input EQL;
input RESET_G;
wire STATE_REG_0_; 
wire STATE_REG_1_; 
wire STATE_REG_2_; 
output USCITE_REG_1_;
output USCITE_REG_2_;
wire _abc_317_new_n15_; 
wire _abc_317_new_n16_; 
wire _abc_317_new_n17_; 
wire _abc_317_new_n18_; 
wire _abc_317_new_n19_; 
wire _abc_317_new_n20_; 
wire _abc_317_new_n21_; 
wire _abc_317_new_n22_; 
wire _abc_317_new_n24_; 
wire _abc_317_new_n25_; 
wire _abc_317_new_n26_; 
wire _abc_317_new_n27_; 
wire _abc_317_new_n29_; 
wire _abc_317_new_n30_; 
wire _abc_317_new_n31_; 
wire _abc_317_new_n32_; 
wire _abc_317_new_n33_; 
wire _abc_317_new_n34_; 
wire _abc_317_new_n35_; 
wire _abc_317_new_n37_; 
wire _abc_317_new_n38_; 
wire _abc_317_new_n39_; 
wire _abc_317_new_n41_; 
wire _abc_317_new_n43_; 
wire _abc_317_new_n45_; 
wire _abc_317_new_n47_; 
wire _abc_317_new_n48_; 
wire _abc_317_new_n49_; 
wire _abc_317_new_n50_; 
wire _auto_iopadmap_cc_368_execute_355; 
wire _auto_iopadmap_cc_368_execute_357; 
wire _auto_iopadmap_cc_368_execute_359; 
wire _auto_iopadmap_cc_368_execute_363; 
wire _auto_iopadmap_cc_368_execute_365; 
input clock;
wire n22; 
wire n26; 
wire n31; 
wire n36; 
wire n41; 
wire n45; 
wire n49; 
wire n53; 
input nRESET_G;
AND2X2 AND2X2_1 ( .A(STATE_REG_1_), .B(EQL), .Y(_abc_317_new_n30_));
AND2X2 AND2X2_2 ( .A(STATE_REG_0_), .B(EQL), .Y(_abc_317_new_n34_));
AND2X2 AND2X2_3 ( .A(_abc_317_new_n30_), .B(_abc_317_new_n20_), .Y(_abc_317_new_n37_));
AOI21X1 AOI21X1_1 ( .A(_abc_317_new_n19_), .B(_abc_317_new_n21_), .C(_abc_317_new_n17_), .Y(_abc_317_new_n22_));
AOI21X1 AOI21X1_2 ( .A(_abc_317_new_n16_), .B(STATE_REG_2_), .C(_abc_317_new_n17_), .Y(_abc_317_new_n27_));
AOI21X1 AOI21X1_3 ( .A(STATE_REG_0_), .B(STATE_REG_2_), .C(_abc_317_new_n38_), .Y(_abc_317_new_n39_));
AOI21X1 AOI21X1_4 ( .A(_abc_317_new_n30_), .B(STATE_REG_2_), .C(_abc_317_new_n17_), .Y(_abc_317_new_n43_));
AOI22X1 AOI22X1_1 ( .A(_abc_317_new_n33_), .B(STATE_REG_1_), .C(_abc_317_new_n32_), .D(_abc_317_new_n34_), .Y(_abc_317_new_n35_));
AOI22X1 AOI22X1_2 ( .A(_abc_317_new_n20_), .B(_abc_317_new_n30_), .C(_abc_317_new_n18_), .D(_abc_317_new_n24_), .Y(_abc_317_new_n41_));
BUFX2 BUFX2_1 ( .A(_auto_iopadmap_cc_368_execute_355), .Y(ACKOUT_REG));
BUFX2 BUFX2_2 ( .A(_auto_iopadmap_cc_368_execute_357), .Y(CC_MUX_REG_1_));
BUFX2 BUFX2_3 ( .A(_auto_iopadmap_cc_368_execute_359), .Y(CC_MUX_REG_2_));
BUFX2 BUFX2_4 ( .A(_auto_iopadmap_cc_368_execute_355), .Y(ENABLE_COUNT_REG));
BUFX2 BUFX2_5 ( .A(_auto_iopadmap_cc_368_execute_363), .Y(USCITE_REG_1_));
BUFX2 BUFX2_6 ( .A(_auto_iopadmap_cc_368_execute_365), .Y(USCITE_REG_2_));
DFFPOSX1 DFFPOSX1_1 ( .CLK(clock), .D(n49), .Q(_auto_iopadmap_cc_368_execute_365));
DFFPOSX1 DFFPOSX1_2 ( .CLK(clock), .D(n41), .Q(_auto_iopadmap_cc_368_execute_359));
DFFPOSX1 DFFPOSX1_3 ( .CLK(clock), .D(n45), .Q(_auto_iopadmap_cc_368_execute_357));
DFFPOSX1 DFFPOSX1_4 ( .CLK(clock), .D(n22), .Q(_auto_iopadmap_cc_368_execute_355));
DFFPOSX1 DFFPOSX1_5 ( .CLK(clock), .D(n53), .Q(_auto_iopadmap_cc_368_execute_363));
DFFPOSX1 DFFPOSX1_6 ( .CLK(clock), .D(n26), .Q(STATE_REG_2_));
DFFPOSX1 DFFPOSX1_7 ( .CLK(clock), .D(n31), .Q(STATE_REG_1_));
DFFPOSX1 DFFPOSX1_8 ( .CLK(clock), .D(n36), .Q(STATE_REG_0_));
INVX1 INVX1_1 ( .A(EQL), .Y(_abc_317_new_n15_));
INVX1 INVX1_2 ( .A(STATE_REG_1_), .Y(_abc_317_new_n18_));
INVX1 INVX1_3 ( .A(STATE_REG_2_), .Y(_abc_317_new_n32_));
INVX1 INVX1_4 ( .A(CONT_EQL), .Y(_abc_317_new_n48_));
INVX2 INVX2_1 ( .A(nRESET_G), .Y(_abc_317_new_n17_));
INVX2 INVX2_2 ( .A(STATE_REG_0_), .Y(_abc_317_new_n20_));
NAND2X1 NAND2X1_1 ( .A(STATE_REG_1_), .B(_abc_317_new_n20_), .Y(_abc_317_new_n21_));
NAND2X1 NAND2X1_2 ( .A(_abc_317_new_n16_), .B(_abc_317_new_n22_), .Y(n36));
NAND2X1 NAND2X1_3 ( .A(_abc_317_new_n25_), .B(_abc_317_new_n24_), .Y(_abc_317_new_n26_));
NAND2X1 NAND2X1_4 ( .A(_abc_317_new_n26_), .B(_abc_317_new_n27_), .Y(n26));
NAND2X1 NAND2X1_5 ( .A(_abc_317_new_n27_), .B(_abc_317_new_n41_), .Y(n41));
NAND2X1 NAND2X1_6 ( .A(_abc_317_new_n29_), .B(_abc_317_new_n43_), .Y(n49));
NAND2X1 NAND2X1_7 ( .A(STATE_REG_0_), .B(STATE_REG_2_), .Y(_abc_317_new_n49_));
NAND3X1 NAND3X1_1 ( .A(_abc_317_new_n20_), .B(STATE_REG_2_), .C(_abc_317_new_n25_), .Y(_abc_317_new_n29_));
NAND3X1 NAND3X1_2 ( .A(_abc_317_new_n29_), .B(_abc_317_new_n31_), .C(_abc_317_new_n35_), .Y(n31));
NAND3X1 NAND3X1_3 ( .A(EQL), .B(nRESET_G), .C(_abc_317_new_n45_), .Y(n53));
NAND3X1 NAND3X1_4 ( .A(STATE_REG_1_), .B(_abc_317_new_n15_), .C(_abc_317_new_n33_), .Y(_abc_317_new_n47_));
NAND3X1 NAND3X1_5 ( .A(nRESET_G), .B(_abc_317_new_n50_), .C(_abc_317_new_n47_), .Y(n22));
NOR2X1 NOR2X1_1 ( .A(STATE_REG_2_), .B(_abc_317_new_n20_), .Y(_abc_317_new_n24_));
NOR2X1 NOR2X1_2 ( .A(STATE_REG_1_), .B(EQL), .Y(_abc_317_new_n25_));
NOR2X1 NOR2X1_3 ( .A(_abc_317_new_n17_), .B(_abc_317_new_n30_), .Y(_abc_317_new_n31_));
NOR2X1 NOR2X1_4 ( .A(STATE_REG_0_), .B(STATE_REG_2_), .Y(_abc_317_new_n33_));
OAI21X1 OAI21X1_1 ( .A(STATE_REG_1_), .B(STATE_REG_0_), .C(_abc_317_new_n15_), .Y(_abc_317_new_n16_));
OAI21X1 OAI21X1_2 ( .A(STATE_REG_0_), .B(STATE_REG_2_), .C(_abc_317_new_n18_), .Y(_abc_317_new_n19_));
OAI21X1 OAI21X1_3 ( .A(STATE_REG_0_), .B(STATE_REG_2_), .C(nRESET_G), .Y(_abc_317_new_n38_));
OAI21X1 OAI21X1_4 ( .A(_abc_317_new_n25_), .B(_abc_317_new_n37_), .C(_abc_317_new_n39_), .Y(n45));
OAI21X1 OAI21X1_5 ( .A(STATE_REG_2_), .B(_abc_317_new_n21_), .C(_abc_317_new_n19_), .Y(_abc_317_new_n45_));
OAI21X1 OAI21X1_6 ( .A(_abc_317_new_n18_), .B(_abc_317_new_n49_), .C(_abc_317_new_n48_), .Y(_abc_317_new_n50_));


endmodule