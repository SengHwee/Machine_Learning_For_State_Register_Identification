module spi_axi_master(CEB, SCLK, DATA, RST, CLK, axi_awready, axi_wready, axi_bvalid, axi_arready, axi_rvalid, \axi_rdata[0] , \axi_rdata[1] , \axi_rdata[2] , \axi_rdata[3] , \axi_rdata[4] , \axi_rdata[5] , \axi_rdata[6] , \axi_rdata[7] , \axi_rdata[8] , \axi_rdata[9] , \axi_rdata[10] , \axi_rdata[11] , \axi_rdata[12] , \axi_rdata[13] , \axi_rdata[14] , \axi_rdata[15] , \axi_rdata[16] , \axi_rdata[17] , \axi_rdata[18] , \axi_rdata[19] , \axi_rdata[20] , \axi_rdata[21] , \axi_rdata[22] , \axi_rdata[23] , \axi_rdata[24] , \axi_rdata[25] , \axi_rdata[26] , \axi_rdata[27] , \axi_rdata[28] , \axi_rdata[29] , \axi_rdata[30] , \axi_rdata[31] , DOUT, PICORV_RST, axi_awvalid, \axi_awaddr[0] , \axi_awaddr[1] , \axi_awaddr[2] , \axi_awaddr[3] , \axi_awaddr[4] , \axi_awaddr[5] , \axi_awaddr[6] , \axi_awaddr[7] , \axi_awaddr[8] , \axi_awaddr[9] , \axi_awaddr[10] , \axi_awaddr[11] , \axi_awaddr[12] , \axi_awaddr[13] , \axi_awaddr[14] , \axi_awaddr[15] , \axi_awaddr[16] , \axi_awaddr[17] , \axi_awaddr[18] , \axi_awaddr[19] , \axi_awaddr[20] , \axi_awaddr[21] , \axi_awaddr[22] , \axi_awaddr[23] , \axi_awaddr[24] , \axi_awaddr[25] , \axi_awaddr[26] , \axi_awaddr[27] , \axi_awaddr[28] , \axi_awaddr[29] , \axi_awaddr[30] , \axi_awaddr[31] , \axi_awprot[0] , \axi_awprot[1] , \axi_awprot[2] , axi_wvalid, \axi_wdata[0] , \axi_wdata[1] , \axi_wdata[2] , \axi_wdata[3] , \axi_wdata[4] , \axi_wdata[5] , \axi_wdata[6] , \axi_wdata[7] , \axi_wdata[8] , \axi_wdata[9] , \axi_wdata[10] , \axi_wdata[11] , \axi_wdata[12] , \axi_wdata[13] , \axi_wdata[14] , \axi_wdata[15] , \axi_wdata[16] , \axi_wdata[17] , \axi_wdata[18] , \axi_wdata[19] , \axi_wdata[20] , \axi_wdata[21] , \axi_wdata[22] , \axi_wdata[23] , \axi_wdata[24] , \axi_wdata[25] , \axi_wdata[26] , \axi_wdata[27] , \axi_wdata[28] , \axi_wdata[29] , \axi_wdata[30] , \axi_wdata[31] , \axi_wstrb[0] , \axi_wstrb[1] , \axi_wstrb[2] , \axi_wstrb[3] , axi_bready, axi_arvalid, \axi_araddr[0] , \axi_araddr[1] , \axi_araddr[2] , \axi_araddr[3] , \axi_araddr[4] , \axi_araddr[5] , \axi_araddr[6] , \axi_araddr[7] , \axi_araddr[8] , \axi_araddr[9] , \axi_araddr[10] , \axi_araddr[11] , \axi_araddr[12] , \axi_araddr[13] , \axi_araddr[14] , \axi_araddr[15] , \axi_araddr[16] , \axi_araddr[17] , \axi_araddr[18] , \axi_araddr[19] , \axi_araddr[20] , \axi_araddr[21] , \axi_araddr[22] , \axi_araddr[23] , \axi_araddr[24] , \axi_araddr[25] , \axi_araddr[26] , \axi_araddr[27] , \axi_araddr[28] , \axi_araddr[29] , \axi_araddr[30] , \axi_araddr[31] , \axi_arprot[0] , \axi_arprot[1] , \axi_arprot[2] , axi_rready);

wire A_ADDR_0_; 
wire A_ADDR_10_; 
wire A_ADDR_11_; 
wire A_ADDR_12_; 
wire A_ADDR_13_; 
wire A_ADDR_14_; 
wire A_ADDR_15_; 
wire A_ADDR_16_; 
wire A_ADDR_17_; 
wire A_ADDR_18_; 
wire A_ADDR_19_; 
wire A_ADDR_1_; 
wire A_ADDR_20_; 
wire A_ADDR_21_; 
wire A_ADDR_22_; 
wire A_ADDR_23_; 
wire A_ADDR_24_; 
wire A_ADDR_25_; 
wire A_ADDR_26_; 
wire A_ADDR_27_; 
wire A_ADDR_28_; 
wire A_ADDR_29_; 
wire A_ADDR_2_; 
wire A_ADDR_30_; 
wire A_ADDR_31_; 
wire A_ADDR_3_; 
wire A_ADDR_4_; 
wire A_ADDR_5_; 
wire A_ADDR_6_; 
wire A_ADDR_7_; 
wire A_ADDR_8_; 
wire A_ADDR_9_; 
input CEB;
input CLK;
input DATA;
output DOUT;
output PICORV_RST;
wire PICORV_RST_SPI; 
input RST;
input SCLK;
wire WDATA_0_; 
wire WDATA_10_; 
wire WDATA_11_; 
wire WDATA_12_; 
wire WDATA_13_; 
wire WDATA_14_; 
wire WDATA_15_; 
wire WDATA_16_; 
wire WDATA_17_; 
wire WDATA_18_; 
wire WDATA_19_; 
wire WDATA_1_; 
wire WDATA_20_; 
wire WDATA_21_; 
wire WDATA_22_; 
wire WDATA_23_; 
wire WDATA_24_; 
wire WDATA_25_; 
wire WDATA_26_; 
wire WDATA_27_; 
wire WDATA_28_; 
wire WDATA_29_; 
wire WDATA_2_; 
wire WDATA_30_; 
wire WDATA_31_; 
wire WDATA_3_; 
wire WDATA_4_; 
wire WDATA_5_; 
wire WDATA_6_; 
wire WDATA_7_; 
wire WDATA_8_; 
wire WDATA_9_; 
wire _0A_ADDR_31_0__0_; 
wire _0A_ADDR_31_0__10_; 
wire _0A_ADDR_31_0__11_; 
wire _0A_ADDR_31_0__12_; 
wire _0A_ADDR_31_0__13_; 
wire _0A_ADDR_31_0__14_; 
wire _0A_ADDR_31_0__15_; 
wire _0A_ADDR_31_0__16_; 
wire _0A_ADDR_31_0__17_; 
wire _0A_ADDR_31_0__18_; 
wire _0A_ADDR_31_0__19_; 
wire _0A_ADDR_31_0__1_; 
wire _0A_ADDR_31_0__20_; 
wire _0A_ADDR_31_0__21_; 
wire _0A_ADDR_31_0__22_; 
wire _0A_ADDR_31_0__23_; 
wire _0A_ADDR_31_0__24_; 
wire _0A_ADDR_31_0__25_; 
wire _0A_ADDR_31_0__26_; 
wire _0A_ADDR_31_0__27_; 
wire _0A_ADDR_31_0__28_; 
wire _0A_ADDR_31_0__29_; 
wire _0A_ADDR_31_0__2_; 
wire _0A_ADDR_31_0__30_; 
wire _0A_ADDR_31_0__31_; 
wire _0A_ADDR_31_0__3_; 
wire _0A_ADDR_31_0__4_; 
wire _0A_ADDR_31_0__5_; 
wire _0A_ADDR_31_0__6_; 
wire _0A_ADDR_31_0__7_; 
wire _0A_ADDR_31_0__8_; 
wire _0A_ADDR_31_0__9_; 
wire _0PICORV_RST_SPI_0_0_; 
wire _0WDATA_31_0__0_; 
wire _0WDATA_31_0__10_; 
wire _0WDATA_31_0__11_; 
wire _0WDATA_31_0__12_; 
wire _0WDATA_31_0__13_; 
wire _0WDATA_31_0__14_; 
wire _0WDATA_31_0__15_; 
wire _0WDATA_31_0__16_; 
wire _0WDATA_31_0__17_; 
wire _0WDATA_31_0__18_; 
wire _0WDATA_31_0__19_; 
wire _0WDATA_31_0__1_; 
wire _0WDATA_31_0__20_; 
wire _0WDATA_31_0__21_; 
wire _0WDATA_31_0__22_; 
wire _0WDATA_31_0__23_; 
wire _0WDATA_31_0__24_; 
wire _0WDATA_31_0__25_; 
wire _0WDATA_31_0__26_; 
wire _0WDATA_31_0__27_; 
wire _0WDATA_31_0__28_; 
wire _0WDATA_31_0__29_; 
wire _0WDATA_31_0__2_; 
wire _0WDATA_31_0__30_; 
wire _0WDATA_31_0__31_; 
wire _0WDATA_31_0__3_; 
wire _0WDATA_31_0__4_; 
wire _0WDATA_31_0__5_; 
wire _0WDATA_31_0__6_; 
wire _0WDATA_31_0__7_; 
wire _0WDATA_31_0__8_; 
wire _0WDATA_31_0__9_; 
wire _0bus_cap_31_0__0_; 
wire _0bus_cap_31_0__10_; 
wire _0bus_cap_31_0__11_; 
wire _0bus_cap_31_0__12_; 
wire _0bus_cap_31_0__13_; 
wire _0bus_cap_31_0__14_; 
wire _0bus_cap_31_0__15_; 
wire _0bus_cap_31_0__16_; 
wire _0bus_cap_31_0__17_; 
wire _0bus_cap_31_0__18_; 
wire _0bus_cap_31_0__19_; 
wire _0bus_cap_31_0__1_; 
wire _0bus_cap_31_0__20_; 
wire _0bus_cap_31_0__21_; 
wire _0bus_cap_31_0__22_; 
wire _0bus_cap_31_0__23_; 
wire _0bus_cap_31_0__24_; 
wire _0bus_cap_31_0__25_; 
wire _0bus_cap_31_0__26_; 
wire _0bus_cap_31_0__27_; 
wire _0bus_cap_31_0__28_; 
wire _0bus_cap_31_0__29_; 
wire _0bus_cap_31_0__2_; 
wire _0bus_cap_31_0__30_; 
wire _0bus_cap_31_0__31_; 
wire _0bus_cap_31_0__3_; 
wire _0bus_cap_31_0__4_; 
wire _0bus_cap_31_0__5_; 
wire _0bus_cap_31_0__6_; 
wire _0bus_cap_31_0__7_; 
wire _0bus_cap_31_0__8_; 
wire _0bus_cap_31_0__9_; 
wire _0counter_65_0__0_; 
wire _0counter_65_0__10_; 
wire _0counter_65_0__11_; 
wire _0counter_65_0__12_; 
wire _0counter_65_0__13_; 
wire _0counter_65_0__14_; 
wire _0counter_65_0__15_; 
wire _0counter_65_0__16_; 
wire _0counter_65_0__17_; 
wire _0counter_65_0__18_; 
wire _0counter_65_0__19_; 
wire _0counter_65_0__1_; 
wire _0counter_65_0__20_; 
wire _0counter_65_0__21_; 
wire _0counter_65_0__22_; 
wire _0counter_65_0__23_; 
wire _0counter_65_0__24_; 
wire _0counter_65_0__25_; 
wire _0counter_65_0__26_; 
wire _0counter_65_0__27_; 
wire _0counter_65_0__28_; 
wire _0counter_65_0__29_; 
wire _0counter_65_0__2_; 
wire _0counter_65_0__30_; 
wire _0counter_65_0__31_; 
wire _0counter_65_0__32_; 
wire _0counter_65_0__33_; 
wire _0counter_65_0__34_; 
wire _0counter_65_0__35_; 
wire _0counter_65_0__36_; 
wire _0counter_65_0__37_; 
wire _0counter_65_0__38_; 
wire _0counter_65_0__39_; 
wire _0counter_65_0__3_; 
wire _0counter_65_0__40_; 
wire _0counter_65_0__41_; 
wire _0counter_65_0__42_; 
wire _0counter_65_0__43_; 
wire _0counter_65_0__44_; 
wire _0counter_65_0__45_; 
wire _0counter_65_0__46_; 
wire _0counter_65_0__47_; 
wire _0counter_65_0__48_; 
wire _0counter_65_0__49_; 
wire _0counter_65_0__4_; 
wire _0counter_65_0__50_; 
wire _0counter_65_0__51_; 
wire _0counter_65_0__52_; 
wire _0counter_65_0__53_; 
wire _0counter_65_0__54_; 
wire _0counter_65_0__55_; 
wire _0counter_65_0__56_; 
wire _0counter_65_0__57_; 
wire _0counter_65_0__58_; 
wire _0counter_65_0__59_; 
wire _0counter_65_0__5_; 
wire _0counter_65_0__60_; 
wire _0counter_65_0__61_; 
wire _0counter_65_0__62_; 
wire _0counter_65_0__63_; 
wire _0counter_65_0__64_; 
wire _0counter_65_0__65_; 
wire _0counter_65_0__6_; 
wire _0counter_65_0__7_; 
wire _0counter_65_0__8_; 
wire _0counter_65_0__9_; 
wire _0fini_spi_0_0_; 
wire _0rdata_31_0__0_; 
wire _0rdata_31_0__10_; 
wire _0rdata_31_0__11_; 
wire _0rdata_31_0__12_; 
wire _0rdata_31_0__13_; 
wire _0rdata_31_0__14_; 
wire _0rdata_31_0__15_; 
wire _0rdata_31_0__16_; 
wire _0rdata_31_0__17_; 
wire _0rdata_31_0__18_; 
wire _0rdata_31_0__19_; 
wire _0rdata_31_0__1_; 
wire _0rdata_31_0__20_; 
wire _0rdata_31_0__21_; 
wire _0rdata_31_0__22_; 
wire _0rdata_31_0__23_; 
wire _0rdata_31_0__24_; 
wire _0rdata_31_0__25_; 
wire _0rdata_31_0__26_; 
wire _0rdata_31_0__27_; 
wire _0rdata_31_0__28_; 
wire _0rdata_31_0__29_; 
wire _0rdata_31_0__2_; 
wire _0rdata_31_0__30_; 
wire _0rdata_31_0__31_; 
wire _0rdata_31_0__3_; 
wire _0rdata_31_0__4_; 
wire _0rdata_31_0__5_; 
wire _0rdata_31_0__6_; 
wire _0rdata_31_0__7_; 
wire _0rdata_31_0__8_; 
wire _0rdata_31_0__9_; 
wire _0re_0_0_; 
wire _0sft_reg_65_0__0_; 
wire _0sft_reg_65_0__10_; 
wire _0sft_reg_65_0__11_; 
wire _0sft_reg_65_0__12_; 
wire _0sft_reg_65_0__13_; 
wire _0sft_reg_65_0__14_; 
wire _0sft_reg_65_0__15_; 
wire _0sft_reg_65_0__16_; 
wire _0sft_reg_65_0__17_; 
wire _0sft_reg_65_0__18_; 
wire _0sft_reg_65_0__19_; 
wire _0sft_reg_65_0__1_; 
wire _0sft_reg_65_0__20_; 
wire _0sft_reg_65_0__21_; 
wire _0sft_reg_65_0__22_; 
wire _0sft_reg_65_0__23_; 
wire _0sft_reg_65_0__24_; 
wire _0sft_reg_65_0__25_; 
wire _0sft_reg_65_0__26_; 
wire _0sft_reg_65_0__27_; 
wire _0sft_reg_65_0__28_; 
wire _0sft_reg_65_0__29_; 
wire _0sft_reg_65_0__2_; 
wire _0sft_reg_65_0__30_; 
wire _0sft_reg_65_0__3_; 
wire _0sft_reg_65_0__4_; 
wire _0sft_reg_65_0__5_; 
wire _0sft_reg_65_0__6_; 
wire _0sft_reg_65_0__7_; 
wire _0sft_reg_65_0__8_; 
wire _0sft_reg_65_0__9_; 
wire _0we_0_0_; 
wire _abc_2903_auto_fsm_map_cc_118_implement_pattern_cache_430; 
wire _abc_2903_auto_fsm_map_cc_118_implement_pattern_cache_479; 
wire _abc_2903_auto_fsm_map_cc_170_map_fsm_402_0_; 
wire _abc_2903_auto_fsm_map_cc_170_map_fsm_402_1_; 
wire _abc_2903_auto_fsm_map_cc_170_map_fsm_402_3_; 
wire _abc_2903_auto_fsm_map_cc_170_map_fsm_402_4_; 
wire _abc_2903_auto_fsm_map_cc_170_map_fsm_402_5_; 
wire _abc_2903_auto_fsm_map_cc_170_map_fsm_402_6_; 
wire _abc_2903_auto_fsm_map_cc_170_map_fsm_402_7_; 
wire _abc_4169_new_n1001_; 
wire _abc_4169_new_n1002_; 
wire _abc_4169_new_n1004_; 
wire _abc_4169_new_n1005_; 
wire _abc_4169_new_n1007_; 
wire _abc_4169_new_n1008_; 
wire _abc_4169_new_n1010_; 
wire _abc_4169_new_n1011_; 
wire _abc_4169_new_n1013_; 
wire _abc_4169_new_n1014_; 
wire _abc_4169_new_n1016_; 
wire _abc_4169_new_n1017_; 
wire _abc_4169_new_n1019_; 
wire _abc_4169_new_n1020_; 
wire _abc_4169_new_n1022_; 
wire _abc_4169_new_n1023_; 
wire _abc_4169_new_n1025_; 
wire _abc_4169_new_n1026_; 
wire _abc_4169_new_n1028_; 
wire _abc_4169_new_n1029_; 
wire _abc_4169_new_n1031_; 
wire _abc_4169_new_n1032_; 
wire _abc_4169_new_n1034_; 
wire _abc_4169_new_n1035_; 
wire _abc_4169_new_n1036_; 
wire _abc_4169_new_n1037_; 
wire _abc_4169_new_n1038_; 
wire _abc_4169_new_n1040_; 
wire _abc_4169_new_n1041_; 
wire _abc_4169_new_n1043_; 
wire _abc_4169_new_n1044_; 
wire _abc_4169_new_n1046_; 
wire _abc_4169_new_n1047_; 
wire _abc_4169_new_n1049_; 
wire _abc_4169_new_n1050_; 
wire _abc_4169_new_n1052_; 
wire _abc_4169_new_n1053_; 
wire _abc_4169_new_n1055_; 
wire _abc_4169_new_n1056_; 
wire _abc_4169_new_n1058_; 
wire _abc_4169_new_n1059_; 
wire _abc_4169_new_n1061_; 
wire _abc_4169_new_n1062_; 
wire _abc_4169_new_n1064_; 
wire _abc_4169_new_n1065_; 
wire _abc_4169_new_n1067_; 
wire _abc_4169_new_n1068_; 
wire _abc_4169_new_n1070_; 
wire _abc_4169_new_n1071_; 
wire _abc_4169_new_n1073_; 
wire _abc_4169_new_n1074_; 
wire _abc_4169_new_n1076_; 
wire _abc_4169_new_n1077_; 
wire _abc_4169_new_n1079_; 
wire _abc_4169_new_n1080_; 
wire _abc_4169_new_n1082_; 
wire _abc_4169_new_n1083_; 
wire _abc_4169_new_n1085_; 
wire _abc_4169_new_n1086_; 
wire _abc_4169_new_n1088_; 
wire _abc_4169_new_n1089_; 
wire _abc_4169_new_n1091_; 
wire _abc_4169_new_n1092_; 
wire _abc_4169_new_n1094_; 
wire _abc_4169_new_n1095_; 
wire _abc_4169_new_n1097_; 
wire _abc_4169_new_n1098_; 
wire _abc_4169_new_n1100_; 
wire _abc_4169_new_n1101_; 
wire _abc_4169_new_n1103_; 
wire _abc_4169_new_n1104_; 
wire _abc_4169_new_n1106_; 
wire _abc_4169_new_n1107_; 
wire _abc_4169_new_n1109_; 
wire _abc_4169_new_n1110_; 
wire _abc_4169_new_n1112_; 
wire _abc_4169_new_n1113_; 
wire _abc_4169_new_n1115_; 
wire _abc_4169_new_n1116_; 
wire _abc_4169_new_n1118_; 
wire _abc_4169_new_n1119_; 
wire _abc_4169_new_n1121_; 
wire _abc_4169_new_n1122_; 
wire _abc_4169_new_n1124_; 
wire _abc_4169_new_n1125_; 
wire _abc_4169_new_n1127_; 
wire _abc_4169_new_n1128_; 
wire _abc_4169_new_n1130_; 
wire _abc_4169_new_n1131_; 
wire _abc_4169_new_n1133_; 
wire _abc_4169_new_n1134_; 
wire _abc_4169_new_n1136_; 
wire _abc_4169_new_n1138_; 
wire _abc_4169_new_n1139_; 
wire _abc_4169_new_n1141_; 
wire _abc_4169_new_n1143_; 
wire _abc_4169_new_n1144_; 
wire _abc_4169_new_n1146_; 
wire _abc_4169_new_n1148_; 
wire _abc_4169_new_n1149_; 
wire _abc_4169_new_n1151_; 
wire _abc_4169_new_n1153_; 
wire _abc_4169_new_n1154_; 
wire _abc_4169_new_n1156_; 
wire _abc_4169_new_n1158_; 
wire _abc_4169_new_n1159_; 
wire _abc_4169_new_n1161_; 
wire _abc_4169_new_n1163_; 
wire _abc_4169_new_n1164_; 
wire _abc_4169_new_n1166_; 
wire _abc_4169_new_n1168_; 
wire _abc_4169_new_n1169_; 
wire _abc_4169_new_n1171_; 
wire _abc_4169_new_n1173_; 
wire _abc_4169_new_n1174_; 
wire _abc_4169_new_n1176_; 
wire _abc_4169_new_n1178_; 
wire _abc_4169_new_n1179_; 
wire _abc_4169_new_n1181_; 
wire _abc_4169_new_n1183_; 
wire _abc_4169_new_n1184_; 
wire _abc_4169_new_n1186_; 
wire _abc_4169_new_n1188_; 
wire _abc_4169_new_n1189_; 
wire _abc_4169_new_n1191_; 
wire _abc_4169_new_n1193_; 
wire _abc_4169_new_n1194_; 
wire _abc_4169_new_n1196_; 
wire _abc_4169_new_n1198_; 
wire _abc_4169_new_n1199_; 
wire _abc_4169_new_n1201_; 
wire _abc_4169_new_n1203_; 
wire _abc_4169_new_n1204_; 
wire _abc_4169_new_n1206_; 
wire _abc_4169_new_n1208_; 
wire _abc_4169_new_n1209_; 
wire _abc_4169_new_n1212_; 
wire _abc_4169_new_n1217_; 
wire _abc_4169_new_n1219_; 
wire _abc_4169_new_n1223_; 
wire _abc_4169_new_n1225_; 
wire _abc_4169_new_n1227_; 
wire _abc_4169_new_n1229_; 
wire _abc_4169_new_n1231_; 
wire _abc_4169_new_n1233_; 
wire _abc_4169_new_n1235_; 
wire _abc_4169_new_n1237_; 
wire _abc_4169_new_n1239_; 
wire _abc_4169_new_n1241_; 
wire _abc_4169_new_n1245_; 
wire _abc_4169_new_n1247_; 
wire _abc_4169_new_n1249_; 
wire _abc_4169_new_n1251_; 
wire _abc_4169_new_n1253_; 
wire _abc_4169_new_n1255_; 
wire _abc_4169_new_n1257_; 
wire _abc_4169_new_n1259_; 
wire _abc_4169_new_n1261_; 
wire _abc_4169_new_n1263_; 
wire _abc_4169_new_n1265_; 
wire _abc_4169_new_n1267_; 
wire _abc_4169_new_n1269_; 
wire _abc_4169_new_n1272_; 
wire _abc_4169_new_n1274_; 
wire _abc_4169_new_n1276_; 
wire _abc_4169_new_n1278_; 
wire _abc_4169_new_n1280_; 
wire _abc_4169_new_n1282_; 
wire _abc_4169_new_n1284_; 
wire _abc_4169_new_n1286_; 
wire _abc_4169_new_n1288_; 
wire _abc_4169_new_n1290_; 
wire _abc_4169_new_n1292_; 
wire _abc_4169_new_n1294_; 
wire _abc_4169_new_n1296_; 
wire _abc_4169_new_n1298_; 
wire _abc_4169_new_n1300_; 
wire _abc_4169_new_n1302_; 
wire _abc_4169_new_n1304_; 
wire _abc_4169_new_n1306_; 
wire _abc_4169_new_n1308_; 
wire _abc_4169_new_n1310_; 
wire _abc_4169_new_n1312_; 
wire _abc_4169_new_n1314_; 
wire _abc_4169_new_n1316_; 
wire _abc_4169_new_n1318_; 
wire _abc_4169_new_n1320_; 
wire _abc_4169_new_n1322_; 
wire _abc_4169_new_n1324_; 
wire _abc_4169_new_n1326_; 
wire _abc_4169_new_n1328_; 
wire _abc_4169_new_n1330_; 
wire _abc_4169_new_n1332_; 
wire _abc_4169_new_n1334_; 
wire _abc_4169_new_n1335_; 
wire _abc_4169_new_n1336_; 
wire _abc_4169_new_n1337_; 
wire _abc_4169_new_n1339_; 
wire _abc_4169_new_n1340_; 
wire _abc_4169_new_n1341_; 
wire _abc_4169_new_n1343_; 
wire _abc_4169_new_n1344_; 
wire _abc_4169_new_n1346_; 
wire _abc_4169_new_n1348_; 
wire _abc_4169_new_n558_; 
wire _abc_4169_new_n559_; 
wire _abc_4169_new_n560_; 
wire _abc_4169_new_n562_; 
wire _abc_4169_new_n564_; 
wire _abc_4169_new_n565_; 
wire _abc_4169_new_n566_; 
wire _abc_4169_new_n568_; 
wire _abc_4169_new_n569_; 
wire _abc_4169_new_n571_; 
wire _abc_4169_new_n572_; 
wire _abc_4169_new_n573_; 
wire _abc_4169_new_n574_; 
wire _abc_4169_new_n575_; 
wire _abc_4169_new_n576_; 
wire _abc_4169_new_n578_; 
wire _abc_4169_new_n579_; 
wire _abc_4169_new_n581_; 
wire _abc_4169_new_n583_; 
wire _abc_4169_new_n585_; 
wire _abc_4169_new_n586_; 
wire _abc_4169_new_n587_; 
wire _abc_4169_new_n589_; 
wire _abc_4169_new_n590_; 
wire _abc_4169_new_n591_; 
wire _abc_4169_new_n593_; 
wire _abc_4169_new_n594_; 
wire _abc_4169_new_n595_; 
wire _abc_4169_new_n597_; 
wire _abc_4169_new_n598_; 
wire _abc_4169_new_n599_; 
wire _abc_4169_new_n600_; 
wire _abc_4169_new_n601_; 
wire _abc_4169_new_n602_; 
wire _abc_4169_new_n603_; 
wire _abc_4169_new_n604_; 
wire _abc_4169_new_n605_; 
wire _abc_4169_new_n606_; 
wire _abc_4169_new_n607_; 
wire _abc_4169_new_n608_; 
wire _abc_4169_new_n609_; 
wire _abc_4169_new_n610_; 
wire _abc_4169_new_n611_; 
wire _abc_4169_new_n612_; 
wire _abc_4169_new_n613_; 
wire _abc_4169_new_n614_; 
wire _abc_4169_new_n615_; 
wire _abc_4169_new_n616_; 
wire _abc_4169_new_n617_; 
wire _abc_4169_new_n618_; 
wire _abc_4169_new_n619_; 
wire _abc_4169_new_n620_; 
wire _abc_4169_new_n621_; 
wire _abc_4169_new_n622_; 
wire _abc_4169_new_n623_; 
wire _abc_4169_new_n624_; 
wire _abc_4169_new_n625_; 
wire _abc_4169_new_n626_; 
wire _abc_4169_new_n627_; 
wire _abc_4169_new_n628_; 
wire _abc_4169_new_n629_; 
wire _abc_4169_new_n630_; 
wire _abc_4169_new_n631_; 
wire _abc_4169_new_n632_; 
wire _abc_4169_new_n633_; 
wire _abc_4169_new_n634_; 
wire _abc_4169_new_n635_; 
wire _abc_4169_new_n636_; 
wire _abc_4169_new_n637_; 
wire _abc_4169_new_n638_; 
wire _abc_4169_new_n639_; 
wire _abc_4169_new_n640_; 
wire _abc_4169_new_n641_; 
wire _abc_4169_new_n642_; 
wire _abc_4169_new_n643_; 
wire _abc_4169_new_n644_; 
wire _abc_4169_new_n645_; 
wire _abc_4169_new_n646_; 
wire _abc_4169_new_n648_; 
wire _abc_4169_new_n649_; 
wire _abc_4169_new_n650_; 
wire _abc_4169_new_n651_; 
wire _abc_4169_new_n652_; 
wire _abc_4169_new_n653_; 
wire _abc_4169_new_n654_; 
wire _abc_4169_new_n655_; 
wire _abc_4169_new_n656_; 
wire _abc_4169_new_n658_; 
wire _abc_4169_new_n659_; 
wire _abc_4169_new_n660_; 
wire _abc_4169_new_n661_; 
wire _abc_4169_new_n662_; 
wire _abc_4169_new_n663_; 
wire _abc_4169_new_n665_; 
wire _abc_4169_new_n666_; 
wire _abc_4169_new_n667_; 
wire _abc_4169_new_n668_; 
wire _abc_4169_new_n669_; 
wire _abc_4169_new_n671_; 
wire _abc_4169_new_n672_; 
wire _abc_4169_new_n673_; 
wire _abc_4169_new_n674_; 
wire _abc_4169_new_n675_; 
wire _abc_4169_new_n677_; 
wire _abc_4169_new_n678_; 
wire _abc_4169_new_n679_; 
wire _abc_4169_new_n680_; 
wire _abc_4169_new_n681_; 
wire _abc_4169_new_n683_; 
wire _abc_4169_new_n684_; 
wire _abc_4169_new_n685_; 
wire _abc_4169_new_n686_; 
wire _abc_4169_new_n687_; 
wire _abc_4169_new_n689_; 
wire _abc_4169_new_n690_; 
wire _abc_4169_new_n691_; 
wire _abc_4169_new_n692_; 
wire _abc_4169_new_n693_; 
wire _abc_4169_new_n695_; 
wire _abc_4169_new_n696_; 
wire _abc_4169_new_n697_; 
wire _abc_4169_new_n698_; 
wire _abc_4169_new_n699_; 
wire _abc_4169_new_n701_; 
wire _abc_4169_new_n702_; 
wire _abc_4169_new_n703_; 
wire _abc_4169_new_n704_; 
wire _abc_4169_new_n705_; 
wire _abc_4169_new_n707_; 
wire _abc_4169_new_n708_; 
wire _abc_4169_new_n709_; 
wire _abc_4169_new_n710_; 
wire _abc_4169_new_n711_; 
wire _abc_4169_new_n713_; 
wire _abc_4169_new_n714_; 
wire _abc_4169_new_n715_; 
wire _abc_4169_new_n716_; 
wire _abc_4169_new_n717_; 
wire _abc_4169_new_n719_; 
wire _abc_4169_new_n720_; 
wire _abc_4169_new_n721_; 
wire _abc_4169_new_n722_; 
wire _abc_4169_new_n723_; 
wire _abc_4169_new_n725_; 
wire _abc_4169_new_n726_; 
wire _abc_4169_new_n727_; 
wire _abc_4169_new_n728_; 
wire _abc_4169_new_n729_; 
wire _abc_4169_new_n731_; 
wire _abc_4169_new_n732_; 
wire _abc_4169_new_n733_; 
wire _abc_4169_new_n734_; 
wire _abc_4169_new_n735_; 
wire _abc_4169_new_n737_; 
wire _abc_4169_new_n738_; 
wire _abc_4169_new_n739_; 
wire _abc_4169_new_n740_; 
wire _abc_4169_new_n741_; 
wire _abc_4169_new_n743_; 
wire _abc_4169_new_n744_; 
wire _abc_4169_new_n745_; 
wire _abc_4169_new_n746_; 
wire _abc_4169_new_n747_; 
wire _abc_4169_new_n749_; 
wire _abc_4169_new_n750_; 
wire _abc_4169_new_n751_; 
wire _abc_4169_new_n752_; 
wire _abc_4169_new_n753_; 
wire _abc_4169_new_n755_; 
wire _abc_4169_new_n756_; 
wire _abc_4169_new_n757_; 
wire _abc_4169_new_n758_; 
wire _abc_4169_new_n759_; 
wire _abc_4169_new_n761_; 
wire _abc_4169_new_n762_; 
wire _abc_4169_new_n763_; 
wire _abc_4169_new_n764_; 
wire _abc_4169_new_n765_; 
wire _abc_4169_new_n767_; 
wire _abc_4169_new_n768_; 
wire _abc_4169_new_n769_; 
wire _abc_4169_new_n770_; 
wire _abc_4169_new_n771_; 
wire _abc_4169_new_n773_; 
wire _abc_4169_new_n774_; 
wire _abc_4169_new_n775_; 
wire _abc_4169_new_n776_; 
wire _abc_4169_new_n777_; 
wire _abc_4169_new_n779_; 
wire _abc_4169_new_n780_; 
wire _abc_4169_new_n781_; 
wire _abc_4169_new_n782_; 
wire _abc_4169_new_n783_; 
wire _abc_4169_new_n785_; 
wire _abc_4169_new_n786_; 
wire _abc_4169_new_n787_; 
wire _abc_4169_new_n788_; 
wire _abc_4169_new_n789_; 
wire _abc_4169_new_n791_; 
wire _abc_4169_new_n792_; 
wire _abc_4169_new_n793_; 
wire _abc_4169_new_n794_; 
wire _abc_4169_new_n795_; 
wire _abc_4169_new_n797_; 
wire _abc_4169_new_n798_; 
wire _abc_4169_new_n799_; 
wire _abc_4169_new_n800_; 
wire _abc_4169_new_n801_; 
wire _abc_4169_new_n803_; 
wire _abc_4169_new_n804_; 
wire _abc_4169_new_n805_; 
wire _abc_4169_new_n806_; 
wire _abc_4169_new_n807_; 
wire _abc_4169_new_n809_; 
wire _abc_4169_new_n810_; 
wire _abc_4169_new_n811_; 
wire _abc_4169_new_n812_; 
wire _abc_4169_new_n813_; 
wire _abc_4169_new_n815_; 
wire _abc_4169_new_n816_; 
wire _abc_4169_new_n817_; 
wire _abc_4169_new_n818_; 
wire _abc_4169_new_n819_; 
wire _abc_4169_new_n821_; 
wire _abc_4169_new_n822_; 
wire _abc_4169_new_n823_; 
wire _abc_4169_new_n824_; 
wire _abc_4169_new_n825_; 
wire _abc_4169_new_n827_; 
wire _abc_4169_new_n828_; 
wire _abc_4169_new_n829_; 
wire _abc_4169_new_n830_; 
wire _abc_4169_new_n831_; 
wire _abc_4169_new_n833_; 
wire _abc_4169_new_n834_; 
wire _abc_4169_new_n835_; 
wire _abc_4169_new_n836_; 
wire _abc_4169_new_n837_; 
wire _abc_4169_new_n839_; 
wire _abc_4169_new_n840_; 
wire _abc_4169_new_n841_; 
wire _abc_4169_new_n843_; 
wire _abc_4169_new_n844_; 
wire _abc_4169_new_n846_; 
wire _abc_4169_new_n847_; 
wire _abc_4169_new_n849_; 
wire _abc_4169_new_n850_; 
wire _abc_4169_new_n852_; 
wire _abc_4169_new_n853_; 
wire _abc_4169_new_n855_; 
wire _abc_4169_new_n856_; 
wire _abc_4169_new_n858_; 
wire _abc_4169_new_n859_; 
wire _abc_4169_new_n861_; 
wire _abc_4169_new_n862_; 
wire _abc_4169_new_n864_; 
wire _abc_4169_new_n865_; 
wire _abc_4169_new_n867_; 
wire _abc_4169_new_n868_; 
wire _abc_4169_new_n870_; 
wire _abc_4169_new_n871_; 
wire _abc_4169_new_n873_; 
wire _abc_4169_new_n874_; 
wire _abc_4169_new_n876_; 
wire _abc_4169_new_n877_; 
wire _abc_4169_new_n879_; 
wire _abc_4169_new_n880_; 
wire _abc_4169_new_n882_; 
wire _abc_4169_new_n883_; 
wire _abc_4169_new_n885_; 
wire _abc_4169_new_n886_; 
wire _abc_4169_new_n888_; 
wire _abc_4169_new_n889_; 
wire _abc_4169_new_n891_; 
wire _abc_4169_new_n892_; 
wire _abc_4169_new_n894_; 
wire _abc_4169_new_n895_; 
wire _abc_4169_new_n897_; 
wire _abc_4169_new_n898_; 
wire _abc_4169_new_n900_; 
wire _abc_4169_new_n901_; 
wire _abc_4169_new_n903_; 
wire _abc_4169_new_n904_; 
wire _abc_4169_new_n906_; 
wire _abc_4169_new_n907_; 
wire _abc_4169_new_n909_; 
wire _abc_4169_new_n910_; 
wire _abc_4169_new_n912_; 
wire _abc_4169_new_n913_; 
wire _abc_4169_new_n915_; 
wire _abc_4169_new_n916_; 
wire _abc_4169_new_n918_; 
wire _abc_4169_new_n919_; 
wire _abc_4169_new_n921_; 
wire _abc_4169_new_n922_; 
wire _abc_4169_new_n924_; 
wire _abc_4169_new_n925_; 
wire _abc_4169_new_n927_; 
wire _abc_4169_new_n928_; 
wire _abc_4169_new_n930_; 
wire _abc_4169_new_n931_; 
wire _abc_4169_new_n933_; 
wire _abc_4169_new_n934_; 
wire _abc_4169_new_n936_; 
wire _abc_4169_new_n937_; 
wire _abc_4169_new_n938_; 
wire _abc_4169_new_n939_; 
wire _abc_4169_new_n941_; 
wire _abc_4169_new_n942_; 
wire _abc_4169_new_n944_; 
wire _abc_4169_new_n945_; 
wire _abc_4169_new_n947_; 
wire _abc_4169_new_n948_; 
wire _abc_4169_new_n950_; 
wire _abc_4169_new_n951_; 
wire _abc_4169_new_n953_; 
wire _abc_4169_new_n954_; 
wire _abc_4169_new_n956_; 
wire _abc_4169_new_n957_; 
wire _abc_4169_new_n959_; 
wire _abc_4169_new_n960_; 
wire _abc_4169_new_n962_; 
wire _abc_4169_new_n963_; 
wire _abc_4169_new_n965_; 
wire _abc_4169_new_n966_; 
wire _abc_4169_new_n968_; 
wire _abc_4169_new_n969_; 
wire _abc_4169_new_n971_; 
wire _abc_4169_new_n972_; 
wire _abc_4169_new_n974_; 
wire _abc_4169_new_n975_; 
wire _abc_4169_new_n977_; 
wire _abc_4169_new_n978_; 
wire _abc_4169_new_n980_; 
wire _abc_4169_new_n981_; 
wire _abc_4169_new_n983_; 
wire _abc_4169_new_n984_; 
wire _abc_4169_new_n986_; 
wire _abc_4169_new_n987_; 
wire _abc_4169_new_n989_; 
wire _abc_4169_new_n990_; 
wire _abc_4169_new_n992_; 
wire _abc_4169_new_n993_; 
wire _abc_4169_new_n995_; 
wire _abc_4169_new_n996_; 
wire _abc_4169_new_n998_; 
wire _abc_4169_new_n999_; 
output \axi_araddr[0] ;
output \axi_araddr[10] ;
output \axi_araddr[11] ;
output \axi_araddr[12] ;
output \axi_araddr[13] ;
output \axi_araddr[14] ;
output \axi_araddr[15] ;
output \axi_araddr[16] ;
output \axi_araddr[17] ;
output \axi_araddr[18] ;
output \axi_araddr[19] ;
output \axi_araddr[1] ;
output \axi_araddr[20] ;
output \axi_araddr[21] ;
output \axi_araddr[22] ;
output \axi_araddr[23] ;
output \axi_araddr[24] ;
output \axi_araddr[25] ;
output \axi_araddr[26] ;
output \axi_araddr[27] ;
output \axi_araddr[28] ;
output \axi_araddr[29] ;
output \axi_araddr[2] ;
output \axi_araddr[30] ;
output \axi_araddr[31] ;
output \axi_araddr[3] ;
output \axi_araddr[4] ;
output \axi_araddr[5] ;
output \axi_araddr[6] ;
output \axi_araddr[7] ;
output \axi_araddr[8] ;
output \axi_araddr[9] ;
output \axi_arprot[0] ;
output \axi_arprot[1] ;
output \axi_arprot[2] ;
input axi_arready;
output axi_arvalid;
output \axi_awaddr[0] ;
output \axi_awaddr[10] ;
output \axi_awaddr[11] ;
output \axi_awaddr[12] ;
output \axi_awaddr[13] ;
output \axi_awaddr[14] ;
output \axi_awaddr[15] ;
output \axi_awaddr[16] ;
output \axi_awaddr[17] ;
output \axi_awaddr[18] ;
output \axi_awaddr[19] ;
output \axi_awaddr[1] ;
output \axi_awaddr[20] ;
output \axi_awaddr[21] ;
output \axi_awaddr[22] ;
output \axi_awaddr[23] ;
output \axi_awaddr[24] ;
output \axi_awaddr[25] ;
output \axi_awaddr[26] ;
output \axi_awaddr[27] ;
output \axi_awaddr[28] ;
output \axi_awaddr[29] ;
output \axi_awaddr[2] ;
output \axi_awaddr[30] ;
output \axi_awaddr[31] ;
output \axi_awaddr[3] ;
output \axi_awaddr[4] ;
output \axi_awaddr[5] ;
output \axi_awaddr[6] ;
output \axi_awaddr[7] ;
output \axi_awaddr[8] ;
output \axi_awaddr[9] ;
output \axi_awprot[0] ;
output \axi_awprot[1] ;
output \axi_awprot[2] ;
input axi_awready;
output axi_awvalid;
output axi_bready;
input axi_bvalid;
input \axi_rdata[0] ;
input \axi_rdata[10] ;
input \axi_rdata[11] ;
input \axi_rdata[12] ;
input \axi_rdata[13] ;
input \axi_rdata[14] ;
input \axi_rdata[15] ;
input \axi_rdata[16] ;
input \axi_rdata[17] ;
input \axi_rdata[18] ;
input \axi_rdata[19] ;
input \axi_rdata[1] ;
input \axi_rdata[20] ;
input \axi_rdata[21] ;
input \axi_rdata[22] ;
input \axi_rdata[23] ;
input \axi_rdata[24] ;
input \axi_rdata[25] ;
input \axi_rdata[26] ;
input \axi_rdata[27] ;
input \axi_rdata[28] ;
input \axi_rdata[29] ;
input \axi_rdata[2] ;
input \axi_rdata[30] ;
input \axi_rdata[31] ;
input \axi_rdata[3] ;
input \axi_rdata[4] ;
input \axi_rdata[5] ;
input \axi_rdata[6] ;
input \axi_rdata[7] ;
input \axi_rdata[8] ;
input \axi_rdata[9] ;
output axi_rready;
input axi_rvalid;
output \axi_wdata[0] ;
output \axi_wdata[10] ;
output \axi_wdata[11] ;
output \axi_wdata[12] ;
output \axi_wdata[13] ;
output \axi_wdata[14] ;
output \axi_wdata[15] ;
output \axi_wdata[16] ;
output \axi_wdata[17] ;
output \axi_wdata[18] ;
output \axi_wdata[19] ;
output \axi_wdata[1] ;
output \axi_wdata[20] ;
output \axi_wdata[21] ;
output \axi_wdata[22] ;
output \axi_wdata[23] ;
output \axi_wdata[24] ;
output \axi_wdata[25] ;
output \axi_wdata[26] ;
output \axi_wdata[27] ;
output \axi_wdata[28] ;
output \axi_wdata[29] ;
output \axi_wdata[2] ;
output \axi_wdata[30] ;
output \axi_wdata[31] ;
output \axi_wdata[3] ;
output \axi_wdata[4] ;
output \axi_wdata[5] ;
output \axi_wdata[6] ;
output \axi_wdata[7] ;
output \axi_wdata[8] ;
output \axi_wdata[9] ;
input axi_wready;
output \axi_wstrb[0] ;
output \axi_wstrb[1] ;
output \axi_wstrb[2] ;
output \axi_wstrb[3] ;
output axi_wvalid;
wire bus_cap_0_; 
wire bus_cap_10_; 
wire bus_cap_11_; 
wire bus_cap_12_; 
wire bus_cap_13_; 
wire bus_cap_14_; 
wire bus_cap_15_; 
wire bus_cap_16_; 
wire bus_cap_17_; 
wire bus_cap_18_; 
wire bus_cap_19_; 
wire bus_cap_1_; 
wire bus_cap_20_; 
wire bus_cap_21_; 
wire bus_cap_22_; 
wire bus_cap_23_; 
wire bus_cap_24_; 
wire bus_cap_25_; 
wire bus_cap_26_; 
wire bus_cap_27_; 
wire bus_cap_28_; 
wire bus_cap_29_; 
wire bus_cap_2_; 
wire bus_cap_30_; 
wire bus_cap_3_; 
wire bus_cap_4_; 
wire bus_cap_5_; 
wire bus_cap_6_; 
wire bus_cap_7_; 
wire bus_cap_8_; 
wire bus_cap_9_; 
wire bus_sync_axi_bus_ECLK1; 
wire bus_sync_axi_bus_EECLK1; 
wire bus_sync_axi_bus_NCLK2; 
wire bus_sync_axi_bus__0ECLK1_0_0_; 
wire bus_sync_axi_bus__0EECLK1_0_0_; 
wire bus_sync_axi_bus__0reg_data1_63_0__0_; 
wire bus_sync_axi_bus__0reg_data1_63_0__10_; 
wire bus_sync_axi_bus__0reg_data1_63_0__11_; 
wire bus_sync_axi_bus__0reg_data1_63_0__12_; 
wire bus_sync_axi_bus__0reg_data1_63_0__13_; 
wire bus_sync_axi_bus__0reg_data1_63_0__14_; 
wire bus_sync_axi_bus__0reg_data1_63_0__15_; 
wire bus_sync_axi_bus__0reg_data1_63_0__16_; 
wire bus_sync_axi_bus__0reg_data1_63_0__17_; 
wire bus_sync_axi_bus__0reg_data1_63_0__18_; 
wire bus_sync_axi_bus__0reg_data1_63_0__19_; 
wire bus_sync_axi_bus__0reg_data1_63_0__1_; 
wire bus_sync_axi_bus__0reg_data1_63_0__20_; 
wire bus_sync_axi_bus__0reg_data1_63_0__21_; 
wire bus_sync_axi_bus__0reg_data1_63_0__22_; 
wire bus_sync_axi_bus__0reg_data1_63_0__23_; 
wire bus_sync_axi_bus__0reg_data1_63_0__24_; 
wire bus_sync_axi_bus__0reg_data1_63_0__25_; 
wire bus_sync_axi_bus__0reg_data1_63_0__26_; 
wire bus_sync_axi_bus__0reg_data1_63_0__27_; 
wire bus_sync_axi_bus__0reg_data1_63_0__28_; 
wire bus_sync_axi_bus__0reg_data1_63_0__29_; 
wire bus_sync_axi_bus__0reg_data1_63_0__2_; 
wire bus_sync_axi_bus__0reg_data1_63_0__30_; 
wire bus_sync_axi_bus__0reg_data1_63_0__31_; 
wire bus_sync_axi_bus__0reg_data1_63_0__32_; 
wire bus_sync_axi_bus__0reg_data1_63_0__33_; 
wire bus_sync_axi_bus__0reg_data1_63_0__34_; 
wire bus_sync_axi_bus__0reg_data1_63_0__35_; 
wire bus_sync_axi_bus__0reg_data1_63_0__36_; 
wire bus_sync_axi_bus__0reg_data1_63_0__37_; 
wire bus_sync_axi_bus__0reg_data1_63_0__38_; 
wire bus_sync_axi_bus__0reg_data1_63_0__39_; 
wire bus_sync_axi_bus__0reg_data1_63_0__3_; 
wire bus_sync_axi_bus__0reg_data1_63_0__40_; 
wire bus_sync_axi_bus__0reg_data1_63_0__41_; 
wire bus_sync_axi_bus__0reg_data1_63_0__42_; 
wire bus_sync_axi_bus__0reg_data1_63_0__43_; 
wire bus_sync_axi_bus__0reg_data1_63_0__44_; 
wire bus_sync_axi_bus__0reg_data1_63_0__45_; 
wire bus_sync_axi_bus__0reg_data1_63_0__46_; 
wire bus_sync_axi_bus__0reg_data1_63_0__47_; 
wire bus_sync_axi_bus__0reg_data1_63_0__48_; 
wire bus_sync_axi_bus__0reg_data1_63_0__49_; 
wire bus_sync_axi_bus__0reg_data1_63_0__4_; 
wire bus_sync_axi_bus__0reg_data1_63_0__50_; 
wire bus_sync_axi_bus__0reg_data1_63_0__51_; 
wire bus_sync_axi_bus__0reg_data1_63_0__52_; 
wire bus_sync_axi_bus__0reg_data1_63_0__53_; 
wire bus_sync_axi_bus__0reg_data1_63_0__54_; 
wire bus_sync_axi_bus__0reg_data1_63_0__55_; 
wire bus_sync_axi_bus__0reg_data1_63_0__56_; 
wire bus_sync_axi_bus__0reg_data1_63_0__57_; 
wire bus_sync_axi_bus__0reg_data1_63_0__58_; 
wire bus_sync_axi_bus__0reg_data1_63_0__59_; 
wire bus_sync_axi_bus__0reg_data1_63_0__5_; 
wire bus_sync_axi_bus__0reg_data1_63_0__60_; 
wire bus_sync_axi_bus__0reg_data1_63_0__61_; 
wire bus_sync_axi_bus__0reg_data1_63_0__62_; 
wire bus_sync_axi_bus__0reg_data1_63_0__63_; 
wire bus_sync_axi_bus__0reg_data1_63_0__6_; 
wire bus_sync_axi_bus__0reg_data1_63_0__7_; 
wire bus_sync_axi_bus__0reg_data1_63_0__8_; 
wire bus_sync_axi_bus__0reg_data1_63_0__9_; 
wire bus_sync_axi_bus__0reg_data2_63_0__0_; 
wire bus_sync_axi_bus__0reg_data2_63_0__10_; 
wire bus_sync_axi_bus__0reg_data2_63_0__11_; 
wire bus_sync_axi_bus__0reg_data2_63_0__12_; 
wire bus_sync_axi_bus__0reg_data2_63_0__13_; 
wire bus_sync_axi_bus__0reg_data2_63_0__14_; 
wire bus_sync_axi_bus__0reg_data2_63_0__15_; 
wire bus_sync_axi_bus__0reg_data2_63_0__16_; 
wire bus_sync_axi_bus__0reg_data2_63_0__17_; 
wire bus_sync_axi_bus__0reg_data2_63_0__18_; 
wire bus_sync_axi_bus__0reg_data2_63_0__19_; 
wire bus_sync_axi_bus__0reg_data2_63_0__1_; 
wire bus_sync_axi_bus__0reg_data2_63_0__20_; 
wire bus_sync_axi_bus__0reg_data2_63_0__21_; 
wire bus_sync_axi_bus__0reg_data2_63_0__22_; 
wire bus_sync_axi_bus__0reg_data2_63_0__23_; 
wire bus_sync_axi_bus__0reg_data2_63_0__24_; 
wire bus_sync_axi_bus__0reg_data2_63_0__25_; 
wire bus_sync_axi_bus__0reg_data2_63_0__26_; 
wire bus_sync_axi_bus__0reg_data2_63_0__27_; 
wire bus_sync_axi_bus__0reg_data2_63_0__28_; 
wire bus_sync_axi_bus__0reg_data2_63_0__29_; 
wire bus_sync_axi_bus__0reg_data2_63_0__2_; 
wire bus_sync_axi_bus__0reg_data2_63_0__30_; 
wire bus_sync_axi_bus__0reg_data2_63_0__31_; 
wire bus_sync_axi_bus__0reg_data2_63_0__32_; 
wire bus_sync_axi_bus__0reg_data2_63_0__33_; 
wire bus_sync_axi_bus__0reg_data2_63_0__34_; 
wire bus_sync_axi_bus__0reg_data2_63_0__35_; 
wire bus_sync_axi_bus__0reg_data2_63_0__36_; 
wire bus_sync_axi_bus__0reg_data2_63_0__37_; 
wire bus_sync_axi_bus__0reg_data2_63_0__38_; 
wire bus_sync_axi_bus__0reg_data2_63_0__39_; 
wire bus_sync_axi_bus__0reg_data2_63_0__3_; 
wire bus_sync_axi_bus__0reg_data2_63_0__40_; 
wire bus_sync_axi_bus__0reg_data2_63_0__41_; 
wire bus_sync_axi_bus__0reg_data2_63_0__42_; 
wire bus_sync_axi_bus__0reg_data2_63_0__43_; 
wire bus_sync_axi_bus__0reg_data2_63_0__44_; 
wire bus_sync_axi_bus__0reg_data2_63_0__45_; 
wire bus_sync_axi_bus__0reg_data2_63_0__46_; 
wire bus_sync_axi_bus__0reg_data2_63_0__47_; 
wire bus_sync_axi_bus__0reg_data2_63_0__48_; 
wire bus_sync_axi_bus__0reg_data2_63_0__49_; 
wire bus_sync_axi_bus__0reg_data2_63_0__4_; 
wire bus_sync_axi_bus__0reg_data2_63_0__50_; 
wire bus_sync_axi_bus__0reg_data2_63_0__51_; 
wire bus_sync_axi_bus__0reg_data2_63_0__52_; 
wire bus_sync_axi_bus__0reg_data2_63_0__53_; 
wire bus_sync_axi_bus__0reg_data2_63_0__54_; 
wire bus_sync_axi_bus__0reg_data2_63_0__55_; 
wire bus_sync_axi_bus__0reg_data2_63_0__56_; 
wire bus_sync_axi_bus__0reg_data2_63_0__57_; 
wire bus_sync_axi_bus__0reg_data2_63_0__58_; 
wire bus_sync_axi_bus__0reg_data2_63_0__59_; 
wire bus_sync_axi_bus__0reg_data2_63_0__5_; 
wire bus_sync_axi_bus__0reg_data2_63_0__60_; 
wire bus_sync_axi_bus__0reg_data2_63_0__61_; 
wire bus_sync_axi_bus__0reg_data2_63_0__62_; 
wire bus_sync_axi_bus__0reg_data2_63_0__63_; 
wire bus_sync_axi_bus__0reg_data2_63_0__6_; 
wire bus_sync_axi_bus__0reg_data2_63_0__7_; 
wire bus_sync_axi_bus__0reg_data2_63_0__8_; 
wire bus_sync_axi_bus__0reg_data2_63_0__9_; 
wire bus_sync_axi_bus__0reg_data3_63_0__0_; 
wire bus_sync_axi_bus__0reg_data3_63_0__10_; 
wire bus_sync_axi_bus__0reg_data3_63_0__11_; 
wire bus_sync_axi_bus__0reg_data3_63_0__12_; 
wire bus_sync_axi_bus__0reg_data3_63_0__13_; 
wire bus_sync_axi_bus__0reg_data3_63_0__14_; 
wire bus_sync_axi_bus__0reg_data3_63_0__15_; 
wire bus_sync_axi_bus__0reg_data3_63_0__16_; 
wire bus_sync_axi_bus__0reg_data3_63_0__17_; 
wire bus_sync_axi_bus__0reg_data3_63_0__18_; 
wire bus_sync_axi_bus__0reg_data3_63_0__19_; 
wire bus_sync_axi_bus__0reg_data3_63_0__1_; 
wire bus_sync_axi_bus__0reg_data3_63_0__20_; 
wire bus_sync_axi_bus__0reg_data3_63_0__21_; 
wire bus_sync_axi_bus__0reg_data3_63_0__22_; 
wire bus_sync_axi_bus__0reg_data3_63_0__23_; 
wire bus_sync_axi_bus__0reg_data3_63_0__24_; 
wire bus_sync_axi_bus__0reg_data3_63_0__25_; 
wire bus_sync_axi_bus__0reg_data3_63_0__26_; 
wire bus_sync_axi_bus__0reg_data3_63_0__27_; 
wire bus_sync_axi_bus__0reg_data3_63_0__28_; 
wire bus_sync_axi_bus__0reg_data3_63_0__29_; 
wire bus_sync_axi_bus__0reg_data3_63_0__2_; 
wire bus_sync_axi_bus__0reg_data3_63_0__30_; 
wire bus_sync_axi_bus__0reg_data3_63_0__31_; 
wire bus_sync_axi_bus__0reg_data3_63_0__32_; 
wire bus_sync_axi_bus__0reg_data3_63_0__33_; 
wire bus_sync_axi_bus__0reg_data3_63_0__34_; 
wire bus_sync_axi_bus__0reg_data3_63_0__35_; 
wire bus_sync_axi_bus__0reg_data3_63_0__36_; 
wire bus_sync_axi_bus__0reg_data3_63_0__37_; 
wire bus_sync_axi_bus__0reg_data3_63_0__38_; 
wire bus_sync_axi_bus__0reg_data3_63_0__39_; 
wire bus_sync_axi_bus__0reg_data3_63_0__3_; 
wire bus_sync_axi_bus__0reg_data3_63_0__40_; 
wire bus_sync_axi_bus__0reg_data3_63_0__41_; 
wire bus_sync_axi_bus__0reg_data3_63_0__42_; 
wire bus_sync_axi_bus__0reg_data3_63_0__43_; 
wire bus_sync_axi_bus__0reg_data3_63_0__44_; 
wire bus_sync_axi_bus__0reg_data3_63_0__45_; 
wire bus_sync_axi_bus__0reg_data3_63_0__46_; 
wire bus_sync_axi_bus__0reg_data3_63_0__47_; 
wire bus_sync_axi_bus__0reg_data3_63_0__48_; 
wire bus_sync_axi_bus__0reg_data3_63_0__49_; 
wire bus_sync_axi_bus__0reg_data3_63_0__4_; 
wire bus_sync_axi_bus__0reg_data3_63_0__50_; 
wire bus_sync_axi_bus__0reg_data3_63_0__51_; 
wire bus_sync_axi_bus__0reg_data3_63_0__52_; 
wire bus_sync_axi_bus__0reg_data3_63_0__53_; 
wire bus_sync_axi_bus__0reg_data3_63_0__54_; 
wire bus_sync_axi_bus__0reg_data3_63_0__55_; 
wire bus_sync_axi_bus__0reg_data3_63_0__56_; 
wire bus_sync_axi_bus__0reg_data3_63_0__57_; 
wire bus_sync_axi_bus__0reg_data3_63_0__58_; 
wire bus_sync_axi_bus__0reg_data3_63_0__59_; 
wire bus_sync_axi_bus__0reg_data3_63_0__5_; 
wire bus_sync_axi_bus__0reg_data3_63_0__60_; 
wire bus_sync_axi_bus__0reg_data3_63_0__61_; 
wire bus_sync_axi_bus__0reg_data3_63_0__62_; 
wire bus_sync_axi_bus__0reg_data3_63_0__63_; 
wire bus_sync_axi_bus__0reg_data3_63_0__6_; 
wire bus_sync_axi_bus__0reg_data3_63_0__7_; 
wire bus_sync_axi_bus__0reg_data3_63_0__8_; 
wire bus_sync_axi_bus__0reg_data3_63_0__9_; 
wire bus_sync_axi_bus__abc_3843_new_n393_; 
wire bus_sync_axi_bus__abc_3843_new_n394_; 
wire bus_sync_axi_bus__abc_3843_new_n395_; 
wire bus_sync_axi_bus__abc_3843_new_n396_; 
wire bus_sync_axi_bus__abc_3843_new_n398_; 
wire bus_sync_axi_bus__abc_3843_new_n399_; 
wire bus_sync_axi_bus__abc_3843_new_n401_; 
wire bus_sync_axi_bus__abc_3843_new_n402_; 
wire bus_sync_axi_bus__abc_3843_new_n404_; 
wire bus_sync_axi_bus__abc_3843_new_n405_; 
wire bus_sync_axi_bus__abc_3843_new_n407_; 
wire bus_sync_axi_bus__abc_3843_new_n408_; 
wire bus_sync_axi_bus__abc_3843_new_n410_; 
wire bus_sync_axi_bus__abc_3843_new_n411_; 
wire bus_sync_axi_bus__abc_3843_new_n413_; 
wire bus_sync_axi_bus__abc_3843_new_n414_; 
wire bus_sync_axi_bus__abc_3843_new_n416_; 
wire bus_sync_axi_bus__abc_3843_new_n417_; 
wire bus_sync_axi_bus__abc_3843_new_n419_; 
wire bus_sync_axi_bus__abc_3843_new_n420_; 
wire bus_sync_axi_bus__abc_3843_new_n422_; 
wire bus_sync_axi_bus__abc_3843_new_n423_; 
wire bus_sync_axi_bus__abc_3843_new_n425_; 
wire bus_sync_axi_bus__abc_3843_new_n426_; 
wire bus_sync_axi_bus__abc_3843_new_n428_; 
wire bus_sync_axi_bus__abc_3843_new_n429_; 
wire bus_sync_axi_bus__abc_3843_new_n431_; 
wire bus_sync_axi_bus__abc_3843_new_n432_; 
wire bus_sync_axi_bus__abc_3843_new_n434_; 
wire bus_sync_axi_bus__abc_3843_new_n435_; 
wire bus_sync_axi_bus__abc_3843_new_n437_; 
wire bus_sync_axi_bus__abc_3843_new_n438_; 
wire bus_sync_axi_bus__abc_3843_new_n440_; 
wire bus_sync_axi_bus__abc_3843_new_n441_; 
wire bus_sync_axi_bus__abc_3843_new_n443_; 
wire bus_sync_axi_bus__abc_3843_new_n444_; 
wire bus_sync_axi_bus__abc_3843_new_n446_; 
wire bus_sync_axi_bus__abc_3843_new_n447_; 
wire bus_sync_axi_bus__abc_3843_new_n449_; 
wire bus_sync_axi_bus__abc_3843_new_n450_; 
wire bus_sync_axi_bus__abc_3843_new_n452_; 
wire bus_sync_axi_bus__abc_3843_new_n453_; 
wire bus_sync_axi_bus__abc_3843_new_n455_; 
wire bus_sync_axi_bus__abc_3843_new_n456_; 
wire bus_sync_axi_bus__abc_3843_new_n458_; 
wire bus_sync_axi_bus__abc_3843_new_n459_; 
wire bus_sync_axi_bus__abc_3843_new_n461_; 
wire bus_sync_axi_bus__abc_3843_new_n462_; 
wire bus_sync_axi_bus__abc_3843_new_n464_; 
wire bus_sync_axi_bus__abc_3843_new_n465_; 
wire bus_sync_axi_bus__abc_3843_new_n467_; 
wire bus_sync_axi_bus__abc_3843_new_n468_; 
wire bus_sync_axi_bus__abc_3843_new_n470_; 
wire bus_sync_axi_bus__abc_3843_new_n471_; 
wire bus_sync_axi_bus__abc_3843_new_n473_; 
wire bus_sync_axi_bus__abc_3843_new_n474_; 
wire bus_sync_axi_bus__abc_3843_new_n476_; 
wire bus_sync_axi_bus__abc_3843_new_n477_; 
wire bus_sync_axi_bus__abc_3843_new_n479_; 
wire bus_sync_axi_bus__abc_3843_new_n480_; 
wire bus_sync_axi_bus__abc_3843_new_n482_; 
wire bus_sync_axi_bus__abc_3843_new_n483_; 
wire bus_sync_axi_bus__abc_3843_new_n485_; 
wire bus_sync_axi_bus__abc_3843_new_n486_; 
wire bus_sync_axi_bus__abc_3843_new_n488_; 
wire bus_sync_axi_bus__abc_3843_new_n489_; 
wire bus_sync_axi_bus__abc_3843_new_n491_; 
wire bus_sync_axi_bus__abc_3843_new_n492_; 
wire bus_sync_axi_bus__abc_3843_new_n494_; 
wire bus_sync_axi_bus__abc_3843_new_n495_; 
wire bus_sync_axi_bus__abc_3843_new_n497_; 
wire bus_sync_axi_bus__abc_3843_new_n498_; 
wire bus_sync_axi_bus__abc_3843_new_n500_; 
wire bus_sync_axi_bus__abc_3843_new_n501_; 
wire bus_sync_axi_bus__abc_3843_new_n503_; 
wire bus_sync_axi_bus__abc_3843_new_n504_; 
wire bus_sync_axi_bus__abc_3843_new_n506_; 
wire bus_sync_axi_bus__abc_3843_new_n507_; 
wire bus_sync_axi_bus__abc_3843_new_n509_; 
wire bus_sync_axi_bus__abc_3843_new_n510_; 
wire bus_sync_axi_bus__abc_3843_new_n512_; 
wire bus_sync_axi_bus__abc_3843_new_n513_; 
wire bus_sync_axi_bus__abc_3843_new_n515_; 
wire bus_sync_axi_bus__abc_3843_new_n516_; 
wire bus_sync_axi_bus__abc_3843_new_n518_; 
wire bus_sync_axi_bus__abc_3843_new_n519_; 
wire bus_sync_axi_bus__abc_3843_new_n521_; 
wire bus_sync_axi_bus__abc_3843_new_n522_; 
wire bus_sync_axi_bus__abc_3843_new_n524_; 
wire bus_sync_axi_bus__abc_3843_new_n525_; 
wire bus_sync_axi_bus__abc_3843_new_n527_; 
wire bus_sync_axi_bus__abc_3843_new_n528_; 
wire bus_sync_axi_bus__abc_3843_new_n530_; 
wire bus_sync_axi_bus__abc_3843_new_n531_; 
wire bus_sync_axi_bus__abc_3843_new_n533_; 
wire bus_sync_axi_bus__abc_3843_new_n534_; 
wire bus_sync_axi_bus__abc_3843_new_n536_; 
wire bus_sync_axi_bus__abc_3843_new_n537_; 
wire bus_sync_axi_bus__abc_3843_new_n539_; 
wire bus_sync_axi_bus__abc_3843_new_n540_; 
wire bus_sync_axi_bus__abc_3843_new_n542_; 
wire bus_sync_axi_bus__abc_3843_new_n543_; 
wire bus_sync_axi_bus__abc_3843_new_n545_; 
wire bus_sync_axi_bus__abc_3843_new_n546_; 
wire bus_sync_axi_bus__abc_3843_new_n548_; 
wire bus_sync_axi_bus__abc_3843_new_n549_; 
wire bus_sync_axi_bus__abc_3843_new_n551_; 
wire bus_sync_axi_bus__abc_3843_new_n552_; 
wire bus_sync_axi_bus__abc_3843_new_n554_; 
wire bus_sync_axi_bus__abc_3843_new_n555_; 
wire bus_sync_axi_bus__abc_3843_new_n557_; 
wire bus_sync_axi_bus__abc_3843_new_n558_; 
wire bus_sync_axi_bus__abc_3843_new_n560_; 
wire bus_sync_axi_bus__abc_3843_new_n561_; 
wire bus_sync_axi_bus__abc_3843_new_n563_; 
wire bus_sync_axi_bus__abc_3843_new_n564_; 
wire bus_sync_axi_bus__abc_3843_new_n566_; 
wire bus_sync_axi_bus__abc_3843_new_n567_; 
wire bus_sync_axi_bus__abc_3843_new_n569_; 
wire bus_sync_axi_bus__abc_3843_new_n570_; 
wire bus_sync_axi_bus__abc_3843_new_n572_; 
wire bus_sync_axi_bus__abc_3843_new_n573_; 
wire bus_sync_axi_bus__abc_3843_new_n575_; 
wire bus_sync_axi_bus__abc_3843_new_n576_; 
wire bus_sync_axi_bus__abc_3843_new_n578_; 
wire bus_sync_axi_bus__abc_3843_new_n579_; 
wire bus_sync_axi_bus__abc_3843_new_n581_; 
wire bus_sync_axi_bus__abc_3843_new_n582_; 
wire bus_sync_axi_bus__abc_3843_new_n584_; 
wire bus_sync_axi_bus__abc_3843_new_n585_; 
wire bus_sync_axi_bus_reg_data1_0_; 
wire bus_sync_axi_bus_reg_data1_10_; 
wire bus_sync_axi_bus_reg_data1_11_; 
wire bus_sync_axi_bus_reg_data1_12_; 
wire bus_sync_axi_bus_reg_data1_13_; 
wire bus_sync_axi_bus_reg_data1_14_; 
wire bus_sync_axi_bus_reg_data1_15_; 
wire bus_sync_axi_bus_reg_data1_16_; 
wire bus_sync_axi_bus_reg_data1_17_; 
wire bus_sync_axi_bus_reg_data1_18_; 
wire bus_sync_axi_bus_reg_data1_19_; 
wire bus_sync_axi_bus_reg_data1_1_; 
wire bus_sync_axi_bus_reg_data1_20_; 
wire bus_sync_axi_bus_reg_data1_21_; 
wire bus_sync_axi_bus_reg_data1_22_; 
wire bus_sync_axi_bus_reg_data1_23_; 
wire bus_sync_axi_bus_reg_data1_24_; 
wire bus_sync_axi_bus_reg_data1_25_; 
wire bus_sync_axi_bus_reg_data1_26_; 
wire bus_sync_axi_bus_reg_data1_27_; 
wire bus_sync_axi_bus_reg_data1_28_; 
wire bus_sync_axi_bus_reg_data1_29_; 
wire bus_sync_axi_bus_reg_data1_2_; 
wire bus_sync_axi_bus_reg_data1_30_; 
wire bus_sync_axi_bus_reg_data1_31_; 
wire bus_sync_axi_bus_reg_data1_32_; 
wire bus_sync_axi_bus_reg_data1_33_; 
wire bus_sync_axi_bus_reg_data1_34_; 
wire bus_sync_axi_bus_reg_data1_35_; 
wire bus_sync_axi_bus_reg_data1_36_; 
wire bus_sync_axi_bus_reg_data1_37_; 
wire bus_sync_axi_bus_reg_data1_38_; 
wire bus_sync_axi_bus_reg_data1_39_; 
wire bus_sync_axi_bus_reg_data1_3_; 
wire bus_sync_axi_bus_reg_data1_40_; 
wire bus_sync_axi_bus_reg_data1_41_; 
wire bus_sync_axi_bus_reg_data1_42_; 
wire bus_sync_axi_bus_reg_data1_43_; 
wire bus_sync_axi_bus_reg_data1_44_; 
wire bus_sync_axi_bus_reg_data1_45_; 
wire bus_sync_axi_bus_reg_data1_46_; 
wire bus_sync_axi_bus_reg_data1_47_; 
wire bus_sync_axi_bus_reg_data1_48_; 
wire bus_sync_axi_bus_reg_data1_49_; 
wire bus_sync_axi_bus_reg_data1_4_; 
wire bus_sync_axi_bus_reg_data1_50_; 
wire bus_sync_axi_bus_reg_data1_51_; 
wire bus_sync_axi_bus_reg_data1_52_; 
wire bus_sync_axi_bus_reg_data1_53_; 
wire bus_sync_axi_bus_reg_data1_54_; 
wire bus_sync_axi_bus_reg_data1_55_; 
wire bus_sync_axi_bus_reg_data1_56_; 
wire bus_sync_axi_bus_reg_data1_57_; 
wire bus_sync_axi_bus_reg_data1_58_; 
wire bus_sync_axi_bus_reg_data1_59_; 
wire bus_sync_axi_bus_reg_data1_5_; 
wire bus_sync_axi_bus_reg_data1_60_; 
wire bus_sync_axi_bus_reg_data1_61_; 
wire bus_sync_axi_bus_reg_data1_62_; 
wire bus_sync_axi_bus_reg_data1_63_; 
wire bus_sync_axi_bus_reg_data1_6_; 
wire bus_sync_axi_bus_reg_data1_7_; 
wire bus_sync_axi_bus_reg_data1_8_; 
wire bus_sync_axi_bus_reg_data1_9_; 
wire bus_sync_axi_bus_reg_data2_0_; 
wire bus_sync_axi_bus_reg_data2_10_; 
wire bus_sync_axi_bus_reg_data2_11_; 
wire bus_sync_axi_bus_reg_data2_12_; 
wire bus_sync_axi_bus_reg_data2_13_; 
wire bus_sync_axi_bus_reg_data2_14_; 
wire bus_sync_axi_bus_reg_data2_15_; 
wire bus_sync_axi_bus_reg_data2_16_; 
wire bus_sync_axi_bus_reg_data2_17_; 
wire bus_sync_axi_bus_reg_data2_18_; 
wire bus_sync_axi_bus_reg_data2_19_; 
wire bus_sync_axi_bus_reg_data2_1_; 
wire bus_sync_axi_bus_reg_data2_20_; 
wire bus_sync_axi_bus_reg_data2_21_; 
wire bus_sync_axi_bus_reg_data2_22_; 
wire bus_sync_axi_bus_reg_data2_23_; 
wire bus_sync_axi_bus_reg_data2_24_; 
wire bus_sync_axi_bus_reg_data2_25_; 
wire bus_sync_axi_bus_reg_data2_26_; 
wire bus_sync_axi_bus_reg_data2_27_; 
wire bus_sync_axi_bus_reg_data2_28_; 
wire bus_sync_axi_bus_reg_data2_29_; 
wire bus_sync_axi_bus_reg_data2_2_; 
wire bus_sync_axi_bus_reg_data2_30_; 
wire bus_sync_axi_bus_reg_data2_31_; 
wire bus_sync_axi_bus_reg_data2_32_; 
wire bus_sync_axi_bus_reg_data2_33_; 
wire bus_sync_axi_bus_reg_data2_34_; 
wire bus_sync_axi_bus_reg_data2_35_; 
wire bus_sync_axi_bus_reg_data2_36_; 
wire bus_sync_axi_bus_reg_data2_37_; 
wire bus_sync_axi_bus_reg_data2_38_; 
wire bus_sync_axi_bus_reg_data2_39_; 
wire bus_sync_axi_bus_reg_data2_3_; 
wire bus_sync_axi_bus_reg_data2_40_; 
wire bus_sync_axi_bus_reg_data2_41_; 
wire bus_sync_axi_bus_reg_data2_42_; 
wire bus_sync_axi_bus_reg_data2_43_; 
wire bus_sync_axi_bus_reg_data2_44_; 
wire bus_sync_axi_bus_reg_data2_45_; 
wire bus_sync_axi_bus_reg_data2_46_; 
wire bus_sync_axi_bus_reg_data2_47_; 
wire bus_sync_axi_bus_reg_data2_48_; 
wire bus_sync_axi_bus_reg_data2_49_; 
wire bus_sync_axi_bus_reg_data2_4_; 
wire bus_sync_axi_bus_reg_data2_50_; 
wire bus_sync_axi_bus_reg_data2_51_; 
wire bus_sync_axi_bus_reg_data2_52_; 
wire bus_sync_axi_bus_reg_data2_53_; 
wire bus_sync_axi_bus_reg_data2_54_; 
wire bus_sync_axi_bus_reg_data2_55_; 
wire bus_sync_axi_bus_reg_data2_56_; 
wire bus_sync_axi_bus_reg_data2_57_; 
wire bus_sync_axi_bus_reg_data2_58_; 
wire bus_sync_axi_bus_reg_data2_59_; 
wire bus_sync_axi_bus_reg_data2_5_; 
wire bus_sync_axi_bus_reg_data2_60_; 
wire bus_sync_axi_bus_reg_data2_61_; 
wire bus_sync_axi_bus_reg_data2_62_; 
wire bus_sync_axi_bus_reg_data2_63_; 
wire bus_sync_axi_bus_reg_data2_6_; 
wire bus_sync_axi_bus_reg_data2_7_; 
wire bus_sync_axi_bus_reg_data2_8_; 
wire bus_sync_axi_bus_reg_data2_9_; 
wire bus_sync_rdata_ECLK2; 
wire bus_sync_rdata_EECLK2; 
wire bus_sync_rdata_NCLK1; 
wire bus_sync_rdata__0ECLK2_0_0_; 
wire bus_sync_rdata__0EECLK2_0_0_; 
wire bus_sync_rdata__0reg_data1_31_0__0_; 
wire bus_sync_rdata__0reg_data1_31_0__10_; 
wire bus_sync_rdata__0reg_data1_31_0__11_; 
wire bus_sync_rdata__0reg_data1_31_0__12_; 
wire bus_sync_rdata__0reg_data1_31_0__13_; 
wire bus_sync_rdata__0reg_data1_31_0__14_; 
wire bus_sync_rdata__0reg_data1_31_0__15_; 
wire bus_sync_rdata__0reg_data1_31_0__16_; 
wire bus_sync_rdata__0reg_data1_31_0__17_; 
wire bus_sync_rdata__0reg_data1_31_0__18_; 
wire bus_sync_rdata__0reg_data1_31_0__19_; 
wire bus_sync_rdata__0reg_data1_31_0__1_; 
wire bus_sync_rdata__0reg_data1_31_0__20_; 
wire bus_sync_rdata__0reg_data1_31_0__21_; 
wire bus_sync_rdata__0reg_data1_31_0__22_; 
wire bus_sync_rdata__0reg_data1_31_0__23_; 
wire bus_sync_rdata__0reg_data1_31_0__24_; 
wire bus_sync_rdata__0reg_data1_31_0__25_; 
wire bus_sync_rdata__0reg_data1_31_0__26_; 
wire bus_sync_rdata__0reg_data1_31_0__27_; 
wire bus_sync_rdata__0reg_data1_31_0__28_; 
wire bus_sync_rdata__0reg_data1_31_0__29_; 
wire bus_sync_rdata__0reg_data1_31_0__2_; 
wire bus_sync_rdata__0reg_data1_31_0__30_; 
wire bus_sync_rdata__0reg_data1_31_0__31_; 
wire bus_sync_rdata__0reg_data1_31_0__3_; 
wire bus_sync_rdata__0reg_data1_31_0__4_; 
wire bus_sync_rdata__0reg_data1_31_0__5_; 
wire bus_sync_rdata__0reg_data1_31_0__6_; 
wire bus_sync_rdata__0reg_data1_31_0__7_; 
wire bus_sync_rdata__0reg_data1_31_0__8_; 
wire bus_sync_rdata__0reg_data1_31_0__9_; 
wire bus_sync_rdata__0reg_data2_31_0__0_; 
wire bus_sync_rdata__0reg_data2_31_0__10_; 
wire bus_sync_rdata__0reg_data2_31_0__11_; 
wire bus_sync_rdata__0reg_data2_31_0__12_; 
wire bus_sync_rdata__0reg_data2_31_0__13_; 
wire bus_sync_rdata__0reg_data2_31_0__14_; 
wire bus_sync_rdata__0reg_data2_31_0__15_; 
wire bus_sync_rdata__0reg_data2_31_0__16_; 
wire bus_sync_rdata__0reg_data2_31_0__17_; 
wire bus_sync_rdata__0reg_data2_31_0__18_; 
wire bus_sync_rdata__0reg_data2_31_0__19_; 
wire bus_sync_rdata__0reg_data2_31_0__1_; 
wire bus_sync_rdata__0reg_data2_31_0__20_; 
wire bus_sync_rdata__0reg_data2_31_0__21_; 
wire bus_sync_rdata__0reg_data2_31_0__22_; 
wire bus_sync_rdata__0reg_data2_31_0__23_; 
wire bus_sync_rdata__0reg_data2_31_0__24_; 
wire bus_sync_rdata__0reg_data2_31_0__25_; 
wire bus_sync_rdata__0reg_data2_31_0__26_; 
wire bus_sync_rdata__0reg_data2_31_0__27_; 
wire bus_sync_rdata__0reg_data2_31_0__28_; 
wire bus_sync_rdata__0reg_data2_31_0__29_; 
wire bus_sync_rdata__0reg_data2_31_0__2_; 
wire bus_sync_rdata__0reg_data2_31_0__30_; 
wire bus_sync_rdata__0reg_data2_31_0__31_; 
wire bus_sync_rdata__0reg_data2_31_0__3_; 
wire bus_sync_rdata__0reg_data2_31_0__4_; 
wire bus_sync_rdata__0reg_data2_31_0__5_; 
wire bus_sync_rdata__0reg_data2_31_0__6_; 
wire bus_sync_rdata__0reg_data2_31_0__7_; 
wire bus_sync_rdata__0reg_data2_31_0__8_; 
wire bus_sync_rdata__0reg_data2_31_0__9_; 
wire bus_sync_rdata__0reg_data3_31_0__0_; 
wire bus_sync_rdata__0reg_data3_31_0__10_; 
wire bus_sync_rdata__0reg_data3_31_0__11_; 
wire bus_sync_rdata__0reg_data3_31_0__12_; 
wire bus_sync_rdata__0reg_data3_31_0__13_; 
wire bus_sync_rdata__0reg_data3_31_0__14_; 
wire bus_sync_rdata__0reg_data3_31_0__15_; 
wire bus_sync_rdata__0reg_data3_31_0__16_; 
wire bus_sync_rdata__0reg_data3_31_0__17_; 
wire bus_sync_rdata__0reg_data3_31_0__18_; 
wire bus_sync_rdata__0reg_data3_31_0__19_; 
wire bus_sync_rdata__0reg_data3_31_0__1_; 
wire bus_sync_rdata__0reg_data3_31_0__20_; 
wire bus_sync_rdata__0reg_data3_31_0__21_; 
wire bus_sync_rdata__0reg_data3_31_0__22_; 
wire bus_sync_rdata__0reg_data3_31_0__23_; 
wire bus_sync_rdata__0reg_data3_31_0__24_; 
wire bus_sync_rdata__0reg_data3_31_0__25_; 
wire bus_sync_rdata__0reg_data3_31_0__26_; 
wire bus_sync_rdata__0reg_data3_31_0__27_; 
wire bus_sync_rdata__0reg_data3_31_0__28_; 
wire bus_sync_rdata__0reg_data3_31_0__29_; 
wire bus_sync_rdata__0reg_data3_31_0__2_; 
wire bus_sync_rdata__0reg_data3_31_0__30_; 
wire bus_sync_rdata__0reg_data3_31_0__31_; 
wire bus_sync_rdata__0reg_data3_31_0__3_; 
wire bus_sync_rdata__0reg_data3_31_0__4_; 
wire bus_sync_rdata__0reg_data3_31_0__5_; 
wire bus_sync_rdata__0reg_data3_31_0__6_; 
wire bus_sync_rdata__0reg_data3_31_0__7_; 
wire bus_sync_rdata__0reg_data3_31_0__8_; 
wire bus_sync_rdata__0reg_data3_31_0__9_; 
wire bus_sync_rdata__abc_3651_new_n265_; 
wire bus_sync_rdata__abc_3651_new_n266_; 
wire bus_sync_rdata__abc_3651_new_n267_; 
wire bus_sync_rdata__abc_3651_new_n268_; 
wire bus_sync_rdata__abc_3651_new_n270_; 
wire bus_sync_rdata__abc_3651_new_n271_; 
wire bus_sync_rdata__abc_3651_new_n273_; 
wire bus_sync_rdata__abc_3651_new_n274_; 
wire bus_sync_rdata__abc_3651_new_n276_; 
wire bus_sync_rdata__abc_3651_new_n277_; 
wire bus_sync_rdata__abc_3651_new_n279_; 
wire bus_sync_rdata__abc_3651_new_n280_; 
wire bus_sync_rdata__abc_3651_new_n282_; 
wire bus_sync_rdata__abc_3651_new_n283_; 
wire bus_sync_rdata__abc_3651_new_n285_; 
wire bus_sync_rdata__abc_3651_new_n286_; 
wire bus_sync_rdata__abc_3651_new_n288_; 
wire bus_sync_rdata__abc_3651_new_n289_; 
wire bus_sync_rdata__abc_3651_new_n291_; 
wire bus_sync_rdata__abc_3651_new_n292_; 
wire bus_sync_rdata__abc_3651_new_n294_; 
wire bus_sync_rdata__abc_3651_new_n295_; 
wire bus_sync_rdata__abc_3651_new_n297_; 
wire bus_sync_rdata__abc_3651_new_n298_; 
wire bus_sync_rdata__abc_3651_new_n300_; 
wire bus_sync_rdata__abc_3651_new_n301_; 
wire bus_sync_rdata__abc_3651_new_n303_; 
wire bus_sync_rdata__abc_3651_new_n304_; 
wire bus_sync_rdata__abc_3651_new_n306_; 
wire bus_sync_rdata__abc_3651_new_n307_; 
wire bus_sync_rdata__abc_3651_new_n309_; 
wire bus_sync_rdata__abc_3651_new_n310_; 
wire bus_sync_rdata__abc_3651_new_n312_; 
wire bus_sync_rdata__abc_3651_new_n313_; 
wire bus_sync_rdata__abc_3651_new_n315_; 
wire bus_sync_rdata__abc_3651_new_n316_; 
wire bus_sync_rdata__abc_3651_new_n318_; 
wire bus_sync_rdata__abc_3651_new_n319_; 
wire bus_sync_rdata__abc_3651_new_n321_; 
wire bus_sync_rdata__abc_3651_new_n322_; 
wire bus_sync_rdata__abc_3651_new_n324_; 
wire bus_sync_rdata__abc_3651_new_n325_; 
wire bus_sync_rdata__abc_3651_new_n327_; 
wire bus_sync_rdata__abc_3651_new_n328_; 
wire bus_sync_rdata__abc_3651_new_n330_; 
wire bus_sync_rdata__abc_3651_new_n331_; 
wire bus_sync_rdata__abc_3651_new_n333_; 
wire bus_sync_rdata__abc_3651_new_n334_; 
wire bus_sync_rdata__abc_3651_new_n336_; 
wire bus_sync_rdata__abc_3651_new_n337_; 
wire bus_sync_rdata__abc_3651_new_n339_; 
wire bus_sync_rdata__abc_3651_new_n340_; 
wire bus_sync_rdata__abc_3651_new_n342_; 
wire bus_sync_rdata__abc_3651_new_n343_; 
wire bus_sync_rdata__abc_3651_new_n345_; 
wire bus_sync_rdata__abc_3651_new_n346_; 
wire bus_sync_rdata__abc_3651_new_n348_; 
wire bus_sync_rdata__abc_3651_new_n349_; 
wire bus_sync_rdata__abc_3651_new_n351_; 
wire bus_sync_rdata__abc_3651_new_n352_; 
wire bus_sync_rdata__abc_3651_new_n354_; 
wire bus_sync_rdata__abc_3651_new_n355_; 
wire bus_sync_rdata__abc_3651_new_n357_; 
wire bus_sync_rdata__abc_3651_new_n358_; 
wire bus_sync_rdata__abc_3651_new_n360_; 
wire bus_sync_rdata__abc_3651_new_n361_; 
wire bus_sync_rdata_data_in_0_; 
wire bus_sync_rdata_data_in_10_; 
wire bus_sync_rdata_data_in_11_; 
wire bus_sync_rdata_data_in_12_; 
wire bus_sync_rdata_data_in_13_; 
wire bus_sync_rdata_data_in_14_; 
wire bus_sync_rdata_data_in_15_; 
wire bus_sync_rdata_data_in_16_; 
wire bus_sync_rdata_data_in_17_; 
wire bus_sync_rdata_data_in_18_; 
wire bus_sync_rdata_data_in_19_; 
wire bus_sync_rdata_data_in_1_; 
wire bus_sync_rdata_data_in_20_; 
wire bus_sync_rdata_data_in_21_; 
wire bus_sync_rdata_data_in_22_; 
wire bus_sync_rdata_data_in_23_; 
wire bus_sync_rdata_data_in_24_; 
wire bus_sync_rdata_data_in_25_; 
wire bus_sync_rdata_data_in_26_; 
wire bus_sync_rdata_data_in_27_; 
wire bus_sync_rdata_data_in_28_; 
wire bus_sync_rdata_data_in_29_; 
wire bus_sync_rdata_data_in_2_; 
wire bus_sync_rdata_data_in_30_; 
wire bus_sync_rdata_data_in_31_; 
wire bus_sync_rdata_data_in_3_; 
wire bus_sync_rdata_data_in_4_; 
wire bus_sync_rdata_data_in_5_; 
wire bus_sync_rdata_data_in_6_; 
wire bus_sync_rdata_data_in_7_; 
wire bus_sync_rdata_data_in_8_; 
wire bus_sync_rdata_data_in_9_; 
wire bus_sync_rdata_data_out_0_; 
wire bus_sync_rdata_data_out_10_; 
wire bus_sync_rdata_data_out_11_; 
wire bus_sync_rdata_data_out_12_; 
wire bus_sync_rdata_data_out_13_; 
wire bus_sync_rdata_data_out_14_; 
wire bus_sync_rdata_data_out_15_; 
wire bus_sync_rdata_data_out_16_; 
wire bus_sync_rdata_data_out_17_; 
wire bus_sync_rdata_data_out_18_; 
wire bus_sync_rdata_data_out_19_; 
wire bus_sync_rdata_data_out_1_; 
wire bus_sync_rdata_data_out_20_; 
wire bus_sync_rdata_data_out_21_; 
wire bus_sync_rdata_data_out_22_; 
wire bus_sync_rdata_data_out_23_; 
wire bus_sync_rdata_data_out_24_; 
wire bus_sync_rdata_data_out_25_; 
wire bus_sync_rdata_data_out_26_; 
wire bus_sync_rdata_data_out_27_; 
wire bus_sync_rdata_data_out_28_; 
wire bus_sync_rdata_data_out_29_; 
wire bus_sync_rdata_data_out_2_; 
wire bus_sync_rdata_data_out_30_; 
wire bus_sync_rdata_data_out_31_; 
wire bus_sync_rdata_data_out_3_; 
wire bus_sync_rdata_data_out_4_; 
wire bus_sync_rdata_data_out_5_; 
wire bus_sync_rdata_data_out_6_; 
wire bus_sync_rdata_data_out_7_; 
wire bus_sync_rdata_data_out_8_; 
wire bus_sync_rdata_data_out_9_; 
wire bus_sync_rdata_reg_data1_0_; 
wire bus_sync_rdata_reg_data1_10_; 
wire bus_sync_rdata_reg_data1_11_; 
wire bus_sync_rdata_reg_data1_12_; 
wire bus_sync_rdata_reg_data1_13_; 
wire bus_sync_rdata_reg_data1_14_; 
wire bus_sync_rdata_reg_data1_15_; 
wire bus_sync_rdata_reg_data1_16_; 
wire bus_sync_rdata_reg_data1_17_; 
wire bus_sync_rdata_reg_data1_18_; 
wire bus_sync_rdata_reg_data1_19_; 
wire bus_sync_rdata_reg_data1_1_; 
wire bus_sync_rdata_reg_data1_20_; 
wire bus_sync_rdata_reg_data1_21_; 
wire bus_sync_rdata_reg_data1_22_; 
wire bus_sync_rdata_reg_data1_23_; 
wire bus_sync_rdata_reg_data1_24_; 
wire bus_sync_rdata_reg_data1_25_; 
wire bus_sync_rdata_reg_data1_26_; 
wire bus_sync_rdata_reg_data1_27_; 
wire bus_sync_rdata_reg_data1_28_; 
wire bus_sync_rdata_reg_data1_29_; 
wire bus_sync_rdata_reg_data1_2_; 
wire bus_sync_rdata_reg_data1_30_; 
wire bus_sync_rdata_reg_data1_31_; 
wire bus_sync_rdata_reg_data1_3_; 
wire bus_sync_rdata_reg_data1_4_; 
wire bus_sync_rdata_reg_data1_5_; 
wire bus_sync_rdata_reg_data1_6_; 
wire bus_sync_rdata_reg_data1_7_; 
wire bus_sync_rdata_reg_data1_8_; 
wire bus_sync_rdata_reg_data1_9_; 
wire bus_sync_rdata_reg_data2_0_; 
wire bus_sync_rdata_reg_data2_10_; 
wire bus_sync_rdata_reg_data2_11_; 
wire bus_sync_rdata_reg_data2_12_; 
wire bus_sync_rdata_reg_data2_13_; 
wire bus_sync_rdata_reg_data2_14_; 
wire bus_sync_rdata_reg_data2_15_; 
wire bus_sync_rdata_reg_data2_16_; 
wire bus_sync_rdata_reg_data2_17_; 
wire bus_sync_rdata_reg_data2_18_; 
wire bus_sync_rdata_reg_data2_19_; 
wire bus_sync_rdata_reg_data2_1_; 
wire bus_sync_rdata_reg_data2_20_; 
wire bus_sync_rdata_reg_data2_21_; 
wire bus_sync_rdata_reg_data2_22_; 
wire bus_sync_rdata_reg_data2_23_; 
wire bus_sync_rdata_reg_data2_24_; 
wire bus_sync_rdata_reg_data2_25_; 
wire bus_sync_rdata_reg_data2_26_; 
wire bus_sync_rdata_reg_data2_27_; 
wire bus_sync_rdata_reg_data2_28_; 
wire bus_sync_rdata_reg_data2_29_; 
wire bus_sync_rdata_reg_data2_2_; 
wire bus_sync_rdata_reg_data2_30_; 
wire bus_sync_rdata_reg_data2_31_; 
wire bus_sync_rdata_reg_data2_3_; 
wire bus_sync_rdata_reg_data2_4_; 
wire bus_sync_rdata_reg_data2_5_; 
wire bus_sync_rdata_reg_data2_6_; 
wire bus_sync_rdata_reg_data2_7_; 
wire bus_sync_rdata_reg_data2_8_; 
wire bus_sync_rdata_reg_data2_9_; 
wire bus_sync_state_machine_ECLK1; 
wire bus_sync_state_machine_EECLK1; 
wire bus_sync_state_machine_NCLK2; 
wire bus_sync_state_machine__0ECLK1_0_0_; 
wire bus_sync_state_machine__0EECLK1_0_0_; 
wire bus_sync_state_machine__0reg_data1_3_0__0_; 
wire bus_sync_state_machine__0reg_data1_3_0__1_; 
wire bus_sync_state_machine__0reg_data1_3_0__2_; 
wire bus_sync_state_machine__0reg_data1_3_0__3_; 
wire bus_sync_state_machine__0reg_data2_3_0__0_; 
wire bus_sync_state_machine__0reg_data2_3_0__1_; 
wire bus_sync_state_machine__0reg_data2_3_0__2_; 
wire bus_sync_state_machine__0reg_data2_3_0__3_; 
wire bus_sync_state_machine__0reg_data3_3_0__0_; 
wire bus_sync_state_machine__0reg_data3_3_0__1_; 
wire bus_sync_state_machine__0reg_data3_3_0__2_; 
wire bus_sync_state_machine__0reg_data3_3_0__3_; 
wire bus_sync_state_machine__abc_3817_new_n33_; 
wire bus_sync_state_machine__abc_3817_new_n34_; 
wire bus_sync_state_machine__abc_3817_new_n35_; 
wire bus_sync_state_machine__abc_3817_new_n36_; 
wire bus_sync_state_machine__abc_3817_new_n38_; 
wire bus_sync_state_machine__abc_3817_new_n39_; 
wire bus_sync_state_machine__abc_3817_new_n41_; 
wire bus_sync_state_machine__abc_3817_new_n42_; 
wire bus_sync_state_machine__abc_3817_new_n44_; 
wire bus_sync_state_machine__abc_3817_new_n45_; 
wire bus_sync_state_machine_reg_data1_0_; 
wire bus_sync_state_machine_reg_data1_1_; 
wire bus_sync_state_machine_reg_data1_2_; 
wire bus_sync_state_machine_reg_data1_3_; 
wire bus_sync_state_machine_reg_data2_0_; 
wire bus_sync_state_machine_reg_data2_1_; 
wire bus_sync_state_machine_reg_data2_2_; 
wire bus_sync_state_machine_reg_data2_3_; 
wire bus_sync_status_ECLK2; 
wire bus_sync_status_EECLK2; 
wire bus_sync_status_NCLK1; 
wire bus_sync_status__0ECLK2_0_0_; 
wire bus_sync_status__0EECLK2_0_0_; 
wire bus_sync_status__0reg_data1_2_0__0_; 
wire bus_sync_status__0reg_data1_2_0__1_; 
wire bus_sync_status__0reg_data1_2_0__2_; 
wire bus_sync_status__0reg_data2_2_0__0_; 
wire bus_sync_status__0reg_data2_2_0__1_; 
wire bus_sync_status__0reg_data2_2_0__2_; 
wire bus_sync_status__0reg_data3_2_0__0_; 
wire bus_sync_status__0reg_data3_2_0__1_; 
wire bus_sync_status__0reg_data3_2_0__2_; 
wire bus_sync_status__abc_3630_new_n27_; 
wire bus_sync_status__abc_3630_new_n28_; 
wire bus_sync_status__abc_3630_new_n29_; 
wire bus_sync_status__abc_3630_new_n30_; 
wire bus_sync_status__abc_3630_new_n32_; 
wire bus_sync_status__abc_3630_new_n33_; 
wire bus_sync_status__abc_3630_new_n35_; 
wire bus_sync_status__abc_3630_new_n36_; 
wire bus_sync_status_data_out_0_; 
wire bus_sync_status_data_out_1_; 
wire bus_sync_status_data_out_2_; 
wire bus_sync_status_reg_data1_0_; 
wire bus_sync_status_reg_data1_1_; 
wire bus_sync_status_reg_data1_2_; 
wire bus_sync_status_reg_data2_0_; 
wire bus_sync_status_reg_data2_1_; 
wire bus_sync_status_reg_data2_2_; 
wire busy; 
wire counter_0_; 
wire counter_10_; 
wire counter_11_; 
wire counter_12_; 
wire counter_13_; 
wire counter_14_; 
wire counter_15_; 
wire counter_16_; 
wire counter_17_; 
wire counter_18_; 
wire counter_19_; 
wire counter_1_; 
wire counter_20_; 
wire counter_21_; 
wire counter_22_; 
wire counter_23_; 
wire counter_24_; 
wire counter_25_; 
wire counter_26_; 
wire counter_27_; 
wire counter_28_; 
wire counter_29_; 
wire counter_2_; 
wire counter_30_; 
wire counter_31_; 
wire counter_32_; 
wire counter_33_; 
wire counter_34_; 
wire counter_35_; 
wire counter_36_; 
wire counter_37_; 
wire counter_38_; 
wire counter_39_; 
wire counter_3_; 
wire counter_40_; 
wire counter_41_; 
wire counter_42_; 
wire counter_43_; 
wire counter_44_; 
wire counter_45_; 
wire counter_46_; 
wire counter_47_; 
wire counter_48_; 
wire counter_49_; 
wire counter_4_; 
wire counter_50_; 
wire counter_51_; 
wire counter_52_; 
wire counter_53_; 
wire counter_54_; 
wire counter_55_; 
wire counter_56_; 
wire counter_57_; 
wire counter_58_; 
wire counter_59_; 
wire counter_5_; 
wire counter_60_; 
wire counter_61_; 
wire counter_62_; 
wire counter_63_; 
wire counter_64_; 
wire counter_65_; 
wire counter_6_; 
wire counter_7_; 
wire counter_8_; 
wire counter_9_; 
wire fini_spi; 
wire fini_spi_clk; 
wire re; 
wire re_clk; 
wire sft_reg_0_; 
wire sft_reg_10_; 
wire sft_reg_11_; 
wire sft_reg_12_; 
wire sft_reg_13_; 
wire sft_reg_14_; 
wire sft_reg_15_; 
wire sft_reg_16_; 
wire sft_reg_17_; 
wire sft_reg_18_; 
wire sft_reg_19_; 
wire sft_reg_1_; 
wire sft_reg_20_; 
wire sft_reg_21_; 
wire sft_reg_22_; 
wire sft_reg_23_; 
wire sft_reg_24_; 
wire sft_reg_25_; 
wire sft_reg_26_; 
wire sft_reg_27_; 
wire sft_reg_28_; 
wire sft_reg_29_; 
wire sft_reg_2_; 
wire sft_reg_30_; 
wire sft_reg_3_; 
wire sft_reg_4_; 
wire sft_reg_5_; 
wire sft_reg_6_; 
wire sft_reg_7_; 
wire sft_reg_8_; 
wire sft_reg_9_; 
wire state_0_; 
wire state_1_; 
wire state_3_; 
wire state_4_; 
wire state_5_; 
wire state_6_; 
wire state_7_; 
wire we; 
wire we_clk; 
AND2X2 AND2X2_1 ( .A(_abc_4169_new_n560_), .B(RST), .Y(_abc_2903_auto_fsm_map_cc_170_map_fsm_402_7_));
AND2X2 AND2X2_10 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_2_), .Y(bus_sync_axi_bus__0reg_data3_63_0__2_));
AND2X2 AND2X2_100 ( .A(RST), .B(WDATA_28_), .Y(bus_sync_axi_bus__0reg_data1_63_0__28_));
AND2X2 AND2X2_101 ( .A(RST), .B(WDATA_29_), .Y(bus_sync_axi_bus__0reg_data1_63_0__29_));
AND2X2 AND2X2_102 ( .A(RST), .B(WDATA_30_), .Y(bus_sync_axi_bus__0reg_data1_63_0__30_));
AND2X2 AND2X2_103 ( .A(RST), .B(WDATA_31_), .Y(bus_sync_axi_bus__0reg_data1_63_0__31_));
AND2X2 AND2X2_104 ( .A(RST), .B(A_ADDR_0_), .Y(bus_sync_axi_bus__0reg_data1_63_0__32_));
AND2X2 AND2X2_105 ( .A(RST), .B(A_ADDR_1_), .Y(bus_sync_axi_bus__0reg_data1_63_0__33_));
AND2X2 AND2X2_106 ( .A(RST), .B(A_ADDR_2_), .Y(bus_sync_axi_bus__0reg_data1_63_0__34_));
AND2X2 AND2X2_107 ( .A(RST), .B(A_ADDR_3_), .Y(bus_sync_axi_bus__0reg_data1_63_0__35_));
AND2X2 AND2X2_108 ( .A(RST), .B(A_ADDR_4_), .Y(bus_sync_axi_bus__0reg_data1_63_0__36_));
AND2X2 AND2X2_109 ( .A(RST), .B(A_ADDR_5_), .Y(bus_sync_axi_bus__0reg_data1_63_0__37_));
AND2X2 AND2X2_11 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_3_), .Y(bus_sync_axi_bus__0reg_data3_63_0__3_));
AND2X2 AND2X2_110 ( .A(RST), .B(A_ADDR_6_), .Y(bus_sync_axi_bus__0reg_data1_63_0__38_));
AND2X2 AND2X2_111 ( .A(RST), .B(A_ADDR_7_), .Y(bus_sync_axi_bus__0reg_data1_63_0__39_));
AND2X2 AND2X2_112 ( .A(RST), .B(A_ADDR_8_), .Y(bus_sync_axi_bus__0reg_data1_63_0__40_));
AND2X2 AND2X2_113 ( .A(RST), .B(A_ADDR_9_), .Y(bus_sync_axi_bus__0reg_data1_63_0__41_));
AND2X2 AND2X2_114 ( .A(RST), .B(A_ADDR_10_), .Y(bus_sync_axi_bus__0reg_data1_63_0__42_));
AND2X2 AND2X2_115 ( .A(RST), .B(A_ADDR_11_), .Y(bus_sync_axi_bus__0reg_data1_63_0__43_));
AND2X2 AND2X2_116 ( .A(RST), .B(A_ADDR_12_), .Y(bus_sync_axi_bus__0reg_data1_63_0__44_));
AND2X2 AND2X2_117 ( .A(RST), .B(A_ADDR_13_), .Y(bus_sync_axi_bus__0reg_data1_63_0__45_));
AND2X2 AND2X2_118 ( .A(RST), .B(A_ADDR_14_), .Y(bus_sync_axi_bus__0reg_data1_63_0__46_));
AND2X2 AND2X2_119 ( .A(RST), .B(A_ADDR_15_), .Y(bus_sync_axi_bus__0reg_data1_63_0__47_));
AND2X2 AND2X2_12 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_4_), .Y(bus_sync_axi_bus__0reg_data3_63_0__4_));
AND2X2 AND2X2_120 ( .A(RST), .B(A_ADDR_16_), .Y(bus_sync_axi_bus__0reg_data1_63_0__48_));
AND2X2 AND2X2_121 ( .A(RST), .B(A_ADDR_17_), .Y(bus_sync_axi_bus__0reg_data1_63_0__49_));
AND2X2 AND2X2_122 ( .A(RST), .B(A_ADDR_18_), .Y(bus_sync_axi_bus__0reg_data1_63_0__50_));
AND2X2 AND2X2_123 ( .A(RST), .B(A_ADDR_19_), .Y(bus_sync_axi_bus__0reg_data1_63_0__51_));
AND2X2 AND2X2_124 ( .A(RST), .B(A_ADDR_20_), .Y(bus_sync_axi_bus__0reg_data1_63_0__52_));
AND2X2 AND2X2_125 ( .A(RST), .B(A_ADDR_21_), .Y(bus_sync_axi_bus__0reg_data1_63_0__53_));
AND2X2 AND2X2_126 ( .A(RST), .B(A_ADDR_22_), .Y(bus_sync_axi_bus__0reg_data1_63_0__54_));
AND2X2 AND2X2_127 ( .A(RST), .B(A_ADDR_23_), .Y(bus_sync_axi_bus__0reg_data1_63_0__55_));
AND2X2 AND2X2_128 ( .A(RST), .B(A_ADDR_24_), .Y(bus_sync_axi_bus__0reg_data1_63_0__56_));
AND2X2 AND2X2_129 ( .A(RST), .B(A_ADDR_25_), .Y(bus_sync_axi_bus__0reg_data1_63_0__57_));
AND2X2 AND2X2_13 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_5_), .Y(bus_sync_axi_bus__0reg_data3_63_0__5_));
AND2X2 AND2X2_130 ( .A(RST), .B(A_ADDR_26_), .Y(bus_sync_axi_bus__0reg_data1_63_0__58_));
AND2X2 AND2X2_131 ( .A(RST), .B(A_ADDR_27_), .Y(bus_sync_axi_bus__0reg_data1_63_0__59_));
AND2X2 AND2X2_132 ( .A(RST), .B(A_ADDR_28_), .Y(bus_sync_axi_bus__0reg_data1_63_0__60_));
AND2X2 AND2X2_133 ( .A(RST), .B(A_ADDR_29_), .Y(bus_sync_axi_bus__0reg_data1_63_0__61_));
AND2X2 AND2X2_134 ( .A(RST), .B(A_ADDR_30_), .Y(bus_sync_axi_bus__0reg_data1_63_0__62_));
AND2X2 AND2X2_135 ( .A(RST), .B(A_ADDR_31_), .Y(bus_sync_axi_bus__0reg_data1_63_0__63_));
AND2X2 AND2X2_136 ( .A(RST), .B(SCLK), .Y(bus_sync_axi_bus__0ECLK1_0_0_));
AND2X2 AND2X2_137 ( .A(RST), .B(bus_sync_axi_bus_ECLK1), .Y(bus_sync_axi_bus__0EECLK1_0_0_));
AND2X2 AND2X2_138 ( .A(RST), .B(bus_sync_rdata_data_in_0_), .Y(bus_sync_rdata__0reg_data1_31_0__0_));
AND2X2 AND2X2_139 ( .A(RST), .B(bus_sync_rdata_data_in_1_), .Y(bus_sync_rdata__0reg_data1_31_0__1_));
AND2X2 AND2X2_14 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_6_), .Y(bus_sync_axi_bus__0reg_data3_63_0__6_));
AND2X2 AND2X2_140 ( .A(RST), .B(bus_sync_rdata_data_in_2_), .Y(bus_sync_rdata__0reg_data1_31_0__2_));
AND2X2 AND2X2_141 ( .A(RST), .B(bus_sync_rdata_data_in_3_), .Y(bus_sync_rdata__0reg_data1_31_0__3_));
AND2X2 AND2X2_142 ( .A(RST), .B(bus_sync_rdata_data_in_4_), .Y(bus_sync_rdata__0reg_data1_31_0__4_));
AND2X2 AND2X2_143 ( .A(RST), .B(bus_sync_rdata_data_in_5_), .Y(bus_sync_rdata__0reg_data1_31_0__5_));
AND2X2 AND2X2_144 ( .A(RST), .B(bus_sync_rdata_data_in_6_), .Y(bus_sync_rdata__0reg_data1_31_0__6_));
AND2X2 AND2X2_145 ( .A(RST), .B(bus_sync_rdata_data_in_7_), .Y(bus_sync_rdata__0reg_data1_31_0__7_));
AND2X2 AND2X2_146 ( .A(RST), .B(bus_sync_rdata_data_in_8_), .Y(bus_sync_rdata__0reg_data1_31_0__8_));
AND2X2 AND2X2_147 ( .A(RST), .B(bus_sync_rdata_data_in_9_), .Y(bus_sync_rdata__0reg_data1_31_0__9_));
AND2X2 AND2X2_148 ( .A(RST), .B(bus_sync_rdata_data_in_10_), .Y(bus_sync_rdata__0reg_data1_31_0__10_));
AND2X2 AND2X2_149 ( .A(RST), .B(bus_sync_rdata_data_in_11_), .Y(bus_sync_rdata__0reg_data1_31_0__11_));
AND2X2 AND2X2_15 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_7_), .Y(bus_sync_axi_bus__0reg_data3_63_0__7_));
AND2X2 AND2X2_150 ( .A(RST), .B(bus_sync_rdata_data_in_12_), .Y(bus_sync_rdata__0reg_data1_31_0__12_));
AND2X2 AND2X2_151 ( .A(RST), .B(bus_sync_rdata_data_in_13_), .Y(bus_sync_rdata__0reg_data1_31_0__13_));
AND2X2 AND2X2_152 ( .A(RST), .B(bus_sync_rdata_data_in_14_), .Y(bus_sync_rdata__0reg_data1_31_0__14_));
AND2X2 AND2X2_153 ( .A(RST), .B(bus_sync_rdata_data_in_15_), .Y(bus_sync_rdata__0reg_data1_31_0__15_));
AND2X2 AND2X2_154 ( .A(RST), .B(bus_sync_rdata_data_in_16_), .Y(bus_sync_rdata__0reg_data1_31_0__16_));
AND2X2 AND2X2_155 ( .A(RST), .B(bus_sync_rdata_data_in_17_), .Y(bus_sync_rdata__0reg_data1_31_0__17_));
AND2X2 AND2X2_156 ( .A(RST), .B(bus_sync_rdata_data_in_18_), .Y(bus_sync_rdata__0reg_data1_31_0__18_));
AND2X2 AND2X2_157 ( .A(RST), .B(bus_sync_rdata_data_in_19_), .Y(bus_sync_rdata__0reg_data1_31_0__19_));
AND2X2 AND2X2_158 ( .A(RST), .B(bus_sync_rdata_data_in_20_), .Y(bus_sync_rdata__0reg_data1_31_0__20_));
AND2X2 AND2X2_159 ( .A(RST), .B(bus_sync_rdata_data_in_21_), .Y(bus_sync_rdata__0reg_data1_31_0__21_));
AND2X2 AND2X2_16 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_8_), .Y(bus_sync_axi_bus__0reg_data3_63_0__8_));
AND2X2 AND2X2_160 ( .A(RST), .B(bus_sync_rdata_data_in_22_), .Y(bus_sync_rdata__0reg_data1_31_0__22_));
AND2X2 AND2X2_161 ( .A(RST), .B(bus_sync_rdata_data_in_23_), .Y(bus_sync_rdata__0reg_data1_31_0__23_));
AND2X2 AND2X2_162 ( .A(RST), .B(bus_sync_rdata_data_in_24_), .Y(bus_sync_rdata__0reg_data1_31_0__24_));
AND2X2 AND2X2_163 ( .A(RST), .B(bus_sync_rdata_data_in_25_), .Y(bus_sync_rdata__0reg_data1_31_0__25_));
AND2X2 AND2X2_164 ( .A(RST), .B(bus_sync_rdata_data_in_26_), .Y(bus_sync_rdata__0reg_data1_31_0__26_));
AND2X2 AND2X2_165 ( .A(RST), .B(bus_sync_rdata_data_in_27_), .Y(bus_sync_rdata__0reg_data1_31_0__27_));
AND2X2 AND2X2_166 ( .A(RST), .B(bus_sync_rdata_data_in_28_), .Y(bus_sync_rdata__0reg_data1_31_0__28_));
AND2X2 AND2X2_167 ( .A(RST), .B(bus_sync_rdata_data_in_29_), .Y(bus_sync_rdata__0reg_data1_31_0__29_));
AND2X2 AND2X2_168 ( .A(RST), .B(bus_sync_rdata_data_in_30_), .Y(bus_sync_rdata__0reg_data1_31_0__30_));
AND2X2 AND2X2_169 ( .A(RST), .B(bus_sync_rdata_data_in_31_), .Y(bus_sync_rdata__0reg_data1_31_0__31_));
AND2X2 AND2X2_17 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_9_), .Y(bus_sync_axi_bus__0reg_data3_63_0__9_));
AND2X2 AND2X2_170 ( .A(RST), .B(bus_sync_rdata_reg_data2_0_), .Y(bus_sync_rdata__0reg_data3_31_0__0_));
AND2X2 AND2X2_171 ( .A(RST), .B(bus_sync_rdata_reg_data2_1_), .Y(bus_sync_rdata__0reg_data3_31_0__1_));
AND2X2 AND2X2_172 ( .A(RST), .B(bus_sync_rdata_reg_data2_2_), .Y(bus_sync_rdata__0reg_data3_31_0__2_));
AND2X2 AND2X2_173 ( .A(RST), .B(bus_sync_rdata_reg_data2_3_), .Y(bus_sync_rdata__0reg_data3_31_0__3_));
AND2X2 AND2X2_174 ( .A(RST), .B(bus_sync_rdata_reg_data2_4_), .Y(bus_sync_rdata__0reg_data3_31_0__4_));
AND2X2 AND2X2_175 ( .A(RST), .B(bus_sync_rdata_reg_data2_5_), .Y(bus_sync_rdata__0reg_data3_31_0__5_));
AND2X2 AND2X2_176 ( .A(RST), .B(bus_sync_rdata_reg_data2_6_), .Y(bus_sync_rdata__0reg_data3_31_0__6_));
AND2X2 AND2X2_177 ( .A(RST), .B(bus_sync_rdata_reg_data2_7_), .Y(bus_sync_rdata__0reg_data3_31_0__7_));
AND2X2 AND2X2_178 ( .A(RST), .B(bus_sync_rdata_reg_data2_8_), .Y(bus_sync_rdata__0reg_data3_31_0__8_));
AND2X2 AND2X2_179 ( .A(RST), .B(bus_sync_rdata_reg_data2_9_), .Y(bus_sync_rdata__0reg_data3_31_0__9_));
AND2X2 AND2X2_18 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_10_), .Y(bus_sync_axi_bus__0reg_data3_63_0__10_));
AND2X2 AND2X2_180 ( .A(RST), .B(bus_sync_rdata_reg_data2_10_), .Y(bus_sync_rdata__0reg_data3_31_0__10_));
AND2X2 AND2X2_181 ( .A(RST), .B(bus_sync_rdata_reg_data2_11_), .Y(bus_sync_rdata__0reg_data3_31_0__11_));
AND2X2 AND2X2_182 ( .A(RST), .B(bus_sync_rdata_reg_data2_12_), .Y(bus_sync_rdata__0reg_data3_31_0__12_));
AND2X2 AND2X2_183 ( .A(RST), .B(bus_sync_rdata_reg_data2_13_), .Y(bus_sync_rdata__0reg_data3_31_0__13_));
AND2X2 AND2X2_184 ( .A(RST), .B(bus_sync_rdata_reg_data2_14_), .Y(bus_sync_rdata__0reg_data3_31_0__14_));
AND2X2 AND2X2_185 ( .A(RST), .B(bus_sync_rdata_reg_data2_15_), .Y(bus_sync_rdata__0reg_data3_31_0__15_));
AND2X2 AND2X2_186 ( .A(RST), .B(bus_sync_rdata_reg_data2_16_), .Y(bus_sync_rdata__0reg_data3_31_0__16_));
AND2X2 AND2X2_187 ( .A(RST), .B(bus_sync_rdata_reg_data2_17_), .Y(bus_sync_rdata__0reg_data3_31_0__17_));
AND2X2 AND2X2_188 ( .A(RST), .B(bus_sync_rdata_reg_data2_18_), .Y(bus_sync_rdata__0reg_data3_31_0__18_));
AND2X2 AND2X2_189 ( .A(RST), .B(bus_sync_rdata_reg_data2_19_), .Y(bus_sync_rdata__0reg_data3_31_0__19_));
AND2X2 AND2X2_19 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_11_), .Y(bus_sync_axi_bus__0reg_data3_63_0__11_));
AND2X2 AND2X2_190 ( .A(RST), .B(bus_sync_rdata_reg_data2_20_), .Y(bus_sync_rdata__0reg_data3_31_0__20_));
AND2X2 AND2X2_191 ( .A(RST), .B(bus_sync_rdata_reg_data2_21_), .Y(bus_sync_rdata__0reg_data3_31_0__21_));
AND2X2 AND2X2_192 ( .A(RST), .B(bus_sync_rdata_reg_data2_22_), .Y(bus_sync_rdata__0reg_data3_31_0__22_));
AND2X2 AND2X2_193 ( .A(RST), .B(bus_sync_rdata_reg_data2_23_), .Y(bus_sync_rdata__0reg_data3_31_0__23_));
AND2X2 AND2X2_194 ( .A(RST), .B(bus_sync_rdata_reg_data2_24_), .Y(bus_sync_rdata__0reg_data3_31_0__24_));
AND2X2 AND2X2_195 ( .A(RST), .B(bus_sync_rdata_reg_data2_25_), .Y(bus_sync_rdata__0reg_data3_31_0__25_));
AND2X2 AND2X2_196 ( .A(RST), .B(bus_sync_rdata_reg_data2_26_), .Y(bus_sync_rdata__0reg_data3_31_0__26_));
AND2X2 AND2X2_197 ( .A(RST), .B(bus_sync_rdata_reg_data2_27_), .Y(bus_sync_rdata__0reg_data3_31_0__27_));
AND2X2 AND2X2_198 ( .A(RST), .B(bus_sync_rdata_reg_data2_28_), .Y(bus_sync_rdata__0reg_data3_31_0__28_));
AND2X2 AND2X2_199 ( .A(RST), .B(bus_sync_rdata_reg_data2_29_), .Y(bus_sync_rdata__0reg_data3_31_0__29_));
AND2X2 AND2X2_2 ( .A(_abc_4169_new_n598_), .B(bus_sync_status_data_out_0_), .Y(_abc_4169_new_n643_));
AND2X2 AND2X2_20 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_12_), .Y(bus_sync_axi_bus__0reg_data3_63_0__12_));
AND2X2 AND2X2_200 ( .A(RST), .B(bus_sync_rdata_reg_data2_30_), .Y(bus_sync_rdata__0reg_data3_31_0__30_));
AND2X2 AND2X2_201 ( .A(RST), .B(bus_sync_rdata_reg_data2_31_), .Y(bus_sync_rdata__0reg_data3_31_0__31_));
AND2X2 AND2X2_202 ( .A(RST), .B(SCLK), .Y(bus_sync_rdata__0ECLK2_0_0_));
AND2X2 AND2X2_203 ( .A(RST), .B(bus_sync_rdata_ECLK2), .Y(bus_sync_rdata__0EECLK2_0_0_));
AND2X2 AND2X2_204 ( .A(RST), .B(bus_sync_state_machine_reg_data2_0_), .Y(bus_sync_state_machine__0reg_data3_3_0__0_));
AND2X2 AND2X2_205 ( .A(RST), .B(bus_sync_state_machine_reg_data2_1_), .Y(bus_sync_state_machine__0reg_data3_3_0__1_));
AND2X2 AND2X2_206 ( .A(RST), .B(bus_sync_state_machine_reg_data2_2_), .Y(bus_sync_state_machine__0reg_data3_3_0__2_));
AND2X2 AND2X2_207 ( .A(RST), .B(bus_sync_state_machine_reg_data2_3_), .Y(bus_sync_state_machine__0reg_data3_3_0__3_));
AND2X2 AND2X2_208 ( .A(RST), .B(fini_spi), .Y(bus_sync_state_machine__0reg_data1_3_0__0_));
AND2X2 AND2X2_209 ( .A(RST), .B(re), .Y(bus_sync_state_machine__0reg_data1_3_0__1_));
AND2X2 AND2X2_21 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_13_), .Y(bus_sync_axi_bus__0reg_data3_63_0__13_));
AND2X2 AND2X2_210 ( .A(RST), .B(we), .Y(bus_sync_state_machine__0reg_data1_3_0__2_));
AND2X2 AND2X2_211 ( .A(RST), .B(PICORV_RST_SPI), .Y(bus_sync_state_machine__0reg_data1_3_0__3_));
AND2X2 AND2X2_212 ( .A(RST), .B(SCLK), .Y(bus_sync_state_machine__0ECLK1_0_0_));
AND2X2 AND2X2_213 ( .A(RST), .B(bus_sync_state_machine_ECLK1), .Y(bus_sync_state_machine__0EECLK1_0_0_));
AND2X2 AND2X2_214 ( .A(RST), .B(bus_sync_status_reg_data2_0_), .Y(bus_sync_status__0reg_data3_2_0__0_));
AND2X2 AND2X2_215 ( .A(RST), .B(bus_sync_status_reg_data2_1_), .Y(bus_sync_status__0reg_data3_2_0__1_));
AND2X2 AND2X2_216 ( .A(RST), .B(bus_sync_status_reg_data2_2_), .Y(bus_sync_status__0reg_data3_2_0__2_));
AND2X2 AND2X2_217 ( .A(RST), .B(busy), .Y(bus_sync_status__0reg_data1_2_0__0_));
AND2X2 AND2X2_218 ( .A(RST), .B(axi_awvalid), .Y(bus_sync_status__0reg_data1_2_0__1_));
AND2X2 AND2X2_219 ( .A(RST), .B(axi_arvalid), .Y(bus_sync_status__0reg_data1_2_0__2_));
AND2X2 AND2X2_22 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_14_), .Y(bus_sync_axi_bus__0reg_data3_63_0__14_));
AND2X2 AND2X2_220 ( .A(RST), .B(bus_sync_status_ECLK2), .Y(bus_sync_status__0EECLK2_0_0_));
AND2X2 AND2X2_221 ( .A(RST), .B(SCLK), .Y(bus_sync_status__0ECLK2_0_0_));
AND2X2 AND2X2_23 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_15_), .Y(bus_sync_axi_bus__0reg_data3_63_0__15_));
AND2X2 AND2X2_24 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_16_), .Y(bus_sync_axi_bus__0reg_data3_63_0__16_));
AND2X2 AND2X2_25 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_17_), .Y(bus_sync_axi_bus__0reg_data3_63_0__17_));
AND2X2 AND2X2_26 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_18_), .Y(bus_sync_axi_bus__0reg_data3_63_0__18_));
AND2X2 AND2X2_27 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_19_), .Y(bus_sync_axi_bus__0reg_data3_63_0__19_));
AND2X2 AND2X2_28 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_20_), .Y(bus_sync_axi_bus__0reg_data3_63_0__20_));
AND2X2 AND2X2_29 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_21_), .Y(bus_sync_axi_bus__0reg_data3_63_0__21_));
AND2X2 AND2X2_3 ( .A(_abc_4169_new_n615_), .B(_abc_4169_new_n622_), .Y(_abc_4169_new_n649_));
AND2X2 AND2X2_30 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_22_), .Y(bus_sync_axi_bus__0reg_data3_63_0__22_));
AND2X2 AND2X2_31 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_23_), .Y(bus_sync_axi_bus__0reg_data3_63_0__23_));
AND2X2 AND2X2_32 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_24_), .Y(bus_sync_axi_bus__0reg_data3_63_0__24_));
AND2X2 AND2X2_33 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_25_), .Y(bus_sync_axi_bus__0reg_data3_63_0__25_));
AND2X2 AND2X2_34 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_26_), .Y(bus_sync_axi_bus__0reg_data3_63_0__26_));
AND2X2 AND2X2_35 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_27_), .Y(bus_sync_axi_bus__0reg_data3_63_0__27_));
AND2X2 AND2X2_36 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_28_), .Y(bus_sync_axi_bus__0reg_data3_63_0__28_));
AND2X2 AND2X2_37 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_29_), .Y(bus_sync_axi_bus__0reg_data3_63_0__29_));
AND2X2 AND2X2_38 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_30_), .Y(bus_sync_axi_bus__0reg_data3_63_0__30_));
AND2X2 AND2X2_39 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_31_), .Y(bus_sync_axi_bus__0reg_data3_63_0__31_));
AND2X2 AND2X2_4 ( .A(_abc_4169_new_n631_), .B(_abc_4169_new_n639_), .Y(_abc_4169_new_n650_));
AND2X2 AND2X2_40 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_32_), .Y(bus_sync_axi_bus__0reg_data3_63_0__32_));
AND2X2 AND2X2_41 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_33_), .Y(bus_sync_axi_bus__0reg_data3_63_0__33_));
AND2X2 AND2X2_42 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_34_), .Y(bus_sync_axi_bus__0reg_data3_63_0__34_));
AND2X2 AND2X2_43 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_35_), .Y(bus_sync_axi_bus__0reg_data3_63_0__35_));
AND2X2 AND2X2_44 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_36_), .Y(bus_sync_axi_bus__0reg_data3_63_0__36_));
AND2X2 AND2X2_45 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_37_), .Y(bus_sync_axi_bus__0reg_data3_63_0__37_));
AND2X2 AND2X2_46 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_38_), .Y(bus_sync_axi_bus__0reg_data3_63_0__38_));
AND2X2 AND2X2_47 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_39_), .Y(bus_sync_axi_bus__0reg_data3_63_0__39_));
AND2X2 AND2X2_48 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_40_), .Y(bus_sync_axi_bus__0reg_data3_63_0__40_));
AND2X2 AND2X2_49 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_41_), .Y(bus_sync_axi_bus__0reg_data3_63_0__41_));
AND2X2 AND2X2_5 ( .A(_abc_4169_new_n598_), .B(bus_sync_status_data_out_1_), .Y(_abc_4169_new_n653_));
AND2X2 AND2X2_50 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_42_), .Y(bus_sync_axi_bus__0reg_data3_63_0__42_));
AND2X2 AND2X2_51 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_43_), .Y(bus_sync_axi_bus__0reg_data3_63_0__43_));
AND2X2 AND2X2_52 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_44_), .Y(bus_sync_axi_bus__0reg_data3_63_0__44_));
AND2X2 AND2X2_53 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_45_), .Y(bus_sync_axi_bus__0reg_data3_63_0__45_));
AND2X2 AND2X2_54 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_46_), .Y(bus_sync_axi_bus__0reg_data3_63_0__46_));
AND2X2 AND2X2_55 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_47_), .Y(bus_sync_axi_bus__0reg_data3_63_0__47_));
AND2X2 AND2X2_56 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_48_), .Y(bus_sync_axi_bus__0reg_data3_63_0__48_));
AND2X2 AND2X2_57 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_49_), .Y(bus_sync_axi_bus__0reg_data3_63_0__49_));
AND2X2 AND2X2_58 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_50_), .Y(bus_sync_axi_bus__0reg_data3_63_0__50_));
AND2X2 AND2X2_59 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_51_), .Y(bus_sync_axi_bus__0reg_data3_63_0__51_));
AND2X2 AND2X2_6 ( .A(_abc_4169_new_n598_), .B(bus_sync_status_data_out_2_), .Y(_abc_4169_new_n660_));
AND2X2 AND2X2_60 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_52_), .Y(bus_sync_axi_bus__0reg_data3_63_0__52_));
AND2X2 AND2X2_61 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_53_), .Y(bus_sync_axi_bus__0reg_data3_63_0__53_));
AND2X2 AND2X2_62 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_54_), .Y(bus_sync_axi_bus__0reg_data3_63_0__54_));
AND2X2 AND2X2_63 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_55_), .Y(bus_sync_axi_bus__0reg_data3_63_0__55_));
AND2X2 AND2X2_64 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_56_), .Y(bus_sync_axi_bus__0reg_data3_63_0__56_));
AND2X2 AND2X2_65 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_57_), .Y(bus_sync_axi_bus__0reg_data3_63_0__57_));
AND2X2 AND2X2_66 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_58_), .Y(bus_sync_axi_bus__0reg_data3_63_0__58_));
AND2X2 AND2X2_67 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_59_), .Y(bus_sync_axi_bus__0reg_data3_63_0__59_));
AND2X2 AND2X2_68 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_60_), .Y(bus_sync_axi_bus__0reg_data3_63_0__60_));
AND2X2 AND2X2_69 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_61_), .Y(bus_sync_axi_bus__0reg_data3_63_0__61_));
AND2X2 AND2X2_7 ( .A(RST), .B(counter_65_), .Y(_0fini_spi_0_0_));
AND2X2 AND2X2_70 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_62_), .Y(bus_sync_axi_bus__0reg_data3_63_0__62_));
AND2X2 AND2X2_71 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_63_), .Y(bus_sync_axi_bus__0reg_data3_63_0__63_));
AND2X2 AND2X2_72 ( .A(RST), .B(WDATA_0_), .Y(bus_sync_axi_bus__0reg_data1_63_0__0_));
AND2X2 AND2X2_73 ( .A(RST), .B(WDATA_1_), .Y(bus_sync_axi_bus__0reg_data1_63_0__1_));
AND2X2 AND2X2_74 ( .A(RST), .B(WDATA_2_), .Y(bus_sync_axi_bus__0reg_data1_63_0__2_));
AND2X2 AND2X2_75 ( .A(RST), .B(WDATA_3_), .Y(bus_sync_axi_bus__0reg_data1_63_0__3_));
AND2X2 AND2X2_76 ( .A(RST), .B(WDATA_4_), .Y(bus_sync_axi_bus__0reg_data1_63_0__4_));
AND2X2 AND2X2_77 ( .A(RST), .B(WDATA_5_), .Y(bus_sync_axi_bus__0reg_data1_63_0__5_));
AND2X2 AND2X2_78 ( .A(RST), .B(WDATA_6_), .Y(bus_sync_axi_bus__0reg_data1_63_0__6_));
AND2X2 AND2X2_79 ( .A(RST), .B(WDATA_7_), .Y(bus_sync_axi_bus__0reg_data1_63_0__7_));
AND2X2 AND2X2_8 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_0_), .Y(bus_sync_axi_bus__0reg_data3_63_0__0_));
AND2X2 AND2X2_80 ( .A(RST), .B(WDATA_8_), .Y(bus_sync_axi_bus__0reg_data1_63_0__8_));
AND2X2 AND2X2_81 ( .A(RST), .B(WDATA_9_), .Y(bus_sync_axi_bus__0reg_data1_63_0__9_));
AND2X2 AND2X2_82 ( .A(RST), .B(WDATA_10_), .Y(bus_sync_axi_bus__0reg_data1_63_0__10_));
AND2X2 AND2X2_83 ( .A(RST), .B(WDATA_11_), .Y(bus_sync_axi_bus__0reg_data1_63_0__11_));
AND2X2 AND2X2_84 ( .A(RST), .B(WDATA_12_), .Y(bus_sync_axi_bus__0reg_data1_63_0__12_));
AND2X2 AND2X2_85 ( .A(RST), .B(WDATA_13_), .Y(bus_sync_axi_bus__0reg_data1_63_0__13_));
AND2X2 AND2X2_86 ( .A(RST), .B(WDATA_14_), .Y(bus_sync_axi_bus__0reg_data1_63_0__14_));
AND2X2 AND2X2_87 ( .A(RST), .B(WDATA_15_), .Y(bus_sync_axi_bus__0reg_data1_63_0__15_));
AND2X2 AND2X2_88 ( .A(RST), .B(WDATA_16_), .Y(bus_sync_axi_bus__0reg_data1_63_0__16_));
AND2X2 AND2X2_89 ( .A(RST), .B(WDATA_17_), .Y(bus_sync_axi_bus__0reg_data1_63_0__17_));
AND2X2 AND2X2_9 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_1_), .Y(bus_sync_axi_bus__0reg_data3_63_0__1_));
AND2X2 AND2X2_90 ( .A(RST), .B(WDATA_18_), .Y(bus_sync_axi_bus__0reg_data1_63_0__18_));
AND2X2 AND2X2_91 ( .A(RST), .B(WDATA_19_), .Y(bus_sync_axi_bus__0reg_data1_63_0__19_));
AND2X2 AND2X2_92 ( .A(RST), .B(WDATA_20_), .Y(bus_sync_axi_bus__0reg_data1_63_0__20_));
AND2X2 AND2X2_93 ( .A(RST), .B(WDATA_21_), .Y(bus_sync_axi_bus__0reg_data1_63_0__21_));
AND2X2 AND2X2_94 ( .A(RST), .B(WDATA_22_), .Y(bus_sync_axi_bus__0reg_data1_63_0__22_));
AND2X2 AND2X2_95 ( .A(RST), .B(WDATA_23_), .Y(bus_sync_axi_bus__0reg_data1_63_0__23_));
AND2X2 AND2X2_96 ( .A(RST), .B(WDATA_24_), .Y(bus_sync_axi_bus__0reg_data1_63_0__24_));
AND2X2 AND2X2_97 ( .A(RST), .B(WDATA_25_), .Y(bus_sync_axi_bus__0reg_data1_63_0__25_));
AND2X2 AND2X2_98 ( .A(RST), .B(WDATA_26_), .Y(bus_sync_axi_bus__0reg_data1_63_0__26_));
AND2X2 AND2X2_99 ( .A(RST), .B(WDATA_27_), .Y(bus_sync_axi_bus__0reg_data1_63_0__27_));
AOI21X1 AOI21X1_1 ( .A(_abc_4169_new_n568_), .B(_abc_4169_new_n569_), .C(_abc_4169_new_n564_), .Y(_abc_2903_auto_fsm_map_cc_170_map_fsm_402_1_));
AOI21X1 AOI21X1_10 ( .A(_abc_4169_new_n651_), .B(bus_cap_3_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n672_));
AOI21X1 AOI21X1_100 ( .A(_abc_4169_new_n944_), .B(_abc_4169_new_n938_), .C(_abc_4169_new_n945_), .Y(_0WDATA_31_0__2_));
AOI21X1 AOI21X1_101 ( .A(_abc_4169_new_n947_), .B(_abc_4169_new_n938_), .C(_abc_4169_new_n948_), .Y(_0WDATA_31_0__3_));
AOI21X1 AOI21X1_102 ( .A(_abc_4169_new_n950_), .B(_abc_4169_new_n938_), .C(_abc_4169_new_n951_), .Y(_0WDATA_31_0__4_));
AOI21X1 AOI21X1_103 ( .A(_abc_4169_new_n953_), .B(_abc_4169_new_n938_), .C(_abc_4169_new_n954_), .Y(_0WDATA_31_0__5_));
AOI21X1 AOI21X1_104 ( .A(_abc_4169_new_n956_), .B(_abc_4169_new_n938_), .C(_abc_4169_new_n957_), .Y(_0WDATA_31_0__6_));
AOI21X1 AOI21X1_105 ( .A(_abc_4169_new_n959_), .B(_abc_4169_new_n938_), .C(_abc_4169_new_n960_), .Y(_0WDATA_31_0__7_));
AOI21X1 AOI21X1_106 ( .A(_abc_4169_new_n962_), .B(_abc_4169_new_n938_), .C(_abc_4169_new_n963_), .Y(_0WDATA_31_0__8_));
AOI21X1 AOI21X1_107 ( .A(_abc_4169_new_n965_), .B(_abc_4169_new_n938_), .C(_abc_4169_new_n966_), .Y(_0WDATA_31_0__9_));
AOI21X1 AOI21X1_108 ( .A(_abc_4169_new_n968_), .B(_abc_4169_new_n938_), .C(_abc_4169_new_n969_), .Y(_0WDATA_31_0__10_));
AOI21X1 AOI21X1_109 ( .A(_abc_4169_new_n971_), .B(_abc_4169_new_n938_), .C(_abc_4169_new_n972_), .Y(_0WDATA_31_0__11_));
AOI21X1 AOI21X1_11 ( .A(_abc_4169_new_n672_), .B(_abc_4169_new_n671_), .C(_abc_4169_new_n675_), .Y(_0bus_cap_31_0__4_));
AOI21X1 AOI21X1_110 ( .A(_abc_4169_new_n974_), .B(_abc_4169_new_n938_), .C(_abc_4169_new_n975_), .Y(_0WDATA_31_0__12_));
AOI21X1 AOI21X1_111 ( .A(_abc_4169_new_n977_), .B(_abc_4169_new_n938_), .C(_abc_4169_new_n978_), .Y(_0WDATA_31_0__13_));
AOI21X1 AOI21X1_112 ( .A(_abc_4169_new_n980_), .B(_abc_4169_new_n938_), .C(_abc_4169_new_n981_), .Y(_0WDATA_31_0__14_));
AOI21X1 AOI21X1_113 ( .A(_abc_4169_new_n983_), .B(_abc_4169_new_n938_), .C(_abc_4169_new_n984_), .Y(_0WDATA_31_0__15_));
AOI21X1 AOI21X1_114 ( .A(_abc_4169_new_n986_), .B(_abc_4169_new_n938_), .C(_abc_4169_new_n987_), .Y(_0WDATA_31_0__16_));
AOI21X1 AOI21X1_115 ( .A(_abc_4169_new_n989_), .B(_abc_4169_new_n938_), .C(_abc_4169_new_n990_), .Y(_0WDATA_31_0__17_));
AOI21X1 AOI21X1_116 ( .A(_abc_4169_new_n992_), .B(_abc_4169_new_n938_), .C(_abc_4169_new_n993_), .Y(_0WDATA_31_0__18_));
AOI21X1 AOI21X1_117 ( .A(_abc_4169_new_n995_), .B(_abc_4169_new_n938_), .C(_abc_4169_new_n996_), .Y(_0WDATA_31_0__19_));
AOI21X1 AOI21X1_118 ( .A(_abc_4169_new_n998_), .B(_abc_4169_new_n938_), .C(_abc_4169_new_n999_), .Y(_0WDATA_31_0__20_));
AOI21X1 AOI21X1_119 ( .A(_abc_4169_new_n1001_), .B(_abc_4169_new_n938_), .C(_abc_4169_new_n1002_), .Y(_0WDATA_31_0__21_));
AOI21X1 AOI21X1_12 ( .A(_abc_4169_new_n651_), .B(bus_cap_4_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n678_));
AOI21X1 AOI21X1_120 ( .A(_abc_4169_new_n1004_), .B(_abc_4169_new_n938_), .C(_abc_4169_new_n1005_), .Y(_0WDATA_31_0__22_));
AOI21X1 AOI21X1_121 ( .A(_abc_4169_new_n1007_), .B(_abc_4169_new_n938_), .C(_abc_4169_new_n1008_), .Y(_0WDATA_31_0__23_));
AOI21X1 AOI21X1_122 ( .A(_abc_4169_new_n1010_), .B(_abc_4169_new_n938_), .C(_abc_4169_new_n1011_), .Y(_0WDATA_31_0__24_));
AOI21X1 AOI21X1_123 ( .A(_abc_4169_new_n1013_), .B(_abc_4169_new_n938_), .C(_abc_4169_new_n1014_), .Y(_0WDATA_31_0__25_));
AOI21X1 AOI21X1_124 ( .A(_abc_4169_new_n1016_), .B(_abc_4169_new_n938_), .C(_abc_4169_new_n1017_), .Y(_0WDATA_31_0__26_));
AOI21X1 AOI21X1_125 ( .A(_abc_4169_new_n1019_), .B(_abc_4169_new_n938_), .C(_abc_4169_new_n1020_), .Y(_0WDATA_31_0__27_));
AOI21X1 AOI21X1_126 ( .A(_abc_4169_new_n1022_), .B(_abc_4169_new_n938_), .C(_abc_4169_new_n1023_), .Y(_0WDATA_31_0__28_));
AOI21X1 AOI21X1_127 ( .A(_abc_4169_new_n1025_), .B(_abc_4169_new_n938_), .C(_abc_4169_new_n1026_), .Y(_0WDATA_31_0__29_));
AOI21X1 AOI21X1_128 ( .A(_abc_4169_new_n1028_), .B(_abc_4169_new_n938_), .C(_abc_4169_new_n1029_), .Y(_0WDATA_31_0__30_));
AOI21X1 AOI21X1_129 ( .A(_abc_4169_new_n1031_), .B(_abc_4169_new_n938_), .C(_abc_4169_new_n1032_), .Y(_0WDATA_31_0__31_));
AOI21X1 AOI21X1_13 ( .A(_abc_4169_new_n678_), .B(_abc_4169_new_n677_), .C(_abc_4169_new_n681_), .Y(_0bus_cap_31_0__5_));
AOI21X1 AOI21X1_130 ( .A(_abc_4169_new_n1034_), .B(_abc_4169_new_n1037_), .C(_abc_4169_new_n1038_), .Y(_0A_ADDR_31_0__0_));
AOI21X1 AOI21X1_131 ( .A(_abc_4169_new_n1040_), .B(_abc_4169_new_n1037_), .C(_abc_4169_new_n1041_), .Y(_0A_ADDR_31_0__1_));
AOI21X1 AOI21X1_132 ( .A(_abc_4169_new_n1043_), .B(_abc_4169_new_n1037_), .C(_abc_4169_new_n1044_), .Y(_0A_ADDR_31_0__2_));
AOI21X1 AOI21X1_133 ( .A(_abc_4169_new_n1046_), .B(_abc_4169_new_n1037_), .C(_abc_4169_new_n1047_), .Y(_0A_ADDR_31_0__3_));
AOI21X1 AOI21X1_134 ( .A(_abc_4169_new_n1049_), .B(_abc_4169_new_n1037_), .C(_abc_4169_new_n1050_), .Y(_0A_ADDR_31_0__4_));
AOI21X1 AOI21X1_135 ( .A(_abc_4169_new_n1052_), .B(_abc_4169_new_n1037_), .C(_abc_4169_new_n1053_), .Y(_0A_ADDR_31_0__5_));
AOI21X1 AOI21X1_136 ( .A(_abc_4169_new_n1055_), .B(_abc_4169_new_n1037_), .C(_abc_4169_new_n1056_), .Y(_0A_ADDR_31_0__6_));
AOI21X1 AOI21X1_137 ( .A(_abc_4169_new_n1058_), .B(_abc_4169_new_n1037_), .C(_abc_4169_new_n1059_), .Y(_0A_ADDR_31_0__7_));
AOI21X1 AOI21X1_138 ( .A(_abc_4169_new_n1061_), .B(_abc_4169_new_n1037_), .C(_abc_4169_new_n1062_), .Y(_0A_ADDR_31_0__8_));
AOI21X1 AOI21X1_139 ( .A(_abc_4169_new_n1064_), .B(_abc_4169_new_n1037_), .C(_abc_4169_new_n1065_), .Y(_0A_ADDR_31_0__9_));
AOI21X1 AOI21X1_14 ( .A(_abc_4169_new_n651_), .B(bus_cap_5_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n684_));
AOI21X1 AOI21X1_140 ( .A(_abc_4169_new_n1067_), .B(_abc_4169_new_n1037_), .C(_abc_4169_new_n1068_), .Y(_0A_ADDR_31_0__10_));
AOI21X1 AOI21X1_141 ( .A(_abc_4169_new_n1070_), .B(_abc_4169_new_n1037_), .C(_abc_4169_new_n1071_), .Y(_0A_ADDR_31_0__11_));
AOI21X1 AOI21X1_142 ( .A(_abc_4169_new_n1073_), .B(_abc_4169_new_n1037_), .C(_abc_4169_new_n1074_), .Y(_0A_ADDR_31_0__12_));
AOI21X1 AOI21X1_143 ( .A(_abc_4169_new_n1076_), .B(_abc_4169_new_n1037_), .C(_abc_4169_new_n1077_), .Y(_0A_ADDR_31_0__13_));
AOI21X1 AOI21X1_144 ( .A(_abc_4169_new_n1079_), .B(_abc_4169_new_n1037_), .C(_abc_4169_new_n1080_), .Y(_0A_ADDR_31_0__14_));
AOI21X1 AOI21X1_145 ( .A(_abc_4169_new_n1082_), .B(_abc_4169_new_n1037_), .C(_abc_4169_new_n1083_), .Y(_0A_ADDR_31_0__15_));
AOI21X1 AOI21X1_146 ( .A(_abc_4169_new_n1085_), .B(_abc_4169_new_n1037_), .C(_abc_4169_new_n1086_), .Y(_0A_ADDR_31_0__16_));
AOI21X1 AOI21X1_147 ( .A(_abc_4169_new_n1088_), .B(_abc_4169_new_n1037_), .C(_abc_4169_new_n1089_), .Y(_0A_ADDR_31_0__17_));
AOI21X1 AOI21X1_148 ( .A(_abc_4169_new_n1091_), .B(_abc_4169_new_n1037_), .C(_abc_4169_new_n1092_), .Y(_0A_ADDR_31_0__18_));
AOI21X1 AOI21X1_149 ( .A(_abc_4169_new_n1094_), .B(_abc_4169_new_n1037_), .C(_abc_4169_new_n1095_), .Y(_0A_ADDR_31_0__19_));
AOI21X1 AOI21X1_15 ( .A(_abc_4169_new_n684_), .B(_abc_4169_new_n683_), .C(_abc_4169_new_n687_), .Y(_0bus_cap_31_0__6_));
AOI21X1 AOI21X1_150 ( .A(_abc_4169_new_n1097_), .B(_abc_4169_new_n1037_), .C(_abc_4169_new_n1098_), .Y(_0A_ADDR_31_0__20_));
AOI21X1 AOI21X1_151 ( .A(_abc_4169_new_n1100_), .B(_abc_4169_new_n1037_), .C(_abc_4169_new_n1101_), .Y(_0A_ADDR_31_0__21_));
AOI21X1 AOI21X1_152 ( .A(_abc_4169_new_n1103_), .B(_abc_4169_new_n1037_), .C(_abc_4169_new_n1104_), .Y(_0A_ADDR_31_0__22_));
AOI21X1 AOI21X1_153 ( .A(_abc_4169_new_n1106_), .B(_abc_4169_new_n1037_), .C(_abc_4169_new_n1107_), .Y(_0A_ADDR_31_0__23_));
AOI21X1 AOI21X1_154 ( .A(_abc_4169_new_n1109_), .B(_abc_4169_new_n1037_), .C(_abc_4169_new_n1110_), .Y(_0A_ADDR_31_0__24_));
AOI21X1 AOI21X1_155 ( .A(_abc_4169_new_n1112_), .B(_abc_4169_new_n1037_), .C(_abc_4169_new_n1113_), .Y(_0A_ADDR_31_0__25_));
AOI21X1 AOI21X1_156 ( .A(_abc_4169_new_n1115_), .B(_abc_4169_new_n1037_), .C(_abc_4169_new_n1116_), .Y(_0A_ADDR_31_0__26_));
AOI21X1 AOI21X1_157 ( .A(_abc_4169_new_n1118_), .B(_abc_4169_new_n1037_), .C(_abc_4169_new_n1119_), .Y(_0A_ADDR_31_0__27_));
AOI21X1 AOI21X1_158 ( .A(_abc_4169_new_n1121_), .B(_abc_4169_new_n1037_), .C(_abc_4169_new_n1122_), .Y(_0A_ADDR_31_0__28_));
AOI21X1 AOI21X1_159 ( .A(_abc_4169_new_n1124_), .B(_abc_4169_new_n1037_), .C(_abc_4169_new_n1125_), .Y(_0A_ADDR_31_0__29_));
AOI21X1 AOI21X1_16 ( .A(_abc_4169_new_n651_), .B(bus_cap_6_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n690_));
AOI21X1 AOI21X1_160 ( .A(_abc_4169_new_n1127_), .B(_abc_4169_new_n1037_), .C(_abc_4169_new_n1128_), .Y(_0A_ADDR_31_0__30_));
AOI21X1 AOI21X1_161 ( .A(_abc_4169_new_n1130_), .B(_abc_4169_new_n1037_), .C(_abc_4169_new_n1131_), .Y(_0A_ADDR_31_0__31_));
AOI21X1 AOI21X1_162 ( .A(CEB), .B(_abc_4169_new_n1133_), .C(_abc_4169_new_n1134_), .Y(_0sft_reg_65_0__0_));
AOI21X1 AOI21X1_163 ( .A(_abc_4169_new_n937_), .B(_abc_4169_new_n1133_), .C(_abc_4169_new_n1136_), .Y(_0sft_reg_65_0__1_));
AOI21X1 AOI21X1_164 ( .A(CEB), .B(_abc_4169_new_n1138_), .C(_abc_4169_new_n1139_), .Y(_0sft_reg_65_0__2_));
AOI21X1 AOI21X1_165 ( .A(_abc_4169_new_n937_), .B(_abc_4169_new_n1138_), .C(_abc_4169_new_n1141_), .Y(_0sft_reg_65_0__3_));
AOI21X1 AOI21X1_166 ( .A(CEB), .B(_abc_4169_new_n1143_), .C(_abc_4169_new_n1144_), .Y(_0sft_reg_65_0__4_));
AOI21X1 AOI21X1_167 ( .A(_abc_4169_new_n937_), .B(_abc_4169_new_n1143_), .C(_abc_4169_new_n1146_), .Y(_0sft_reg_65_0__5_));
AOI21X1 AOI21X1_168 ( .A(CEB), .B(_abc_4169_new_n1148_), .C(_abc_4169_new_n1149_), .Y(_0sft_reg_65_0__6_));
AOI21X1 AOI21X1_169 ( .A(_abc_4169_new_n937_), .B(_abc_4169_new_n1148_), .C(_abc_4169_new_n1151_), .Y(_0sft_reg_65_0__7_));
AOI21X1 AOI21X1_17 ( .A(_abc_4169_new_n690_), .B(_abc_4169_new_n689_), .C(_abc_4169_new_n693_), .Y(_0bus_cap_31_0__7_));
AOI21X1 AOI21X1_170 ( .A(CEB), .B(_abc_4169_new_n1153_), .C(_abc_4169_new_n1154_), .Y(_0sft_reg_65_0__8_));
AOI21X1 AOI21X1_171 ( .A(_abc_4169_new_n937_), .B(_abc_4169_new_n1153_), .C(_abc_4169_new_n1156_), .Y(_0sft_reg_65_0__9_));
AOI21X1 AOI21X1_172 ( .A(CEB), .B(_abc_4169_new_n1158_), .C(_abc_4169_new_n1159_), .Y(_0sft_reg_65_0__10_));
AOI21X1 AOI21X1_173 ( .A(_abc_4169_new_n937_), .B(_abc_4169_new_n1158_), .C(_abc_4169_new_n1161_), .Y(_0sft_reg_65_0__11_));
AOI21X1 AOI21X1_174 ( .A(CEB), .B(_abc_4169_new_n1163_), .C(_abc_4169_new_n1164_), .Y(_0sft_reg_65_0__12_));
AOI21X1 AOI21X1_175 ( .A(_abc_4169_new_n937_), .B(_abc_4169_new_n1163_), .C(_abc_4169_new_n1166_), .Y(_0sft_reg_65_0__13_));
AOI21X1 AOI21X1_176 ( .A(CEB), .B(_abc_4169_new_n1168_), .C(_abc_4169_new_n1169_), .Y(_0sft_reg_65_0__14_));
AOI21X1 AOI21X1_177 ( .A(_abc_4169_new_n937_), .B(_abc_4169_new_n1168_), .C(_abc_4169_new_n1171_), .Y(_0sft_reg_65_0__15_));
AOI21X1 AOI21X1_178 ( .A(CEB), .B(_abc_4169_new_n1173_), .C(_abc_4169_new_n1174_), .Y(_0sft_reg_65_0__16_));
AOI21X1 AOI21X1_179 ( .A(_abc_4169_new_n937_), .B(_abc_4169_new_n1173_), .C(_abc_4169_new_n1176_), .Y(_0sft_reg_65_0__17_));
AOI21X1 AOI21X1_18 ( .A(_abc_4169_new_n651_), .B(bus_cap_7_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n696_));
AOI21X1 AOI21X1_180 ( .A(CEB), .B(_abc_4169_new_n1178_), .C(_abc_4169_new_n1179_), .Y(_0sft_reg_65_0__18_));
AOI21X1 AOI21X1_181 ( .A(_abc_4169_new_n937_), .B(_abc_4169_new_n1178_), .C(_abc_4169_new_n1181_), .Y(_0sft_reg_65_0__19_));
AOI21X1 AOI21X1_182 ( .A(CEB), .B(_abc_4169_new_n1183_), .C(_abc_4169_new_n1184_), .Y(_0sft_reg_65_0__20_));
AOI21X1 AOI21X1_183 ( .A(_abc_4169_new_n937_), .B(_abc_4169_new_n1183_), .C(_abc_4169_new_n1186_), .Y(_0sft_reg_65_0__21_));
AOI21X1 AOI21X1_184 ( .A(CEB), .B(_abc_4169_new_n1188_), .C(_abc_4169_new_n1189_), .Y(_0sft_reg_65_0__22_));
AOI21X1 AOI21X1_185 ( .A(_abc_4169_new_n937_), .B(_abc_4169_new_n1188_), .C(_abc_4169_new_n1191_), .Y(_0sft_reg_65_0__23_));
AOI21X1 AOI21X1_186 ( .A(CEB), .B(_abc_4169_new_n1193_), .C(_abc_4169_new_n1194_), .Y(_0sft_reg_65_0__24_));
AOI21X1 AOI21X1_187 ( .A(_abc_4169_new_n937_), .B(_abc_4169_new_n1193_), .C(_abc_4169_new_n1196_), .Y(_0sft_reg_65_0__25_));
AOI21X1 AOI21X1_188 ( .A(CEB), .B(_abc_4169_new_n1198_), .C(_abc_4169_new_n1199_), .Y(_0sft_reg_65_0__26_));
AOI21X1 AOI21X1_189 ( .A(_abc_4169_new_n937_), .B(_abc_4169_new_n1198_), .C(_abc_4169_new_n1201_), .Y(_0sft_reg_65_0__27_));
AOI21X1 AOI21X1_19 ( .A(_abc_4169_new_n696_), .B(_abc_4169_new_n695_), .C(_abc_4169_new_n699_), .Y(_0bus_cap_31_0__8_));
AOI21X1 AOI21X1_190 ( .A(CEB), .B(_abc_4169_new_n1203_), .C(_abc_4169_new_n1204_), .Y(_0sft_reg_65_0__28_));
AOI21X1 AOI21X1_191 ( .A(_abc_4169_new_n937_), .B(_abc_4169_new_n1203_), .C(_abc_4169_new_n1206_), .Y(_0sft_reg_65_0__29_));
AOI21X1 AOI21X1_192 ( .A(CEB), .B(_abc_4169_new_n1208_), .C(_abc_4169_new_n1209_), .Y(_0sft_reg_65_0__30_));
AOI21X1 AOI21X1_193 ( .A(_abc_4169_new_n1334_), .B(_abc_4169_new_n1336_), .C(_abc_4169_new_n1337_), .Y(_0PICORV_RST_SPI_0_0_));
AOI21X1 AOI21X1_194 ( .A(_abc_4169_new_n604_), .B(_abc_4169_new_n1339_), .C(_abc_4169_new_n1341_), .Y(_0re_0_0_));
AOI21X1 AOI21X1_195 ( .A(_abc_4169_new_n605_), .B(_abc_4169_new_n1343_), .C(_abc_4169_new_n1344_), .Y(_0we_0_0_));
AOI21X1 AOI21X1_196 ( .A(bus_sync_axi_bus__abc_3843_new_n395_), .B(bus_sync_axi_bus__abc_3843_new_n396_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__0_));
AOI21X1 AOI21X1_197 ( .A(bus_sync_axi_bus__abc_3843_new_n398_), .B(bus_sync_axi_bus__abc_3843_new_n399_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__1_));
AOI21X1 AOI21X1_198 ( .A(bus_sync_axi_bus__abc_3843_new_n401_), .B(bus_sync_axi_bus__abc_3843_new_n402_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__2_));
AOI21X1 AOI21X1_199 ( .A(bus_sync_axi_bus__abc_3843_new_n404_), .B(bus_sync_axi_bus__abc_3843_new_n405_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__3_));
AOI21X1 AOI21X1_2 ( .A(_abc_4169_new_n590_), .B(state_1_), .C(_abc_4169_new_n564_), .Y(_abc_4169_new_n591_));
AOI21X1 AOI21X1_20 ( .A(_abc_4169_new_n651_), .B(bus_cap_8_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n702_));
AOI21X1 AOI21X1_200 ( .A(bus_sync_axi_bus__abc_3843_new_n407_), .B(bus_sync_axi_bus__abc_3843_new_n408_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__4_));
AOI21X1 AOI21X1_201 ( .A(bus_sync_axi_bus__abc_3843_new_n410_), .B(bus_sync_axi_bus__abc_3843_new_n411_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__5_));
AOI21X1 AOI21X1_202 ( .A(bus_sync_axi_bus__abc_3843_new_n413_), .B(bus_sync_axi_bus__abc_3843_new_n414_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__6_));
AOI21X1 AOI21X1_203 ( .A(bus_sync_axi_bus__abc_3843_new_n416_), .B(bus_sync_axi_bus__abc_3843_new_n417_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__7_));
AOI21X1 AOI21X1_204 ( .A(bus_sync_axi_bus__abc_3843_new_n419_), .B(bus_sync_axi_bus__abc_3843_new_n420_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__8_));
AOI21X1 AOI21X1_205 ( .A(bus_sync_axi_bus__abc_3843_new_n422_), .B(bus_sync_axi_bus__abc_3843_new_n423_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__9_));
AOI21X1 AOI21X1_206 ( .A(bus_sync_axi_bus__abc_3843_new_n425_), .B(bus_sync_axi_bus__abc_3843_new_n426_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__10_));
AOI21X1 AOI21X1_207 ( .A(bus_sync_axi_bus__abc_3843_new_n428_), .B(bus_sync_axi_bus__abc_3843_new_n429_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__11_));
AOI21X1 AOI21X1_208 ( .A(bus_sync_axi_bus__abc_3843_new_n431_), .B(bus_sync_axi_bus__abc_3843_new_n432_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__12_));
AOI21X1 AOI21X1_209 ( .A(bus_sync_axi_bus__abc_3843_new_n434_), .B(bus_sync_axi_bus__abc_3843_new_n435_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__13_));
AOI21X1 AOI21X1_21 ( .A(_abc_4169_new_n702_), .B(_abc_4169_new_n701_), .C(_abc_4169_new_n705_), .Y(_0bus_cap_31_0__9_));
AOI21X1 AOI21X1_210 ( .A(bus_sync_axi_bus__abc_3843_new_n437_), .B(bus_sync_axi_bus__abc_3843_new_n438_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__14_));
AOI21X1 AOI21X1_211 ( .A(bus_sync_axi_bus__abc_3843_new_n440_), .B(bus_sync_axi_bus__abc_3843_new_n441_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__15_));
AOI21X1 AOI21X1_212 ( .A(bus_sync_axi_bus__abc_3843_new_n443_), .B(bus_sync_axi_bus__abc_3843_new_n444_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__16_));
AOI21X1 AOI21X1_213 ( .A(bus_sync_axi_bus__abc_3843_new_n446_), .B(bus_sync_axi_bus__abc_3843_new_n447_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__17_));
AOI21X1 AOI21X1_214 ( .A(bus_sync_axi_bus__abc_3843_new_n449_), .B(bus_sync_axi_bus__abc_3843_new_n450_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__18_));
AOI21X1 AOI21X1_215 ( .A(bus_sync_axi_bus__abc_3843_new_n452_), .B(bus_sync_axi_bus__abc_3843_new_n453_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__19_));
AOI21X1 AOI21X1_216 ( .A(bus_sync_axi_bus__abc_3843_new_n455_), .B(bus_sync_axi_bus__abc_3843_new_n456_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__20_));
AOI21X1 AOI21X1_217 ( .A(bus_sync_axi_bus__abc_3843_new_n458_), .B(bus_sync_axi_bus__abc_3843_new_n459_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__21_));
AOI21X1 AOI21X1_218 ( .A(bus_sync_axi_bus__abc_3843_new_n461_), .B(bus_sync_axi_bus__abc_3843_new_n462_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__22_));
AOI21X1 AOI21X1_219 ( .A(bus_sync_axi_bus__abc_3843_new_n464_), .B(bus_sync_axi_bus__abc_3843_new_n465_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__23_));
AOI21X1 AOI21X1_22 ( .A(_abc_4169_new_n651_), .B(bus_cap_9_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n708_));
AOI21X1 AOI21X1_220 ( .A(bus_sync_axi_bus__abc_3843_new_n467_), .B(bus_sync_axi_bus__abc_3843_new_n468_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__24_));
AOI21X1 AOI21X1_221 ( .A(bus_sync_axi_bus__abc_3843_new_n470_), .B(bus_sync_axi_bus__abc_3843_new_n471_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__25_));
AOI21X1 AOI21X1_222 ( .A(bus_sync_axi_bus__abc_3843_new_n473_), .B(bus_sync_axi_bus__abc_3843_new_n474_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__26_));
AOI21X1 AOI21X1_223 ( .A(bus_sync_axi_bus__abc_3843_new_n476_), .B(bus_sync_axi_bus__abc_3843_new_n477_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__27_));
AOI21X1 AOI21X1_224 ( .A(bus_sync_axi_bus__abc_3843_new_n479_), .B(bus_sync_axi_bus__abc_3843_new_n480_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__28_));
AOI21X1 AOI21X1_225 ( .A(bus_sync_axi_bus__abc_3843_new_n482_), .B(bus_sync_axi_bus__abc_3843_new_n483_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__29_));
AOI21X1 AOI21X1_226 ( .A(bus_sync_axi_bus__abc_3843_new_n485_), .B(bus_sync_axi_bus__abc_3843_new_n486_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__30_));
AOI21X1 AOI21X1_227 ( .A(bus_sync_axi_bus__abc_3843_new_n488_), .B(bus_sync_axi_bus__abc_3843_new_n489_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__31_));
AOI21X1 AOI21X1_228 ( .A(bus_sync_axi_bus__abc_3843_new_n491_), .B(bus_sync_axi_bus__abc_3843_new_n492_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__32_));
AOI21X1 AOI21X1_229 ( .A(bus_sync_axi_bus__abc_3843_new_n494_), .B(bus_sync_axi_bus__abc_3843_new_n495_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__33_));
AOI21X1 AOI21X1_23 ( .A(_abc_4169_new_n708_), .B(_abc_4169_new_n707_), .C(_abc_4169_new_n711_), .Y(_0bus_cap_31_0__10_));
AOI21X1 AOI21X1_230 ( .A(bus_sync_axi_bus__abc_3843_new_n497_), .B(bus_sync_axi_bus__abc_3843_new_n498_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__34_));
AOI21X1 AOI21X1_231 ( .A(bus_sync_axi_bus__abc_3843_new_n500_), .B(bus_sync_axi_bus__abc_3843_new_n501_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__35_));
AOI21X1 AOI21X1_232 ( .A(bus_sync_axi_bus__abc_3843_new_n503_), .B(bus_sync_axi_bus__abc_3843_new_n504_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__36_));
AOI21X1 AOI21X1_233 ( .A(bus_sync_axi_bus__abc_3843_new_n506_), .B(bus_sync_axi_bus__abc_3843_new_n507_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__37_));
AOI21X1 AOI21X1_234 ( .A(bus_sync_axi_bus__abc_3843_new_n509_), .B(bus_sync_axi_bus__abc_3843_new_n510_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__38_));
AOI21X1 AOI21X1_235 ( .A(bus_sync_axi_bus__abc_3843_new_n512_), .B(bus_sync_axi_bus__abc_3843_new_n513_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__39_));
AOI21X1 AOI21X1_236 ( .A(bus_sync_axi_bus__abc_3843_new_n515_), .B(bus_sync_axi_bus__abc_3843_new_n516_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__40_));
AOI21X1 AOI21X1_237 ( .A(bus_sync_axi_bus__abc_3843_new_n518_), .B(bus_sync_axi_bus__abc_3843_new_n519_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__41_));
AOI21X1 AOI21X1_238 ( .A(bus_sync_axi_bus__abc_3843_new_n521_), .B(bus_sync_axi_bus__abc_3843_new_n522_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__42_));
AOI21X1 AOI21X1_239 ( .A(bus_sync_axi_bus__abc_3843_new_n524_), .B(bus_sync_axi_bus__abc_3843_new_n525_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__43_));
AOI21X1 AOI21X1_24 ( .A(_abc_4169_new_n651_), .B(bus_cap_10_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n714_));
AOI21X1 AOI21X1_240 ( .A(bus_sync_axi_bus__abc_3843_new_n527_), .B(bus_sync_axi_bus__abc_3843_new_n528_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__44_));
AOI21X1 AOI21X1_241 ( .A(bus_sync_axi_bus__abc_3843_new_n530_), .B(bus_sync_axi_bus__abc_3843_new_n531_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__45_));
AOI21X1 AOI21X1_242 ( .A(bus_sync_axi_bus__abc_3843_new_n533_), .B(bus_sync_axi_bus__abc_3843_new_n534_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__46_));
AOI21X1 AOI21X1_243 ( .A(bus_sync_axi_bus__abc_3843_new_n536_), .B(bus_sync_axi_bus__abc_3843_new_n537_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__47_));
AOI21X1 AOI21X1_244 ( .A(bus_sync_axi_bus__abc_3843_new_n539_), .B(bus_sync_axi_bus__abc_3843_new_n540_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__48_));
AOI21X1 AOI21X1_245 ( .A(bus_sync_axi_bus__abc_3843_new_n542_), .B(bus_sync_axi_bus__abc_3843_new_n543_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__49_));
AOI21X1 AOI21X1_246 ( .A(bus_sync_axi_bus__abc_3843_new_n545_), .B(bus_sync_axi_bus__abc_3843_new_n546_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__50_));
AOI21X1 AOI21X1_247 ( .A(bus_sync_axi_bus__abc_3843_new_n548_), .B(bus_sync_axi_bus__abc_3843_new_n549_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__51_));
AOI21X1 AOI21X1_248 ( .A(bus_sync_axi_bus__abc_3843_new_n551_), .B(bus_sync_axi_bus__abc_3843_new_n552_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__52_));
AOI21X1 AOI21X1_249 ( .A(bus_sync_axi_bus__abc_3843_new_n554_), .B(bus_sync_axi_bus__abc_3843_new_n555_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__53_));
AOI21X1 AOI21X1_25 ( .A(_abc_4169_new_n714_), .B(_abc_4169_new_n713_), .C(_abc_4169_new_n717_), .Y(_0bus_cap_31_0__11_));
AOI21X1 AOI21X1_250 ( .A(bus_sync_axi_bus__abc_3843_new_n557_), .B(bus_sync_axi_bus__abc_3843_new_n558_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__54_));
AOI21X1 AOI21X1_251 ( .A(bus_sync_axi_bus__abc_3843_new_n560_), .B(bus_sync_axi_bus__abc_3843_new_n561_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__55_));
AOI21X1 AOI21X1_252 ( .A(bus_sync_axi_bus__abc_3843_new_n563_), .B(bus_sync_axi_bus__abc_3843_new_n564_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__56_));
AOI21X1 AOI21X1_253 ( .A(bus_sync_axi_bus__abc_3843_new_n566_), .B(bus_sync_axi_bus__abc_3843_new_n567_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__57_));
AOI21X1 AOI21X1_254 ( .A(bus_sync_axi_bus__abc_3843_new_n569_), .B(bus_sync_axi_bus__abc_3843_new_n570_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__58_));
AOI21X1 AOI21X1_255 ( .A(bus_sync_axi_bus__abc_3843_new_n572_), .B(bus_sync_axi_bus__abc_3843_new_n573_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__59_));
AOI21X1 AOI21X1_256 ( .A(bus_sync_axi_bus__abc_3843_new_n575_), .B(bus_sync_axi_bus__abc_3843_new_n576_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__60_));
AOI21X1 AOI21X1_257 ( .A(bus_sync_axi_bus__abc_3843_new_n578_), .B(bus_sync_axi_bus__abc_3843_new_n579_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__61_));
AOI21X1 AOI21X1_258 ( .A(bus_sync_axi_bus__abc_3843_new_n581_), .B(bus_sync_axi_bus__abc_3843_new_n582_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__62_));
AOI21X1 AOI21X1_259 ( .A(bus_sync_axi_bus__abc_3843_new_n584_), .B(bus_sync_axi_bus__abc_3843_new_n585_), .C(bus_sync_axi_bus__abc_3843_new_n393_), .Y(bus_sync_axi_bus__0reg_data2_63_0__63_));
AOI21X1 AOI21X1_26 ( .A(_abc_4169_new_n651_), .B(bus_cap_11_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n720_));
AOI21X1 AOI21X1_260 ( .A(bus_sync_rdata__abc_3651_new_n267_), .B(bus_sync_rdata__abc_3651_new_n268_), .C(bus_sync_rdata__abc_3651_new_n265_), .Y(bus_sync_rdata__0reg_data2_31_0__0_));
AOI21X1 AOI21X1_261 ( .A(bus_sync_rdata__abc_3651_new_n270_), .B(bus_sync_rdata__abc_3651_new_n271_), .C(bus_sync_rdata__abc_3651_new_n265_), .Y(bus_sync_rdata__0reg_data2_31_0__1_));
AOI21X1 AOI21X1_262 ( .A(bus_sync_rdata__abc_3651_new_n273_), .B(bus_sync_rdata__abc_3651_new_n274_), .C(bus_sync_rdata__abc_3651_new_n265_), .Y(bus_sync_rdata__0reg_data2_31_0__2_));
AOI21X1 AOI21X1_263 ( .A(bus_sync_rdata__abc_3651_new_n276_), .B(bus_sync_rdata__abc_3651_new_n277_), .C(bus_sync_rdata__abc_3651_new_n265_), .Y(bus_sync_rdata__0reg_data2_31_0__3_));
AOI21X1 AOI21X1_264 ( .A(bus_sync_rdata__abc_3651_new_n279_), .B(bus_sync_rdata__abc_3651_new_n280_), .C(bus_sync_rdata__abc_3651_new_n265_), .Y(bus_sync_rdata__0reg_data2_31_0__4_));
AOI21X1 AOI21X1_265 ( .A(bus_sync_rdata__abc_3651_new_n282_), .B(bus_sync_rdata__abc_3651_new_n283_), .C(bus_sync_rdata__abc_3651_new_n265_), .Y(bus_sync_rdata__0reg_data2_31_0__5_));
AOI21X1 AOI21X1_266 ( .A(bus_sync_rdata__abc_3651_new_n285_), .B(bus_sync_rdata__abc_3651_new_n286_), .C(bus_sync_rdata__abc_3651_new_n265_), .Y(bus_sync_rdata__0reg_data2_31_0__6_));
AOI21X1 AOI21X1_267 ( .A(bus_sync_rdata__abc_3651_new_n288_), .B(bus_sync_rdata__abc_3651_new_n289_), .C(bus_sync_rdata__abc_3651_new_n265_), .Y(bus_sync_rdata__0reg_data2_31_0__7_));
AOI21X1 AOI21X1_268 ( .A(bus_sync_rdata__abc_3651_new_n291_), .B(bus_sync_rdata__abc_3651_new_n292_), .C(bus_sync_rdata__abc_3651_new_n265_), .Y(bus_sync_rdata__0reg_data2_31_0__8_));
AOI21X1 AOI21X1_269 ( .A(bus_sync_rdata__abc_3651_new_n294_), .B(bus_sync_rdata__abc_3651_new_n295_), .C(bus_sync_rdata__abc_3651_new_n265_), .Y(bus_sync_rdata__0reg_data2_31_0__9_));
AOI21X1 AOI21X1_27 ( .A(_abc_4169_new_n720_), .B(_abc_4169_new_n719_), .C(_abc_4169_new_n723_), .Y(_0bus_cap_31_0__12_));
AOI21X1 AOI21X1_270 ( .A(bus_sync_rdata__abc_3651_new_n297_), .B(bus_sync_rdata__abc_3651_new_n298_), .C(bus_sync_rdata__abc_3651_new_n265_), .Y(bus_sync_rdata__0reg_data2_31_0__10_));
AOI21X1 AOI21X1_271 ( .A(bus_sync_rdata__abc_3651_new_n300_), .B(bus_sync_rdata__abc_3651_new_n301_), .C(bus_sync_rdata__abc_3651_new_n265_), .Y(bus_sync_rdata__0reg_data2_31_0__11_));
AOI21X1 AOI21X1_272 ( .A(bus_sync_rdata__abc_3651_new_n303_), .B(bus_sync_rdata__abc_3651_new_n304_), .C(bus_sync_rdata__abc_3651_new_n265_), .Y(bus_sync_rdata__0reg_data2_31_0__12_));
AOI21X1 AOI21X1_273 ( .A(bus_sync_rdata__abc_3651_new_n306_), .B(bus_sync_rdata__abc_3651_new_n307_), .C(bus_sync_rdata__abc_3651_new_n265_), .Y(bus_sync_rdata__0reg_data2_31_0__13_));
AOI21X1 AOI21X1_274 ( .A(bus_sync_rdata__abc_3651_new_n309_), .B(bus_sync_rdata__abc_3651_new_n310_), .C(bus_sync_rdata__abc_3651_new_n265_), .Y(bus_sync_rdata__0reg_data2_31_0__14_));
AOI21X1 AOI21X1_275 ( .A(bus_sync_rdata__abc_3651_new_n312_), .B(bus_sync_rdata__abc_3651_new_n313_), .C(bus_sync_rdata__abc_3651_new_n265_), .Y(bus_sync_rdata__0reg_data2_31_0__15_));
AOI21X1 AOI21X1_276 ( .A(bus_sync_rdata__abc_3651_new_n315_), .B(bus_sync_rdata__abc_3651_new_n316_), .C(bus_sync_rdata__abc_3651_new_n265_), .Y(bus_sync_rdata__0reg_data2_31_0__16_));
AOI21X1 AOI21X1_277 ( .A(bus_sync_rdata__abc_3651_new_n318_), .B(bus_sync_rdata__abc_3651_new_n319_), .C(bus_sync_rdata__abc_3651_new_n265_), .Y(bus_sync_rdata__0reg_data2_31_0__17_));
AOI21X1 AOI21X1_278 ( .A(bus_sync_rdata__abc_3651_new_n321_), .B(bus_sync_rdata__abc_3651_new_n322_), .C(bus_sync_rdata__abc_3651_new_n265_), .Y(bus_sync_rdata__0reg_data2_31_0__18_));
AOI21X1 AOI21X1_279 ( .A(bus_sync_rdata__abc_3651_new_n324_), .B(bus_sync_rdata__abc_3651_new_n325_), .C(bus_sync_rdata__abc_3651_new_n265_), .Y(bus_sync_rdata__0reg_data2_31_0__19_));
AOI21X1 AOI21X1_28 ( .A(_abc_4169_new_n651_), .B(bus_cap_12_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n726_));
AOI21X1 AOI21X1_280 ( .A(bus_sync_rdata__abc_3651_new_n327_), .B(bus_sync_rdata__abc_3651_new_n328_), .C(bus_sync_rdata__abc_3651_new_n265_), .Y(bus_sync_rdata__0reg_data2_31_0__20_));
AOI21X1 AOI21X1_281 ( .A(bus_sync_rdata__abc_3651_new_n330_), .B(bus_sync_rdata__abc_3651_new_n331_), .C(bus_sync_rdata__abc_3651_new_n265_), .Y(bus_sync_rdata__0reg_data2_31_0__21_));
AOI21X1 AOI21X1_282 ( .A(bus_sync_rdata__abc_3651_new_n333_), .B(bus_sync_rdata__abc_3651_new_n334_), .C(bus_sync_rdata__abc_3651_new_n265_), .Y(bus_sync_rdata__0reg_data2_31_0__22_));
AOI21X1 AOI21X1_283 ( .A(bus_sync_rdata__abc_3651_new_n336_), .B(bus_sync_rdata__abc_3651_new_n337_), .C(bus_sync_rdata__abc_3651_new_n265_), .Y(bus_sync_rdata__0reg_data2_31_0__23_));
AOI21X1 AOI21X1_284 ( .A(bus_sync_rdata__abc_3651_new_n339_), .B(bus_sync_rdata__abc_3651_new_n340_), .C(bus_sync_rdata__abc_3651_new_n265_), .Y(bus_sync_rdata__0reg_data2_31_0__24_));
AOI21X1 AOI21X1_285 ( .A(bus_sync_rdata__abc_3651_new_n342_), .B(bus_sync_rdata__abc_3651_new_n343_), .C(bus_sync_rdata__abc_3651_new_n265_), .Y(bus_sync_rdata__0reg_data2_31_0__25_));
AOI21X1 AOI21X1_286 ( .A(bus_sync_rdata__abc_3651_new_n345_), .B(bus_sync_rdata__abc_3651_new_n346_), .C(bus_sync_rdata__abc_3651_new_n265_), .Y(bus_sync_rdata__0reg_data2_31_0__26_));
AOI21X1 AOI21X1_287 ( .A(bus_sync_rdata__abc_3651_new_n348_), .B(bus_sync_rdata__abc_3651_new_n349_), .C(bus_sync_rdata__abc_3651_new_n265_), .Y(bus_sync_rdata__0reg_data2_31_0__27_));
AOI21X1 AOI21X1_288 ( .A(bus_sync_rdata__abc_3651_new_n351_), .B(bus_sync_rdata__abc_3651_new_n352_), .C(bus_sync_rdata__abc_3651_new_n265_), .Y(bus_sync_rdata__0reg_data2_31_0__28_));
AOI21X1 AOI21X1_289 ( .A(bus_sync_rdata__abc_3651_new_n354_), .B(bus_sync_rdata__abc_3651_new_n355_), .C(bus_sync_rdata__abc_3651_new_n265_), .Y(bus_sync_rdata__0reg_data2_31_0__29_));
AOI21X1 AOI21X1_29 ( .A(_abc_4169_new_n726_), .B(_abc_4169_new_n725_), .C(_abc_4169_new_n729_), .Y(_0bus_cap_31_0__13_));
AOI21X1 AOI21X1_290 ( .A(bus_sync_rdata__abc_3651_new_n357_), .B(bus_sync_rdata__abc_3651_new_n358_), .C(bus_sync_rdata__abc_3651_new_n265_), .Y(bus_sync_rdata__0reg_data2_31_0__30_));
AOI21X1 AOI21X1_291 ( .A(bus_sync_rdata__abc_3651_new_n360_), .B(bus_sync_rdata__abc_3651_new_n361_), .C(bus_sync_rdata__abc_3651_new_n265_), .Y(bus_sync_rdata__0reg_data2_31_0__31_));
AOI21X1 AOI21X1_292 ( .A(bus_sync_state_machine__abc_3817_new_n35_), .B(bus_sync_state_machine__abc_3817_new_n36_), .C(bus_sync_state_machine__abc_3817_new_n33_), .Y(bus_sync_state_machine__0reg_data2_3_0__0_));
AOI21X1 AOI21X1_293 ( .A(bus_sync_state_machine__abc_3817_new_n38_), .B(bus_sync_state_machine__abc_3817_new_n39_), .C(bus_sync_state_machine__abc_3817_new_n33_), .Y(bus_sync_state_machine__0reg_data2_3_0__1_));
AOI21X1 AOI21X1_294 ( .A(bus_sync_state_machine__abc_3817_new_n41_), .B(bus_sync_state_machine__abc_3817_new_n42_), .C(bus_sync_state_machine__abc_3817_new_n33_), .Y(bus_sync_state_machine__0reg_data2_3_0__2_));
AOI21X1 AOI21X1_295 ( .A(bus_sync_state_machine__abc_3817_new_n44_), .B(bus_sync_state_machine__abc_3817_new_n45_), .C(bus_sync_state_machine__abc_3817_new_n33_), .Y(bus_sync_state_machine__0reg_data2_3_0__3_));
AOI21X1 AOI21X1_296 ( .A(bus_sync_status__abc_3630_new_n29_), .B(bus_sync_status__abc_3630_new_n30_), .C(bus_sync_status__abc_3630_new_n27_), .Y(bus_sync_status__0reg_data2_2_0__0_));
AOI21X1 AOI21X1_297 ( .A(bus_sync_status__abc_3630_new_n32_), .B(bus_sync_status__abc_3630_new_n33_), .C(bus_sync_status__abc_3630_new_n27_), .Y(bus_sync_status__0reg_data2_2_0__1_));
AOI21X1 AOI21X1_298 ( .A(bus_sync_status__abc_3630_new_n35_), .B(bus_sync_status__abc_3630_new_n36_), .C(bus_sync_status__abc_3630_new_n27_), .Y(bus_sync_status__0reg_data2_2_0__2_));
AOI21X1 AOI21X1_3 ( .A(_abc_4169_new_n642_), .B(_abc_4169_new_n602_), .C(_abc_4169_new_n646_), .Y(_0bus_cap_31_0__0_));
AOI21X1 AOI21X1_30 ( .A(_abc_4169_new_n651_), .B(bus_cap_13_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n732_));
AOI21X1 AOI21X1_31 ( .A(_abc_4169_new_n732_), .B(_abc_4169_new_n731_), .C(_abc_4169_new_n735_), .Y(_0bus_cap_31_0__14_));
AOI21X1 AOI21X1_32 ( .A(_abc_4169_new_n651_), .B(bus_cap_14_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n738_));
AOI21X1 AOI21X1_33 ( .A(_abc_4169_new_n738_), .B(_abc_4169_new_n737_), .C(_abc_4169_new_n741_), .Y(_0bus_cap_31_0__15_));
AOI21X1 AOI21X1_34 ( .A(_abc_4169_new_n651_), .B(bus_cap_15_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n744_));
AOI21X1 AOI21X1_35 ( .A(_abc_4169_new_n744_), .B(_abc_4169_new_n743_), .C(_abc_4169_new_n747_), .Y(_0bus_cap_31_0__16_));
AOI21X1 AOI21X1_36 ( .A(_abc_4169_new_n651_), .B(bus_cap_16_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n750_));
AOI21X1 AOI21X1_37 ( .A(_abc_4169_new_n750_), .B(_abc_4169_new_n749_), .C(_abc_4169_new_n753_), .Y(_0bus_cap_31_0__17_));
AOI21X1 AOI21X1_38 ( .A(_abc_4169_new_n651_), .B(bus_cap_17_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n756_));
AOI21X1 AOI21X1_39 ( .A(_abc_4169_new_n756_), .B(_abc_4169_new_n755_), .C(_abc_4169_new_n759_), .Y(_0bus_cap_31_0__18_));
AOI21X1 AOI21X1_4 ( .A(_abc_4169_new_n651_), .B(bus_cap_0_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n652_));
AOI21X1 AOI21X1_40 ( .A(_abc_4169_new_n651_), .B(bus_cap_18_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n762_));
AOI21X1 AOI21X1_41 ( .A(_abc_4169_new_n762_), .B(_abc_4169_new_n761_), .C(_abc_4169_new_n765_), .Y(_0bus_cap_31_0__19_));
AOI21X1 AOI21X1_42 ( .A(_abc_4169_new_n651_), .B(bus_cap_19_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n768_));
AOI21X1 AOI21X1_43 ( .A(_abc_4169_new_n768_), .B(_abc_4169_new_n767_), .C(_abc_4169_new_n771_), .Y(_0bus_cap_31_0__20_));
AOI21X1 AOI21X1_44 ( .A(_abc_4169_new_n651_), .B(bus_cap_20_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n774_));
AOI21X1 AOI21X1_45 ( .A(_abc_4169_new_n774_), .B(_abc_4169_new_n773_), .C(_abc_4169_new_n777_), .Y(_0bus_cap_31_0__21_));
AOI21X1 AOI21X1_46 ( .A(_abc_4169_new_n651_), .B(bus_cap_21_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n780_));
AOI21X1 AOI21X1_47 ( .A(_abc_4169_new_n780_), .B(_abc_4169_new_n779_), .C(_abc_4169_new_n783_), .Y(_0bus_cap_31_0__22_));
AOI21X1 AOI21X1_48 ( .A(_abc_4169_new_n651_), .B(bus_cap_22_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n786_));
AOI21X1 AOI21X1_49 ( .A(_abc_4169_new_n786_), .B(_abc_4169_new_n785_), .C(_abc_4169_new_n789_), .Y(_0bus_cap_31_0__23_));
AOI21X1 AOI21X1_5 ( .A(_abc_4169_new_n652_), .B(_abc_4169_new_n648_), .C(_abc_4169_new_n656_), .Y(_0bus_cap_31_0__1_));
AOI21X1 AOI21X1_50 ( .A(_abc_4169_new_n651_), .B(bus_cap_23_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n792_));
AOI21X1 AOI21X1_51 ( .A(_abc_4169_new_n792_), .B(_abc_4169_new_n791_), .C(_abc_4169_new_n795_), .Y(_0bus_cap_31_0__24_));
AOI21X1 AOI21X1_52 ( .A(_abc_4169_new_n651_), .B(bus_cap_24_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n798_));
AOI21X1 AOI21X1_53 ( .A(_abc_4169_new_n798_), .B(_abc_4169_new_n797_), .C(_abc_4169_new_n801_), .Y(_0bus_cap_31_0__25_));
AOI21X1 AOI21X1_54 ( .A(_abc_4169_new_n651_), .B(bus_cap_25_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n804_));
AOI21X1 AOI21X1_55 ( .A(_abc_4169_new_n804_), .B(_abc_4169_new_n803_), .C(_abc_4169_new_n807_), .Y(_0bus_cap_31_0__26_));
AOI21X1 AOI21X1_56 ( .A(_abc_4169_new_n651_), .B(bus_cap_26_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n810_));
AOI21X1 AOI21X1_57 ( .A(_abc_4169_new_n810_), .B(_abc_4169_new_n809_), .C(_abc_4169_new_n813_), .Y(_0bus_cap_31_0__27_));
AOI21X1 AOI21X1_58 ( .A(_abc_4169_new_n651_), .B(bus_cap_27_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n816_));
AOI21X1 AOI21X1_59 ( .A(_abc_4169_new_n816_), .B(_abc_4169_new_n815_), .C(_abc_4169_new_n819_), .Y(_0bus_cap_31_0__28_));
AOI21X1 AOI21X1_6 ( .A(_abc_4169_new_n651_), .B(bus_cap_1_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n659_));
AOI21X1 AOI21X1_60 ( .A(_abc_4169_new_n651_), .B(bus_cap_28_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n822_));
AOI21X1 AOI21X1_61 ( .A(_abc_4169_new_n822_), .B(_abc_4169_new_n821_), .C(_abc_4169_new_n825_), .Y(_0bus_cap_31_0__29_));
AOI21X1 AOI21X1_62 ( .A(_abc_4169_new_n651_), .B(bus_cap_29_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n828_));
AOI21X1 AOI21X1_63 ( .A(_abc_4169_new_n828_), .B(_abc_4169_new_n827_), .C(_abc_4169_new_n831_), .Y(_0bus_cap_31_0__30_));
AOI21X1 AOI21X1_64 ( .A(_abc_4169_new_n651_), .B(bus_cap_30_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n834_));
AOI21X1 AOI21X1_65 ( .A(_abc_4169_new_n834_), .B(_abc_4169_new_n833_), .C(_abc_4169_new_n837_), .Y(_0bus_cap_31_0__31_));
AOI21X1 AOI21X1_66 ( .A(_abc_4169_new_n839_), .B(_abc_4169_new_n840_), .C(_abc_4169_new_n841_), .Y(_0rdata_31_0__0_));
AOI21X1 AOI21X1_67 ( .A(_abc_4169_new_n839_), .B(_abc_4169_new_n843_), .C(_abc_4169_new_n844_), .Y(_0rdata_31_0__1_));
AOI21X1 AOI21X1_68 ( .A(_abc_4169_new_n839_), .B(_abc_4169_new_n846_), .C(_abc_4169_new_n847_), .Y(_0rdata_31_0__2_));
AOI21X1 AOI21X1_69 ( .A(_abc_4169_new_n839_), .B(_abc_4169_new_n849_), .C(_abc_4169_new_n850_), .Y(_0rdata_31_0__3_));
AOI21X1 AOI21X1_7 ( .A(_abc_4169_new_n659_), .B(_abc_4169_new_n658_), .C(_abc_4169_new_n663_), .Y(_0bus_cap_31_0__2_));
AOI21X1 AOI21X1_70 ( .A(_abc_4169_new_n839_), .B(_abc_4169_new_n852_), .C(_abc_4169_new_n853_), .Y(_0rdata_31_0__4_));
AOI21X1 AOI21X1_71 ( .A(_abc_4169_new_n839_), .B(_abc_4169_new_n855_), .C(_abc_4169_new_n856_), .Y(_0rdata_31_0__5_));
AOI21X1 AOI21X1_72 ( .A(_abc_4169_new_n839_), .B(_abc_4169_new_n858_), .C(_abc_4169_new_n859_), .Y(_0rdata_31_0__6_));
AOI21X1 AOI21X1_73 ( .A(_abc_4169_new_n839_), .B(_abc_4169_new_n861_), .C(_abc_4169_new_n862_), .Y(_0rdata_31_0__7_));
AOI21X1 AOI21X1_74 ( .A(_abc_4169_new_n839_), .B(_abc_4169_new_n864_), .C(_abc_4169_new_n865_), .Y(_0rdata_31_0__8_));
AOI21X1 AOI21X1_75 ( .A(_abc_4169_new_n839_), .B(_abc_4169_new_n867_), .C(_abc_4169_new_n868_), .Y(_0rdata_31_0__9_));
AOI21X1 AOI21X1_76 ( .A(_abc_4169_new_n839_), .B(_abc_4169_new_n870_), .C(_abc_4169_new_n871_), .Y(_0rdata_31_0__10_));
AOI21X1 AOI21X1_77 ( .A(_abc_4169_new_n839_), .B(_abc_4169_new_n873_), .C(_abc_4169_new_n874_), .Y(_0rdata_31_0__11_));
AOI21X1 AOI21X1_78 ( .A(_abc_4169_new_n839_), .B(_abc_4169_new_n876_), .C(_abc_4169_new_n877_), .Y(_0rdata_31_0__12_));
AOI21X1 AOI21X1_79 ( .A(_abc_4169_new_n839_), .B(_abc_4169_new_n879_), .C(_abc_4169_new_n880_), .Y(_0rdata_31_0__13_));
AOI21X1 AOI21X1_8 ( .A(_abc_4169_new_n651_), .B(bus_cap_2_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n666_));
AOI21X1 AOI21X1_80 ( .A(_abc_4169_new_n839_), .B(_abc_4169_new_n882_), .C(_abc_4169_new_n883_), .Y(_0rdata_31_0__14_));
AOI21X1 AOI21X1_81 ( .A(_abc_4169_new_n839_), .B(_abc_4169_new_n885_), .C(_abc_4169_new_n886_), .Y(_0rdata_31_0__15_));
AOI21X1 AOI21X1_82 ( .A(_abc_4169_new_n839_), .B(_abc_4169_new_n888_), .C(_abc_4169_new_n889_), .Y(_0rdata_31_0__16_));
AOI21X1 AOI21X1_83 ( .A(_abc_4169_new_n839_), .B(_abc_4169_new_n891_), .C(_abc_4169_new_n892_), .Y(_0rdata_31_0__17_));
AOI21X1 AOI21X1_84 ( .A(_abc_4169_new_n839_), .B(_abc_4169_new_n894_), .C(_abc_4169_new_n895_), .Y(_0rdata_31_0__18_));
AOI21X1 AOI21X1_85 ( .A(_abc_4169_new_n839_), .B(_abc_4169_new_n897_), .C(_abc_4169_new_n898_), .Y(_0rdata_31_0__19_));
AOI21X1 AOI21X1_86 ( .A(_abc_4169_new_n839_), .B(_abc_4169_new_n900_), .C(_abc_4169_new_n901_), .Y(_0rdata_31_0__20_));
AOI21X1 AOI21X1_87 ( .A(_abc_4169_new_n839_), .B(_abc_4169_new_n903_), .C(_abc_4169_new_n904_), .Y(_0rdata_31_0__21_));
AOI21X1 AOI21X1_88 ( .A(_abc_4169_new_n839_), .B(_abc_4169_new_n906_), .C(_abc_4169_new_n907_), .Y(_0rdata_31_0__22_));
AOI21X1 AOI21X1_89 ( .A(_abc_4169_new_n839_), .B(_abc_4169_new_n909_), .C(_abc_4169_new_n910_), .Y(_0rdata_31_0__23_));
AOI21X1 AOI21X1_9 ( .A(_abc_4169_new_n666_), .B(_abc_4169_new_n665_), .C(_abc_4169_new_n669_), .Y(_0bus_cap_31_0__3_));
AOI21X1 AOI21X1_90 ( .A(_abc_4169_new_n839_), .B(_abc_4169_new_n912_), .C(_abc_4169_new_n913_), .Y(_0rdata_31_0__24_));
AOI21X1 AOI21X1_91 ( .A(_abc_4169_new_n839_), .B(_abc_4169_new_n915_), .C(_abc_4169_new_n916_), .Y(_0rdata_31_0__25_));
AOI21X1 AOI21X1_92 ( .A(_abc_4169_new_n839_), .B(_abc_4169_new_n918_), .C(_abc_4169_new_n919_), .Y(_0rdata_31_0__26_));
AOI21X1 AOI21X1_93 ( .A(_abc_4169_new_n839_), .B(_abc_4169_new_n921_), .C(_abc_4169_new_n922_), .Y(_0rdata_31_0__27_));
AOI21X1 AOI21X1_94 ( .A(_abc_4169_new_n839_), .B(_abc_4169_new_n924_), .C(_abc_4169_new_n925_), .Y(_0rdata_31_0__28_));
AOI21X1 AOI21X1_95 ( .A(_abc_4169_new_n839_), .B(_abc_4169_new_n927_), .C(_abc_4169_new_n928_), .Y(_0rdata_31_0__29_));
AOI21X1 AOI21X1_96 ( .A(_abc_4169_new_n839_), .B(_abc_4169_new_n930_), .C(_abc_4169_new_n931_), .Y(_0rdata_31_0__30_));
AOI21X1 AOI21X1_97 ( .A(_abc_4169_new_n839_), .B(_abc_4169_new_n933_), .C(_abc_4169_new_n934_), .Y(_0rdata_31_0__31_));
AOI21X1 AOI21X1_98 ( .A(_abc_4169_new_n936_), .B(_abc_4169_new_n938_), .C(_abc_4169_new_n939_), .Y(_0WDATA_31_0__0_));
AOI21X1 AOI21X1_99 ( .A(_abc_4169_new_n941_), .B(_abc_4169_new_n938_), .C(_abc_4169_new_n942_), .Y(_0WDATA_31_0__1_));
AOI22X1 AOI22X1_1 ( .A(state_5_), .B(axi_awready), .C(state_3_), .D(_abc_4169_new_n565_), .Y(_abc_4169_new_n566_));
AOI22X1 AOI22X1_2 ( .A(state_5_), .B(_abc_4169_new_n593_), .C(state_0_), .D(_abc_4169_new_n594_), .Y(_abc_4169_new_n595_));
AOI22X1 AOI22X1_3 ( .A(_abc_4169_new_n603_), .B(_abc_4169_new_n606_), .C(_abc_4169_new_n649_), .D(_abc_4169_new_n650_), .Y(_abc_4169_new_n651_));
DFFPOSX1 DFFPOSX1_1 ( .CLK(SCLK), .D(_0counter_65_0__0_), .Q(counter_0_));
DFFPOSX1 DFFPOSX1_10 ( .CLK(SCLK), .D(_0counter_65_0__9_), .Q(counter_9_));
DFFPOSX1 DFFPOSX1_100 ( .CLK(CLK), .D(_0rdata_31_0__0_), .Q(bus_sync_rdata_data_in_0_));
DFFPOSX1 DFFPOSX1_101 ( .CLK(CLK), .D(_0rdata_31_0__1_), .Q(bus_sync_rdata_data_in_1_));
DFFPOSX1 DFFPOSX1_102 ( .CLK(CLK), .D(_0rdata_31_0__2_), .Q(bus_sync_rdata_data_in_2_));
DFFPOSX1 DFFPOSX1_103 ( .CLK(CLK), .D(_0rdata_31_0__3_), .Q(bus_sync_rdata_data_in_3_));
DFFPOSX1 DFFPOSX1_104 ( .CLK(CLK), .D(_0rdata_31_0__4_), .Q(bus_sync_rdata_data_in_4_));
DFFPOSX1 DFFPOSX1_105 ( .CLK(CLK), .D(_0rdata_31_0__5_), .Q(bus_sync_rdata_data_in_5_));
DFFPOSX1 DFFPOSX1_106 ( .CLK(CLK), .D(_0rdata_31_0__6_), .Q(bus_sync_rdata_data_in_6_));
DFFPOSX1 DFFPOSX1_107 ( .CLK(CLK), .D(_0rdata_31_0__7_), .Q(bus_sync_rdata_data_in_7_));
DFFPOSX1 DFFPOSX1_108 ( .CLK(CLK), .D(_0rdata_31_0__8_), .Q(bus_sync_rdata_data_in_8_));
DFFPOSX1 DFFPOSX1_109 ( .CLK(CLK), .D(_0rdata_31_0__9_), .Q(bus_sync_rdata_data_in_9_));
DFFPOSX1 DFFPOSX1_11 ( .CLK(SCLK), .D(_0counter_65_0__10_), .Q(counter_10_));
DFFPOSX1 DFFPOSX1_110 ( .CLK(CLK), .D(_0rdata_31_0__10_), .Q(bus_sync_rdata_data_in_10_));
DFFPOSX1 DFFPOSX1_111 ( .CLK(CLK), .D(_0rdata_31_0__11_), .Q(bus_sync_rdata_data_in_11_));
DFFPOSX1 DFFPOSX1_112 ( .CLK(CLK), .D(_0rdata_31_0__12_), .Q(bus_sync_rdata_data_in_12_));
DFFPOSX1 DFFPOSX1_113 ( .CLK(CLK), .D(_0rdata_31_0__13_), .Q(bus_sync_rdata_data_in_13_));
DFFPOSX1 DFFPOSX1_114 ( .CLK(CLK), .D(_0rdata_31_0__14_), .Q(bus_sync_rdata_data_in_14_));
DFFPOSX1 DFFPOSX1_115 ( .CLK(CLK), .D(_0rdata_31_0__15_), .Q(bus_sync_rdata_data_in_15_));
DFFPOSX1 DFFPOSX1_116 ( .CLK(CLK), .D(_0rdata_31_0__16_), .Q(bus_sync_rdata_data_in_16_));
DFFPOSX1 DFFPOSX1_117 ( .CLK(CLK), .D(_0rdata_31_0__17_), .Q(bus_sync_rdata_data_in_17_));
DFFPOSX1 DFFPOSX1_118 ( .CLK(CLK), .D(_0rdata_31_0__18_), .Q(bus_sync_rdata_data_in_18_));
DFFPOSX1 DFFPOSX1_119 ( .CLK(CLK), .D(_0rdata_31_0__19_), .Q(bus_sync_rdata_data_in_19_));
DFFPOSX1 DFFPOSX1_12 ( .CLK(SCLK), .D(_0counter_65_0__11_), .Q(counter_11_));
DFFPOSX1 DFFPOSX1_120 ( .CLK(CLK), .D(_0rdata_31_0__20_), .Q(bus_sync_rdata_data_in_20_));
DFFPOSX1 DFFPOSX1_121 ( .CLK(CLK), .D(_0rdata_31_0__21_), .Q(bus_sync_rdata_data_in_21_));
DFFPOSX1 DFFPOSX1_122 ( .CLK(CLK), .D(_0rdata_31_0__22_), .Q(bus_sync_rdata_data_in_22_));
DFFPOSX1 DFFPOSX1_123 ( .CLK(CLK), .D(_0rdata_31_0__23_), .Q(bus_sync_rdata_data_in_23_));
DFFPOSX1 DFFPOSX1_124 ( .CLK(CLK), .D(_0rdata_31_0__24_), .Q(bus_sync_rdata_data_in_24_));
DFFPOSX1 DFFPOSX1_125 ( .CLK(CLK), .D(_0rdata_31_0__25_), .Q(bus_sync_rdata_data_in_25_));
DFFPOSX1 DFFPOSX1_126 ( .CLK(CLK), .D(_0rdata_31_0__26_), .Q(bus_sync_rdata_data_in_26_));
DFFPOSX1 DFFPOSX1_127 ( .CLK(CLK), .D(_0rdata_31_0__27_), .Q(bus_sync_rdata_data_in_27_));
DFFPOSX1 DFFPOSX1_128 ( .CLK(CLK), .D(_0rdata_31_0__28_), .Q(bus_sync_rdata_data_in_28_));
DFFPOSX1 DFFPOSX1_129 ( .CLK(CLK), .D(_0rdata_31_0__29_), .Q(bus_sync_rdata_data_in_29_));
DFFPOSX1 DFFPOSX1_13 ( .CLK(SCLK), .D(_0counter_65_0__12_), .Q(counter_12_));
DFFPOSX1 DFFPOSX1_130 ( .CLK(CLK), .D(_0rdata_31_0__30_), .Q(bus_sync_rdata_data_in_30_));
DFFPOSX1 DFFPOSX1_131 ( .CLK(CLK), .D(_0rdata_31_0__31_), .Q(bus_sync_rdata_data_in_31_));
DFFPOSX1 DFFPOSX1_132 ( .CLK(SCLK), .D(_0A_ADDR_31_0__0_), .Q(A_ADDR_0_));
DFFPOSX1 DFFPOSX1_133 ( .CLK(SCLK), .D(_0A_ADDR_31_0__1_), .Q(A_ADDR_1_));
DFFPOSX1 DFFPOSX1_134 ( .CLK(SCLK), .D(_0A_ADDR_31_0__2_), .Q(A_ADDR_2_));
DFFPOSX1 DFFPOSX1_135 ( .CLK(SCLK), .D(_0A_ADDR_31_0__3_), .Q(A_ADDR_3_));
DFFPOSX1 DFFPOSX1_136 ( .CLK(SCLK), .D(_0A_ADDR_31_0__4_), .Q(A_ADDR_4_));
DFFPOSX1 DFFPOSX1_137 ( .CLK(SCLK), .D(_0A_ADDR_31_0__5_), .Q(A_ADDR_5_));
DFFPOSX1 DFFPOSX1_138 ( .CLK(SCLK), .D(_0A_ADDR_31_0__6_), .Q(A_ADDR_6_));
DFFPOSX1 DFFPOSX1_139 ( .CLK(SCLK), .D(_0A_ADDR_31_0__7_), .Q(A_ADDR_7_));
DFFPOSX1 DFFPOSX1_14 ( .CLK(SCLK), .D(_0counter_65_0__13_), .Q(counter_13_));
DFFPOSX1 DFFPOSX1_140 ( .CLK(SCLK), .D(_0A_ADDR_31_0__8_), .Q(A_ADDR_8_));
DFFPOSX1 DFFPOSX1_141 ( .CLK(SCLK), .D(_0A_ADDR_31_0__9_), .Q(A_ADDR_9_));
DFFPOSX1 DFFPOSX1_142 ( .CLK(SCLK), .D(_0A_ADDR_31_0__10_), .Q(A_ADDR_10_));
DFFPOSX1 DFFPOSX1_143 ( .CLK(SCLK), .D(_0A_ADDR_31_0__11_), .Q(A_ADDR_11_));
DFFPOSX1 DFFPOSX1_144 ( .CLK(SCLK), .D(_0A_ADDR_31_0__12_), .Q(A_ADDR_12_));
DFFPOSX1 DFFPOSX1_145 ( .CLK(SCLK), .D(_0A_ADDR_31_0__13_), .Q(A_ADDR_13_));
DFFPOSX1 DFFPOSX1_146 ( .CLK(SCLK), .D(_0A_ADDR_31_0__14_), .Q(A_ADDR_14_));
DFFPOSX1 DFFPOSX1_147 ( .CLK(SCLK), .D(_0A_ADDR_31_0__15_), .Q(A_ADDR_15_));
DFFPOSX1 DFFPOSX1_148 ( .CLK(SCLK), .D(_0A_ADDR_31_0__16_), .Q(A_ADDR_16_));
DFFPOSX1 DFFPOSX1_149 ( .CLK(SCLK), .D(_0A_ADDR_31_0__17_), .Q(A_ADDR_17_));
DFFPOSX1 DFFPOSX1_15 ( .CLK(SCLK), .D(_0counter_65_0__14_), .Q(counter_14_));
DFFPOSX1 DFFPOSX1_150 ( .CLK(SCLK), .D(_0A_ADDR_31_0__18_), .Q(A_ADDR_18_));
DFFPOSX1 DFFPOSX1_151 ( .CLK(SCLK), .D(_0A_ADDR_31_0__19_), .Q(A_ADDR_19_));
DFFPOSX1 DFFPOSX1_152 ( .CLK(SCLK), .D(_0A_ADDR_31_0__20_), .Q(A_ADDR_20_));
DFFPOSX1 DFFPOSX1_153 ( .CLK(SCLK), .D(_0A_ADDR_31_0__21_), .Q(A_ADDR_21_));
DFFPOSX1 DFFPOSX1_154 ( .CLK(SCLK), .D(_0A_ADDR_31_0__22_), .Q(A_ADDR_22_));
DFFPOSX1 DFFPOSX1_155 ( .CLK(SCLK), .D(_0A_ADDR_31_0__23_), .Q(A_ADDR_23_));
DFFPOSX1 DFFPOSX1_156 ( .CLK(SCLK), .D(_0A_ADDR_31_0__24_), .Q(A_ADDR_24_));
DFFPOSX1 DFFPOSX1_157 ( .CLK(SCLK), .D(_0A_ADDR_31_0__25_), .Q(A_ADDR_25_));
DFFPOSX1 DFFPOSX1_158 ( .CLK(SCLK), .D(_0A_ADDR_31_0__26_), .Q(A_ADDR_26_));
DFFPOSX1 DFFPOSX1_159 ( .CLK(SCLK), .D(_0A_ADDR_31_0__27_), .Q(A_ADDR_27_));
DFFPOSX1 DFFPOSX1_16 ( .CLK(SCLK), .D(_0counter_65_0__15_), .Q(counter_15_));
DFFPOSX1 DFFPOSX1_160 ( .CLK(SCLK), .D(_0A_ADDR_31_0__28_), .Q(A_ADDR_28_));
DFFPOSX1 DFFPOSX1_161 ( .CLK(SCLK), .D(_0A_ADDR_31_0__29_), .Q(A_ADDR_29_));
DFFPOSX1 DFFPOSX1_162 ( .CLK(SCLK), .D(_0A_ADDR_31_0__30_), .Q(A_ADDR_30_));
DFFPOSX1 DFFPOSX1_163 ( .CLK(SCLK), .D(_0A_ADDR_31_0__31_), .Q(A_ADDR_31_));
DFFPOSX1 DFFPOSX1_164 ( .CLK(SCLK), .D(_0WDATA_31_0__0_), .Q(WDATA_0_));
DFFPOSX1 DFFPOSX1_165 ( .CLK(SCLK), .D(_0WDATA_31_0__1_), .Q(WDATA_1_));
DFFPOSX1 DFFPOSX1_166 ( .CLK(SCLK), .D(_0WDATA_31_0__2_), .Q(WDATA_2_));
DFFPOSX1 DFFPOSX1_167 ( .CLK(SCLK), .D(_0WDATA_31_0__3_), .Q(WDATA_3_));
DFFPOSX1 DFFPOSX1_168 ( .CLK(SCLK), .D(_0WDATA_31_0__4_), .Q(WDATA_4_));
DFFPOSX1 DFFPOSX1_169 ( .CLK(SCLK), .D(_0WDATA_31_0__5_), .Q(WDATA_5_));
DFFPOSX1 DFFPOSX1_17 ( .CLK(SCLK), .D(_0counter_65_0__16_), .Q(counter_16_));
DFFPOSX1 DFFPOSX1_170 ( .CLK(SCLK), .D(_0WDATA_31_0__6_), .Q(WDATA_6_));
DFFPOSX1 DFFPOSX1_171 ( .CLK(SCLK), .D(_0WDATA_31_0__7_), .Q(WDATA_7_));
DFFPOSX1 DFFPOSX1_172 ( .CLK(SCLK), .D(_0WDATA_31_0__8_), .Q(WDATA_8_));
DFFPOSX1 DFFPOSX1_173 ( .CLK(SCLK), .D(_0WDATA_31_0__9_), .Q(WDATA_9_));
DFFPOSX1 DFFPOSX1_174 ( .CLK(SCLK), .D(_0WDATA_31_0__10_), .Q(WDATA_10_));
DFFPOSX1 DFFPOSX1_175 ( .CLK(SCLK), .D(_0WDATA_31_0__11_), .Q(WDATA_11_));
DFFPOSX1 DFFPOSX1_176 ( .CLK(SCLK), .D(_0WDATA_31_0__12_), .Q(WDATA_12_));
DFFPOSX1 DFFPOSX1_177 ( .CLK(SCLK), .D(_0WDATA_31_0__13_), .Q(WDATA_13_));
DFFPOSX1 DFFPOSX1_178 ( .CLK(SCLK), .D(_0WDATA_31_0__14_), .Q(WDATA_14_));
DFFPOSX1 DFFPOSX1_179 ( .CLK(SCLK), .D(_0WDATA_31_0__15_), .Q(WDATA_15_));
DFFPOSX1 DFFPOSX1_18 ( .CLK(SCLK), .D(_0counter_65_0__17_), .Q(counter_17_));
DFFPOSX1 DFFPOSX1_180 ( .CLK(SCLK), .D(_0WDATA_31_0__16_), .Q(WDATA_16_));
DFFPOSX1 DFFPOSX1_181 ( .CLK(SCLK), .D(_0WDATA_31_0__17_), .Q(WDATA_17_));
DFFPOSX1 DFFPOSX1_182 ( .CLK(SCLK), .D(_0WDATA_31_0__18_), .Q(WDATA_18_));
DFFPOSX1 DFFPOSX1_183 ( .CLK(SCLK), .D(_0WDATA_31_0__19_), .Q(WDATA_19_));
DFFPOSX1 DFFPOSX1_184 ( .CLK(SCLK), .D(_0WDATA_31_0__20_), .Q(WDATA_20_));
DFFPOSX1 DFFPOSX1_185 ( .CLK(SCLK), .D(_0WDATA_31_0__21_), .Q(WDATA_21_));
DFFPOSX1 DFFPOSX1_186 ( .CLK(SCLK), .D(_0WDATA_31_0__22_), .Q(WDATA_22_));
DFFPOSX1 DFFPOSX1_187 ( .CLK(SCLK), .D(_0WDATA_31_0__23_), .Q(WDATA_23_));
DFFPOSX1 DFFPOSX1_188 ( .CLK(SCLK), .D(_0WDATA_31_0__24_), .Q(WDATA_24_));
DFFPOSX1 DFFPOSX1_189 ( .CLK(SCLK), .D(_0WDATA_31_0__25_), .Q(WDATA_25_));
DFFPOSX1 DFFPOSX1_19 ( .CLK(SCLK), .D(_0counter_65_0__18_), .Q(counter_18_));
DFFPOSX1 DFFPOSX1_190 ( .CLK(SCLK), .D(_0WDATA_31_0__26_), .Q(WDATA_26_));
DFFPOSX1 DFFPOSX1_191 ( .CLK(SCLK), .D(_0WDATA_31_0__27_), .Q(WDATA_27_));
DFFPOSX1 DFFPOSX1_192 ( .CLK(SCLK), .D(_0WDATA_31_0__28_), .Q(WDATA_28_));
DFFPOSX1 DFFPOSX1_193 ( .CLK(SCLK), .D(_0WDATA_31_0__29_), .Q(WDATA_29_));
DFFPOSX1 DFFPOSX1_194 ( .CLK(SCLK), .D(_0WDATA_31_0__30_), .Q(WDATA_30_));
DFFPOSX1 DFFPOSX1_195 ( .CLK(SCLK), .D(_0WDATA_31_0__31_), .Q(WDATA_31_));
DFFPOSX1 DFFPOSX1_196 ( .CLK(SCLK), .D(_0PICORV_RST_SPI_0_0_), .Q(PICORV_RST_SPI));
DFFPOSX1 DFFPOSX1_197 ( .CLK(SCLK), .D(_0we_0_0_), .Q(we));
DFFPOSX1 DFFPOSX1_198 ( .CLK(SCLK), .D(_0re_0_0_), .Q(re));
DFFPOSX1 DFFPOSX1_199 ( .CLK(SCLK), .D(_0sft_reg_65_0__0_), .Q(sft_reg_0_));
DFFPOSX1 DFFPOSX1_2 ( .CLK(SCLK), .D(_0counter_65_0__1_), .Q(counter_1_));
DFFPOSX1 DFFPOSX1_20 ( .CLK(SCLK), .D(_0counter_65_0__19_), .Q(counter_19_));
DFFPOSX1 DFFPOSX1_200 ( .CLK(SCLK), .D(_0sft_reg_65_0__1_), .Q(sft_reg_1_));
DFFPOSX1 DFFPOSX1_201 ( .CLK(SCLK), .D(_0sft_reg_65_0__2_), .Q(sft_reg_2_));
DFFPOSX1 DFFPOSX1_202 ( .CLK(SCLK), .D(_0sft_reg_65_0__3_), .Q(sft_reg_3_));
DFFPOSX1 DFFPOSX1_203 ( .CLK(SCLK), .D(_0sft_reg_65_0__4_), .Q(sft_reg_4_));
DFFPOSX1 DFFPOSX1_204 ( .CLK(SCLK), .D(_0sft_reg_65_0__5_), .Q(sft_reg_5_));
DFFPOSX1 DFFPOSX1_205 ( .CLK(SCLK), .D(_0sft_reg_65_0__6_), .Q(sft_reg_6_));
DFFPOSX1 DFFPOSX1_206 ( .CLK(SCLK), .D(_0sft_reg_65_0__7_), .Q(sft_reg_7_));
DFFPOSX1 DFFPOSX1_207 ( .CLK(SCLK), .D(_0sft_reg_65_0__8_), .Q(sft_reg_8_));
DFFPOSX1 DFFPOSX1_208 ( .CLK(SCLK), .D(_0sft_reg_65_0__9_), .Q(sft_reg_9_));
DFFPOSX1 DFFPOSX1_209 ( .CLK(SCLK), .D(_0sft_reg_65_0__10_), .Q(sft_reg_10_));
DFFPOSX1 DFFPOSX1_21 ( .CLK(SCLK), .D(_0counter_65_0__20_), .Q(counter_20_));
DFFPOSX1 DFFPOSX1_210 ( .CLK(SCLK), .D(_0sft_reg_65_0__11_), .Q(sft_reg_11_));
DFFPOSX1 DFFPOSX1_211 ( .CLK(SCLK), .D(_0sft_reg_65_0__12_), .Q(sft_reg_12_));
DFFPOSX1 DFFPOSX1_212 ( .CLK(SCLK), .D(_0sft_reg_65_0__13_), .Q(sft_reg_13_));
DFFPOSX1 DFFPOSX1_213 ( .CLK(SCLK), .D(_0sft_reg_65_0__14_), .Q(sft_reg_14_));
DFFPOSX1 DFFPOSX1_214 ( .CLK(SCLK), .D(_0sft_reg_65_0__15_), .Q(sft_reg_15_));
DFFPOSX1 DFFPOSX1_215 ( .CLK(SCLK), .D(_0sft_reg_65_0__16_), .Q(sft_reg_16_));
DFFPOSX1 DFFPOSX1_216 ( .CLK(SCLK), .D(_0sft_reg_65_0__17_), .Q(sft_reg_17_));
DFFPOSX1 DFFPOSX1_217 ( .CLK(SCLK), .D(_0sft_reg_65_0__18_), .Q(sft_reg_18_));
DFFPOSX1 DFFPOSX1_218 ( .CLK(SCLK), .D(_0sft_reg_65_0__19_), .Q(sft_reg_19_));
DFFPOSX1 DFFPOSX1_219 ( .CLK(SCLK), .D(_0sft_reg_65_0__20_), .Q(sft_reg_20_));
DFFPOSX1 DFFPOSX1_22 ( .CLK(SCLK), .D(_0counter_65_0__21_), .Q(counter_21_));
DFFPOSX1 DFFPOSX1_220 ( .CLK(SCLK), .D(_0sft_reg_65_0__21_), .Q(sft_reg_21_));
DFFPOSX1 DFFPOSX1_221 ( .CLK(SCLK), .D(_0sft_reg_65_0__22_), .Q(sft_reg_22_));
DFFPOSX1 DFFPOSX1_222 ( .CLK(SCLK), .D(_0sft_reg_65_0__23_), .Q(sft_reg_23_));
DFFPOSX1 DFFPOSX1_223 ( .CLK(SCLK), .D(_0sft_reg_65_0__24_), .Q(sft_reg_24_));
DFFPOSX1 DFFPOSX1_224 ( .CLK(SCLK), .D(_0sft_reg_65_0__25_), .Q(sft_reg_25_));
DFFPOSX1 DFFPOSX1_225 ( .CLK(SCLK), .D(_0sft_reg_65_0__26_), .Q(sft_reg_26_));
DFFPOSX1 DFFPOSX1_226 ( .CLK(SCLK), .D(_0sft_reg_65_0__27_), .Q(sft_reg_27_));
DFFPOSX1 DFFPOSX1_227 ( .CLK(SCLK), .D(_0sft_reg_65_0__28_), .Q(sft_reg_28_));
DFFPOSX1 DFFPOSX1_228 ( .CLK(SCLK), .D(_0sft_reg_65_0__29_), .Q(sft_reg_29_));
DFFPOSX1 DFFPOSX1_229 ( .CLK(SCLK), .D(_0sft_reg_65_0__30_), .Q(sft_reg_30_));
DFFPOSX1 DFFPOSX1_23 ( .CLK(SCLK), .D(_0counter_65_0__22_), .Q(counter_22_));
DFFPOSX1 DFFPOSX1_230 ( .CLK(CLK), .D(_abc_2903_auto_fsm_map_cc_170_map_fsm_402_0_), .Q(state_0_));
DFFPOSX1 DFFPOSX1_231 ( .CLK(CLK), .D(_abc_2903_auto_fsm_map_cc_170_map_fsm_402_1_), .Q(state_1_));
DFFPOSX1 DFFPOSX1_232 ( .CLK(CLK), .D(_abc_2903_auto_fsm_map_cc_118_implement_pattern_cache_430), .Q(axi_bready));
DFFPOSX1 DFFPOSX1_233 ( .CLK(CLK), .D(_abc_2903_auto_fsm_map_cc_170_map_fsm_402_3_), .Q(state_3_));
DFFPOSX1 DFFPOSX1_234 ( .CLK(CLK), .D(_abc_2903_auto_fsm_map_cc_170_map_fsm_402_4_), .Q(state_4_));
DFFPOSX1 DFFPOSX1_235 ( .CLK(CLK), .D(_abc_2903_auto_fsm_map_cc_170_map_fsm_402_5_), .Q(state_5_));
DFFPOSX1 DFFPOSX1_236 ( .CLK(CLK), .D(_abc_2903_auto_fsm_map_cc_170_map_fsm_402_6_), .Q(state_6_));
DFFPOSX1 DFFPOSX1_237 ( .CLK(CLK), .D(_abc_2903_auto_fsm_map_cc_170_map_fsm_402_7_), .Q(state_7_));
DFFPOSX1 DFFPOSX1_238 ( .CLK(CLK), .D(_abc_2903_auto_fsm_map_cc_118_implement_pattern_cache_479), .Q(axi_rready));
DFFPOSX1 DFFPOSX1_239 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__0_), .Q(bus_sync_axi_bus_reg_data2_0_));
DFFPOSX1 DFFPOSX1_24 ( .CLK(SCLK), .D(_0counter_65_0__23_), .Q(counter_23_));
DFFPOSX1 DFFPOSX1_240 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__1_), .Q(bus_sync_axi_bus_reg_data2_1_));
DFFPOSX1 DFFPOSX1_241 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__2_), .Q(bus_sync_axi_bus_reg_data2_2_));
DFFPOSX1 DFFPOSX1_242 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__3_), .Q(bus_sync_axi_bus_reg_data2_3_));
DFFPOSX1 DFFPOSX1_243 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__4_), .Q(bus_sync_axi_bus_reg_data2_4_));
DFFPOSX1 DFFPOSX1_244 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__5_), .Q(bus_sync_axi_bus_reg_data2_5_));
DFFPOSX1 DFFPOSX1_245 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__6_), .Q(bus_sync_axi_bus_reg_data2_6_));
DFFPOSX1 DFFPOSX1_246 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__7_), .Q(bus_sync_axi_bus_reg_data2_7_));
DFFPOSX1 DFFPOSX1_247 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__8_), .Q(bus_sync_axi_bus_reg_data2_8_));
DFFPOSX1 DFFPOSX1_248 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__9_), .Q(bus_sync_axi_bus_reg_data2_9_));
DFFPOSX1 DFFPOSX1_249 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__10_), .Q(bus_sync_axi_bus_reg_data2_10_));
DFFPOSX1 DFFPOSX1_25 ( .CLK(SCLK), .D(_0counter_65_0__24_), .Q(counter_24_));
DFFPOSX1 DFFPOSX1_250 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__11_), .Q(bus_sync_axi_bus_reg_data2_11_));
DFFPOSX1 DFFPOSX1_251 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__12_), .Q(bus_sync_axi_bus_reg_data2_12_));
DFFPOSX1 DFFPOSX1_252 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__13_), .Q(bus_sync_axi_bus_reg_data2_13_));
DFFPOSX1 DFFPOSX1_253 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__14_), .Q(bus_sync_axi_bus_reg_data2_14_));
DFFPOSX1 DFFPOSX1_254 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__15_), .Q(bus_sync_axi_bus_reg_data2_15_));
DFFPOSX1 DFFPOSX1_255 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__16_), .Q(bus_sync_axi_bus_reg_data2_16_));
DFFPOSX1 DFFPOSX1_256 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__17_), .Q(bus_sync_axi_bus_reg_data2_17_));
DFFPOSX1 DFFPOSX1_257 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__18_), .Q(bus_sync_axi_bus_reg_data2_18_));
DFFPOSX1 DFFPOSX1_258 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__19_), .Q(bus_sync_axi_bus_reg_data2_19_));
DFFPOSX1 DFFPOSX1_259 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__20_), .Q(bus_sync_axi_bus_reg_data2_20_));
DFFPOSX1 DFFPOSX1_26 ( .CLK(SCLK), .D(_0counter_65_0__25_), .Q(counter_25_));
DFFPOSX1 DFFPOSX1_260 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__21_), .Q(bus_sync_axi_bus_reg_data2_21_));
DFFPOSX1 DFFPOSX1_261 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__22_), .Q(bus_sync_axi_bus_reg_data2_22_));
DFFPOSX1 DFFPOSX1_262 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__23_), .Q(bus_sync_axi_bus_reg_data2_23_));
DFFPOSX1 DFFPOSX1_263 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__24_), .Q(bus_sync_axi_bus_reg_data2_24_));
DFFPOSX1 DFFPOSX1_264 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__25_), .Q(bus_sync_axi_bus_reg_data2_25_));
DFFPOSX1 DFFPOSX1_265 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__26_), .Q(bus_sync_axi_bus_reg_data2_26_));
DFFPOSX1 DFFPOSX1_266 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__27_), .Q(bus_sync_axi_bus_reg_data2_27_));
DFFPOSX1 DFFPOSX1_267 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__28_), .Q(bus_sync_axi_bus_reg_data2_28_));
DFFPOSX1 DFFPOSX1_268 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__29_), .Q(bus_sync_axi_bus_reg_data2_29_));
DFFPOSX1 DFFPOSX1_269 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__30_), .Q(bus_sync_axi_bus_reg_data2_30_));
DFFPOSX1 DFFPOSX1_27 ( .CLK(SCLK), .D(_0counter_65_0__26_), .Q(counter_26_));
DFFPOSX1 DFFPOSX1_270 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__31_), .Q(bus_sync_axi_bus_reg_data2_31_));
DFFPOSX1 DFFPOSX1_271 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__32_), .Q(bus_sync_axi_bus_reg_data2_32_));
DFFPOSX1 DFFPOSX1_272 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__33_), .Q(bus_sync_axi_bus_reg_data2_33_));
DFFPOSX1 DFFPOSX1_273 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__34_), .Q(bus_sync_axi_bus_reg_data2_34_));
DFFPOSX1 DFFPOSX1_274 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__35_), .Q(bus_sync_axi_bus_reg_data2_35_));
DFFPOSX1 DFFPOSX1_275 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__36_), .Q(bus_sync_axi_bus_reg_data2_36_));
DFFPOSX1 DFFPOSX1_276 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__37_), .Q(bus_sync_axi_bus_reg_data2_37_));
DFFPOSX1 DFFPOSX1_277 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__38_), .Q(bus_sync_axi_bus_reg_data2_38_));
DFFPOSX1 DFFPOSX1_278 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__39_), .Q(bus_sync_axi_bus_reg_data2_39_));
DFFPOSX1 DFFPOSX1_279 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__40_), .Q(bus_sync_axi_bus_reg_data2_40_));
DFFPOSX1 DFFPOSX1_28 ( .CLK(SCLK), .D(_0counter_65_0__27_), .Q(counter_27_));
DFFPOSX1 DFFPOSX1_280 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__41_), .Q(bus_sync_axi_bus_reg_data2_41_));
DFFPOSX1 DFFPOSX1_281 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__42_), .Q(bus_sync_axi_bus_reg_data2_42_));
DFFPOSX1 DFFPOSX1_282 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__43_), .Q(bus_sync_axi_bus_reg_data2_43_));
DFFPOSX1 DFFPOSX1_283 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__44_), .Q(bus_sync_axi_bus_reg_data2_44_));
DFFPOSX1 DFFPOSX1_284 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__45_), .Q(bus_sync_axi_bus_reg_data2_45_));
DFFPOSX1 DFFPOSX1_285 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__46_), .Q(bus_sync_axi_bus_reg_data2_46_));
DFFPOSX1 DFFPOSX1_286 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__47_), .Q(bus_sync_axi_bus_reg_data2_47_));
DFFPOSX1 DFFPOSX1_287 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__48_), .Q(bus_sync_axi_bus_reg_data2_48_));
DFFPOSX1 DFFPOSX1_288 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__49_), .Q(bus_sync_axi_bus_reg_data2_49_));
DFFPOSX1 DFFPOSX1_289 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__50_), .Q(bus_sync_axi_bus_reg_data2_50_));
DFFPOSX1 DFFPOSX1_29 ( .CLK(SCLK), .D(_0counter_65_0__28_), .Q(counter_28_));
DFFPOSX1 DFFPOSX1_290 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__51_), .Q(bus_sync_axi_bus_reg_data2_51_));
DFFPOSX1 DFFPOSX1_291 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__52_), .Q(bus_sync_axi_bus_reg_data2_52_));
DFFPOSX1 DFFPOSX1_292 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__53_), .Q(bus_sync_axi_bus_reg_data2_53_));
DFFPOSX1 DFFPOSX1_293 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__54_), .Q(bus_sync_axi_bus_reg_data2_54_));
DFFPOSX1 DFFPOSX1_294 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__55_), .Q(bus_sync_axi_bus_reg_data2_55_));
DFFPOSX1 DFFPOSX1_295 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__56_), .Q(bus_sync_axi_bus_reg_data2_56_));
DFFPOSX1 DFFPOSX1_296 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__57_), .Q(bus_sync_axi_bus_reg_data2_57_));
DFFPOSX1 DFFPOSX1_297 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__58_), .Q(bus_sync_axi_bus_reg_data2_58_));
DFFPOSX1 DFFPOSX1_298 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__59_), .Q(bus_sync_axi_bus_reg_data2_59_));
DFFPOSX1 DFFPOSX1_299 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__60_), .Q(bus_sync_axi_bus_reg_data2_60_));
DFFPOSX1 DFFPOSX1_3 ( .CLK(SCLK), .D(_0counter_65_0__2_), .Q(counter_2_));
DFFPOSX1 DFFPOSX1_30 ( .CLK(SCLK), .D(_0counter_65_0__29_), .Q(counter_29_));
DFFPOSX1 DFFPOSX1_300 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__61_), .Q(bus_sync_axi_bus_reg_data2_61_));
DFFPOSX1 DFFPOSX1_301 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__62_), .Q(bus_sync_axi_bus_reg_data2_62_));
DFFPOSX1 DFFPOSX1_302 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__63_), .Q(bus_sync_axi_bus_reg_data2_63_));
DFFPOSX1 DFFPOSX1_303 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__0_), .Q(\axi_wdata[0] ));
DFFPOSX1 DFFPOSX1_304 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__1_), .Q(\axi_wdata[1] ));
DFFPOSX1 DFFPOSX1_305 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__2_), .Q(\axi_wdata[2] ));
DFFPOSX1 DFFPOSX1_306 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__3_), .Q(\axi_wdata[3] ));
DFFPOSX1 DFFPOSX1_307 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__4_), .Q(\axi_wdata[4] ));
DFFPOSX1 DFFPOSX1_308 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__5_), .Q(\axi_wdata[5] ));
DFFPOSX1 DFFPOSX1_309 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__6_), .Q(\axi_wdata[6] ));
DFFPOSX1 DFFPOSX1_31 ( .CLK(SCLK), .D(_0counter_65_0__30_), .Q(counter_30_));
DFFPOSX1 DFFPOSX1_310 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__7_), .Q(\axi_wdata[7] ));
DFFPOSX1 DFFPOSX1_311 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__8_), .Q(\axi_wdata[8] ));
DFFPOSX1 DFFPOSX1_312 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__9_), .Q(\axi_wdata[9] ));
DFFPOSX1 DFFPOSX1_313 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__10_), .Q(\axi_wdata[10] ));
DFFPOSX1 DFFPOSX1_314 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__11_), .Q(\axi_wdata[11] ));
DFFPOSX1 DFFPOSX1_315 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__12_), .Q(\axi_wdata[12] ));
DFFPOSX1 DFFPOSX1_316 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__13_), .Q(\axi_wdata[13] ));
DFFPOSX1 DFFPOSX1_317 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__14_), .Q(\axi_wdata[14] ));
DFFPOSX1 DFFPOSX1_318 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__15_), .Q(\axi_wdata[15] ));
DFFPOSX1 DFFPOSX1_319 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__16_), .Q(\axi_wdata[16] ));
DFFPOSX1 DFFPOSX1_32 ( .CLK(SCLK), .D(_0counter_65_0__31_), .Q(counter_31_));
DFFPOSX1 DFFPOSX1_320 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__17_), .Q(\axi_wdata[17] ));
DFFPOSX1 DFFPOSX1_321 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__18_), .Q(\axi_wdata[18] ));
DFFPOSX1 DFFPOSX1_322 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__19_), .Q(\axi_wdata[19] ));
DFFPOSX1 DFFPOSX1_323 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__20_), .Q(\axi_wdata[20] ));
DFFPOSX1 DFFPOSX1_324 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__21_), .Q(\axi_wdata[21] ));
DFFPOSX1 DFFPOSX1_325 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__22_), .Q(\axi_wdata[22] ));
DFFPOSX1 DFFPOSX1_326 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__23_), .Q(\axi_wdata[23] ));
DFFPOSX1 DFFPOSX1_327 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__24_), .Q(\axi_wdata[24] ));
DFFPOSX1 DFFPOSX1_328 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__25_), .Q(\axi_wdata[25] ));
DFFPOSX1 DFFPOSX1_329 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__26_), .Q(\axi_wdata[26] ));
DFFPOSX1 DFFPOSX1_33 ( .CLK(SCLK), .D(_0counter_65_0__32_), .Q(counter_32_));
DFFPOSX1 DFFPOSX1_330 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__27_), .Q(\axi_wdata[27] ));
DFFPOSX1 DFFPOSX1_331 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__28_), .Q(\axi_wdata[28] ));
DFFPOSX1 DFFPOSX1_332 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__29_), .Q(\axi_wdata[29] ));
DFFPOSX1 DFFPOSX1_333 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__30_), .Q(\axi_wdata[30] ));
DFFPOSX1 DFFPOSX1_334 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__31_), .Q(\axi_wdata[31] ));
DFFPOSX1 DFFPOSX1_335 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__32_), .Q(\axi_araddr[0] ));
DFFPOSX1 DFFPOSX1_336 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__33_), .Q(\axi_araddr[1] ));
DFFPOSX1 DFFPOSX1_337 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__34_), .Q(\axi_araddr[2] ));
DFFPOSX1 DFFPOSX1_338 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__35_), .Q(\axi_araddr[3] ));
DFFPOSX1 DFFPOSX1_339 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__36_), .Q(\axi_araddr[4] ));
DFFPOSX1 DFFPOSX1_34 ( .CLK(SCLK), .D(_0counter_65_0__33_), .Q(counter_33_));
DFFPOSX1 DFFPOSX1_340 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__37_), .Q(\axi_araddr[5] ));
DFFPOSX1 DFFPOSX1_341 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__38_), .Q(\axi_araddr[6] ));
DFFPOSX1 DFFPOSX1_342 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__39_), .Q(\axi_araddr[7] ));
DFFPOSX1 DFFPOSX1_343 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__40_), .Q(\axi_araddr[8] ));
DFFPOSX1 DFFPOSX1_344 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__41_), .Q(\axi_araddr[9] ));
DFFPOSX1 DFFPOSX1_345 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__42_), .Q(\axi_araddr[10] ));
DFFPOSX1 DFFPOSX1_346 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__43_), .Q(\axi_araddr[11] ));
DFFPOSX1 DFFPOSX1_347 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__44_), .Q(\axi_araddr[12] ));
DFFPOSX1 DFFPOSX1_348 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__45_), .Q(\axi_araddr[13] ));
DFFPOSX1 DFFPOSX1_349 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__46_), .Q(\axi_araddr[14] ));
DFFPOSX1 DFFPOSX1_35 ( .CLK(SCLK), .D(_0counter_65_0__34_), .Q(counter_34_));
DFFPOSX1 DFFPOSX1_350 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__47_), .Q(\axi_araddr[15] ));
DFFPOSX1 DFFPOSX1_351 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__48_), .Q(\axi_araddr[16] ));
DFFPOSX1 DFFPOSX1_352 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__49_), .Q(\axi_araddr[17] ));
DFFPOSX1 DFFPOSX1_353 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__50_), .Q(\axi_araddr[18] ));
DFFPOSX1 DFFPOSX1_354 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__51_), .Q(\axi_araddr[19] ));
DFFPOSX1 DFFPOSX1_355 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__52_), .Q(\axi_araddr[20] ));
DFFPOSX1 DFFPOSX1_356 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__53_), .Q(\axi_araddr[21] ));
DFFPOSX1 DFFPOSX1_357 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__54_), .Q(\axi_araddr[22] ));
DFFPOSX1 DFFPOSX1_358 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__55_), .Q(\axi_araddr[23] ));
DFFPOSX1 DFFPOSX1_359 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__56_), .Q(\axi_araddr[24] ));
DFFPOSX1 DFFPOSX1_36 ( .CLK(SCLK), .D(_0counter_65_0__35_), .Q(counter_35_));
DFFPOSX1 DFFPOSX1_360 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__57_), .Q(\axi_araddr[25] ));
DFFPOSX1 DFFPOSX1_361 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__58_), .Q(\axi_araddr[26] ));
DFFPOSX1 DFFPOSX1_362 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__59_), .Q(\axi_araddr[27] ));
DFFPOSX1 DFFPOSX1_363 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__60_), .Q(\axi_araddr[28] ));
DFFPOSX1 DFFPOSX1_364 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__61_), .Q(\axi_araddr[29] ));
DFFPOSX1 DFFPOSX1_365 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__62_), .Q(\axi_araddr[30] ));
DFFPOSX1 DFFPOSX1_366 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__63_), .Q(\axi_araddr[31] ));
DFFPOSX1 DFFPOSX1_367 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__0_), .Q(bus_sync_axi_bus_reg_data1_0_));
DFFPOSX1 DFFPOSX1_368 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__1_), .Q(bus_sync_axi_bus_reg_data1_1_));
DFFPOSX1 DFFPOSX1_369 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__2_), .Q(bus_sync_axi_bus_reg_data1_2_));
DFFPOSX1 DFFPOSX1_37 ( .CLK(SCLK), .D(_0counter_65_0__36_), .Q(counter_36_));
DFFPOSX1 DFFPOSX1_370 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__3_), .Q(bus_sync_axi_bus_reg_data1_3_));
DFFPOSX1 DFFPOSX1_371 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__4_), .Q(bus_sync_axi_bus_reg_data1_4_));
DFFPOSX1 DFFPOSX1_372 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__5_), .Q(bus_sync_axi_bus_reg_data1_5_));
DFFPOSX1 DFFPOSX1_373 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__6_), .Q(bus_sync_axi_bus_reg_data1_6_));
DFFPOSX1 DFFPOSX1_374 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__7_), .Q(bus_sync_axi_bus_reg_data1_7_));
DFFPOSX1 DFFPOSX1_375 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__8_), .Q(bus_sync_axi_bus_reg_data1_8_));
DFFPOSX1 DFFPOSX1_376 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__9_), .Q(bus_sync_axi_bus_reg_data1_9_));
DFFPOSX1 DFFPOSX1_377 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__10_), .Q(bus_sync_axi_bus_reg_data1_10_));
DFFPOSX1 DFFPOSX1_378 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__11_), .Q(bus_sync_axi_bus_reg_data1_11_));
DFFPOSX1 DFFPOSX1_379 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__12_), .Q(bus_sync_axi_bus_reg_data1_12_));
DFFPOSX1 DFFPOSX1_38 ( .CLK(SCLK), .D(_0counter_65_0__37_), .Q(counter_37_));
DFFPOSX1 DFFPOSX1_380 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__13_), .Q(bus_sync_axi_bus_reg_data1_13_));
DFFPOSX1 DFFPOSX1_381 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__14_), .Q(bus_sync_axi_bus_reg_data1_14_));
DFFPOSX1 DFFPOSX1_382 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__15_), .Q(bus_sync_axi_bus_reg_data1_15_));
DFFPOSX1 DFFPOSX1_383 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__16_), .Q(bus_sync_axi_bus_reg_data1_16_));
DFFPOSX1 DFFPOSX1_384 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__17_), .Q(bus_sync_axi_bus_reg_data1_17_));
DFFPOSX1 DFFPOSX1_385 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__18_), .Q(bus_sync_axi_bus_reg_data1_18_));
DFFPOSX1 DFFPOSX1_386 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__19_), .Q(bus_sync_axi_bus_reg_data1_19_));
DFFPOSX1 DFFPOSX1_387 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__20_), .Q(bus_sync_axi_bus_reg_data1_20_));
DFFPOSX1 DFFPOSX1_388 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__21_), .Q(bus_sync_axi_bus_reg_data1_21_));
DFFPOSX1 DFFPOSX1_389 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__22_), .Q(bus_sync_axi_bus_reg_data1_22_));
DFFPOSX1 DFFPOSX1_39 ( .CLK(SCLK), .D(_0counter_65_0__38_), .Q(counter_38_));
DFFPOSX1 DFFPOSX1_390 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__23_), .Q(bus_sync_axi_bus_reg_data1_23_));
DFFPOSX1 DFFPOSX1_391 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__24_), .Q(bus_sync_axi_bus_reg_data1_24_));
DFFPOSX1 DFFPOSX1_392 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__25_), .Q(bus_sync_axi_bus_reg_data1_25_));
DFFPOSX1 DFFPOSX1_393 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__26_), .Q(bus_sync_axi_bus_reg_data1_26_));
DFFPOSX1 DFFPOSX1_394 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__27_), .Q(bus_sync_axi_bus_reg_data1_27_));
DFFPOSX1 DFFPOSX1_395 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__28_), .Q(bus_sync_axi_bus_reg_data1_28_));
DFFPOSX1 DFFPOSX1_396 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__29_), .Q(bus_sync_axi_bus_reg_data1_29_));
DFFPOSX1 DFFPOSX1_397 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__30_), .Q(bus_sync_axi_bus_reg_data1_30_));
DFFPOSX1 DFFPOSX1_398 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__31_), .Q(bus_sync_axi_bus_reg_data1_31_));
DFFPOSX1 DFFPOSX1_399 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__32_), .Q(bus_sync_axi_bus_reg_data1_32_));
DFFPOSX1 DFFPOSX1_4 ( .CLK(SCLK), .D(_0counter_65_0__3_), .Q(counter_3_));
DFFPOSX1 DFFPOSX1_40 ( .CLK(SCLK), .D(_0counter_65_0__39_), .Q(counter_39_));
DFFPOSX1 DFFPOSX1_400 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__33_), .Q(bus_sync_axi_bus_reg_data1_33_));
DFFPOSX1 DFFPOSX1_401 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__34_), .Q(bus_sync_axi_bus_reg_data1_34_));
DFFPOSX1 DFFPOSX1_402 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__35_), .Q(bus_sync_axi_bus_reg_data1_35_));
DFFPOSX1 DFFPOSX1_403 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__36_), .Q(bus_sync_axi_bus_reg_data1_36_));
DFFPOSX1 DFFPOSX1_404 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__37_), .Q(bus_sync_axi_bus_reg_data1_37_));
DFFPOSX1 DFFPOSX1_405 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__38_), .Q(bus_sync_axi_bus_reg_data1_38_));
DFFPOSX1 DFFPOSX1_406 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__39_), .Q(bus_sync_axi_bus_reg_data1_39_));
DFFPOSX1 DFFPOSX1_407 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__40_), .Q(bus_sync_axi_bus_reg_data1_40_));
DFFPOSX1 DFFPOSX1_408 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__41_), .Q(bus_sync_axi_bus_reg_data1_41_));
DFFPOSX1 DFFPOSX1_409 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__42_), .Q(bus_sync_axi_bus_reg_data1_42_));
DFFPOSX1 DFFPOSX1_41 ( .CLK(SCLK), .D(_0counter_65_0__40_), .Q(counter_40_));
DFFPOSX1 DFFPOSX1_410 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__43_), .Q(bus_sync_axi_bus_reg_data1_43_));
DFFPOSX1 DFFPOSX1_411 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__44_), .Q(bus_sync_axi_bus_reg_data1_44_));
DFFPOSX1 DFFPOSX1_412 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__45_), .Q(bus_sync_axi_bus_reg_data1_45_));
DFFPOSX1 DFFPOSX1_413 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__46_), .Q(bus_sync_axi_bus_reg_data1_46_));
DFFPOSX1 DFFPOSX1_414 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__47_), .Q(bus_sync_axi_bus_reg_data1_47_));
DFFPOSX1 DFFPOSX1_415 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__48_), .Q(bus_sync_axi_bus_reg_data1_48_));
DFFPOSX1 DFFPOSX1_416 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__49_), .Q(bus_sync_axi_bus_reg_data1_49_));
DFFPOSX1 DFFPOSX1_417 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__50_), .Q(bus_sync_axi_bus_reg_data1_50_));
DFFPOSX1 DFFPOSX1_418 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__51_), .Q(bus_sync_axi_bus_reg_data1_51_));
DFFPOSX1 DFFPOSX1_419 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__52_), .Q(bus_sync_axi_bus_reg_data1_52_));
DFFPOSX1 DFFPOSX1_42 ( .CLK(SCLK), .D(_0counter_65_0__41_), .Q(counter_41_));
DFFPOSX1 DFFPOSX1_420 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__53_), .Q(bus_sync_axi_bus_reg_data1_53_));
DFFPOSX1 DFFPOSX1_421 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__54_), .Q(bus_sync_axi_bus_reg_data1_54_));
DFFPOSX1 DFFPOSX1_422 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__55_), .Q(bus_sync_axi_bus_reg_data1_55_));
DFFPOSX1 DFFPOSX1_423 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__56_), .Q(bus_sync_axi_bus_reg_data1_56_));
DFFPOSX1 DFFPOSX1_424 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__57_), .Q(bus_sync_axi_bus_reg_data1_57_));
DFFPOSX1 DFFPOSX1_425 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__58_), .Q(bus_sync_axi_bus_reg_data1_58_));
DFFPOSX1 DFFPOSX1_426 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__59_), .Q(bus_sync_axi_bus_reg_data1_59_));
DFFPOSX1 DFFPOSX1_427 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__60_), .Q(bus_sync_axi_bus_reg_data1_60_));
DFFPOSX1 DFFPOSX1_428 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__61_), .Q(bus_sync_axi_bus_reg_data1_61_));
DFFPOSX1 DFFPOSX1_429 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__62_), .Q(bus_sync_axi_bus_reg_data1_62_));
DFFPOSX1 DFFPOSX1_43 ( .CLK(SCLK), .D(_0counter_65_0__42_), .Q(counter_42_));
DFFPOSX1 DFFPOSX1_430 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__63_), .Q(bus_sync_axi_bus_reg_data1_63_));
DFFPOSX1 DFFPOSX1_431 ( .CLK(bus_sync_axi_bus_NCLK2), .D(bus_sync_axi_bus__0ECLK1_0_0_), .Q(bus_sync_axi_bus_ECLK1));
DFFPOSX1 DFFPOSX1_432 ( .CLK(bus_sync_axi_bus_NCLK2), .D(bus_sync_axi_bus__0EECLK1_0_0_), .Q(bus_sync_axi_bus_EECLK1));
DFFPOSX1 DFFPOSX1_433 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__0_), .Q(bus_sync_rdata_data_out_0_));
DFFPOSX1 DFFPOSX1_434 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__1_), .Q(bus_sync_rdata_data_out_1_));
DFFPOSX1 DFFPOSX1_435 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__2_), .Q(bus_sync_rdata_data_out_2_));
DFFPOSX1 DFFPOSX1_436 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__3_), .Q(bus_sync_rdata_data_out_3_));
DFFPOSX1 DFFPOSX1_437 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__4_), .Q(bus_sync_rdata_data_out_4_));
DFFPOSX1 DFFPOSX1_438 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__5_), .Q(bus_sync_rdata_data_out_5_));
DFFPOSX1 DFFPOSX1_439 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__6_), .Q(bus_sync_rdata_data_out_6_));
DFFPOSX1 DFFPOSX1_44 ( .CLK(SCLK), .D(_0counter_65_0__43_), .Q(counter_43_));
DFFPOSX1 DFFPOSX1_440 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__7_), .Q(bus_sync_rdata_data_out_7_));
DFFPOSX1 DFFPOSX1_441 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__8_), .Q(bus_sync_rdata_data_out_8_));
DFFPOSX1 DFFPOSX1_442 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__9_), .Q(bus_sync_rdata_data_out_9_));
DFFPOSX1 DFFPOSX1_443 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__10_), .Q(bus_sync_rdata_data_out_10_));
DFFPOSX1 DFFPOSX1_444 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__11_), .Q(bus_sync_rdata_data_out_11_));
DFFPOSX1 DFFPOSX1_445 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__12_), .Q(bus_sync_rdata_data_out_12_));
DFFPOSX1 DFFPOSX1_446 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__13_), .Q(bus_sync_rdata_data_out_13_));
DFFPOSX1 DFFPOSX1_447 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__14_), .Q(bus_sync_rdata_data_out_14_));
DFFPOSX1 DFFPOSX1_448 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__15_), .Q(bus_sync_rdata_data_out_15_));
DFFPOSX1 DFFPOSX1_449 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__16_), .Q(bus_sync_rdata_data_out_16_));
DFFPOSX1 DFFPOSX1_45 ( .CLK(SCLK), .D(_0counter_65_0__44_), .Q(counter_44_));
DFFPOSX1 DFFPOSX1_450 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__17_), .Q(bus_sync_rdata_data_out_17_));
DFFPOSX1 DFFPOSX1_451 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__18_), .Q(bus_sync_rdata_data_out_18_));
DFFPOSX1 DFFPOSX1_452 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__19_), .Q(bus_sync_rdata_data_out_19_));
DFFPOSX1 DFFPOSX1_453 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__20_), .Q(bus_sync_rdata_data_out_20_));
DFFPOSX1 DFFPOSX1_454 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__21_), .Q(bus_sync_rdata_data_out_21_));
DFFPOSX1 DFFPOSX1_455 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__22_), .Q(bus_sync_rdata_data_out_22_));
DFFPOSX1 DFFPOSX1_456 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__23_), .Q(bus_sync_rdata_data_out_23_));
DFFPOSX1 DFFPOSX1_457 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__24_), .Q(bus_sync_rdata_data_out_24_));
DFFPOSX1 DFFPOSX1_458 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__25_), .Q(bus_sync_rdata_data_out_25_));
DFFPOSX1 DFFPOSX1_459 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__26_), .Q(bus_sync_rdata_data_out_26_));
DFFPOSX1 DFFPOSX1_46 ( .CLK(SCLK), .D(_0counter_65_0__45_), .Q(counter_45_));
DFFPOSX1 DFFPOSX1_460 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__27_), .Q(bus_sync_rdata_data_out_27_));
DFFPOSX1 DFFPOSX1_461 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__28_), .Q(bus_sync_rdata_data_out_28_));
DFFPOSX1 DFFPOSX1_462 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__29_), .Q(bus_sync_rdata_data_out_29_));
DFFPOSX1 DFFPOSX1_463 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__30_), .Q(bus_sync_rdata_data_out_30_));
DFFPOSX1 DFFPOSX1_464 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__31_), .Q(bus_sync_rdata_data_out_31_));
DFFPOSX1 DFFPOSX1_465 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__0_), .Q(bus_sync_rdata_reg_data1_0_));
DFFPOSX1 DFFPOSX1_466 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__1_), .Q(bus_sync_rdata_reg_data1_1_));
DFFPOSX1 DFFPOSX1_467 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__2_), .Q(bus_sync_rdata_reg_data1_2_));
DFFPOSX1 DFFPOSX1_468 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__3_), .Q(bus_sync_rdata_reg_data1_3_));
DFFPOSX1 DFFPOSX1_469 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__4_), .Q(bus_sync_rdata_reg_data1_4_));
DFFPOSX1 DFFPOSX1_47 ( .CLK(SCLK), .D(_0counter_65_0__46_), .Q(counter_46_));
DFFPOSX1 DFFPOSX1_470 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__5_), .Q(bus_sync_rdata_reg_data1_5_));
DFFPOSX1 DFFPOSX1_471 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__6_), .Q(bus_sync_rdata_reg_data1_6_));
DFFPOSX1 DFFPOSX1_472 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__7_), .Q(bus_sync_rdata_reg_data1_7_));
DFFPOSX1 DFFPOSX1_473 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__8_), .Q(bus_sync_rdata_reg_data1_8_));
DFFPOSX1 DFFPOSX1_474 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__9_), .Q(bus_sync_rdata_reg_data1_9_));
DFFPOSX1 DFFPOSX1_475 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__10_), .Q(bus_sync_rdata_reg_data1_10_));
DFFPOSX1 DFFPOSX1_476 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__11_), .Q(bus_sync_rdata_reg_data1_11_));
DFFPOSX1 DFFPOSX1_477 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__12_), .Q(bus_sync_rdata_reg_data1_12_));
DFFPOSX1 DFFPOSX1_478 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__13_), .Q(bus_sync_rdata_reg_data1_13_));
DFFPOSX1 DFFPOSX1_479 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__14_), .Q(bus_sync_rdata_reg_data1_14_));
DFFPOSX1 DFFPOSX1_48 ( .CLK(SCLK), .D(_0counter_65_0__47_), .Q(counter_47_));
DFFPOSX1 DFFPOSX1_480 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__15_), .Q(bus_sync_rdata_reg_data1_15_));
DFFPOSX1 DFFPOSX1_481 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__16_), .Q(bus_sync_rdata_reg_data1_16_));
DFFPOSX1 DFFPOSX1_482 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__17_), .Q(bus_sync_rdata_reg_data1_17_));
DFFPOSX1 DFFPOSX1_483 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__18_), .Q(bus_sync_rdata_reg_data1_18_));
DFFPOSX1 DFFPOSX1_484 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__19_), .Q(bus_sync_rdata_reg_data1_19_));
DFFPOSX1 DFFPOSX1_485 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__20_), .Q(bus_sync_rdata_reg_data1_20_));
DFFPOSX1 DFFPOSX1_486 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__21_), .Q(bus_sync_rdata_reg_data1_21_));
DFFPOSX1 DFFPOSX1_487 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__22_), .Q(bus_sync_rdata_reg_data1_22_));
DFFPOSX1 DFFPOSX1_488 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__23_), .Q(bus_sync_rdata_reg_data1_23_));
DFFPOSX1 DFFPOSX1_489 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__24_), .Q(bus_sync_rdata_reg_data1_24_));
DFFPOSX1 DFFPOSX1_49 ( .CLK(SCLK), .D(_0counter_65_0__48_), .Q(counter_48_));
DFFPOSX1 DFFPOSX1_490 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__25_), .Q(bus_sync_rdata_reg_data1_25_));
DFFPOSX1 DFFPOSX1_491 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__26_), .Q(bus_sync_rdata_reg_data1_26_));
DFFPOSX1 DFFPOSX1_492 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__27_), .Q(bus_sync_rdata_reg_data1_27_));
DFFPOSX1 DFFPOSX1_493 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__28_), .Q(bus_sync_rdata_reg_data1_28_));
DFFPOSX1 DFFPOSX1_494 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__29_), .Q(bus_sync_rdata_reg_data1_29_));
DFFPOSX1 DFFPOSX1_495 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__30_), .Q(bus_sync_rdata_reg_data1_30_));
DFFPOSX1 DFFPOSX1_496 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__31_), .Q(bus_sync_rdata_reg_data1_31_));
DFFPOSX1 DFFPOSX1_497 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__0_), .Q(bus_sync_rdata_reg_data2_0_));
DFFPOSX1 DFFPOSX1_498 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__1_), .Q(bus_sync_rdata_reg_data2_1_));
DFFPOSX1 DFFPOSX1_499 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__2_), .Q(bus_sync_rdata_reg_data2_2_));
DFFPOSX1 DFFPOSX1_5 ( .CLK(SCLK), .D(_0counter_65_0__4_), .Q(counter_4_));
DFFPOSX1 DFFPOSX1_50 ( .CLK(SCLK), .D(_0counter_65_0__49_), .Q(counter_49_));
DFFPOSX1 DFFPOSX1_500 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__3_), .Q(bus_sync_rdata_reg_data2_3_));
DFFPOSX1 DFFPOSX1_501 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__4_), .Q(bus_sync_rdata_reg_data2_4_));
DFFPOSX1 DFFPOSX1_502 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__5_), .Q(bus_sync_rdata_reg_data2_5_));
DFFPOSX1 DFFPOSX1_503 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__6_), .Q(bus_sync_rdata_reg_data2_6_));
DFFPOSX1 DFFPOSX1_504 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__7_), .Q(bus_sync_rdata_reg_data2_7_));
DFFPOSX1 DFFPOSX1_505 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__8_), .Q(bus_sync_rdata_reg_data2_8_));
DFFPOSX1 DFFPOSX1_506 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__9_), .Q(bus_sync_rdata_reg_data2_9_));
DFFPOSX1 DFFPOSX1_507 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__10_), .Q(bus_sync_rdata_reg_data2_10_));
DFFPOSX1 DFFPOSX1_508 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__11_), .Q(bus_sync_rdata_reg_data2_11_));
DFFPOSX1 DFFPOSX1_509 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__12_), .Q(bus_sync_rdata_reg_data2_12_));
DFFPOSX1 DFFPOSX1_51 ( .CLK(SCLK), .D(_0counter_65_0__50_), .Q(counter_50_));
DFFPOSX1 DFFPOSX1_510 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__13_), .Q(bus_sync_rdata_reg_data2_13_));
DFFPOSX1 DFFPOSX1_511 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__14_), .Q(bus_sync_rdata_reg_data2_14_));
DFFPOSX1 DFFPOSX1_512 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__15_), .Q(bus_sync_rdata_reg_data2_15_));
DFFPOSX1 DFFPOSX1_513 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__16_), .Q(bus_sync_rdata_reg_data2_16_));
DFFPOSX1 DFFPOSX1_514 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__17_), .Q(bus_sync_rdata_reg_data2_17_));
DFFPOSX1 DFFPOSX1_515 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__18_), .Q(bus_sync_rdata_reg_data2_18_));
DFFPOSX1 DFFPOSX1_516 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__19_), .Q(bus_sync_rdata_reg_data2_19_));
DFFPOSX1 DFFPOSX1_517 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__20_), .Q(bus_sync_rdata_reg_data2_20_));
DFFPOSX1 DFFPOSX1_518 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__21_), .Q(bus_sync_rdata_reg_data2_21_));
DFFPOSX1 DFFPOSX1_519 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__22_), .Q(bus_sync_rdata_reg_data2_22_));
DFFPOSX1 DFFPOSX1_52 ( .CLK(SCLK), .D(_0counter_65_0__51_), .Q(counter_51_));
DFFPOSX1 DFFPOSX1_520 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__23_), .Q(bus_sync_rdata_reg_data2_23_));
DFFPOSX1 DFFPOSX1_521 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__24_), .Q(bus_sync_rdata_reg_data2_24_));
DFFPOSX1 DFFPOSX1_522 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__25_), .Q(bus_sync_rdata_reg_data2_25_));
DFFPOSX1 DFFPOSX1_523 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__26_), .Q(bus_sync_rdata_reg_data2_26_));
DFFPOSX1 DFFPOSX1_524 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__27_), .Q(bus_sync_rdata_reg_data2_27_));
DFFPOSX1 DFFPOSX1_525 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__28_), .Q(bus_sync_rdata_reg_data2_28_));
DFFPOSX1 DFFPOSX1_526 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__29_), .Q(bus_sync_rdata_reg_data2_29_));
DFFPOSX1 DFFPOSX1_527 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__30_), .Q(bus_sync_rdata_reg_data2_30_));
DFFPOSX1 DFFPOSX1_528 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__31_), .Q(bus_sync_rdata_reg_data2_31_));
DFFPOSX1 DFFPOSX1_529 ( .CLK(bus_sync_rdata_NCLK1), .D(bus_sync_rdata__0EECLK2_0_0_), .Q(bus_sync_rdata_EECLK2));
DFFPOSX1 DFFPOSX1_53 ( .CLK(SCLK), .D(_0counter_65_0__52_), .Q(counter_52_));
DFFPOSX1 DFFPOSX1_530 ( .CLK(bus_sync_rdata_NCLK1), .D(bus_sync_rdata__0ECLK2_0_0_), .Q(bus_sync_rdata_ECLK2));
DFFPOSX1 DFFPOSX1_531 ( .CLK(CLK), .D(bus_sync_state_machine__0reg_data2_3_0__0_), .Q(bus_sync_state_machine_reg_data2_0_));
DFFPOSX1 DFFPOSX1_532 ( .CLK(CLK), .D(bus_sync_state_machine__0reg_data2_3_0__1_), .Q(bus_sync_state_machine_reg_data2_1_));
DFFPOSX1 DFFPOSX1_533 ( .CLK(CLK), .D(bus_sync_state_machine__0reg_data2_3_0__2_), .Q(bus_sync_state_machine_reg_data2_2_));
DFFPOSX1 DFFPOSX1_534 ( .CLK(CLK), .D(bus_sync_state_machine__0reg_data2_3_0__3_), .Q(bus_sync_state_machine_reg_data2_3_));
DFFPOSX1 DFFPOSX1_535 ( .CLK(CLK), .D(bus_sync_state_machine__0reg_data3_3_0__0_), .Q(fini_spi_clk));
DFFPOSX1 DFFPOSX1_536 ( .CLK(CLK), .D(bus_sync_state_machine__0reg_data3_3_0__1_), .Q(re_clk));
DFFPOSX1 DFFPOSX1_537 ( .CLK(CLK), .D(bus_sync_state_machine__0reg_data3_3_0__2_), .Q(we_clk));
DFFPOSX1 DFFPOSX1_538 ( .CLK(CLK), .D(bus_sync_state_machine__0reg_data3_3_0__3_), .Q(PICORV_RST));
DFFPOSX1 DFFPOSX1_539 ( .CLK(SCLK), .D(bus_sync_state_machine__0reg_data1_3_0__0_), .Q(bus_sync_state_machine_reg_data1_0_));
DFFPOSX1 DFFPOSX1_54 ( .CLK(SCLK), .D(_0counter_65_0__53_), .Q(counter_53_));
DFFPOSX1 DFFPOSX1_540 ( .CLK(SCLK), .D(bus_sync_state_machine__0reg_data1_3_0__1_), .Q(bus_sync_state_machine_reg_data1_1_));
DFFPOSX1 DFFPOSX1_541 ( .CLK(SCLK), .D(bus_sync_state_machine__0reg_data1_3_0__2_), .Q(bus_sync_state_machine_reg_data1_2_));
DFFPOSX1 DFFPOSX1_542 ( .CLK(SCLK), .D(bus_sync_state_machine__0reg_data1_3_0__3_), .Q(bus_sync_state_machine_reg_data1_3_));
DFFPOSX1 DFFPOSX1_543 ( .CLK(bus_sync_state_machine_NCLK2), .D(bus_sync_state_machine__0ECLK1_0_0_), .Q(bus_sync_state_machine_ECLK1));
DFFPOSX1 DFFPOSX1_544 ( .CLK(bus_sync_state_machine_NCLK2), .D(bus_sync_state_machine__0EECLK1_0_0_), .Q(bus_sync_state_machine_EECLK1));
DFFPOSX1 DFFPOSX1_545 ( .CLK(SCLK), .D(bus_sync_status__0reg_data3_2_0__0_), .Q(bus_sync_status_data_out_0_));
DFFPOSX1 DFFPOSX1_546 ( .CLK(SCLK), .D(bus_sync_status__0reg_data3_2_0__1_), .Q(bus_sync_status_data_out_1_));
DFFPOSX1 DFFPOSX1_547 ( .CLK(SCLK), .D(bus_sync_status__0reg_data3_2_0__2_), .Q(bus_sync_status_data_out_2_));
DFFPOSX1 DFFPOSX1_548 ( .CLK(CLK), .D(bus_sync_status__0reg_data1_2_0__0_), .Q(bus_sync_status_reg_data1_0_));
DFFPOSX1 DFFPOSX1_549 ( .CLK(CLK), .D(bus_sync_status__0reg_data1_2_0__1_), .Q(bus_sync_status_reg_data1_1_));
DFFPOSX1 DFFPOSX1_55 ( .CLK(SCLK), .D(_0counter_65_0__54_), .Q(counter_54_));
DFFPOSX1 DFFPOSX1_550 ( .CLK(CLK), .D(bus_sync_status__0reg_data1_2_0__2_), .Q(bus_sync_status_reg_data1_2_));
DFFPOSX1 DFFPOSX1_551 ( .CLK(CLK), .D(bus_sync_status__0reg_data2_2_0__0_), .Q(bus_sync_status_reg_data2_0_));
DFFPOSX1 DFFPOSX1_552 ( .CLK(CLK), .D(bus_sync_status__0reg_data2_2_0__1_), .Q(bus_sync_status_reg_data2_1_));
DFFPOSX1 DFFPOSX1_553 ( .CLK(CLK), .D(bus_sync_status__0reg_data2_2_0__2_), .Q(bus_sync_status_reg_data2_2_));
DFFPOSX1 DFFPOSX1_554 ( .CLK(bus_sync_status_NCLK1), .D(bus_sync_status__0EECLK2_0_0_), .Q(bus_sync_status_EECLK2));
DFFPOSX1 DFFPOSX1_555 ( .CLK(bus_sync_status_NCLK1), .D(bus_sync_status__0ECLK2_0_0_), .Q(bus_sync_status_ECLK2));
DFFPOSX1 DFFPOSX1_56 ( .CLK(SCLK), .D(_0counter_65_0__55_), .Q(counter_55_));
DFFPOSX1 DFFPOSX1_57 ( .CLK(SCLK), .D(_0counter_65_0__56_), .Q(counter_56_));
DFFPOSX1 DFFPOSX1_58 ( .CLK(SCLK), .D(_0counter_65_0__57_), .Q(counter_57_));
DFFPOSX1 DFFPOSX1_59 ( .CLK(SCLK), .D(_0counter_65_0__58_), .Q(counter_58_));
DFFPOSX1 DFFPOSX1_6 ( .CLK(SCLK), .D(_0counter_65_0__5_), .Q(counter_5_));
DFFPOSX1 DFFPOSX1_60 ( .CLK(SCLK), .D(_0counter_65_0__59_), .Q(counter_59_));
DFFPOSX1 DFFPOSX1_61 ( .CLK(SCLK), .D(_0counter_65_0__60_), .Q(counter_60_));
DFFPOSX1 DFFPOSX1_62 ( .CLK(SCLK), .D(_0counter_65_0__61_), .Q(counter_61_));
DFFPOSX1 DFFPOSX1_63 ( .CLK(SCLK), .D(_0counter_65_0__62_), .Q(counter_62_));
DFFPOSX1 DFFPOSX1_64 ( .CLK(SCLK), .D(_0counter_65_0__63_), .Q(counter_63_));
DFFPOSX1 DFFPOSX1_65 ( .CLK(SCLK), .D(_0counter_65_0__64_), .Q(counter_64_));
DFFPOSX1 DFFPOSX1_66 ( .CLK(SCLK), .D(_0counter_65_0__65_), .Q(counter_65_));
DFFPOSX1 DFFPOSX1_67 ( .CLK(SCLK), .D(_0fini_spi_0_0_), .Q(fini_spi));
DFFPOSX1 DFFPOSX1_68 ( .CLK(SCLK), .D(_0bus_cap_31_0__0_), .Q(bus_cap_0_));
DFFPOSX1 DFFPOSX1_69 ( .CLK(SCLK), .D(_0bus_cap_31_0__1_), .Q(bus_cap_1_));
DFFPOSX1 DFFPOSX1_7 ( .CLK(SCLK), .D(_0counter_65_0__6_), .Q(counter_6_));
DFFPOSX1 DFFPOSX1_70 ( .CLK(SCLK), .D(_0bus_cap_31_0__2_), .Q(bus_cap_2_));
DFFPOSX1 DFFPOSX1_71 ( .CLK(SCLK), .D(_0bus_cap_31_0__3_), .Q(bus_cap_3_));
DFFPOSX1 DFFPOSX1_72 ( .CLK(SCLK), .D(_0bus_cap_31_0__4_), .Q(bus_cap_4_));
DFFPOSX1 DFFPOSX1_73 ( .CLK(SCLK), .D(_0bus_cap_31_0__5_), .Q(bus_cap_5_));
DFFPOSX1 DFFPOSX1_74 ( .CLK(SCLK), .D(_0bus_cap_31_0__6_), .Q(bus_cap_6_));
DFFPOSX1 DFFPOSX1_75 ( .CLK(SCLK), .D(_0bus_cap_31_0__7_), .Q(bus_cap_7_));
DFFPOSX1 DFFPOSX1_76 ( .CLK(SCLK), .D(_0bus_cap_31_0__8_), .Q(bus_cap_8_));
DFFPOSX1 DFFPOSX1_77 ( .CLK(SCLK), .D(_0bus_cap_31_0__9_), .Q(bus_cap_9_));
DFFPOSX1 DFFPOSX1_78 ( .CLK(SCLK), .D(_0bus_cap_31_0__10_), .Q(bus_cap_10_));
DFFPOSX1 DFFPOSX1_79 ( .CLK(SCLK), .D(_0bus_cap_31_0__11_), .Q(bus_cap_11_));
DFFPOSX1 DFFPOSX1_8 ( .CLK(SCLK), .D(_0counter_65_0__7_), .Q(counter_7_));
DFFPOSX1 DFFPOSX1_80 ( .CLK(SCLK), .D(_0bus_cap_31_0__12_), .Q(bus_cap_12_));
DFFPOSX1 DFFPOSX1_81 ( .CLK(SCLK), .D(_0bus_cap_31_0__13_), .Q(bus_cap_13_));
DFFPOSX1 DFFPOSX1_82 ( .CLK(SCLK), .D(_0bus_cap_31_0__14_), .Q(bus_cap_14_));
DFFPOSX1 DFFPOSX1_83 ( .CLK(SCLK), .D(_0bus_cap_31_0__15_), .Q(bus_cap_15_));
DFFPOSX1 DFFPOSX1_84 ( .CLK(SCLK), .D(_0bus_cap_31_0__16_), .Q(bus_cap_16_));
DFFPOSX1 DFFPOSX1_85 ( .CLK(SCLK), .D(_0bus_cap_31_0__17_), .Q(bus_cap_17_));
DFFPOSX1 DFFPOSX1_86 ( .CLK(SCLK), .D(_0bus_cap_31_0__18_), .Q(bus_cap_18_));
DFFPOSX1 DFFPOSX1_87 ( .CLK(SCLK), .D(_0bus_cap_31_0__19_), .Q(bus_cap_19_));
DFFPOSX1 DFFPOSX1_88 ( .CLK(SCLK), .D(_0bus_cap_31_0__20_), .Q(bus_cap_20_));
DFFPOSX1 DFFPOSX1_89 ( .CLK(SCLK), .D(_0bus_cap_31_0__21_), .Q(bus_cap_21_));
DFFPOSX1 DFFPOSX1_9 ( .CLK(SCLK), .D(_0counter_65_0__8_), .Q(counter_8_));
DFFPOSX1 DFFPOSX1_90 ( .CLK(SCLK), .D(_0bus_cap_31_0__22_), .Q(bus_cap_22_));
DFFPOSX1 DFFPOSX1_91 ( .CLK(SCLK), .D(_0bus_cap_31_0__23_), .Q(bus_cap_23_));
DFFPOSX1 DFFPOSX1_92 ( .CLK(SCLK), .D(_0bus_cap_31_0__24_), .Q(bus_cap_24_));
DFFPOSX1 DFFPOSX1_93 ( .CLK(SCLK), .D(_0bus_cap_31_0__25_), .Q(bus_cap_25_));
DFFPOSX1 DFFPOSX1_94 ( .CLK(SCLK), .D(_0bus_cap_31_0__26_), .Q(bus_cap_26_));
DFFPOSX1 DFFPOSX1_95 ( .CLK(SCLK), .D(_0bus_cap_31_0__27_), .Q(bus_cap_27_));
DFFPOSX1 DFFPOSX1_96 ( .CLK(SCLK), .D(_0bus_cap_31_0__28_), .Q(bus_cap_28_));
DFFPOSX1 DFFPOSX1_97 ( .CLK(SCLK), .D(_0bus_cap_31_0__29_), .Q(bus_cap_29_));
DFFPOSX1 DFFPOSX1_98 ( .CLK(SCLK), .D(_0bus_cap_31_0__30_), .Q(bus_cap_30_));
DFFPOSX1 DFFPOSX1_99 ( .CLK(SCLK), .D(_0bus_cap_31_0__31_), .Q(DOUT));
INVX1 INVX1_1 ( .A(state_7_), .Y(_abc_4169_new_n558_));
INVX1 INVX1_10 ( .A(_abc_4169_new_n601_), .Y(_abc_4169_new_n602_));
INVX1 INVX1_100 ( .A(WDATA_15_), .Y(_abc_4169_new_n983_));
INVX1 INVX1_101 ( .A(WDATA_16_), .Y(_abc_4169_new_n986_));
INVX1 INVX1_102 ( .A(WDATA_17_), .Y(_abc_4169_new_n989_));
INVX1 INVX1_103 ( .A(WDATA_18_), .Y(_abc_4169_new_n992_));
INVX1 INVX1_104 ( .A(WDATA_19_), .Y(_abc_4169_new_n995_));
INVX1 INVX1_105 ( .A(WDATA_20_), .Y(_abc_4169_new_n998_));
INVX1 INVX1_106 ( .A(WDATA_21_), .Y(_abc_4169_new_n1001_));
INVX1 INVX1_107 ( .A(WDATA_22_), .Y(_abc_4169_new_n1004_));
INVX1 INVX1_108 ( .A(WDATA_23_), .Y(_abc_4169_new_n1007_));
INVX1 INVX1_109 ( .A(WDATA_24_), .Y(_abc_4169_new_n1010_));
INVX1 INVX1_11 ( .A(re), .Y(_abc_4169_new_n604_));
INVX1 INVX1_110 ( .A(WDATA_25_), .Y(_abc_4169_new_n1013_));
INVX1 INVX1_111 ( .A(WDATA_26_), .Y(_abc_4169_new_n1016_));
INVX1 INVX1_112 ( .A(WDATA_27_), .Y(_abc_4169_new_n1019_));
INVX1 INVX1_113 ( .A(WDATA_28_), .Y(_abc_4169_new_n1022_));
INVX1 INVX1_114 ( .A(WDATA_29_), .Y(_abc_4169_new_n1025_));
INVX1 INVX1_115 ( .A(WDATA_30_), .Y(_abc_4169_new_n1028_));
INVX1 INVX1_116 ( .A(WDATA_31_), .Y(_abc_4169_new_n1031_));
INVX1 INVX1_117 ( .A(A_ADDR_0_), .Y(_abc_4169_new_n1034_));
INVX1 INVX1_118 ( .A(counter_33_), .Y(_abc_4169_new_n1035_));
INVX1 INVX1_119 ( .A(A_ADDR_1_), .Y(_abc_4169_new_n1040_));
INVX1 INVX1_12 ( .A(we), .Y(_abc_4169_new_n605_));
INVX1 INVX1_120 ( .A(A_ADDR_2_), .Y(_abc_4169_new_n1043_));
INVX1 INVX1_121 ( .A(A_ADDR_3_), .Y(_abc_4169_new_n1046_));
INVX1 INVX1_122 ( .A(A_ADDR_4_), .Y(_abc_4169_new_n1049_));
INVX1 INVX1_123 ( .A(A_ADDR_5_), .Y(_abc_4169_new_n1052_));
INVX1 INVX1_124 ( .A(A_ADDR_6_), .Y(_abc_4169_new_n1055_));
INVX1 INVX1_125 ( .A(A_ADDR_7_), .Y(_abc_4169_new_n1058_));
INVX1 INVX1_126 ( .A(A_ADDR_8_), .Y(_abc_4169_new_n1061_));
INVX1 INVX1_127 ( .A(A_ADDR_9_), .Y(_abc_4169_new_n1064_));
INVX1 INVX1_128 ( .A(A_ADDR_10_), .Y(_abc_4169_new_n1067_));
INVX1 INVX1_129 ( .A(A_ADDR_11_), .Y(_abc_4169_new_n1070_));
INVX1 INVX1_13 ( .A(counter_2_), .Y(_abc_4169_new_n611_));
INVX1 INVX1_130 ( .A(A_ADDR_12_), .Y(_abc_4169_new_n1073_));
INVX1 INVX1_131 ( .A(A_ADDR_13_), .Y(_abc_4169_new_n1076_));
INVX1 INVX1_132 ( .A(A_ADDR_14_), .Y(_abc_4169_new_n1079_));
INVX1 INVX1_133 ( .A(A_ADDR_15_), .Y(_abc_4169_new_n1082_));
INVX1 INVX1_134 ( .A(A_ADDR_16_), .Y(_abc_4169_new_n1085_));
INVX1 INVX1_135 ( .A(A_ADDR_17_), .Y(_abc_4169_new_n1088_));
INVX1 INVX1_136 ( .A(A_ADDR_18_), .Y(_abc_4169_new_n1091_));
INVX1 INVX1_137 ( .A(A_ADDR_19_), .Y(_abc_4169_new_n1094_));
INVX1 INVX1_138 ( .A(A_ADDR_20_), .Y(_abc_4169_new_n1097_));
INVX1 INVX1_139 ( .A(A_ADDR_21_), .Y(_abc_4169_new_n1100_));
INVX1 INVX1_14 ( .A(counter_3_), .Y(_abc_4169_new_n612_));
INVX1 INVX1_140 ( .A(A_ADDR_22_), .Y(_abc_4169_new_n1103_));
INVX1 INVX1_141 ( .A(A_ADDR_23_), .Y(_abc_4169_new_n1106_));
INVX1 INVX1_142 ( .A(A_ADDR_24_), .Y(_abc_4169_new_n1109_));
INVX1 INVX1_143 ( .A(A_ADDR_25_), .Y(_abc_4169_new_n1112_));
INVX1 INVX1_144 ( .A(A_ADDR_26_), .Y(_abc_4169_new_n1115_));
INVX1 INVX1_145 ( .A(A_ADDR_27_), .Y(_abc_4169_new_n1118_));
INVX1 INVX1_146 ( .A(A_ADDR_28_), .Y(_abc_4169_new_n1121_));
INVX1 INVX1_147 ( .A(A_ADDR_29_), .Y(_abc_4169_new_n1124_));
INVX1 INVX1_148 ( .A(A_ADDR_30_), .Y(_abc_4169_new_n1127_));
INVX1 INVX1_149 ( .A(A_ADDR_31_), .Y(_abc_4169_new_n1130_));
INVX1 INVX1_15 ( .A(counter_6_), .Y(_abc_4169_new_n627_));
INVX1 INVX1_150 ( .A(sft_reg_0_), .Y(_abc_4169_new_n1133_));
INVX1 INVX1_151 ( .A(sft_reg_2_), .Y(_abc_4169_new_n1138_));
INVX1 INVX1_152 ( .A(sft_reg_4_), .Y(_abc_4169_new_n1143_));
INVX1 INVX1_153 ( .A(sft_reg_6_), .Y(_abc_4169_new_n1148_));
INVX1 INVX1_154 ( .A(sft_reg_8_), .Y(_abc_4169_new_n1153_));
INVX1 INVX1_155 ( .A(sft_reg_10_), .Y(_abc_4169_new_n1158_));
INVX1 INVX1_156 ( .A(sft_reg_12_), .Y(_abc_4169_new_n1163_));
INVX1 INVX1_157 ( .A(sft_reg_14_), .Y(_abc_4169_new_n1168_));
INVX1 INVX1_158 ( .A(sft_reg_16_), .Y(_abc_4169_new_n1173_));
INVX1 INVX1_159 ( .A(sft_reg_18_), .Y(_abc_4169_new_n1178_));
INVX1 INVX1_16 ( .A(counter_7_), .Y(_abc_4169_new_n628_));
INVX1 INVX1_160 ( .A(sft_reg_20_), .Y(_abc_4169_new_n1183_));
INVX1 INVX1_161 ( .A(sft_reg_22_), .Y(_abc_4169_new_n1188_));
INVX1 INVX1_162 ( .A(sft_reg_24_), .Y(_abc_4169_new_n1193_));
INVX1 INVX1_163 ( .A(sft_reg_26_), .Y(_abc_4169_new_n1198_));
INVX1 INVX1_164 ( .A(sft_reg_28_), .Y(_abc_4169_new_n1203_));
INVX1 INVX1_165 ( .A(sft_reg_30_), .Y(_abc_4169_new_n1208_));
INVX1 INVX1_166 ( .A(counter_0_), .Y(_abc_4169_new_n1212_));
INVX1 INVX1_167 ( .A(counter_4_), .Y(_abc_4169_new_n1217_));
INVX1 INVX1_168 ( .A(counter_5_), .Y(_abc_4169_new_n1219_));
INVX1 INVX1_169 ( .A(counter_8_), .Y(_abc_4169_new_n1223_));
INVX1 INVX1_17 ( .A(counter_18_), .Y(_abc_4169_new_n635_));
INVX1 INVX1_170 ( .A(counter_9_), .Y(_abc_4169_new_n1225_));
INVX1 INVX1_171 ( .A(counter_10_), .Y(_abc_4169_new_n1227_));
INVX1 INVX1_172 ( .A(counter_11_), .Y(_abc_4169_new_n1229_));
INVX1 INVX1_173 ( .A(counter_12_), .Y(_abc_4169_new_n1231_));
INVX1 INVX1_174 ( .A(counter_13_), .Y(_abc_4169_new_n1233_));
INVX1 INVX1_175 ( .A(counter_14_), .Y(_abc_4169_new_n1235_));
INVX1 INVX1_176 ( .A(counter_15_), .Y(_abc_4169_new_n1237_));
INVX1 INVX1_177 ( .A(counter_16_), .Y(_abc_4169_new_n1239_));
INVX1 INVX1_178 ( .A(counter_17_), .Y(_abc_4169_new_n1241_));
INVX1 INVX1_179 ( .A(counter_20_), .Y(_abc_4169_new_n1245_));
INVX1 INVX1_18 ( .A(counter_19_), .Y(_abc_4169_new_n636_));
INVX1 INVX1_180 ( .A(counter_21_), .Y(_abc_4169_new_n1247_));
INVX1 INVX1_181 ( .A(counter_22_), .Y(_abc_4169_new_n1249_));
INVX1 INVX1_182 ( .A(counter_23_), .Y(_abc_4169_new_n1251_));
INVX1 INVX1_183 ( .A(counter_24_), .Y(_abc_4169_new_n1253_));
INVX1 INVX1_184 ( .A(counter_25_), .Y(_abc_4169_new_n1255_));
INVX1 INVX1_185 ( .A(counter_26_), .Y(_abc_4169_new_n1257_));
INVX1 INVX1_186 ( .A(counter_27_), .Y(_abc_4169_new_n1259_));
INVX1 INVX1_187 ( .A(counter_28_), .Y(_abc_4169_new_n1261_));
INVX1 INVX1_188 ( .A(counter_29_), .Y(_abc_4169_new_n1263_));
INVX1 INVX1_189 ( .A(counter_30_), .Y(_abc_4169_new_n1265_));
INVX1 INVX1_19 ( .A(bus_sync_rdata_data_out_0_), .Y(_abc_4169_new_n644_));
INVX1 INVX1_190 ( .A(counter_31_), .Y(_abc_4169_new_n1267_));
INVX1 INVX1_191 ( .A(counter_32_), .Y(_abc_4169_new_n1269_));
INVX1 INVX1_192 ( .A(counter_34_), .Y(_abc_4169_new_n1272_));
INVX1 INVX1_193 ( .A(counter_35_), .Y(_abc_4169_new_n1274_));
INVX1 INVX1_194 ( .A(counter_36_), .Y(_abc_4169_new_n1276_));
INVX1 INVX1_195 ( .A(counter_37_), .Y(_abc_4169_new_n1278_));
INVX1 INVX1_196 ( .A(counter_38_), .Y(_abc_4169_new_n1280_));
INVX1 INVX1_197 ( .A(counter_39_), .Y(_abc_4169_new_n1282_));
INVX1 INVX1_198 ( .A(counter_40_), .Y(_abc_4169_new_n1284_));
INVX1 INVX1_199 ( .A(counter_41_), .Y(_abc_4169_new_n1286_));
INVX1 INVX1_2 ( .A(RST), .Y(_abc_4169_new_n564_));
INVX1 INVX1_20 ( .A(bus_sync_rdata_data_out_1_), .Y(_abc_4169_new_n654_));
INVX1 INVX1_200 ( .A(counter_42_), .Y(_abc_4169_new_n1288_));
INVX1 INVX1_201 ( .A(counter_43_), .Y(_abc_4169_new_n1290_));
INVX1 INVX1_202 ( .A(counter_44_), .Y(_abc_4169_new_n1292_));
INVX1 INVX1_203 ( .A(counter_45_), .Y(_abc_4169_new_n1294_));
INVX1 INVX1_204 ( .A(counter_46_), .Y(_abc_4169_new_n1296_));
INVX1 INVX1_205 ( .A(counter_47_), .Y(_abc_4169_new_n1298_));
INVX1 INVX1_206 ( .A(counter_48_), .Y(_abc_4169_new_n1300_));
INVX1 INVX1_207 ( .A(counter_49_), .Y(_abc_4169_new_n1302_));
INVX1 INVX1_208 ( .A(counter_50_), .Y(_abc_4169_new_n1304_));
INVX1 INVX1_209 ( .A(counter_51_), .Y(_abc_4169_new_n1306_));
INVX1 INVX1_21 ( .A(bus_sync_rdata_data_out_2_), .Y(_abc_4169_new_n661_));
INVX1 INVX1_210 ( .A(counter_52_), .Y(_abc_4169_new_n1308_));
INVX1 INVX1_211 ( .A(counter_53_), .Y(_abc_4169_new_n1310_));
INVX1 INVX1_212 ( .A(counter_54_), .Y(_abc_4169_new_n1312_));
INVX1 INVX1_213 ( .A(counter_55_), .Y(_abc_4169_new_n1314_));
INVX1 INVX1_214 ( .A(counter_56_), .Y(_abc_4169_new_n1316_));
INVX1 INVX1_215 ( .A(counter_57_), .Y(_abc_4169_new_n1318_));
INVX1 INVX1_216 ( .A(counter_58_), .Y(_abc_4169_new_n1320_));
INVX1 INVX1_217 ( .A(counter_59_), .Y(_abc_4169_new_n1322_));
INVX1 INVX1_218 ( .A(counter_60_), .Y(_abc_4169_new_n1324_));
INVX1 INVX1_219 ( .A(counter_61_), .Y(_abc_4169_new_n1326_));
INVX1 INVX1_22 ( .A(bus_sync_rdata_data_out_3_), .Y(_abc_4169_new_n667_));
INVX1 INVX1_220 ( .A(counter_62_), .Y(_abc_4169_new_n1328_));
INVX1 INVX1_221 ( .A(counter_63_), .Y(_abc_4169_new_n1330_));
INVX1 INVX1_222 ( .A(counter_64_), .Y(_abc_4169_new_n1332_));
INVX1 INVX1_223 ( .A(PICORV_RST_SPI), .Y(_abc_4169_new_n1334_));
INVX1 INVX1_224 ( .A(_abc_4169_new_n606_), .Y(_abc_4169_new_n1335_));
INVX1 INVX1_225 ( .A(_abc_4169_new_n1346_), .Y(_abc_2903_auto_fsm_map_cc_118_implement_pattern_cache_479));
INVX1 INVX1_226 ( .A(_abc_4169_new_n1348_), .Y(_abc_2903_auto_fsm_map_cc_118_implement_pattern_cache_430));
INVX1 INVX1_227 ( .A(RST), .Y(bus_sync_axi_bus__abc_3843_new_n393_));
INVX1 INVX1_228 ( .A(bus_sync_axi_bus_EECLK1), .Y(bus_sync_axi_bus__abc_3843_new_n394_));
INVX1 INVX1_229 ( .A(CLK), .Y(bus_sync_axi_bus_NCLK2));
INVX1 INVX1_23 ( .A(bus_sync_rdata_data_out_4_), .Y(_abc_4169_new_n673_));
INVX1 INVX1_230 ( .A(RST), .Y(bus_sync_rdata__abc_3651_new_n265_));
INVX1 INVX1_231 ( .A(bus_sync_rdata_EECLK2), .Y(bus_sync_rdata__abc_3651_new_n266_));
INVX1 INVX1_232 ( .A(CLK), .Y(bus_sync_rdata_NCLK1));
INVX1 INVX1_233 ( .A(RST), .Y(bus_sync_state_machine__abc_3817_new_n33_));
INVX1 INVX1_234 ( .A(bus_sync_state_machine_EECLK1), .Y(bus_sync_state_machine__abc_3817_new_n34_));
INVX1 INVX1_235 ( .A(CLK), .Y(bus_sync_state_machine_NCLK2));
INVX1 INVX1_236 ( .A(RST), .Y(bus_sync_status__abc_3630_new_n27_));
INVX1 INVX1_237 ( .A(bus_sync_status_EECLK2), .Y(bus_sync_status__abc_3630_new_n28_));
INVX1 INVX1_238 ( .A(CLK), .Y(bus_sync_status_NCLK1));
INVX1 INVX1_24 ( .A(bus_sync_rdata_data_out_5_), .Y(_abc_4169_new_n679_));
INVX1 INVX1_25 ( .A(bus_sync_rdata_data_out_6_), .Y(_abc_4169_new_n685_));
INVX1 INVX1_26 ( .A(bus_sync_rdata_data_out_7_), .Y(_abc_4169_new_n691_));
INVX1 INVX1_27 ( .A(bus_sync_rdata_data_out_8_), .Y(_abc_4169_new_n697_));
INVX1 INVX1_28 ( .A(bus_sync_rdata_data_out_9_), .Y(_abc_4169_new_n703_));
INVX1 INVX1_29 ( .A(bus_sync_rdata_data_out_10_), .Y(_abc_4169_new_n709_));
INVX1 INVX1_3 ( .A(axi_wready), .Y(_abc_4169_new_n565_));
INVX1 INVX1_30 ( .A(bus_sync_rdata_data_out_11_), .Y(_abc_4169_new_n715_));
INVX1 INVX1_31 ( .A(bus_sync_rdata_data_out_12_), .Y(_abc_4169_new_n721_));
INVX1 INVX1_32 ( .A(bus_sync_rdata_data_out_13_), .Y(_abc_4169_new_n727_));
INVX1 INVX1_33 ( .A(bus_sync_rdata_data_out_14_), .Y(_abc_4169_new_n733_));
INVX1 INVX1_34 ( .A(bus_sync_rdata_data_out_15_), .Y(_abc_4169_new_n739_));
INVX1 INVX1_35 ( .A(bus_sync_rdata_data_out_16_), .Y(_abc_4169_new_n745_));
INVX1 INVX1_36 ( .A(bus_sync_rdata_data_out_17_), .Y(_abc_4169_new_n751_));
INVX1 INVX1_37 ( .A(bus_sync_rdata_data_out_18_), .Y(_abc_4169_new_n757_));
INVX1 INVX1_38 ( .A(bus_sync_rdata_data_out_19_), .Y(_abc_4169_new_n763_));
INVX1 INVX1_39 ( .A(bus_sync_rdata_data_out_20_), .Y(_abc_4169_new_n769_));
INVX1 INVX1_4 ( .A(axi_arready), .Y(_abc_4169_new_n578_));
INVX1 INVX1_40 ( .A(bus_sync_rdata_data_out_21_), .Y(_abc_4169_new_n775_));
INVX1 INVX1_41 ( .A(bus_sync_rdata_data_out_22_), .Y(_abc_4169_new_n781_));
INVX1 INVX1_42 ( .A(bus_sync_rdata_data_out_23_), .Y(_abc_4169_new_n787_));
INVX1 INVX1_43 ( .A(bus_sync_rdata_data_out_24_), .Y(_abc_4169_new_n793_));
INVX1 INVX1_44 ( .A(bus_sync_rdata_data_out_25_), .Y(_abc_4169_new_n799_));
INVX1 INVX1_45 ( .A(bus_sync_rdata_data_out_26_), .Y(_abc_4169_new_n805_));
INVX1 INVX1_46 ( .A(bus_sync_rdata_data_out_27_), .Y(_abc_4169_new_n811_));
INVX1 INVX1_47 ( .A(bus_sync_rdata_data_out_28_), .Y(_abc_4169_new_n817_));
INVX1 INVX1_48 ( .A(bus_sync_rdata_data_out_29_), .Y(_abc_4169_new_n823_));
INVX1 INVX1_49 ( .A(bus_sync_rdata_data_out_30_), .Y(_abc_4169_new_n829_));
INVX1 INVX1_5 ( .A(_abc_4169_new_n562_), .Y(_abc_4169_new_n586_));
INVX1 INVX1_50 ( .A(bus_sync_rdata_data_out_31_), .Y(_abc_4169_new_n835_));
INVX1 INVX1_51 ( .A(axi_rready), .Y(_abc_4169_new_n839_));
INVX1 INVX1_52 ( .A(bus_sync_rdata_data_in_0_), .Y(_abc_4169_new_n840_));
INVX1 INVX1_53 ( .A(bus_sync_rdata_data_in_1_), .Y(_abc_4169_new_n843_));
INVX1 INVX1_54 ( .A(bus_sync_rdata_data_in_2_), .Y(_abc_4169_new_n846_));
INVX1 INVX1_55 ( .A(bus_sync_rdata_data_in_3_), .Y(_abc_4169_new_n849_));
INVX1 INVX1_56 ( .A(bus_sync_rdata_data_in_4_), .Y(_abc_4169_new_n852_));
INVX1 INVX1_57 ( .A(bus_sync_rdata_data_in_5_), .Y(_abc_4169_new_n855_));
INVX1 INVX1_58 ( .A(bus_sync_rdata_data_in_6_), .Y(_abc_4169_new_n858_));
INVX1 INVX1_59 ( .A(bus_sync_rdata_data_in_7_), .Y(_abc_4169_new_n861_));
INVX1 INVX1_6 ( .A(fini_spi_clk), .Y(_abc_4169_new_n590_));
INVX1 INVX1_60 ( .A(bus_sync_rdata_data_in_8_), .Y(_abc_4169_new_n864_));
INVX1 INVX1_61 ( .A(bus_sync_rdata_data_in_9_), .Y(_abc_4169_new_n867_));
INVX1 INVX1_62 ( .A(bus_sync_rdata_data_in_10_), .Y(_abc_4169_new_n870_));
INVX1 INVX1_63 ( .A(bus_sync_rdata_data_in_11_), .Y(_abc_4169_new_n873_));
INVX1 INVX1_64 ( .A(bus_sync_rdata_data_in_12_), .Y(_abc_4169_new_n876_));
INVX1 INVX1_65 ( .A(bus_sync_rdata_data_in_13_), .Y(_abc_4169_new_n879_));
INVX1 INVX1_66 ( .A(bus_sync_rdata_data_in_14_), .Y(_abc_4169_new_n882_));
INVX1 INVX1_67 ( .A(bus_sync_rdata_data_in_15_), .Y(_abc_4169_new_n885_));
INVX1 INVX1_68 ( .A(bus_sync_rdata_data_in_16_), .Y(_abc_4169_new_n888_));
INVX1 INVX1_69 ( .A(bus_sync_rdata_data_in_17_), .Y(_abc_4169_new_n891_));
INVX1 INVX1_7 ( .A(axi_awready), .Y(_abc_4169_new_n593_));
INVX1 INVX1_70 ( .A(bus_sync_rdata_data_in_18_), .Y(_abc_4169_new_n894_));
INVX1 INVX1_71 ( .A(bus_sync_rdata_data_in_19_), .Y(_abc_4169_new_n897_));
INVX1 INVX1_72 ( .A(bus_sync_rdata_data_in_20_), .Y(_abc_4169_new_n900_));
INVX1 INVX1_73 ( .A(bus_sync_rdata_data_in_21_), .Y(_abc_4169_new_n903_));
INVX1 INVX1_74 ( .A(bus_sync_rdata_data_in_22_), .Y(_abc_4169_new_n906_));
INVX1 INVX1_75 ( .A(bus_sync_rdata_data_in_23_), .Y(_abc_4169_new_n909_));
INVX1 INVX1_76 ( .A(bus_sync_rdata_data_in_24_), .Y(_abc_4169_new_n912_));
INVX1 INVX1_77 ( .A(bus_sync_rdata_data_in_25_), .Y(_abc_4169_new_n915_));
INVX1 INVX1_78 ( .A(bus_sync_rdata_data_in_26_), .Y(_abc_4169_new_n918_));
INVX1 INVX1_79 ( .A(bus_sync_rdata_data_in_27_), .Y(_abc_4169_new_n921_));
INVX1 INVX1_8 ( .A(counter_1_), .Y(_abc_4169_new_n597_));
INVX1 INVX1_80 ( .A(bus_sync_rdata_data_in_28_), .Y(_abc_4169_new_n924_));
INVX1 INVX1_81 ( .A(bus_sync_rdata_data_in_29_), .Y(_abc_4169_new_n927_));
INVX1 INVX1_82 ( .A(bus_sync_rdata_data_in_30_), .Y(_abc_4169_new_n930_));
INVX1 INVX1_83 ( .A(bus_sync_rdata_data_in_31_), .Y(_abc_4169_new_n933_));
INVX1 INVX1_84 ( .A(WDATA_0_), .Y(_abc_4169_new_n936_));
INVX1 INVX1_85 ( .A(CEB), .Y(_abc_4169_new_n937_));
INVX1 INVX1_86 ( .A(WDATA_1_), .Y(_abc_4169_new_n941_));
INVX1 INVX1_87 ( .A(WDATA_2_), .Y(_abc_4169_new_n944_));
INVX1 INVX1_88 ( .A(WDATA_3_), .Y(_abc_4169_new_n947_));
INVX1 INVX1_89 ( .A(WDATA_4_), .Y(_abc_4169_new_n950_));
INVX1 INVX1_9 ( .A(_abc_4169_new_n599_), .Y(_abc_4169_new_n600_));
INVX1 INVX1_90 ( .A(WDATA_5_), .Y(_abc_4169_new_n953_));
INVX1 INVX1_91 ( .A(WDATA_6_), .Y(_abc_4169_new_n956_));
INVX1 INVX1_92 ( .A(WDATA_7_), .Y(_abc_4169_new_n959_));
INVX1 INVX1_93 ( .A(WDATA_8_), .Y(_abc_4169_new_n962_));
INVX1 INVX1_94 ( .A(WDATA_9_), .Y(_abc_4169_new_n965_));
INVX1 INVX1_95 ( .A(WDATA_10_), .Y(_abc_4169_new_n968_));
INVX1 INVX1_96 ( .A(WDATA_11_), .Y(_abc_4169_new_n971_));
INVX1 INVX1_97 ( .A(WDATA_12_), .Y(_abc_4169_new_n974_));
INVX1 INVX1_98 ( .A(WDATA_13_), .Y(_abc_4169_new_n977_));
INVX1 INVX1_99 ( .A(WDATA_14_), .Y(_abc_4169_new_n980_));
NAND2X1 NAND2X1_1 ( .A(state_3_), .B(axi_wready), .Y(_abc_4169_new_n559_));
NAND2X1 NAND2X1_10 ( .A(re), .B(we), .Y(_abc_4169_new_n603_));
NAND2X1 NAND2X1_100 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_7_), .Y(bus_sync_axi_bus__abc_3843_new_n417_));
NAND2X1 NAND2X1_101 ( .A(bus_sync_axi_bus_reg_data2_8_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n419_));
NAND2X1 NAND2X1_102 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_8_), .Y(bus_sync_axi_bus__abc_3843_new_n420_));
NAND2X1 NAND2X1_103 ( .A(bus_sync_axi_bus_reg_data2_9_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n422_));
NAND2X1 NAND2X1_104 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_9_), .Y(bus_sync_axi_bus__abc_3843_new_n423_));
NAND2X1 NAND2X1_105 ( .A(bus_sync_axi_bus_reg_data2_10_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n425_));
NAND2X1 NAND2X1_106 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_10_), .Y(bus_sync_axi_bus__abc_3843_new_n426_));
NAND2X1 NAND2X1_107 ( .A(bus_sync_axi_bus_reg_data2_11_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n428_));
NAND2X1 NAND2X1_108 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_11_), .Y(bus_sync_axi_bus__abc_3843_new_n429_));
NAND2X1 NAND2X1_109 ( .A(bus_sync_axi_bus_reg_data2_12_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n431_));
NAND2X1 NAND2X1_11 ( .A(_abc_4169_new_n604_), .B(_abc_4169_new_n605_), .Y(_abc_4169_new_n606_));
NAND2X1 NAND2X1_110 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_12_), .Y(bus_sync_axi_bus__abc_3843_new_n432_));
NAND2X1 NAND2X1_111 ( .A(bus_sync_axi_bus_reg_data2_13_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n434_));
NAND2X1 NAND2X1_112 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_13_), .Y(bus_sync_axi_bus__abc_3843_new_n435_));
NAND2X1 NAND2X1_113 ( .A(bus_sync_axi_bus_reg_data2_14_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n437_));
NAND2X1 NAND2X1_114 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_14_), .Y(bus_sync_axi_bus__abc_3843_new_n438_));
NAND2X1 NAND2X1_115 ( .A(bus_sync_axi_bus_reg_data2_15_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n440_));
NAND2X1 NAND2X1_116 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_15_), .Y(bus_sync_axi_bus__abc_3843_new_n441_));
NAND2X1 NAND2X1_117 ( .A(bus_sync_axi_bus_reg_data2_16_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n443_));
NAND2X1 NAND2X1_118 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_16_), .Y(bus_sync_axi_bus__abc_3843_new_n444_));
NAND2X1 NAND2X1_119 ( .A(bus_sync_axi_bus_reg_data2_17_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n446_));
NAND2X1 NAND2X1_12 ( .A(_abc_4169_new_n603_), .B(_abc_4169_new_n606_), .Y(_abc_4169_new_n607_));
NAND2X1 NAND2X1_120 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_17_), .Y(bus_sync_axi_bus__abc_3843_new_n447_));
NAND2X1 NAND2X1_121 ( .A(bus_sync_axi_bus_reg_data2_18_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n449_));
NAND2X1 NAND2X1_122 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_18_), .Y(bus_sync_axi_bus__abc_3843_new_n450_));
NAND2X1 NAND2X1_123 ( .A(bus_sync_axi_bus_reg_data2_19_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n452_));
NAND2X1 NAND2X1_124 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_19_), .Y(bus_sync_axi_bus__abc_3843_new_n453_));
NAND2X1 NAND2X1_125 ( .A(bus_sync_axi_bus_reg_data2_20_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n455_));
NAND2X1 NAND2X1_126 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_20_), .Y(bus_sync_axi_bus__abc_3843_new_n456_));
NAND2X1 NAND2X1_127 ( .A(bus_sync_axi_bus_reg_data2_21_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n458_));
NAND2X1 NAND2X1_128 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_21_), .Y(bus_sync_axi_bus__abc_3843_new_n459_));
NAND2X1 NAND2X1_129 ( .A(bus_sync_axi_bus_reg_data2_22_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n461_));
NAND2X1 NAND2X1_13 ( .A(_abc_4169_new_n608_), .B(_abc_4169_new_n609_), .Y(_abc_4169_new_n610_));
NAND2X1 NAND2X1_130 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_22_), .Y(bus_sync_axi_bus__abc_3843_new_n462_));
NAND2X1 NAND2X1_131 ( .A(bus_sync_axi_bus_reg_data2_23_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n464_));
NAND2X1 NAND2X1_132 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_23_), .Y(bus_sync_axi_bus__abc_3843_new_n465_));
NAND2X1 NAND2X1_133 ( .A(bus_sync_axi_bus_reg_data2_24_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n467_));
NAND2X1 NAND2X1_134 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_24_), .Y(bus_sync_axi_bus__abc_3843_new_n468_));
NAND2X1 NAND2X1_135 ( .A(bus_sync_axi_bus_reg_data2_25_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n470_));
NAND2X1 NAND2X1_136 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_25_), .Y(bus_sync_axi_bus__abc_3843_new_n471_));
NAND2X1 NAND2X1_137 ( .A(bus_sync_axi_bus_reg_data2_26_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n473_));
NAND2X1 NAND2X1_138 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_26_), .Y(bus_sync_axi_bus__abc_3843_new_n474_));
NAND2X1 NAND2X1_139 ( .A(bus_sync_axi_bus_reg_data2_27_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n476_));
NAND2X1 NAND2X1_14 ( .A(_abc_4169_new_n616_), .B(_abc_4169_new_n617_), .Y(_abc_4169_new_n618_));
NAND2X1 NAND2X1_140 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_27_), .Y(bus_sync_axi_bus__abc_3843_new_n477_));
NAND2X1 NAND2X1_141 ( .A(bus_sync_axi_bus_reg_data2_28_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n479_));
NAND2X1 NAND2X1_142 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_28_), .Y(bus_sync_axi_bus__abc_3843_new_n480_));
NAND2X1 NAND2X1_143 ( .A(bus_sync_axi_bus_reg_data2_29_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n482_));
NAND2X1 NAND2X1_144 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_29_), .Y(bus_sync_axi_bus__abc_3843_new_n483_));
NAND2X1 NAND2X1_145 ( .A(bus_sync_axi_bus_reg_data2_30_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n485_));
NAND2X1 NAND2X1_146 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_30_), .Y(bus_sync_axi_bus__abc_3843_new_n486_));
NAND2X1 NAND2X1_147 ( .A(bus_sync_axi_bus_reg_data2_31_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n488_));
NAND2X1 NAND2X1_148 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_31_), .Y(bus_sync_axi_bus__abc_3843_new_n489_));
NAND2X1 NAND2X1_149 ( .A(bus_sync_axi_bus_reg_data2_32_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n491_));
NAND2X1 NAND2X1_15 ( .A(_abc_4169_new_n619_), .B(_abc_4169_new_n620_), .Y(_abc_4169_new_n621_));
NAND2X1 NAND2X1_150 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_32_), .Y(bus_sync_axi_bus__abc_3843_new_n492_));
NAND2X1 NAND2X1_151 ( .A(bus_sync_axi_bus_reg_data2_33_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n494_));
NAND2X1 NAND2X1_152 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_33_), .Y(bus_sync_axi_bus__abc_3843_new_n495_));
NAND2X1 NAND2X1_153 ( .A(bus_sync_axi_bus_reg_data2_34_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n497_));
NAND2X1 NAND2X1_154 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_34_), .Y(bus_sync_axi_bus__abc_3843_new_n498_));
NAND2X1 NAND2X1_155 ( .A(bus_sync_axi_bus_reg_data2_35_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n500_));
NAND2X1 NAND2X1_156 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_35_), .Y(bus_sync_axi_bus__abc_3843_new_n501_));
NAND2X1 NAND2X1_157 ( .A(bus_sync_axi_bus_reg_data2_36_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n503_));
NAND2X1 NAND2X1_158 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_36_), .Y(bus_sync_axi_bus__abc_3843_new_n504_));
NAND2X1 NAND2X1_159 ( .A(bus_sync_axi_bus_reg_data2_37_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n506_));
NAND2X1 NAND2X1_16 ( .A(_abc_4169_new_n622_), .B(_abc_4169_new_n615_), .Y(_abc_4169_new_n623_));
NAND2X1 NAND2X1_160 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_37_), .Y(bus_sync_axi_bus__abc_3843_new_n507_));
NAND2X1 NAND2X1_161 ( .A(bus_sync_axi_bus_reg_data2_38_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n509_));
NAND2X1 NAND2X1_162 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_38_), .Y(bus_sync_axi_bus__abc_3843_new_n510_));
NAND2X1 NAND2X1_163 ( .A(bus_sync_axi_bus_reg_data2_39_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n512_));
NAND2X1 NAND2X1_164 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_39_), .Y(bus_sync_axi_bus__abc_3843_new_n513_));
NAND2X1 NAND2X1_165 ( .A(bus_sync_axi_bus_reg_data2_40_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n515_));
NAND2X1 NAND2X1_166 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_40_), .Y(bus_sync_axi_bus__abc_3843_new_n516_));
NAND2X1 NAND2X1_167 ( .A(bus_sync_axi_bus_reg_data2_41_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n518_));
NAND2X1 NAND2X1_168 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_41_), .Y(bus_sync_axi_bus__abc_3843_new_n519_));
NAND2X1 NAND2X1_169 ( .A(bus_sync_axi_bus_reg_data2_42_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n521_));
NAND2X1 NAND2X1_17 ( .A(_abc_4169_new_n624_), .B(_abc_4169_new_n625_), .Y(_abc_4169_new_n626_));
NAND2X1 NAND2X1_170 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_42_), .Y(bus_sync_axi_bus__abc_3843_new_n522_));
NAND2X1 NAND2X1_171 ( .A(bus_sync_axi_bus_reg_data2_43_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n524_));
NAND2X1 NAND2X1_172 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_43_), .Y(bus_sync_axi_bus__abc_3843_new_n525_));
NAND2X1 NAND2X1_173 ( .A(bus_sync_axi_bus_reg_data2_44_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n527_));
NAND2X1 NAND2X1_174 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_44_), .Y(bus_sync_axi_bus__abc_3843_new_n528_));
NAND2X1 NAND2X1_175 ( .A(bus_sync_axi_bus_reg_data2_45_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n530_));
NAND2X1 NAND2X1_176 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_45_), .Y(bus_sync_axi_bus__abc_3843_new_n531_));
NAND2X1 NAND2X1_177 ( .A(bus_sync_axi_bus_reg_data2_46_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n533_));
NAND2X1 NAND2X1_178 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_46_), .Y(bus_sync_axi_bus__abc_3843_new_n534_));
NAND2X1 NAND2X1_179 ( .A(bus_sync_axi_bus_reg_data2_47_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n536_));
NAND2X1 NAND2X1_18 ( .A(_abc_4169_new_n632_), .B(_abc_4169_new_n633_), .Y(_abc_4169_new_n634_));
NAND2X1 NAND2X1_180 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_47_), .Y(bus_sync_axi_bus__abc_3843_new_n537_));
NAND2X1 NAND2X1_181 ( .A(bus_sync_axi_bus_reg_data2_48_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n539_));
NAND2X1 NAND2X1_182 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_48_), .Y(bus_sync_axi_bus__abc_3843_new_n540_));
NAND2X1 NAND2X1_183 ( .A(bus_sync_axi_bus_reg_data2_49_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n542_));
NAND2X1 NAND2X1_184 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_49_), .Y(bus_sync_axi_bus__abc_3843_new_n543_));
NAND2X1 NAND2X1_185 ( .A(bus_sync_axi_bus_reg_data2_50_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n545_));
NAND2X1 NAND2X1_186 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_50_), .Y(bus_sync_axi_bus__abc_3843_new_n546_));
NAND2X1 NAND2X1_187 ( .A(bus_sync_axi_bus_reg_data2_51_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n548_));
NAND2X1 NAND2X1_188 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_51_), .Y(bus_sync_axi_bus__abc_3843_new_n549_));
NAND2X1 NAND2X1_189 ( .A(bus_sync_axi_bus_reg_data2_52_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n551_));
NAND2X1 NAND2X1_19 ( .A(_abc_4169_new_n631_), .B(_abc_4169_new_n639_), .Y(_abc_4169_new_n640_));
NAND2X1 NAND2X1_190 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_52_), .Y(bus_sync_axi_bus__abc_3843_new_n552_));
NAND2X1 NAND2X1_191 ( .A(bus_sync_axi_bus_reg_data2_53_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n554_));
NAND2X1 NAND2X1_192 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_53_), .Y(bus_sync_axi_bus__abc_3843_new_n555_));
NAND2X1 NAND2X1_193 ( .A(bus_sync_axi_bus_reg_data2_54_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n557_));
NAND2X1 NAND2X1_194 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_54_), .Y(bus_sync_axi_bus__abc_3843_new_n558_));
NAND2X1 NAND2X1_195 ( .A(bus_sync_axi_bus_reg_data2_55_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n560_));
NAND2X1 NAND2X1_196 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_55_), .Y(bus_sync_axi_bus__abc_3843_new_n561_));
NAND2X1 NAND2X1_197 ( .A(bus_sync_axi_bus_reg_data2_56_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n563_));
NAND2X1 NAND2X1_198 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_56_), .Y(bus_sync_axi_bus__abc_3843_new_n564_));
NAND2X1 NAND2X1_199 ( .A(bus_sync_axi_bus_reg_data2_57_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n566_));
NAND2X1 NAND2X1_2 ( .A(_abc_4169_new_n558_), .B(_abc_4169_new_n562_), .Y(axi_wvalid));
NAND2X1 NAND2X1_20 ( .A(bus_cap_0_), .B(_abc_4169_new_n641_), .Y(_abc_4169_new_n642_));
NAND2X1 NAND2X1_200 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_57_), .Y(bus_sync_axi_bus__abc_3843_new_n567_));
NAND2X1 NAND2X1_201 ( .A(bus_sync_axi_bus_reg_data2_58_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n569_));
NAND2X1 NAND2X1_202 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_58_), .Y(bus_sync_axi_bus__abc_3843_new_n570_));
NAND2X1 NAND2X1_203 ( .A(bus_sync_axi_bus_reg_data2_59_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n572_));
NAND2X1 NAND2X1_204 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_59_), .Y(bus_sync_axi_bus__abc_3843_new_n573_));
NAND2X1 NAND2X1_205 ( .A(bus_sync_axi_bus_reg_data2_60_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n575_));
NAND2X1 NAND2X1_206 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_60_), .Y(bus_sync_axi_bus__abc_3843_new_n576_));
NAND2X1 NAND2X1_207 ( .A(bus_sync_axi_bus_reg_data2_61_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n578_));
NAND2X1 NAND2X1_208 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_61_), .Y(bus_sync_axi_bus__abc_3843_new_n579_));
NAND2X1 NAND2X1_209 ( .A(bus_sync_axi_bus_reg_data2_62_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n581_));
NAND2X1 NAND2X1_21 ( .A(bus_cap_1_), .B(_abc_4169_new_n641_), .Y(_abc_4169_new_n648_));
NAND2X1 NAND2X1_210 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_62_), .Y(bus_sync_axi_bus__abc_3843_new_n582_));
NAND2X1 NAND2X1_211 ( .A(bus_sync_axi_bus_reg_data2_63_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n584_));
NAND2X1 NAND2X1_212 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_63_), .Y(bus_sync_axi_bus__abc_3843_new_n585_));
NAND2X1 NAND2X1_213 ( .A(bus_sync_rdata_reg_data2_0_), .B(bus_sync_rdata__abc_3651_new_n266_), .Y(bus_sync_rdata__abc_3651_new_n267_));
NAND2X1 NAND2X1_214 ( .A(bus_sync_rdata_reg_data1_0_), .B(bus_sync_rdata_EECLK2), .Y(bus_sync_rdata__abc_3651_new_n268_));
NAND2X1 NAND2X1_215 ( .A(bus_sync_rdata_reg_data2_1_), .B(bus_sync_rdata__abc_3651_new_n266_), .Y(bus_sync_rdata__abc_3651_new_n270_));
NAND2X1 NAND2X1_216 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_1_), .Y(bus_sync_rdata__abc_3651_new_n271_));
NAND2X1 NAND2X1_217 ( .A(bus_sync_rdata_reg_data2_2_), .B(bus_sync_rdata__abc_3651_new_n266_), .Y(bus_sync_rdata__abc_3651_new_n273_));
NAND2X1 NAND2X1_218 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_2_), .Y(bus_sync_rdata__abc_3651_new_n274_));
NAND2X1 NAND2X1_219 ( .A(bus_sync_rdata_reg_data2_3_), .B(bus_sync_rdata__abc_3651_new_n266_), .Y(bus_sync_rdata__abc_3651_new_n276_));
NAND2X1 NAND2X1_22 ( .A(bus_cap_2_), .B(_abc_4169_new_n641_), .Y(_abc_4169_new_n658_));
NAND2X1 NAND2X1_220 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_3_), .Y(bus_sync_rdata__abc_3651_new_n277_));
NAND2X1 NAND2X1_221 ( .A(bus_sync_rdata_reg_data2_4_), .B(bus_sync_rdata__abc_3651_new_n266_), .Y(bus_sync_rdata__abc_3651_new_n279_));
NAND2X1 NAND2X1_222 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_4_), .Y(bus_sync_rdata__abc_3651_new_n280_));
NAND2X1 NAND2X1_223 ( .A(bus_sync_rdata_reg_data2_5_), .B(bus_sync_rdata__abc_3651_new_n266_), .Y(bus_sync_rdata__abc_3651_new_n282_));
NAND2X1 NAND2X1_224 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_5_), .Y(bus_sync_rdata__abc_3651_new_n283_));
NAND2X1 NAND2X1_225 ( .A(bus_sync_rdata_reg_data2_6_), .B(bus_sync_rdata__abc_3651_new_n266_), .Y(bus_sync_rdata__abc_3651_new_n285_));
NAND2X1 NAND2X1_226 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_6_), .Y(bus_sync_rdata__abc_3651_new_n286_));
NAND2X1 NAND2X1_227 ( .A(bus_sync_rdata_reg_data2_7_), .B(bus_sync_rdata__abc_3651_new_n266_), .Y(bus_sync_rdata__abc_3651_new_n288_));
NAND2X1 NAND2X1_228 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_7_), .Y(bus_sync_rdata__abc_3651_new_n289_));
NAND2X1 NAND2X1_229 ( .A(bus_sync_rdata_reg_data2_8_), .B(bus_sync_rdata__abc_3651_new_n266_), .Y(bus_sync_rdata__abc_3651_new_n291_));
NAND2X1 NAND2X1_23 ( .A(bus_cap_3_), .B(_abc_4169_new_n641_), .Y(_abc_4169_new_n665_));
NAND2X1 NAND2X1_230 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_8_), .Y(bus_sync_rdata__abc_3651_new_n292_));
NAND2X1 NAND2X1_231 ( .A(bus_sync_rdata_reg_data2_9_), .B(bus_sync_rdata__abc_3651_new_n266_), .Y(bus_sync_rdata__abc_3651_new_n294_));
NAND2X1 NAND2X1_232 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_9_), .Y(bus_sync_rdata__abc_3651_new_n295_));
NAND2X1 NAND2X1_233 ( .A(bus_sync_rdata_reg_data2_10_), .B(bus_sync_rdata__abc_3651_new_n266_), .Y(bus_sync_rdata__abc_3651_new_n297_));
NAND2X1 NAND2X1_234 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_10_), .Y(bus_sync_rdata__abc_3651_new_n298_));
NAND2X1 NAND2X1_235 ( .A(bus_sync_rdata_reg_data2_11_), .B(bus_sync_rdata__abc_3651_new_n266_), .Y(bus_sync_rdata__abc_3651_new_n300_));
NAND2X1 NAND2X1_236 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_11_), .Y(bus_sync_rdata__abc_3651_new_n301_));
NAND2X1 NAND2X1_237 ( .A(bus_sync_rdata_reg_data2_12_), .B(bus_sync_rdata__abc_3651_new_n266_), .Y(bus_sync_rdata__abc_3651_new_n303_));
NAND2X1 NAND2X1_238 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_12_), .Y(bus_sync_rdata__abc_3651_new_n304_));
NAND2X1 NAND2X1_239 ( .A(bus_sync_rdata_reg_data2_13_), .B(bus_sync_rdata__abc_3651_new_n266_), .Y(bus_sync_rdata__abc_3651_new_n306_));
NAND2X1 NAND2X1_24 ( .A(RST), .B(_abc_4169_new_n668_), .Y(_abc_4169_new_n669_));
NAND2X1 NAND2X1_240 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_13_), .Y(bus_sync_rdata__abc_3651_new_n307_));
NAND2X1 NAND2X1_241 ( .A(bus_sync_rdata_reg_data2_14_), .B(bus_sync_rdata__abc_3651_new_n266_), .Y(bus_sync_rdata__abc_3651_new_n309_));
NAND2X1 NAND2X1_242 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_14_), .Y(bus_sync_rdata__abc_3651_new_n310_));
NAND2X1 NAND2X1_243 ( .A(bus_sync_rdata_reg_data2_15_), .B(bus_sync_rdata__abc_3651_new_n266_), .Y(bus_sync_rdata__abc_3651_new_n312_));
NAND2X1 NAND2X1_244 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_15_), .Y(bus_sync_rdata__abc_3651_new_n313_));
NAND2X1 NAND2X1_245 ( .A(bus_sync_rdata_reg_data2_16_), .B(bus_sync_rdata__abc_3651_new_n266_), .Y(bus_sync_rdata__abc_3651_new_n315_));
NAND2X1 NAND2X1_246 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_16_), .Y(bus_sync_rdata__abc_3651_new_n316_));
NAND2X1 NAND2X1_247 ( .A(bus_sync_rdata_reg_data2_17_), .B(bus_sync_rdata__abc_3651_new_n266_), .Y(bus_sync_rdata__abc_3651_new_n318_));
NAND2X1 NAND2X1_248 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_17_), .Y(bus_sync_rdata__abc_3651_new_n319_));
NAND2X1 NAND2X1_249 ( .A(bus_sync_rdata_reg_data2_18_), .B(bus_sync_rdata__abc_3651_new_n266_), .Y(bus_sync_rdata__abc_3651_new_n321_));
NAND2X1 NAND2X1_25 ( .A(bus_cap_4_), .B(_abc_4169_new_n641_), .Y(_abc_4169_new_n671_));
NAND2X1 NAND2X1_250 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_18_), .Y(bus_sync_rdata__abc_3651_new_n322_));
NAND2X1 NAND2X1_251 ( .A(bus_sync_rdata_reg_data2_19_), .B(bus_sync_rdata__abc_3651_new_n266_), .Y(bus_sync_rdata__abc_3651_new_n324_));
NAND2X1 NAND2X1_252 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_19_), .Y(bus_sync_rdata__abc_3651_new_n325_));
NAND2X1 NAND2X1_253 ( .A(bus_sync_rdata_reg_data2_20_), .B(bus_sync_rdata__abc_3651_new_n266_), .Y(bus_sync_rdata__abc_3651_new_n327_));
NAND2X1 NAND2X1_254 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_20_), .Y(bus_sync_rdata__abc_3651_new_n328_));
NAND2X1 NAND2X1_255 ( .A(bus_sync_rdata_reg_data2_21_), .B(bus_sync_rdata__abc_3651_new_n266_), .Y(bus_sync_rdata__abc_3651_new_n330_));
NAND2X1 NAND2X1_256 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_21_), .Y(bus_sync_rdata__abc_3651_new_n331_));
NAND2X1 NAND2X1_257 ( .A(bus_sync_rdata_reg_data2_22_), .B(bus_sync_rdata__abc_3651_new_n266_), .Y(bus_sync_rdata__abc_3651_new_n333_));
NAND2X1 NAND2X1_258 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_22_), .Y(bus_sync_rdata__abc_3651_new_n334_));
NAND2X1 NAND2X1_259 ( .A(bus_sync_rdata_reg_data2_23_), .B(bus_sync_rdata__abc_3651_new_n266_), .Y(bus_sync_rdata__abc_3651_new_n336_));
NAND2X1 NAND2X1_26 ( .A(RST), .B(_abc_4169_new_n674_), .Y(_abc_4169_new_n675_));
NAND2X1 NAND2X1_260 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_23_), .Y(bus_sync_rdata__abc_3651_new_n337_));
NAND2X1 NAND2X1_261 ( .A(bus_sync_rdata_reg_data2_24_), .B(bus_sync_rdata__abc_3651_new_n266_), .Y(bus_sync_rdata__abc_3651_new_n339_));
NAND2X1 NAND2X1_262 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_24_), .Y(bus_sync_rdata__abc_3651_new_n340_));
NAND2X1 NAND2X1_263 ( .A(bus_sync_rdata_reg_data2_25_), .B(bus_sync_rdata__abc_3651_new_n266_), .Y(bus_sync_rdata__abc_3651_new_n342_));
NAND2X1 NAND2X1_264 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_25_), .Y(bus_sync_rdata__abc_3651_new_n343_));
NAND2X1 NAND2X1_265 ( .A(bus_sync_rdata_reg_data2_26_), .B(bus_sync_rdata__abc_3651_new_n266_), .Y(bus_sync_rdata__abc_3651_new_n345_));
NAND2X1 NAND2X1_266 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_26_), .Y(bus_sync_rdata__abc_3651_new_n346_));
NAND2X1 NAND2X1_267 ( .A(bus_sync_rdata_reg_data2_27_), .B(bus_sync_rdata__abc_3651_new_n266_), .Y(bus_sync_rdata__abc_3651_new_n348_));
NAND2X1 NAND2X1_268 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_27_), .Y(bus_sync_rdata__abc_3651_new_n349_));
NAND2X1 NAND2X1_269 ( .A(bus_sync_rdata_reg_data2_28_), .B(bus_sync_rdata__abc_3651_new_n266_), .Y(bus_sync_rdata__abc_3651_new_n351_));
NAND2X1 NAND2X1_27 ( .A(bus_cap_5_), .B(_abc_4169_new_n641_), .Y(_abc_4169_new_n677_));
NAND2X1 NAND2X1_270 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_28_), .Y(bus_sync_rdata__abc_3651_new_n352_));
NAND2X1 NAND2X1_271 ( .A(bus_sync_rdata_reg_data2_29_), .B(bus_sync_rdata__abc_3651_new_n266_), .Y(bus_sync_rdata__abc_3651_new_n354_));
NAND2X1 NAND2X1_272 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_29_), .Y(bus_sync_rdata__abc_3651_new_n355_));
NAND2X1 NAND2X1_273 ( .A(bus_sync_rdata_reg_data2_30_), .B(bus_sync_rdata__abc_3651_new_n266_), .Y(bus_sync_rdata__abc_3651_new_n357_));
NAND2X1 NAND2X1_274 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_30_), .Y(bus_sync_rdata__abc_3651_new_n358_));
NAND2X1 NAND2X1_275 ( .A(bus_sync_rdata_reg_data2_31_), .B(bus_sync_rdata__abc_3651_new_n266_), .Y(bus_sync_rdata__abc_3651_new_n360_));
NAND2X1 NAND2X1_276 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_31_), .Y(bus_sync_rdata__abc_3651_new_n361_));
NAND2X1 NAND2X1_277 ( .A(bus_sync_state_machine_reg_data2_0_), .B(bus_sync_state_machine__abc_3817_new_n34_), .Y(bus_sync_state_machine__abc_3817_new_n35_));
NAND2X1 NAND2X1_278 ( .A(bus_sync_state_machine_reg_data1_0_), .B(bus_sync_state_machine_EECLK1), .Y(bus_sync_state_machine__abc_3817_new_n36_));
NAND2X1 NAND2X1_279 ( .A(bus_sync_state_machine_reg_data2_1_), .B(bus_sync_state_machine__abc_3817_new_n34_), .Y(bus_sync_state_machine__abc_3817_new_n38_));
NAND2X1 NAND2X1_28 ( .A(RST), .B(_abc_4169_new_n680_), .Y(_abc_4169_new_n681_));
NAND2X1 NAND2X1_280 ( .A(bus_sync_state_machine_EECLK1), .B(bus_sync_state_machine_reg_data1_1_), .Y(bus_sync_state_machine__abc_3817_new_n39_));
NAND2X1 NAND2X1_281 ( .A(bus_sync_state_machine_reg_data2_2_), .B(bus_sync_state_machine__abc_3817_new_n34_), .Y(bus_sync_state_machine__abc_3817_new_n41_));
NAND2X1 NAND2X1_282 ( .A(bus_sync_state_machine_EECLK1), .B(bus_sync_state_machine_reg_data1_2_), .Y(bus_sync_state_machine__abc_3817_new_n42_));
NAND2X1 NAND2X1_283 ( .A(bus_sync_state_machine_reg_data2_3_), .B(bus_sync_state_machine__abc_3817_new_n34_), .Y(bus_sync_state_machine__abc_3817_new_n44_));
NAND2X1 NAND2X1_284 ( .A(bus_sync_state_machine_EECLK1), .B(bus_sync_state_machine_reg_data1_3_), .Y(bus_sync_state_machine__abc_3817_new_n45_));
NAND2X1 NAND2X1_285 ( .A(bus_sync_status_reg_data2_0_), .B(bus_sync_status__abc_3630_new_n28_), .Y(bus_sync_status__abc_3630_new_n29_));
NAND2X1 NAND2X1_286 ( .A(bus_sync_status_reg_data1_0_), .B(bus_sync_status_EECLK2), .Y(bus_sync_status__abc_3630_new_n30_));
NAND2X1 NAND2X1_287 ( .A(bus_sync_status_reg_data2_1_), .B(bus_sync_status__abc_3630_new_n28_), .Y(bus_sync_status__abc_3630_new_n32_));
NAND2X1 NAND2X1_288 ( .A(bus_sync_status_EECLK2), .B(bus_sync_status_reg_data1_1_), .Y(bus_sync_status__abc_3630_new_n33_));
NAND2X1 NAND2X1_289 ( .A(bus_sync_status_reg_data2_2_), .B(bus_sync_status__abc_3630_new_n28_), .Y(bus_sync_status__abc_3630_new_n35_));
NAND2X1 NAND2X1_29 ( .A(bus_cap_6_), .B(_abc_4169_new_n641_), .Y(_abc_4169_new_n683_));
NAND2X1 NAND2X1_290 ( .A(bus_sync_status_EECLK2), .B(bus_sync_status_reg_data1_2_), .Y(bus_sync_status__abc_3630_new_n36_));
NAND2X1 NAND2X1_3 ( .A(state_1_), .B(fini_spi_clk), .Y(_abc_4169_new_n569_));
NAND2X1 NAND2X1_30 ( .A(RST), .B(_abc_4169_new_n686_), .Y(_abc_4169_new_n687_));
NAND2X1 NAND2X1_31 ( .A(bus_cap_7_), .B(_abc_4169_new_n641_), .Y(_abc_4169_new_n689_));
NAND2X1 NAND2X1_32 ( .A(RST), .B(_abc_4169_new_n692_), .Y(_abc_4169_new_n693_));
NAND2X1 NAND2X1_33 ( .A(bus_cap_8_), .B(_abc_4169_new_n641_), .Y(_abc_4169_new_n695_));
NAND2X1 NAND2X1_34 ( .A(RST), .B(_abc_4169_new_n698_), .Y(_abc_4169_new_n699_));
NAND2X1 NAND2X1_35 ( .A(bus_cap_9_), .B(_abc_4169_new_n641_), .Y(_abc_4169_new_n701_));
NAND2X1 NAND2X1_36 ( .A(RST), .B(_abc_4169_new_n704_), .Y(_abc_4169_new_n705_));
NAND2X1 NAND2X1_37 ( .A(bus_cap_10_), .B(_abc_4169_new_n641_), .Y(_abc_4169_new_n707_));
NAND2X1 NAND2X1_38 ( .A(RST), .B(_abc_4169_new_n710_), .Y(_abc_4169_new_n711_));
NAND2X1 NAND2X1_39 ( .A(bus_cap_11_), .B(_abc_4169_new_n641_), .Y(_abc_4169_new_n713_));
NAND2X1 NAND2X1_4 ( .A(RST), .B(state_6_), .Y(_abc_4169_new_n571_));
NAND2X1 NAND2X1_40 ( .A(RST), .B(_abc_4169_new_n716_), .Y(_abc_4169_new_n717_));
NAND2X1 NAND2X1_41 ( .A(bus_cap_12_), .B(_abc_4169_new_n641_), .Y(_abc_4169_new_n719_));
NAND2X1 NAND2X1_42 ( .A(RST), .B(_abc_4169_new_n722_), .Y(_abc_4169_new_n723_));
NAND2X1 NAND2X1_43 ( .A(bus_cap_13_), .B(_abc_4169_new_n641_), .Y(_abc_4169_new_n725_));
NAND2X1 NAND2X1_44 ( .A(RST), .B(_abc_4169_new_n728_), .Y(_abc_4169_new_n729_));
NAND2X1 NAND2X1_45 ( .A(bus_cap_14_), .B(_abc_4169_new_n641_), .Y(_abc_4169_new_n731_));
NAND2X1 NAND2X1_46 ( .A(RST), .B(_abc_4169_new_n734_), .Y(_abc_4169_new_n735_));
NAND2X1 NAND2X1_47 ( .A(bus_cap_15_), .B(_abc_4169_new_n641_), .Y(_abc_4169_new_n737_));
NAND2X1 NAND2X1_48 ( .A(RST), .B(_abc_4169_new_n740_), .Y(_abc_4169_new_n741_));
NAND2X1 NAND2X1_49 ( .A(bus_cap_16_), .B(_abc_4169_new_n641_), .Y(_abc_4169_new_n743_));
NAND2X1 NAND2X1_5 ( .A(fini_spi_clk), .B(we_clk), .Y(_abc_4169_new_n572_));
NAND2X1 NAND2X1_50 ( .A(RST), .B(_abc_4169_new_n746_), .Y(_abc_4169_new_n747_));
NAND2X1 NAND2X1_51 ( .A(bus_cap_17_), .B(_abc_4169_new_n641_), .Y(_abc_4169_new_n749_));
NAND2X1 NAND2X1_52 ( .A(RST), .B(_abc_4169_new_n752_), .Y(_abc_4169_new_n753_));
NAND2X1 NAND2X1_53 ( .A(bus_cap_18_), .B(_abc_4169_new_n641_), .Y(_abc_4169_new_n755_));
NAND2X1 NAND2X1_54 ( .A(RST), .B(_abc_4169_new_n758_), .Y(_abc_4169_new_n759_));
NAND2X1 NAND2X1_55 ( .A(bus_cap_19_), .B(_abc_4169_new_n641_), .Y(_abc_4169_new_n761_));
NAND2X1 NAND2X1_56 ( .A(RST), .B(_abc_4169_new_n764_), .Y(_abc_4169_new_n765_));
NAND2X1 NAND2X1_57 ( .A(bus_cap_20_), .B(_abc_4169_new_n641_), .Y(_abc_4169_new_n767_));
NAND2X1 NAND2X1_58 ( .A(RST), .B(_abc_4169_new_n770_), .Y(_abc_4169_new_n771_));
NAND2X1 NAND2X1_59 ( .A(bus_cap_21_), .B(_abc_4169_new_n641_), .Y(_abc_4169_new_n773_));
NAND2X1 NAND2X1_6 ( .A(fini_spi_clk), .B(re_clk), .Y(_abc_4169_new_n574_));
NAND2X1 NAND2X1_60 ( .A(RST), .B(_abc_4169_new_n776_), .Y(_abc_4169_new_n777_));
NAND2X1 NAND2X1_61 ( .A(bus_cap_22_), .B(_abc_4169_new_n641_), .Y(_abc_4169_new_n779_));
NAND2X1 NAND2X1_62 ( .A(RST), .B(_abc_4169_new_n782_), .Y(_abc_4169_new_n783_));
NAND2X1 NAND2X1_63 ( .A(bus_cap_23_), .B(_abc_4169_new_n641_), .Y(_abc_4169_new_n785_));
NAND2X1 NAND2X1_64 ( .A(RST), .B(_abc_4169_new_n788_), .Y(_abc_4169_new_n789_));
NAND2X1 NAND2X1_65 ( .A(bus_cap_24_), .B(_abc_4169_new_n641_), .Y(_abc_4169_new_n791_));
NAND2X1 NAND2X1_66 ( .A(RST), .B(_abc_4169_new_n794_), .Y(_abc_4169_new_n795_));
NAND2X1 NAND2X1_67 ( .A(bus_cap_25_), .B(_abc_4169_new_n641_), .Y(_abc_4169_new_n797_));
NAND2X1 NAND2X1_68 ( .A(RST), .B(_abc_4169_new_n800_), .Y(_abc_4169_new_n801_));
NAND2X1 NAND2X1_69 ( .A(bus_cap_26_), .B(_abc_4169_new_n641_), .Y(_abc_4169_new_n803_));
NAND2X1 NAND2X1_7 ( .A(state_0_), .B(_abc_4169_new_n575_), .Y(_abc_4169_new_n576_));
NAND2X1 NAND2X1_70 ( .A(RST), .B(_abc_4169_new_n806_), .Y(_abc_4169_new_n807_));
NAND2X1 NAND2X1_71 ( .A(bus_cap_27_), .B(_abc_4169_new_n641_), .Y(_abc_4169_new_n809_));
NAND2X1 NAND2X1_72 ( .A(RST), .B(_abc_4169_new_n812_), .Y(_abc_4169_new_n813_));
NAND2X1 NAND2X1_73 ( .A(bus_cap_28_), .B(_abc_4169_new_n641_), .Y(_abc_4169_new_n815_));
NAND2X1 NAND2X1_74 ( .A(RST), .B(_abc_4169_new_n818_), .Y(_abc_4169_new_n819_));
NAND2X1 NAND2X1_75 ( .A(bus_cap_29_), .B(_abc_4169_new_n641_), .Y(_abc_4169_new_n821_));
NAND2X1 NAND2X1_76 ( .A(RST), .B(_abc_4169_new_n824_), .Y(_abc_4169_new_n825_));
NAND2X1 NAND2X1_77 ( .A(bus_cap_30_), .B(_abc_4169_new_n641_), .Y(_abc_4169_new_n827_));
NAND2X1 NAND2X1_78 ( .A(RST), .B(_abc_4169_new_n830_), .Y(_abc_4169_new_n831_));
NAND2X1 NAND2X1_79 ( .A(DOUT), .B(_abc_4169_new_n641_), .Y(_abc_4169_new_n833_));
NAND2X1 NAND2X1_8 ( .A(RST), .B(state_4_), .Y(_abc_4169_new_n579_));
NAND2X1 NAND2X1_80 ( .A(RST), .B(_abc_4169_new_n836_), .Y(_abc_4169_new_n837_));
NAND2X1 NAND2X1_81 ( .A(_abc_4169_new_n937_), .B(_abc_4169_new_n1036_), .Y(_abc_4169_new_n1037_));
NAND2X1 NAND2X1_82 ( .A(RST), .B(_abc_4169_new_n937_), .Y(_0counter_65_0__0_));
NAND2X1 NAND2X1_83 ( .A(counter_1_), .B(_abc_4169_new_n937_), .Y(_abc_4169_new_n1339_));
NAND2X1 NAND2X1_84 ( .A(counter_0_), .B(_abc_4169_new_n937_), .Y(_abc_4169_new_n1343_));
NAND2X1 NAND2X1_85 ( .A(bus_sync_axi_bus_reg_data2_0_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n395_));
NAND2X1 NAND2X1_86 ( .A(bus_sync_axi_bus_reg_data1_0_), .B(bus_sync_axi_bus_EECLK1), .Y(bus_sync_axi_bus__abc_3843_new_n396_));
NAND2X1 NAND2X1_87 ( .A(bus_sync_axi_bus_reg_data2_1_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n398_));
NAND2X1 NAND2X1_88 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_1_), .Y(bus_sync_axi_bus__abc_3843_new_n399_));
NAND2X1 NAND2X1_89 ( .A(bus_sync_axi_bus_reg_data2_2_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n401_));
NAND2X1 NAND2X1_9 ( .A(_abc_4169_new_n562_), .B(_abc_4169_new_n583_), .Y(axi_awvalid));
NAND2X1 NAND2X1_90 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_2_), .Y(bus_sync_axi_bus__abc_3843_new_n402_));
NAND2X1 NAND2X1_91 ( .A(bus_sync_axi_bus_reg_data2_3_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n404_));
NAND2X1 NAND2X1_92 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_3_), .Y(bus_sync_axi_bus__abc_3843_new_n405_));
NAND2X1 NAND2X1_93 ( .A(bus_sync_axi_bus_reg_data2_4_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n407_));
NAND2X1 NAND2X1_94 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_4_), .Y(bus_sync_axi_bus__abc_3843_new_n408_));
NAND2X1 NAND2X1_95 ( .A(bus_sync_axi_bus_reg_data2_5_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n410_));
NAND2X1 NAND2X1_96 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_5_), .Y(bus_sync_axi_bus__abc_3843_new_n411_));
NAND2X1 NAND2X1_97 ( .A(bus_sync_axi_bus_reg_data2_6_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n413_));
NAND2X1 NAND2X1_98 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_6_), .Y(bus_sync_axi_bus__abc_3843_new_n414_));
NAND2X1 NAND2X1_99 ( .A(bus_sync_axi_bus_reg_data2_7_), .B(bus_sync_axi_bus__abc_3843_new_n394_), .Y(bus_sync_axi_bus__abc_3843_new_n416_));
NAND3X1 NAND3X1_1 ( .A(_abc_4169_new_n583_), .B(_abc_4169_new_n585_), .C(_abc_4169_new_n587_), .Y(busy));
NAND3X1 NAND3X1_2 ( .A(we), .B(DATA), .C(counter_1_), .Y(_abc_4169_new_n598_));
NAND3X1 NAND3X1_3 ( .A(_abc_4169_new_n611_), .B(_abc_4169_new_n612_), .C(_abc_4169_new_n613_), .Y(_abc_4169_new_n614_));
NAND3X1 NAND3X1_4 ( .A(_abc_4169_new_n627_), .B(_abc_4169_new_n628_), .C(_abc_4169_new_n629_), .Y(_abc_4169_new_n630_));
NAND3X1 NAND3X1_5 ( .A(_abc_4169_new_n635_), .B(_abc_4169_new_n636_), .C(_abc_4169_new_n637_), .Y(_abc_4169_new_n638_));
NAND3X1 NAND3X1_6 ( .A(we), .B(counter_65_), .C(_abc_4169_new_n937_), .Y(_abc_4169_new_n938_));
NAND3X1 NAND3X1_7 ( .A(counter_65_), .B(_abc_4169_new_n937_), .C(_abc_4169_new_n1335_), .Y(_abc_4169_new_n1336_));
NAND3X1 NAND3X1_8 ( .A(RST), .B(state_4_), .C(axi_rvalid), .Y(_abc_4169_new_n1346_));
NAND3X1 NAND3X1_9 ( .A(state_7_), .B(RST), .C(axi_bvalid), .Y(_abc_4169_new_n1348_));
NOR2X1 NOR2X1_1 ( .A(state_3_), .B(axi_bready), .Y(_abc_4169_new_n562_));
NOR2X1 NOR2X1_10 ( .A(we), .B(DATA), .Y(_abc_4169_new_n599_));
NOR2X1 NOR2X1_11 ( .A(counter_16_), .B(counter_17_), .Y(_abc_4169_new_n608_));
NOR2X1 NOR2X1_12 ( .A(counter_14_), .B(counter_15_), .Y(_abc_4169_new_n609_));
NOR2X1 NOR2X1_13 ( .A(counter_4_), .B(counter_5_), .Y(_abc_4169_new_n613_));
NOR2X1 NOR2X1_14 ( .A(_abc_4169_new_n610_), .B(_abc_4169_new_n614_), .Y(_abc_4169_new_n615_));
NOR2X1 NOR2X1_15 ( .A(counter_28_), .B(counter_29_), .Y(_abc_4169_new_n616_));
NOR2X1 NOR2X1_16 ( .A(counter_26_), .B(counter_27_), .Y(_abc_4169_new_n617_));
NOR2X1 NOR2X1_17 ( .A(counter_24_), .B(counter_25_), .Y(_abc_4169_new_n619_));
NOR2X1 NOR2X1_18 ( .A(counter_22_), .B(counter_23_), .Y(_abc_4169_new_n620_));
NOR2X1 NOR2X1_19 ( .A(_abc_4169_new_n618_), .B(_abc_4169_new_n621_), .Y(_abc_4169_new_n622_));
NOR2X1 NOR2X1_2 ( .A(_abc_4169_new_n564_), .B(_abc_4169_new_n566_), .Y(_abc_2903_auto_fsm_map_cc_170_map_fsm_402_3_));
NOR2X1 NOR2X1_20 ( .A(counter_12_), .B(counter_13_), .Y(_abc_4169_new_n624_));
NOR2X1 NOR2X1_21 ( .A(counter_10_), .B(counter_11_), .Y(_abc_4169_new_n625_));
NOR2X1 NOR2X1_22 ( .A(counter_8_), .B(counter_9_), .Y(_abc_4169_new_n629_));
NOR2X1 NOR2X1_23 ( .A(_abc_4169_new_n626_), .B(_abc_4169_new_n630_), .Y(_abc_4169_new_n631_));
NOR2X1 NOR2X1_24 ( .A(counter_32_), .B(counter_33_), .Y(_abc_4169_new_n632_));
NOR2X1 NOR2X1_25 ( .A(counter_30_), .B(counter_31_), .Y(_abc_4169_new_n633_));
NOR2X1 NOR2X1_26 ( .A(counter_20_), .B(counter_21_), .Y(_abc_4169_new_n637_));
NOR2X1 NOR2X1_27 ( .A(_abc_4169_new_n634_), .B(_abc_4169_new_n638_), .Y(_abc_4169_new_n639_));
NOR2X1 NOR2X1_28 ( .A(_abc_4169_new_n1035_), .B(_abc_4169_new_n607_), .Y(_abc_4169_new_n1036_));
NOR2X1 NOR2X1_29 ( .A(_abc_4169_new_n1212_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__1_));
NOR2X1 NOR2X1_3 ( .A(axi_bready), .B(axi_rready), .Y(_abc_4169_new_n568_));
NOR2X1 NOR2X1_30 ( .A(_abc_4169_new_n597_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__2_));
NOR2X1 NOR2X1_31 ( .A(_abc_4169_new_n611_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__3_));
NOR2X1 NOR2X1_32 ( .A(_abc_4169_new_n612_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__4_));
NOR2X1 NOR2X1_33 ( .A(_abc_4169_new_n1217_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__5_));
NOR2X1 NOR2X1_34 ( .A(_abc_4169_new_n1219_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__6_));
NOR2X1 NOR2X1_35 ( .A(_abc_4169_new_n627_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__7_));
NOR2X1 NOR2X1_36 ( .A(_abc_4169_new_n628_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__8_));
NOR2X1 NOR2X1_37 ( .A(_abc_4169_new_n1223_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__9_));
NOR2X1 NOR2X1_38 ( .A(_abc_4169_new_n1225_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__10_));
NOR2X1 NOR2X1_39 ( .A(_abc_4169_new_n1227_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__11_));
NOR2X1 NOR2X1_4 ( .A(we_clk), .B(_abc_4169_new_n574_), .Y(_abc_4169_new_n575_));
NOR2X1 NOR2X1_40 ( .A(_abc_4169_new_n1229_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__12_));
NOR2X1 NOR2X1_41 ( .A(_abc_4169_new_n1231_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__13_));
NOR2X1 NOR2X1_42 ( .A(_abc_4169_new_n1233_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__14_));
NOR2X1 NOR2X1_43 ( .A(_abc_4169_new_n1235_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__15_));
NOR2X1 NOR2X1_44 ( .A(_abc_4169_new_n1237_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__16_));
NOR2X1 NOR2X1_45 ( .A(_abc_4169_new_n1239_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__17_));
NOR2X1 NOR2X1_46 ( .A(_abc_4169_new_n1241_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__18_));
NOR2X1 NOR2X1_47 ( .A(_abc_4169_new_n635_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__19_));
NOR2X1 NOR2X1_48 ( .A(_abc_4169_new_n636_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__20_));
NOR2X1 NOR2X1_49 ( .A(_abc_4169_new_n1245_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__21_));
NOR2X1 NOR2X1_5 ( .A(state_7_), .B(state_5_), .Y(_abc_4169_new_n583_));
NOR2X1 NOR2X1_50 ( .A(_abc_4169_new_n1247_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__22_));
NOR2X1 NOR2X1_51 ( .A(_abc_4169_new_n1249_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__23_));
NOR2X1 NOR2X1_52 ( .A(_abc_4169_new_n1251_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__24_));
NOR2X1 NOR2X1_53 ( .A(_abc_4169_new_n1253_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__25_));
NOR2X1 NOR2X1_54 ( .A(_abc_4169_new_n1255_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__26_));
NOR2X1 NOR2X1_55 ( .A(_abc_4169_new_n1257_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__27_));
NOR2X1 NOR2X1_56 ( .A(_abc_4169_new_n1259_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__28_));
NOR2X1 NOR2X1_57 ( .A(_abc_4169_new_n1261_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__29_));
NOR2X1 NOR2X1_58 ( .A(_abc_4169_new_n1263_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__30_));
NOR2X1 NOR2X1_59 ( .A(_abc_4169_new_n1265_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__31_));
NOR2X1 NOR2X1_6 ( .A(state_1_), .B(state_4_), .Y(_abc_4169_new_n585_));
NOR2X1 NOR2X1_60 ( .A(_abc_4169_new_n1267_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__32_));
NOR2X1 NOR2X1_61 ( .A(_abc_4169_new_n1269_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__33_));
NOR2X1 NOR2X1_62 ( .A(_abc_4169_new_n1035_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__34_));
NOR2X1 NOR2X1_63 ( .A(_abc_4169_new_n1272_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__35_));
NOR2X1 NOR2X1_64 ( .A(_abc_4169_new_n1274_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__36_));
NOR2X1 NOR2X1_65 ( .A(_abc_4169_new_n1276_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__37_));
NOR2X1 NOR2X1_66 ( .A(_abc_4169_new_n1278_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__38_));
NOR2X1 NOR2X1_67 ( .A(_abc_4169_new_n1280_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__39_));
NOR2X1 NOR2X1_68 ( .A(_abc_4169_new_n1282_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__40_));
NOR2X1 NOR2X1_69 ( .A(_abc_4169_new_n1284_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__41_));
NOR2X1 NOR2X1_7 ( .A(_abc_4169_new_n581_), .B(_abc_4169_new_n586_), .Y(_abc_4169_new_n587_));
NOR2X1 NOR2X1_70 ( .A(_abc_4169_new_n1286_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__42_));
NOR2X1 NOR2X1_71 ( .A(_abc_4169_new_n1288_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__43_));
NOR2X1 NOR2X1_72 ( .A(_abc_4169_new_n1290_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__44_));
NOR2X1 NOR2X1_73 ( .A(_abc_4169_new_n1292_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__45_));
NOR2X1 NOR2X1_74 ( .A(_abc_4169_new_n1294_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__46_));
NOR2X1 NOR2X1_75 ( .A(_abc_4169_new_n1296_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__47_));
NOR2X1 NOR2X1_76 ( .A(_abc_4169_new_n1298_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__48_));
NOR2X1 NOR2X1_77 ( .A(_abc_4169_new_n1300_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__49_));
NOR2X1 NOR2X1_78 ( .A(_abc_4169_new_n1302_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__50_));
NOR2X1 NOR2X1_79 ( .A(_abc_4169_new_n1304_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__51_));
NOR2X1 NOR2X1_8 ( .A(re_clk), .B(_abc_4169_new_n572_), .Y(_abc_4169_new_n594_));
NOR2X1 NOR2X1_80 ( .A(_abc_4169_new_n1306_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__52_));
NOR2X1 NOR2X1_81 ( .A(_abc_4169_new_n1308_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__53_));
NOR2X1 NOR2X1_82 ( .A(_abc_4169_new_n1310_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__54_));
NOR2X1 NOR2X1_83 ( .A(_abc_4169_new_n1312_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__55_));
NOR2X1 NOR2X1_84 ( .A(_abc_4169_new_n1314_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__56_));
NOR2X1 NOR2X1_85 ( .A(_abc_4169_new_n1316_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__57_));
NOR2X1 NOR2X1_86 ( .A(_abc_4169_new_n1318_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__58_));
NOR2X1 NOR2X1_87 ( .A(_abc_4169_new_n1320_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__59_));
NOR2X1 NOR2X1_88 ( .A(_abc_4169_new_n1322_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__60_));
NOR2X1 NOR2X1_89 ( .A(_abc_4169_new_n1324_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__61_));
NOR2X1 NOR2X1_9 ( .A(_abc_4169_new_n564_), .B(_abc_4169_new_n595_), .Y(_abc_2903_auto_fsm_map_cc_170_map_fsm_402_5_));
NOR2X1 NOR2X1_90 ( .A(_abc_4169_new_n1326_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__62_));
NOR2X1 NOR2X1_91 ( .A(_abc_4169_new_n1328_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__63_));
NOR2X1 NOR2X1_92 ( .A(_abc_4169_new_n1330_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__64_));
NOR2X1 NOR2X1_93 ( .A(_abc_4169_new_n1332_), .B(_0counter_65_0__0_), .Y(_0counter_65_0__65_));
OAI21X1 OAI21X1_1 ( .A(axi_bvalid), .B(_abc_4169_new_n558_), .C(_abc_4169_new_n559_), .Y(_abc_4169_new_n560_));
OAI21X1 OAI21X1_10 ( .A(_abc_4169_new_n653_), .B(_abc_4169_new_n655_), .C(RST), .Y(_abc_4169_new_n656_));
OAI21X1 OAI21X1_100 ( .A(sft_reg_25_), .B(_abc_4169_new_n938_), .C(RST), .Y(_abc_4169_new_n1017_));
OAI21X1 OAI21X1_101 ( .A(sft_reg_26_), .B(_abc_4169_new_n938_), .C(RST), .Y(_abc_4169_new_n1020_));
OAI21X1 OAI21X1_102 ( .A(sft_reg_27_), .B(_abc_4169_new_n938_), .C(RST), .Y(_abc_4169_new_n1023_));
OAI21X1 OAI21X1_103 ( .A(sft_reg_28_), .B(_abc_4169_new_n938_), .C(RST), .Y(_abc_4169_new_n1026_));
OAI21X1 OAI21X1_104 ( .A(sft_reg_29_), .B(_abc_4169_new_n938_), .C(RST), .Y(_abc_4169_new_n1029_));
OAI21X1 OAI21X1_105 ( .A(sft_reg_30_), .B(_abc_4169_new_n938_), .C(RST), .Y(_abc_4169_new_n1032_));
OAI21X1 OAI21X1_106 ( .A(DATA), .B(_abc_4169_new_n1037_), .C(RST), .Y(_abc_4169_new_n1038_));
OAI21X1 OAI21X1_107 ( .A(sft_reg_0_), .B(_abc_4169_new_n1037_), .C(RST), .Y(_abc_4169_new_n1041_));
OAI21X1 OAI21X1_108 ( .A(sft_reg_1_), .B(_abc_4169_new_n1037_), .C(RST), .Y(_abc_4169_new_n1044_));
OAI21X1 OAI21X1_109 ( .A(sft_reg_2_), .B(_abc_4169_new_n1037_), .C(RST), .Y(_abc_4169_new_n1047_));
OAI21X1 OAI21X1_11 ( .A(_abc_4169_new_n661_), .B(_abc_4169_new_n598_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n662_));
OAI21X1 OAI21X1_110 ( .A(sft_reg_3_), .B(_abc_4169_new_n1037_), .C(RST), .Y(_abc_4169_new_n1050_));
OAI21X1 OAI21X1_111 ( .A(sft_reg_4_), .B(_abc_4169_new_n1037_), .C(RST), .Y(_abc_4169_new_n1053_));
OAI21X1 OAI21X1_112 ( .A(sft_reg_5_), .B(_abc_4169_new_n1037_), .C(RST), .Y(_abc_4169_new_n1056_));
OAI21X1 OAI21X1_113 ( .A(sft_reg_6_), .B(_abc_4169_new_n1037_), .C(RST), .Y(_abc_4169_new_n1059_));
OAI21X1 OAI21X1_114 ( .A(sft_reg_7_), .B(_abc_4169_new_n1037_), .C(RST), .Y(_abc_4169_new_n1062_));
OAI21X1 OAI21X1_115 ( .A(sft_reg_8_), .B(_abc_4169_new_n1037_), .C(RST), .Y(_abc_4169_new_n1065_));
OAI21X1 OAI21X1_116 ( .A(sft_reg_9_), .B(_abc_4169_new_n1037_), .C(RST), .Y(_abc_4169_new_n1068_));
OAI21X1 OAI21X1_117 ( .A(sft_reg_10_), .B(_abc_4169_new_n1037_), .C(RST), .Y(_abc_4169_new_n1071_));
OAI21X1 OAI21X1_118 ( .A(sft_reg_11_), .B(_abc_4169_new_n1037_), .C(RST), .Y(_abc_4169_new_n1074_));
OAI21X1 OAI21X1_119 ( .A(sft_reg_12_), .B(_abc_4169_new_n1037_), .C(RST), .Y(_abc_4169_new_n1077_));
OAI21X1 OAI21X1_12 ( .A(_abc_4169_new_n660_), .B(_abc_4169_new_n662_), .C(RST), .Y(_abc_4169_new_n663_));
OAI21X1 OAI21X1_120 ( .A(sft_reg_13_), .B(_abc_4169_new_n1037_), .C(RST), .Y(_abc_4169_new_n1080_));
OAI21X1 OAI21X1_121 ( .A(sft_reg_14_), .B(_abc_4169_new_n1037_), .C(RST), .Y(_abc_4169_new_n1083_));
OAI21X1 OAI21X1_122 ( .A(sft_reg_15_), .B(_abc_4169_new_n1037_), .C(RST), .Y(_abc_4169_new_n1086_));
OAI21X1 OAI21X1_123 ( .A(sft_reg_16_), .B(_abc_4169_new_n1037_), .C(RST), .Y(_abc_4169_new_n1089_));
OAI21X1 OAI21X1_124 ( .A(sft_reg_17_), .B(_abc_4169_new_n1037_), .C(RST), .Y(_abc_4169_new_n1092_));
OAI21X1 OAI21X1_125 ( .A(sft_reg_18_), .B(_abc_4169_new_n1037_), .C(RST), .Y(_abc_4169_new_n1095_));
OAI21X1 OAI21X1_126 ( .A(sft_reg_19_), .B(_abc_4169_new_n1037_), .C(RST), .Y(_abc_4169_new_n1098_));
OAI21X1 OAI21X1_127 ( .A(sft_reg_20_), .B(_abc_4169_new_n1037_), .C(RST), .Y(_abc_4169_new_n1101_));
OAI21X1 OAI21X1_128 ( .A(sft_reg_21_), .B(_abc_4169_new_n1037_), .C(RST), .Y(_abc_4169_new_n1104_));
OAI21X1 OAI21X1_129 ( .A(sft_reg_22_), .B(_abc_4169_new_n1037_), .C(RST), .Y(_abc_4169_new_n1107_));
OAI21X1 OAI21X1_13 ( .A(_abc_4169_new_n667_), .B(_abc_4169_new_n598_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n668_));
OAI21X1 OAI21X1_130 ( .A(sft_reg_23_), .B(_abc_4169_new_n1037_), .C(RST), .Y(_abc_4169_new_n1110_));
OAI21X1 OAI21X1_131 ( .A(sft_reg_24_), .B(_abc_4169_new_n1037_), .C(RST), .Y(_abc_4169_new_n1113_));
OAI21X1 OAI21X1_132 ( .A(sft_reg_25_), .B(_abc_4169_new_n1037_), .C(RST), .Y(_abc_4169_new_n1116_));
OAI21X1 OAI21X1_133 ( .A(sft_reg_26_), .B(_abc_4169_new_n1037_), .C(RST), .Y(_abc_4169_new_n1119_));
OAI21X1 OAI21X1_134 ( .A(sft_reg_27_), .B(_abc_4169_new_n1037_), .C(RST), .Y(_abc_4169_new_n1122_));
OAI21X1 OAI21X1_135 ( .A(sft_reg_28_), .B(_abc_4169_new_n1037_), .C(RST), .Y(_abc_4169_new_n1125_));
OAI21X1 OAI21X1_136 ( .A(sft_reg_29_), .B(_abc_4169_new_n1037_), .C(RST), .Y(_abc_4169_new_n1128_));
OAI21X1 OAI21X1_137 ( .A(sft_reg_30_), .B(_abc_4169_new_n1037_), .C(RST), .Y(_abc_4169_new_n1131_));
OAI21X1 OAI21X1_138 ( .A(DATA), .B(CEB), .C(RST), .Y(_abc_4169_new_n1134_));
OAI21X1 OAI21X1_139 ( .A(sft_reg_1_), .B(_abc_4169_new_n937_), .C(RST), .Y(_abc_4169_new_n1136_));
OAI21X1 OAI21X1_14 ( .A(_abc_4169_new_n673_), .B(_abc_4169_new_n598_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n674_));
OAI21X1 OAI21X1_140 ( .A(CEB), .B(sft_reg_1_), .C(RST), .Y(_abc_4169_new_n1139_));
OAI21X1 OAI21X1_141 ( .A(sft_reg_3_), .B(_abc_4169_new_n937_), .C(RST), .Y(_abc_4169_new_n1141_));
OAI21X1 OAI21X1_142 ( .A(CEB), .B(sft_reg_3_), .C(RST), .Y(_abc_4169_new_n1144_));
OAI21X1 OAI21X1_143 ( .A(sft_reg_5_), .B(_abc_4169_new_n937_), .C(RST), .Y(_abc_4169_new_n1146_));
OAI21X1 OAI21X1_144 ( .A(CEB), .B(sft_reg_5_), .C(RST), .Y(_abc_4169_new_n1149_));
OAI21X1 OAI21X1_145 ( .A(sft_reg_7_), .B(_abc_4169_new_n937_), .C(RST), .Y(_abc_4169_new_n1151_));
OAI21X1 OAI21X1_146 ( .A(CEB), .B(sft_reg_7_), .C(RST), .Y(_abc_4169_new_n1154_));
OAI21X1 OAI21X1_147 ( .A(sft_reg_9_), .B(_abc_4169_new_n937_), .C(RST), .Y(_abc_4169_new_n1156_));
OAI21X1 OAI21X1_148 ( .A(CEB), .B(sft_reg_9_), .C(RST), .Y(_abc_4169_new_n1159_));
OAI21X1 OAI21X1_149 ( .A(sft_reg_11_), .B(_abc_4169_new_n937_), .C(RST), .Y(_abc_4169_new_n1161_));
OAI21X1 OAI21X1_15 ( .A(_abc_4169_new_n679_), .B(_abc_4169_new_n598_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n680_));
OAI21X1 OAI21X1_150 ( .A(CEB), .B(sft_reg_11_), .C(RST), .Y(_abc_4169_new_n1164_));
OAI21X1 OAI21X1_151 ( .A(sft_reg_13_), .B(_abc_4169_new_n937_), .C(RST), .Y(_abc_4169_new_n1166_));
OAI21X1 OAI21X1_152 ( .A(CEB), .B(sft_reg_13_), .C(RST), .Y(_abc_4169_new_n1169_));
OAI21X1 OAI21X1_153 ( .A(sft_reg_15_), .B(_abc_4169_new_n937_), .C(RST), .Y(_abc_4169_new_n1171_));
OAI21X1 OAI21X1_154 ( .A(CEB), .B(sft_reg_15_), .C(RST), .Y(_abc_4169_new_n1174_));
OAI21X1 OAI21X1_155 ( .A(sft_reg_17_), .B(_abc_4169_new_n937_), .C(RST), .Y(_abc_4169_new_n1176_));
OAI21X1 OAI21X1_156 ( .A(CEB), .B(sft_reg_17_), .C(RST), .Y(_abc_4169_new_n1179_));
OAI21X1 OAI21X1_157 ( .A(sft_reg_19_), .B(_abc_4169_new_n937_), .C(RST), .Y(_abc_4169_new_n1181_));
OAI21X1 OAI21X1_158 ( .A(CEB), .B(sft_reg_19_), .C(RST), .Y(_abc_4169_new_n1184_));
OAI21X1 OAI21X1_159 ( .A(sft_reg_21_), .B(_abc_4169_new_n937_), .C(RST), .Y(_abc_4169_new_n1186_));
OAI21X1 OAI21X1_16 ( .A(_abc_4169_new_n685_), .B(_abc_4169_new_n598_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n686_));
OAI21X1 OAI21X1_160 ( .A(CEB), .B(sft_reg_21_), .C(RST), .Y(_abc_4169_new_n1189_));
OAI21X1 OAI21X1_161 ( .A(sft_reg_23_), .B(_abc_4169_new_n937_), .C(RST), .Y(_abc_4169_new_n1191_));
OAI21X1 OAI21X1_162 ( .A(CEB), .B(sft_reg_23_), .C(RST), .Y(_abc_4169_new_n1194_));
OAI21X1 OAI21X1_163 ( .A(sft_reg_25_), .B(_abc_4169_new_n937_), .C(RST), .Y(_abc_4169_new_n1196_));
OAI21X1 OAI21X1_164 ( .A(CEB), .B(sft_reg_25_), .C(RST), .Y(_abc_4169_new_n1199_));
OAI21X1 OAI21X1_165 ( .A(sft_reg_27_), .B(_abc_4169_new_n937_), .C(RST), .Y(_abc_4169_new_n1201_));
OAI21X1 OAI21X1_166 ( .A(CEB), .B(sft_reg_27_), .C(RST), .Y(_abc_4169_new_n1204_));
OAI21X1 OAI21X1_167 ( .A(sft_reg_29_), .B(_abc_4169_new_n937_), .C(RST), .Y(_abc_4169_new_n1206_));
OAI21X1 OAI21X1_168 ( .A(CEB), .B(sft_reg_29_), .C(RST), .Y(_abc_4169_new_n1209_));
OAI21X1 OAI21X1_169 ( .A(DATA), .B(_abc_4169_new_n1336_), .C(RST), .Y(_abc_4169_new_n1337_));
OAI21X1 OAI21X1_17 ( .A(_abc_4169_new_n691_), .B(_abc_4169_new_n598_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n692_));
OAI21X1 OAI21X1_170 ( .A(_abc_4169_new_n597_), .B(_abc_4169_new_n1340_), .C(RST), .Y(_abc_4169_new_n1341_));
OAI21X1 OAI21X1_171 ( .A(_abc_4169_new_n1212_), .B(_abc_4169_new_n1340_), .C(RST), .Y(_abc_4169_new_n1344_));
OAI21X1 OAI21X1_18 ( .A(_abc_4169_new_n697_), .B(_abc_4169_new_n598_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n698_));
OAI21X1 OAI21X1_19 ( .A(_abc_4169_new_n703_), .B(_abc_4169_new_n598_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n704_));
OAI21X1 OAI21X1_2 ( .A(re_clk), .B(_abc_4169_new_n572_), .C(RST), .Y(_abc_4169_new_n573_));
OAI21X1 OAI21X1_20 ( .A(_abc_4169_new_n709_), .B(_abc_4169_new_n598_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n710_));
OAI21X1 OAI21X1_21 ( .A(_abc_4169_new_n715_), .B(_abc_4169_new_n598_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n716_));
OAI21X1 OAI21X1_22 ( .A(_abc_4169_new_n721_), .B(_abc_4169_new_n598_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n722_));
OAI21X1 OAI21X1_23 ( .A(_abc_4169_new_n727_), .B(_abc_4169_new_n598_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n728_));
OAI21X1 OAI21X1_24 ( .A(_abc_4169_new_n733_), .B(_abc_4169_new_n598_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n734_));
OAI21X1 OAI21X1_25 ( .A(_abc_4169_new_n739_), .B(_abc_4169_new_n598_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n740_));
OAI21X1 OAI21X1_26 ( .A(_abc_4169_new_n745_), .B(_abc_4169_new_n598_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n746_));
OAI21X1 OAI21X1_27 ( .A(_abc_4169_new_n751_), .B(_abc_4169_new_n598_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n752_));
OAI21X1 OAI21X1_28 ( .A(_abc_4169_new_n757_), .B(_abc_4169_new_n598_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n758_));
OAI21X1 OAI21X1_29 ( .A(_abc_4169_new_n763_), .B(_abc_4169_new_n598_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n764_));
OAI21X1 OAI21X1_3 ( .A(we_clk), .B(_abc_4169_new_n574_), .C(state_0_), .Y(_abc_4169_new_n589_));
OAI21X1 OAI21X1_30 ( .A(_abc_4169_new_n769_), .B(_abc_4169_new_n598_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n770_));
OAI21X1 OAI21X1_31 ( .A(_abc_4169_new_n775_), .B(_abc_4169_new_n598_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n776_));
OAI21X1 OAI21X1_32 ( .A(_abc_4169_new_n781_), .B(_abc_4169_new_n598_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n782_));
OAI21X1 OAI21X1_33 ( .A(_abc_4169_new_n787_), .B(_abc_4169_new_n598_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n788_));
OAI21X1 OAI21X1_34 ( .A(_abc_4169_new_n793_), .B(_abc_4169_new_n598_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n794_));
OAI21X1 OAI21X1_35 ( .A(_abc_4169_new_n799_), .B(_abc_4169_new_n598_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n800_));
OAI21X1 OAI21X1_36 ( .A(_abc_4169_new_n805_), .B(_abc_4169_new_n598_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n806_));
OAI21X1 OAI21X1_37 ( .A(_abc_4169_new_n811_), .B(_abc_4169_new_n598_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n812_));
OAI21X1 OAI21X1_38 ( .A(_abc_4169_new_n817_), .B(_abc_4169_new_n598_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n818_));
OAI21X1 OAI21X1_39 ( .A(_abc_4169_new_n823_), .B(_abc_4169_new_n598_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n824_));
OAI21X1 OAI21X1_4 ( .A(_abc_4169_new_n573_), .B(_abc_4169_new_n589_), .C(_abc_4169_new_n591_), .Y(_abc_2903_auto_fsm_map_cc_170_map_fsm_402_0_));
OAI21X1 OAI21X1_40 ( .A(_abc_4169_new_n829_), .B(_abc_4169_new_n598_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n830_));
OAI21X1 OAI21X1_41 ( .A(_abc_4169_new_n835_), .B(_abc_4169_new_n598_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n836_));
OAI21X1 OAI21X1_42 ( .A(\axi_rdata[0] ), .B(_abc_4169_new_n839_), .C(RST), .Y(_abc_4169_new_n841_));
OAI21X1 OAI21X1_43 ( .A(\axi_rdata[1] ), .B(_abc_4169_new_n839_), .C(RST), .Y(_abc_4169_new_n844_));
OAI21X1 OAI21X1_44 ( .A(\axi_rdata[2] ), .B(_abc_4169_new_n839_), .C(RST), .Y(_abc_4169_new_n847_));
OAI21X1 OAI21X1_45 ( .A(\axi_rdata[3] ), .B(_abc_4169_new_n839_), .C(RST), .Y(_abc_4169_new_n850_));
OAI21X1 OAI21X1_46 ( .A(\axi_rdata[4] ), .B(_abc_4169_new_n839_), .C(RST), .Y(_abc_4169_new_n853_));
OAI21X1 OAI21X1_47 ( .A(\axi_rdata[5] ), .B(_abc_4169_new_n839_), .C(RST), .Y(_abc_4169_new_n856_));
OAI21X1 OAI21X1_48 ( .A(\axi_rdata[6] ), .B(_abc_4169_new_n839_), .C(RST), .Y(_abc_4169_new_n859_));
OAI21X1 OAI21X1_49 ( .A(\axi_rdata[7] ), .B(_abc_4169_new_n839_), .C(RST), .Y(_abc_4169_new_n862_));
OAI21X1 OAI21X1_5 ( .A(_abc_4169_new_n597_), .B(_abc_4169_new_n600_), .C(_abc_4169_new_n598_), .Y(_abc_4169_new_n601_));
OAI21X1 OAI21X1_50 ( .A(\axi_rdata[8] ), .B(_abc_4169_new_n839_), .C(RST), .Y(_abc_4169_new_n865_));
OAI21X1 OAI21X1_51 ( .A(\axi_rdata[9] ), .B(_abc_4169_new_n839_), .C(RST), .Y(_abc_4169_new_n868_));
OAI21X1 OAI21X1_52 ( .A(\axi_rdata[10] ), .B(_abc_4169_new_n839_), .C(RST), .Y(_abc_4169_new_n871_));
OAI21X1 OAI21X1_53 ( .A(\axi_rdata[11] ), .B(_abc_4169_new_n839_), .C(RST), .Y(_abc_4169_new_n874_));
OAI21X1 OAI21X1_54 ( .A(\axi_rdata[12] ), .B(_abc_4169_new_n839_), .C(RST), .Y(_abc_4169_new_n877_));
OAI21X1 OAI21X1_55 ( .A(\axi_rdata[13] ), .B(_abc_4169_new_n839_), .C(RST), .Y(_abc_4169_new_n880_));
OAI21X1 OAI21X1_56 ( .A(\axi_rdata[14] ), .B(_abc_4169_new_n839_), .C(RST), .Y(_abc_4169_new_n883_));
OAI21X1 OAI21X1_57 ( .A(\axi_rdata[15] ), .B(_abc_4169_new_n839_), .C(RST), .Y(_abc_4169_new_n886_));
OAI21X1 OAI21X1_58 ( .A(\axi_rdata[16] ), .B(_abc_4169_new_n839_), .C(RST), .Y(_abc_4169_new_n889_));
OAI21X1 OAI21X1_59 ( .A(\axi_rdata[17] ), .B(_abc_4169_new_n839_), .C(RST), .Y(_abc_4169_new_n892_));
OAI21X1 OAI21X1_6 ( .A(_abc_4169_new_n623_), .B(_abc_4169_new_n640_), .C(_abc_4169_new_n607_), .Y(_abc_4169_new_n641_));
OAI21X1 OAI21X1_60 ( .A(\axi_rdata[18] ), .B(_abc_4169_new_n839_), .C(RST), .Y(_abc_4169_new_n895_));
OAI21X1 OAI21X1_61 ( .A(\axi_rdata[19] ), .B(_abc_4169_new_n839_), .C(RST), .Y(_abc_4169_new_n898_));
OAI21X1 OAI21X1_62 ( .A(\axi_rdata[20] ), .B(_abc_4169_new_n839_), .C(RST), .Y(_abc_4169_new_n901_));
OAI21X1 OAI21X1_63 ( .A(\axi_rdata[21] ), .B(_abc_4169_new_n839_), .C(RST), .Y(_abc_4169_new_n904_));
OAI21X1 OAI21X1_64 ( .A(\axi_rdata[22] ), .B(_abc_4169_new_n839_), .C(RST), .Y(_abc_4169_new_n907_));
OAI21X1 OAI21X1_65 ( .A(\axi_rdata[23] ), .B(_abc_4169_new_n839_), .C(RST), .Y(_abc_4169_new_n910_));
OAI21X1 OAI21X1_66 ( .A(\axi_rdata[24] ), .B(_abc_4169_new_n839_), .C(RST), .Y(_abc_4169_new_n913_));
OAI21X1 OAI21X1_67 ( .A(\axi_rdata[25] ), .B(_abc_4169_new_n839_), .C(RST), .Y(_abc_4169_new_n916_));
OAI21X1 OAI21X1_68 ( .A(\axi_rdata[26] ), .B(_abc_4169_new_n839_), .C(RST), .Y(_abc_4169_new_n919_));
OAI21X1 OAI21X1_69 ( .A(\axi_rdata[27] ), .B(_abc_4169_new_n839_), .C(RST), .Y(_abc_4169_new_n922_));
OAI21X1 OAI21X1_7 ( .A(_abc_4169_new_n644_), .B(_abc_4169_new_n598_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n645_));
OAI21X1 OAI21X1_70 ( .A(\axi_rdata[28] ), .B(_abc_4169_new_n839_), .C(RST), .Y(_abc_4169_new_n925_));
OAI21X1 OAI21X1_71 ( .A(\axi_rdata[29] ), .B(_abc_4169_new_n839_), .C(RST), .Y(_abc_4169_new_n928_));
OAI21X1 OAI21X1_72 ( .A(\axi_rdata[30] ), .B(_abc_4169_new_n839_), .C(RST), .Y(_abc_4169_new_n931_));
OAI21X1 OAI21X1_73 ( .A(\axi_rdata[31] ), .B(_abc_4169_new_n839_), .C(RST), .Y(_abc_4169_new_n934_));
OAI21X1 OAI21X1_74 ( .A(DATA), .B(_abc_4169_new_n938_), .C(RST), .Y(_abc_4169_new_n939_));
OAI21X1 OAI21X1_75 ( .A(sft_reg_0_), .B(_abc_4169_new_n938_), .C(RST), .Y(_abc_4169_new_n942_));
OAI21X1 OAI21X1_76 ( .A(sft_reg_1_), .B(_abc_4169_new_n938_), .C(RST), .Y(_abc_4169_new_n945_));
OAI21X1 OAI21X1_77 ( .A(sft_reg_2_), .B(_abc_4169_new_n938_), .C(RST), .Y(_abc_4169_new_n948_));
OAI21X1 OAI21X1_78 ( .A(sft_reg_3_), .B(_abc_4169_new_n938_), .C(RST), .Y(_abc_4169_new_n951_));
OAI21X1 OAI21X1_79 ( .A(sft_reg_4_), .B(_abc_4169_new_n938_), .C(RST), .Y(_abc_4169_new_n954_));
OAI21X1 OAI21X1_8 ( .A(_abc_4169_new_n643_), .B(_abc_4169_new_n645_), .C(RST), .Y(_abc_4169_new_n646_));
OAI21X1 OAI21X1_80 ( .A(sft_reg_5_), .B(_abc_4169_new_n938_), .C(RST), .Y(_abc_4169_new_n957_));
OAI21X1 OAI21X1_81 ( .A(sft_reg_6_), .B(_abc_4169_new_n938_), .C(RST), .Y(_abc_4169_new_n960_));
OAI21X1 OAI21X1_82 ( .A(sft_reg_7_), .B(_abc_4169_new_n938_), .C(RST), .Y(_abc_4169_new_n963_));
OAI21X1 OAI21X1_83 ( .A(sft_reg_8_), .B(_abc_4169_new_n938_), .C(RST), .Y(_abc_4169_new_n966_));
OAI21X1 OAI21X1_84 ( .A(sft_reg_9_), .B(_abc_4169_new_n938_), .C(RST), .Y(_abc_4169_new_n969_));
OAI21X1 OAI21X1_85 ( .A(sft_reg_10_), .B(_abc_4169_new_n938_), .C(RST), .Y(_abc_4169_new_n972_));
OAI21X1 OAI21X1_86 ( .A(sft_reg_11_), .B(_abc_4169_new_n938_), .C(RST), .Y(_abc_4169_new_n975_));
OAI21X1 OAI21X1_87 ( .A(sft_reg_12_), .B(_abc_4169_new_n938_), .C(RST), .Y(_abc_4169_new_n978_));
OAI21X1 OAI21X1_88 ( .A(sft_reg_13_), .B(_abc_4169_new_n938_), .C(RST), .Y(_abc_4169_new_n981_));
OAI21X1 OAI21X1_89 ( .A(sft_reg_14_), .B(_abc_4169_new_n938_), .C(RST), .Y(_abc_4169_new_n984_));
OAI21X1 OAI21X1_9 ( .A(_abc_4169_new_n654_), .B(_abc_4169_new_n598_), .C(_abc_4169_new_n601_), .Y(_abc_4169_new_n655_));
OAI21X1 OAI21X1_90 ( .A(sft_reg_15_), .B(_abc_4169_new_n938_), .C(RST), .Y(_abc_4169_new_n987_));
OAI21X1 OAI21X1_91 ( .A(sft_reg_16_), .B(_abc_4169_new_n938_), .C(RST), .Y(_abc_4169_new_n990_));
OAI21X1 OAI21X1_92 ( .A(sft_reg_17_), .B(_abc_4169_new_n938_), .C(RST), .Y(_abc_4169_new_n993_));
OAI21X1 OAI21X1_93 ( .A(sft_reg_18_), .B(_abc_4169_new_n938_), .C(RST), .Y(_abc_4169_new_n996_));
OAI21X1 OAI21X1_94 ( .A(sft_reg_19_), .B(_abc_4169_new_n938_), .C(RST), .Y(_abc_4169_new_n999_));
OAI21X1 OAI21X1_95 ( .A(sft_reg_20_), .B(_abc_4169_new_n938_), .C(RST), .Y(_abc_4169_new_n1002_));
OAI21X1 OAI21X1_96 ( .A(sft_reg_21_), .B(_abc_4169_new_n938_), .C(RST), .Y(_abc_4169_new_n1005_));
OAI21X1 OAI21X1_97 ( .A(sft_reg_22_), .B(_abc_4169_new_n938_), .C(RST), .Y(_abc_4169_new_n1008_));
OAI21X1 OAI21X1_98 ( .A(sft_reg_23_), .B(_abc_4169_new_n938_), .C(RST), .Y(_abc_4169_new_n1011_));
OAI21X1 OAI21X1_99 ( .A(sft_reg_24_), .B(_abc_4169_new_n938_), .C(RST), .Y(_abc_4169_new_n1014_));
OAI22X1 OAI22X1_1 ( .A(axi_arready), .B(_abc_4169_new_n571_), .C(_abc_4169_new_n573_), .D(_abc_4169_new_n576_), .Y(_abc_2903_auto_fsm_map_cc_170_map_fsm_402_6_));
OAI22X1 OAI22X1_2 ( .A(_abc_4169_new_n578_), .B(_abc_4169_new_n571_), .C(axi_rvalid), .D(_abc_4169_new_n579_), .Y(_abc_2903_auto_fsm_map_cc_170_map_fsm_402_4_));
OR2X2 OR2X2_1 ( .A(axi_rready), .B(state_6_), .Y(_abc_4169_new_n581_));
OR2X2 OR2X2_2 ( .A(_abc_4169_new_n581_), .B(state_4_), .Y(axi_arvalid));
OR2X2 OR2X2_3 ( .A(DATA), .B(CEB), .Y(_abc_4169_new_n1340_));

assign \axi_arprot[0]  = 1'h0;
assign \axi_arprot[1]  = 1'h0;
assign \axi_arprot[2]  = 1'h0;
assign \axi_awprot[0]  = 1'h0;
assign \axi_awprot[1]  = 1'h0;
assign \axi_awprot[2]  = 1'h0;
assign \axi_wstrb[0]  = 1'h1;
assign \axi_wstrb[1]  = 1'h1;
assign \axi_wstrb[2]  = 1'h1;
assign \axi_wstrb[3]  = 1'h1;

endmodule