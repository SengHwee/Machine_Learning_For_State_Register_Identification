module sha1_core(clk, reset_n, init, next, \block[0] , \block[1] , \block[2] , \block[3] , \block[4] , \block[5] , \block[6] , \block[7] , \block[8] , \block[9] , \block[10] , \block[11] , \block[12] , \block[13] , \block[14] , \block[15] , \block[16] , \block[17] , \block[18] , \block[19] , \block[20] , \block[21] , \block[22] , \block[23] , \block[24] , \block[25] , \block[26] , \block[27] , \block[28] , \block[29] , \block[30] , \block[31] , \block[32] , \block[33] , \block[34] , \block[35] , \block[36] , \block[37] , \block[38] , \block[39] , \block[40] , \block[41] , \block[42] , \block[43] , \block[44] , \block[45] , \block[46] , \block[47] , \block[48] , \block[49] , \block[50] , \block[51] , \block[52] , \block[53] , \block[54] , \block[55] , \block[56] , \block[57] , \block[58] , \block[59] , \block[60] , \block[61] , \block[62] , \block[63] , \block[64] , \block[65] , \block[66] , \block[67] , \block[68] , \block[69] , \block[70] , \block[71] , \block[72] , \block[73] , \block[74] , \block[75] , \block[76] , \block[77] , \block[78] , \block[79] , \block[80] , \block[81] , \block[82] , \block[83] , \block[84] , \block[85] , \block[86] , \block[87] , \block[88] , \block[89] , \block[90] , \block[91] , \block[92] , \block[93] , \block[94] , \block[95] , \block[96] , \block[97] , \block[98] , \block[99] , \block[100] , \block[101] , \block[102] , \block[103] , \block[104] , \block[105] , \block[106] , \block[107] , \block[108] , \block[109] , \block[110] , \block[111] , \block[112] , \block[113] , \block[114] , \block[115] , \block[116] , \block[117] , \block[118] , \block[119] , \block[120] , \block[121] , \block[122] , \block[123] , \block[124] , \block[125] , \block[126] , \block[127] , \block[128] , \block[129] , \block[130] , \block[131] , \block[132] , \block[133] , \block[134] , \block[135] , \block[136] , \block[137] , \block[138] , \block[139] , \block[140] , \block[141] , \block[142] , \block[143] , \block[144] , \block[145] , \block[146] , \block[147] , \block[148] , \block[149] , \block[150] , \block[151] , \block[152] , \block[153] , \block[154] , \block[155] , \block[156] , \block[157] , \block[158] , \block[159] , \block[160] , \block[161] , \block[162] , \block[163] , \block[164] , \block[165] , \block[166] , \block[167] , \block[168] , \block[169] , \block[170] , \block[171] , \block[172] , \block[173] , \block[174] , \block[175] , \block[176] , \block[177] , \block[178] , \block[179] , \block[180] , \block[181] , \block[182] , \block[183] , \block[184] , \block[185] , \block[186] , \block[187] , \block[188] , \block[189] , \block[190] , \block[191] , \block[192] , \block[193] , \block[194] , \block[195] , \block[196] , \block[197] , \block[198] , \block[199] , \block[200] , \block[201] , \block[202] , \block[203] , \block[204] , \block[205] , \block[206] , \block[207] , \block[208] , \block[209] , \block[210] , \block[211] , \block[212] , \block[213] , \block[214] , \block[215] , \block[216] , \block[217] , \block[218] , \block[219] , \block[220] , \block[221] , \block[222] , \block[223] , \block[224] , \block[225] , \block[226] , \block[227] , \block[228] , \block[229] , \block[230] , \block[231] , \block[232] , \block[233] , \block[234] , \block[235] , \block[236] , \block[237] , \block[238] , \block[239] , \block[240] , \block[241] , \block[242] , \block[243] , \block[244] , \block[245] , \block[246] , \block[247] , \block[248] , \block[249] , \block[250] , \block[251] , \block[252] , \block[253] , \block[254] , \block[255] , \block[256] , \block[257] , \block[258] , \block[259] , \block[260] , \block[261] , \block[262] , \block[263] , \block[264] , \block[265] , \block[266] , \block[267] , \block[268] , \block[269] , \block[270] , \block[271] , \block[272] , \block[273] , \block[274] , \block[275] , \block[276] , \block[277] , \block[278] , \block[279] , \block[280] , \block[281] , \block[282] , \block[283] , \block[284] , \block[285] , \block[286] , \block[287] , \block[288] , \block[289] , \block[290] , \block[291] , \block[292] , \block[293] , \block[294] , \block[295] , \block[296] , \block[297] , \block[298] , \block[299] , \block[300] , \block[301] , \block[302] , \block[303] , \block[304] , \block[305] , \block[306] , \block[307] , \block[308] , \block[309] , \block[310] , \block[311] , \block[312] , \block[313] , \block[314] , \block[315] , \block[316] , \block[317] , \block[318] , \block[319] , \block[320] , \block[321] , \block[322] , \block[323] , \block[324] , \block[325] , \block[326] , \block[327] , \block[328] , \block[329] , \block[330] , \block[331] , \block[332] , \block[333] , \block[334] , \block[335] , \block[336] , \block[337] , \block[338] , \block[339] , \block[340] , \block[341] , \block[342] , \block[343] , \block[344] , \block[345] , \block[346] , \block[347] , \block[348] , \block[349] , \block[350] , \block[351] , \block[352] , \block[353] , \block[354] , \block[355] , \block[356] , \block[357] , \block[358] , \block[359] , \block[360] , \block[361] , \block[362] , \block[363] , \block[364] , \block[365] , \block[366] , \block[367] , \block[368] , \block[369] , \block[370] , \block[371] , \block[372] , \block[373] , \block[374] , \block[375] , \block[376] , \block[377] , \block[378] , \block[379] , \block[380] , \block[381] , \block[382] , \block[383] , \block[384] , \block[385] , \block[386] , \block[387] , \block[388] , \block[389] , \block[390] , \block[391] , \block[392] , \block[393] , \block[394] , \block[395] , \block[396] , \block[397] , \block[398] , \block[399] , \block[400] , \block[401] , \block[402] , \block[403] , \block[404] , \block[405] , \block[406] , \block[407] , \block[408] , \block[409] , \block[410] , \block[411] , \block[412] , \block[413] , \block[414] , \block[415] , \block[416] , \block[417] , \block[418] , \block[419] , \block[420] , \block[421] , \block[422] , \block[423] , \block[424] , \block[425] , \block[426] , \block[427] , \block[428] , \block[429] , \block[430] , \block[431] , \block[432] , \block[433] , \block[434] , \block[435] , \block[436] , \block[437] , \block[438] , \block[439] , \block[440] , \block[441] , \block[442] , \block[443] , \block[444] , \block[445] , \block[446] , \block[447] , \block[448] , \block[449] , \block[450] , \block[451] , \block[452] , \block[453] , \block[454] , \block[455] , \block[456] , \block[457] , \block[458] , \block[459] , \block[460] , \block[461] , \block[462] , \block[463] , \block[464] , \block[465] , \block[466] , \block[467] , \block[468] , \block[469] , \block[470] , \block[471] , \block[472] , \block[473] , \block[474] , \block[475] , \block[476] , \block[477] , \block[478] , \block[479] , \block[480] , \block[481] , \block[482] , \block[483] , \block[484] , \block[485] , \block[486] , \block[487] , \block[488] , \block[489] , \block[490] , \block[491] , \block[492] , \block[493] , \block[494] , \block[495] , \block[496] , \block[497] , \block[498] , \block[499] , \block[500] , \block[501] , \block[502] , \block[503] , \block[504] , \block[505] , \block[506] , \block[507] , \block[508] , \block[509] , \block[510] , \block[511] , ready, \digest[0] , \digest[1] , \digest[2] , \digest[3] , \digest[4] , \digest[5] , \digest[6] , \digest[7] , \digest[8] , \digest[9] , \digest[10] , \digest[11] , \digest[12] , \digest[13] , \digest[14] , \digest[15] , \digest[16] , \digest[17] , \digest[18] , \digest[19] , \digest[20] , \digest[21] , \digest[22] , \digest[23] , \digest[24] , \digest[25] , \digest[26] , \digest[27] , \digest[28] , \digest[29] , \digest[30] , \digest[31] , \digest[32] , \digest[33] , \digest[34] , \digest[35] , \digest[36] , \digest[37] , \digest[38] , \digest[39] , \digest[40] , \digest[41] , \digest[42] , \digest[43] , \digest[44] , \digest[45] , \digest[46] , \digest[47] , \digest[48] , \digest[49] , \digest[50] , \digest[51] , \digest[52] , \digest[53] , \digest[54] , \digest[55] , \digest[56] , \digest[57] , \digest[58] , \digest[59] , \digest[60] , \digest[61] , \digest[62] , \digest[63] , \digest[64] , \digest[65] , \digest[66] , \digest[67] , \digest[68] , \digest[69] , \digest[70] , \digest[71] , \digest[72] , \digest[73] , \digest[74] , \digest[75] , \digest[76] , \digest[77] , \digest[78] , \digest[79] , \digest[80] , \digest[81] , \digest[82] , \digest[83] , \digest[84] , \digest[85] , \digest[86] , \digest[87] , \digest[88] , \digest[89] , \digest[90] , \digest[91] , \digest[92] , \digest[93] , \digest[94] , \digest[95] , \digest[96] , \digest[97] , \digest[98] , \digest[99] , \digest[100] , \digest[101] , \digest[102] , \digest[103] , \digest[104] , \digest[105] , \digest[106] , \digest[107] , \digest[108] , \digest[109] , \digest[110] , \digest[111] , \digest[112] , \digest[113] , \digest[114] , \digest[115] , \digest[116] , \digest[117] , \digest[118] , \digest[119] , \digest[120] , \digest[121] , \digest[122] , \digest[123] , \digest[124] , \digest[125] , \digest[126] , \digest[127] , \digest[128] , \digest[129] , \digest[130] , \digest[131] , \digest[132] , \digest[133] , \digest[134] , \digest[135] , \digest[136] , \digest[137] , \digest[138] , \digest[139] , \digest[140] , \digest[141] , \digest[142] , \digest[143] , \digest[144] , \digest[145] , \digest[146] , \digest[147] , \digest[148] , \digest[149] , \digest[150] , \digest[151] , \digest[152] , \digest[153] , \digest[154] , \digest[155] , \digest[156] , \digest[157] , \digest[158] , \digest[159] , digest_valid);

wire _0H0_reg_31_0__0_; 
wire _0H0_reg_31_0__10_; 
wire _0H0_reg_31_0__11_; 
wire _0H0_reg_31_0__12_; 
wire _0H0_reg_31_0__13_; 
wire _0H0_reg_31_0__14_; 
wire _0H0_reg_31_0__15_; 
wire _0H0_reg_31_0__16_; 
wire _0H0_reg_31_0__17_; 
wire _0H0_reg_31_0__18_; 
wire _0H0_reg_31_0__19_; 
wire _0H0_reg_31_0__1_; 
wire _0H0_reg_31_0__20_; 
wire _0H0_reg_31_0__21_; 
wire _0H0_reg_31_0__22_; 
wire _0H0_reg_31_0__23_; 
wire _0H0_reg_31_0__24_; 
wire _0H0_reg_31_0__25_; 
wire _0H0_reg_31_0__26_; 
wire _0H0_reg_31_0__27_; 
wire _0H0_reg_31_0__28_; 
wire _0H0_reg_31_0__29_; 
wire _0H0_reg_31_0__2_; 
wire _0H0_reg_31_0__30_; 
wire _0H0_reg_31_0__31_; 
wire _0H0_reg_31_0__3_; 
wire _0H0_reg_31_0__4_; 
wire _0H0_reg_31_0__5_; 
wire _0H0_reg_31_0__6_; 
wire _0H0_reg_31_0__7_; 
wire _0H0_reg_31_0__8_; 
wire _0H0_reg_31_0__9_; 
wire _0H1_reg_31_0__0_; 
wire _0H1_reg_31_0__10_; 
wire _0H1_reg_31_0__11_; 
wire _0H1_reg_31_0__12_; 
wire _0H1_reg_31_0__13_; 
wire _0H1_reg_31_0__14_; 
wire _0H1_reg_31_0__15_; 
wire _0H1_reg_31_0__16_; 
wire _0H1_reg_31_0__17_; 
wire _0H1_reg_31_0__18_; 
wire _0H1_reg_31_0__19_; 
wire _0H1_reg_31_0__1_; 
wire _0H1_reg_31_0__20_; 
wire _0H1_reg_31_0__21_; 
wire _0H1_reg_31_0__22_; 
wire _0H1_reg_31_0__23_; 
wire _0H1_reg_31_0__24_; 
wire _0H1_reg_31_0__25_; 
wire _0H1_reg_31_0__26_; 
wire _0H1_reg_31_0__27_; 
wire _0H1_reg_31_0__28_; 
wire _0H1_reg_31_0__29_; 
wire _0H1_reg_31_0__2_; 
wire _0H1_reg_31_0__30_; 
wire _0H1_reg_31_0__31_; 
wire _0H1_reg_31_0__3_; 
wire _0H1_reg_31_0__4_; 
wire _0H1_reg_31_0__5_; 
wire _0H1_reg_31_0__6_; 
wire _0H1_reg_31_0__7_; 
wire _0H1_reg_31_0__8_; 
wire _0H1_reg_31_0__9_; 
wire _0H2_reg_31_0__0_; 
wire _0H2_reg_31_0__10_; 
wire _0H2_reg_31_0__11_; 
wire _0H2_reg_31_0__12_; 
wire _0H2_reg_31_0__13_; 
wire _0H2_reg_31_0__14_; 
wire _0H2_reg_31_0__15_; 
wire _0H2_reg_31_0__16_; 
wire _0H2_reg_31_0__17_; 
wire _0H2_reg_31_0__18_; 
wire _0H2_reg_31_0__19_; 
wire _0H2_reg_31_0__1_; 
wire _0H2_reg_31_0__20_; 
wire _0H2_reg_31_0__21_; 
wire _0H2_reg_31_0__22_; 
wire _0H2_reg_31_0__23_; 
wire _0H2_reg_31_0__24_; 
wire _0H2_reg_31_0__25_; 
wire _0H2_reg_31_0__26_; 
wire _0H2_reg_31_0__27_; 
wire _0H2_reg_31_0__28_; 
wire _0H2_reg_31_0__29_; 
wire _0H2_reg_31_0__2_; 
wire _0H2_reg_31_0__30_; 
wire _0H2_reg_31_0__31_; 
wire _0H2_reg_31_0__3_; 
wire _0H2_reg_31_0__4_; 
wire _0H2_reg_31_0__5_; 
wire _0H2_reg_31_0__6_; 
wire _0H2_reg_31_0__7_; 
wire _0H2_reg_31_0__8_; 
wire _0H2_reg_31_0__9_; 
wire _0H3_reg_31_0__0_; 
wire _0H3_reg_31_0__10_; 
wire _0H3_reg_31_0__11_; 
wire _0H3_reg_31_0__12_; 
wire _0H3_reg_31_0__13_; 
wire _0H3_reg_31_0__14_; 
wire _0H3_reg_31_0__15_; 
wire _0H3_reg_31_0__16_; 
wire _0H3_reg_31_0__17_; 
wire _0H3_reg_31_0__18_; 
wire _0H3_reg_31_0__19_; 
wire _0H3_reg_31_0__1_; 
wire _0H3_reg_31_0__20_; 
wire _0H3_reg_31_0__21_; 
wire _0H3_reg_31_0__22_; 
wire _0H3_reg_31_0__23_; 
wire _0H3_reg_31_0__24_; 
wire _0H3_reg_31_0__25_; 
wire _0H3_reg_31_0__26_; 
wire _0H3_reg_31_0__27_; 
wire _0H3_reg_31_0__28_; 
wire _0H3_reg_31_0__29_; 
wire _0H3_reg_31_0__2_; 
wire _0H3_reg_31_0__30_; 
wire _0H3_reg_31_0__31_; 
wire _0H3_reg_31_0__3_; 
wire _0H3_reg_31_0__4_; 
wire _0H3_reg_31_0__5_; 
wire _0H3_reg_31_0__6_; 
wire _0H3_reg_31_0__7_; 
wire _0H3_reg_31_0__8_; 
wire _0H3_reg_31_0__9_; 
wire _0H4_reg_31_0__0_; 
wire _0H4_reg_31_0__10_; 
wire _0H4_reg_31_0__11_; 
wire _0H4_reg_31_0__12_; 
wire _0H4_reg_31_0__13_; 
wire _0H4_reg_31_0__14_; 
wire _0H4_reg_31_0__15_; 
wire _0H4_reg_31_0__16_; 
wire _0H4_reg_31_0__17_; 
wire _0H4_reg_31_0__18_; 
wire _0H4_reg_31_0__19_; 
wire _0H4_reg_31_0__1_; 
wire _0H4_reg_31_0__20_; 
wire _0H4_reg_31_0__21_; 
wire _0H4_reg_31_0__22_; 
wire _0H4_reg_31_0__23_; 
wire _0H4_reg_31_0__24_; 
wire _0H4_reg_31_0__25_; 
wire _0H4_reg_31_0__26_; 
wire _0H4_reg_31_0__27_; 
wire _0H4_reg_31_0__28_; 
wire _0H4_reg_31_0__29_; 
wire _0H4_reg_31_0__2_; 
wire _0H4_reg_31_0__30_; 
wire _0H4_reg_31_0__31_; 
wire _0H4_reg_31_0__3_; 
wire _0H4_reg_31_0__4_; 
wire _0H4_reg_31_0__5_; 
wire _0H4_reg_31_0__6_; 
wire _0H4_reg_31_0__7_; 
wire _0H4_reg_31_0__8_; 
wire _0H4_reg_31_0__9_; 
wire _0a_reg_31_0__0_; 
wire _0a_reg_31_0__10_; 
wire _0a_reg_31_0__11_; 
wire _0a_reg_31_0__12_; 
wire _0a_reg_31_0__13_; 
wire _0a_reg_31_0__14_; 
wire _0a_reg_31_0__15_; 
wire _0a_reg_31_0__16_; 
wire _0a_reg_31_0__17_; 
wire _0a_reg_31_0__18_; 
wire _0a_reg_31_0__19_; 
wire _0a_reg_31_0__1_; 
wire _0a_reg_31_0__20_; 
wire _0a_reg_31_0__21_; 
wire _0a_reg_31_0__22_; 
wire _0a_reg_31_0__23_; 
wire _0a_reg_31_0__24_; 
wire _0a_reg_31_0__25_; 
wire _0a_reg_31_0__26_; 
wire _0a_reg_31_0__27_; 
wire _0a_reg_31_0__28_; 
wire _0a_reg_31_0__29_; 
wire _0a_reg_31_0__2_; 
wire _0a_reg_31_0__30_; 
wire _0a_reg_31_0__31_; 
wire _0a_reg_31_0__3_; 
wire _0a_reg_31_0__4_; 
wire _0a_reg_31_0__5_; 
wire _0a_reg_31_0__6_; 
wire _0a_reg_31_0__7_; 
wire _0a_reg_31_0__8_; 
wire _0a_reg_31_0__9_; 
wire _0b_reg_31_0__0_; 
wire _0b_reg_31_0__10_; 
wire _0b_reg_31_0__11_; 
wire _0b_reg_31_0__12_; 
wire _0b_reg_31_0__13_; 
wire _0b_reg_31_0__14_; 
wire _0b_reg_31_0__15_; 
wire _0b_reg_31_0__16_; 
wire _0b_reg_31_0__17_; 
wire _0b_reg_31_0__18_; 
wire _0b_reg_31_0__19_; 
wire _0b_reg_31_0__1_; 
wire _0b_reg_31_0__20_; 
wire _0b_reg_31_0__21_; 
wire _0b_reg_31_0__22_; 
wire _0b_reg_31_0__23_; 
wire _0b_reg_31_0__24_; 
wire _0b_reg_31_0__25_; 
wire _0b_reg_31_0__26_; 
wire _0b_reg_31_0__27_; 
wire _0b_reg_31_0__28_; 
wire _0b_reg_31_0__29_; 
wire _0b_reg_31_0__2_; 
wire _0b_reg_31_0__30_; 
wire _0b_reg_31_0__31_; 
wire _0b_reg_31_0__3_; 
wire _0b_reg_31_0__4_; 
wire _0b_reg_31_0__5_; 
wire _0b_reg_31_0__6_; 
wire _0b_reg_31_0__7_; 
wire _0b_reg_31_0__8_; 
wire _0b_reg_31_0__9_; 
wire _0c_reg_31_0__0_; 
wire _0c_reg_31_0__10_; 
wire _0c_reg_31_0__11_; 
wire _0c_reg_31_0__12_; 
wire _0c_reg_31_0__13_; 
wire _0c_reg_31_0__14_; 
wire _0c_reg_31_0__15_; 
wire _0c_reg_31_0__16_; 
wire _0c_reg_31_0__17_; 
wire _0c_reg_31_0__18_; 
wire _0c_reg_31_0__19_; 
wire _0c_reg_31_0__1_; 
wire _0c_reg_31_0__20_; 
wire _0c_reg_31_0__21_; 
wire _0c_reg_31_0__22_; 
wire _0c_reg_31_0__23_; 
wire _0c_reg_31_0__24_; 
wire _0c_reg_31_0__25_; 
wire _0c_reg_31_0__26_; 
wire _0c_reg_31_0__27_; 
wire _0c_reg_31_0__28_; 
wire _0c_reg_31_0__29_; 
wire _0c_reg_31_0__2_; 
wire _0c_reg_31_0__30_; 
wire _0c_reg_31_0__31_; 
wire _0c_reg_31_0__3_; 
wire _0c_reg_31_0__4_; 
wire _0c_reg_31_0__5_; 
wire _0c_reg_31_0__6_; 
wire _0c_reg_31_0__7_; 
wire _0c_reg_31_0__8_; 
wire _0c_reg_31_0__9_; 
wire _0d_reg_31_0__0_; 
wire _0d_reg_31_0__10_; 
wire _0d_reg_31_0__11_; 
wire _0d_reg_31_0__12_; 
wire _0d_reg_31_0__13_; 
wire _0d_reg_31_0__14_; 
wire _0d_reg_31_0__15_; 
wire _0d_reg_31_0__16_; 
wire _0d_reg_31_0__17_; 
wire _0d_reg_31_0__18_; 
wire _0d_reg_31_0__19_; 
wire _0d_reg_31_0__1_; 
wire _0d_reg_31_0__20_; 
wire _0d_reg_31_0__21_; 
wire _0d_reg_31_0__22_; 
wire _0d_reg_31_0__23_; 
wire _0d_reg_31_0__24_; 
wire _0d_reg_31_0__25_; 
wire _0d_reg_31_0__26_; 
wire _0d_reg_31_0__27_; 
wire _0d_reg_31_0__28_; 
wire _0d_reg_31_0__29_; 
wire _0d_reg_31_0__2_; 
wire _0d_reg_31_0__30_; 
wire _0d_reg_31_0__31_; 
wire _0d_reg_31_0__3_; 
wire _0d_reg_31_0__4_; 
wire _0d_reg_31_0__5_; 
wire _0d_reg_31_0__6_; 
wire _0d_reg_31_0__7_; 
wire _0d_reg_31_0__8_; 
wire _0d_reg_31_0__9_; 
wire _0digest_valid_reg_0_0_; 
wire _0e_reg_31_0__0_; 
wire _0e_reg_31_0__10_; 
wire _0e_reg_31_0__11_; 
wire _0e_reg_31_0__12_; 
wire _0e_reg_31_0__13_; 
wire _0e_reg_31_0__14_; 
wire _0e_reg_31_0__15_; 
wire _0e_reg_31_0__16_; 
wire _0e_reg_31_0__17_; 
wire _0e_reg_31_0__18_; 
wire _0e_reg_31_0__19_; 
wire _0e_reg_31_0__1_; 
wire _0e_reg_31_0__20_; 
wire _0e_reg_31_0__21_; 
wire _0e_reg_31_0__22_; 
wire _0e_reg_31_0__23_; 
wire _0e_reg_31_0__24_; 
wire _0e_reg_31_0__25_; 
wire _0e_reg_31_0__26_; 
wire _0e_reg_31_0__27_; 
wire _0e_reg_31_0__28_; 
wire _0e_reg_31_0__29_; 
wire _0e_reg_31_0__2_; 
wire _0e_reg_31_0__30_; 
wire _0e_reg_31_0__31_; 
wire _0e_reg_31_0__3_; 
wire _0e_reg_31_0__4_; 
wire _0e_reg_31_0__5_; 
wire _0e_reg_31_0__6_; 
wire _0e_reg_31_0__7_; 
wire _0e_reg_31_0__8_; 
wire _0e_reg_31_0__9_; 
wire _0round_ctr_reg_6_0__0_; 
wire _0round_ctr_reg_6_0__1_; 
wire _0round_ctr_reg_6_0__2_; 
wire _0round_ctr_reg_6_0__3_; 
wire _0round_ctr_reg_6_0__4_; 
wire _0round_ctr_reg_6_0__5_; 
wire _0round_ctr_reg_6_0__6_; 
wire _abc_15497_abc_9717_auto_fsm_map_cc_118_implement_pattern_cache_863; 
wire _abc_15497_abc_9717_auto_fsm_map_cc_170_map_fsm_844_0_; 
wire _abc_15497_abc_9717_auto_fsm_map_cc_170_map_fsm_844_2_; 
wire _abc_15497_new_n1000_; 
wire _abc_15497_new_n1001_; 
wire _abc_15497_new_n1002_; 
wire _abc_15497_new_n1003_; 
wire _abc_15497_new_n1004_; 
wire _abc_15497_new_n1005_; 
wire _abc_15497_new_n1006_; 
wire _abc_15497_new_n1007_; 
wire _abc_15497_new_n1009_; 
wire _abc_15497_new_n1010_; 
wire _abc_15497_new_n1011_; 
wire _abc_15497_new_n1012_; 
wire _abc_15497_new_n1013_; 
wire _abc_15497_new_n1014_; 
wire _abc_15497_new_n1016_; 
wire _abc_15497_new_n1017_; 
wire _abc_15497_new_n1018_; 
wire _abc_15497_new_n1019_; 
wire _abc_15497_new_n1020_; 
wire _abc_15497_new_n1021_; 
wire _abc_15497_new_n1022_; 
wire _abc_15497_new_n1023_; 
wire _abc_15497_new_n1024_; 
wire _abc_15497_new_n1025_; 
wire _abc_15497_new_n1026_; 
wire _abc_15497_new_n1028_; 
wire _abc_15497_new_n1029_; 
wire _abc_15497_new_n1030_; 
wire _abc_15497_new_n1031_; 
wire _abc_15497_new_n1032_; 
wire _abc_15497_new_n1033_; 
wire _abc_15497_new_n1034_; 
wire _abc_15497_new_n1035_; 
wire _abc_15497_new_n1036_; 
wire _abc_15497_new_n1037_; 
wire _abc_15497_new_n1038_; 
wire _abc_15497_new_n1039_; 
wire _abc_15497_new_n1040_; 
wire _abc_15497_new_n1042_; 
wire _abc_15497_new_n1043_; 
wire _abc_15497_new_n1044_; 
wire _abc_15497_new_n1045_; 
wire _abc_15497_new_n1046_; 
wire _abc_15497_new_n1047_; 
wire _abc_15497_new_n1048_; 
wire _abc_15497_new_n1049_; 
wire _abc_15497_new_n1050_; 
wire _abc_15497_new_n1051_; 
wire _abc_15497_new_n1052_; 
wire _abc_15497_new_n1053_; 
wire _abc_15497_new_n1054_; 
wire _abc_15497_new_n1056_; 
wire _abc_15497_new_n1057_; 
wire _abc_15497_new_n1058_; 
wire _abc_15497_new_n1059_; 
wire _abc_15497_new_n1060_; 
wire _abc_15497_new_n1061_; 
wire _abc_15497_new_n1062_; 
wire _abc_15497_new_n1063_; 
wire _abc_15497_new_n1064_; 
wire _abc_15497_new_n1065_; 
wire _abc_15497_new_n1066_; 
wire _abc_15497_new_n1067_; 
wire _abc_15497_new_n1068_; 
wire _abc_15497_new_n1069_; 
wire _abc_15497_new_n1070_; 
wire _abc_15497_new_n1071_; 
wire _abc_15497_new_n1073_; 
wire _abc_15497_new_n1074_; 
wire _abc_15497_new_n1075_; 
wire _abc_15497_new_n1076_; 
wire _abc_15497_new_n1077_; 
wire _abc_15497_new_n1078_; 
wire _abc_15497_new_n1079_; 
wire _abc_15497_new_n1080_; 
wire _abc_15497_new_n1081_; 
wire _abc_15497_new_n1082_; 
wire _abc_15497_new_n1083_; 
wire _abc_15497_new_n1084_; 
wire _abc_15497_new_n1085_; 
wire _abc_15497_new_n1086_; 
wire _abc_15497_new_n1088_; 
wire _abc_15497_new_n1089_; 
wire _abc_15497_new_n1090_; 
wire _abc_15497_new_n1091_; 
wire _abc_15497_new_n1092_; 
wire _abc_15497_new_n1093_; 
wire _abc_15497_new_n1094_; 
wire _abc_15497_new_n1095_; 
wire _abc_15497_new_n1096_; 
wire _abc_15497_new_n1097_; 
wire _abc_15497_new_n1098_; 
wire _abc_15497_new_n1099_; 
wire _abc_15497_new_n1100_; 
wire _abc_15497_new_n1101_; 
wire _abc_15497_new_n1103_; 
wire _abc_15497_new_n1104_; 
wire _abc_15497_new_n1105_; 
wire _abc_15497_new_n1106_; 
wire _abc_15497_new_n1107_; 
wire _abc_15497_new_n1108_; 
wire _abc_15497_new_n1109_; 
wire _abc_15497_new_n1110_; 
wire _abc_15497_new_n1111_; 
wire _abc_15497_new_n1112_; 
wire _abc_15497_new_n1113_; 
wire _abc_15497_new_n1114_; 
wire _abc_15497_new_n1115_; 
wire _abc_15497_new_n1116_; 
wire _abc_15497_new_n1118_; 
wire _abc_15497_new_n1119_; 
wire _abc_15497_new_n1120_; 
wire _abc_15497_new_n1121_; 
wire _abc_15497_new_n1122_; 
wire _abc_15497_new_n1123_; 
wire _abc_15497_new_n1124_; 
wire _abc_15497_new_n1125_; 
wire _abc_15497_new_n1126_; 
wire _abc_15497_new_n1127_; 
wire _abc_15497_new_n1128_; 
wire _abc_15497_new_n1129_; 
wire _abc_15497_new_n1130_; 
wire _abc_15497_new_n1132_; 
wire _abc_15497_new_n1133_; 
wire _abc_15497_new_n1134_; 
wire _abc_15497_new_n1135_; 
wire _abc_15497_new_n1136_; 
wire _abc_15497_new_n1137_; 
wire _abc_15497_new_n1138_; 
wire _abc_15497_new_n1139_; 
wire _abc_15497_new_n1140_; 
wire _abc_15497_new_n1141_; 
wire _abc_15497_new_n1142_; 
wire _abc_15497_new_n1143_; 
wire _abc_15497_new_n1144_; 
wire _abc_15497_new_n1145_; 
wire _abc_15497_new_n1146_; 
wire _abc_15497_new_n1148_; 
wire _abc_15497_new_n1149_; 
wire _abc_15497_new_n1150_; 
wire _abc_15497_new_n1151_; 
wire _abc_15497_new_n1152_; 
wire _abc_15497_new_n1153_; 
wire _abc_15497_new_n1154_; 
wire _abc_15497_new_n1155_; 
wire _abc_15497_new_n1156_; 
wire _abc_15497_new_n1157_; 
wire _abc_15497_new_n1158_; 
wire _abc_15497_new_n1159_; 
wire _abc_15497_new_n1160_; 
wire _abc_15497_new_n1162_; 
wire _abc_15497_new_n1163_; 
wire _abc_15497_new_n1164_; 
wire _abc_15497_new_n1165_; 
wire _abc_15497_new_n1166_; 
wire _abc_15497_new_n1167_; 
wire _abc_15497_new_n1168_; 
wire _abc_15497_new_n1169_; 
wire _abc_15497_new_n1170_; 
wire _abc_15497_new_n1171_; 
wire _abc_15497_new_n1172_; 
wire _abc_15497_new_n1173_; 
wire _abc_15497_new_n1175_; 
wire _abc_15497_new_n1176_; 
wire _abc_15497_new_n1177_; 
wire _abc_15497_new_n1178_; 
wire _abc_15497_new_n1179_; 
wire _abc_15497_new_n1180_; 
wire _abc_15497_new_n1181_; 
wire _abc_15497_new_n1182_; 
wire _abc_15497_new_n1183_; 
wire _abc_15497_new_n1184_; 
wire _abc_15497_new_n1185_; 
wire _abc_15497_new_n1186_; 
wire _abc_15497_new_n1187_; 
wire _abc_15497_new_n1188_; 
wire _abc_15497_new_n1189_; 
wire _abc_15497_new_n1190_; 
wire _abc_15497_new_n1191_; 
wire _abc_15497_new_n1192_; 
wire _abc_15497_new_n1193_; 
wire _abc_15497_new_n1194_; 
wire _abc_15497_new_n1195_; 
wire _abc_15497_new_n1197_; 
wire _abc_15497_new_n1198_; 
wire _abc_15497_new_n1199_; 
wire _abc_15497_new_n1200_; 
wire _abc_15497_new_n1201_; 
wire _abc_15497_new_n1202_; 
wire _abc_15497_new_n1203_; 
wire _abc_15497_new_n1204_; 
wire _abc_15497_new_n1205_; 
wire _abc_15497_new_n1206_; 
wire _abc_15497_new_n1207_; 
wire _abc_15497_new_n1208_; 
wire _abc_15497_new_n1209_; 
wire _abc_15497_new_n1211_; 
wire _abc_15497_new_n1212_; 
wire _abc_15497_new_n1213_; 
wire _abc_15497_new_n1214_; 
wire _abc_15497_new_n1215_; 
wire _abc_15497_new_n1216_; 
wire _abc_15497_new_n1217_; 
wire _abc_15497_new_n1218_; 
wire _abc_15497_new_n1219_; 
wire _abc_15497_new_n1220_; 
wire _abc_15497_new_n1221_; 
wire _abc_15497_new_n1222_; 
wire _abc_15497_new_n1223_; 
wire _abc_15497_new_n1224_; 
wire _abc_15497_new_n1225_; 
wire _abc_15497_new_n1226_; 
wire _abc_15497_new_n1228_; 
wire _abc_15497_new_n1229_; 
wire _abc_15497_new_n1230_; 
wire _abc_15497_new_n1231_; 
wire _abc_15497_new_n1232_; 
wire _abc_15497_new_n1233_; 
wire _abc_15497_new_n1234_; 
wire _abc_15497_new_n1235_; 
wire _abc_15497_new_n1236_; 
wire _abc_15497_new_n1237_; 
wire _abc_15497_new_n1238_; 
wire _abc_15497_new_n1239_; 
wire _abc_15497_new_n1240_; 
wire _abc_15497_new_n1242_; 
wire _abc_15497_new_n1243_; 
wire _abc_15497_new_n1244_; 
wire _abc_15497_new_n1245_; 
wire _abc_15497_new_n1246_; 
wire _abc_15497_new_n1247_; 
wire _abc_15497_new_n1248_; 
wire _abc_15497_new_n1249_; 
wire _abc_15497_new_n1250_; 
wire _abc_15497_new_n1251_; 
wire _abc_15497_new_n1252_; 
wire _abc_15497_new_n1253_; 
wire _abc_15497_new_n1254_; 
wire _abc_15497_new_n1255_; 
wire _abc_15497_new_n1256_; 
wire _abc_15497_new_n1257_; 
wire _abc_15497_new_n1258_; 
wire _abc_15497_new_n1259_; 
wire _abc_15497_new_n1260_; 
wire _abc_15497_new_n1261_; 
wire _abc_15497_new_n1262_; 
wire _abc_15497_new_n1263_; 
wire _abc_15497_new_n1264_; 
wire _abc_15497_new_n1265_; 
wire _abc_15497_new_n1267_; 
wire _abc_15497_new_n1268_; 
wire _abc_15497_new_n1269_; 
wire _abc_15497_new_n1270_; 
wire _abc_15497_new_n1271_; 
wire _abc_15497_new_n1272_; 
wire _abc_15497_new_n1273_; 
wire _abc_15497_new_n1274_; 
wire _abc_15497_new_n1275_; 
wire _abc_15497_new_n1276_; 
wire _abc_15497_new_n1277_; 
wire _abc_15497_new_n1278_; 
wire _abc_15497_new_n1279_; 
wire _abc_15497_new_n1281_; 
wire _abc_15497_new_n1282_; 
wire _abc_15497_new_n1283_; 
wire _abc_15497_new_n1284_; 
wire _abc_15497_new_n1285_; 
wire _abc_15497_new_n1286_; 
wire _abc_15497_new_n1287_; 
wire _abc_15497_new_n1288_; 
wire _abc_15497_new_n1289_; 
wire _abc_15497_new_n1290_; 
wire _abc_15497_new_n1291_; 
wire _abc_15497_new_n1292_; 
wire _abc_15497_new_n1293_; 
wire _abc_15497_new_n1294_; 
wire _abc_15497_new_n1295_; 
wire _abc_15497_new_n1297_; 
wire _abc_15497_new_n1298_; 
wire _abc_15497_new_n1299_; 
wire _abc_15497_new_n1300_; 
wire _abc_15497_new_n1301_; 
wire _abc_15497_new_n1302_; 
wire _abc_15497_new_n1303_; 
wire _abc_15497_new_n1304_; 
wire _abc_15497_new_n1305_; 
wire _abc_15497_new_n1306_; 
wire _abc_15497_new_n1307_; 
wire _abc_15497_new_n1308_; 
wire _abc_15497_new_n1310_; 
wire _abc_15497_new_n1311_; 
wire _abc_15497_new_n1312_; 
wire _abc_15497_new_n1313_; 
wire _abc_15497_new_n1314_; 
wire _abc_15497_new_n1315_; 
wire _abc_15497_new_n1316_; 
wire _abc_15497_new_n1317_; 
wire _abc_15497_new_n1318_; 
wire _abc_15497_new_n1319_; 
wire _abc_15497_new_n1320_; 
wire _abc_15497_new_n1321_; 
wire _abc_15497_new_n1322_; 
wire _abc_15497_new_n1323_; 
wire _abc_15497_new_n1324_; 
wire _abc_15497_new_n1325_; 
wire _abc_15497_new_n1326_; 
wire _abc_15497_new_n1327_; 
wire _abc_15497_new_n1328_; 
wire _abc_15497_new_n1329_; 
wire _abc_15497_new_n1330_; 
wire _abc_15497_new_n1331_; 
wire _abc_15497_new_n1332_; 
wire _abc_15497_new_n1333_; 
wire _abc_15497_new_n1335_; 
wire _abc_15497_new_n1336_; 
wire _abc_15497_new_n1337_; 
wire _abc_15497_new_n1338_; 
wire _abc_15497_new_n1339_; 
wire _abc_15497_new_n1340_; 
wire _abc_15497_new_n1341_; 
wire _abc_15497_new_n1342_; 
wire _abc_15497_new_n1343_; 
wire _abc_15497_new_n1344_; 
wire _abc_15497_new_n1345_; 
wire _abc_15497_new_n1346_; 
wire _abc_15497_new_n1347_; 
wire _abc_15497_new_n1348_; 
wire _abc_15497_new_n1349_; 
wire _abc_15497_new_n1351_; 
wire _abc_15497_new_n1352_; 
wire _abc_15497_new_n1353_; 
wire _abc_15497_new_n1354_; 
wire _abc_15497_new_n1355_; 
wire _abc_15497_new_n1356_; 
wire _abc_15497_new_n1357_; 
wire _abc_15497_new_n1358_; 
wire _abc_15497_new_n1359_; 
wire _abc_15497_new_n1360_; 
wire _abc_15497_new_n1361_; 
wire _abc_15497_new_n1362_; 
wire _abc_15497_new_n1363_; 
wire _abc_15497_new_n1364_; 
wire _abc_15497_new_n1366_; 
wire _abc_15497_new_n1367_; 
wire _abc_15497_new_n1368_; 
wire _abc_15497_new_n1369_; 
wire _abc_15497_new_n1370_; 
wire _abc_15497_new_n1371_; 
wire _abc_15497_new_n1372_; 
wire _abc_15497_new_n1373_; 
wire _abc_15497_new_n1374_; 
wire _abc_15497_new_n1375_; 
wire _abc_15497_new_n1376_; 
wire _abc_15497_new_n1377_; 
wire _abc_15497_new_n1378_; 
wire _abc_15497_new_n1380_; 
wire _abc_15497_new_n1381_; 
wire _abc_15497_new_n1382_; 
wire _abc_15497_new_n1383_; 
wire _abc_15497_new_n1384_; 
wire _abc_15497_new_n1385_; 
wire _abc_15497_new_n1386_; 
wire _abc_15497_new_n1387_; 
wire _abc_15497_new_n1388_; 
wire _abc_15497_new_n1389_; 
wire _abc_15497_new_n1390_; 
wire _abc_15497_new_n1391_; 
wire _abc_15497_new_n1392_; 
wire _abc_15497_new_n1393_; 
wire _abc_15497_new_n1394_; 
wire _abc_15497_new_n1395_; 
wire _abc_15497_new_n1396_; 
wire _abc_15497_new_n1397_; 
wire _abc_15497_new_n1398_; 
wire _abc_15497_new_n1399_; 
wire _abc_15497_new_n1400_; 
wire _abc_15497_new_n1401_; 
wire _abc_15497_new_n1402_; 
wire _abc_15497_new_n1404_; 
wire _abc_15497_new_n1405_; 
wire _abc_15497_new_n1406_; 
wire _abc_15497_new_n1407_; 
wire _abc_15497_new_n1408_; 
wire _abc_15497_new_n1409_; 
wire _abc_15497_new_n1410_; 
wire _abc_15497_new_n1411_; 
wire _abc_15497_new_n1412_; 
wire _abc_15497_new_n1413_; 
wire _abc_15497_new_n1414_; 
wire _abc_15497_new_n1415_; 
wire _abc_15497_new_n1416_; 
wire _abc_15497_new_n1418_; 
wire _abc_15497_new_n1419_; 
wire _abc_15497_new_n1420_; 
wire _abc_15497_new_n1421_; 
wire _abc_15497_new_n1422_; 
wire _abc_15497_new_n1423_; 
wire _abc_15497_new_n1424_; 
wire _abc_15497_new_n1425_; 
wire _abc_15497_new_n1426_; 
wire _abc_15497_new_n1427_; 
wire _abc_15497_new_n1428_; 
wire _abc_15497_new_n1429_; 
wire _abc_15497_new_n1430_; 
wire _abc_15497_new_n1431_; 
wire _abc_15497_new_n1432_; 
wire _abc_15497_new_n1434_; 
wire _abc_15497_new_n1435_; 
wire _abc_15497_new_n1436_; 
wire _abc_15497_new_n1437_; 
wire _abc_15497_new_n1438_; 
wire _abc_15497_new_n1439_; 
wire _abc_15497_new_n1440_; 
wire _abc_15497_new_n1441_; 
wire _abc_15497_new_n1442_; 
wire _abc_15497_new_n1443_; 
wire _abc_15497_new_n1444_; 
wire _abc_15497_new_n1445_; 
wire _abc_15497_new_n1446_; 
wire _abc_15497_new_n1447_; 
wire _abc_15497_new_n1448_; 
wire _abc_15497_new_n1449_; 
wire _abc_15497_new_n1450_; 
wire _abc_15497_new_n1451_; 
wire _abc_15497_new_n1452_; 
wire _abc_15497_new_n1453_; 
wire _abc_15497_new_n1454_; 
wire _abc_15497_new_n1455_; 
wire _abc_15497_new_n1456_; 
wire _abc_15497_new_n1457_; 
wire _abc_15497_new_n1458_; 
wire _abc_15497_new_n1459_; 
wire _abc_15497_new_n1460_; 
wire _abc_15497_new_n1461_; 
wire _abc_15497_new_n1462_; 
wire _abc_15497_new_n1463_; 
wire _abc_15497_new_n1465_; 
wire _abc_15497_new_n1466_; 
wire _abc_15497_new_n1467_; 
wire _abc_15497_new_n1468_; 
wire _abc_15497_new_n1469_; 
wire _abc_15497_new_n1470_; 
wire _abc_15497_new_n1471_; 
wire _abc_15497_new_n1472_; 
wire _abc_15497_new_n1473_; 
wire _abc_15497_new_n1474_; 
wire _abc_15497_new_n1475_; 
wire _abc_15497_new_n1476_; 
wire _abc_15497_new_n1477_; 
wire _abc_15497_new_n1478_; 
wire _abc_15497_new_n1479_; 
wire _abc_15497_new_n1481_; 
wire _abc_15497_new_n1482_; 
wire _abc_15497_new_n1483_; 
wire _abc_15497_new_n1484_; 
wire _abc_15497_new_n1485_; 
wire _abc_15497_new_n1486_; 
wire _abc_15497_new_n1487_; 
wire _abc_15497_new_n1488_; 
wire _abc_15497_new_n1489_; 
wire _abc_15497_new_n1490_; 
wire _abc_15497_new_n1491_; 
wire _abc_15497_new_n1492_; 
wire _abc_15497_new_n1493_; 
wire _abc_15497_new_n1494_; 
wire _abc_15497_new_n1496_; 
wire _abc_15497_new_n1497_; 
wire _abc_15497_new_n1498_; 
wire _abc_15497_new_n1499_; 
wire _abc_15497_new_n1500_; 
wire _abc_15497_new_n1501_; 
wire _abc_15497_new_n1502_; 
wire _abc_15497_new_n1503_; 
wire _abc_15497_new_n1504_; 
wire _abc_15497_new_n1505_; 
wire _abc_15497_new_n1506_; 
wire _abc_15497_new_n1507_; 
wire _abc_15497_new_n1508_; 
wire _abc_15497_new_n1509_; 
wire _abc_15497_new_n1510_; 
wire _abc_15497_new_n1511_; 
wire _abc_15497_new_n1513_; 
wire _abc_15497_new_n1514_; 
wire _abc_15497_new_n1515_; 
wire _abc_15497_new_n1516_; 
wire _abc_15497_new_n1517_; 
wire _abc_15497_new_n1518_; 
wire _abc_15497_new_n1519_; 
wire _abc_15497_new_n1520_; 
wire _abc_15497_new_n1521_; 
wire _abc_15497_new_n1522_; 
wire _abc_15497_new_n1523_; 
wire _abc_15497_new_n1524_; 
wire _abc_15497_new_n1525_; 
wire _abc_15497_new_n1526_; 
wire _abc_15497_new_n1527_; 
wire _abc_15497_new_n1529_; 
wire _abc_15497_new_n1530_; 
wire _abc_15497_new_n1531_; 
wire _abc_15497_new_n1532_; 
wire _abc_15497_new_n1533_; 
wire _abc_15497_new_n1534_; 
wire _abc_15497_new_n1536_; 
wire _abc_15497_new_n1537_; 
wire _abc_15497_new_n1538_; 
wire _abc_15497_new_n1539_; 
wire _abc_15497_new_n1540_; 
wire _abc_15497_new_n1541_; 
wire _abc_15497_new_n1542_; 
wire _abc_15497_new_n1543_; 
wire _abc_15497_new_n1544_; 
wire _abc_15497_new_n1545_; 
wire _abc_15497_new_n1546_; 
wire _abc_15497_new_n1548_; 
wire _abc_15497_new_n1549_; 
wire _abc_15497_new_n1550_; 
wire _abc_15497_new_n1551_; 
wire _abc_15497_new_n1552_; 
wire _abc_15497_new_n1553_; 
wire _abc_15497_new_n1554_; 
wire _abc_15497_new_n1555_; 
wire _abc_15497_new_n1556_; 
wire _abc_15497_new_n1557_; 
wire _abc_15497_new_n1558_; 
wire _abc_15497_new_n1559_; 
wire _abc_15497_new_n1561_; 
wire _abc_15497_new_n1562_; 
wire _abc_15497_new_n1563_; 
wire _abc_15497_new_n1564_; 
wire _abc_15497_new_n1565_; 
wire _abc_15497_new_n1566_; 
wire _abc_15497_new_n1567_; 
wire _abc_15497_new_n1568_; 
wire _abc_15497_new_n1569_; 
wire _abc_15497_new_n1570_; 
wire _abc_15497_new_n1571_; 
wire _abc_15497_new_n1572_; 
wire _abc_15497_new_n1574_; 
wire _abc_15497_new_n1575_; 
wire _abc_15497_new_n1576_; 
wire _abc_15497_new_n1577_; 
wire _abc_15497_new_n1578_; 
wire _abc_15497_new_n1579_; 
wire _abc_15497_new_n1580_; 
wire _abc_15497_new_n1581_; 
wire _abc_15497_new_n1582_; 
wire _abc_15497_new_n1583_; 
wire _abc_15497_new_n1584_; 
wire _abc_15497_new_n1585_; 
wire _abc_15497_new_n1586_; 
wire _abc_15497_new_n1588_; 
wire _abc_15497_new_n1589_; 
wire _abc_15497_new_n1590_; 
wire _abc_15497_new_n1591_; 
wire _abc_15497_new_n1592_; 
wire _abc_15497_new_n1593_; 
wire _abc_15497_new_n1594_; 
wire _abc_15497_new_n1595_; 
wire _abc_15497_new_n1596_; 
wire _abc_15497_new_n1597_; 
wire _abc_15497_new_n1598_; 
wire _abc_15497_new_n1599_; 
wire _abc_15497_new_n1601_; 
wire _abc_15497_new_n1602_; 
wire _abc_15497_new_n1603_; 
wire _abc_15497_new_n1604_; 
wire _abc_15497_new_n1605_; 
wire _abc_15497_new_n1606_; 
wire _abc_15497_new_n1607_; 
wire _abc_15497_new_n1608_; 
wire _abc_15497_new_n1609_; 
wire _abc_15497_new_n1610_; 
wire _abc_15497_new_n1611_; 
wire _abc_15497_new_n1612_; 
wire _abc_15497_new_n1614_; 
wire _abc_15497_new_n1615_; 
wire _abc_15497_new_n1616_; 
wire _abc_15497_new_n1617_; 
wire _abc_15497_new_n1618_; 
wire _abc_15497_new_n1619_; 
wire _abc_15497_new_n1620_; 
wire _abc_15497_new_n1621_; 
wire _abc_15497_new_n1622_; 
wire _abc_15497_new_n1623_; 
wire _abc_15497_new_n1624_; 
wire _abc_15497_new_n1626_; 
wire _abc_15497_new_n1627_; 
wire _abc_15497_new_n1628_; 
wire _abc_15497_new_n1629_; 
wire _abc_15497_new_n1630_; 
wire _abc_15497_new_n1631_; 
wire _abc_15497_new_n1632_; 
wire _abc_15497_new_n1633_; 
wire _abc_15497_new_n1634_; 
wire _abc_15497_new_n1635_; 
wire _abc_15497_new_n1636_; 
wire _abc_15497_new_n1638_; 
wire _abc_15497_new_n1639_; 
wire _abc_15497_new_n1640_; 
wire _abc_15497_new_n1641_; 
wire _abc_15497_new_n1642_; 
wire _abc_15497_new_n1643_; 
wire _abc_15497_new_n1644_; 
wire _abc_15497_new_n1645_; 
wire _abc_15497_new_n1646_; 
wire _abc_15497_new_n1647_; 
wire _abc_15497_new_n1648_; 
wire _abc_15497_new_n1649_; 
wire _abc_15497_new_n1650_; 
wire _abc_15497_new_n1651_; 
wire _abc_15497_new_n1652_; 
wire _abc_15497_new_n1654_; 
wire _abc_15497_new_n1655_; 
wire _abc_15497_new_n1656_; 
wire _abc_15497_new_n1657_; 
wire _abc_15497_new_n1658_; 
wire _abc_15497_new_n1659_; 
wire _abc_15497_new_n1660_; 
wire _abc_15497_new_n1661_; 
wire _abc_15497_new_n1662_; 
wire _abc_15497_new_n1663_; 
wire _abc_15497_new_n1664_; 
wire _abc_15497_new_n1665_; 
wire _abc_15497_new_n1666_; 
wire _abc_15497_new_n1667_; 
wire _abc_15497_new_n1669_; 
wire _abc_15497_new_n1670_; 
wire _abc_15497_new_n1671_; 
wire _abc_15497_new_n1672_; 
wire _abc_15497_new_n1673_; 
wire _abc_15497_new_n1674_; 
wire _abc_15497_new_n1675_; 
wire _abc_15497_new_n1676_; 
wire _abc_15497_new_n1677_; 
wire _abc_15497_new_n1678_; 
wire _abc_15497_new_n1679_; 
wire _abc_15497_new_n1680_; 
wire _abc_15497_new_n1682_; 
wire _abc_15497_new_n1683_; 
wire _abc_15497_new_n1684_; 
wire _abc_15497_new_n1685_; 
wire _abc_15497_new_n1686_; 
wire _abc_15497_new_n1687_; 
wire _abc_15497_new_n1688_; 
wire _abc_15497_new_n1689_; 
wire _abc_15497_new_n1690_; 
wire _abc_15497_new_n1691_; 
wire _abc_15497_new_n1692_; 
wire _abc_15497_new_n1693_; 
wire _abc_15497_new_n1694_; 
wire _abc_15497_new_n1695_; 
wire _abc_15497_new_n1696_; 
wire _abc_15497_new_n1697_; 
wire _abc_15497_new_n1698_; 
wire _abc_15497_new_n1699_; 
wire _abc_15497_new_n1700_; 
wire _abc_15497_new_n1701_; 
wire _abc_15497_new_n1703_; 
wire _abc_15497_new_n1704_; 
wire _abc_15497_new_n1705_; 
wire _abc_15497_new_n1706_; 
wire _abc_15497_new_n1707_; 
wire _abc_15497_new_n1708_; 
wire _abc_15497_new_n1709_; 
wire _abc_15497_new_n1710_; 
wire _abc_15497_new_n1711_; 
wire _abc_15497_new_n1712_; 
wire _abc_15497_new_n1713_; 
wire _abc_15497_new_n1714_; 
wire _abc_15497_new_n1715_; 
wire _abc_15497_new_n1716_; 
wire _abc_15497_new_n1717_; 
wire _abc_15497_new_n1719_; 
wire _abc_15497_new_n1720_; 
wire _abc_15497_new_n1721_; 
wire _abc_15497_new_n1722_; 
wire _abc_15497_new_n1723_; 
wire _abc_15497_new_n1724_; 
wire _abc_15497_new_n1725_; 
wire _abc_15497_new_n1726_; 
wire _abc_15497_new_n1727_; 
wire _abc_15497_new_n1728_; 
wire _abc_15497_new_n1729_; 
wire _abc_15497_new_n1730_; 
wire _abc_15497_new_n1731_; 
wire _abc_15497_new_n1732_; 
wire _abc_15497_new_n1734_; 
wire _abc_15497_new_n1735_; 
wire _abc_15497_new_n1736_; 
wire _abc_15497_new_n1737_; 
wire _abc_15497_new_n1738_; 
wire _abc_15497_new_n1739_; 
wire _abc_15497_new_n1740_; 
wire _abc_15497_new_n1741_; 
wire _abc_15497_new_n1742_; 
wire _abc_15497_new_n1743_; 
wire _abc_15497_new_n1744_; 
wire _abc_15497_new_n1745_; 
wire _abc_15497_new_n1747_; 
wire _abc_15497_new_n1748_; 
wire _abc_15497_new_n1749_; 
wire _abc_15497_new_n1750_; 
wire _abc_15497_new_n1751_; 
wire _abc_15497_new_n1752_; 
wire _abc_15497_new_n1753_; 
wire _abc_15497_new_n1754_; 
wire _abc_15497_new_n1755_; 
wire _abc_15497_new_n1756_; 
wire _abc_15497_new_n1757_; 
wire _abc_15497_new_n1758_; 
wire _abc_15497_new_n1759_; 
wire _abc_15497_new_n1760_; 
wire _abc_15497_new_n1761_; 
wire _abc_15497_new_n1762_; 
wire _abc_15497_new_n1763_; 
wire _abc_15497_new_n1764_; 
wire _abc_15497_new_n1765_; 
wire _abc_15497_new_n1766_; 
wire _abc_15497_new_n1767_; 
wire _abc_15497_new_n1769_; 
wire _abc_15497_new_n1770_; 
wire _abc_15497_new_n1771_; 
wire _abc_15497_new_n1772_; 
wire _abc_15497_new_n1773_; 
wire _abc_15497_new_n1774_; 
wire _abc_15497_new_n1775_; 
wire _abc_15497_new_n1776_; 
wire _abc_15497_new_n1777_; 
wire _abc_15497_new_n1778_; 
wire _abc_15497_new_n1779_; 
wire _abc_15497_new_n1780_; 
wire _abc_15497_new_n1781_; 
wire _abc_15497_new_n1783_; 
wire _abc_15497_new_n1784_; 
wire _abc_15497_new_n1785_; 
wire _abc_15497_new_n1786_; 
wire _abc_15497_new_n1787_; 
wire _abc_15497_new_n1788_; 
wire _abc_15497_new_n1789_; 
wire _abc_15497_new_n1790_; 
wire _abc_15497_new_n1791_; 
wire _abc_15497_new_n1792_; 
wire _abc_15497_new_n1793_; 
wire _abc_15497_new_n1794_; 
wire _abc_15497_new_n1795_; 
wire _abc_15497_new_n1796_; 
wire _abc_15497_new_n1797_; 
wire _abc_15497_new_n1799_; 
wire _abc_15497_new_n1800_; 
wire _abc_15497_new_n1801_; 
wire _abc_15497_new_n1802_; 
wire _abc_15497_new_n1803_; 
wire _abc_15497_new_n1804_; 
wire _abc_15497_new_n1805_; 
wire _abc_15497_new_n1806_; 
wire _abc_15497_new_n1807_; 
wire _abc_15497_new_n1808_; 
wire _abc_15497_new_n1809_; 
wire _abc_15497_new_n1810_; 
wire _abc_15497_new_n1812_; 
wire _abc_15497_new_n1813_; 
wire _abc_15497_new_n1814_; 
wire _abc_15497_new_n1815_; 
wire _abc_15497_new_n1816_; 
wire _abc_15497_new_n1817_; 
wire _abc_15497_new_n1818_; 
wire _abc_15497_new_n1819_; 
wire _abc_15497_new_n1820_; 
wire _abc_15497_new_n1821_; 
wire _abc_15497_new_n1822_; 
wire _abc_15497_new_n1823_; 
wire _abc_15497_new_n1824_; 
wire _abc_15497_new_n1825_; 
wire _abc_15497_new_n1826_; 
wire _abc_15497_new_n1827_; 
wire _abc_15497_new_n1828_; 
wire _abc_15497_new_n1829_; 
wire _abc_15497_new_n1830_; 
wire _abc_15497_new_n1832_; 
wire _abc_15497_new_n1833_; 
wire _abc_15497_new_n1834_; 
wire _abc_15497_new_n1835_; 
wire _abc_15497_new_n1836_; 
wire _abc_15497_new_n1837_; 
wire _abc_15497_new_n1838_; 
wire _abc_15497_new_n1839_; 
wire _abc_15497_new_n1840_; 
wire _abc_15497_new_n1841_; 
wire _abc_15497_new_n1842_; 
wire _abc_15497_new_n1843_; 
wire _abc_15497_new_n1844_; 
wire _abc_15497_new_n1846_; 
wire _abc_15497_new_n1847_; 
wire _abc_15497_new_n1848_; 
wire _abc_15497_new_n1849_; 
wire _abc_15497_new_n1850_; 
wire _abc_15497_new_n1851_; 
wire _abc_15497_new_n1852_; 
wire _abc_15497_new_n1853_; 
wire _abc_15497_new_n1854_; 
wire _abc_15497_new_n1855_; 
wire _abc_15497_new_n1856_; 
wire _abc_15497_new_n1857_; 
wire _abc_15497_new_n1858_; 
wire _abc_15497_new_n1859_; 
wire _abc_15497_new_n1860_; 
wire _abc_15497_new_n1862_; 
wire _abc_15497_new_n1863_; 
wire _abc_15497_new_n1864_; 
wire _abc_15497_new_n1865_; 
wire _abc_15497_new_n1866_; 
wire _abc_15497_new_n1867_; 
wire _abc_15497_new_n1868_; 
wire _abc_15497_new_n1869_; 
wire _abc_15497_new_n1870_; 
wire _abc_15497_new_n1871_; 
wire _abc_15497_new_n1872_; 
wire _abc_15497_new_n1873_; 
wire _abc_15497_new_n1875_; 
wire _abc_15497_new_n1876_; 
wire _abc_15497_new_n1877_; 
wire _abc_15497_new_n1878_; 
wire _abc_15497_new_n1879_; 
wire _abc_15497_new_n1880_; 
wire _abc_15497_new_n1881_; 
wire _abc_15497_new_n1882_; 
wire _abc_15497_new_n1883_; 
wire _abc_15497_new_n1884_; 
wire _abc_15497_new_n1885_; 
wire _abc_15497_new_n1886_; 
wire _abc_15497_new_n1887_; 
wire _abc_15497_new_n1888_; 
wire _abc_15497_new_n1889_; 
wire _abc_15497_new_n1890_; 
wire _abc_15497_new_n1891_; 
wire _abc_15497_new_n1892_; 
wire _abc_15497_new_n1893_; 
wire _abc_15497_new_n1894_; 
wire _abc_15497_new_n1895_; 
wire _abc_15497_new_n1896_; 
wire _abc_15497_new_n1897_; 
wire _abc_15497_new_n1899_; 
wire _abc_15497_new_n1900_; 
wire _abc_15497_new_n1901_; 
wire _abc_15497_new_n1902_; 
wire _abc_15497_new_n1903_; 
wire _abc_15497_new_n1904_; 
wire _abc_15497_new_n1905_; 
wire _abc_15497_new_n1906_; 
wire _abc_15497_new_n1907_; 
wire _abc_15497_new_n1908_; 
wire _abc_15497_new_n1909_; 
wire _abc_15497_new_n1910_; 
wire _abc_15497_new_n1911_; 
wire _abc_15497_new_n1912_; 
wire _abc_15497_new_n1913_; 
wire _abc_15497_new_n1915_; 
wire _abc_15497_new_n1916_; 
wire _abc_15497_new_n1917_; 
wire _abc_15497_new_n1918_; 
wire _abc_15497_new_n1919_; 
wire _abc_15497_new_n1920_; 
wire _abc_15497_new_n1921_; 
wire _abc_15497_new_n1922_; 
wire _abc_15497_new_n1923_; 
wire _abc_15497_new_n1924_; 
wire _abc_15497_new_n1925_; 
wire _abc_15497_new_n1926_; 
wire _abc_15497_new_n1927_; 
wire _abc_15497_new_n1929_; 
wire _abc_15497_new_n1930_; 
wire _abc_15497_new_n1931_; 
wire _abc_15497_new_n1932_; 
wire _abc_15497_new_n1933_; 
wire _abc_15497_new_n1934_; 
wire _abc_15497_new_n1935_; 
wire _abc_15497_new_n1936_; 
wire _abc_15497_new_n1937_; 
wire _abc_15497_new_n1938_; 
wire _abc_15497_new_n1939_; 
wire _abc_15497_new_n1940_; 
wire _abc_15497_new_n1941_; 
wire _abc_15497_new_n1942_; 
wire _abc_15497_new_n1943_; 
wire _abc_15497_new_n1945_; 
wire _abc_15497_new_n1946_; 
wire _abc_15497_new_n1947_; 
wire _abc_15497_new_n1948_; 
wire _abc_15497_new_n1949_; 
wire _abc_15497_new_n1950_; 
wire _abc_15497_new_n1951_; 
wire _abc_15497_new_n1952_; 
wire _abc_15497_new_n1953_; 
wire _abc_15497_new_n1954_; 
wire _abc_15497_new_n1955_; 
wire _abc_15497_new_n1956_; 
wire _abc_15497_new_n1957_; 
wire _abc_15497_new_n1958_; 
wire _abc_15497_new_n1959_; 
wire _abc_15497_new_n1960_; 
wire _abc_15497_new_n1961_; 
wire _abc_15497_new_n1962_; 
wire _abc_15497_new_n1964_; 
wire _abc_15497_new_n1965_; 
wire _abc_15497_new_n1966_; 
wire _abc_15497_new_n1967_; 
wire _abc_15497_new_n1968_; 
wire _abc_15497_new_n1969_; 
wire _abc_15497_new_n1970_; 
wire _abc_15497_new_n1971_; 
wire _abc_15497_new_n1972_; 
wire _abc_15497_new_n1973_; 
wire _abc_15497_new_n1974_; 
wire _abc_15497_new_n1975_; 
wire _abc_15497_new_n1977_; 
wire _abc_15497_new_n1978_; 
wire _abc_15497_new_n1979_; 
wire _abc_15497_new_n1980_; 
wire _abc_15497_new_n1981_; 
wire _abc_15497_new_n1982_; 
wire _abc_15497_new_n1983_; 
wire _abc_15497_new_n1984_; 
wire _abc_15497_new_n1985_; 
wire _abc_15497_new_n1986_; 
wire _abc_15497_new_n1987_; 
wire _abc_15497_new_n1988_; 
wire _abc_15497_new_n1989_; 
wire _abc_15497_new_n1990_; 
wire _abc_15497_new_n1991_; 
wire _abc_15497_new_n1993_; 
wire _abc_15497_new_n1994_; 
wire _abc_15497_new_n1995_; 
wire _abc_15497_new_n1996_; 
wire _abc_15497_new_n1997_; 
wire _abc_15497_new_n1998_; 
wire _abc_15497_new_n1999_; 
wire _abc_15497_new_n2000_; 
wire _abc_15497_new_n2001_; 
wire _abc_15497_new_n2002_; 
wire _abc_15497_new_n2003_; 
wire _abc_15497_new_n2004_; 
wire _abc_15497_new_n2006_; 
wire _abc_15497_new_n2008_; 
wire _abc_15497_new_n2009_; 
wire _abc_15497_new_n2010_; 
wire _abc_15497_new_n2011_; 
wire _abc_15497_new_n2012_; 
wire _abc_15497_new_n2013_; 
wire _abc_15497_new_n2014_; 
wire _abc_15497_new_n2015_; 
wire _abc_15497_new_n2016_; 
wire _abc_15497_new_n2018_; 
wire _abc_15497_new_n2019_; 
wire _abc_15497_new_n2020_; 
wire _abc_15497_new_n2021_; 
wire _abc_15497_new_n2022_; 
wire _abc_15497_new_n2024_; 
wire _abc_15497_new_n2025_; 
wire _abc_15497_new_n2026_; 
wire _abc_15497_new_n2027_; 
wire _abc_15497_new_n2028_; 
wire _abc_15497_new_n2030_; 
wire _abc_15497_new_n2031_; 
wire _abc_15497_new_n2032_; 
wire _abc_15497_new_n2033_; 
wire _abc_15497_new_n2034_; 
wire _abc_15497_new_n2036_; 
wire _abc_15497_new_n2037_; 
wire _abc_15497_new_n2038_; 
wire _abc_15497_new_n2039_; 
wire _abc_15497_new_n2041_; 
wire _abc_15497_new_n2042_; 
wire _abc_15497_new_n2043_; 
wire _abc_15497_new_n2044_; 
wire _abc_15497_new_n2046_; 
wire _abc_15497_new_n2047_; 
wire _abc_15497_new_n2048_; 
wire _abc_15497_new_n2049_; 
wire _abc_15497_new_n2051_; 
wire _abc_15497_new_n2052_; 
wire _abc_15497_new_n2053_; 
wire _abc_15497_new_n2054_; 
wire _abc_15497_new_n2056_; 
wire _abc_15497_new_n2057_; 
wire _abc_15497_new_n2058_; 
wire _abc_15497_new_n2059_; 
wire _abc_15497_new_n2061_; 
wire _abc_15497_new_n2062_; 
wire _abc_15497_new_n2063_; 
wire _abc_15497_new_n2064_; 
wire _abc_15497_new_n2065_; 
wire _abc_15497_new_n2067_; 
wire _abc_15497_new_n2068_; 
wire _abc_15497_new_n2069_; 
wire _abc_15497_new_n2070_; 
wire _abc_15497_new_n2071_; 
wire _abc_15497_new_n2073_; 
wire _abc_15497_new_n2074_; 
wire _abc_15497_new_n2075_; 
wire _abc_15497_new_n2076_; 
wire _abc_15497_new_n2077_; 
wire _abc_15497_new_n2079_; 
wire _abc_15497_new_n2080_; 
wire _abc_15497_new_n2081_; 
wire _abc_15497_new_n2082_; 
wire _abc_15497_new_n2083_; 
wire _abc_15497_new_n2085_; 
wire _abc_15497_new_n2086_; 
wire _abc_15497_new_n2087_; 
wire _abc_15497_new_n2088_; 
wire _abc_15497_new_n2090_; 
wire _abc_15497_new_n2091_; 
wire _abc_15497_new_n2092_; 
wire _abc_15497_new_n2093_; 
wire _abc_15497_new_n2095_; 
wire _abc_15497_new_n2096_; 
wire _abc_15497_new_n2097_; 
wire _abc_15497_new_n2098_; 
wire _abc_15497_new_n2100_; 
wire _abc_15497_new_n2101_; 
wire _abc_15497_new_n2102_; 
wire _abc_15497_new_n2103_; 
wire _abc_15497_new_n2104_; 
wire _abc_15497_new_n2106_; 
wire _abc_15497_new_n2107_; 
wire _abc_15497_new_n2108_; 
wire _abc_15497_new_n2109_; 
wire _abc_15497_new_n2111_; 
wire _abc_15497_new_n2112_; 
wire _abc_15497_new_n2113_; 
wire _abc_15497_new_n2114_; 
wire _abc_15497_new_n2115_; 
wire _abc_15497_new_n2117_; 
wire _abc_15497_new_n2118_; 
wire _abc_15497_new_n2119_; 
wire _abc_15497_new_n2120_; 
wire _abc_15497_new_n2121_; 
wire _abc_15497_new_n2123_; 
wire _abc_15497_new_n2124_; 
wire _abc_15497_new_n2125_; 
wire _abc_15497_new_n2126_; 
wire _abc_15497_new_n2128_; 
wire _abc_15497_new_n2129_; 
wire _abc_15497_new_n2130_; 
wire _abc_15497_new_n2131_; 
wire _abc_15497_new_n2132_; 
wire _abc_15497_new_n2134_; 
wire _abc_15497_new_n2135_; 
wire _abc_15497_new_n2136_; 
wire _abc_15497_new_n2137_; 
wire _abc_15497_new_n2139_; 
wire _abc_15497_new_n2140_; 
wire _abc_15497_new_n2141_; 
wire _abc_15497_new_n2142_; 
wire _abc_15497_new_n2144_; 
wire _abc_15497_new_n2145_; 
wire _abc_15497_new_n2146_; 
wire _abc_15497_new_n2147_; 
wire _abc_15497_new_n2149_; 
wire _abc_15497_new_n2150_; 
wire _abc_15497_new_n2151_; 
wire _abc_15497_new_n2152_; 
wire _abc_15497_new_n2154_; 
wire _abc_15497_new_n2155_; 
wire _abc_15497_new_n2156_; 
wire _abc_15497_new_n2157_; 
wire _abc_15497_new_n2158_; 
wire _abc_15497_new_n2160_; 
wire _abc_15497_new_n2161_; 
wire _abc_15497_new_n2162_; 
wire _abc_15497_new_n2163_; 
wire _abc_15497_new_n2164_; 
wire _abc_15497_new_n2166_; 
wire _abc_15497_new_n2167_; 
wire _abc_15497_new_n2168_; 
wire _abc_15497_new_n2169_; 
wire _abc_15497_new_n2170_; 
wire _abc_15497_new_n2172_; 
wire _abc_15497_new_n2173_; 
wire _abc_15497_new_n2174_; 
wire _abc_15497_new_n2175_; 
wire _abc_15497_new_n2177_; 
wire _abc_15497_new_n2178_; 
wire _abc_15497_new_n2179_; 
wire _abc_15497_new_n2180_; 
wire _abc_15497_new_n2182_; 
wire _abc_15497_new_n2183_; 
wire _abc_15497_new_n2184_; 
wire _abc_15497_new_n2185_; 
wire _abc_15497_new_n2187_; 
wire _abc_15497_new_n2188_; 
wire _abc_15497_new_n2189_; 
wire _abc_15497_new_n2190_; 
wire _abc_15497_new_n2191_; 
wire _abc_15497_new_n2192_; 
wire _abc_15497_new_n2193_; 
wire _abc_15497_new_n2195_; 
wire _abc_15497_new_n2196_; 
wire _abc_15497_new_n2197_; 
wire _abc_15497_new_n2198_; 
wire _abc_15497_new_n2199_; 
wire _abc_15497_new_n2200_; 
wire _abc_15497_new_n2201_; 
wire _abc_15497_new_n2202_; 
wire _abc_15497_new_n2203_; 
wire _abc_15497_new_n2204_; 
wire _abc_15497_new_n2205_; 
wire _abc_15497_new_n2207_; 
wire _abc_15497_new_n2208_; 
wire _abc_15497_new_n2209_; 
wire _abc_15497_new_n2210_; 
wire _abc_15497_new_n2211_; 
wire _abc_15497_new_n2212_; 
wire _abc_15497_new_n2213_; 
wire _abc_15497_new_n2214_; 
wire _abc_15497_new_n2215_; 
wire _abc_15497_new_n2216_; 
wire _abc_15497_new_n2217_; 
wire _abc_15497_new_n2218_; 
wire _abc_15497_new_n2219_; 
wire _abc_15497_new_n2221_; 
wire _abc_15497_new_n2222_; 
wire _abc_15497_new_n2223_; 
wire _abc_15497_new_n2224_; 
wire _abc_15497_new_n2225_; 
wire _abc_15497_new_n2226_; 
wire _abc_15497_new_n2227_; 
wire _abc_15497_new_n2228_; 
wire _abc_15497_new_n2229_; 
wire _abc_15497_new_n2230_; 
wire _abc_15497_new_n2231_; 
wire _abc_15497_new_n2232_; 
wire _abc_15497_new_n2233_; 
wire _abc_15497_new_n2234_; 
wire _abc_15497_new_n2236_; 
wire _abc_15497_new_n2237_; 
wire _abc_15497_new_n2238_; 
wire _abc_15497_new_n2239_; 
wire _abc_15497_new_n2240_; 
wire _abc_15497_new_n2241_; 
wire _abc_15497_new_n2242_; 
wire _abc_15497_new_n2243_; 
wire _abc_15497_new_n2244_; 
wire _abc_15497_new_n2245_; 
wire _abc_15497_new_n2246_; 
wire _abc_15497_new_n2247_; 
wire _abc_15497_new_n2248_; 
wire _abc_15497_new_n2249_; 
wire _abc_15497_new_n2250_; 
wire _abc_15497_new_n2252_; 
wire _abc_15497_new_n2253_; 
wire _abc_15497_new_n2254_; 
wire _abc_15497_new_n2255_; 
wire _abc_15497_new_n2256_; 
wire _abc_15497_new_n2257_; 
wire _abc_15497_new_n2258_; 
wire _abc_15497_new_n2259_; 
wire _abc_15497_new_n2260_; 
wire _abc_15497_new_n2261_; 
wire _abc_15497_new_n2262_; 
wire _abc_15497_new_n2263_; 
wire _abc_15497_new_n2264_; 
wire _abc_15497_new_n2266_; 
wire _abc_15497_new_n2267_; 
wire _abc_15497_new_n2268_; 
wire _abc_15497_new_n2269_; 
wire _abc_15497_new_n2270_; 
wire _abc_15497_new_n2271_; 
wire _abc_15497_new_n2272_; 
wire _abc_15497_new_n2273_; 
wire _abc_15497_new_n2274_; 
wire _abc_15497_new_n2275_; 
wire _abc_15497_new_n2276_; 
wire _abc_15497_new_n2277_; 
wire _abc_15497_new_n2278_; 
wire _abc_15497_new_n2280_; 
wire _abc_15497_new_n2281_; 
wire _abc_15497_new_n2282_; 
wire _abc_15497_new_n2283_; 
wire _abc_15497_new_n2284_; 
wire _abc_15497_new_n2285_; 
wire _abc_15497_new_n2286_; 
wire _abc_15497_new_n2287_; 
wire _abc_15497_new_n2288_; 
wire _abc_15497_new_n2289_; 
wire _abc_15497_new_n2290_; 
wire _abc_15497_new_n2291_; 
wire _abc_15497_new_n2292_; 
wire _abc_15497_new_n2293_; 
wire _abc_15497_new_n2295_; 
wire _abc_15497_new_n2296_; 
wire _abc_15497_new_n2297_; 
wire _abc_15497_new_n2298_; 
wire _abc_15497_new_n2299_; 
wire _abc_15497_new_n2300_; 
wire _abc_15497_new_n2301_; 
wire _abc_15497_new_n2302_; 
wire _abc_15497_new_n2303_; 
wire _abc_15497_new_n2304_; 
wire _abc_15497_new_n2305_; 
wire _abc_15497_new_n2306_; 
wire _abc_15497_new_n2307_; 
wire _abc_15497_new_n2309_; 
wire _abc_15497_new_n2310_; 
wire _abc_15497_new_n2311_; 
wire _abc_15497_new_n2312_; 
wire _abc_15497_new_n2313_; 
wire _abc_15497_new_n2314_; 
wire _abc_15497_new_n2315_; 
wire _abc_15497_new_n2316_; 
wire _abc_15497_new_n2317_; 
wire _abc_15497_new_n2318_; 
wire _abc_15497_new_n2319_; 
wire _abc_15497_new_n2320_; 
wire _abc_15497_new_n2321_; 
wire _abc_15497_new_n2323_; 
wire _abc_15497_new_n2324_; 
wire _abc_15497_new_n2325_; 
wire _abc_15497_new_n2326_; 
wire _abc_15497_new_n2327_; 
wire _abc_15497_new_n2328_; 
wire _abc_15497_new_n2329_; 
wire _abc_15497_new_n2330_; 
wire _abc_15497_new_n2331_; 
wire _abc_15497_new_n2332_; 
wire _abc_15497_new_n2333_; 
wire _abc_15497_new_n2334_; 
wire _abc_15497_new_n2335_; 
wire _abc_15497_new_n2336_; 
wire _abc_15497_new_n2337_; 
wire _abc_15497_new_n2338_; 
wire _abc_15497_new_n2340_; 
wire _abc_15497_new_n2341_; 
wire _abc_15497_new_n2342_; 
wire _abc_15497_new_n2343_; 
wire _abc_15497_new_n2344_; 
wire _abc_15497_new_n2345_; 
wire _abc_15497_new_n2346_; 
wire _abc_15497_new_n2347_; 
wire _abc_15497_new_n2348_; 
wire _abc_15497_new_n2349_; 
wire _abc_15497_new_n2350_; 
wire _abc_15497_new_n2351_; 
wire _abc_15497_new_n2352_; 
wire _abc_15497_new_n2354_; 
wire _abc_15497_new_n2355_; 
wire _abc_15497_new_n2356_; 
wire _abc_15497_new_n2357_; 
wire _abc_15497_new_n2358_; 
wire _abc_15497_new_n2359_; 
wire _abc_15497_new_n2360_; 
wire _abc_15497_new_n2361_; 
wire _abc_15497_new_n2362_; 
wire _abc_15497_new_n2363_; 
wire _abc_15497_new_n2364_; 
wire _abc_15497_new_n2365_; 
wire _abc_15497_new_n2366_; 
wire _abc_15497_new_n2367_; 
wire _abc_15497_new_n2368_; 
wire _abc_15497_new_n2369_; 
wire _abc_15497_new_n2370_; 
wire _abc_15497_new_n2371_; 
wire _abc_15497_new_n2373_; 
wire _abc_15497_new_n2374_; 
wire _abc_15497_new_n2375_; 
wire _abc_15497_new_n2376_; 
wire _abc_15497_new_n2377_; 
wire _abc_15497_new_n2378_; 
wire _abc_15497_new_n2379_; 
wire _abc_15497_new_n2380_; 
wire _abc_15497_new_n2381_; 
wire _abc_15497_new_n2382_; 
wire _abc_15497_new_n2383_; 
wire _abc_15497_new_n2384_; 
wire _abc_15497_new_n2385_; 
wire _abc_15497_new_n2387_; 
wire _abc_15497_new_n2388_; 
wire _abc_15497_new_n2389_; 
wire _abc_15497_new_n2390_; 
wire _abc_15497_new_n2391_; 
wire _abc_15497_new_n2392_; 
wire _abc_15497_new_n2393_; 
wire _abc_15497_new_n2394_; 
wire _abc_15497_new_n2395_; 
wire _abc_15497_new_n2396_; 
wire _abc_15497_new_n2397_; 
wire _abc_15497_new_n2398_; 
wire _abc_15497_new_n2399_; 
wire _abc_15497_new_n2400_; 
wire _abc_15497_new_n2401_; 
wire _abc_15497_new_n2403_; 
wire _abc_15497_new_n2404_; 
wire _abc_15497_new_n2405_; 
wire _abc_15497_new_n2406_; 
wire _abc_15497_new_n2407_; 
wire _abc_15497_new_n2408_; 
wire _abc_15497_new_n2409_; 
wire _abc_15497_new_n2410_; 
wire _abc_15497_new_n2411_; 
wire _abc_15497_new_n2412_; 
wire _abc_15497_new_n2413_; 
wire _abc_15497_new_n2414_; 
wire _abc_15497_new_n2415_; 
wire _abc_15497_new_n2417_; 
wire _abc_15497_new_n2418_; 
wire _abc_15497_new_n2419_; 
wire _abc_15497_new_n2420_; 
wire _abc_15497_new_n2421_; 
wire _abc_15497_new_n2422_; 
wire _abc_15497_new_n2423_; 
wire _abc_15497_new_n2424_; 
wire _abc_15497_new_n2425_; 
wire _abc_15497_new_n2426_; 
wire _abc_15497_new_n2427_; 
wire _abc_15497_new_n2428_; 
wire _abc_15497_new_n2429_; 
wire _abc_15497_new_n2430_; 
wire _abc_15497_new_n2431_; 
wire _abc_15497_new_n2432_; 
wire _abc_15497_new_n2433_; 
wire _abc_15497_new_n2434_; 
wire _abc_15497_new_n2435_; 
wire _abc_15497_new_n2436_; 
wire _abc_15497_new_n2437_; 
wire _abc_15497_new_n2438_; 
wire _abc_15497_new_n2439_; 
wire _abc_15497_new_n2440_; 
wire _abc_15497_new_n2442_; 
wire _abc_15497_new_n2443_; 
wire _abc_15497_new_n2444_; 
wire _abc_15497_new_n2445_; 
wire _abc_15497_new_n2446_; 
wire _abc_15497_new_n2447_; 
wire _abc_15497_new_n2448_; 
wire _abc_15497_new_n2449_; 
wire _abc_15497_new_n2450_; 
wire _abc_15497_new_n2451_; 
wire _abc_15497_new_n2452_; 
wire _abc_15497_new_n2453_; 
wire _abc_15497_new_n2454_; 
wire _abc_15497_new_n2455_; 
wire _abc_15497_new_n2456_; 
wire _abc_15497_new_n2458_; 
wire _abc_15497_new_n2459_; 
wire _abc_15497_new_n2460_; 
wire _abc_15497_new_n2461_; 
wire _abc_15497_new_n2462_; 
wire _abc_15497_new_n2463_; 
wire _abc_15497_new_n2464_; 
wire _abc_15497_new_n2465_; 
wire _abc_15497_new_n2466_; 
wire _abc_15497_new_n2467_; 
wire _abc_15497_new_n2468_; 
wire _abc_15497_new_n2469_; 
wire _abc_15497_new_n2470_; 
wire _abc_15497_new_n2471_; 
wire _abc_15497_new_n2473_; 
wire _abc_15497_new_n2474_; 
wire _abc_15497_new_n2475_; 
wire _abc_15497_new_n2476_; 
wire _abc_15497_new_n2477_; 
wire _abc_15497_new_n2478_; 
wire _abc_15497_new_n2479_; 
wire _abc_15497_new_n2480_; 
wire _abc_15497_new_n2481_; 
wire _abc_15497_new_n2482_; 
wire _abc_15497_new_n2483_; 
wire _abc_15497_new_n2484_; 
wire _abc_15497_new_n2485_; 
wire _abc_15497_new_n2487_; 
wire _abc_15497_new_n2488_; 
wire _abc_15497_new_n2489_; 
wire _abc_15497_new_n2490_; 
wire _abc_15497_new_n2491_; 
wire _abc_15497_new_n2492_; 
wire _abc_15497_new_n2493_; 
wire _abc_15497_new_n2494_; 
wire _abc_15497_new_n2495_; 
wire _abc_15497_new_n2496_; 
wire _abc_15497_new_n2497_; 
wire _abc_15497_new_n2498_; 
wire _abc_15497_new_n2499_; 
wire _abc_15497_new_n2500_; 
wire _abc_15497_new_n2501_; 
wire _abc_15497_new_n2502_; 
wire _abc_15497_new_n2503_; 
wire _abc_15497_new_n2504_; 
wire _abc_15497_new_n2505_; 
wire _abc_15497_new_n2506_; 
wire _abc_15497_new_n2507_; 
wire _abc_15497_new_n2509_; 
wire _abc_15497_new_n2510_; 
wire _abc_15497_new_n2511_; 
wire _abc_15497_new_n2512_; 
wire _abc_15497_new_n2513_; 
wire _abc_15497_new_n2514_; 
wire _abc_15497_new_n2515_; 
wire _abc_15497_new_n2516_; 
wire _abc_15497_new_n2517_; 
wire _abc_15497_new_n2518_; 
wire _abc_15497_new_n2519_; 
wire _abc_15497_new_n2520_; 
wire _abc_15497_new_n2521_; 
wire _abc_15497_new_n2522_; 
wire _abc_15497_new_n2524_; 
wire _abc_15497_new_n2525_; 
wire _abc_15497_new_n2526_; 
wire _abc_15497_new_n2527_; 
wire _abc_15497_new_n2528_; 
wire _abc_15497_new_n2529_; 
wire _abc_15497_new_n2530_; 
wire _abc_15497_new_n2531_; 
wire _abc_15497_new_n2532_; 
wire _abc_15497_new_n2533_; 
wire _abc_15497_new_n2534_; 
wire _abc_15497_new_n2535_; 
wire _abc_15497_new_n2536_; 
wire _abc_15497_new_n2538_; 
wire _abc_15497_new_n2539_; 
wire _abc_15497_new_n2540_; 
wire _abc_15497_new_n2541_; 
wire _abc_15497_new_n2542_; 
wire _abc_15497_new_n2543_; 
wire _abc_15497_new_n2544_; 
wire _abc_15497_new_n2545_; 
wire _abc_15497_new_n2546_; 
wire _abc_15497_new_n2547_; 
wire _abc_15497_new_n2548_; 
wire _abc_15497_new_n2549_; 
wire _abc_15497_new_n2550_; 
wire _abc_15497_new_n2552_; 
wire _abc_15497_new_n2553_; 
wire _abc_15497_new_n2554_; 
wire _abc_15497_new_n2555_; 
wire _abc_15497_new_n2556_; 
wire _abc_15497_new_n2557_; 
wire _abc_15497_new_n2558_; 
wire _abc_15497_new_n2559_; 
wire _abc_15497_new_n2560_; 
wire _abc_15497_new_n2561_; 
wire _abc_15497_new_n2562_; 
wire _abc_15497_new_n2563_; 
wire _abc_15497_new_n2564_; 
wire _abc_15497_new_n2565_; 
wire _abc_15497_new_n2566_; 
wire _abc_15497_new_n2567_; 
wire _abc_15497_new_n2568_; 
wire _abc_15497_new_n2569_; 
wire _abc_15497_new_n2570_; 
wire _abc_15497_new_n2571_; 
wire _abc_15497_new_n2572_; 
wire _abc_15497_new_n2573_; 
wire _abc_15497_new_n2574_; 
wire _abc_15497_new_n2576_; 
wire _abc_15497_new_n2577_; 
wire _abc_15497_new_n2578_; 
wire _abc_15497_new_n2579_; 
wire _abc_15497_new_n2580_; 
wire _abc_15497_new_n2581_; 
wire _abc_15497_new_n2582_; 
wire _abc_15497_new_n2583_; 
wire _abc_15497_new_n2584_; 
wire _abc_15497_new_n2585_; 
wire _abc_15497_new_n2586_; 
wire _abc_15497_new_n2587_; 
wire _abc_15497_new_n2588_; 
wire _abc_15497_new_n2590_; 
wire _abc_15497_new_n2591_; 
wire _abc_15497_new_n2592_; 
wire _abc_15497_new_n2593_; 
wire _abc_15497_new_n2594_; 
wire _abc_15497_new_n2595_; 
wire _abc_15497_new_n2596_; 
wire _abc_15497_new_n2597_; 
wire _abc_15497_new_n2598_; 
wire _abc_15497_new_n2599_; 
wire _abc_15497_new_n2600_; 
wire _abc_15497_new_n2601_; 
wire _abc_15497_new_n2602_; 
wire _abc_15497_new_n2603_; 
wire _abc_15497_new_n2604_; 
wire _abc_15497_new_n2605_; 
wire _abc_15497_new_n2607_; 
wire _abc_15497_new_n2608_; 
wire _abc_15497_new_n2609_; 
wire _abc_15497_new_n2610_; 
wire _abc_15497_new_n2611_; 
wire _abc_15497_new_n2612_; 
wire _abc_15497_new_n2613_; 
wire _abc_15497_new_n2614_; 
wire _abc_15497_new_n2615_; 
wire _abc_15497_new_n2616_; 
wire _abc_15497_new_n2617_; 
wire _abc_15497_new_n2618_; 
wire _abc_15497_new_n2619_; 
wire _abc_15497_new_n2621_; 
wire _abc_15497_new_n2622_; 
wire _abc_15497_new_n2623_; 
wire _abc_15497_new_n2624_; 
wire _abc_15497_new_n2625_; 
wire _abc_15497_new_n2626_; 
wire _abc_15497_new_n2627_; 
wire _abc_15497_new_n2628_; 
wire _abc_15497_new_n2629_; 
wire _abc_15497_new_n2630_; 
wire _abc_15497_new_n2631_; 
wire _abc_15497_new_n2632_; 
wire _abc_15497_new_n2633_; 
wire _abc_15497_new_n2634_; 
wire _abc_15497_new_n2635_; 
wire _abc_15497_new_n2637_; 
wire _abc_15497_new_n2638_; 
wire _abc_15497_new_n2639_; 
wire _abc_15497_new_n2640_; 
wire _abc_15497_new_n2641_; 
wire _abc_15497_new_n2642_; 
wire _abc_15497_new_n2643_; 
wire _abc_15497_new_n2644_; 
wire _abc_15497_new_n2645_; 
wire _abc_15497_new_n2646_; 
wire _abc_15497_new_n2647_; 
wire _abc_15497_new_n2648_; 
wire _abc_15497_new_n2649_; 
wire _abc_15497_new_n2651_; 
wire _abc_15497_new_n2652_; 
wire _abc_15497_new_n2653_; 
wire _abc_15497_new_n2654_; 
wire _abc_15497_new_n2655_; 
wire _abc_15497_new_n2656_; 
wire _abc_15497_new_n2657_; 
wire _abc_15497_new_n2658_; 
wire _abc_15497_new_n2659_; 
wire _abc_15497_new_n2660_; 
wire _abc_15497_new_n2661_; 
wire _abc_15497_new_n2662_; 
wire _abc_15497_new_n2663_; 
wire _abc_15497_new_n2664_; 
wire _abc_15497_new_n2665_; 
wire _abc_15497_new_n2666_; 
wire _abc_15497_new_n2667_; 
wire _abc_15497_new_n2668_; 
wire _abc_15497_new_n2669_; 
wire _abc_15497_new_n2670_; 
wire _abc_15497_new_n2671_; 
wire _abc_15497_new_n2672_; 
wire _abc_15497_new_n2673_; 
wire _abc_15497_new_n2674_; 
wire _abc_15497_new_n2675_; 
wire _abc_15497_new_n2676_; 
wire _abc_15497_new_n2677_; 
wire _abc_15497_new_n2678_; 
wire _abc_15497_new_n2679_; 
wire _abc_15497_new_n2680_; 
wire _abc_15497_new_n2681_; 
wire _abc_15497_new_n2682_; 
wire _abc_15497_new_n2683_; 
wire _abc_15497_new_n2684_; 
wire _abc_15497_new_n2685_; 
wire _abc_15497_new_n2686_; 
wire _abc_15497_new_n2687_; 
wire _abc_15497_new_n2688_; 
wire _abc_15497_new_n2689_; 
wire _abc_15497_new_n2690_; 
wire _abc_15497_new_n2691_; 
wire _abc_15497_new_n2692_; 
wire _abc_15497_new_n2694_; 
wire _abc_15497_new_n2695_; 
wire _abc_15497_new_n2696_; 
wire _abc_15497_new_n2697_; 
wire _abc_15497_new_n2698_; 
wire _abc_15497_new_n2699_; 
wire _abc_15497_new_n2700_; 
wire _abc_15497_new_n2701_; 
wire _abc_15497_new_n2702_; 
wire _abc_15497_new_n2703_; 
wire _abc_15497_new_n2704_; 
wire _abc_15497_new_n2705_; 
wire _abc_15497_new_n2706_; 
wire _abc_15497_new_n2707_; 
wire _abc_15497_new_n2708_; 
wire _abc_15497_new_n2710_; 
wire _abc_15497_new_n2711_; 
wire _abc_15497_new_n2712_; 
wire _abc_15497_new_n2713_; 
wire _abc_15497_new_n2714_; 
wire _abc_15497_new_n2715_; 
wire _abc_15497_new_n2716_; 
wire _abc_15497_new_n2718_; 
wire _abc_15497_new_n2719_; 
wire _abc_15497_new_n2720_; 
wire _abc_15497_new_n2721_; 
wire _abc_15497_new_n2722_; 
wire _abc_15497_new_n2723_; 
wire _abc_15497_new_n2724_; 
wire _abc_15497_new_n2725_; 
wire _abc_15497_new_n2726_; 
wire _abc_15497_new_n2727_; 
wire _abc_15497_new_n2729_; 
wire _abc_15497_new_n2730_; 
wire _abc_15497_new_n2731_; 
wire _abc_15497_new_n2732_; 
wire _abc_15497_new_n2733_; 
wire _abc_15497_new_n2734_; 
wire _abc_15497_new_n2735_; 
wire _abc_15497_new_n2736_; 
wire _abc_15497_new_n2737_; 
wire _abc_15497_new_n2738_; 
wire _abc_15497_new_n2739_; 
wire _abc_15497_new_n2740_; 
wire _abc_15497_new_n2742_; 
wire _abc_15497_new_n2743_; 
wire _abc_15497_new_n2744_; 
wire _abc_15497_new_n2745_; 
wire _abc_15497_new_n2746_; 
wire _abc_15497_new_n2747_; 
wire _abc_15497_new_n2748_; 
wire _abc_15497_new_n2749_; 
wire _abc_15497_new_n2750_; 
wire _abc_15497_new_n2751_; 
wire _abc_15497_new_n2752_; 
wire _abc_15497_new_n2753_; 
wire _abc_15497_new_n2755_; 
wire _abc_15497_new_n2756_; 
wire _abc_15497_new_n2757_; 
wire _abc_15497_new_n2758_; 
wire _abc_15497_new_n2759_; 
wire _abc_15497_new_n2760_; 
wire _abc_15497_new_n2761_; 
wire _abc_15497_new_n2762_; 
wire _abc_15497_new_n2763_; 
wire _abc_15497_new_n2764_; 
wire _abc_15497_new_n2765_; 
wire _abc_15497_new_n2766_; 
wire _abc_15497_new_n2767_; 
wire _abc_15497_new_n2768_; 
wire _abc_15497_new_n2770_; 
wire _abc_15497_new_n2771_; 
wire _abc_15497_new_n2772_; 
wire _abc_15497_new_n2773_; 
wire _abc_15497_new_n2774_; 
wire _abc_15497_new_n2775_; 
wire _abc_15497_new_n2776_; 
wire _abc_15497_new_n2777_; 
wire _abc_15497_new_n2778_; 
wire _abc_15497_new_n2779_; 
wire _abc_15497_new_n2780_; 
wire _abc_15497_new_n2781_; 
wire _abc_15497_new_n2783_; 
wire _abc_15497_new_n2784_; 
wire _abc_15497_new_n2785_; 
wire _abc_15497_new_n2786_; 
wire _abc_15497_new_n2787_; 
wire _abc_15497_new_n2788_; 
wire _abc_15497_new_n2789_; 
wire _abc_15497_new_n2790_; 
wire _abc_15497_new_n2791_; 
wire _abc_15497_new_n2792_; 
wire _abc_15497_new_n2793_; 
wire _abc_15497_new_n2794_; 
wire _abc_15497_new_n2796_; 
wire _abc_15497_new_n2797_; 
wire _abc_15497_new_n2798_; 
wire _abc_15497_new_n2799_; 
wire _abc_15497_new_n2800_; 
wire _abc_15497_new_n2801_; 
wire _abc_15497_new_n2802_; 
wire _abc_15497_new_n2803_; 
wire _abc_15497_new_n2804_; 
wire _abc_15497_new_n2805_; 
wire _abc_15497_new_n2806_; 
wire _abc_15497_new_n2807_; 
wire _abc_15497_new_n2808_; 
wire _abc_15497_new_n2809_; 
wire _abc_15497_new_n2810_; 
wire _abc_15497_new_n2812_; 
wire _abc_15497_new_n2813_; 
wire _abc_15497_new_n2814_; 
wire _abc_15497_new_n2815_; 
wire _abc_15497_new_n2816_; 
wire _abc_15497_new_n2817_; 
wire _abc_15497_new_n2818_; 
wire _abc_15497_new_n2819_; 
wire _abc_15497_new_n2820_; 
wire _abc_15497_new_n2821_; 
wire _abc_15497_new_n2822_; 
wire _abc_15497_new_n2823_; 
wire _abc_15497_new_n2824_; 
wire _abc_15497_new_n2825_; 
wire _abc_15497_new_n2827_; 
wire _abc_15497_new_n2828_; 
wire _abc_15497_new_n2829_; 
wire _abc_15497_new_n2830_; 
wire _abc_15497_new_n2831_; 
wire _abc_15497_new_n2832_; 
wire _abc_15497_new_n2833_; 
wire _abc_15497_new_n2834_; 
wire _abc_15497_new_n2835_; 
wire _abc_15497_new_n2836_; 
wire _abc_15497_new_n2837_; 
wire _abc_15497_new_n2838_; 
wire _abc_15497_new_n2839_; 
wire _abc_15497_new_n2841_; 
wire _abc_15497_new_n2842_; 
wire _abc_15497_new_n2843_; 
wire _abc_15497_new_n2844_; 
wire _abc_15497_new_n2845_; 
wire _abc_15497_new_n2846_; 
wire _abc_15497_new_n2847_; 
wire _abc_15497_new_n2848_; 
wire _abc_15497_new_n2849_; 
wire _abc_15497_new_n2850_; 
wire _abc_15497_new_n2851_; 
wire _abc_15497_new_n2852_; 
wire _abc_15497_new_n2853_; 
wire _abc_15497_new_n2854_; 
wire _abc_15497_new_n2855_; 
wire _abc_15497_new_n2856_; 
wire _abc_15497_new_n2858_; 
wire _abc_15497_new_n2859_; 
wire _abc_15497_new_n2860_; 
wire _abc_15497_new_n2861_; 
wire _abc_15497_new_n2862_; 
wire _abc_15497_new_n2863_; 
wire _abc_15497_new_n2864_; 
wire _abc_15497_new_n2865_; 
wire _abc_15497_new_n2866_; 
wire _abc_15497_new_n2867_; 
wire _abc_15497_new_n2868_; 
wire _abc_15497_new_n2869_; 
wire _abc_15497_new_n2871_; 
wire _abc_15497_new_n2872_; 
wire _abc_15497_new_n2873_; 
wire _abc_15497_new_n2874_; 
wire _abc_15497_new_n2875_; 
wire _abc_15497_new_n2876_; 
wire _abc_15497_new_n2877_; 
wire _abc_15497_new_n2878_; 
wire _abc_15497_new_n2879_; 
wire _abc_15497_new_n2880_; 
wire _abc_15497_new_n2881_; 
wire _abc_15497_new_n2882_; 
wire _abc_15497_new_n2883_; 
wire _abc_15497_new_n2884_; 
wire _abc_15497_new_n2885_; 
wire _abc_15497_new_n2886_; 
wire _abc_15497_new_n2887_; 
wire _abc_15497_new_n2888_; 
wire _abc_15497_new_n2889_; 
wire _abc_15497_new_n2890_; 
wire _abc_15497_new_n2892_; 
wire _abc_15497_new_n2893_; 
wire _abc_15497_new_n2894_; 
wire _abc_15497_new_n2895_; 
wire _abc_15497_new_n2896_; 
wire _abc_15497_new_n2897_; 
wire _abc_15497_new_n2898_; 
wire _abc_15497_new_n2899_; 
wire _abc_15497_new_n2900_; 
wire _abc_15497_new_n2901_; 
wire _abc_15497_new_n2902_; 
wire _abc_15497_new_n2903_; 
wire _abc_15497_new_n2904_; 
wire _abc_15497_new_n2906_; 
wire _abc_15497_new_n2907_; 
wire _abc_15497_new_n2908_; 
wire _abc_15497_new_n2909_; 
wire _abc_15497_new_n2910_; 
wire _abc_15497_new_n2911_; 
wire _abc_15497_new_n2912_; 
wire _abc_15497_new_n2913_; 
wire _abc_15497_new_n2914_; 
wire _abc_15497_new_n2915_; 
wire _abc_15497_new_n2916_; 
wire _abc_15497_new_n2917_; 
wire _abc_15497_new_n2918_; 
wire _abc_15497_new_n2919_; 
wire _abc_15497_new_n2920_; 
wire _abc_15497_new_n2922_; 
wire _abc_15497_new_n2923_; 
wire _abc_15497_new_n2924_; 
wire _abc_15497_new_n2925_; 
wire _abc_15497_new_n2926_; 
wire _abc_15497_new_n2927_; 
wire _abc_15497_new_n2928_; 
wire _abc_15497_new_n2929_; 
wire _abc_15497_new_n2930_; 
wire _abc_15497_new_n2931_; 
wire _abc_15497_new_n2932_; 
wire _abc_15497_new_n2933_; 
wire _abc_15497_new_n2935_; 
wire _abc_15497_new_n2936_; 
wire _abc_15497_new_n2937_; 
wire _abc_15497_new_n2938_; 
wire _abc_15497_new_n2939_; 
wire _abc_15497_new_n2940_; 
wire _abc_15497_new_n2941_; 
wire _abc_15497_new_n2942_; 
wire _abc_15497_new_n2943_; 
wire _abc_15497_new_n2944_; 
wire _abc_15497_new_n2945_; 
wire _abc_15497_new_n2946_; 
wire _abc_15497_new_n2947_; 
wire _abc_15497_new_n2948_; 
wire _abc_15497_new_n2949_; 
wire _abc_15497_new_n2950_; 
wire _abc_15497_new_n2951_; 
wire _abc_15497_new_n2952_; 
wire _abc_15497_new_n2953_; 
wire _abc_15497_new_n2954_; 
wire _abc_15497_new_n2955_; 
wire _abc_15497_new_n2956_; 
wire _abc_15497_new_n2957_; 
wire _abc_15497_new_n2958_; 
wire _abc_15497_new_n2960_; 
wire _abc_15497_new_n2961_; 
wire _abc_15497_new_n2962_; 
wire _abc_15497_new_n2963_; 
wire _abc_15497_new_n2964_; 
wire _abc_15497_new_n2965_; 
wire _abc_15497_new_n2966_; 
wire _abc_15497_new_n2967_; 
wire _abc_15497_new_n2968_; 
wire _abc_15497_new_n2969_; 
wire _abc_15497_new_n2970_; 
wire _abc_15497_new_n2971_; 
wire _abc_15497_new_n2972_; 
wire _abc_15497_new_n2973_; 
wire _abc_15497_new_n2974_; 
wire _abc_15497_new_n2976_; 
wire _abc_15497_new_n2977_; 
wire _abc_15497_new_n2978_; 
wire _abc_15497_new_n2979_; 
wire _abc_15497_new_n2980_; 
wire _abc_15497_new_n2981_; 
wire _abc_15497_new_n2982_; 
wire _abc_15497_new_n2983_; 
wire _abc_15497_new_n2984_; 
wire _abc_15497_new_n2985_; 
wire _abc_15497_new_n2986_; 
wire _abc_15497_new_n2987_; 
wire _abc_15497_new_n2988_; 
wire _abc_15497_new_n2989_; 
wire _abc_15497_new_n2991_; 
wire _abc_15497_new_n2992_; 
wire _abc_15497_new_n2993_; 
wire _abc_15497_new_n2994_; 
wire _abc_15497_new_n2995_; 
wire _abc_15497_new_n2996_; 
wire _abc_15497_new_n2997_; 
wire _abc_15497_new_n2998_; 
wire _abc_15497_new_n2999_; 
wire _abc_15497_new_n3000_; 
wire _abc_15497_new_n3001_; 
wire _abc_15497_new_n3002_; 
wire _abc_15497_new_n3004_; 
wire _abc_15497_new_n3005_; 
wire _abc_15497_new_n3006_; 
wire _abc_15497_new_n3007_; 
wire _abc_15497_new_n3008_; 
wire _abc_15497_new_n3009_; 
wire _abc_15497_new_n3010_; 
wire _abc_15497_new_n3011_; 
wire _abc_15497_new_n3012_; 
wire _abc_15497_new_n3013_; 
wire _abc_15497_new_n3014_; 
wire _abc_15497_new_n3015_; 
wire _abc_15497_new_n3016_; 
wire _abc_15497_new_n3017_; 
wire _abc_15497_new_n3018_; 
wire _abc_15497_new_n3019_; 
wire _abc_15497_new_n3020_; 
wire _abc_15497_new_n3021_; 
wire _abc_15497_new_n3022_; 
wire _abc_15497_new_n3024_; 
wire _abc_15497_new_n3025_; 
wire _abc_15497_new_n3026_; 
wire _abc_15497_new_n3027_; 
wire _abc_15497_new_n3028_; 
wire _abc_15497_new_n3029_; 
wire _abc_15497_new_n3030_; 
wire _abc_15497_new_n3031_; 
wire _abc_15497_new_n3032_; 
wire _abc_15497_new_n3033_; 
wire _abc_15497_new_n3034_; 
wire _abc_15497_new_n3035_; 
wire _abc_15497_new_n3036_; 
wire _abc_15497_new_n3037_; 
wire _abc_15497_new_n3039_; 
wire _abc_15497_new_n3040_; 
wire _abc_15497_new_n3041_; 
wire _abc_15497_new_n3042_; 
wire _abc_15497_new_n3043_; 
wire _abc_15497_new_n3044_; 
wire _abc_15497_new_n3045_; 
wire _abc_15497_new_n3046_; 
wire _abc_15497_new_n3047_; 
wire _abc_15497_new_n3048_; 
wire _abc_15497_new_n3049_; 
wire _abc_15497_new_n3050_; 
wire _abc_15497_new_n3051_; 
wire _abc_15497_new_n3053_; 
wire _abc_15497_new_n3054_; 
wire _abc_15497_new_n3055_; 
wire _abc_15497_new_n3056_; 
wire _abc_15497_new_n3057_; 
wire _abc_15497_new_n3058_; 
wire _abc_15497_new_n3059_; 
wire _abc_15497_new_n3060_; 
wire _abc_15497_new_n3061_; 
wire _abc_15497_new_n3062_; 
wire _abc_15497_new_n3063_; 
wire _abc_15497_new_n3064_; 
wire _abc_15497_new_n3066_; 
wire _abc_15497_new_n3067_; 
wire _abc_15497_new_n3068_; 
wire _abc_15497_new_n3069_; 
wire _abc_15497_new_n3070_; 
wire _abc_15497_new_n3071_; 
wire _abc_15497_new_n3072_; 
wire _abc_15497_new_n3073_; 
wire _abc_15497_new_n3074_; 
wire _abc_15497_new_n3075_; 
wire _abc_15497_new_n3076_; 
wire _abc_15497_new_n3077_; 
wire _abc_15497_new_n3078_; 
wire _abc_15497_new_n3079_; 
wire _abc_15497_new_n3080_; 
wire _abc_15497_new_n3081_; 
wire _abc_15497_new_n3082_; 
wire _abc_15497_new_n3083_; 
wire _abc_15497_new_n3084_; 
wire _abc_15497_new_n3085_; 
wire _abc_15497_new_n3087_; 
wire _abc_15497_new_n3088_; 
wire _abc_15497_new_n3089_; 
wire _abc_15497_new_n3090_; 
wire _abc_15497_new_n3091_; 
wire _abc_15497_new_n3092_; 
wire _abc_15497_new_n3093_; 
wire _abc_15497_new_n3094_; 
wire _abc_15497_new_n3095_; 
wire _abc_15497_new_n3096_; 
wire _abc_15497_new_n3097_; 
wire _abc_15497_new_n3098_; 
wire _abc_15497_new_n3099_; 
wire _abc_15497_new_n3101_; 
wire _abc_15497_new_n3102_; 
wire _abc_15497_new_n3103_; 
wire _abc_15497_new_n3104_; 
wire _abc_15497_new_n3105_; 
wire _abc_15497_new_n3106_; 
wire _abc_15497_new_n3107_; 
wire _abc_15497_new_n3108_; 
wire _abc_15497_new_n3109_; 
wire _abc_15497_new_n3110_; 
wire _abc_15497_new_n3111_; 
wire _abc_15497_new_n3112_; 
wire _abc_15497_new_n3113_; 
wire _abc_15497_new_n3114_; 
wire _abc_15497_new_n3115_; 
wire _abc_15497_new_n3116_; 
wire _abc_15497_new_n3118_; 
wire _abc_15497_new_n3119_; 
wire _abc_15497_new_n3120_; 
wire _abc_15497_new_n3121_; 
wire _abc_15497_new_n3122_; 
wire _abc_15497_new_n3123_; 
wire _abc_15497_new_n3124_; 
wire _abc_15497_new_n3125_; 
wire _abc_15497_new_n3126_; 
wire _abc_15497_new_n3127_; 
wire _abc_15497_new_n3128_; 
wire _abc_15497_new_n3129_; 
wire _abc_15497_new_n3131_; 
wire _abc_15497_new_n3132_; 
wire _abc_15497_new_n3133_; 
wire _abc_15497_new_n3134_; 
wire _abc_15497_new_n3135_; 
wire _abc_15497_new_n3136_; 
wire _abc_15497_new_n3137_; 
wire _abc_15497_new_n3138_; 
wire _abc_15497_new_n3139_; 
wire _abc_15497_new_n3140_; 
wire _abc_15497_new_n3141_; 
wire _abc_15497_new_n3142_; 
wire _abc_15497_new_n3143_; 
wire _abc_15497_new_n3144_; 
wire _abc_15497_new_n3145_; 
wire _abc_15497_new_n3146_; 
wire _abc_15497_new_n3147_; 
wire _abc_15497_new_n3148_; 
wire _abc_15497_new_n3149_; 
wire _abc_15497_new_n3150_; 
wire _abc_15497_new_n3151_; 
wire _abc_15497_new_n3153_; 
wire _abc_15497_new_n3154_; 
wire _abc_15497_new_n3155_; 
wire _abc_15497_new_n3156_; 
wire _abc_15497_new_n3157_; 
wire _abc_15497_new_n3158_; 
wire _abc_15497_new_n3159_; 
wire _abc_15497_new_n3160_; 
wire _abc_15497_new_n3161_; 
wire _abc_15497_new_n3162_; 
wire _abc_15497_new_n3163_; 
wire _abc_15497_new_n3164_; 
wire _abc_15497_new_n3165_; 
wire _abc_15497_new_n3167_; 
wire _abc_15497_new_n3168_; 
wire _abc_15497_new_n3169_; 
wire _abc_15497_new_n3170_; 
wire _abc_15497_new_n3171_; 
wire _abc_15497_new_n3172_; 
wire _abc_15497_new_n3173_; 
wire _abc_15497_new_n3174_; 
wire _abc_15497_new_n3175_; 
wire _abc_15497_new_n3176_; 
wire _abc_15497_new_n3177_; 
wire _abc_15497_new_n3178_; 
wire _abc_15497_new_n3179_; 
wire _abc_15497_new_n3180_; 
wire _abc_15497_new_n3181_; 
wire _abc_15497_new_n3182_; 
wire _abc_15497_new_n3184_; 
wire _abc_15497_new_n3185_; 
wire _abc_15497_new_n3186_; 
wire _abc_15497_new_n3187_; 
wire _abc_15497_new_n3188_; 
wire _abc_15497_new_n3189_; 
wire _abc_15497_new_n3190_; 
wire _abc_15497_new_n3191_; 
wire _abc_15497_new_n3192_; 
wire _abc_15497_new_n3193_; 
wire _abc_15497_new_n3194_; 
wire _abc_15497_new_n3195_; 
wire _abc_15497_new_n3197_; 
wire _abc_15497_new_n3198_; 
wire _abc_15497_new_n3199_; 
wire _abc_15497_new_n3200_; 
wire _abc_15497_new_n3202_; 
wire _abc_15497_new_n3203_; 
wire _abc_15497_new_n3204_; 
wire _abc_15497_new_n3205_; 
wire _abc_15497_new_n3206_; 
wire _abc_15497_new_n3208_; 
wire _abc_15497_new_n3209_; 
wire _abc_15497_new_n3210_; 
wire _abc_15497_new_n3211_; 
wire _abc_15497_new_n3212_; 
wire _abc_15497_new_n3214_; 
wire _abc_15497_new_n3215_; 
wire _abc_15497_new_n3216_; 
wire _abc_15497_new_n3217_; 
wire _abc_15497_new_n3219_; 
wire _abc_15497_new_n3220_; 
wire _abc_15497_new_n3221_; 
wire _abc_15497_new_n3222_; 
wire _abc_15497_new_n3223_; 
wire _abc_15497_new_n3225_; 
wire _abc_15497_new_n3226_; 
wire _abc_15497_new_n3227_; 
wire _abc_15497_new_n3228_; 
wire _abc_15497_new_n3229_; 
wire _abc_15497_new_n3231_; 
wire _abc_15497_new_n3232_; 
wire _abc_15497_new_n3233_; 
wire _abc_15497_new_n3234_; 
wire _abc_15497_new_n3235_; 
wire _abc_15497_new_n3237_; 
wire _abc_15497_new_n3238_; 
wire _abc_15497_new_n3239_; 
wire _abc_15497_new_n3240_; 
wire _abc_15497_new_n3242_; 
wire _abc_15497_new_n3243_; 
wire _abc_15497_new_n3244_; 
wire _abc_15497_new_n3245_; 
wire _abc_15497_new_n3247_; 
wire _abc_15497_new_n3248_; 
wire _abc_15497_new_n3249_; 
wire _abc_15497_new_n3250_; 
wire _abc_15497_new_n3252_; 
wire _abc_15497_new_n3253_; 
wire _abc_15497_new_n3254_; 
wire _abc_15497_new_n3255_; 
wire _abc_15497_new_n3256_; 
wire _abc_15497_new_n3258_; 
wire _abc_15497_new_n3259_; 
wire _abc_15497_new_n3260_; 
wire _abc_15497_new_n3261_; 
wire _abc_15497_new_n3263_; 
wire _abc_15497_new_n3264_; 
wire _abc_15497_new_n3265_; 
wire _abc_15497_new_n3266_; 
wire _abc_15497_new_n3267_; 
wire _abc_15497_new_n3269_; 
wire _abc_15497_new_n3270_; 
wire _abc_15497_new_n3271_; 
wire _abc_15497_new_n3272_; 
wire _abc_15497_new_n3274_; 
wire _abc_15497_new_n3275_; 
wire _abc_15497_new_n3276_; 
wire _abc_15497_new_n3277_; 
wire _abc_15497_new_n3278_; 
wire _abc_15497_new_n3280_; 
wire _abc_15497_new_n3281_; 
wire _abc_15497_new_n3282_; 
wire _abc_15497_new_n3283_; 
wire _abc_15497_new_n3285_; 
wire _abc_15497_new_n3286_; 
wire _abc_15497_new_n3287_; 
wire _abc_15497_new_n3288_; 
wire _abc_15497_new_n3290_; 
wire _abc_15497_new_n3291_; 
wire _abc_15497_new_n3292_; 
wire _abc_15497_new_n3293_; 
wire _abc_15497_new_n3294_; 
wire _abc_15497_new_n3296_; 
wire _abc_15497_new_n3297_; 
wire _abc_15497_new_n3298_; 
wire _abc_15497_new_n3299_; 
wire _abc_15497_new_n3301_; 
wire _abc_15497_new_n3302_; 
wire _abc_15497_new_n3303_; 
wire _abc_15497_new_n3304_; 
wire _abc_15497_new_n3306_; 
wire _abc_15497_new_n3307_; 
wire _abc_15497_new_n3308_; 
wire _abc_15497_new_n3309_; 
wire _abc_15497_new_n3310_; 
wire _abc_15497_new_n3312_; 
wire _abc_15497_new_n3313_; 
wire _abc_15497_new_n3314_; 
wire _abc_15497_new_n3315_; 
wire _abc_15497_new_n3316_; 
wire _abc_15497_new_n3318_; 
wire _abc_15497_new_n3319_; 
wire _abc_15497_new_n3320_; 
wire _abc_15497_new_n3321_; 
wire _abc_15497_new_n3323_; 
wire _abc_15497_new_n3324_; 
wire _abc_15497_new_n3325_; 
wire _abc_15497_new_n3326_; 
wire _abc_15497_new_n3328_; 
wire _abc_15497_new_n3329_; 
wire _abc_15497_new_n3330_; 
wire _abc_15497_new_n3331_; 
wire _abc_15497_new_n3333_; 
wire _abc_15497_new_n3334_; 
wire _abc_15497_new_n3335_; 
wire _abc_15497_new_n3336_; 
wire _abc_15497_new_n3338_; 
wire _abc_15497_new_n3339_; 
wire _abc_15497_new_n3340_; 
wire _abc_15497_new_n3341_; 
wire _abc_15497_new_n3343_; 
wire _abc_15497_new_n3344_; 
wire _abc_15497_new_n3345_; 
wire _abc_15497_new_n3346_; 
wire _abc_15497_new_n3348_; 
wire _abc_15497_new_n3349_; 
wire _abc_15497_new_n3350_; 
wire _abc_15497_new_n3351_; 
wire _abc_15497_new_n3352_; 
wire _abc_15497_new_n3354_; 
wire _abc_15497_new_n3355_; 
wire _abc_15497_new_n3356_; 
wire _abc_15497_new_n3357_; 
wire _abc_15497_new_n3359_; 
wire _abc_15497_new_n3360_; 
wire _abc_15497_new_n3361_; 
wire _abc_15497_new_n3362_; 
wire _abc_15497_new_n3364_; 
wire _abc_15497_new_n3365_; 
wire _abc_15497_new_n3366_; 
wire _abc_15497_new_n3367_; 
wire _abc_15497_new_n3369_; 
wire _abc_15497_new_n3370_; 
wire _abc_15497_new_n3371_; 
wire _abc_15497_new_n3372_; 
wire _abc_15497_new_n3373_; 
wire _abc_15497_new_n3375_; 
wire _abc_15497_new_n3376_; 
wire _abc_15497_new_n3377_; 
wire _abc_15497_new_n3378_; 
wire _abc_15497_new_n3380_; 
wire _abc_15497_new_n3381_; 
wire _abc_15497_new_n3382_; 
wire _abc_15497_new_n3383_; 
wire _abc_15497_new_n3385_; 
wire _abc_15497_new_n3386_; 
wire _abc_15497_new_n3387_; 
wire _abc_15497_new_n3388_; 
wire _abc_15497_new_n3389_; 
wire _abc_15497_new_n3391_; 
wire _abc_15497_new_n3392_; 
wire _abc_15497_new_n3393_; 
wire _abc_15497_new_n3394_; 
wire _abc_15497_new_n3396_; 
wire _abc_15497_new_n3397_; 
wire _abc_15497_new_n3398_; 
wire _abc_15497_new_n3399_; 
wire _abc_15497_new_n3401_; 
wire _abc_15497_new_n3402_; 
wire _abc_15497_new_n3403_; 
wire _abc_15497_new_n3404_; 
wire _abc_15497_new_n3406_; 
wire _abc_15497_new_n3407_; 
wire _abc_15497_new_n3408_; 
wire _abc_15497_new_n3409_; 
wire _abc_15497_new_n3410_; 
wire _abc_15497_new_n3412_; 
wire _abc_15497_new_n3413_; 
wire _abc_15497_new_n3414_; 
wire _abc_15497_new_n3415_; 
wire _abc_15497_new_n3416_; 
wire _abc_15497_new_n3418_; 
wire _abc_15497_new_n3419_; 
wire _abc_15497_new_n3420_; 
wire _abc_15497_new_n3421_; 
wire _abc_15497_new_n3422_; 
wire _abc_15497_new_n3424_; 
wire _abc_15497_new_n3425_; 
wire _abc_15497_new_n3426_; 
wire _abc_15497_new_n3427_; 
wire _abc_15497_new_n3429_; 
wire _abc_15497_new_n3430_; 
wire _abc_15497_new_n3431_; 
wire _abc_15497_new_n3432_; 
wire _abc_15497_new_n3433_; 
wire _abc_15497_new_n3435_; 
wire _abc_15497_new_n3436_; 
wire _abc_15497_new_n3437_; 
wire _abc_15497_new_n3438_; 
wire _abc_15497_new_n3440_; 
wire _abc_15497_new_n3441_; 
wire _abc_15497_new_n3442_; 
wire _abc_15497_new_n3443_; 
wire _abc_15497_new_n3444_; 
wire _abc_15497_new_n3446_; 
wire _abc_15497_new_n3447_; 
wire _abc_15497_new_n3448_; 
wire _abc_15497_new_n3449_; 
wire _abc_15497_new_n3451_; 
wire _abc_15497_new_n3452_; 
wire _abc_15497_new_n3453_; 
wire _abc_15497_new_n3454_; 
wire _abc_15497_new_n3455_; 
wire _abc_15497_new_n3457_; 
wire _abc_15497_new_n3458_; 
wire _abc_15497_new_n3459_; 
wire _abc_15497_new_n3460_; 
wire _abc_15497_new_n3461_; 
wire _abc_15497_new_n3463_; 
wire _abc_15497_new_n3464_; 
wire _abc_15497_new_n3465_; 
wire _abc_15497_new_n3466_; 
wire _abc_15497_new_n3468_; 
wire _abc_15497_new_n3469_; 
wire _abc_15497_new_n3470_; 
wire _abc_15497_new_n3471_; 
wire _abc_15497_new_n3472_; 
wire _abc_15497_new_n3474_; 
wire _abc_15497_new_n3475_; 
wire _abc_15497_new_n3476_; 
wire _abc_15497_new_n3477_; 
wire _abc_15497_new_n3478_; 
wire _abc_15497_new_n3480_; 
wire _abc_15497_new_n3481_; 
wire _abc_15497_new_n3482_; 
wire _abc_15497_new_n3483_; 
wire _abc_15497_new_n3485_; 
wire _abc_15497_new_n3486_; 
wire _abc_15497_new_n3487_; 
wire _abc_15497_new_n3488_; 
wire _abc_15497_new_n3490_; 
wire _abc_15497_new_n3491_; 
wire _abc_15497_new_n3492_; 
wire _abc_15497_new_n3493_; 
wire _abc_15497_new_n3494_; 
wire _abc_15497_new_n3496_; 
wire _abc_15497_new_n3497_; 
wire _abc_15497_new_n3498_; 
wire _abc_15497_new_n3499_; 
wire _abc_15497_new_n3500_; 
wire _abc_15497_new_n3502_; 
wire _abc_15497_new_n3503_; 
wire _abc_15497_new_n3504_; 
wire _abc_15497_new_n3505_; 
wire _abc_15497_new_n3506_; 
wire _abc_15497_new_n3508_; 
wire _abc_15497_new_n3509_; 
wire _abc_15497_new_n3510_; 
wire _abc_15497_new_n3511_; 
wire _abc_15497_new_n3512_; 
wire _abc_15497_new_n3514_; 
wire _abc_15497_new_n3515_; 
wire _abc_15497_new_n3516_; 
wire _abc_15497_new_n3517_; 
wire _abc_15497_new_n3518_; 
wire _abc_15497_new_n3520_; 
wire _abc_15497_new_n3521_; 
wire _abc_15497_new_n3522_; 
wire _abc_15497_new_n3523_; 
wire _abc_15497_new_n3524_; 
wire _abc_15497_new_n3526_; 
wire _abc_15497_new_n3527_; 
wire _abc_15497_new_n3528_; 
wire _abc_15497_new_n3529_; 
wire _abc_15497_new_n3531_; 
wire _abc_15497_new_n3532_; 
wire _abc_15497_new_n3533_; 
wire _abc_15497_new_n3534_; 
wire _abc_15497_new_n3535_; 
wire _abc_15497_new_n3537_; 
wire _abc_15497_new_n3538_; 
wire _abc_15497_new_n3539_; 
wire _abc_15497_new_n3540_; 
wire _abc_15497_new_n3541_; 
wire _abc_15497_new_n3543_; 
wire _abc_15497_new_n3544_; 
wire _abc_15497_new_n3545_; 
wire _abc_15497_new_n3546_; 
wire _abc_15497_new_n3547_; 
wire _abc_15497_new_n3549_; 
wire _abc_15497_new_n3550_; 
wire _abc_15497_new_n3551_; 
wire _abc_15497_new_n3552_; 
wire _abc_15497_new_n3553_; 
wire _abc_15497_new_n3555_; 
wire _abc_15497_new_n3556_; 
wire _abc_15497_new_n3557_; 
wire _abc_15497_new_n3558_; 
wire _abc_15497_new_n3559_; 
wire _abc_15497_new_n3561_; 
wire _abc_15497_new_n3562_; 
wire _abc_15497_new_n3563_; 
wire _abc_15497_new_n3564_; 
wire _abc_15497_new_n3565_; 
wire _abc_15497_new_n3567_; 
wire _abc_15497_new_n3568_; 
wire _abc_15497_new_n3569_; 
wire _abc_15497_new_n3570_; 
wire _abc_15497_new_n3571_; 
wire _abc_15497_new_n3573_; 
wire _abc_15497_new_n3574_; 
wire _abc_15497_new_n3575_; 
wire _abc_15497_new_n3576_; 
wire _abc_15497_new_n3577_; 
wire _abc_15497_new_n3579_; 
wire _abc_15497_new_n3580_; 
wire _abc_15497_new_n3581_; 
wire _abc_15497_new_n3582_; 
wire _abc_15497_new_n3583_; 
wire _abc_15497_new_n3585_; 
wire _abc_15497_new_n3586_; 
wire _abc_15497_new_n3587_; 
wire _abc_15497_new_n3588_; 
wire _abc_15497_new_n3589_; 
wire _abc_15497_new_n3591_; 
wire _abc_15497_new_n3592_; 
wire _abc_15497_new_n3593_; 
wire _abc_15497_new_n3594_; 
wire _abc_15497_new_n3595_; 
wire _abc_15497_new_n3597_; 
wire _abc_15497_new_n3598_; 
wire _abc_15497_new_n3599_; 
wire _abc_15497_new_n3600_; 
wire _abc_15497_new_n3601_; 
wire _abc_15497_new_n3603_; 
wire _abc_15497_new_n3604_; 
wire _abc_15497_new_n3605_; 
wire _abc_15497_new_n3606_; 
wire _abc_15497_new_n3607_; 
wire _abc_15497_new_n3609_; 
wire _abc_15497_new_n3610_; 
wire _abc_15497_new_n3611_; 
wire _abc_15497_new_n3612_; 
wire _abc_15497_new_n3613_; 
wire _abc_15497_new_n3615_; 
wire _abc_15497_new_n3616_; 
wire _abc_15497_new_n3617_; 
wire _abc_15497_new_n3618_; 
wire _abc_15497_new_n3619_; 
wire _abc_15497_new_n3621_; 
wire _abc_15497_new_n3622_; 
wire _abc_15497_new_n3623_; 
wire _abc_15497_new_n3624_; 
wire _abc_15497_new_n3625_; 
wire _abc_15497_new_n3627_; 
wire _abc_15497_new_n3628_; 
wire _abc_15497_new_n3629_; 
wire _abc_15497_new_n3630_; 
wire _abc_15497_new_n3631_; 
wire _abc_15497_new_n3633_; 
wire _abc_15497_new_n3634_; 
wire _abc_15497_new_n3635_; 
wire _abc_15497_new_n3636_; 
wire _abc_15497_new_n3637_; 
wire _abc_15497_new_n3639_; 
wire _abc_15497_new_n3640_; 
wire _abc_15497_new_n3641_; 
wire _abc_15497_new_n3642_; 
wire _abc_15497_new_n3643_; 
wire _abc_15497_new_n3645_; 
wire _abc_15497_new_n3646_; 
wire _abc_15497_new_n3647_; 
wire _abc_15497_new_n3648_; 
wire _abc_15497_new_n3649_; 
wire _abc_15497_new_n3651_; 
wire _abc_15497_new_n3652_; 
wire _abc_15497_new_n3653_; 
wire _abc_15497_new_n3654_; 
wire _abc_15497_new_n3655_; 
wire _abc_15497_new_n3657_; 
wire _abc_15497_new_n3658_; 
wire _abc_15497_new_n3659_; 
wire _abc_15497_new_n3660_; 
wire _abc_15497_new_n3661_; 
wire _abc_15497_new_n3663_; 
wire _abc_15497_new_n3664_; 
wire _abc_15497_new_n3665_; 
wire _abc_15497_new_n3666_; 
wire _abc_15497_new_n3667_; 
wire _abc_15497_new_n3669_; 
wire _abc_15497_new_n3670_; 
wire _abc_15497_new_n3671_; 
wire _abc_15497_new_n3672_; 
wire _abc_15497_new_n3673_; 
wire _abc_15497_new_n3675_; 
wire _abc_15497_new_n3676_; 
wire _abc_15497_new_n3677_; 
wire _abc_15497_new_n3678_; 
wire _abc_15497_new_n3679_; 
wire _abc_15497_new_n3681_; 
wire _abc_15497_new_n3682_; 
wire _abc_15497_new_n3683_; 
wire _abc_15497_new_n3684_; 
wire _abc_15497_new_n3685_; 
wire _abc_15497_new_n3687_; 
wire _abc_15497_new_n3688_; 
wire _abc_15497_new_n3689_; 
wire _abc_15497_new_n3690_; 
wire _abc_15497_new_n3691_; 
wire _abc_15497_new_n3693_; 
wire _abc_15497_new_n3694_; 
wire _abc_15497_new_n3695_; 
wire _abc_15497_new_n3696_; 
wire _abc_15497_new_n3697_; 
wire _abc_15497_new_n3699_; 
wire _abc_15497_new_n3700_; 
wire _abc_15497_new_n3701_; 
wire _abc_15497_new_n3702_; 
wire _abc_15497_new_n3703_; 
wire _abc_15497_new_n3705_; 
wire _abc_15497_new_n3706_; 
wire _abc_15497_new_n3707_; 
wire _abc_15497_new_n3708_; 
wire _abc_15497_new_n3709_; 
wire _abc_15497_new_n3711_; 
wire _abc_15497_new_n3712_; 
wire _abc_15497_new_n3713_; 
wire _abc_15497_new_n3714_; 
wire _abc_15497_new_n3716_; 
wire _abc_15497_new_n3717_; 
wire _abc_15497_new_n3718_; 
wire _abc_15497_new_n3719_; 
wire _abc_15497_new_n3721_; 
wire _abc_15497_new_n3722_; 
wire _abc_15497_new_n3723_; 
wire _abc_15497_new_n3724_; 
wire _abc_15497_new_n3725_; 
wire _abc_15497_new_n3727_; 
wire _abc_15497_new_n3728_; 
wire _abc_15497_new_n3729_; 
wire _abc_15497_new_n3730_; 
wire _abc_15497_new_n3731_; 
wire _abc_15497_new_n3733_; 
wire _abc_15497_new_n3734_; 
wire _abc_15497_new_n3735_; 
wire _abc_15497_new_n3736_; 
wire _abc_15497_new_n3738_; 
wire _abc_15497_new_n3739_; 
wire _abc_15497_new_n3740_; 
wire _abc_15497_new_n3741_; 
wire _abc_15497_new_n3742_; 
wire _abc_15497_new_n3743_; 
wire _abc_15497_new_n3744_; 
wire _abc_15497_new_n3745_; 
wire _abc_15497_new_n3746_; 
wire _abc_15497_new_n3747_; 
wire _abc_15497_new_n3748_; 
wire _abc_15497_new_n3749_; 
wire _abc_15497_new_n3750_; 
wire _abc_15497_new_n3751_; 
wire _abc_15497_new_n3752_; 
wire _abc_15497_new_n3753_; 
wire _abc_15497_new_n3754_; 
wire _abc_15497_new_n3755_; 
wire _abc_15497_new_n3756_; 
wire _abc_15497_new_n3757_; 
wire _abc_15497_new_n3758_; 
wire _abc_15497_new_n3759_; 
wire _abc_15497_new_n3760_; 
wire _abc_15497_new_n3761_; 
wire _abc_15497_new_n3762_; 
wire _abc_15497_new_n3763_; 
wire _abc_15497_new_n3764_; 
wire _abc_15497_new_n3765_; 
wire _abc_15497_new_n3766_; 
wire _abc_15497_new_n3767_; 
wire _abc_15497_new_n3768_; 
wire _abc_15497_new_n3769_; 
wire _abc_15497_new_n3770_; 
wire _abc_15497_new_n3771_; 
wire _abc_15497_new_n3772_; 
wire _abc_15497_new_n3773_; 
wire _abc_15497_new_n3774_; 
wire _abc_15497_new_n3775_; 
wire _abc_15497_new_n3776_; 
wire _abc_15497_new_n3777_; 
wire _abc_15497_new_n3778_; 
wire _abc_15497_new_n3779_; 
wire _abc_15497_new_n3780_; 
wire _abc_15497_new_n3781_; 
wire _abc_15497_new_n3782_; 
wire _abc_15497_new_n3783_; 
wire _abc_15497_new_n3784_; 
wire _abc_15497_new_n3785_; 
wire _abc_15497_new_n3786_; 
wire _abc_15497_new_n3787_; 
wire _abc_15497_new_n3788_; 
wire _abc_15497_new_n3789_; 
wire _abc_15497_new_n3790_; 
wire _abc_15497_new_n3791_; 
wire _abc_15497_new_n3792_; 
wire _abc_15497_new_n3793_; 
wire _abc_15497_new_n3794_; 
wire _abc_15497_new_n3795_; 
wire _abc_15497_new_n3796_; 
wire _abc_15497_new_n3797_; 
wire _abc_15497_new_n3798_; 
wire _abc_15497_new_n3799_; 
wire _abc_15497_new_n3800_; 
wire _abc_15497_new_n3801_; 
wire _abc_15497_new_n3802_; 
wire _abc_15497_new_n3803_; 
wire _abc_15497_new_n3804_; 
wire _abc_15497_new_n3805_; 
wire _abc_15497_new_n3806_; 
wire _abc_15497_new_n3807_; 
wire _abc_15497_new_n3808_; 
wire _abc_15497_new_n3809_; 
wire _abc_15497_new_n3810_; 
wire _abc_15497_new_n3811_; 
wire _abc_15497_new_n3812_; 
wire _abc_15497_new_n3813_; 
wire _abc_15497_new_n3814_; 
wire _abc_15497_new_n3815_; 
wire _abc_15497_new_n3816_; 
wire _abc_15497_new_n3817_; 
wire _abc_15497_new_n3818_; 
wire _abc_15497_new_n3819_; 
wire _abc_15497_new_n3820_; 
wire _abc_15497_new_n3821_; 
wire _abc_15497_new_n3823_; 
wire _abc_15497_new_n3824_; 
wire _abc_15497_new_n3825_; 
wire _abc_15497_new_n3826_; 
wire _abc_15497_new_n3827_; 
wire _abc_15497_new_n3828_; 
wire _abc_15497_new_n3829_; 
wire _abc_15497_new_n3830_; 
wire _abc_15497_new_n3831_; 
wire _abc_15497_new_n3832_; 
wire _abc_15497_new_n3833_; 
wire _abc_15497_new_n3834_; 
wire _abc_15497_new_n3835_; 
wire _abc_15497_new_n3836_; 
wire _abc_15497_new_n3837_; 
wire _abc_15497_new_n3838_; 
wire _abc_15497_new_n3839_; 
wire _abc_15497_new_n3840_; 
wire _abc_15497_new_n3841_; 
wire _abc_15497_new_n3842_; 
wire _abc_15497_new_n3843_; 
wire _abc_15497_new_n3844_; 
wire _abc_15497_new_n3845_; 
wire _abc_15497_new_n3846_; 
wire _abc_15497_new_n3847_; 
wire _abc_15497_new_n3848_; 
wire _abc_15497_new_n3849_; 
wire _abc_15497_new_n3850_; 
wire _abc_15497_new_n3851_; 
wire _abc_15497_new_n3852_; 
wire _abc_15497_new_n3853_; 
wire _abc_15497_new_n3854_; 
wire _abc_15497_new_n3855_; 
wire _abc_15497_new_n3856_; 
wire _abc_15497_new_n3857_; 
wire _abc_15497_new_n3858_; 
wire _abc_15497_new_n3859_; 
wire _abc_15497_new_n3860_; 
wire _abc_15497_new_n3861_; 
wire _abc_15497_new_n3862_; 
wire _abc_15497_new_n3863_; 
wire _abc_15497_new_n3864_; 
wire _abc_15497_new_n3865_; 
wire _abc_15497_new_n3866_; 
wire _abc_15497_new_n3867_; 
wire _abc_15497_new_n3868_; 
wire _abc_15497_new_n3869_; 
wire _abc_15497_new_n3870_; 
wire _abc_15497_new_n3871_; 
wire _abc_15497_new_n3872_; 
wire _abc_15497_new_n3873_; 
wire _abc_15497_new_n3874_; 
wire _abc_15497_new_n3875_; 
wire _abc_15497_new_n3876_; 
wire _abc_15497_new_n3877_; 
wire _abc_15497_new_n3878_; 
wire _abc_15497_new_n3879_; 
wire _abc_15497_new_n3880_; 
wire _abc_15497_new_n3881_; 
wire _abc_15497_new_n3882_; 
wire _abc_15497_new_n3883_; 
wire _abc_15497_new_n3884_; 
wire _abc_15497_new_n3885_; 
wire _abc_15497_new_n3886_; 
wire _abc_15497_new_n3887_; 
wire _abc_15497_new_n3888_; 
wire _abc_15497_new_n3889_; 
wire _abc_15497_new_n3890_; 
wire _abc_15497_new_n3891_; 
wire _abc_15497_new_n3892_; 
wire _abc_15497_new_n3893_; 
wire _abc_15497_new_n3895_; 
wire _abc_15497_new_n3896_; 
wire _abc_15497_new_n3897_; 
wire _abc_15497_new_n3898_; 
wire _abc_15497_new_n3899_; 
wire _abc_15497_new_n3900_; 
wire _abc_15497_new_n3901_; 
wire _abc_15497_new_n3902_; 
wire _abc_15497_new_n3903_; 
wire _abc_15497_new_n3904_; 
wire _abc_15497_new_n3905_; 
wire _abc_15497_new_n3906_; 
wire _abc_15497_new_n3907_; 
wire _abc_15497_new_n3908_; 
wire _abc_15497_new_n3909_; 
wire _abc_15497_new_n3910_; 
wire _abc_15497_new_n3911_; 
wire _abc_15497_new_n3912_; 
wire _abc_15497_new_n3913_; 
wire _abc_15497_new_n3914_; 
wire _abc_15497_new_n3915_; 
wire _abc_15497_new_n3916_; 
wire _abc_15497_new_n3917_; 
wire _abc_15497_new_n3918_; 
wire _abc_15497_new_n3919_; 
wire _abc_15497_new_n3920_; 
wire _abc_15497_new_n3921_; 
wire _abc_15497_new_n3922_; 
wire _abc_15497_new_n3923_; 
wire _abc_15497_new_n3924_; 
wire _abc_15497_new_n3925_; 
wire _abc_15497_new_n3926_; 
wire _abc_15497_new_n3927_; 
wire _abc_15497_new_n3928_; 
wire _abc_15497_new_n3929_; 
wire _abc_15497_new_n3930_; 
wire _abc_15497_new_n3931_; 
wire _abc_15497_new_n3932_; 
wire _abc_15497_new_n3933_; 
wire _abc_15497_new_n3934_; 
wire _abc_15497_new_n3935_; 
wire _abc_15497_new_n3936_; 
wire _abc_15497_new_n3937_; 
wire _abc_15497_new_n3938_; 
wire _abc_15497_new_n3939_; 
wire _abc_15497_new_n3940_; 
wire _abc_15497_new_n3941_; 
wire _abc_15497_new_n3942_; 
wire _abc_15497_new_n3943_; 
wire _abc_15497_new_n3944_; 
wire _abc_15497_new_n3945_; 
wire _abc_15497_new_n3946_; 
wire _abc_15497_new_n3947_; 
wire _abc_15497_new_n3948_; 
wire _abc_15497_new_n3949_; 
wire _abc_15497_new_n3950_; 
wire _abc_15497_new_n3951_; 
wire _abc_15497_new_n3952_; 
wire _abc_15497_new_n3953_; 
wire _abc_15497_new_n3954_; 
wire _abc_15497_new_n3955_; 
wire _abc_15497_new_n3956_; 
wire _abc_15497_new_n3957_; 
wire _abc_15497_new_n3958_; 
wire _abc_15497_new_n3959_; 
wire _abc_15497_new_n3960_; 
wire _abc_15497_new_n3961_; 
wire _abc_15497_new_n3962_; 
wire _abc_15497_new_n3963_; 
wire _abc_15497_new_n3964_; 
wire _abc_15497_new_n3965_; 
wire _abc_15497_new_n3966_; 
wire _abc_15497_new_n3967_; 
wire _abc_15497_new_n3968_; 
wire _abc_15497_new_n3969_; 
wire _abc_15497_new_n3970_; 
wire _abc_15497_new_n3971_; 
wire _abc_15497_new_n3972_; 
wire _abc_15497_new_n3973_; 
wire _abc_15497_new_n3974_; 
wire _abc_15497_new_n3975_; 
wire _abc_15497_new_n3976_; 
wire _abc_15497_new_n3977_; 
wire _abc_15497_new_n3978_; 
wire _abc_15497_new_n3980_; 
wire _abc_15497_new_n3981_; 
wire _abc_15497_new_n3982_; 
wire _abc_15497_new_n3983_; 
wire _abc_15497_new_n3984_; 
wire _abc_15497_new_n3985_; 
wire _abc_15497_new_n3986_; 
wire _abc_15497_new_n3987_; 
wire _abc_15497_new_n3988_; 
wire _abc_15497_new_n3989_; 
wire _abc_15497_new_n3990_; 
wire _abc_15497_new_n3991_; 
wire _abc_15497_new_n3992_; 
wire _abc_15497_new_n3993_; 
wire _abc_15497_new_n3994_; 
wire _abc_15497_new_n3995_; 
wire _abc_15497_new_n3996_; 
wire _abc_15497_new_n3997_; 
wire _abc_15497_new_n3998_; 
wire _abc_15497_new_n3999_; 
wire _abc_15497_new_n4000_; 
wire _abc_15497_new_n4001_; 
wire _abc_15497_new_n4002_; 
wire _abc_15497_new_n4003_; 
wire _abc_15497_new_n4004_; 
wire _abc_15497_new_n4005_; 
wire _abc_15497_new_n4006_; 
wire _abc_15497_new_n4007_; 
wire _abc_15497_new_n4008_; 
wire _abc_15497_new_n4009_; 
wire _abc_15497_new_n4010_; 
wire _abc_15497_new_n4011_; 
wire _abc_15497_new_n4012_; 
wire _abc_15497_new_n4013_; 
wire _abc_15497_new_n4014_; 
wire _abc_15497_new_n4015_; 
wire _abc_15497_new_n4016_; 
wire _abc_15497_new_n4017_; 
wire _abc_15497_new_n4018_; 
wire _abc_15497_new_n4019_; 
wire _abc_15497_new_n4020_; 
wire _abc_15497_new_n4021_; 
wire _abc_15497_new_n4022_; 
wire _abc_15497_new_n4023_; 
wire _abc_15497_new_n4024_; 
wire _abc_15497_new_n4025_; 
wire _abc_15497_new_n4026_; 
wire _abc_15497_new_n4027_; 
wire _abc_15497_new_n4028_; 
wire _abc_15497_new_n4029_; 
wire _abc_15497_new_n4030_; 
wire _abc_15497_new_n4031_; 
wire _abc_15497_new_n4032_; 
wire _abc_15497_new_n4033_; 
wire _abc_15497_new_n4034_; 
wire _abc_15497_new_n4035_; 
wire _abc_15497_new_n4036_; 
wire _abc_15497_new_n4037_; 
wire _abc_15497_new_n4038_; 
wire _abc_15497_new_n4039_; 
wire _abc_15497_new_n4040_; 
wire _abc_15497_new_n4041_; 
wire _abc_15497_new_n4042_; 
wire _abc_15497_new_n4043_; 
wire _abc_15497_new_n4044_; 
wire _abc_15497_new_n4045_; 
wire _abc_15497_new_n4046_; 
wire _abc_15497_new_n4047_; 
wire _abc_15497_new_n4048_; 
wire _abc_15497_new_n4049_; 
wire _abc_15497_new_n4050_; 
wire _abc_15497_new_n4051_; 
wire _abc_15497_new_n4053_; 
wire _abc_15497_new_n4054_; 
wire _abc_15497_new_n4055_; 
wire _abc_15497_new_n4056_; 
wire _abc_15497_new_n4057_; 
wire _abc_15497_new_n4058_; 
wire _abc_15497_new_n4059_; 
wire _abc_15497_new_n4060_; 
wire _abc_15497_new_n4061_; 
wire _abc_15497_new_n4062_; 
wire _abc_15497_new_n4063_; 
wire _abc_15497_new_n4064_; 
wire _abc_15497_new_n4065_; 
wire _abc_15497_new_n4066_; 
wire _abc_15497_new_n4067_; 
wire _abc_15497_new_n4068_; 
wire _abc_15497_new_n4069_; 
wire _abc_15497_new_n4070_; 
wire _abc_15497_new_n4071_; 
wire _abc_15497_new_n4072_; 
wire _abc_15497_new_n4073_; 
wire _abc_15497_new_n4074_; 
wire _abc_15497_new_n4075_; 
wire _abc_15497_new_n4076_; 
wire _abc_15497_new_n4077_; 
wire _abc_15497_new_n4078_; 
wire _abc_15497_new_n4079_; 
wire _abc_15497_new_n4080_; 
wire _abc_15497_new_n4081_; 
wire _abc_15497_new_n4082_; 
wire _abc_15497_new_n4083_; 
wire _abc_15497_new_n4084_; 
wire _abc_15497_new_n4085_; 
wire _abc_15497_new_n4086_; 
wire _abc_15497_new_n4087_; 
wire _abc_15497_new_n4088_; 
wire _abc_15497_new_n4089_; 
wire _abc_15497_new_n4090_; 
wire _abc_15497_new_n4091_; 
wire _abc_15497_new_n4092_; 
wire _abc_15497_new_n4093_; 
wire _abc_15497_new_n4094_; 
wire _abc_15497_new_n4095_; 
wire _abc_15497_new_n4096_; 
wire _abc_15497_new_n4097_; 
wire _abc_15497_new_n4098_; 
wire _abc_15497_new_n4099_; 
wire _abc_15497_new_n4100_; 
wire _abc_15497_new_n4101_; 
wire _abc_15497_new_n4102_; 
wire _abc_15497_new_n4103_; 
wire _abc_15497_new_n4104_; 
wire _abc_15497_new_n4105_; 
wire _abc_15497_new_n4106_; 
wire _abc_15497_new_n4107_; 
wire _abc_15497_new_n4108_; 
wire _abc_15497_new_n4109_; 
wire _abc_15497_new_n4110_; 
wire _abc_15497_new_n4111_; 
wire _abc_15497_new_n4112_; 
wire _abc_15497_new_n4113_; 
wire _abc_15497_new_n4114_; 
wire _abc_15497_new_n4115_; 
wire _abc_15497_new_n4116_; 
wire _abc_15497_new_n4117_; 
wire _abc_15497_new_n4118_; 
wire _abc_15497_new_n4119_; 
wire _abc_15497_new_n4120_; 
wire _abc_15497_new_n4121_; 
wire _abc_15497_new_n4122_; 
wire _abc_15497_new_n4123_; 
wire _abc_15497_new_n4124_; 
wire _abc_15497_new_n4125_; 
wire _abc_15497_new_n4126_; 
wire _abc_15497_new_n4127_; 
wire _abc_15497_new_n4128_; 
wire _abc_15497_new_n4129_; 
wire _abc_15497_new_n4130_; 
wire _abc_15497_new_n4131_; 
wire _abc_15497_new_n4132_; 
wire _abc_15497_new_n4133_; 
wire _abc_15497_new_n4134_; 
wire _abc_15497_new_n4136_; 
wire _abc_15497_new_n4137_; 
wire _abc_15497_new_n4138_; 
wire _abc_15497_new_n4139_; 
wire _abc_15497_new_n4140_; 
wire _abc_15497_new_n4141_; 
wire _abc_15497_new_n4142_; 
wire _abc_15497_new_n4143_; 
wire _abc_15497_new_n4144_; 
wire _abc_15497_new_n4145_; 
wire _abc_15497_new_n4146_; 
wire _abc_15497_new_n4147_; 
wire _abc_15497_new_n4148_; 
wire _abc_15497_new_n4149_; 
wire _abc_15497_new_n4150_; 
wire _abc_15497_new_n4151_; 
wire _abc_15497_new_n4152_; 
wire _abc_15497_new_n4153_; 
wire _abc_15497_new_n4154_; 
wire _abc_15497_new_n4155_; 
wire _abc_15497_new_n4156_; 
wire _abc_15497_new_n4157_; 
wire _abc_15497_new_n4158_; 
wire _abc_15497_new_n4159_; 
wire _abc_15497_new_n4160_; 
wire _abc_15497_new_n4161_; 
wire _abc_15497_new_n4162_; 
wire _abc_15497_new_n4163_; 
wire _abc_15497_new_n4164_; 
wire _abc_15497_new_n4165_; 
wire _abc_15497_new_n4166_; 
wire _abc_15497_new_n4167_; 
wire _abc_15497_new_n4168_; 
wire _abc_15497_new_n4169_; 
wire _abc_15497_new_n4170_; 
wire _abc_15497_new_n4171_; 
wire _abc_15497_new_n4172_; 
wire _abc_15497_new_n4173_; 
wire _abc_15497_new_n4174_; 
wire _abc_15497_new_n4175_; 
wire _abc_15497_new_n4176_; 
wire _abc_15497_new_n4177_; 
wire _abc_15497_new_n4178_; 
wire _abc_15497_new_n4179_; 
wire _abc_15497_new_n4180_; 
wire _abc_15497_new_n4181_; 
wire _abc_15497_new_n4182_; 
wire _abc_15497_new_n4183_; 
wire _abc_15497_new_n4184_; 
wire _abc_15497_new_n4185_; 
wire _abc_15497_new_n4186_; 
wire _abc_15497_new_n4187_; 
wire _abc_15497_new_n4188_; 
wire _abc_15497_new_n4189_; 
wire _abc_15497_new_n4190_; 
wire _abc_15497_new_n4191_; 
wire _abc_15497_new_n4192_; 
wire _abc_15497_new_n4193_; 
wire _abc_15497_new_n4194_; 
wire _abc_15497_new_n4195_; 
wire _abc_15497_new_n4196_; 
wire _abc_15497_new_n4197_; 
wire _abc_15497_new_n4198_; 
wire _abc_15497_new_n4199_; 
wire _abc_15497_new_n4200_; 
wire _abc_15497_new_n4201_; 
wire _abc_15497_new_n4202_; 
wire _abc_15497_new_n4203_; 
wire _abc_15497_new_n4204_; 
wire _abc_15497_new_n4205_; 
wire _abc_15497_new_n4206_; 
wire _abc_15497_new_n4207_; 
wire _abc_15497_new_n4208_; 
wire _abc_15497_new_n4209_; 
wire _abc_15497_new_n4210_; 
wire _abc_15497_new_n4211_; 
wire _abc_15497_new_n4212_; 
wire _abc_15497_new_n4214_; 
wire _abc_15497_new_n4215_; 
wire _abc_15497_new_n4216_; 
wire _abc_15497_new_n4217_; 
wire _abc_15497_new_n4218_; 
wire _abc_15497_new_n4219_; 
wire _abc_15497_new_n4220_; 
wire _abc_15497_new_n4221_; 
wire _abc_15497_new_n4222_; 
wire _abc_15497_new_n4223_; 
wire _abc_15497_new_n4224_; 
wire _abc_15497_new_n4225_; 
wire _abc_15497_new_n4226_; 
wire _abc_15497_new_n4227_; 
wire _abc_15497_new_n4228_; 
wire _abc_15497_new_n4229_; 
wire _abc_15497_new_n4230_; 
wire _abc_15497_new_n4231_; 
wire _abc_15497_new_n4232_; 
wire _abc_15497_new_n4233_; 
wire _abc_15497_new_n4234_; 
wire _abc_15497_new_n4235_; 
wire _abc_15497_new_n4236_; 
wire _abc_15497_new_n4237_; 
wire _abc_15497_new_n4238_; 
wire _abc_15497_new_n4239_; 
wire _abc_15497_new_n4240_; 
wire _abc_15497_new_n4241_; 
wire _abc_15497_new_n4242_; 
wire _abc_15497_new_n4243_; 
wire _abc_15497_new_n4244_; 
wire _abc_15497_new_n4245_; 
wire _abc_15497_new_n4246_; 
wire _abc_15497_new_n4247_; 
wire _abc_15497_new_n4248_; 
wire _abc_15497_new_n4249_; 
wire _abc_15497_new_n4250_; 
wire _abc_15497_new_n4251_; 
wire _abc_15497_new_n4252_; 
wire _abc_15497_new_n4253_; 
wire _abc_15497_new_n4254_; 
wire _abc_15497_new_n4255_; 
wire _abc_15497_new_n4256_; 
wire _abc_15497_new_n4257_; 
wire _abc_15497_new_n4258_; 
wire _abc_15497_new_n4259_; 
wire _abc_15497_new_n4260_; 
wire _abc_15497_new_n4261_; 
wire _abc_15497_new_n4262_; 
wire _abc_15497_new_n4263_; 
wire _abc_15497_new_n4264_; 
wire _abc_15497_new_n4265_; 
wire _abc_15497_new_n4266_; 
wire _abc_15497_new_n4267_; 
wire _abc_15497_new_n4268_; 
wire _abc_15497_new_n4269_; 
wire _abc_15497_new_n4270_; 
wire _abc_15497_new_n4271_; 
wire _abc_15497_new_n4272_; 
wire _abc_15497_new_n4273_; 
wire _abc_15497_new_n4274_; 
wire _abc_15497_new_n4275_; 
wire _abc_15497_new_n4276_; 
wire _abc_15497_new_n4277_; 
wire _abc_15497_new_n4278_; 
wire _abc_15497_new_n4279_; 
wire _abc_15497_new_n4280_; 
wire _abc_15497_new_n4281_; 
wire _abc_15497_new_n4282_; 
wire _abc_15497_new_n4283_; 
wire _abc_15497_new_n4284_; 
wire _abc_15497_new_n4285_; 
wire _abc_15497_new_n4286_; 
wire _abc_15497_new_n4287_; 
wire _abc_15497_new_n4288_; 
wire _abc_15497_new_n4289_; 
wire _abc_15497_new_n4290_; 
wire _abc_15497_new_n4291_; 
wire _abc_15497_new_n4292_; 
wire _abc_15497_new_n4293_; 
wire _abc_15497_new_n4294_; 
wire _abc_15497_new_n4295_; 
wire _abc_15497_new_n4296_; 
wire _abc_15497_new_n4298_; 
wire _abc_15497_new_n4299_; 
wire _abc_15497_new_n4300_; 
wire _abc_15497_new_n4301_; 
wire _abc_15497_new_n4302_; 
wire _abc_15497_new_n4303_; 
wire _abc_15497_new_n4304_; 
wire _abc_15497_new_n4305_; 
wire _abc_15497_new_n4306_; 
wire _abc_15497_new_n4307_; 
wire _abc_15497_new_n4308_; 
wire _abc_15497_new_n4309_; 
wire _abc_15497_new_n4310_; 
wire _abc_15497_new_n4311_; 
wire _abc_15497_new_n4312_; 
wire _abc_15497_new_n4313_; 
wire _abc_15497_new_n4314_; 
wire _abc_15497_new_n4315_; 
wire _abc_15497_new_n4316_; 
wire _abc_15497_new_n4317_; 
wire _abc_15497_new_n4318_; 
wire _abc_15497_new_n4319_; 
wire _abc_15497_new_n4320_; 
wire _abc_15497_new_n4321_; 
wire _abc_15497_new_n4322_; 
wire _abc_15497_new_n4323_; 
wire _abc_15497_new_n4324_; 
wire _abc_15497_new_n4325_; 
wire _abc_15497_new_n4326_; 
wire _abc_15497_new_n4327_; 
wire _abc_15497_new_n4328_; 
wire _abc_15497_new_n4329_; 
wire _abc_15497_new_n4330_; 
wire _abc_15497_new_n4331_; 
wire _abc_15497_new_n4332_; 
wire _abc_15497_new_n4333_; 
wire _abc_15497_new_n4334_; 
wire _abc_15497_new_n4335_; 
wire _abc_15497_new_n4336_; 
wire _abc_15497_new_n4337_; 
wire _abc_15497_new_n4338_; 
wire _abc_15497_new_n4339_; 
wire _abc_15497_new_n4340_; 
wire _abc_15497_new_n4341_; 
wire _abc_15497_new_n4342_; 
wire _abc_15497_new_n4343_; 
wire _abc_15497_new_n4344_; 
wire _abc_15497_new_n4345_; 
wire _abc_15497_new_n4346_; 
wire _abc_15497_new_n4347_; 
wire _abc_15497_new_n4348_; 
wire _abc_15497_new_n4349_; 
wire _abc_15497_new_n4350_; 
wire _abc_15497_new_n4351_; 
wire _abc_15497_new_n4352_; 
wire _abc_15497_new_n4353_; 
wire _abc_15497_new_n4354_; 
wire _abc_15497_new_n4355_; 
wire _abc_15497_new_n4356_; 
wire _abc_15497_new_n4357_; 
wire _abc_15497_new_n4358_; 
wire _abc_15497_new_n4359_; 
wire _abc_15497_new_n4360_; 
wire _abc_15497_new_n4361_; 
wire _abc_15497_new_n4362_; 
wire _abc_15497_new_n4363_; 
wire _abc_15497_new_n4364_; 
wire _abc_15497_new_n4366_; 
wire _abc_15497_new_n4367_; 
wire _abc_15497_new_n4368_; 
wire _abc_15497_new_n4369_; 
wire _abc_15497_new_n4370_; 
wire _abc_15497_new_n4371_; 
wire _abc_15497_new_n4372_; 
wire _abc_15497_new_n4373_; 
wire _abc_15497_new_n4374_; 
wire _abc_15497_new_n4375_; 
wire _abc_15497_new_n4376_; 
wire _abc_15497_new_n4377_; 
wire _abc_15497_new_n4378_; 
wire _abc_15497_new_n4379_; 
wire _abc_15497_new_n4380_; 
wire _abc_15497_new_n4381_; 
wire _abc_15497_new_n4382_; 
wire _abc_15497_new_n4383_; 
wire _abc_15497_new_n4384_; 
wire _abc_15497_new_n4385_; 
wire _abc_15497_new_n4386_; 
wire _abc_15497_new_n4387_; 
wire _abc_15497_new_n4388_; 
wire _abc_15497_new_n4389_; 
wire _abc_15497_new_n4390_; 
wire _abc_15497_new_n4391_; 
wire _abc_15497_new_n4392_; 
wire _abc_15497_new_n4393_; 
wire _abc_15497_new_n4394_; 
wire _abc_15497_new_n4395_; 
wire _abc_15497_new_n4396_; 
wire _abc_15497_new_n4397_; 
wire _abc_15497_new_n4398_; 
wire _abc_15497_new_n4399_; 
wire _abc_15497_new_n4400_; 
wire _abc_15497_new_n4401_; 
wire _abc_15497_new_n4402_; 
wire _abc_15497_new_n4403_; 
wire _abc_15497_new_n4404_; 
wire _abc_15497_new_n4405_; 
wire _abc_15497_new_n4406_; 
wire _abc_15497_new_n4407_; 
wire _abc_15497_new_n4408_; 
wire _abc_15497_new_n4409_; 
wire _abc_15497_new_n4410_; 
wire _abc_15497_new_n4411_; 
wire _abc_15497_new_n4412_; 
wire _abc_15497_new_n4413_; 
wire _abc_15497_new_n4414_; 
wire _abc_15497_new_n4415_; 
wire _abc_15497_new_n4416_; 
wire _abc_15497_new_n4417_; 
wire _abc_15497_new_n4418_; 
wire _abc_15497_new_n4419_; 
wire _abc_15497_new_n4420_; 
wire _abc_15497_new_n4421_; 
wire _abc_15497_new_n4422_; 
wire _abc_15497_new_n4423_; 
wire _abc_15497_new_n4424_; 
wire _abc_15497_new_n4425_; 
wire _abc_15497_new_n4426_; 
wire _abc_15497_new_n4427_; 
wire _abc_15497_new_n4428_; 
wire _abc_15497_new_n4429_; 
wire _abc_15497_new_n4430_; 
wire _abc_15497_new_n4431_; 
wire _abc_15497_new_n4432_; 
wire _abc_15497_new_n4433_; 
wire _abc_15497_new_n4434_; 
wire _abc_15497_new_n4435_; 
wire _abc_15497_new_n4436_; 
wire _abc_15497_new_n4437_; 
wire _abc_15497_new_n4438_; 
wire _abc_15497_new_n4439_; 
wire _abc_15497_new_n4440_; 
wire _abc_15497_new_n4441_; 
wire _abc_15497_new_n4442_; 
wire _abc_15497_new_n4443_; 
wire _abc_15497_new_n4444_; 
wire _abc_15497_new_n4445_; 
wire _abc_15497_new_n4446_; 
wire _abc_15497_new_n4447_; 
wire _abc_15497_new_n4448_; 
wire _abc_15497_new_n4449_; 
wire _abc_15497_new_n4450_; 
wire _abc_15497_new_n4452_; 
wire _abc_15497_new_n4453_; 
wire _abc_15497_new_n4454_; 
wire _abc_15497_new_n4455_; 
wire _abc_15497_new_n4456_; 
wire _abc_15497_new_n4457_; 
wire _abc_15497_new_n4458_; 
wire _abc_15497_new_n4459_; 
wire _abc_15497_new_n4460_; 
wire _abc_15497_new_n4461_; 
wire _abc_15497_new_n4462_; 
wire _abc_15497_new_n4463_; 
wire _abc_15497_new_n4464_; 
wire _abc_15497_new_n4465_; 
wire _abc_15497_new_n4466_; 
wire _abc_15497_new_n4467_; 
wire _abc_15497_new_n4468_; 
wire _abc_15497_new_n4469_; 
wire _abc_15497_new_n4470_; 
wire _abc_15497_new_n4471_; 
wire _abc_15497_new_n4472_; 
wire _abc_15497_new_n4473_; 
wire _abc_15497_new_n4474_; 
wire _abc_15497_new_n4475_; 
wire _abc_15497_new_n4476_; 
wire _abc_15497_new_n4477_; 
wire _abc_15497_new_n4478_; 
wire _abc_15497_new_n4479_; 
wire _abc_15497_new_n4480_; 
wire _abc_15497_new_n4481_; 
wire _abc_15497_new_n4482_; 
wire _abc_15497_new_n4483_; 
wire _abc_15497_new_n4484_; 
wire _abc_15497_new_n4485_; 
wire _abc_15497_new_n4486_; 
wire _abc_15497_new_n4487_; 
wire _abc_15497_new_n4488_; 
wire _abc_15497_new_n4489_; 
wire _abc_15497_new_n4490_; 
wire _abc_15497_new_n4491_; 
wire _abc_15497_new_n4492_; 
wire _abc_15497_new_n4493_; 
wire _abc_15497_new_n4494_; 
wire _abc_15497_new_n4495_; 
wire _abc_15497_new_n4496_; 
wire _abc_15497_new_n4497_; 
wire _abc_15497_new_n4498_; 
wire _abc_15497_new_n4499_; 
wire _abc_15497_new_n4500_; 
wire _abc_15497_new_n4501_; 
wire _abc_15497_new_n4502_; 
wire _abc_15497_new_n4503_; 
wire _abc_15497_new_n4504_; 
wire _abc_15497_new_n4505_; 
wire _abc_15497_new_n4506_; 
wire _abc_15497_new_n4507_; 
wire _abc_15497_new_n4508_; 
wire _abc_15497_new_n4509_; 
wire _abc_15497_new_n4510_; 
wire _abc_15497_new_n4511_; 
wire _abc_15497_new_n4512_; 
wire _abc_15497_new_n4513_; 
wire _abc_15497_new_n4514_; 
wire _abc_15497_new_n4515_; 
wire _abc_15497_new_n4516_; 
wire _abc_15497_new_n4517_; 
wire _abc_15497_new_n4518_; 
wire _abc_15497_new_n4519_; 
wire _abc_15497_new_n4520_; 
wire _abc_15497_new_n4521_; 
wire _abc_15497_new_n4522_; 
wire _abc_15497_new_n4523_; 
wire _abc_15497_new_n4524_; 
wire _abc_15497_new_n4525_; 
wire _abc_15497_new_n4527_; 
wire _abc_15497_new_n4528_; 
wire _abc_15497_new_n4529_; 
wire _abc_15497_new_n4530_; 
wire _abc_15497_new_n4531_; 
wire _abc_15497_new_n4532_; 
wire _abc_15497_new_n4533_; 
wire _abc_15497_new_n4534_; 
wire _abc_15497_new_n4535_; 
wire _abc_15497_new_n4536_; 
wire _abc_15497_new_n4537_; 
wire _abc_15497_new_n4538_; 
wire _abc_15497_new_n4539_; 
wire _abc_15497_new_n4540_; 
wire _abc_15497_new_n4541_; 
wire _abc_15497_new_n4542_; 
wire _abc_15497_new_n4543_; 
wire _abc_15497_new_n4544_; 
wire _abc_15497_new_n4545_; 
wire _abc_15497_new_n4546_; 
wire _abc_15497_new_n4547_; 
wire _abc_15497_new_n4548_; 
wire _abc_15497_new_n4549_; 
wire _abc_15497_new_n4550_; 
wire _abc_15497_new_n4551_; 
wire _abc_15497_new_n4552_; 
wire _abc_15497_new_n4553_; 
wire _abc_15497_new_n4554_; 
wire _abc_15497_new_n4555_; 
wire _abc_15497_new_n4556_; 
wire _abc_15497_new_n4557_; 
wire _abc_15497_new_n4558_; 
wire _abc_15497_new_n4559_; 
wire _abc_15497_new_n4560_; 
wire _abc_15497_new_n4561_; 
wire _abc_15497_new_n4562_; 
wire _abc_15497_new_n4563_; 
wire _abc_15497_new_n4564_; 
wire _abc_15497_new_n4565_; 
wire _abc_15497_new_n4566_; 
wire _abc_15497_new_n4567_; 
wire _abc_15497_new_n4568_; 
wire _abc_15497_new_n4569_; 
wire _abc_15497_new_n4570_; 
wire _abc_15497_new_n4571_; 
wire _abc_15497_new_n4572_; 
wire _abc_15497_new_n4573_; 
wire _abc_15497_new_n4574_; 
wire _abc_15497_new_n4575_; 
wire _abc_15497_new_n4576_; 
wire _abc_15497_new_n4577_; 
wire _abc_15497_new_n4578_; 
wire _abc_15497_new_n4579_; 
wire _abc_15497_new_n4580_; 
wire _abc_15497_new_n4581_; 
wire _abc_15497_new_n4582_; 
wire _abc_15497_new_n4583_; 
wire _abc_15497_new_n4584_; 
wire _abc_15497_new_n4585_; 
wire _abc_15497_new_n4586_; 
wire _abc_15497_new_n4587_; 
wire _abc_15497_new_n4588_; 
wire _abc_15497_new_n4589_; 
wire _abc_15497_new_n4590_; 
wire _abc_15497_new_n4591_; 
wire _abc_15497_new_n4592_; 
wire _abc_15497_new_n4593_; 
wire _abc_15497_new_n4594_; 
wire _abc_15497_new_n4595_; 
wire _abc_15497_new_n4596_; 
wire _abc_15497_new_n4597_; 
wire _abc_15497_new_n4598_; 
wire _abc_15497_new_n4599_; 
wire _abc_15497_new_n4600_; 
wire _abc_15497_new_n4601_; 
wire _abc_15497_new_n4602_; 
wire _abc_15497_new_n4603_; 
wire _abc_15497_new_n4604_; 
wire _abc_15497_new_n4605_; 
wire _abc_15497_new_n4606_; 
wire _abc_15497_new_n4607_; 
wire _abc_15497_new_n4608_; 
wire _abc_15497_new_n4609_; 
wire _abc_15497_new_n4611_; 
wire _abc_15497_new_n4612_; 
wire _abc_15497_new_n4613_; 
wire _abc_15497_new_n4614_; 
wire _abc_15497_new_n4615_; 
wire _abc_15497_new_n4616_; 
wire _abc_15497_new_n4617_; 
wire _abc_15497_new_n4618_; 
wire _abc_15497_new_n4619_; 
wire _abc_15497_new_n4620_; 
wire _abc_15497_new_n4621_; 
wire _abc_15497_new_n4622_; 
wire _abc_15497_new_n4623_; 
wire _abc_15497_new_n4624_; 
wire _abc_15497_new_n4625_; 
wire _abc_15497_new_n4626_; 
wire _abc_15497_new_n4627_; 
wire _abc_15497_new_n4628_; 
wire _abc_15497_new_n4629_; 
wire _abc_15497_new_n4630_; 
wire _abc_15497_new_n4631_; 
wire _abc_15497_new_n4632_; 
wire _abc_15497_new_n4633_; 
wire _abc_15497_new_n4634_; 
wire _abc_15497_new_n4635_; 
wire _abc_15497_new_n4636_; 
wire _abc_15497_new_n4637_; 
wire _abc_15497_new_n4638_; 
wire _abc_15497_new_n4639_; 
wire _abc_15497_new_n4640_; 
wire _abc_15497_new_n4641_; 
wire _abc_15497_new_n4642_; 
wire _abc_15497_new_n4643_; 
wire _abc_15497_new_n4644_; 
wire _abc_15497_new_n4645_; 
wire _abc_15497_new_n4646_; 
wire _abc_15497_new_n4647_; 
wire _abc_15497_new_n4648_; 
wire _abc_15497_new_n4649_; 
wire _abc_15497_new_n4650_; 
wire _abc_15497_new_n4651_; 
wire _abc_15497_new_n4652_; 
wire _abc_15497_new_n4653_; 
wire _abc_15497_new_n4654_; 
wire _abc_15497_new_n4655_; 
wire _abc_15497_new_n4656_; 
wire _abc_15497_new_n4657_; 
wire _abc_15497_new_n4658_; 
wire _abc_15497_new_n4659_; 
wire _abc_15497_new_n4660_; 
wire _abc_15497_new_n4661_; 
wire _abc_15497_new_n4662_; 
wire _abc_15497_new_n4663_; 
wire _abc_15497_new_n4664_; 
wire _abc_15497_new_n4665_; 
wire _abc_15497_new_n4666_; 
wire _abc_15497_new_n4667_; 
wire _abc_15497_new_n4668_; 
wire _abc_15497_new_n4669_; 
wire _abc_15497_new_n4670_; 
wire _abc_15497_new_n4671_; 
wire _abc_15497_new_n4672_; 
wire _abc_15497_new_n4673_; 
wire _abc_15497_new_n4674_; 
wire _abc_15497_new_n4675_; 
wire _abc_15497_new_n4676_; 
wire _abc_15497_new_n4677_; 
wire _abc_15497_new_n4678_; 
wire _abc_15497_new_n4679_; 
wire _abc_15497_new_n4680_; 
wire _abc_15497_new_n4681_; 
wire _abc_15497_new_n4682_; 
wire _abc_15497_new_n4683_; 
wire _abc_15497_new_n4684_; 
wire _abc_15497_new_n4685_; 
wire _abc_15497_new_n4686_; 
wire _abc_15497_new_n4688_; 
wire _abc_15497_new_n4689_; 
wire _abc_15497_new_n4690_; 
wire _abc_15497_new_n4691_; 
wire _abc_15497_new_n4692_; 
wire _abc_15497_new_n4693_; 
wire _abc_15497_new_n4694_; 
wire _abc_15497_new_n4695_; 
wire _abc_15497_new_n4696_; 
wire _abc_15497_new_n4697_; 
wire _abc_15497_new_n4698_; 
wire _abc_15497_new_n4699_; 
wire _abc_15497_new_n4700_; 
wire _abc_15497_new_n4701_; 
wire _abc_15497_new_n4702_; 
wire _abc_15497_new_n4703_; 
wire _abc_15497_new_n4704_; 
wire _abc_15497_new_n4705_; 
wire _abc_15497_new_n4706_; 
wire _abc_15497_new_n4707_; 
wire _abc_15497_new_n4708_; 
wire _abc_15497_new_n4709_; 
wire _abc_15497_new_n4710_; 
wire _abc_15497_new_n4711_; 
wire _abc_15497_new_n4712_; 
wire _abc_15497_new_n4713_; 
wire _abc_15497_new_n4714_; 
wire _abc_15497_new_n4715_; 
wire _abc_15497_new_n4716_; 
wire _abc_15497_new_n4717_; 
wire _abc_15497_new_n4718_; 
wire _abc_15497_new_n4719_; 
wire _abc_15497_new_n4720_; 
wire _abc_15497_new_n4721_; 
wire _abc_15497_new_n4722_; 
wire _abc_15497_new_n4723_; 
wire _abc_15497_new_n4724_; 
wire _abc_15497_new_n4725_; 
wire _abc_15497_new_n4726_; 
wire _abc_15497_new_n4727_; 
wire _abc_15497_new_n4728_; 
wire _abc_15497_new_n4729_; 
wire _abc_15497_new_n4730_; 
wire _abc_15497_new_n4731_; 
wire _abc_15497_new_n4732_; 
wire _abc_15497_new_n4733_; 
wire _abc_15497_new_n4734_; 
wire _abc_15497_new_n4735_; 
wire _abc_15497_new_n4736_; 
wire _abc_15497_new_n4737_; 
wire _abc_15497_new_n4738_; 
wire _abc_15497_new_n4739_; 
wire _abc_15497_new_n4740_; 
wire _abc_15497_new_n4741_; 
wire _abc_15497_new_n4742_; 
wire _abc_15497_new_n4743_; 
wire _abc_15497_new_n4744_; 
wire _abc_15497_new_n4745_; 
wire _abc_15497_new_n4746_; 
wire _abc_15497_new_n4747_; 
wire _abc_15497_new_n4748_; 
wire _abc_15497_new_n4749_; 
wire _abc_15497_new_n4750_; 
wire _abc_15497_new_n4751_; 
wire _abc_15497_new_n4752_; 
wire _abc_15497_new_n4753_; 
wire _abc_15497_new_n4754_; 
wire _abc_15497_new_n4755_; 
wire _abc_15497_new_n4756_; 
wire _abc_15497_new_n4757_; 
wire _abc_15497_new_n4758_; 
wire _abc_15497_new_n4759_; 
wire _abc_15497_new_n4760_; 
wire _abc_15497_new_n4761_; 
wire _abc_15497_new_n4762_; 
wire _abc_15497_new_n4763_; 
wire _abc_15497_new_n4764_; 
wire _abc_15497_new_n4765_; 
wire _abc_15497_new_n4766_; 
wire _abc_15497_new_n4767_; 
wire _abc_15497_new_n4768_; 
wire _abc_15497_new_n4769_; 
wire _abc_15497_new_n4771_; 
wire _abc_15497_new_n4772_; 
wire _abc_15497_new_n4773_; 
wire _abc_15497_new_n4774_; 
wire _abc_15497_new_n4775_; 
wire _abc_15497_new_n4776_; 
wire _abc_15497_new_n4777_; 
wire _abc_15497_new_n4778_; 
wire _abc_15497_new_n4779_; 
wire _abc_15497_new_n4780_; 
wire _abc_15497_new_n4781_; 
wire _abc_15497_new_n4782_; 
wire _abc_15497_new_n4783_; 
wire _abc_15497_new_n4784_; 
wire _abc_15497_new_n4785_; 
wire _abc_15497_new_n4786_; 
wire _abc_15497_new_n4787_; 
wire _abc_15497_new_n4788_; 
wire _abc_15497_new_n4789_; 
wire _abc_15497_new_n4790_; 
wire _abc_15497_new_n4791_; 
wire _abc_15497_new_n4792_; 
wire _abc_15497_new_n4793_; 
wire _abc_15497_new_n4794_; 
wire _abc_15497_new_n4795_; 
wire _abc_15497_new_n4796_; 
wire _abc_15497_new_n4797_; 
wire _abc_15497_new_n4798_; 
wire _abc_15497_new_n4799_; 
wire _abc_15497_new_n4800_; 
wire _abc_15497_new_n4801_; 
wire _abc_15497_new_n4802_; 
wire _abc_15497_new_n4803_; 
wire _abc_15497_new_n4804_; 
wire _abc_15497_new_n4805_; 
wire _abc_15497_new_n4806_; 
wire _abc_15497_new_n4807_; 
wire _abc_15497_new_n4808_; 
wire _abc_15497_new_n4809_; 
wire _abc_15497_new_n4810_; 
wire _abc_15497_new_n4811_; 
wire _abc_15497_new_n4812_; 
wire _abc_15497_new_n4813_; 
wire _abc_15497_new_n4814_; 
wire _abc_15497_new_n4815_; 
wire _abc_15497_new_n4816_; 
wire _abc_15497_new_n4817_; 
wire _abc_15497_new_n4818_; 
wire _abc_15497_new_n4819_; 
wire _abc_15497_new_n4820_; 
wire _abc_15497_new_n4821_; 
wire _abc_15497_new_n4822_; 
wire _abc_15497_new_n4823_; 
wire _abc_15497_new_n4824_; 
wire _abc_15497_new_n4825_; 
wire _abc_15497_new_n4826_; 
wire _abc_15497_new_n4827_; 
wire _abc_15497_new_n4828_; 
wire _abc_15497_new_n4829_; 
wire _abc_15497_new_n4830_; 
wire _abc_15497_new_n4831_; 
wire _abc_15497_new_n4832_; 
wire _abc_15497_new_n4833_; 
wire _abc_15497_new_n4834_; 
wire _abc_15497_new_n4835_; 
wire _abc_15497_new_n4836_; 
wire _abc_15497_new_n4837_; 
wire _abc_15497_new_n4838_; 
wire _abc_15497_new_n4839_; 
wire _abc_15497_new_n4840_; 
wire _abc_15497_new_n4841_; 
wire _abc_15497_new_n4842_; 
wire _abc_15497_new_n4844_; 
wire _abc_15497_new_n4845_; 
wire _abc_15497_new_n4846_; 
wire _abc_15497_new_n4847_; 
wire _abc_15497_new_n4848_; 
wire _abc_15497_new_n4849_; 
wire _abc_15497_new_n4850_; 
wire _abc_15497_new_n4851_; 
wire _abc_15497_new_n4852_; 
wire _abc_15497_new_n4853_; 
wire _abc_15497_new_n4854_; 
wire _abc_15497_new_n4855_; 
wire _abc_15497_new_n4856_; 
wire _abc_15497_new_n4857_; 
wire _abc_15497_new_n4858_; 
wire _abc_15497_new_n4859_; 
wire _abc_15497_new_n4860_; 
wire _abc_15497_new_n4861_; 
wire _abc_15497_new_n4862_; 
wire _abc_15497_new_n4863_; 
wire _abc_15497_new_n4864_; 
wire _abc_15497_new_n4865_; 
wire _abc_15497_new_n4866_; 
wire _abc_15497_new_n4867_; 
wire _abc_15497_new_n4868_; 
wire _abc_15497_new_n4869_; 
wire _abc_15497_new_n4870_; 
wire _abc_15497_new_n4871_; 
wire _abc_15497_new_n4872_; 
wire _abc_15497_new_n4873_; 
wire _abc_15497_new_n4874_; 
wire _abc_15497_new_n4875_; 
wire _abc_15497_new_n4876_; 
wire _abc_15497_new_n4877_; 
wire _abc_15497_new_n4878_; 
wire _abc_15497_new_n4879_; 
wire _abc_15497_new_n4880_; 
wire _abc_15497_new_n4881_; 
wire _abc_15497_new_n4882_; 
wire _abc_15497_new_n4883_; 
wire _abc_15497_new_n4884_; 
wire _abc_15497_new_n4885_; 
wire _abc_15497_new_n4886_; 
wire _abc_15497_new_n4887_; 
wire _abc_15497_new_n4888_; 
wire _abc_15497_new_n4889_; 
wire _abc_15497_new_n4890_; 
wire _abc_15497_new_n4891_; 
wire _abc_15497_new_n4892_; 
wire _abc_15497_new_n4893_; 
wire _abc_15497_new_n4894_; 
wire _abc_15497_new_n4895_; 
wire _abc_15497_new_n4896_; 
wire _abc_15497_new_n4897_; 
wire _abc_15497_new_n4898_; 
wire _abc_15497_new_n4899_; 
wire _abc_15497_new_n4900_; 
wire _abc_15497_new_n4901_; 
wire _abc_15497_new_n4902_; 
wire _abc_15497_new_n4903_; 
wire _abc_15497_new_n4904_; 
wire _abc_15497_new_n4905_; 
wire _abc_15497_new_n4906_; 
wire _abc_15497_new_n4907_; 
wire _abc_15497_new_n4908_; 
wire _abc_15497_new_n4909_; 
wire _abc_15497_new_n4910_; 
wire _abc_15497_new_n4911_; 
wire _abc_15497_new_n4912_; 
wire _abc_15497_new_n4913_; 
wire _abc_15497_new_n4914_; 
wire _abc_15497_new_n4915_; 
wire _abc_15497_new_n4916_; 
wire _abc_15497_new_n4917_; 
wire _abc_15497_new_n4918_; 
wire _abc_15497_new_n4919_; 
wire _abc_15497_new_n4920_; 
wire _abc_15497_new_n4921_; 
wire _abc_15497_new_n4923_; 
wire _abc_15497_new_n4924_; 
wire _abc_15497_new_n4925_; 
wire _abc_15497_new_n4926_; 
wire _abc_15497_new_n4927_; 
wire _abc_15497_new_n4928_; 
wire _abc_15497_new_n4929_; 
wire _abc_15497_new_n4930_; 
wire _abc_15497_new_n4931_; 
wire _abc_15497_new_n4932_; 
wire _abc_15497_new_n4933_; 
wire _abc_15497_new_n4934_; 
wire _abc_15497_new_n4935_; 
wire _abc_15497_new_n4936_; 
wire _abc_15497_new_n4937_; 
wire _abc_15497_new_n4938_; 
wire _abc_15497_new_n4939_; 
wire _abc_15497_new_n4940_; 
wire _abc_15497_new_n4941_; 
wire _abc_15497_new_n4942_; 
wire _abc_15497_new_n4943_; 
wire _abc_15497_new_n4944_; 
wire _abc_15497_new_n4945_; 
wire _abc_15497_new_n4946_; 
wire _abc_15497_new_n4947_; 
wire _abc_15497_new_n4948_; 
wire _abc_15497_new_n4949_; 
wire _abc_15497_new_n4950_; 
wire _abc_15497_new_n4951_; 
wire _abc_15497_new_n4952_; 
wire _abc_15497_new_n4953_; 
wire _abc_15497_new_n4954_; 
wire _abc_15497_new_n4955_; 
wire _abc_15497_new_n4956_; 
wire _abc_15497_new_n4957_; 
wire _abc_15497_new_n4958_; 
wire _abc_15497_new_n4959_; 
wire _abc_15497_new_n4960_; 
wire _abc_15497_new_n4961_; 
wire _abc_15497_new_n4962_; 
wire _abc_15497_new_n4963_; 
wire _abc_15497_new_n4964_; 
wire _abc_15497_new_n4965_; 
wire _abc_15497_new_n4966_; 
wire _abc_15497_new_n4967_; 
wire _abc_15497_new_n4968_; 
wire _abc_15497_new_n4969_; 
wire _abc_15497_new_n4970_; 
wire _abc_15497_new_n4971_; 
wire _abc_15497_new_n4972_; 
wire _abc_15497_new_n4973_; 
wire _abc_15497_new_n4974_; 
wire _abc_15497_new_n4975_; 
wire _abc_15497_new_n4976_; 
wire _abc_15497_new_n4977_; 
wire _abc_15497_new_n4978_; 
wire _abc_15497_new_n4979_; 
wire _abc_15497_new_n4980_; 
wire _abc_15497_new_n4981_; 
wire _abc_15497_new_n4982_; 
wire _abc_15497_new_n4983_; 
wire _abc_15497_new_n4984_; 
wire _abc_15497_new_n4985_; 
wire _abc_15497_new_n4986_; 
wire _abc_15497_new_n4987_; 
wire _abc_15497_new_n4988_; 
wire _abc_15497_new_n4989_; 
wire _abc_15497_new_n4990_; 
wire _abc_15497_new_n4991_; 
wire _abc_15497_new_n4992_; 
wire _abc_15497_new_n4993_; 
wire _abc_15497_new_n4994_; 
wire _abc_15497_new_n4996_; 
wire _abc_15497_new_n4997_; 
wire _abc_15497_new_n4998_; 
wire _abc_15497_new_n4999_; 
wire _abc_15497_new_n5000_; 
wire _abc_15497_new_n5001_; 
wire _abc_15497_new_n5002_; 
wire _abc_15497_new_n5003_; 
wire _abc_15497_new_n5004_; 
wire _abc_15497_new_n5005_; 
wire _abc_15497_new_n5006_; 
wire _abc_15497_new_n5007_; 
wire _abc_15497_new_n5008_; 
wire _abc_15497_new_n5009_; 
wire _abc_15497_new_n5010_; 
wire _abc_15497_new_n5011_; 
wire _abc_15497_new_n5012_; 
wire _abc_15497_new_n5013_; 
wire _abc_15497_new_n5014_; 
wire _abc_15497_new_n5015_; 
wire _abc_15497_new_n5016_; 
wire _abc_15497_new_n5017_; 
wire _abc_15497_new_n5018_; 
wire _abc_15497_new_n5019_; 
wire _abc_15497_new_n5020_; 
wire _abc_15497_new_n5021_; 
wire _abc_15497_new_n5022_; 
wire _abc_15497_new_n5023_; 
wire _abc_15497_new_n5024_; 
wire _abc_15497_new_n5025_; 
wire _abc_15497_new_n5026_; 
wire _abc_15497_new_n5027_; 
wire _abc_15497_new_n5028_; 
wire _abc_15497_new_n5029_; 
wire _abc_15497_new_n5030_; 
wire _abc_15497_new_n5031_; 
wire _abc_15497_new_n5032_; 
wire _abc_15497_new_n5033_; 
wire _abc_15497_new_n5034_; 
wire _abc_15497_new_n5035_; 
wire _abc_15497_new_n5036_; 
wire _abc_15497_new_n5037_; 
wire _abc_15497_new_n5038_; 
wire _abc_15497_new_n5039_; 
wire _abc_15497_new_n5040_; 
wire _abc_15497_new_n5041_; 
wire _abc_15497_new_n5042_; 
wire _abc_15497_new_n5043_; 
wire _abc_15497_new_n5044_; 
wire _abc_15497_new_n5045_; 
wire _abc_15497_new_n5046_; 
wire _abc_15497_new_n5047_; 
wire _abc_15497_new_n5048_; 
wire _abc_15497_new_n5049_; 
wire _abc_15497_new_n5050_; 
wire _abc_15497_new_n5051_; 
wire _abc_15497_new_n5052_; 
wire _abc_15497_new_n5053_; 
wire _abc_15497_new_n5054_; 
wire _abc_15497_new_n5055_; 
wire _abc_15497_new_n5056_; 
wire _abc_15497_new_n5057_; 
wire _abc_15497_new_n5058_; 
wire _abc_15497_new_n5059_; 
wire _abc_15497_new_n5060_; 
wire _abc_15497_new_n5061_; 
wire _abc_15497_new_n5062_; 
wire _abc_15497_new_n5063_; 
wire _abc_15497_new_n5064_; 
wire _abc_15497_new_n5065_; 
wire _abc_15497_new_n5066_; 
wire _abc_15497_new_n5067_; 
wire _abc_15497_new_n5068_; 
wire _abc_15497_new_n5069_; 
wire _abc_15497_new_n5070_; 
wire _abc_15497_new_n5071_; 
wire _abc_15497_new_n5072_; 
wire _abc_15497_new_n5073_; 
wire _abc_15497_new_n5074_; 
wire _abc_15497_new_n5076_; 
wire _abc_15497_new_n5077_; 
wire _abc_15497_new_n5078_; 
wire _abc_15497_new_n5079_; 
wire _abc_15497_new_n5080_; 
wire _abc_15497_new_n5081_; 
wire _abc_15497_new_n5082_; 
wire _abc_15497_new_n5083_; 
wire _abc_15497_new_n5084_; 
wire _abc_15497_new_n5085_; 
wire _abc_15497_new_n5086_; 
wire _abc_15497_new_n5087_; 
wire _abc_15497_new_n5088_; 
wire _abc_15497_new_n5089_; 
wire _abc_15497_new_n5090_; 
wire _abc_15497_new_n5091_; 
wire _abc_15497_new_n5092_; 
wire _abc_15497_new_n5093_; 
wire _abc_15497_new_n5094_; 
wire _abc_15497_new_n5095_; 
wire _abc_15497_new_n5096_; 
wire _abc_15497_new_n5097_; 
wire _abc_15497_new_n5098_; 
wire _abc_15497_new_n5099_; 
wire _abc_15497_new_n5100_; 
wire _abc_15497_new_n5101_; 
wire _abc_15497_new_n5102_; 
wire _abc_15497_new_n5103_; 
wire _abc_15497_new_n5104_; 
wire _abc_15497_new_n5105_; 
wire _abc_15497_new_n5106_; 
wire _abc_15497_new_n5107_; 
wire _abc_15497_new_n5108_; 
wire _abc_15497_new_n5109_; 
wire _abc_15497_new_n5110_; 
wire _abc_15497_new_n5111_; 
wire _abc_15497_new_n5112_; 
wire _abc_15497_new_n5113_; 
wire _abc_15497_new_n5114_; 
wire _abc_15497_new_n5115_; 
wire _abc_15497_new_n5116_; 
wire _abc_15497_new_n5117_; 
wire _abc_15497_new_n5118_; 
wire _abc_15497_new_n5119_; 
wire _abc_15497_new_n5120_; 
wire _abc_15497_new_n5121_; 
wire _abc_15497_new_n5122_; 
wire _abc_15497_new_n5123_; 
wire _abc_15497_new_n5124_; 
wire _abc_15497_new_n5125_; 
wire _abc_15497_new_n5126_; 
wire _abc_15497_new_n5127_; 
wire _abc_15497_new_n5128_; 
wire _abc_15497_new_n5129_; 
wire _abc_15497_new_n5130_; 
wire _abc_15497_new_n5131_; 
wire _abc_15497_new_n5132_; 
wire _abc_15497_new_n5133_; 
wire _abc_15497_new_n5134_; 
wire _abc_15497_new_n5135_; 
wire _abc_15497_new_n5136_; 
wire _abc_15497_new_n5137_; 
wire _abc_15497_new_n5138_; 
wire _abc_15497_new_n5139_; 
wire _abc_15497_new_n5140_; 
wire _abc_15497_new_n5141_; 
wire _abc_15497_new_n5142_; 
wire _abc_15497_new_n5143_; 
wire _abc_15497_new_n5144_; 
wire _abc_15497_new_n5146_; 
wire _abc_15497_new_n5147_; 
wire _abc_15497_new_n5148_; 
wire _abc_15497_new_n5149_; 
wire _abc_15497_new_n5150_; 
wire _abc_15497_new_n5151_; 
wire _abc_15497_new_n5152_; 
wire _abc_15497_new_n5153_; 
wire _abc_15497_new_n5154_; 
wire _abc_15497_new_n5155_; 
wire _abc_15497_new_n5156_; 
wire _abc_15497_new_n5157_; 
wire _abc_15497_new_n5158_; 
wire _abc_15497_new_n5159_; 
wire _abc_15497_new_n5160_; 
wire _abc_15497_new_n5161_; 
wire _abc_15497_new_n5162_; 
wire _abc_15497_new_n5163_; 
wire _abc_15497_new_n5164_; 
wire _abc_15497_new_n5165_; 
wire _abc_15497_new_n5166_; 
wire _abc_15497_new_n5167_; 
wire _abc_15497_new_n5168_; 
wire _abc_15497_new_n5169_; 
wire _abc_15497_new_n5170_; 
wire _abc_15497_new_n5171_; 
wire _abc_15497_new_n5172_; 
wire _abc_15497_new_n5173_; 
wire _abc_15497_new_n5174_; 
wire _abc_15497_new_n5175_; 
wire _abc_15497_new_n5176_; 
wire _abc_15497_new_n5177_; 
wire _abc_15497_new_n5178_; 
wire _abc_15497_new_n5179_; 
wire _abc_15497_new_n5180_; 
wire _abc_15497_new_n5181_; 
wire _abc_15497_new_n5182_; 
wire _abc_15497_new_n5183_; 
wire _abc_15497_new_n5184_; 
wire _abc_15497_new_n5185_; 
wire _abc_15497_new_n5186_; 
wire _abc_15497_new_n5187_; 
wire _abc_15497_new_n5188_; 
wire _abc_15497_new_n5189_; 
wire _abc_15497_new_n5190_; 
wire _abc_15497_new_n5191_; 
wire _abc_15497_new_n5192_; 
wire _abc_15497_new_n5193_; 
wire _abc_15497_new_n5194_; 
wire _abc_15497_new_n5195_; 
wire _abc_15497_new_n5196_; 
wire _abc_15497_new_n5197_; 
wire _abc_15497_new_n5198_; 
wire _abc_15497_new_n5199_; 
wire _abc_15497_new_n5200_; 
wire _abc_15497_new_n5201_; 
wire _abc_15497_new_n5202_; 
wire _abc_15497_new_n5203_; 
wire _abc_15497_new_n5204_; 
wire _abc_15497_new_n5205_; 
wire _abc_15497_new_n5206_; 
wire _abc_15497_new_n5207_; 
wire _abc_15497_new_n5208_; 
wire _abc_15497_new_n5209_; 
wire _abc_15497_new_n5210_; 
wire _abc_15497_new_n5211_; 
wire _abc_15497_new_n5212_; 
wire _abc_15497_new_n5213_; 
wire _abc_15497_new_n5215_; 
wire _abc_15497_new_n5216_; 
wire _abc_15497_new_n5217_; 
wire _abc_15497_new_n5218_; 
wire _abc_15497_new_n5219_; 
wire _abc_15497_new_n5220_; 
wire _abc_15497_new_n5221_; 
wire _abc_15497_new_n5222_; 
wire _abc_15497_new_n5223_; 
wire _abc_15497_new_n5224_; 
wire _abc_15497_new_n5225_; 
wire _abc_15497_new_n5226_; 
wire _abc_15497_new_n5227_; 
wire _abc_15497_new_n5228_; 
wire _abc_15497_new_n5229_; 
wire _abc_15497_new_n5230_; 
wire _abc_15497_new_n5231_; 
wire _abc_15497_new_n5232_; 
wire _abc_15497_new_n5233_; 
wire _abc_15497_new_n5234_; 
wire _abc_15497_new_n5235_; 
wire _abc_15497_new_n5236_; 
wire _abc_15497_new_n5237_; 
wire _abc_15497_new_n5238_; 
wire _abc_15497_new_n5239_; 
wire _abc_15497_new_n5240_; 
wire _abc_15497_new_n5241_; 
wire _abc_15497_new_n5242_; 
wire _abc_15497_new_n5243_; 
wire _abc_15497_new_n5244_; 
wire _abc_15497_new_n5245_; 
wire _abc_15497_new_n5246_; 
wire _abc_15497_new_n5247_; 
wire _abc_15497_new_n5248_; 
wire _abc_15497_new_n5249_; 
wire _abc_15497_new_n5250_; 
wire _abc_15497_new_n5251_; 
wire _abc_15497_new_n5252_; 
wire _abc_15497_new_n5253_; 
wire _abc_15497_new_n5254_; 
wire _abc_15497_new_n5255_; 
wire _abc_15497_new_n5256_; 
wire _abc_15497_new_n5257_; 
wire _abc_15497_new_n5258_; 
wire _abc_15497_new_n5259_; 
wire _abc_15497_new_n5260_; 
wire _abc_15497_new_n5261_; 
wire _abc_15497_new_n5262_; 
wire _abc_15497_new_n5263_; 
wire _abc_15497_new_n5264_; 
wire _abc_15497_new_n5265_; 
wire _abc_15497_new_n5266_; 
wire _abc_15497_new_n5267_; 
wire _abc_15497_new_n5268_; 
wire _abc_15497_new_n5269_; 
wire _abc_15497_new_n5270_; 
wire _abc_15497_new_n5271_; 
wire _abc_15497_new_n5272_; 
wire _abc_15497_new_n5273_; 
wire _abc_15497_new_n5274_; 
wire _abc_15497_new_n5275_; 
wire _abc_15497_new_n5276_; 
wire _abc_15497_new_n5277_; 
wire _abc_15497_new_n5278_; 
wire _abc_15497_new_n5279_; 
wire _abc_15497_new_n5280_; 
wire _abc_15497_new_n5281_; 
wire _abc_15497_new_n5282_; 
wire _abc_15497_new_n5284_; 
wire _abc_15497_new_n5285_; 
wire _abc_15497_new_n5286_; 
wire _abc_15497_new_n5287_; 
wire _abc_15497_new_n5288_; 
wire _abc_15497_new_n5289_; 
wire _abc_15497_new_n5290_; 
wire _abc_15497_new_n5291_; 
wire _abc_15497_new_n5292_; 
wire _abc_15497_new_n5293_; 
wire _abc_15497_new_n5294_; 
wire _abc_15497_new_n5295_; 
wire _abc_15497_new_n5296_; 
wire _abc_15497_new_n5297_; 
wire _abc_15497_new_n5298_; 
wire _abc_15497_new_n5299_; 
wire _abc_15497_new_n5300_; 
wire _abc_15497_new_n5301_; 
wire _abc_15497_new_n5302_; 
wire _abc_15497_new_n5303_; 
wire _abc_15497_new_n5304_; 
wire _abc_15497_new_n5305_; 
wire _abc_15497_new_n5306_; 
wire _abc_15497_new_n5307_; 
wire _abc_15497_new_n5308_; 
wire _abc_15497_new_n5309_; 
wire _abc_15497_new_n5310_; 
wire _abc_15497_new_n5311_; 
wire _abc_15497_new_n5312_; 
wire _abc_15497_new_n5313_; 
wire _abc_15497_new_n5314_; 
wire _abc_15497_new_n5315_; 
wire _abc_15497_new_n5316_; 
wire _abc_15497_new_n5317_; 
wire _abc_15497_new_n5318_; 
wire _abc_15497_new_n5319_; 
wire _abc_15497_new_n5320_; 
wire _abc_15497_new_n5321_; 
wire _abc_15497_new_n5322_; 
wire _abc_15497_new_n5323_; 
wire _abc_15497_new_n5324_; 
wire _abc_15497_new_n5325_; 
wire _abc_15497_new_n5326_; 
wire _abc_15497_new_n5327_; 
wire _abc_15497_new_n5328_; 
wire _abc_15497_new_n5329_; 
wire _abc_15497_new_n5330_; 
wire _abc_15497_new_n5331_; 
wire _abc_15497_new_n5332_; 
wire _abc_15497_new_n5333_; 
wire _abc_15497_new_n5334_; 
wire _abc_15497_new_n5335_; 
wire _abc_15497_new_n5336_; 
wire _abc_15497_new_n5337_; 
wire _abc_15497_new_n5338_; 
wire _abc_15497_new_n5339_; 
wire _abc_15497_new_n5340_; 
wire _abc_15497_new_n5341_; 
wire _abc_15497_new_n5342_; 
wire _abc_15497_new_n5343_; 
wire _abc_15497_new_n5344_; 
wire _abc_15497_new_n5345_; 
wire _abc_15497_new_n5346_; 
wire _abc_15497_new_n5347_; 
wire _abc_15497_new_n5348_; 
wire _abc_15497_new_n5349_; 
wire _abc_15497_new_n5350_; 
wire _abc_15497_new_n5351_; 
wire _abc_15497_new_n5352_; 
wire _abc_15497_new_n5353_; 
wire _abc_15497_new_n5354_; 
wire _abc_15497_new_n5355_; 
wire _abc_15497_new_n5356_; 
wire _abc_15497_new_n5357_; 
wire _abc_15497_new_n5358_; 
wire _abc_15497_new_n5359_; 
wire _abc_15497_new_n5360_; 
wire _abc_15497_new_n5361_; 
wire _abc_15497_new_n5362_; 
wire _abc_15497_new_n5363_; 
wire _abc_15497_new_n5365_; 
wire _abc_15497_new_n5366_; 
wire _abc_15497_new_n5367_; 
wire _abc_15497_new_n5368_; 
wire _abc_15497_new_n5369_; 
wire _abc_15497_new_n5370_; 
wire _abc_15497_new_n5371_; 
wire _abc_15497_new_n5372_; 
wire _abc_15497_new_n5373_; 
wire _abc_15497_new_n5374_; 
wire _abc_15497_new_n5375_; 
wire _abc_15497_new_n5376_; 
wire _abc_15497_new_n5377_; 
wire _abc_15497_new_n5378_; 
wire _abc_15497_new_n5379_; 
wire _abc_15497_new_n5380_; 
wire _abc_15497_new_n5381_; 
wire _abc_15497_new_n5382_; 
wire _abc_15497_new_n5383_; 
wire _abc_15497_new_n5384_; 
wire _abc_15497_new_n5385_; 
wire _abc_15497_new_n5386_; 
wire _abc_15497_new_n5387_; 
wire _abc_15497_new_n5388_; 
wire _abc_15497_new_n5389_; 
wire _abc_15497_new_n5390_; 
wire _abc_15497_new_n5391_; 
wire _abc_15497_new_n5392_; 
wire _abc_15497_new_n5393_; 
wire _abc_15497_new_n5394_; 
wire _abc_15497_new_n5395_; 
wire _abc_15497_new_n5396_; 
wire _abc_15497_new_n5397_; 
wire _abc_15497_new_n5398_; 
wire _abc_15497_new_n5399_; 
wire _abc_15497_new_n5400_; 
wire _abc_15497_new_n5401_; 
wire _abc_15497_new_n5402_; 
wire _abc_15497_new_n5403_; 
wire _abc_15497_new_n5404_; 
wire _abc_15497_new_n5405_; 
wire _abc_15497_new_n5406_; 
wire _abc_15497_new_n5407_; 
wire _abc_15497_new_n5408_; 
wire _abc_15497_new_n5409_; 
wire _abc_15497_new_n5410_; 
wire _abc_15497_new_n5411_; 
wire _abc_15497_new_n5412_; 
wire _abc_15497_new_n5413_; 
wire _abc_15497_new_n5414_; 
wire _abc_15497_new_n5415_; 
wire _abc_15497_new_n5416_; 
wire _abc_15497_new_n5417_; 
wire _abc_15497_new_n5418_; 
wire _abc_15497_new_n5419_; 
wire _abc_15497_new_n5420_; 
wire _abc_15497_new_n5421_; 
wire _abc_15497_new_n5422_; 
wire _abc_15497_new_n5423_; 
wire _abc_15497_new_n5424_; 
wire _abc_15497_new_n5425_; 
wire _abc_15497_new_n5426_; 
wire _abc_15497_new_n5427_; 
wire _abc_15497_new_n5428_; 
wire _abc_15497_new_n5429_; 
wire _abc_15497_new_n5430_; 
wire _abc_15497_new_n5431_; 
wire _abc_15497_new_n5432_; 
wire _abc_15497_new_n5433_; 
wire _abc_15497_new_n5435_; 
wire _abc_15497_new_n5436_; 
wire _abc_15497_new_n5437_; 
wire _abc_15497_new_n5438_; 
wire _abc_15497_new_n5439_; 
wire _abc_15497_new_n5440_; 
wire _abc_15497_new_n5441_; 
wire _abc_15497_new_n5442_; 
wire _abc_15497_new_n5443_; 
wire _abc_15497_new_n5444_; 
wire _abc_15497_new_n5445_; 
wire _abc_15497_new_n5446_; 
wire _abc_15497_new_n5447_; 
wire _abc_15497_new_n5448_; 
wire _abc_15497_new_n5449_; 
wire _abc_15497_new_n5450_; 
wire _abc_15497_new_n5451_; 
wire _abc_15497_new_n5452_; 
wire _abc_15497_new_n5453_; 
wire _abc_15497_new_n5454_; 
wire _abc_15497_new_n5455_; 
wire _abc_15497_new_n5456_; 
wire _abc_15497_new_n5457_; 
wire _abc_15497_new_n5458_; 
wire _abc_15497_new_n5459_; 
wire _abc_15497_new_n5460_; 
wire _abc_15497_new_n5461_; 
wire _abc_15497_new_n5462_; 
wire _abc_15497_new_n5463_; 
wire _abc_15497_new_n5464_; 
wire _abc_15497_new_n5465_; 
wire _abc_15497_new_n5466_; 
wire _abc_15497_new_n5467_; 
wire _abc_15497_new_n5468_; 
wire _abc_15497_new_n5469_; 
wire _abc_15497_new_n5470_; 
wire _abc_15497_new_n5471_; 
wire _abc_15497_new_n5472_; 
wire _abc_15497_new_n5473_; 
wire _abc_15497_new_n5474_; 
wire _abc_15497_new_n5475_; 
wire _abc_15497_new_n5476_; 
wire _abc_15497_new_n5477_; 
wire _abc_15497_new_n5478_; 
wire _abc_15497_new_n5479_; 
wire _abc_15497_new_n5480_; 
wire _abc_15497_new_n5481_; 
wire _abc_15497_new_n5482_; 
wire _abc_15497_new_n5483_; 
wire _abc_15497_new_n5484_; 
wire _abc_15497_new_n5485_; 
wire _abc_15497_new_n5486_; 
wire _abc_15497_new_n5487_; 
wire _abc_15497_new_n5488_; 
wire _abc_15497_new_n5489_; 
wire _abc_15497_new_n5490_; 
wire _abc_15497_new_n5491_; 
wire _abc_15497_new_n5492_; 
wire _abc_15497_new_n5493_; 
wire _abc_15497_new_n5494_; 
wire _abc_15497_new_n5495_; 
wire _abc_15497_new_n5496_; 
wire _abc_15497_new_n5497_; 
wire _abc_15497_new_n5498_; 
wire _abc_15497_new_n5499_; 
wire _abc_15497_new_n5500_; 
wire _abc_15497_new_n5501_; 
wire _abc_15497_new_n5502_; 
wire _abc_15497_new_n5503_; 
wire _abc_15497_new_n5504_; 
wire _abc_15497_new_n5505_; 
wire _abc_15497_new_n5506_; 
wire _abc_15497_new_n5507_; 
wire _abc_15497_new_n5508_; 
wire _abc_15497_new_n5510_; 
wire _abc_15497_new_n5511_; 
wire _abc_15497_new_n5512_; 
wire _abc_15497_new_n5513_; 
wire _abc_15497_new_n5514_; 
wire _abc_15497_new_n5515_; 
wire _abc_15497_new_n5516_; 
wire _abc_15497_new_n5517_; 
wire _abc_15497_new_n5518_; 
wire _abc_15497_new_n5519_; 
wire _abc_15497_new_n5520_; 
wire _abc_15497_new_n5521_; 
wire _abc_15497_new_n5522_; 
wire _abc_15497_new_n5523_; 
wire _abc_15497_new_n5524_; 
wire _abc_15497_new_n5525_; 
wire _abc_15497_new_n5526_; 
wire _abc_15497_new_n5527_; 
wire _abc_15497_new_n5528_; 
wire _abc_15497_new_n5529_; 
wire _abc_15497_new_n5530_; 
wire _abc_15497_new_n5531_; 
wire _abc_15497_new_n5532_; 
wire _abc_15497_new_n5533_; 
wire _abc_15497_new_n5534_; 
wire _abc_15497_new_n5535_; 
wire _abc_15497_new_n5536_; 
wire _abc_15497_new_n5537_; 
wire _abc_15497_new_n5538_; 
wire _abc_15497_new_n5539_; 
wire _abc_15497_new_n5540_; 
wire _abc_15497_new_n5541_; 
wire _abc_15497_new_n5542_; 
wire _abc_15497_new_n5543_; 
wire _abc_15497_new_n5544_; 
wire _abc_15497_new_n5545_; 
wire _abc_15497_new_n5546_; 
wire _abc_15497_new_n5547_; 
wire _abc_15497_new_n5548_; 
wire _abc_15497_new_n5549_; 
wire _abc_15497_new_n5550_; 
wire _abc_15497_new_n5551_; 
wire _abc_15497_new_n5552_; 
wire _abc_15497_new_n5553_; 
wire _abc_15497_new_n5554_; 
wire _abc_15497_new_n5555_; 
wire _abc_15497_new_n5556_; 
wire _abc_15497_new_n5557_; 
wire _abc_15497_new_n5558_; 
wire _abc_15497_new_n5559_; 
wire _abc_15497_new_n5560_; 
wire _abc_15497_new_n5561_; 
wire _abc_15497_new_n5562_; 
wire _abc_15497_new_n5563_; 
wire _abc_15497_new_n5564_; 
wire _abc_15497_new_n5565_; 
wire _abc_15497_new_n5566_; 
wire _abc_15497_new_n5567_; 
wire _abc_15497_new_n5568_; 
wire _abc_15497_new_n5569_; 
wire _abc_15497_new_n5570_; 
wire _abc_15497_new_n5571_; 
wire _abc_15497_new_n5572_; 
wire _abc_15497_new_n5573_; 
wire _abc_15497_new_n5574_; 
wire _abc_15497_new_n5575_; 
wire _abc_15497_new_n5576_; 
wire _abc_15497_new_n5577_; 
wire _abc_15497_new_n5579_; 
wire _abc_15497_new_n5580_; 
wire _abc_15497_new_n5581_; 
wire _abc_15497_new_n5582_; 
wire _abc_15497_new_n5583_; 
wire _abc_15497_new_n5584_; 
wire _abc_15497_new_n5585_; 
wire _abc_15497_new_n5586_; 
wire _abc_15497_new_n5587_; 
wire _abc_15497_new_n5588_; 
wire _abc_15497_new_n5589_; 
wire _abc_15497_new_n5590_; 
wire _abc_15497_new_n5591_; 
wire _abc_15497_new_n5592_; 
wire _abc_15497_new_n5593_; 
wire _abc_15497_new_n5594_; 
wire _abc_15497_new_n5595_; 
wire _abc_15497_new_n5596_; 
wire _abc_15497_new_n5597_; 
wire _abc_15497_new_n5598_; 
wire _abc_15497_new_n5599_; 
wire _abc_15497_new_n5600_; 
wire _abc_15497_new_n5601_; 
wire _abc_15497_new_n5602_; 
wire _abc_15497_new_n5603_; 
wire _abc_15497_new_n5604_; 
wire _abc_15497_new_n5605_; 
wire _abc_15497_new_n5606_; 
wire _abc_15497_new_n5607_; 
wire _abc_15497_new_n5608_; 
wire _abc_15497_new_n5609_; 
wire _abc_15497_new_n5610_; 
wire _abc_15497_new_n5611_; 
wire _abc_15497_new_n5612_; 
wire _abc_15497_new_n5613_; 
wire _abc_15497_new_n5614_; 
wire _abc_15497_new_n5615_; 
wire _abc_15497_new_n5616_; 
wire _abc_15497_new_n5617_; 
wire _abc_15497_new_n5618_; 
wire _abc_15497_new_n5619_; 
wire _abc_15497_new_n5620_; 
wire _abc_15497_new_n5621_; 
wire _abc_15497_new_n5622_; 
wire _abc_15497_new_n5623_; 
wire _abc_15497_new_n5624_; 
wire _abc_15497_new_n5625_; 
wire _abc_15497_new_n5626_; 
wire _abc_15497_new_n5627_; 
wire _abc_15497_new_n5628_; 
wire _abc_15497_new_n5629_; 
wire _abc_15497_new_n5630_; 
wire _abc_15497_new_n5631_; 
wire _abc_15497_new_n5632_; 
wire _abc_15497_new_n5633_; 
wire _abc_15497_new_n5634_; 
wire _abc_15497_new_n5635_; 
wire _abc_15497_new_n5636_; 
wire _abc_15497_new_n5637_; 
wire _abc_15497_new_n5638_; 
wire _abc_15497_new_n5639_; 
wire _abc_15497_new_n5640_; 
wire _abc_15497_new_n5641_; 
wire _abc_15497_new_n5642_; 
wire _abc_15497_new_n5643_; 
wire _abc_15497_new_n5644_; 
wire _abc_15497_new_n5645_; 
wire _abc_15497_new_n5646_; 
wire _abc_15497_new_n5647_; 
wire _abc_15497_new_n5648_; 
wire _abc_15497_new_n5649_; 
wire _abc_15497_new_n5650_; 
wire _abc_15497_new_n5651_; 
wire _abc_15497_new_n5652_; 
wire _abc_15497_new_n5653_; 
wire _abc_15497_new_n5654_; 
wire _abc_15497_new_n5655_; 
wire _abc_15497_new_n5656_; 
wire _abc_15497_new_n5658_; 
wire _abc_15497_new_n5659_; 
wire _abc_15497_new_n5660_; 
wire _abc_15497_new_n5661_; 
wire _abc_15497_new_n5662_; 
wire _abc_15497_new_n5663_; 
wire _abc_15497_new_n5664_; 
wire _abc_15497_new_n5665_; 
wire _abc_15497_new_n5666_; 
wire _abc_15497_new_n5667_; 
wire _abc_15497_new_n5668_; 
wire _abc_15497_new_n5669_; 
wire _abc_15497_new_n5670_; 
wire _abc_15497_new_n5671_; 
wire _abc_15497_new_n5672_; 
wire _abc_15497_new_n5673_; 
wire _abc_15497_new_n5674_; 
wire _abc_15497_new_n5675_; 
wire _abc_15497_new_n5676_; 
wire _abc_15497_new_n5677_; 
wire _abc_15497_new_n5678_; 
wire _abc_15497_new_n5679_; 
wire _abc_15497_new_n5680_; 
wire _abc_15497_new_n5681_; 
wire _abc_15497_new_n5682_; 
wire _abc_15497_new_n5683_; 
wire _abc_15497_new_n5684_; 
wire _abc_15497_new_n5685_; 
wire _abc_15497_new_n5686_; 
wire _abc_15497_new_n5687_; 
wire _abc_15497_new_n5688_; 
wire _abc_15497_new_n5689_; 
wire _abc_15497_new_n5690_; 
wire _abc_15497_new_n5691_; 
wire _abc_15497_new_n5692_; 
wire _abc_15497_new_n5693_; 
wire _abc_15497_new_n5694_; 
wire _abc_15497_new_n5695_; 
wire _abc_15497_new_n5696_; 
wire _abc_15497_new_n5697_; 
wire _abc_15497_new_n5698_; 
wire _abc_15497_new_n5699_; 
wire _abc_15497_new_n5700_; 
wire _abc_15497_new_n5701_; 
wire _abc_15497_new_n5702_; 
wire _abc_15497_new_n5703_; 
wire _abc_15497_new_n5704_; 
wire _abc_15497_new_n5705_; 
wire _abc_15497_new_n5706_; 
wire _abc_15497_new_n5707_; 
wire _abc_15497_new_n5708_; 
wire _abc_15497_new_n5709_; 
wire _abc_15497_new_n5710_; 
wire _abc_15497_new_n5711_; 
wire _abc_15497_new_n5712_; 
wire _abc_15497_new_n5713_; 
wire _abc_15497_new_n5714_; 
wire _abc_15497_new_n5715_; 
wire _abc_15497_new_n5716_; 
wire _abc_15497_new_n5717_; 
wire _abc_15497_new_n5718_; 
wire _abc_15497_new_n5719_; 
wire _abc_15497_new_n5720_; 
wire _abc_15497_new_n5722_; 
wire _abc_15497_new_n5723_; 
wire _abc_15497_new_n5724_; 
wire _abc_15497_new_n5725_; 
wire _abc_15497_new_n5726_; 
wire _abc_15497_new_n5727_; 
wire _abc_15497_new_n5728_; 
wire _abc_15497_new_n5729_; 
wire _abc_15497_new_n5730_; 
wire _abc_15497_new_n5731_; 
wire _abc_15497_new_n5732_; 
wire _abc_15497_new_n5733_; 
wire _abc_15497_new_n5734_; 
wire _abc_15497_new_n5735_; 
wire _abc_15497_new_n5736_; 
wire _abc_15497_new_n5737_; 
wire _abc_15497_new_n5738_; 
wire _abc_15497_new_n5739_; 
wire _abc_15497_new_n5740_; 
wire _abc_15497_new_n5741_; 
wire _abc_15497_new_n5742_; 
wire _abc_15497_new_n5743_; 
wire _abc_15497_new_n5744_; 
wire _abc_15497_new_n5745_; 
wire _abc_15497_new_n5746_; 
wire _abc_15497_new_n5747_; 
wire _abc_15497_new_n5748_; 
wire _abc_15497_new_n5749_; 
wire _abc_15497_new_n5750_; 
wire _abc_15497_new_n5751_; 
wire _abc_15497_new_n5752_; 
wire _abc_15497_new_n5753_; 
wire _abc_15497_new_n5754_; 
wire _abc_15497_new_n5755_; 
wire _abc_15497_new_n5756_; 
wire _abc_15497_new_n5757_; 
wire _abc_15497_new_n5758_; 
wire _abc_15497_new_n5759_; 
wire _abc_15497_new_n5760_; 
wire _abc_15497_new_n5761_; 
wire _abc_15497_new_n5762_; 
wire _abc_15497_new_n5763_; 
wire _abc_15497_new_n5764_; 
wire _abc_15497_new_n5765_; 
wire _abc_15497_new_n5766_; 
wire _abc_15497_new_n5767_; 
wire _abc_15497_new_n5768_; 
wire _abc_15497_new_n5769_; 
wire _abc_15497_new_n5770_; 
wire _abc_15497_new_n5771_; 
wire _abc_15497_new_n5772_; 
wire _abc_15497_new_n5773_; 
wire _abc_15497_new_n5774_; 
wire _abc_15497_new_n5775_; 
wire _abc_15497_new_n5776_; 
wire _abc_15497_new_n5777_; 
wire _abc_15497_new_n5778_; 
wire _abc_15497_new_n5779_; 
wire _abc_15497_new_n5780_; 
wire _abc_15497_new_n5781_; 
wire _abc_15497_new_n5782_; 
wire _abc_15497_new_n5783_; 
wire _abc_15497_new_n5784_; 
wire _abc_15497_new_n5785_; 
wire _abc_15497_new_n5786_; 
wire _abc_15497_new_n5787_; 
wire _abc_15497_new_n5788_; 
wire _abc_15497_new_n5789_; 
wire _abc_15497_new_n5790_; 
wire _abc_15497_new_n5791_; 
wire _abc_15497_new_n5792_; 
wire _abc_15497_new_n5793_; 
wire _abc_15497_new_n5795_; 
wire _abc_15497_new_n5796_; 
wire _abc_15497_new_n5797_; 
wire _abc_15497_new_n5798_; 
wire _abc_15497_new_n5799_; 
wire _abc_15497_new_n5800_; 
wire _abc_15497_new_n5801_; 
wire _abc_15497_new_n5802_; 
wire _abc_15497_new_n5803_; 
wire _abc_15497_new_n5804_; 
wire _abc_15497_new_n5805_; 
wire _abc_15497_new_n5806_; 
wire _abc_15497_new_n5807_; 
wire _abc_15497_new_n5808_; 
wire _abc_15497_new_n5809_; 
wire _abc_15497_new_n5810_; 
wire _abc_15497_new_n5811_; 
wire _abc_15497_new_n5812_; 
wire _abc_15497_new_n5813_; 
wire _abc_15497_new_n5814_; 
wire _abc_15497_new_n5815_; 
wire _abc_15497_new_n5816_; 
wire _abc_15497_new_n5817_; 
wire _abc_15497_new_n5818_; 
wire _abc_15497_new_n5819_; 
wire _abc_15497_new_n5820_; 
wire _abc_15497_new_n5821_; 
wire _abc_15497_new_n5822_; 
wire _abc_15497_new_n5823_; 
wire _abc_15497_new_n5824_; 
wire _abc_15497_new_n5825_; 
wire _abc_15497_new_n5826_; 
wire _abc_15497_new_n5827_; 
wire _abc_15497_new_n5828_; 
wire _abc_15497_new_n5829_; 
wire _abc_15497_new_n5830_; 
wire _abc_15497_new_n5831_; 
wire _abc_15497_new_n5832_; 
wire _abc_15497_new_n5833_; 
wire _abc_15497_new_n5834_; 
wire _abc_15497_new_n5835_; 
wire _abc_15497_new_n5836_; 
wire _abc_15497_new_n5837_; 
wire _abc_15497_new_n5838_; 
wire _abc_15497_new_n5839_; 
wire _abc_15497_new_n5840_; 
wire _abc_15497_new_n5841_; 
wire _abc_15497_new_n5842_; 
wire _abc_15497_new_n5843_; 
wire _abc_15497_new_n5844_; 
wire _abc_15497_new_n5845_; 
wire _abc_15497_new_n5846_; 
wire _abc_15497_new_n5847_; 
wire _abc_15497_new_n5848_; 
wire _abc_15497_new_n5849_; 
wire _abc_15497_new_n5850_; 
wire _abc_15497_new_n5851_; 
wire _abc_15497_new_n5852_; 
wire _abc_15497_new_n5853_; 
wire _abc_15497_new_n5854_; 
wire _abc_15497_new_n5855_; 
wire _abc_15497_new_n5856_; 
wire _abc_15497_new_n5857_; 
wire _abc_15497_new_n5858_; 
wire _abc_15497_new_n5860_; 
wire _abc_15497_new_n5861_; 
wire _abc_15497_new_n5862_; 
wire _abc_15497_new_n5863_; 
wire _abc_15497_new_n5864_; 
wire _abc_15497_new_n5865_; 
wire _abc_15497_new_n5866_; 
wire _abc_15497_new_n5867_; 
wire _abc_15497_new_n5868_; 
wire _abc_15497_new_n5869_; 
wire _abc_15497_new_n5870_; 
wire _abc_15497_new_n5871_; 
wire _abc_15497_new_n5872_; 
wire _abc_15497_new_n5873_; 
wire _abc_15497_new_n5874_; 
wire _abc_15497_new_n5875_; 
wire _abc_15497_new_n5876_; 
wire _abc_15497_new_n5877_; 
wire _abc_15497_new_n5878_; 
wire _abc_15497_new_n5879_; 
wire _abc_15497_new_n5880_; 
wire _abc_15497_new_n5881_; 
wire _abc_15497_new_n5882_; 
wire _abc_15497_new_n5883_; 
wire _abc_15497_new_n5884_; 
wire _abc_15497_new_n5885_; 
wire _abc_15497_new_n5886_; 
wire _abc_15497_new_n5887_; 
wire _abc_15497_new_n5888_; 
wire _abc_15497_new_n5889_; 
wire _abc_15497_new_n5890_; 
wire _abc_15497_new_n5891_; 
wire _abc_15497_new_n5892_; 
wire _abc_15497_new_n5893_; 
wire _abc_15497_new_n5894_; 
wire _abc_15497_new_n5895_; 
wire _abc_15497_new_n5896_; 
wire _abc_15497_new_n5897_; 
wire _abc_15497_new_n5898_; 
wire _abc_15497_new_n5899_; 
wire _abc_15497_new_n5900_; 
wire _abc_15497_new_n5901_; 
wire _abc_15497_new_n5902_; 
wire _abc_15497_new_n5903_; 
wire _abc_15497_new_n5904_; 
wire _abc_15497_new_n5905_; 
wire _abc_15497_new_n5906_; 
wire _abc_15497_new_n5907_; 
wire _abc_15497_new_n5908_; 
wire _abc_15497_new_n5909_; 
wire _abc_15497_new_n5910_; 
wire _abc_15497_new_n5911_; 
wire _abc_15497_new_n5912_; 
wire _abc_15497_new_n5913_; 
wire _abc_15497_new_n5914_; 
wire _abc_15497_new_n5915_; 
wire _abc_15497_new_n5916_; 
wire _abc_15497_new_n5917_; 
wire _abc_15497_new_n5918_; 
wire _abc_15497_new_n5919_; 
wire _abc_15497_new_n5920_; 
wire _abc_15497_new_n5921_; 
wire _abc_15497_new_n5922_; 
wire _abc_15497_new_n5923_; 
wire _abc_15497_new_n5924_; 
wire _abc_15497_new_n5925_; 
wire _abc_15497_new_n5926_; 
wire _abc_15497_new_n5927_; 
wire _abc_15497_new_n5928_; 
wire _abc_15497_new_n5929_; 
wire _abc_15497_new_n5930_; 
wire _abc_15497_new_n5931_; 
wire _abc_15497_new_n5932_; 
wire _abc_15497_new_n5933_; 
wire _abc_15497_new_n5934_; 
wire _abc_15497_new_n5935_; 
wire _abc_15497_new_n5936_; 
wire _abc_15497_new_n5938_; 
wire _abc_15497_new_n5939_; 
wire _abc_15497_new_n5940_; 
wire _abc_15497_new_n5941_; 
wire _abc_15497_new_n5942_; 
wire _abc_15497_new_n5943_; 
wire _abc_15497_new_n5944_; 
wire _abc_15497_new_n5945_; 
wire _abc_15497_new_n5946_; 
wire _abc_15497_new_n5947_; 
wire _abc_15497_new_n5948_; 
wire _abc_15497_new_n5949_; 
wire _abc_15497_new_n5950_; 
wire _abc_15497_new_n5951_; 
wire _abc_15497_new_n5952_; 
wire _abc_15497_new_n5953_; 
wire _abc_15497_new_n5954_; 
wire _abc_15497_new_n5955_; 
wire _abc_15497_new_n5956_; 
wire _abc_15497_new_n5957_; 
wire _abc_15497_new_n5958_; 
wire _abc_15497_new_n5959_; 
wire _abc_15497_new_n5960_; 
wire _abc_15497_new_n5961_; 
wire _abc_15497_new_n5962_; 
wire _abc_15497_new_n5963_; 
wire _abc_15497_new_n5964_; 
wire _abc_15497_new_n5965_; 
wire _abc_15497_new_n5966_; 
wire _abc_15497_new_n5967_; 
wire _abc_15497_new_n5968_; 
wire _abc_15497_new_n5969_; 
wire _abc_15497_new_n5970_; 
wire _abc_15497_new_n5971_; 
wire _abc_15497_new_n5972_; 
wire _abc_15497_new_n5973_; 
wire _abc_15497_new_n5974_; 
wire _abc_15497_new_n5975_; 
wire _abc_15497_new_n5976_; 
wire _abc_15497_new_n5977_; 
wire _abc_15497_new_n5978_; 
wire _abc_15497_new_n5979_; 
wire _abc_15497_new_n5980_; 
wire _abc_15497_new_n5981_; 
wire _abc_15497_new_n5982_; 
wire _abc_15497_new_n5983_; 
wire _abc_15497_new_n5984_; 
wire _abc_15497_new_n5985_; 
wire _abc_15497_new_n5986_; 
wire _abc_15497_new_n5987_; 
wire _abc_15497_new_n5988_; 
wire _abc_15497_new_n5989_; 
wire _abc_15497_new_n5990_; 
wire _abc_15497_new_n5991_; 
wire _abc_15497_new_n5992_; 
wire _abc_15497_new_n5993_; 
wire _abc_15497_new_n5994_; 
wire _abc_15497_new_n5995_; 
wire _abc_15497_new_n5996_; 
wire _abc_15497_new_n5997_; 
wire _abc_15497_new_n5998_; 
wire _abc_15497_new_n5999_; 
wire _abc_15497_new_n6000_; 
wire _abc_15497_new_n6001_; 
wire _abc_15497_new_n6002_; 
wire _abc_15497_new_n6003_; 
wire _abc_15497_new_n6004_; 
wire _abc_15497_new_n6005_; 
wire _abc_15497_new_n6007_; 
wire _abc_15497_new_n6008_; 
wire _abc_15497_new_n6009_; 
wire _abc_15497_new_n6010_; 
wire _abc_15497_new_n6011_; 
wire _abc_15497_new_n6012_; 
wire _abc_15497_new_n6013_; 
wire _abc_15497_new_n6014_; 
wire _abc_15497_new_n6015_; 
wire _abc_15497_new_n6016_; 
wire _abc_15497_new_n6017_; 
wire _abc_15497_new_n6018_; 
wire _abc_15497_new_n6019_; 
wire _abc_15497_new_n6020_; 
wire _abc_15497_new_n6021_; 
wire _abc_15497_new_n6022_; 
wire _abc_15497_new_n6023_; 
wire _abc_15497_new_n6024_; 
wire _abc_15497_new_n6025_; 
wire _abc_15497_new_n6026_; 
wire _abc_15497_new_n6027_; 
wire _abc_15497_new_n6028_; 
wire _abc_15497_new_n6029_; 
wire _abc_15497_new_n6030_; 
wire _abc_15497_new_n6031_; 
wire _abc_15497_new_n6032_; 
wire _abc_15497_new_n6033_; 
wire _abc_15497_new_n6034_; 
wire _abc_15497_new_n6035_; 
wire _abc_15497_new_n6036_; 
wire _abc_15497_new_n6037_; 
wire _abc_15497_new_n6038_; 
wire _abc_15497_new_n6039_; 
wire _abc_15497_new_n6040_; 
wire _abc_15497_new_n6041_; 
wire _abc_15497_new_n6042_; 
wire _abc_15497_new_n6043_; 
wire _abc_15497_new_n6044_; 
wire _abc_15497_new_n6045_; 
wire _abc_15497_new_n6046_; 
wire _abc_15497_new_n6047_; 
wire _abc_15497_new_n6048_; 
wire _abc_15497_new_n6049_; 
wire _abc_15497_new_n6050_; 
wire _abc_15497_new_n6051_; 
wire _abc_15497_new_n6052_; 
wire _abc_15497_new_n6053_; 
wire _abc_15497_new_n6054_; 
wire _abc_15497_new_n6055_; 
wire _abc_15497_new_n6056_; 
wire _abc_15497_new_n6057_; 
wire _abc_15497_new_n6058_; 
wire _abc_15497_new_n6059_; 
wire _abc_15497_new_n6060_; 
wire _abc_15497_new_n6061_; 
wire _abc_15497_new_n6062_; 
wire _abc_15497_new_n6063_; 
wire _abc_15497_new_n6064_; 
wire _abc_15497_new_n6065_; 
wire _abc_15497_new_n6066_; 
wire _abc_15497_new_n6067_; 
wire _abc_15497_new_n6068_; 
wire _abc_15497_new_n6069_; 
wire _abc_15497_new_n6070_; 
wire _abc_15497_new_n6071_; 
wire _abc_15497_new_n6072_; 
wire _abc_15497_new_n6073_; 
wire _abc_15497_new_n6074_; 
wire _abc_15497_new_n6075_; 
wire _abc_15497_new_n6076_; 
wire _abc_15497_new_n6077_; 
wire _abc_15497_new_n6078_; 
wire _abc_15497_new_n6079_; 
wire _abc_15497_new_n6081_; 
wire _abc_15497_new_n6082_; 
wire _abc_15497_new_n6083_; 
wire _abc_15497_new_n6084_; 
wire _abc_15497_new_n6085_; 
wire _abc_15497_new_n6086_; 
wire _abc_15497_new_n6087_; 
wire _abc_15497_new_n6088_; 
wire _abc_15497_new_n6089_; 
wire _abc_15497_new_n6090_; 
wire _abc_15497_new_n6091_; 
wire _abc_15497_new_n6092_; 
wire _abc_15497_new_n6093_; 
wire _abc_15497_new_n6094_; 
wire _abc_15497_new_n6095_; 
wire _abc_15497_new_n6096_; 
wire _abc_15497_new_n6097_; 
wire _abc_15497_new_n6098_; 
wire _abc_15497_new_n6099_; 
wire _abc_15497_new_n6100_; 
wire _abc_15497_new_n6101_; 
wire _abc_15497_new_n6102_; 
wire _abc_15497_new_n6103_; 
wire _abc_15497_new_n6104_; 
wire _abc_15497_new_n6105_; 
wire _abc_15497_new_n6106_; 
wire _abc_15497_new_n6107_; 
wire _abc_15497_new_n6108_; 
wire _abc_15497_new_n6109_; 
wire _abc_15497_new_n6110_; 
wire _abc_15497_new_n6111_; 
wire _abc_15497_new_n6112_; 
wire _abc_15497_new_n6113_; 
wire _abc_15497_new_n6114_; 
wire _abc_15497_new_n6115_; 
wire _abc_15497_new_n6116_; 
wire _abc_15497_new_n6117_; 
wire _abc_15497_new_n6118_; 
wire _abc_15497_new_n6119_; 
wire _abc_15497_new_n6120_; 
wire _abc_15497_new_n6121_; 
wire _abc_15497_new_n6122_; 
wire _abc_15497_new_n6123_; 
wire _abc_15497_new_n6124_; 
wire _abc_15497_new_n6125_; 
wire _abc_15497_new_n6126_; 
wire _abc_15497_new_n6127_; 
wire _abc_15497_new_n6128_; 
wire _abc_15497_new_n6129_; 
wire _abc_15497_new_n6130_; 
wire _abc_15497_new_n6131_; 
wire _abc_15497_new_n6132_; 
wire _abc_15497_new_n6133_; 
wire _abc_15497_new_n6134_; 
wire _abc_15497_new_n6135_; 
wire _abc_15497_new_n6136_; 
wire _abc_15497_new_n6137_; 
wire _abc_15497_new_n6138_; 
wire _abc_15497_new_n6139_; 
wire _abc_15497_new_n6140_; 
wire _abc_15497_new_n6141_; 
wire _abc_15497_new_n6142_; 
wire _abc_15497_new_n6143_; 
wire _abc_15497_new_n6144_; 
wire _abc_15497_new_n6145_; 
wire _abc_15497_new_n6146_; 
wire _abc_15497_new_n6148_; 
wire _abc_15497_new_n6149_; 
wire _abc_15497_new_n6150_; 
wire _abc_15497_new_n6151_; 
wire _abc_15497_new_n6153_; 
wire _abc_15497_new_n6154_; 
wire _abc_15497_new_n6155_; 
wire _abc_15497_new_n6156_; 
wire _abc_15497_new_n6157_; 
wire _abc_15497_new_n6159_; 
wire _abc_15497_new_n6161_; 
wire _abc_15497_new_n6162_; 
wire _abc_15497_new_n6163_; 
wire _abc_15497_new_n6165_; 
wire _abc_15497_new_n6166_; 
wire _abc_15497_new_n6167_; 
wire _abc_15497_new_n6168_; 
wire _abc_15497_new_n6169_; 
wire _abc_15497_new_n6171_; 
wire _abc_15497_new_n6172_; 
wire _abc_15497_new_n6173_; 
wire _abc_15497_new_n6174_; 
wire _abc_15497_new_n6175_; 
wire _abc_15497_new_n6176_; 
wire _abc_15497_new_n6178_; 
wire _abc_15497_new_n6179_; 
wire _abc_15497_new_n6180_; 
wire _abc_15497_new_n6181_; 
wire _abc_15497_new_n6182_; 
wire _abc_15497_new_n6183_; 
wire _abc_15497_new_n6185_; 
wire _abc_15497_new_n6186_; 
wire _abc_15497_new_n6187_; 
wire _abc_15497_new_n6188_; 
wire _abc_15497_new_n6190_; 
wire _abc_15497_new_n6191_; 
wire _abc_15497_new_n6192_; 
wire _abc_15497_new_n6193_; 
wire _abc_15497_new_n6194_; 
wire _abc_15497_new_n6196_; 
wire _abc_15497_new_n6197_; 
wire _abc_15497_new_n6198_; 
wire _abc_15497_new_n6200_; 
wire _abc_15497_new_n6202_; 
wire _abc_15497_new_n6203_; 
wire _abc_15497_new_n6204_; 
wire _abc_15497_new_n6205_; 
wire _abc_15497_new_n6207_; 
wire _abc_15497_new_n6208_; 
wire _abc_15497_new_n6209_; 
wire _abc_15497_new_n6210_; 
wire _abc_15497_new_n6212_; 
wire _abc_15497_new_n6213_; 
wire _abc_15497_new_n6214_; 
wire _abc_15497_new_n6215_; 
wire _abc_15497_new_n6217_; 
wire _abc_15497_new_n6218_; 
wire _abc_15497_new_n6219_; 
wire _abc_15497_new_n6220_; 
wire _abc_15497_new_n6221_; 
wire _abc_15497_new_n6222_; 
wire _abc_15497_new_n6223_; 
wire _abc_15497_new_n6225_; 
wire _abc_15497_new_n6226_; 
wire _abc_15497_new_n6227_; 
wire _abc_15497_new_n6228_; 
wire _abc_15497_new_n6230_; 
wire _abc_15497_new_n6231_; 
wire _abc_15497_new_n6232_; 
wire _abc_15497_new_n6233_; 
wire _abc_15497_new_n6234_; 
wire _abc_15497_new_n6235_; 
wire _abc_15497_new_n6236_; 
wire _abc_15497_new_n6238_; 
wire _abc_15497_new_n6239_; 
wire _abc_15497_new_n6240_; 
wire _abc_15497_new_n6241_; 
wire _abc_15497_new_n6242_; 
wire _abc_15497_new_n6243_; 
wire _abc_15497_new_n6245_; 
wire _abc_15497_new_n6246_; 
wire _abc_15497_new_n6247_; 
wire _abc_15497_new_n6248_; 
wire _abc_15497_new_n6249_; 
wire _abc_15497_new_n6250_; 
wire _abc_15497_new_n6251_; 
wire _abc_15497_new_n6252_; 
wire _abc_15497_new_n6254_; 
wire _abc_15497_new_n6255_; 
wire _abc_15497_new_n6256_; 
wire _abc_15497_new_n6257_; 
wire _abc_15497_new_n6258_; 
wire _abc_15497_new_n6259_; 
wire _abc_15497_new_n6261_; 
wire _abc_15497_new_n6262_; 
wire _abc_15497_new_n6263_; 
wire _abc_15497_new_n6264_; 
wire _abc_15497_new_n6265_; 
wire _abc_15497_new_n6266_; 
wire _abc_15497_new_n6267_; 
wire _abc_15497_new_n6268_; 
wire _abc_15497_new_n6270_; 
wire _abc_15497_new_n6271_; 
wire _abc_15497_new_n6272_; 
wire _abc_15497_new_n6273_; 
wire _abc_15497_new_n6274_; 
wire _abc_15497_new_n6275_; 
wire _abc_15497_new_n6277_; 
wire _abc_15497_new_n6278_; 
wire _abc_15497_new_n6279_; 
wire _abc_15497_new_n6280_; 
wire _abc_15497_new_n6281_; 
wire _abc_15497_new_n6282_; 
wire _abc_15497_new_n6283_; 
wire _abc_15497_new_n6284_; 
wire _abc_15497_new_n6286_; 
wire _abc_15497_new_n6287_; 
wire _abc_15497_new_n6288_; 
wire _abc_15497_new_n6289_; 
wire _abc_15497_new_n6290_; 
wire _abc_15497_new_n6291_; 
wire _abc_15497_new_n6293_; 
wire _abc_15497_new_n6294_; 
wire _abc_15497_new_n6295_; 
wire _abc_15497_new_n6296_; 
wire _abc_15497_new_n6297_; 
wire _abc_15497_new_n6298_; 
wire _abc_15497_new_n6299_; 
wire _abc_15497_new_n6301_; 
wire _abc_15497_new_n6302_; 
wire _abc_15497_new_n6303_; 
wire _abc_15497_new_n6304_; 
wire _abc_15497_new_n6305_; 
wire _abc_15497_new_n6306_; 
wire _abc_15497_new_n6307_; 
wire _abc_15497_new_n6308_; 
wire _abc_15497_new_n6310_; 
wire _abc_15497_new_n6311_; 
wire _abc_15497_new_n6312_; 
wire _abc_15497_new_n6313_; 
wire _abc_15497_new_n6314_; 
wire _abc_15497_new_n6315_; 
wire _abc_15497_new_n6316_; 
wire _abc_15497_new_n6317_; 
wire _abc_15497_new_n6319_; 
wire _abc_15497_new_n6320_; 
wire _abc_15497_new_n6321_; 
wire _abc_15497_new_n6322_; 
wire _abc_15497_new_n6323_; 
wire _abc_15497_new_n6324_; 
wire _abc_15497_new_n6326_; 
wire _abc_15497_new_n6327_; 
wire _abc_15497_new_n6328_; 
wire _abc_15497_new_n6329_; 
wire _abc_15497_new_n6330_; 
wire _abc_15497_new_n6331_; 
wire _abc_15497_new_n6332_; 
wire _abc_15497_new_n6334_; 
wire _abc_15497_new_n6335_; 
wire _abc_15497_new_n6336_; 
wire _abc_15497_new_n6337_; 
wire _abc_15497_new_n6338_; 
wire _abc_15497_new_n6339_; 
wire _abc_15497_new_n6340_; 
wire _abc_15497_new_n6341_; 
wire _abc_15497_new_n6343_; 
wire _abc_15497_new_n6344_; 
wire _abc_15497_new_n6345_; 
wire _abc_15497_new_n6346_; 
wire _abc_15497_new_n6347_; 
wire _abc_15497_new_n6348_; 
wire _abc_15497_new_n6349_; 
wire _abc_15497_new_n6350_; 
wire _abc_15497_new_n6352_; 
wire _abc_15497_new_n6353_; 
wire _abc_15497_new_n6354_; 
wire _abc_15497_new_n6355_; 
wire _abc_15497_new_n6356_; 
wire _abc_15497_new_n6357_; 
wire _abc_15497_new_n6358_; 
wire _abc_15497_new_n6359_; 
wire _abc_15497_new_n6361_; 
wire _abc_15497_new_n6362_; 
wire _abc_15497_new_n6363_; 
wire _abc_15497_new_n6364_; 
wire _abc_15497_new_n6365_; 
wire _abc_15497_new_n6366_; 
wire _abc_15497_new_n6367_; 
wire _abc_15497_new_n6369_; 
wire _abc_15497_new_n6370_; 
wire _abc_15497_new_n6371_; 
wire _abc_15497_new_n6372_; 
wire _abc_15497_new_n6373_; 
wire _abc_15497_new_n6374_; 
wire _abc_15497_new_n6375_; 
wire _abc_15497_new_n6376_; 
wire _abc_15497_new_n6378_; 
wire _abc_15497_new_n6379_; 
wire _abc_15497_new_n6380_; 
wire _abc_15497_new_n6381_; 
wire _abc_15497_new_n6382_; 
wire _abc_15497_new_n6383_; 
wire _abc_15497_new_n6384_; 
wire _abc_15497_new_n6385_; 
wire _abc_15497_new_n6387_; 
wire _abc_15497_new_n6388_; 
wire _abc_15497_new_n6389_; 
wire _abc_15497_new_n6390_; 
wire _abc_15497_new_n6391_; 
wire _abc_15497_new_n6392_; 
wire _abc_15497_new_n6394_; 
wire _abc_15497_new_n6395_; 
wire _abc_15497_new_n6396_; 
wire _abc_15497_new_n6397_; 
wire _abc_15497_new_n6398_; 
wire _abc_15497_new_n6399_; 
wire _abc_15497_new_n6400_; 
wire _abc_15497_new_n6401_; 
wire _abc_15497_new_n698_; 
wire _abc_15497_new_n699_; 
wire _abc_15497_new_n700_; 
wire _abc_15497_new_n701_; 
wire _abc_15497_new_n702_; 
wire _abc_15497_new_n703_; 
wire _abc_15497_new_n704_; 
wire _abc_15497_new_n705_; 
wire _abc_15497_new_n706_; 
wire _abc_15497_new_n707_; 
wire _abc_15497_new_n708_; 
wire _abc_15497_new_n709_; 
wire _abc_15497_new_n710_; 
wire _abc_15497_new_n711_; 
wire _abc_15497_new_n712_; 
wire _abc_15497_new_n713_; 
wire _abc_15497_new_n714_; 
wire _abc_15497_new_n715_; 
wire _abc_15497_new_n716_; 
wire _abc_15497_new_n717_; 
wire _abc_15497_new_n718_; 
wire _abc_15497_new_n719_; 
wire _abc_15497_new_n720_; 
wire _abc_15497_new_n721_; 
wire _abc_15497_new_n722_; 
wire _abc_15497_new_n723_; 
wire _abc_15497_new_n724_; 
wire _abc_15497_new_n725_; 
wire _abc_15497_new_n726_; 
wire _abc_15497_new_n727_; 
wire _abc_15497_new_n728_; 
wire _abc_15497_new_n729_; 
wire _abc_15497_new_n730_; 
wire _abc_15497_new_n731_; 
wire _abc_15497_new_n732_; 
wire _abc_15497_new_n733_; 
wire _abc_15497_new_n734_; 
wire _abc_15497_new_n735_; 
wire _abc_15497_new_n736_; 
wire _abc_15497_new_n737_; 
wire _abc_15497_new_n738_; 
wire _abc_15497_new_n739_; 
wire _abc_15497_new_n740_; 
wire _abc_15497_new_n741_; 
wire _abc_15497_new_n742_; 
wire _abc_15497_new_n743_; 
wire _abc_15497_new_n744_; 
wire _abc_15497_new_n745_; 
wire _abc_15497_new_n746_; 
wire _abc_15497_new_n747_; 
wire _abc_15497_new_n748_; 
wire _abc_15497_new_n749_; 
wire _abc_15497_new_n750_; 
wire _abc_15497_new_n751_; 
wire _abc_15497_new_n752_; 
wire _abc_15497_new_n753_; 
wire _abc_15497_new_n754_; 
wire _abc_15497_new_n755_; 
wire _abc_15497_new_n756_; 
wire _abc_15497_new_n757_; 
wire _abc_15497_new_n758_; 
wire _abc_15497_new_n759_; 
wire _abc_15497_new_n760_; 
wire _abc_15497_new_n761_; 
wire _abc_15497_new_n762_; 
wire _abc_15497_new_n763_; 
wire _abc_15497_new_n764_; 
wire _abc_15497_new_n765_; 
wire _abc_15497_new_n766_; 
wire _abc_15497_new_n767_; 
wire _abc_15497_new_n768_; 
wire _abc_15497_new_n769_; 
wire _abc_15497_new_n770_; 
wire _abc_15497_new_n771_; 
wire _abc_15497_new_n772_; 
wire _abc_15497_new_n773_; 
wire _abc_15497_new_n774_; 
wire _abc_15497_new_n775_; 
wire _abc_15497_new_n776_; 
wire _abc_15497_new_n777_; 
wire _abc_15497_new_n778_; 
wire _abc_15497_new_n779_; 
wire _abc_15497_new_n780_; 
wire _abc_15497_new_n781_; 
wire _abc_15497_new_n782_; 
wire _abc_15497_new_n783_; 
wire _abc_15497_new_n784_; 
wire _abc_15497_new_n785_; 
wire _abc_15497_new_n786_; 
wire _abc_15497_new_n787_; 
wire _abc_15497_new_n788_; 
wire _abc_15497_new_n789_; 
wire _abc_15497_new_n790_; 
wire _abc_15497_new_n791_; 
wire _abc_15497_new_n792_; 
wire _abc_15497_new_n793_; 
wire _abc_15497_new_n794_; 
wire _abc_15497_new_n795_; 
wire _abc_15497_new_n796_; 
wire _abc_15497_new_n797_; 
wire _abc_15497_new_n798_; 
wire _abc_15497_new_n799_; 
wire _abc_15497_new_n800_; 
wire _abc_15497_new_n801_; 
wire _abc_15497_new_n802_; 
wire _abc_15497_new_n803_; 
wire _abc_15497_new_n804_; 
wire _abc_15497_new_n805_; 
wire _abc_15497_new_n806_; 
wire _abc_15497_new_n807_; 
wire _abc_15497_new_n808_; 
wire _abc_15497_new_n809_; 
wire _abc_15497_new_n810_; 
wire _abc_15497_new_n811_; 
wire _abc_15497_new_n812_; 
wire _abc_15497_new_n813_; 
wire _abc_15497_new_n814_; 
wire _abc_15497_new_n815_; 
wire _abc_15497_new_n816_; 
wire _abc_15497_new_n817_; 
wire _abc_15497_new_n818_; 
wire _abc_15497_new_n819_; 
wire _abc_15497_new_n820_; 
wire _abc_15497_new_n821_; 
wire _abc_15497_new_n822_; 
wire _abc_15497_new_n823_; 
wire _abc_15497_new_n824_; 
wire _abc_15497_new_n825_; 
wire _abc_15497_new_n826_; 
wire _abc_15497_new_n827_; 
wire _abc_15497_new_n828_; 
wire _abc_15497_new_n829_; 
wire _abc_15497_new_n830_; 
wire _abc_15497_new_n831_; 
wire _abc_15497_new_n832_; 
wire _abc_15497_new_n833_; 
wire _abc_15497_new_n834_; 
wire _abc_15497_new_n835_; 
wire _abc_15497_new_n836_; 
wire _abc_15497_new_n837_; 
wire _abc_15497_new_n838_; 
wire _abc_15497_new_n839_; 
wire _abc_15497_new_n840_; 
wire _abc_15497_new_n841_; 
wire _abc_15497_new_n842_; 
wire _abc_15497_new_n843_; 
wire _abc_15497_new_n844_; 
wire _abc_15497_new_n845_; 
wire _abc_15497_new_n846_; 
wire _abc_15497_new_n847_; 
wire _abc_15497_new_n848_; 
wire _abc_15497_new_n849_; 
wire _abc_15497_new_n850_; 
wire _abc_15497_new_n851_; 
wire _abc_15497_new_n852_; 
wire _abc_15497_new_n853_; 
wire _abc_15497_new_n854_; 
wire _abc_15497_new_n855_; 
wire _abc_15497_new_n856_; 
wire _abc_15497_new_n857_; 
wire _abc_15497_new_n858_; 
wire _abc_15497_new_n859_; 
wire _abc_15497_new_n860_; 
wire _abc_15497_new_n861_; 
wire _abc_15497_new_n862_; 
wire _abc_15497_new_n863_; 
wire _abc_15497_new_n864_; 
wire _abc_15497_new_n865_; 
wire _abc_15497_new_n866_; 
wire _abc_15497_new_n867_; 
wire _abc_15497_new_n868_; 
wire _abc_15497_new_n869_; 
wire _abc_15497_new_n870_; 
wire _abc_15497_new_n871_; 
wire _abc_15497_new_n872_; 
wire _abc_15497_new_n873_; 
wire _abc_15497_new_n874_; 
wire _abc_15497_new_n875_; 
wire _abc_15497_new_n876_; 
wire _abc_15497_new_n877_; 
wire _abc_15497_new_n878_; 
wire _abc_15497_new_n879_; 
wire _abc_15497_new_n880_; 
wire _abc_15497_new_n881_; 
wire _abc_15497_new_n883_; 
wire _abc_15497_new_n884_; 
wire _abc_15497_new_n885_; 
wire _abc_15497_new_n886_; 
wire _abc_15497_new_n887_; 
wire _abc_15497_new_n888_; 
wire _abc_15497_new_n889_; 
wire _abc_15497_new_n890_; 
wire _abc_15497_new_n891_; 
wire _abc_15497_new_n892_; 
wire _abc_15497_new_n893_; 
wire _abc_15497_new_n894_; 
wire _abc_15497_new_n895_; 
wire _abc_15497_new_n897_; 
wire _abc_15497_new_n898_; 
wire _abc_15497_new_n899_; 
wire _abc_15497_new_n900_; 
wire _abc_15497_new_n901_; 
wire _abc_15497_new_n902_; 
wire _abc_15497_new_n903_; 
wire _abc_15497_new_n904_; 
wire _abc_15497_new_n905_; 
wire _abc_15497_new_n906_; 
wire _abc_15497_new_n907_; 
wire _abc_15497_new_n908_; 
wire _abc_15497_new_n909_; 
wire _abc_15497_new_n910_; 
wire _abc_15497_new_n911_; 
wire _abc_15497_new_n912_; 
wire _abc_15497_new_n914_; 
wire _abc_15497_new_n915_; 
wire _abc_15497_new_n916_; 
wire _abc_15497_new_n917_; 
wire _abc_15497_new_n918_; 
wire _abc_15497_new_n919_; 
wire _abc_15497_new_n920_; 
wire _abc_15497_new_n921_; 
wire _abc_15497_new_n922_; 
wire _abc_15497_new_n923_; 
wire _abc_15497_new_n924_; 
wire _abc_15497_new_n925_; 
wire _abc_15497_new_n927_; 
wire _abc_15497_new_n928_; 
wire _abc_15497_new_n929_; 
wire _abc_15497_new_n930_; 
wire _abc_15497_new_n931_; 
wire _abc_15497_new_n932_; 
wire _abc_15497_new_n933_; 
wire _abc_15497_new_n934_; 
wire _abc_15497_new_n935_; 
wire _abc_15497_new_n936_; 
wire _abc_15497_new_n937_; 
wire _abc_15497_new_n938_; 
wire _abc_15497_new_n939_; 
wire _abc_15497_new_n940_; 
wire _abc_15497_new_n941_; 
wire _abc_15497_new_n942_; 
wire _abc_15497_new_n943_; 
wire _abc_15497_new_n944_; 
wire _abc_15497_new_n945_; 
wire _abc_15497_new_n946_; 
wire _abc_15497_new_n947_; 
wire _abc_15497_new_n948_; 
wire _abc_15497_new_n949_; 
wire _abc_15497_new_n950_; 
wire _abc_15497_new_n951_; 
wire _abc_15497_new_n952_; 
wire _abc_15497_new_n953_; 
wire _abc_15497_new_n954_; 
wire _abc_15497_new_n955_; 
wire _abc_15497_new_n956_; 
wire _abc_15497_new_n957_; 
wire _abc_15497_new_n958_; 
wire _abc_15497_new_n959_; 
wire _abc_15497_new_n960_; 
wire _abc_15497_new_n961_; 
wire _abc_15497_new_n962_; 
wire _abc_15497_new_n963_; 
wire _abc_15497_new_n964_; 
wire _abc_15497_new_n965_; 
wire _abc_15497_new_n966_; 
wire _abc_15497_new_n967_; 
wire _abc_15497_new_n968_; 
wire _abc_15497_new_n969_; 
wire _abc_15497_new_n970_; 
wire _abc_15497_new_n971_; 
wire _abc_15497_new_n972_; 
wire _abc_15497_new_n973_; 
wire _abc_15497_new_n974_; 
wire _abc_15497_new_n975_; 
wire _abc_15497_new_n976_; 
wire _abc_15497_new_n977_; 
wire _abc_15497_new_n978_; 
wire _abc_15497_new_n979_; 
wire _abc_15497_new_n980_; 
wire _abc_15497_new_n981_; 
wire _abc_15497_new_n982_; 
wire _abc_15497_new_n983_; 
wire _abc_15497_new_n984_; 
wire _abc_15497_new_n985_; 
wire _abc_15497_new_n986_; 
wire _abc_15497_new_n987_; 
wire _abc_15497_new_n988_; 
wire _abc_15497_new_n989_; 
wire _abc_15497_new_n990_; 
wire _abc_15497_new_n991_; 
wire _abc_15497_new_n993_; 
wire _abc_15497_new_n994_; 
wire _abc_15497_new_n995_; 
wire _abc_15497_new_n996_; 
wire _abc_15497_new_n997_; 
wire _abc_15497_new_n998_; 
wire _abc_15497_new_n999_; 
wire a_reg_0_; 
wire a_reg_10_; 
wire a_reg_11_; 
wire a_reg_12_; 
wire a_reg_13_; 
wire a_reg_14_; 
wire a_reg_15_; 
wire a_reg_16_; 
wire a_reg_17_; 
wire a_reg_18_; 
wire a_reg_19_; 
wire a_reg_1_; 
wire a_reg_20_; 
wire a_reg_21_; 
wire a_reg_22_; 
wire a_reg_23_; 
wire a_reg_24_; 
wire a_reg_25_; 
wire a_reg_26_; 
wire a_reg_27_; 
wire a_reg_28_; 
wire a_reg_29_; 
wire a_reg_2_; 
wire a_reg_30_; 
wire a_reg_31_; 
wire a_reg_3_; 
wire a_reg_4_; 
wire a_reg_5_; 
wire a_reg_6_; 
wire a_reg_7_; 
wire a_reg_8_; 
wire a_reg_9_; 
wire b_reg_0_; 
wire b_reg_10_; 
wire b_reg_11_; 
wire b_reg_12_; 
wire b_reg_13_; 
wire b_reg_14_; 
wire b_reg_15_; 
wire b_reg_16_; 
wire b_reg_17_; 
wire b_reg_18_; 
wire b_reg_19_; 
wire b_reg_1_; 
wire b_reg_20_; 
wire b_reg_21_; 
wire b_reg_22_; 
wire b_reg_23_; 
wire b_reg_24_; 
wire b_reg_25_; 
wire b_reg_26_; 
wire b_reg_27_; 
wire b_reg_28_; 
wire b_reg_29_; 
wire b_reg_2_; 
wire b_reg_30_; 
wire b_reg_31_; 
wire b_reg_3_; 
wire b_reg_4_; 
wire b_reg_5_; 
wire b_reg_6_; 
wire b_reg_7_; 
wire b_reg_8_; 
wire b_reg_9_; 
input \block[0] ;
input \block[100] ;
input \block[101] ;
input \block[102] ;
input \block[103] ;
input \block[104] ;
input \block[105] ;
input \block[106] ;
input \block[107] ;
input \block[108] ;
input \block[109] ;
input \block[10] ;
input \block[110] ;
input \block[111] ;
input \block[112] ;
input \block[113] ;
input \block[114] ;
input \block[115] ;
input \block[116] ;
input \block[117] ;
input \block[118] ;
input \block[119] ;
input \block[11] ;
input \block[120] ;
input \block[121] ;
input \block[122] ;
input \block[123] ;
input \block[124] ;
input \block[125] ;
input \block[126] ;
input \block[127] ;
input \block[128] ;
input \block[129] ;
input \block[12] ;
input \block[130] ;
input \block[131] ;
input \block[132] ;
input \block[133] ;
input \block[134] ;
input \block[135] ;
input \block[136] ;
input \block[137] ;
input \block[138] ;
input \block[139] ;
input \block[13] ;
input \block[140] ;
input \block[141] ;
input \block[142] ;
input \block[143] ;
input \block[144] ;
input \block[145] ;
input \block[146] ;
input \block[147] ;
input \block[148] ;
input \block[149] ;
input \block[14] ;
input \block[150] ;
input \block[151] ;
input \block[152] ;
input \block[153] ;
input \block[154] ;
input \block[155] ;
input \block[156] ;
input \block[157] ;
input \block[158] ;
input \block[159] ;
input \block[15] ;
input \block[160] ;
input \block[161] ;
input \block[162] ;
input \block[163] ;
input \block[164] ;
input \block[165] ;
input \block[166] ;
input \block[167] ;
input \block[168] ;
input \block[169] ;
input \block[16] ;
input \block[170] ;
input \block[171] ;
input \block[172] ;
input \block[173] ;
input \block[174] ;
input \block[175] ;
input \block[176] ;
input \block[177] ;
input \block[178] ;
input \block[179] ;
input \block[17] ;
input \block[180] ;
input \block[181] ;
input \block[182] ;
input \block[183] ;
input \block[184] ;
input \block[185] ;
input \block[186] ;
input \block[187] ;
input \block[188] ;
input \block[189] ;
input \block[18] ;
input \block[190] ;
input \block[191] ;
input \block[192] ;
input \block[193] ;
input \block[194] ;
input \block[195] ;
input \block[196] ;
input \block[197] ;
input \block[198] ;
input \block[199] ;
input \block[19] ;
input \block[1] ;
input \block[200] ;
input \block[201] ;
input \block[202] ;
input \block[203] ;
input \block[204] ;
input \block[205] ;
input \block[206] ;
input \block[207] ;
input \block[208] ;
input \block[209] ;
input \block[20] ;
input \block[210] ;
input \block[211] ;
input \block[212] ;
input \block[213] ;
input \block[214] ;
input \block[215] ;
input \block[216] ;
input \block[217] ;
input \block[218] ;
input \block[219] ;
input \block[21] ;
input \block[220] ;
input \block[221] ;
input \block[222] ;
input \block[223] ;
input \block[224] ;
input \block[225] ;
input \block[226] ;
input \block[227] ;
input \block[228] ;
input \block[229] ;
input \block[22] ;
input \block[230] ;
input \block[231] ;
input \block[232] ;
input \block[233] ;
input \block[234] ;
input \block[235] ;
input \block[236] ;
input \block[237] ;
input \block[238] ;
input \block[239] ;
input \block[23] ;
input \block[240] ;
input \block[241] ;
input \block[242] ;
input \block[243] ;
input \block[244] ;
input \block[245] ;
input \block[246] ;
input \block[247] ;
input \block[248] ;
input \block[249] ;
input \block[24] ;
input \block[250] ;
input \block[251] ;
input \block[252] ;
input \block[253] ;
input \block[254] ;
input \block[255] ;
input \block[256] ;
input \block[257] ;
input \block[258] ;
input \block[259] ;
input \block[25] ;
input \block[260] ;
input \block[261] ;
input \block[262] ;
input \block[263] ;
input \block[264] ;
input \block[265] ;
input \block[266] ;
input \block[267] ;
input \block[268] ;
input \block[269] ;
input \block[26] ;
input \block[270] ;
input \block[271] ;
input \block[272] ;
input \block[273] ;
input \block[274] ;
input \block[275] ;
input \block[276] ;
input \block[277] ;
input \block[278] ;
input \block[279] ;
input \block[27] ;
input \block[280] ;
input \block[281] ;
input \block[282] ;
input \block[283] ;
input \block[284] ;
input \block[285] ;
input \block[286] ;
input \block[287] ;
input \block[288] ;
input \block[289] ;
input \block[28] ;
input \block[290] ;
input \block[291] ;
input \block[292] ;
input \block[293] ;
input \block[294] ;
input \block[295] ;
input \block[296] ;
input \block[297] ;
input \block[298] ;
input \block[299] ;
input \block[29] ;
input \block[2] ;
input \block[300] ;
input \block[301] ;
input \block[302] ;
input \block[303] ;
input \block[304] ;
input \block[305] ;
input \block[306] ;
input \block[307] ;
input \block[308] ;
input \block[309] ;
input \block[30] ;
input \block[310] ;
input \block[311] ;
input \block[312] ;
input \block[313] ;
input \block[314] ;
input \block[315] ;
input \block[316] ;
input \block[317] ;
input \block[318] ;
input \block[319] ;
input \block[31] ;
input \block[320] ;
input \block[321] ;
input \block[322] ;
input \block[323] ;
input \block[324] ;
input \block[325] ;
input \block[326] ;
input \block[327] ;
input \block[328] ;
input \block[329] ;
input \block[32] ;
input \block[330] ;
input \block[331] ;
input \block[332] ;
input \block[333] ;
input \block[334] ;
input \block[335] ;
input \block[336] ;
input \block[337] ;
input \block[338] ;
input \block[339] ;
input \block[33] ;
input \block[340] ;
input \block[341] ;
input \block[342] ;
input \block[343] ;
input \block[344] ;
input \block[345] ;
input \block[346] ;
input \block[347] ;
input \block[348] ;
input \block[349] ;
input \block[34] ;
input \block[350] ;
input \block[351] ;
input \block[352] ;
input \block[353] ;
input \block[354] ;
input \block[355] ;
input \block[356] ;
input \block[357] ;
input \block[358] ;
input \block[359] ;
input \block[35] ;
input \block[360] ;
input \block[361] ;
input \block[362] ;
input \block[363] ;
input \block[364] ;
input \block[365] ;
input \block[366] ;
input \block[367] ;
input \block[368] ;
input \block[369] ;
input \block[36] ;
input \block[370] ;
input \block[371] ;
input \block[372] ;
input \block[373] ;
input \block[374] ;
input \block[375] ;
input \block[376] ;
input \block[377] ;
input \block[378] ;
input \block[379] ;
input \block[37] ;
input \block[380] ;
input \block[381] ;
input \block[382] ;
input \block[383] ;
input \block[384] ;
input \block[385] ;
input \block[386] ;
input \block[387] ;
input \block[388] ;
input \block[389] ;
input \block[38] ;
input \block[390] ;
input \block[391] ;
input \block[392] ;
input \block[393] ;
input \block[394] ;
input \block[395] ;
input \block[396] ;
input \block[397] ;
input \block[398] ;
input \block[399] ;
input \block[39] ;
input \block[3] ;
input \block[400] ;
input \block[401] ;
input \block[402] ;
input \block[403] ;
input \block[404] ;
input \block[405] ;
input \block[406] ;
input \block[407] ;
input \block[408] ;
input \block[409] ;
input \block[40] ;
input \block[410] ;
input \block[411] ;
input \block[412] ;
input \block[413] ;
input \block[414] ;
input \block[415] ;
input \block[416] ;
input \block[417] ;
input \block[418] ;
input \block[419] ;
input \block[41] ;
input \block[420] ;
input \block[421] ;
input \block[422] ;
input \block[423] ;
input \block[424] ;
input \block[425] ;
input \block[426] ;
input \block[427] ;
input \block[428] ;
input \block[429] ;
input \block[42] ;
input \block[430] ;
input \block[431] ;
input \block[432] ;
input \block[433] ;
input \block[434] ;
input \block[435] ;
input \block[436] ;
input \block[437] ;
input \block[438] ;
input \block[439] ;
input \block[43] ;
input \block[440] ;
input \block[441] ;
input \block[442] ;
input \block[443] ;
input \block[444] ;
input \block[445] ;
input \block[446] ;
input \block[447] ;
input \block[448] ;
input \block[449] ;
input \block[44] ;
input \block[450] ;
input \block[451] ;
input \block[452] ;
input \block[453] ;
input \block[454] ;
input \block[455] ;
input \block[456] ;
input \block[457] ;
input \block[458] ;
input \block[459] ;
input \block[45] ;
input \block[460] ;
input \block[461] ;
input \block[462] ;
input \block[463] ;
input \block[464] ;
input \block[465] ;
input \block[466] ;
input \block[467] ;
input \block[468] ;
input \block[469] ;
input \block[46] ;
input \block[470] ;
input \block[471] ;
input \block[472] ;
input \block[473] ;
input \block[474] ;
input \block[475] ;
input \block[476] ;
input \block[477] ;
input \block[478] ;
input \block[479] ;
input \block[47] ;
input \block[480] ;
input \block[481] ;
input \block[482] ;
input \block[483] ;
input \block[484] ;
input \block[485] ;
input \block[486] ;
input \block[487] ;
input \block[488] ;
input \block[489] ;
input \block[48] ;
input \block[490] ;
input \block[491] ;
input \block[492] ;
input \block[493] ;
input \block[494] ;
input \block[495] ;
input \block[496] ;
input \block[497] ;
input \block[498] ;
input \block[499] ;
input \block[49] ;
input \block[4] ;
input \block[500] ;
input \block[501] ;
input \block[502] ;
input \block[503] ;
input \block[504] ;
input \block[505] ;
input \block[506] ;
input \block[507] ;
input \block[508] ;
input \block[509] ;
input \block[50] ;
input \block[510] ;
input \block[511] ;
input \block[51] ;
input \block[52] ;
input \block[53] ;
input \block[54] ;
input \block[55] ;
input \block[56] ;
input \block[57] ;
input \block[58] ;
input \block[59] ;
input \block[5] ;
input \block[60] ;
input \block[61] ;
input \block[62] ;
input \block[63] ;
input \block[64] ;
input \block[65] ;
input \block[66] ;
input \block[67] ;
input \block[68] ;
input \block[69] ;
input \block[6] ;
input \block[70] ;
input \block[71] ;
input \block[72] ;
input \block[73] ;
input \block[74] ;
input \block[75] ;
input \block[76] ;
input \block[77] ;
input \block[78] ;
input \block[79] ;
input \block[7] ;
input \block[80] ;
input \block[81] ;
input \block[82] ;
input \block[83] ;
input \block[84] ;
input \block[85] ;
input \block[86] ;
input \block[87] ;
input \block[88] ;
input \block[89] ;
input \block[8] ;
input \block[90] ;
input \block[91] ;
input \block[92] ;
input \block[93] ;
input \block[94] ;
input \block[95] ;
input \block[96] ;
input \block[97] ;
input \block[98] ;
input \block[99] ;
input \block[9] ;
wire c_reg_0_; 
wire c_reg_10_; 
wire c_reg_11_; 
wire c_reg_12_; 
wire c_reg_13_; 
wire c_reg_14_; 
wire c_reg_15_; 
wire c_reg_16_; 
wire c_reg_17_; 
wire c_reg_18_; 
wire c_reg_19_; 
wire c_reg_1_; 
wire c_reg_20_; 
wire c_reg_21_; 
wire c_reg_22_; 
wire c_reg_23_; 
wire c_reg_24_; 
wire c_reg_25_; 
wire c_reg_26_; 
wire c_reg_27_; 
wire c_reg_28_; 
wire c_reg_29_; 
wire c_reg_2_; 
wire c_reg_30_; 
wire c_reg_31_; 
wire c_reg_3_; 
wire c_reg_4_; 
wire c_reg_5_; 
wire c_reg_6_; 
wire c_reg_7_; 
wire c_reg_8_; 
wire c_reg_9_; 
input clk;
wire d_reg_0_; 
wire d_reg_10_; 
wire d_reg_11_; 
wire d_reg_12_; 
wire d_reg_13_; 
wire d_reg_14_; 
wire d_reg_15_; 
wire d_reg_16_; 
wire d_reg_17_; 
wire d_reg_18_; 
wire d_reg_19_; 
wire d_reg_1_; 
wire d_reg_20_; 
wire d_reg_21_; 
wire d_reg_22_; 
wire d_reg_23_; 
wire d_reg_24_; 
wire d_reg_25_; 
wire d_reg_26_; 
wire d_reg_27_; 
wire d_reg_28_; 
wire d_reg_29_; 
wire d_reg_2_; 
wire d_reg_30_; 
wire d_reg_31_; 
wire d_reg_3_; 
wire d_reg_4_; 
wire d_reg_5_; 
wire d_reg_6_; 
wire d_reg_7_; 
wire d_reg_8_; 
wire d_reg_9_; 
output \digest[0] ;
output \digest[100] ;
output \digest[101] ;
output \digest[102] ;
output \digest[103] ;
output \digest[104] ;
output \digest[105] ;
output \digest[106] ;
output \digest[107] ;
output \digest[108] ;
output \digest[109] ;
output \digest[10] ;
output \digest[110] ;
output \digest[111] ;
output \digest[112] ;
output \digest[113] ;
output \digest[114] ;
output \digest[115] ;
output \digest[116] ;
output \digest[117] ;
output \digest[118] ;
output \digest[119] ;
output \digest[11] ;
output \digest[120] ;
output \digest[121] ;
output \digest[122] ;
output \digest[123] ;
output \digest[124] ;
output \digest[125] ;
output \digest[126] ;
output \digest[127] ;
output \digest[128] ;
output \digest[129] ;
output \digest[12] ;
output \digest[130] ;
output \digest[131] ;
output \digest[132] ;
output \digest[133] ;
output \digest[134] ;
output \digest[135] ;
output \digest[136] ;
output \digest[137] ;
output \digest[138] ;
output \digest[139] ;
output \digest[13] ;
output \digest[140] ;
output \digest[141] ;
output \digest[142] ;
output \digest[143] ;
output \digest[144] ;
output \digest[145] ;
output \digest[146] ;
output \digest[147] ;
output \digest[148] ;
output \digest[149] ;
output \digest[14] ;
output \digest[150] ;
output \digest[151] ;
output \digest[152] ;
output \digest[153] ;
output \digest[154] ;
output \digest[155] ;
output \digest[156] ;
output \digest[157] ;
output \digest[158] ;
output \digest[159] ;
output \digest[15] ;
output \digest[16] ;
output \digest[17] ;
output \digest[18] ;
output \digest[19] ;
output \digest[1] ;
output \digest[20] ;
output \digest[21] ;
output \digest[22] ;
output \digest[23] ;
output \digest[24] ;
output \digest[25] ;
output \digest[26] ;
output \digest[27] ;
output \digest[28] ;
output \digest[29] ;
output \digest[2] ;
output \digest[30] ;
output \digest[31] ;
output \digest[32] ;
output \digest[33] ;
output \digest[34] ;
output \digest[35] ;
output \digest[36] ;
output \digest[37] ;
output \digest[38] ;
output \digest[39] ;
output \digest[3] ;
output \digest[40] ;
output \digest[41] ;
output \digest[42] ;
output \digest[43] ;
output \digest[44] ;
output \digest[45] ;
output \digest[46] ;
output \digest[47] ;
output \digest[48] ;
output \digest[49] ;
output \digest[4] ;
output \digest[50] ;
output \digest[51] ;
output \digest[52] ;
output \digest[53] ;
output \digest[54] ;
output \digest[55] ;
output \digest[56] ;
output \digest[57] ;
output \digest[58] ;
output \digest[59] ;
output \digest[5] ;
output \digest[60] ;
output \digest[61] ;
output \digest[62] ;
output \digest[63] ;
output \digest[64] ;
output \digest[65] ;
output \digest[66] ;
output \digest[67] ;
output \digest[68] ;
output \digest[69] ;
output \digest[6] ;
output \digest[70] ;
output \digest[71] ;
output \digest[72] ;
output \digest[73] ;
output \digest[74] ;
output \digest[75] ;
output \digest[76] ;
output \digest[77] ;
output \digest[78] ;
output \digest[79] ;
output \digest[7] ;
output \digest[80] ;
output \digest[81] ;
output \digest[82] ;
output \digest[83] ;
output \digest[84] ;
output \digest[85] ;
output \digest[86] ;
output \digest[87] ;
output \digest[88] ;
output \digest[89] ;
output \digest[8] ;
output \digest[90] ;
output \digest[91] ;
output \digest[92] ;
output \digest[93] ;
output \digest[94] ;
output \digest[95] ;
output \digest[96] ;
output \digest[97] ;
output \digest[98] ;
output \digest[99] ;
output \digest[9] ;
wire digest_update; 
output digest_valid;
wire e_reg_0_; 
wire e_reg_10_; 
wire e_reg_11_; 
wire e_reg_12_; 
wire e_reg_13_; 
wire e_reg_14_; 
wire e_reg_15_; 
wire e_reg_16_; 
wire e_reg_17_; 
wire e_reg_18_; 
wire e_reg_19_; 
wire e_reg_1_; 
wire e_reg_20_; 
wire e_reg_21_; 
wire e_reg_22_; 
wire e_reg_23_; 
wire e_reg_24_; 
wire e_reg_25_; 
wire e_reg_26_; 
wire e_reg_27_; 
wire e_reg_28_; 
wire e_reg_29_; 
wire e_reg_2_; 
wire e_reg_30_; 
wire e_reg_31_; 
wire e_reg_3_; 
wire e_reg_4_; 
wire e_reg_5_; 
wire e_reg_6_; 
wire e_reg_7_; 
wire e_reg_8_; 
wire e_reg_9_; 
input init;
input next;
output ready;
input reset_n;
wire round_ctr_inc; 
wire round_ctr_reg_0_; 
wire round_ctr_reg_1_; 
wire round_ctr_reg_2_; 
wire round_ctr_reg_3_; 
wire round_ctr_reg_4_; 
wire round_ctr_reg_5_; 
wire round_ctr_reg_6_; 
wire round_ctr_rst; 
wire w_0_; 
wire w_10_; 
wire w_11_; 
wire w_12_; 
wire w_13_; 
wire w_14_; 
wire w_15_; 
wire w_16_; 
wire w_17_; 
wire w_18_; 
wire w_19_; 
wire w_1_; 
wire w_20_; 
wire w_21_; 
wire w_22_; 
wire w_23_; 
wire w_24_; 
wire w_25_; 
wire w_26_; 
wire w_27_; 
wire w_28_; 
wire w_29_; 
wire w_2_; 
wire w_30_; 
wire w_31_; 
wire w_3_; 
wire w_4_; 
wire w_5_; 
wire w_6_; 
wire w_7_; 
wire w_8_; 
wire w_9_; 
wire w_mem_inst__0w_ctr_reg_6_0__0_; 
wire w_mem_inst__0w_ctr_reg_6_0__1_; 
wire w_mem_inst__0w_ctr_reg_6_0__2_; 
wire w_mem_inst__0w_ctr_reg_6_0__3_; 
wire w_mem_inst__0w_ctr_reg_6_0__4_; 
wire w_mem_inst__0w_ctr_reg_6_0__5_; 
wire w_mem_inst__0w_ctr_reg_6_0__6_; 
wire w_mem_inst__0w_mem_0__31_0__0_; 
wire w_mem_inst__0w_mem_0__31_0__10_; 
wire w_mem_inst__0w_mem_0__31_0__11_; 
wire w_mem_inst__0w_mem_0__31_0__12_; 
wire w_mem_inst__0w_mem_0__31_0__13_; 
wire w_mem_inst__0w_mem_0__31_0__14_; 
wire w_mem_inst__0w_mem_0__31_0__15_; 
wire w_mem_inst__0w_mem_0__31_0__16_; 
wire w_mem_inst__0w_mem_0__31_0__17_; 
wire w_mem_inst__0w_mem_0__31_0__18_; 
wire w_mem_inst__0w_mem_0__31_0__19_; 
wire w_mem_inst__0w_mem_0__31_0__1_; 
wire w_mem_inst__0w_mem_0__31_0__20_; 
wire w_mem_inst__0w_mem_0__31_0__21_; 
wire w_mem_inst__0w_mem_0__31_0__22_; 
wire w_mem_inst__0w_mem_0__31_0__23_; 
wire w_mem_inst__0w_mem_0__31_0__24_; 
wire w_mem_inst__0w_mem_0__31_0__25_; 
wire w_mem_inst__0w_mem_0__31_0__26_; 
wire w_mem_inst__0w_mem_0__31_0__27_; 
wire w_mem_inst__0w_mem_0__31_0__28_; 
wire w_mem_inst__0w_mem_0__31_0__29_; 
wire w_mem_inst__0w_mem_0__31_0__2_; 
wire w_mem_inst__0w_mem_0__31_0__30_; 
wire w_mem_inst__0w_mem_0__31_0__31_; 
wire w_mem_inst__0w_mem_0__31_0__3_; 
wire w_mem_inst__0w_mem_0__31_0__4_; 
wire w_mem_inst__0w_mem_0__31_0__5_; 
wire w_mem_inst__0w_mem_0__31_0__6_; 
wire w_mem_inst__0w_mem_0__31_0__7_; 
wire w_mem_inst__0w_mem_0__31_0__8_; 
wire w_mem_inst__0w_mem_0__31_0__9_; 
wire w_mem_inst__0w_mem_10__31_0__0_; 
wire w_mem_inst__0w_mem_10__31_0__10_; 
wire w_mem_inst__0w_mem_10__31_0__11_; 
wire w_mem_inst__0w_mem_10__31_0__12_; 
wire w_mem_inst__0w_mem_10__31_0__13_; 
wire w_mem_inst__0w_mem_10__31_0__14_; 
wire w_mem_inst__0w_mem_10__31_0__15_; 
wire w_mem_inst__0w_mem_10__31_0__16_; 
wire w_mem_inst__0w_mem_10__31_0__17_; 
wire w_mem_inst__0w_mem_10__31_0__18_; 
wire w_mem_inst__0w_mem_10__31_0__19_; 
wire w_mem_inst__0w_mem_10__31_0__1_; 
wire w_mem_inst__0w_mem_10__31_0__20_; 
wire w_mem_inst__0w_mem_10__31_0__21_; 
wire w_mem_inst__0w_mem_10__31_0__22_; 
wire w_mem_inst__0w_mem_10__31_0__23_; 
wire w_mem_inst__0w_mem_10__31_0__24_; 
wire w_mem_inst__0w_mem_10__31_0__25_; 
wire w_mem_inst__0w_mem_10__31_0__26_; 
wire w_mem_inst__0w_mem_10__31_0__27_; 
wire w_mem_inst__0w_mem_10__31_0__28_; 
wire w_mem_inst__0w_mem_10__31_0__29_; 
wire w_mem_inst__0w_mem_10__31_0__2_; 
wire w_mem_inst__0w_mem_10__31_0__30_; 
wire w_mem_inst__0w_mem_10__31_0__31_; 
wire w_mem_inst__0w_mem_10__31_0__3_; 
wire w_mem_inst__0w_mem_10__31_0__4_; 
wire w_mem_inst__0w_mem_10__31_0__5_; 
wire w_mem_inst__0w_mem_10__31_0__6_; 
wire w_mem_inst__0w_mem_10__31_0__7_; 
wire w_mem_inst__0w_mem_10__31_0__8_; 
wire w_mem_inst__0w_mem_10__31_0__9_; 
wire w_mem_inst__0w_mem_11__31_0__0_; 
wire w_mem_inst__0w_mem_11__31_0__10_; 
wire w_mem_inst__0w_mem_11__31_0__11_; 
wire w_mem_inst__0w_mem_11__31_0__12_; 
wire w_mem_inst__0w_mem_11__31_0__13_; 
wire w_mem_inst__0w_mem_11__31_0__14_; 
wire w_mem_inst__0w_mem_11__31_0__15_; 
wire w_mem_inst__0w_mem_11__31_0__16_; 
wire w_mem_inst__0w_mem_11__31_0__17_; 
wire w_mem_inst__0w_mem_11__31_0__18_; 
wire w_mem_inst__0w_mem_11__31_0__19_; 
wire w_mem_inst__0w_mem_11__31_0__1_; 
wire w_mem_inst__0w_mem_11__31_0__20_; 
wire w_mem_inst__0w_mem_11__31_0__21_; 
wire w_mem_inst__0w_mem_11__31_0__22_; 
wire w_mem_inst__0w_mem_11__31_0__23_; 
wire w_mem_inst__0w_mem_11__31_0__24_; 
wire w_mem_inst__0w_mem_11__31_0__25_; 
wire w_mem_inst__0w_mem_11__31_0__26_; 
wire w_mem_inst__0w_mem_11__31_0__27_; 
wire w_mem_inst__0w_mem_11__31_0__28_; 
wire w_mem_inst__0w_mem_11__31_0__29_; 
wire w_mem_inst__0w_mem_11__31_0__2_; 
wire w_mem_inst__0w_mem_11__31_0__30_; 
wire w_mem_inst__0w_mem_11__31_0__31_; 
wire w_mem_inst__0w_mem_11__31_0__3_; 
wire w_mem_inst__0w_mem_11__31_0__4_; 
wire w_mem_inst__0w_mem_11__31_0__5_; 
wire w_mem_inst__0w_mem_11__31_0__6_; 
wire w_mem_inst__0w_mem_11__31_0__7_; 
wire w_mem_inst__0w_mem_11__31_0__8_; 
wire w_mem_inst__0w_mem_11__31_0__9_; 
wire w_mem_inst__0w_mem_12__31_0__0_; 
wire w_mem_inst__0w_mem_12__31_0__10_; 
wire w_mem_inst__0w_mem_12__31_0__11_; 
wire w_mem_inst__0w_mem_12__31_0__12_; 
wire w_mem_inst__0w_mem_12__31_0__13_; 
wire w_mem_inst__0w_mem_12__31_0__14_; 
wire w_mem_inst__0w_mem_12__31_0__15_; 
wire w_mem_inst__0w_mem_12__31_0__16_; 
wire w_mem_inst__0w_mem_12__31_0__17_; 
wire w_mem_inst__0w_mem_12__31_0__18_; 
wire w_mem_inst__0w_mem_12__31_0__19_; 
wire w_mem_inst__0w_mem_12__31_0__1_; 
wire w_mem_inst__0w_mem_12__31_0__20_; 
wire w_mem_inst__0w_mem_12__31_0__21_; 
wire w_mem_inst__0w_mem_12__31_0__22_; 
wire w_mem_inst__0w_mem_12__31_0__23_; 
wire w_mem_inst__0w_mem_12__31_0__24_; 
wire w_mem_inst__0w_mem_12__31_0__25_; 
wire w_mem_inst__0w_mem_12__31_0__26_; 
wire w_mem_inst__0w_mem_12__31_0__27_; 
wire w_mem_inst__0w_mem_12__31_0__28_; 
wire w_mem_inst__0w_mem_12__31_0__29_; 
wire w_mem_inst__0w_mem_12__31_0__2_; 
wire w_mem_inst__0w_mem_12__31_0__30_; 
wire w_mem_inst__0w_mem_12__31_0__31_; 
wire w_mem_inst__0w_mem_12__31_0__3_; 
wire w_mem_inst__0w_mem_12__31_0__4_; 
wire w_mem_inst__0w_mem_12__31_0__5_; 
wire w_mem_inst__0w_mem_12__31_0__6_; 
wire w_mem_inst__0w_mem_12__31_0__7_; 
wire w_mem_inst__0w_mem_12__31_0__8_; 
wire w_mem_inst__0w_mem_12__31_0__9_; 
wire w_mem_inst__0w_mem_13__31_0__0_; 
wire w_mem_inst__0w_mem_13__31_0__10_; 
wire w_mem_inst__0w_mem_13__31_0__11_; 
wire w_mem_inst__0w_mem_13__31_0__12_; 
wire w_mem_inst__0w_mem_13__31_0__13_; 
wire w_mem_inst__0w_mem_13__31_0__14_; 
wire w_mem_inst__0w_mem_13__31_0__15_; 
wire w_mem_inst__0w_mem_13__31_0__16_; 
wire w_mem_inst__0w_mem_13__31_0__17_; 
wire w_mem_inst__0w_mem_13__31_0__18_; 
wire w_mem_inst__0w_mem_13__31_0__19_; 
wire w_mem_inst__0w_mem_13__31_0__1_; 
wire w_mem_inst__0w_mem_13__31_0__20_; 
wire w_mem_inst__0w_mem_13__31_0__21_; 
wire w_mem_inst__0w_mem_13__31_0__22_; 
wire w_mem_inst__0w_mem_13__31_0__23_; 
wire w_mem_inst__0w_mem_13__31_0__24_; 
wire w_mem_inst__0w_mem_13__31_0__25_; 
wire w_mem_inst__0w_mem_13__31_0__26_; 
wire w_mem_inst__0w_mem_13__31_0__27_; 
wire w_mem_inst__0w_mem_13__31_0__28_; 
wire w_mem_inst__0w_mem_13__31_0__29_; 
wire w_mem_inst__0w_mem_13__31_0__2_; 
wire w_mem_inst__0w_mem_13__31_0__30_; 
wire w_mem_inst__0w_mem_13__31_0__31_; 
wire w_mem_inst__0w_mem_13__31_0__3_; 
wire w_mem_inst__0w_mem_13__31_0__4_; 
wire w_mem_inst__0w_mem_13__31_0__5_; 
wire w_mem_inst__0w_mem_13__31_0__6_; 
wire w_mem_inst__0w_mem_13__31_0__7_; 
wire w_mem_inst__0w_mem_13__31_0__8_; 
wire w_mem_inst__0w_mem_13__31_0__9_; 
wire w_mem_inst__0w_mem_14__31_0__0_; 
wire w_mem_inst__0w_mem_14__31_0__10_; 
wire w_mem_inst__0w_mem_14__31_0__11_; 
wire w_mem_inst__0w_mem_14__31_0__12_; 
wire w_mem_inst__0w_mem_14__31_0__13_; 
wire w_mem_inst__0w_mem_14__31_0__14_; 
wire w_mem_inst__0w_mem_14__31_0__15_; 
wire w_mem_inst__0w_mem_14__31_0__16_; 
wire w_mem_inst__0w_mem_14__31_0__17_; 
wire w_mem_inst__0w_mem_14__31_0__18_; 
wire w_mem_inst__0w_mem_14__31_0__19_; 
wire w_mem_inst__0w_mem_14__31_0__1_; 
wire w_mem_inst__0w_mem_14__31_0__20_; 
wire w_mem_inst__0w_mem_14__31_0__21_; 
wire w_mem_inst__0w_mem_14__31_0__22_; 
wire w_mem_inst__0w_mem_14__31_0__23_; 
wire w_mem_inst__0w_mem_14__31_0__24_; 
wire w_mem_inst__0w_mem_14__31_0__25_; 
wire w_mem_inst__0w_mem_14__31_0__26_; 
wire w_mem_inst__0w_mem_14__31_0__27_; 
wire w_mem_inst__0w_mem_14__31_0__28_; 
wire w_mem_inst__0w_mem_14__31_0__29_; 
wire w_mem_inst__0w_mem_14__31_0__2_; 
wire w_mem_inst__0w_mem_14__31_0__30_; 
wire w_mem_inst__0w_mem_14__31_0__31_; 
wire w_mem_inst__0w_mem_14__31_0__3_; 
wire w_mem_inst__0w_mem_14__31_0__4_; 
wire w_mem_inst__0w_mem_14__31_0__5_; 
wire w_mem_inst__0w_mem_14__31_0__6_; 
wire w_mem_inst__0w_mem_14__31_0__7_; 
wire w_mem_inst__0w_mem_14__31_0__8_; 
wire w_mem_inst__0w_mem_14__31_0__9_; 
wire w_mem_inst__0w_mem_15__31_0__0_; 
wire w_mem_inst__0w_mem_15__31_0__10_; 
wire w_mem_inst__0w_mem_15__31_0__11_; 
wire w_mem_inst__0w_mem_15__31_0__12_; 
wire w_mem_inst__0w_mem_15__31_0__13_; 
wire w_mem_inst__0w_mem_15__31_0__14_; 
wire w_mem_inst__0w_mem_15__31_0__15_; 
wire w_mem_inst__0w_mem_15__31_0__16_; 
wire w_mem_inst__0w_mem_15__31_0__17_; 
wire w_mem_inst__0w_mem_15__31_0__18_; 
wire w_mem_inst__0w_mem_15__31_0__19_; 
wire w_mem_inst__0w_mem_15__31_0__1_; 
wire w_mem_inst__0w_mem_15__31_0__20_; 
wire w_mem_inst__0w_mem_15__31_0__21_; 
wire w_mem_inst__0w_mem_15__31_0__22_; 
wire w_mem_inst__0w_mem_15__31_0__23_; 
wire w_mem_inst__0w_mem_15__31_0__24_; 
wire w_mem_inst__0w_mem_15__31_0__25_; 
wire w_mem_inst__0w_mem_15__31_0__26_; 
wire w_mem_inst__0w_mem_15__31_0__27_; 
wire w_mem_inst__0w_mem_15__31_0__28_; 
wire w_mem_inst__0w_mem_15__31_0__29_; 
wire w_mem_inst__0w_mem_15__31_0__2_; 
wire w_mem_inst__0w_mem_15__31_0__30_; 
wire w_mem_inst__0w_mem_15__31_0__31_; 
wire w_mem_inst__0w_mem_15__31_0__3_; 
wire w_mem_inst__0w_mem_15__31_0__4_; 
wire w_mem_inst__0w_mem_15__31_0__5_; 
wire w_mem_inst__0w_mem_15__31_0__6_; 
wire w_mem_inst__0w_mem_15__31_0__7_; 
wire w_mem_inst__0w_mem_15__31_0__8_; 
wire w_mem_inst__0w_mem_15__31_0__9_; 
wire w_mem_inst__0w_mem_1__31_0__0_; 
wire w_mem_inst__0w_mem_1__31_0__10_; 
wire w_mem_inst__0w_mem_1__31_0__11_; 
wire w_mem_inst__0w_mem_1__31_0__12_; 
wire w_mem_inst__0w_mem_1__31_0__13_; 
wire w_mem_inst__0w_mem_1__31_0__14_; 
wire w_mem_inst__0w_mem_1__31_0__15_; 
wire w_mem_inst__0w_mem_1__31_0__16_; 
wire w_mem_inst__0w_mem_1__31_0__17_; 
wire w_mem_inst__0w_mem_1__31_0__18_; 
wire w_mem_inst__0w_mem_1__31_0__19_; 
wire w_mem_inst__0w_mem_1__31_0__1_; 
wire w_mem_inst__0w_mem_1__31_0__20_; 
wire w_mem_inst__0w_mem_1__31_0__21_; 
wire w_mem_inst__0w_mem_1__31_0__22_; 
wire w_mem_inst__0w_mem_1__31_0__23_; 
wire w_mem_inst__0w_mem_1__31_0__24_; 
wire w_mem_inst__0w_mem_1__31_0__25_; 
wire w_mem_inst__0w_mem_1__31_0__26_; 
wire w_mem_inst__0w_mem_1__31_0__27_; 
wire w_mem_inst__0w_mem_1__31_0__28_; 
wire w_mem_inst__0w_mem_1__31_0__29_; 
wire w_mem_inst__0w_mem_1__31_0__2_; 
wire w_mem_inst__0w_mem_1__31_0__30_; 
wire w_mem_inst__0w_mem_1__31_0__31_; 
wire w_mem_inst__0w_mem_1__31_0__3_; 
wire w_mem_inst__0w_mem_1__31_0__4_; 
wire w_mem_inst__0w_mem_1__31_0__5_; 
wire w_mem_inst__0w_mem_1__31_0__6_; 
wire w_mem_inst__0w_mem_1__31_0__7_; 
wire w_mem_inst__0w_mem_1__31_0__8_; 
wire w_mem_inst__0w_mem_1__31_0__9_; 
wire w_mem_inst__0w_mem_2__31_0__0_; 
wire w_mem_inst__0w_mem_2__31_0__10_; 
wire w_mem_inst__0w_mem_2__31_0__11_; 
wire w_mem_inst__0w_mem_2__31_0__12_; 
wire w_mem_inst__0w_mem_2__31_0__13_; 
wire w_mem_inst__0w_mem_2__31_0__14_; 
wire w_mem_inst__0w_mem_2__31_0__15_; 
wire w_mem_inst__0w_mem_2__31_0__16_; 
wire w_mem_inst__0w_mem_2__31_0__17_; 
wire w_mem_inst__0w_mem_2__31_0__18_; 
wire w_mem_inst__0w_mem_2__31_0__19_; 
wire w_mem_inst__0w_mem_2__31_0__1_; 
wire w_mem_inst__0w_mem_2__31_0__20_; 
wire w_mem_inst__0w_mem_2__31_0__21_; 
wire w_mem_inst__0w_mem_2__31_0__22_; 
wire w_mem_inst__0w_mem_2__31_0__23_; 
wire w_mem_inst__0w_mem_2__31_0__24_; 
wire w_mem_inst__0w_mem_2__31_0__25_; 
wire w_mem_inst__0w_mem_2__31_0__26_; 
wire w_mem_inst__0w_mem_2__31_0__27_; 
wire w_mem_inst__0w_mem_2__31_0__28_; 
wire w_mem_inst__0w_mem_2__31_0__29_; 
wire w_mem_inst__0w_mem_2__31_0__2_; 
wire w_mem_inst__0w_mem_2__31_0__30_; 
wire w_mem_inst__0w_mem_2__31_0__31_; 
wire w_mem_inst__0w_mem_2__31_0__3_; 
wire w_mem_inst__0w_mem_2__31_0__4_; 
wire w_mem_inst__0w_mem_2__31_0__5_; 
wire w_mem_inst__0w_mem_2__31_0__6_; 
wire w_mem_inst__0w_mem_2__31_0__7_; 
wire w_mem_inst__0w_mem_2__31_0__8_; 
wire w_mem_inst__0w_mem_2__31_0__9_; 
wire w_mem_inst__0w_mem_3__31_0__0_; 
wire w_mem_inst__0w_mem_3__31_0__10_; 
wire w_mem_inst__0w_mem_3__31_0__11_; 
wire w_mem_inst__0w_mem_3__31_0__12_; 
wire w_mem_inst__0w_mem_3__31_0__13_; 
wire w_mem_inst__0w_mem_3__31_0__14_; 
wire w_mem_inst__0w_mem_3__31_0__15_; 
wire w_mem_inst__0w_mem_3__31_0__16_; 
wire w_mem_inst__0w_mem_3__31_0__17_; 
wire w_mem_inst__0w_mem_3__31_0__18_; 
wire w_mem_inst__0w_mem_3__31_0__19_; 
wire w_mem_inst__0w_mem_3__31_0__1_; 
wire w_mem_inst__0w_mem_3__31_0__20_; 
wire w_mem_inst__0w_mem_3__31_0__21_; 
wire w_mem_inst__0w_mem_3__31_0__22_; 
wire w_mem_inst__0w_mem_3__31_0__23_; 
wire w_mem_inst__0w_mem_3__31_0__24_; 
wire w_mem_inst__0w_mem_3__31_0__25_; 
wire w_mem_inst__0w_mem_3__31_0__26_; 
wire w_mem_inst__0w_mem_3__31_0__27_; 
wire w_mem_inst__0w_mem_3__31_0__28_; 
wire w_mem_inst__0w_mem_3__31_0__29_; 
wire w_mem_inst__0w_mem_3__31_0__2_; 
wire w_mem_inst__0w_mem_3__31_0__30_; 
wire w_mem_inst__0w_mem_3__31_0__31_; 
wire w_mem_inst__0w_mem_3__31_0__3_; 
wire w_mem_inst__0w_mem_3__31_0__4_; 
wire w_mem_inst__0w_mem_3__31_0__5_; 
wire w_mem_inst__0w_mem_3__31_0__6_; 
wire w_mem_inst__0w_mem_3__31_0__7_; 
wire w_mem_inst__0w_mem_3__31_0__8_; 
wire w_mem_inst__0w_mem_3__31_0__9_; 
wire w_mem_inst__0w_mem_4__31_0__0_; 
wire w_mem_inst__0w_mem_4__31_0__10_; 
wire w_mem_inst__0w_mem_4__31_0__11_; 
wire w_mem_inst__0w_mem_4__31_0__12_; 
wire w_mem_inst__0w_mem_4__31_0__13_; 
wire w_mem_inst__0w_mem_4__31_0__14_; 
wire w_mem_inst__0w_mem_4__31_0__15_; 
wire w_mem_inst__0w_mem_4__31_0__16_; 
wire w_mem_inst__0w_mem_4__31_0__17_; 
wire w_mem_inst__0w_mem_4__31_0__18_; 
wire w_mem_inst__0w_mem_4__31_0__19_; 
wire w_mem_inst__0w_mem_4__31_0__1_; 
wire w_mem_inst__0w_mem_4__31_0__20_; 
wire w_mem_inst__0w_mem_4__31_0__21_; 
wire w_mem_inst__0w_mem_4__31_0__22_; 
wire w_mem_inst__0w_mem_4__31_0__23_; 
wire w_mem_inst__0w_mem_4__31_0__24_; 
wire w_mem_inst__0w_mem_4__31_0__25_; 
wire w_mem_inst__0w_mem_4__31_0__26_; 
wire w_mem_inst__0w_mem_4__31_0__27_; 
wire w_mem_inst__0w_mem_4__31_0__28_; 
wire w_mem_inst__0w_mem_4__31_0__29_; 
wire w_mem_inst__0w_mem_4__31_0__2_; 
wire w_mem_inst__0w_mem_4__31_0__30_; 
wire w_mem_inst__0w_mem_4__31_0__31_; 
wire w_mem_inst__0w_mem_4__31_0__3_; 
wire w_mem_inst__0w_mem_4__31_0__4_; 
wire w_mem_inst__0w_mem_4__31_0__5_; 
wire w_mem_inst__0w_mem_4__31_0__6_; 
wire w_mem_inst__0w_mem_4__31_0__7_; 
wire w_mem_inst__0w_mem_4__31_0__8_; 
wire w_mem_inst__0w_mem_4__31_0__9_; 
wire w_mem_inst__0w_mem_5__31_0__0_; 
wire w_mem_inst__0w_mem_5__31_0__10_; 
wire w_mem_inst__0w_mem_5__31_0__11_; 
wire w_mem_inst__0w_mem_5__31_0__12_; 
wire w_mem_inst__0w_mem_5__31_0__13_; 
wire w_mem_inst__0w_mem_5__31_0__14_; 
wire w_mem_inst__0w_mem_5__31_0__15_; 
wire w_mem_inst__0w_mem_5__31_0__16_; 
wire w_mem_inst__0w_mem_5__31_0__17_; 
wire w_mem_inst__0w_mem_5__31_0__18_; 
wire w_mem_inst__0w_mem_5__31_0__19_; 
wire w_mem_inst__0w_mem_5__31_0__1_; 
wire w_mem_inst__0w_mem_5__31_0__20_; 
wire w_mem_inst__0w_mem_5__31_0__21_; 
wire w_mem_inst__0w_mem_5__31_0__22_; 
wire w_mem_inst__0w_mem_5__31_0__23_; 
wire w_mem_inst__0w_mem_5__31_0__24_; 
wire w_mem_inst__0w_mem_5__31_0__25_; 
wire w_mem_inst__0w_mem_5__31_0__26_; 
wire w_mem_inst__0w_mem_5__31_0__27_; 
wire w_mem_inst__0w_mem_5__31_0__28_; 
wire w_mem_inst__0w_mem_5__31_0__29_; 
wire w_mem_inst__0w_mem_5__31_0__2_; 
wire w_mem_inst__0w_mem_5__31_0__30_; 
wire w_mem_inst__0w_mem_5__31_0__31_; 
wire w_mem_inst__0w_mem_5__31_0__3_; 
wire w_mem_inst__0w_mem_5__31_0__4_; 
wire w_mem_inst__0w_mem_5__31_0__5_; 
wire w_mem_inst__0w_mem_5__31_0__6_; 
wire w_mem_inst__0w_mem_5__31_0__7_; 
wire w_mem_inst__0w_mem_5__31_0__8_; 
wire w_mem_inst__0w_mem_5__31_0__9_; 
wire w_mem_inst__0w_mem_6__31_0__0_; 
wire w_mem_inst__0w_mem_6__31_0__10_; 
wire w_mem_inst__0w_mem_6__31_0__11_; 
wire w_mem_inst__0w_mem_6__31_0__12_; 
wire w_mem_inst__0w_mem_6__31_0__13_; 
wire w_mem_inst__0w_mem_6__31_0__14_; 
wire w_mem_inst__0w_mem_6__31_0__15_; 
wire w_mem_inst__0w_mem_6__31_0__16_; 
wire w_mem_inst__0w_mem_6__31_0__17_; 
wire w_mem_inst__0w_mem_6__31_0__18_; 
wire w_mem_inst__0w_mem_6__31_0__19_; 
wire w_mem_inst__0w_mem_6__31_0__1_; 
wire w_mem_inst__0w_mem_6__31_0__20_; 
wire w_mem_inst__0w_mem_6__31_0__21_; 
wire w_mem_inst__0w_mem_6__31_0__22_; 
wire w_mem_inst__0w_mem_6__31_0__23_; 
wire w_mem_inst__0w_mem_6__31_0__24_; 
wire w_mem_inst__0w_mem_6__31_0__25_; 
wire w_mem_inst__0w_mem_6__31_0__26_; 
wire w_mem_inst__0w_mem_6__31_0__27_; 
wire w_mem_inst__0w_mem_6__31_0__28_; 
wire w_mem_inst__0w_mem_6__31_0__29_; 
wire w_mem_inst__0w_mem_6__31_0__2_; 
wire w_mem_inst__0w_mem_6__31_0__30_; 
wire w_mem_inst__0w_mem_6__31_0__31_; 
wire w_mem_inst__0w_mem_6__31_0__3_; 
wire w_mem_inst__0w_mem_6__31_0__4_; 
wire w_mem_inst__0w_mem_6__31_0__5_; 
wire w_mem_inst__0w_mem_6__31_0__6_; 
wire w_mem_inst__0w_mem_6__31_0__7_; 
wire w_mem_inst__0w_mem_6__31_0__8_; 
wire w_mem_inst__0w_mem_6__31_0__9_; 
wire w_mem_inst__0w_mem_7__31_0__0_; 
wire w_mem_inst__0w_mem_7__31_0__10_; 
wire w_mem_inst__0w_mem_7__31_0__11_; 
wire w_mem_inst__0w_mem_7__31_0__12_; 
wire w_mem_inst__0w_mem_7__31_0__13_; 
wire w_mem_inst__0w_mem_7__31_0__14_; 
wire w_mem_inst__0w_mem_7__31_0__15_; 
wire w_mem_inst__0w_mem_7__31_0__16_; 
wire w_mem_inst__0w_mem_7__31_0__17_; 
wire w_mem_inst__0w_mem_7__31_0__18_; 
wire w_mem_inst__0w_mem_7__31_0__19_; 
wire w_mem_inst__0w_mem_7__31_0__1_; 
wire w_mem_inst__0w_mem_7__31_0__20_; 
wire w_mem_inst__0w_mem_7__31_0__21_; 
wire w_mem_inst__0w_mem_7__31_0__22_; 
wire w_mem_inst__0w_mem_7__31_0__23_; 
wire w_mem_inst__0w_mem_7__31_0__24_; 
wire w_mem_inst__0w_mem_7__31_0__25_; 
wire w_mem_inst__0w_mem_7__31_0__26_; 
wire w_mem_inst__0w_mem_7__31_0__27_; 
wire w_mem_inst__0w_mem_7__31_0__28_; 
wire w_mem_inst__0w_mem_7__31_0__29_; 
wire w_mem_inst__0w_mem_7__31_0__2_; 
wire w_mem_inst__0w_mem_7__31_0__30_; 
wire w_mem_inst__0w_mem_7__31_0__31_; 
wire w_mem_inst__0w_mem_7__31_0__3_; 
wire w_mem_inst__0w_mem_7__31_0__4_; 
wire w_mem_inst__0w_mem_7__31_0__5_; 
wire w_mem_inst__0w_mem_7__31_0__6_; 
wire w_mem_inst__0w_mem_7__31_0__7_; 
wire w_mem_inst__0w_mem_7__31_0__8_; 
wire w_mem_inst__0w_mem_7__31_0__9_; 
wire w_mem_inst__0w_mem_8__31_0__0_; 
wire w_mem_inst__0w_mem_8__31_0__10_; 
wire w_mem_inst__0w_mem_8__31_0__11_; 
wire w_mem_inst__0w_mem_8__31_0__12_; 
wire w_mem_inst__0w_mem_8__31_0__13_; 
wire w_mem_inst__0w_mem_8__31_0__14_; 
wire w_mem_inst__0w_mem_8__31_0__15_; 
wire w_mem_inst__0w_mem_8__31_0__16_; 
wire w_mem_inst__0w_mem_8__31_0__17_; 
wire w_mem_inst__0w_mem_8__31_0__18_; 
wire w_mem_inst__0w_mem_8__31_0__19_; 
wire w_mem_inst__0w_mem_8__31_0__1_; 
wire w_mem_inst__0w_mem_8__31_0__20_; 
wire w_mem_inst__0w_mem_8__31_0__21_; 
wire w_mem_inst__0w_mem_8__31_0__22_; 
wire w_mem_inst__0w_mem_8__31_0__23_; 
wire w_mem_inst__0w_mem_8__31_0__24_; 
wire w_mem_inst__0w_mem_8__31_0__25_; 
wire w_mem_inst__0w_mem_8__31_0__26_; 
wire w_mem_inst__0w_mem_8__31_0__27_; 
wire w_mem_inst__0w_mem_8__31_0__28_; 
wire w_mem_inst__0w_mem_8__31_0__29_; 
wire w_mem_inst__0w_mem_8__31_0__2_; 
wire w_mem_inst__0w_mem_8__31_0__30_; 
wire w_mem_inst__0w_mem_8__31_0__31_; 
wire w_mem_inst__0w_mem_8__31_0__3_; 
wire w_mem_inst__0w_mem_8__31_0__4_; 
wire w_mem_inst__0w_mem_8__31_0__5_; 
wire w_mem_inst__0w_mem_8__31_0__6_; 
wire w_mem_inst__0w_mem_8__31_0__7_; 
wire w_mem_inst__0w_mem_8__31_0__8_; 
wire w_mem_inst__0w_mem_8__31_0__9_; 
wire w_mem_inst__0w_mem_9__31_0__0_; 
wire w_mem_inst__0w_mem_9__31_0__10_; 
wire w_mem_inst__0w_mem_9__31_0__11_; 
wire w_mem_inst__0w_mem_9__31_0__12_; 
wire w_mem_inst__0w_mem_9__31_0__13_; 
wire w_mem_inst__0w_mem_9__31_0__14_; 
wire w_mem_inst__0w_mem_9__31_0__15_; 
wire w_mem_inst__0w_mem_9__31_0__16_; 
wire w_mem_inst__0w_mem_9__31_0__17_; 
wire w_mem_inst__0w_mem_9__31_0__18_; 
wire w_mem_inst__0w_mem_9__31_0__19_; 
wire w_mem_inst__0w_mem_9__31_0__1_; 
wire w_mem_inst__0w_mem_9__31_0__20_; 
wire w_mem_inst__0w_mem_9__31_0__21_; 
wire w_mem_inst__0w_mem_9__31_0__22_; 
wire w_mem_inst__0w_mem_9__31_0__23_; 
wire w_mem_inst__0w_mem_9__31_0__24_; 
wire w_mem_inst__0w_mem_9__31_0__25_; 
wire w_mem_inst__0w_mem_9__31_0__26_; 
wire w_mem_inst__0w_mem_9__31_0__27_; 
wire w_mem_inst__0w_mem_9__31_0__28_; 
wire w_mem_inst__0w_mem_9__31_0__29_; 
wire w_mem_inst__0w_mem_9__31_0__2_; 
wire w_mem_inst__0w_mem_9__31_0__30_; 
wire w_mem_inst__0w_mem_9__31_0__31_; 
wire w_mem_inst__0w_mem_9__31_0__3_; 
wire w_mem_inst__0w_mem_9__31_0__4_; 
wire w_mem_inst__0w_mem_9__31_0__5_; 
wire w_mem_inst__0w_mem_9__31_0__6_; 
wire w_mem_inst__0w_mem_9__31_0__7_; 
wire w_mem_inst__0w_mem_9__31_0__8_; 
wire w_mem_inst__0w_mem_9__31_0__9_; 
wire w_mem_inst__abc_21203_new_n1585_; 
wire w_mem_inst__abc_21203_new_n1586_; 
wire w_mem_inst__abc_21203_new_n1587_; 
wire w_mem_inst__abc_21203_new_n1588_; 
wire w_mem_inst__abc_21203_new_n1589_; 
wire w_mem_inst__abc_21203_new_n1590_; 
wire w_mem_inst__abc_21203_new_n1591_; 
wire w_mem_inst__abc_21203_new_n1592_; 
wire w_mem_inst__abc_21203_new_n1593_; 
wire w_mem_inst__abc_21203_new_n1594_; 
wire w_mem_inst__abc_21203_new_n1595_; 
wire w_mem_inst__abc_21203_new_n1596_; 
wire w_mem_inst__abc_21203_new_n1597_; 
wire w_mem_inst__abc_21203_new_n1598_; 
wire w_mem_inst__abc_21203_new_n1599_; 
wire w_mem_inst__abc_21203_new_n1600_; 
wire w_mem_inst__abc_21203_new_n1601_; 
wire w_mem_inst__abc_21203_new_n1602_; 
wire w_mem_inst__abc_21203_new_n1603_; 
wire w_mem_inst__abc_21203_new_n1604_; 
wire w_mem_inst__abc_21203_new_n1605_; 
wire w_mem_inst__abc_21203_new_n1606_; 
wire w_mem_inst__abc_21203_new_n1607_; 
wire w_mem_inst__abc_21203_new_n1608_; 
wire w_mem_inst__abc_21203_new_n1609_; 
wire w_mem_inst__abc_21203_new_n1610_; 
wire w_mem_inst__abc_21203_new_n1611_; 
wire w_mem_inst__abc_21203_new_n1612_; 
wire w_mem_inst__abc_21203_new_n1613_; 
wire w_mem_inst__abc_21203_new_n1614_; 
wire w_mem_inst__abc_21203_new_n1615_; 
wire w_mem_inst__abc_21203_new_n1616_; 
wire w_mem_inst__abc_21203_new_n1617_; 
wire w_mem_inst__abc_21203_new_n1618_; 
wire w_mem_inst__abc_21203_new_n1619_; 
wire w_mem_inst__abc_21203_new_n1620_; 
wire w_mem_inst__abc_21203_new_n1621_; 
wire w_mem_inst__abc_21203_new_n1622_; 
wire w_mem_inst__abc_21203_new_n1623_; 
wire w_mem_inst__abc_21203_new_n1624_; 
wire w_mem_inst__abc_21203_new_n1625_; 
wire w_mem_inst__abc_21203_new_n1626_; 
wire w_mem_inst__abc_21203_new_n1627_; 
wire w_mem_inst__abc_21203_new_n1628_; 
wire w_mem_inst__abc_21203_new_n1629_; 
wire w_mem_inst__abc_21203_new_n1630_; 
wire w_mem_inst__abc_21203_new_n1631_; 
wire w_mem_inst__abc_21203_new_n1632_; 
wire w_mem_inst__abc_21203_new_n1633_; 
wire w_mem_inst__abc_21203_new_n1634_; 
wire w_mem_inst__abc_21203_new_n1635_; 
wire w_mem_inst__abc_21203_new_n1636_; 
wire w_mem_inst__abc_21203_new_n1637_; 
wire w_mem_inst__abc_21203_new_n1638_; 
wire w_mem_inst__abc_21203_new_n1639_; 
wire w_mem_inst__abc_21203_new_n1640_; 
wire w_mem_inst__abc_21203_new_n1641_; 
wire w_mem_inst__abc_21203_new_n1642_; 
wire w_mem_inst__abc_21203_new_n1643_; 
wire w_mem_inst__abc_21203_new_n1644_; 
wire w_mem_inst__abc_21203_new_n1645_; 
wire w_mem_inst__abc_21203_new_n1646_; 
wire w_mem_inst__abc_21203_new_n1647_; 
wire w_mem_inst__abc_21203_new_n1648_; 
wire w_mem_inst__abc_21203_new_n1649_; 
wire w_mem_inst__abc_21203_new_n1650_; 
wire w_mem_inst__abc_21203_new_n1651_; 
wire w_mem_inst__abc_21203_new_n1652_; 
wire w_mem_inst__abc_21203_new_n1653_; 
wire w_mem_inst__abc_21203_new_n1654_; 
wire w_mem_inst__abc_21203_new_n1655_; 
wire w_mem_inst__abc_21203_new_n1656_; 
wire w_mem_inst__abc_21203_new_n1657_; 
wire w_mem_inst__abc_21203_new_n1658_; 
wire w_mem_inst__abc_21203_new_n1659_; 
wire w_mem_inst__abc_21203_new_n1660_; 
wire w_mem_inst__abc_21203_new_n1661_; 
wire w_mem_inst__abc_21203_new_n1662_; 
wire w_mem_inst__abc_21203_new_n1664_; 
wire w_mem_inst__abc_21203_new_n1665_; 
wire w_mem_inst__abc_21203_new_n1666_; 
wire w_mem_inst__abc_21203_new_n1667_; 
wire w_mem_inst__abc_21203_new_n1668_; 
wire w_mem_inst__abc_21203_new_n1669_; 
wire w_mem_inst__abc_21203_new_n1670_; 
wire w_mem_inst__abc_21203_new_n1671_; 
wire w_mem_inst__abc_21203_new_n1672_; 
wire w_mem_inst__abc_21203_new_n1673_; 
wire w_mem_inst__abc_21203_new_n1674_; 
wire w_mem_inst__abc_21203_new_n1675_; 
wire w_mem_inst__abc_21203_new_n1676_; 
wire w_mem_inst__abc_21203_new_n1677_; 
wire w_mem_inst__abc_21203_new_n1678_; 
wire w_mem_inst__abc_21203_new_n1679_; 
wire w_mem_inst__abc_21203_new_n1680_; 
wire w_mem_inst__abc_21203_new_n1681_; 
wire w_mem_inst__abc_21203_new_n1682_; 
wire w_mem_inst__abc_21203_new_n1683_; 
wire w_mem_inst__abc_21203_new_n1684_; 
wire w_mem_inst__abc_21203_new_n1685_; 
wire w_mem_inst__abc_21203_new_n1686_; 
wire w_mem_inst__abc_21203_new_n1687_; 
wire w_mem_inst__abc_21203_new_n1688_; 
wire w_mem_inst__abc_21203_new_n1689_; 
wire w_mem_inst__abc_21203_new_n1690_; 
wire w_mem_inst__abc_21203_new_n1691_; 
wire w_mem_inst__abc_21203_new_n1692_; 
wire w_mem_inst__abc_21203_new_n1693_; 
wire w_mem_inst__abc_21203_new_n1694_; 
wire w_mem_inst__abc_21203_new_n1695_; 
wire w_mem_inst__abc_21203_new_n1696_; 
wire w_mem_inst__abc_21203_new_n1697_; 
wire w_mem_inst__abc_21203_new_n1698_; 
wire w_mem_inst__abc_21203_new_n1699_; 
wire w_mem_inst__abc_21203_new_n1700_; 
wire w_mem_inst__abc_21203_new_n1701_; 
wire w_mem_inst__abc_21203_new_n1702_; 
wire w_mem_inst__abc_21203_new_n1703_; 
wire w_mem_inst__abc_21203_new_n1704_; 
wire w_mem_inst__abc_21203_new_n1705_; 
wire w_mem_inst__abc_21203_new_n1706_; 
wire w_mem_inst__abc_21203_new_n1707_; 
wire w_mem_inst__abc_21203_new_n1708_; 
wire w_mem_inst__abc_21203_new_n1709_; 
wire w_mem_inst__abc_21203_new_n1710_; 
wire w_mem_inst__abc_21203_new_n1712_; 
wire w_mem_inst__abc_21203_new_n1713_; 
wire w_mem_inst__abc_21203_new_n1714_; 
wire w_mem_inst__abc_21203_new_n1715_; 
wire w_mem_inst__abc_21203_new_n1716_; 
wire w_mem_inst__abc_21203_new_n1717_; 
wire w_mem_inst__abc_21203_new_n1718_; 
wire w_mem_inst__abc_21203_new_n1719_; 
wire w_mem_inst__abc_21203_new_n1720_; 
wire w_mem_inst__abc_21203_new_n1721_; 
wire w_mem_inst__abc_21203_new_n1722_; 
wire w_mem_inst__abc_21203_new_n1723_; 
wire w_mem_inst__abc_21203_new_n1724_; 
wire w_mem_inst__abc_21203_new_n1725_; 
wire w_mem_inst__abc_21203_new_n1726_; 
wire w_mem_inst__abc_21203_new_n1727_; 
wire w_mem_inst__abc_21203_new_n1728_; 
wire w_mem_inst__abc_21203_new_n1729_; 
wire w_mem_inst__abc_21203_new_n1730_; 
wire w_mem_inst__abc_21203_new_n1731_; 
wire w_mem_inst__abc_21203_new_n1732_; 
wire w_mem_inst__abc_21203_new_n1733_; 
wire w_mem_inst__abc_21203_new_n1734_; 
wire w_mem_inst__abc_21203_new_n1735_; 
wire w_mem_inst__abc_21203_new_n1736_; 
wire w_mem_inst__abc_21203_new_n1737_; 
wire w_mem_inst__abc_21203_new_n1738_; 
wire w_mem_inst__abc_21203_new_n1739_; 
wire w_mem_inst__abc_21203_new_n1740_; 
wire w_mem_inst__abc_21203_new_n1741_; 
wire w_mem_inst__abc_21203_new_n1742_; 
wire w_mem_inst__abc_21203_new_n1743_; 
wire w_mem_inst__abc_21203_new_n1744_; 
wire w_mem_inst__abc_21203_new_n1745_; 
wire w_mem_inst__abc_21203_new_n1746_; 
wire w_mem_inst__abc_21203_new_n1747_; 
wire w_mem_inst__abc_21203_new_n1748_; 
wire w_mem_inst__abc_21203_new_n1749_; 
wire w_mem_inst__abc_21203_new_n1750_; 
wire w_mem_inst__abc_21203_new_n1751_; 
wire w_mem_inst__abc_21203_new_n1752_; 
wire w_mem_inst__abc_21203_new_n1753_; 
wire w_mem_inst__abc_21203_new_n1754_; 
wire w_mem_inst__abc_21203_new_n1755_; 
wire w_mem_inst__abc_21203_new_n1756_; 
wire w_mem_inst__abc_21203_new_n1757_; 
wire w_mem_inst__abc_21203_new_n1758_; 
wire w_mem_inst__abc_21203_new_n1760_; 
wire w_mem_inst__abc_21203_new_n1761_; 
wire w_mem_inst__abc_21203_new_n1762_; 
wire w_mem_inst__abc_21203_new_n1763_; 
wire w_mem_inst__abc_21203_new_n1764_; 
wire w_mem_inst__abc_21203_new_n1765_; 
wire w_mem_inst__abc_21203_new_n1766_; 
wire w_mem_inst__abc_21203_new_n1767_; 
wire w_mem_inst__abc_21203_new_n1768_; 
wire w_mem_inst__abc_21203_new_n1769_; 
wire w_mem_inst__abc_21203_new_n1770_; 
wire w_mem_inst__abc_21203_new_n1771_; 
wire w_mem_inst__abc_21203_new_n1772_; 
wire w_mem_inst__abc_21203_new_n1773_; 
wire w_mem_inst__abc_21203_new_n1774_; 
wire w_mem_inst__abc_21203_new_n1775_; 
wire w_mem_inst__abc_21203_new_n1776_; 
wire w_mem_inst__abc_21203_new_n1777_; 
wire w_mem_inst__abc_21203_new_n1778_; 
wire w_mem_inst__abc_21203_new_n1779_; 
wire w_mem_inst__abc_21203_new_n1780_; 
wire w_mem_inst__abc_21203_new_n1781_; 
wire w_mem_inst__abc_21203_new_n1782_; 
wire w_mem_inst__abc_21203_new_n1783_; 
wire w_mem_inst__abc_21203_new_n1784_; 
wire w_mem_inst__abc_21203_new_n1785_; 
wire w_mem_inst__abc_21203_new_n1786_; 
wire w_mem_inst__abc_21203_new_n1787_; 
wire w_mem_inst__abc_21203_new_n1788_; 
wire w_mem_inst__abc_21203_new_n1789_; 
wire w_mem_inst__abc_21203_new_n1790_; 
wire w_mem_inst__abc_21203_new_n1791_; 
wire w_mem_inst__abc_21203_new_n1792_; 
wire w_mem_inst__abc_21203_new_n1793_; 
wire w_mem_inst__abc_21203_new_n1794_; 
wire w_mem_inst__abc_21203_new_n1795_; 
wire w_mem_inst__abc_21203_new_n1796_; 
wire w_mem_inst__abc_21203_new_n1797_; 
wire w_mem_inst__abc_21203_new_n1798_; 
wire w_mem_inst__abc_21203_new_n1799_; 
wire w_mem_inst__abc_21203_new_n1800_; 
wire w_mem_inst__abc_21203_new_n1801_; 
wire w_mem_inst__abc_21203_new_n1802_; 
wire w_mem_inst__abc_21203_new_n1803_; 
wire w_mem_inst__abc_21203_new_n1804_; 
wire w_mem_inst__abc_21203_new_n1805_; 
wire w_mem_inst__abc_21203_new_n1806_; 
wire w_mem_inst__abc_21203_new_n1808_; 
wire w_mem_inst__abc_21203_new_n1809_; 
wire w_mem_inst__abc_21203_new_n1810_; 
wire w_mem_inst__abc_21203_new_n1811_; 
wire w_mem_inst__abc_21203_new_n1812_; 
wire w_mem_inst__abc_21203_new_n1813_; 
wire w_mem_inst__abc_21203_new_n1814_; 
wire w_mem_inst__abc_21203_new_n1815_; 
wire w_mem_inst__abc_21203_new_n1816_; 
wire w_mem_inst__abc_21203_new_n1817_; 
wire w_mem_inst__abc_21203_new_n1818_; 
wire w_mem_inst__abc_21203_new_n1819_; 
wire w_mem_inst__abc_21203_new_n1820_; 
wire w_mem_inst__abc_21203_new_n1821_; 
wire w_mem_inst__abc_21203_new_n1822_; 
wire w_mem_inst__abc_21203_new_n1823_; 
wire w_mem_inst__abc_21203_new_n1824_; 
wire w_mem_inst__abc_21203_new_n1825_; 
wire w_mem_inst__abc_21203_new_n1826_; 
wire w_mem_inst__abc_21203_new_n1827_; 
wire w_mem_inst__abc_21203_new_n1828_; 
wire w_mem_inst__abc_21203_new_n1829_; 
wire w_mem_inst__abc_21203_new_n1830_; 
wire w_mem_inst__abc_21203_new_n1831_; 
wire w_mem_inst__abc_21203_new_n1832_; 
wire w_mem_inst__abc_21203_new_n1833_; 
wire w_mem_inst__abc_21203_new_n1834_; 
wire w_mem_inst__abc_21203_new_n1835_; 
wire w_mem_inst__abc_21203_new_n1836_; 
wire w_mem_inst__abc_21203_new_n1837_; 
wire w_mem_inst__abc_21203_new_n1838_; 
wire w_mem_inst__abc_21203_new_n1839_; 
wire w_mem_inst__abc_21203_new_n1840_; 
wire w_mem_inst__abc_21203_new_n1841_; 
wire w_mem_inst__abc_21203_new_n1842_; 
wire w_mem_inst__abc_21203_new_n1843_; 
wire w_mem_inst__abc_21203_new_n1844_; 
wire w_mem_inst__abc_21203_new_n1845_; 
wire w_mem_inst__abc_21203_new_n1846_; 
wire w_mem_inst__abc_21203_new_n1847_; 
wire w_mem_inst__abc_21203_new_n1848_; 
wire w_mem_inst__abc_21203_new_n1849_; 
wire w_mem_inst__abc_21203_new_n1850_; 
wire w_mem_inst__abc_21203_new_n1851_; 
wire w_mem_inst__abc_21203_new_n1852_; 
wire w_mem_inst__abc_21203_new_n1853_; 
wire w_mem_inst__abc_21203_new_n1854_; 
wire w_mem_inst__abc_21203_new_n1856_; 
wire w_mem_inst__abc_21203_new_n1857_; 
wire w_mem_inst__abc_21203_new_n1858_; 
wire w_mem_inst__abc_21203_new_n1859_; 
wire w_mem_inst__abc_21203_new_n1860_; 
wire w_mem_inst__abc_21203_new_n1861_; 
wire w_mem_inst__abc_21203_new_n1862_; 
wire w_mem_inst__abc_21203_new_n1863_; 
wire w_mem_inst__abc_21203_new_n1864_; 
wire w_mem_inst__abc_21203_new_n1865_; 
wire w_mem_inst__abc_21203_new_n1866_; 
wire w_mem_inst__abc_21203_new_n1867_; 
wire w_mem_inst__abc_21203_new_n1868_; 
wire w_mem_inst__abc_21203_new_n1869_; 
wire w_mem_inst__abc_21203_new_n1870_; 
wire w_mem_inst__abc_21203_new_n1871_; 
wire w_mem_inst__abc_21203_new_n1872_; 
wire w_mem_inst__abc_21203_new_n1873_; 
wire w_mem_inst__abc_21203_new_n1874_; 
wire w_mem_inst__abc_21203_new_n1875_; 
wire w_mem_inst__abc_21203_new_n1876_; 
wire w_mem_inst__abc_21203_new_n1877_; 
wire w_mem_inst__abc_21203_new_n1878_; 
wire w_mem_inst__abc_21203_new_n1879_; 
wire w_mem_inst__abc_21203_new_n1880_; 
wire w_mem_inst__abc_21203_new_n1881_; 
wire w_mem_inst__abc_21203_new_n1882_; 
wire w_mem_inst__abc_21203_new_n1883_; 
wire w_mem_inst__abc_21203_new_n1884_; 
wire w_mem_inst__abc_21203_new_n1885_; 
wire w_mem_inst__abc_21203_new_n1886_; 
wire w_mem_inst__abc_21203_new_n1887_; 
wire w_mem_inst__abc_21203_new_n1888_; 
wire w_mem_inst__abc_21203_new_n1889_; 
wire w_mem_inst__abc_21203_new_n1890_; 
wire w_mem_inst__abc_21203_new_n1891_; 
wire w_mem_inst__abc_21203_new_n1892_; 
wire w_mem_inst__abc_21203_new_n1893_; 
wire w_mem_inst__abc_21203_new_n1894_; 
wire w_mem_inst__abc_21203_new_n1895_; 
wire w_mem_inst__abc_21203_new_n1896_; 
wire w_mem_inst__abc_21203_new_n1897_; 
wire w_mem_inst__abc_21203_new_n1898_; 
wire w_mem_inst__abc_21203_new_n1899_; 
wire w_mem_inst__abc_21203_new_n1900_; 
wire w_mem_inst__abc_21203_new_n1901_; 
wire w_mem_inst__abc_21203_new_n1902_; 
wire w_mem_inst__abc_21203_new_n1904_; 
wire w_mem_inst__abc_21203_new_n1905_; 
wire w_mem_inst__abc_21203_new_n1906_; 
wire w_mem_inst__abc_21203_new_n1907_; 
wire w_mem_inst__abc_21203_new_n1908_; 
wire w_mem_inst__abc_21203_new_n1909_; 
wire w_mem_inst__abc_21203_new_n1910_; 
wire w_mem_inst__abc_21203_new_n1911_; 
wire w_mem_inst__abc_21203_new_n1912_; 
wire w_mem_inst__abc_21203_new_n1913_; 
wire w_mem_inst__abc_21203_new_n1914_; 
wire w_mem_inst__abc_21203_new_n1915_; 
wire w_mem_inst__abc_21203_new_n1916_; 
wire w_mem_inst__abc_21203_new_n1917_; 
wire w_mem_inst__abc_21203_new_n1918_; 
wire w_mem_inst__abc_21203_new_n1919_; 
wire w_mem_inst__abc_21203_new_n1920_; 
wire w_mem_inst__abc_21203_new_n1921_; 
wire w_mem_inst__abc_21203_new_n1922_; 
wire w_mem_inst__abc_21203_new_n1923_; 
wire w_mem_inst__abc_21203_new_n1924_; 
wire w_mem_inst__abc_21203_new_n1925_; 
wire w_mem_inst__abc_21203_new_n1926_; 
wire w_mem_inst__abc_21203_new_n1927_; 
wire w_mem_inst__abc_21203_new_n1928_; 
wire w_mem_inst__abc_21203_new_n1929_; 
wire w_mem_inst__abc_21203_new_n1930_; 
wire w_mem_inst__abc_21203_new_n1931_; 
wire w_mem_inst__abc_21203_new_n1932_; 
wire w_mem_inst__abc_21203_new_n1933_; 
wire w_mem_inst__abc_21203_new_n1934_; 
wire w_mem_inst__abc_21203_new_n1935_; 
wire w_mem_inst__abc_21203_new_n1936_; 
wire w_mem_inst__abc_21203_new_n1937_; 
wire w_mem_inst__abc_21203_new_n1938_; 
wire w_mem_inst__abc_21203_new_n1939_; 
wire w_mem_inst__abc_21203_new_n1940_; 
wire w_mem_inst__abc_21203_new_n1941_; 
wire w_mem_inst__abc_21203_new_n1942_; 
wire w_mem_inst__abc_21203_new_n1943_; 
wire w_mem_inst__abc_21203_new_n1944_; 
wire w_mem_inst__abc_21203_new_n1945_; 
wire w_mem_inst__abc_21203_new_n1946_; 
wire w_mem_inst__abc_21203_new_n1947_; 
wire w_mem_inst__abc_21203_new_n1948_; 
wire w_mem_inst__abc_21203_new_n1949_; 
wire w_mem_inst__abc_21203_new_n1950_; 
wire w_mem_inst__abc_21203_new_n1952_; 
wire w_mem_inst__abc_21203_new_n1953_; 
wire w_mem_inst__abc_21203_new_n1954_; 
wire w_mem_inst__abc_21203_new_n1955_; 
wire w_mem_inst__abc_21203_new_n1956_; 
wire w_mem_inst__abc_21203_new_n1957_; 
wire w_mem_inst__abc_21203_new_n1958_; 
wire w_mem_inst__abc_21203_new_n1959_; 
wire w_mem_inst__abc_21203_new_n1960_; 
wire w_mem_inst__abc_21203_new_n1961_; 
wire w_mem_inst__abc_21203_new_n1962_; 
wire w_mem_inst__abc_21203_new_n1963_; 
wire w_mem_inst__abc_21203_new_n1964_; 
wire w_mem_inst__abc_21203_new_n1965_; 
wire w_mem_inst__abc_21203_new_n1966_; 
wire w_mem_inst__abc_21203_new_n1967_; 
wire w_mem_inst__abc_21203_new_n1968_; 
wire w_mem_inst__abc_21203_new_n1969_; 
wire w_mem_inst__abc_21203_new_n1970_; 
wire w_mem_inst__abc_21203_new_n1971_; 
wire w_mem_inst__abc_21203_new_n1972_; 
wire w_mem_inst__abc_21203_new_n1973_; 
wire w_mem_inst__abc_21203_new_n1974_; 
wire w_mem_inst__abc_21203_new_n1975_; 
wire w_mem_inst__abc_21203_new_n1976_; 
wire w_mem_inst__abc_21203_new_n1977_; 
wire w_mem_inst__abc_21203_new_n1978_; 
wire w_mem_inst__abc_21203_new_n1979_; 
wire w_mem_inst__abc_21203_new_n1980_; 
wire w_mem_inst__abc_21203_new_n1981_; 
wire w_mem_inst__abc_21203_new_n1982_; 
wire w_mem_inst__abc_21203_new_n1983_; 
wire w_mem_inst__abc_21203_new_n1984_; 
wire w_mem_inst__abc_21203_new_n1985_; 
wire w_mem_inst__abc_21203_new_n1986_; 
wire w_mem_inst__abc_21203_new_n1987_; 
wire w_mem_inst__abc_21203_new_n1988_; 
wire w_mem_inst__abc_21203_new_n1989_; 
wire w_mem_inst__abc_21203_new_n1990_; 
wire w_mem_inst__abc_21203_new_n1991_; 
wire w_mem_inst__abc_21203_new_n1992_; 
wire w_mem_inst__abc_21203_new_n1993_; 
wire w_mem_inst__abc_21203_new_n1994_; 
wire w_mem_inst__abc_21203_new_n1995_; 
wire w_mem_inst__abc_21203_new_n1996_; 
wire w_mem_inst__abc_21203_new_n1997_; 
wire w_mem_inst__abc_21203_new_n1998_; 
wire w_mem_inst__abc_21203_new_n2000_; 
wire w_mem_inst__abc_21203_new_n2001_; 
wire w_mem_inst__abc_21203_new_n2002_; 
wire w_mem_inst__abc_21203_new_n2003_; 
wire w_mem_inst__abc_21203_new_n2004_; 
wire w_mem_inst__abc_21203_new_n2005_; 
wire w_mem_inst__abc_21203_new_n2006_; 
wire w_mem_inst__abc_21203_new_n2007_; 
wire w_mem_inst__abc_21203_new_n2008_; 
wire w_mem_inst__abc_21203_new_n2009_; 
wire w_mem_inst__abc_21203_new_n2010_; 
wire w_mem_inst__abc_21203_new_n2011_; 
wire w_mem_inst__abc_21203_new_n2012_; 
wire w_mem_inst__abc_21203_new_n2013_; 
wire w_mem_inst__abc_21203_new_n2014_; 
wire w_mem_inst__abc_21203_new_n2015_; 
wire w_mem_inst__abc_21203_new_n2016_; 
wire w_mem_inst__abc_21203_new_n2017_; 
wire w_mem_inst__abc_21203_new_n2018_; 
wire w_mem_inst__abc_21203_new_n2019_; 
wire w_mem_inst__abc_21203_new_n2020_; 
wire w_mem_inst__abc_21203_new_n2021_; 
wire w_mem_inst__abc_21203_new_n2022_; 
wire w_mem_inst__abc_21203_new_n2023_; 
wire w_mem_inst__abc_21203_new_n2024_; 
wire w_mem_inst__abc_21203_new_n2025_; 
wire w_mem_inst__abc_21203_new_n2026_; 
wire w_mem_inst__abc_21203_new_n2027_; 
wire w_mem_inst__abc_21203_new_n2028_; 
wire w_mem_inst__abc_21203_new_n2029_; 
wire w_mem_inst__abc_21203_new_n2030_; 
wire w_mem_inst__abc_21203_new_n2031_; 
wire w_mem_inst__abc_21203_new_n2032_; 
wire w_mem_inst__abc_21203_new_n2033_; 
wire w_mem_inst__abc_21203_new_n2034_; 
wire w_mem_inst__abc_21203_new_n2035_; 
wire w_mem_inst__abc_21203_new_n2036_; 
wire w_mem_inst__abc_21203_new_n2037_; 
wire w_mem_inst__abc_21203_new_n2038_; 
wire w_mem_inst__abc_21203_new_n2039_; 
wire w_mem_inst__abc_21203_new_n2040_; 
wire w_mem_inst__abc_21203_new_n2041_; 
wire w_mem_inst__abc_21203_new_n2042_; 
wire w_mem_inst__abc_21203_new_n2043_; 
wire w_mem_inst__abc_21203_new_n2044_; 
wire w_mem_inst__abc_21203_new_n2045_; 
wire w_mem_inst__abc_21203_new_n2046_; 
wire w_mem_inst__abc_21203_new_n2048_; 
wire w_mem_inst__abc_21203_new_n2049_; 
wire w_mem_inst__abc_21203_new_n2050_; 
wire w_mem_inst__abc_21203_new_n2051_; 
wire w_mem_inst__abc_21203_new_n2052_; 
wire w_mem_inst__abc_21203_new_n2053_; 
wire w_mem_inst__abc_21203_new_n2054_; 
wire w_mem_inst__abc_21203_new_n2055_; 
wire w_mem_inst__abc_21203_new_n2056_; 
wire w_mem_inst__abc_21203_new_n2057_; 
wire w_mem_inst__abc_21203_new_n2058_; 
wire w_mem_inst__abc_21203_new_n2059_; 
wire w_mem_inst__abc_21203_new_n2060_; 
wire w_mem_inst__abc_21203_new_n2061_; 
wire w_mem_inst__abc_21203_new_n2062_; 
wire w_mem_inst__abc_21203_new_n2063_; 
wire w_mem_inst__abc_21203_new_n2064_; 
wire w_mem_inst__abc_21203_new_n2065_; 
wire w_mem_inst__abc_21203_new_n2066_; 
wire w_mem_inst__abc_21203_new_n2067_; 
wire w_mem_inst__abc_21203_new_n2068_; 
wire w_mem_inst__abc_21203_new_n2069_; 
wire w_mem_inst__abc_21203_new_n2070_; 
wire w_mem_inst__abc_21203_new_n2071_; 
wire w_mem_inst__abc_21203_new_n2072_; 
wire w_mem_inst__abc_21203_new_n2073_; 
wire w_mem_inst__abc_21203_new_n2074_; 
wire w_mem_inst__abc_21203_new_n2075_; 
wire w_mem_inst__abc_21203_new_n2076_; 
wire w_mem_inst__abc_21203_new_n2077_; 
wire w_mem_inst__abc_21203_new_n2078_; 
wire w_mem_inst__abc_21203_new_n2079_; 
wire w_mem_inst__abc_21203_new_n2080_; 
wire w_mem_inst__abc_21203_new_n2081_; 
wire w_mem_inst__abc_21203_new_n2082_; 
wire w_mem_inst__abc_21203_new_n2083_; 
wire w_mem_inst__abc_21203_new_n2084_; 
wire w_mem_inst__abc_21203_new_n2085_; 
wire w_mem_inst__abc_21203_new_n2086_; 
wire w_mem_inst__abc_21203_new_n2087_; 
wire w_mem_inst__abc_21203_new_n2088_; 
wire w_mem_inst__abc_21203_new_n2089_; 
wire w_mem_inst__abc_21203_new_n2090_; 
wire w_mem_inst__abc_21203_new_n2091_; 
wire w_mem_inst__abc_21203_new_n2092_; 
wire w_mem_inst__abc_21203_new_n2093_; 
wire w_mem_inst__abc_21203_new_n2094_; 
wire w_mem_inst__abc_21203_new_n2096_; 
wire w_mem_inst__abc_21203_new_n2097_; 
wire w_mem_inst__abc_21203_new_n2098_; 
wire w_mem_inst__abc_21203_new_n2099_; 
wire w_mem_inst__abc_21203_new_n2100_; 
wire w_mem_inst__abc_21203_new_n2101_; 
wire w_mem_inst__abc_21203_new_n2102_; 
wire w_mem_inst__abc_21203_new_n2103_; 
wire w_mem_inst__abc_21203_new_n2104_; 
wire w_mem_inst__abc_21203_new_n2105_; 
wire w_mem_inst__abc_21203_new_n2106_; 
wire w_mem_inst__abc_21203_new_n2107_; 
wire w_mem_inst__abc_21203_new_n2108_; 
wire w_mem_inst__abc_21203_new_n2109_; 
wire w_mem_inst__abc_21203_new_n2110_; 
wire w_mem_inst__abc_21203_new_n2111_; 
wire w_mem_inst__abc_21203_new_n2112_; 
wire w_mem_inst__abc_21203_new_n2113_; 
wire w_mem_inst__abc_21203_new_n2114_; 
wire w_mem_inst__abc_21203_new_n2115_; 
wire w_mem_inst__abc_21203_new_n2116_; 
wire w_mem_inst__abc_21203_new_n2117_; 
wire w_mem_inst__abc_21203_new_n2118_; 
wire w_mem_inst__abc_21203_new_n2119_; 
wire w_mem_inst__abc_21203_new_n2120_; 
wire w_mem_inst__abc_21203_new_n2121_; 
wire w_mem_inst__abc_21203_new_n2122_; 
wire w_mem_inst__abc_21203_new_n2123_; 
wire w_mem_inst__abc_21203_new_n2124_; 
wire w_mem_inst__abc_21203_new_n2125_; 
wire w_mem_inst__abc_21203_new_n2126_; 
wire w_mem_inst__abc_21203_new_n2127_; 
wire w_mem_inst__abc_21203_new_n2128_; 
wire w_mem_inst__abc_21203_new_n2129_; 
wire w_mem_inst__abc_21203_new_n2130_; 
wire w_mem_inst__abc_21203_new_n2131_; 
wire w_mem_inst__abc_21203_new_n2132_; 
wire w_mem_inst__abc_21203_new_n2133_; 
wire w_mem_inst__abc_21203_new_n2134_; 
wire w_mem_inst__abc_21203_new_n2135_; 
wire w_mem_inst__abc_21203_new_n2136_; 
wire w_mem_inst__abc_21203_new_n2137_; 
wire w_mem_inst__abc_21203_new_n2138_; 
wire w_mem_inst__abc_21203_new_n2139_; 
wire w_mem_inst__abc_21203_new_n2140_; 
wire w_mem_inst__abc_21203_new_n2141_; 
wire w_mem_inst__abc_21203_new_n2142_; 
wire w_mem_inst__abc_21203_new_n2144_; 
wire w_mem_inst__abc_21203_new_n2145_; 
wire w_mem_inst__abc_21203_new_n2146_; 
wire w_mem_inst__abc_21203_new_n2147_; 
wire w_mem_inst__abc_21203_new_n2148_; 
wire w_mem_inst__abc_21203_new_n2149_; 
wire w_mem_inst__abc_21203_new_n2150_; 
wire w_mem_inst__abc_21203_new_n2151_; 
wire w_mem_inst__abc_21203_new_n2152_; 
wire w_mem_inst__abc_21203_new_n2153_; 
wire w_mem_inst__abc_21203_new_n2154_; 
wire w_mem_inst__abc_21203_new_n2155_; 
wire w_mem_inst__abc_21203_new_n2156_; 
wire w_mem_inst__abc_21203_new_n2157_; 
wire w_mem_inst__abc_21203_new_n2158_; 
wire w_mem_inst__abc_21203_new_n2159_; 
wire w_mem_inst__abc_21203_new_n2160_; 
wire w_mem_inst__abc_21203_new_n2161_; 
wire w_mem_inst__abc_21203_new_n2162_; 
wire w_mem_inst__abc_21203_new_n2163_; 
wire w_mem_inst__abc_21203_new_n2164_; 
wire w_mem_inst__abc_21203_new_n2165_; 
wire w_mem_inst__abc_21203_new_n2166_; 
wire w_mem_inst__abc_21203_new_n2167_; 
wire w_mem_inst__abc_21203_new_n2168_; 
wire w_mem_inst__abc_21203_new_n2169_; 
wire w_mem_inst__abc_21203_new_n2170_; 
wire w_mem_inst__abc_21203_new_n2171_; 
wire w_mem_inst__abc_21203_new_n2172_; 
wire w_mem_inst__abc_21203_new_n2173_; 
wire w_mem_inst__abc_21203_new_n2174_; 
wire w_mem_inst__abc_21203_new_n2175_; 
wire w_mem_inst__abc_21203_new_n2176_; 
wire w_mem_inst__abc_21203_new_n2177_; 
wire w_mem_inst__abc_21203_new_n2178_; 
wire w_mem_inst__abc_21203_new_n2179_; 
wire w_mem_inst__abc_21203_new_n2180_; 
wire w_mem_inst__abc_21203_new_n2181_; 
wire w_mem_inst__abc_21203_new_n2182_; 
wire w_mem_inst__abc_21203_new_n2183_; 
wire w_mem_inst__abc_21203_new_n2184_; 
wire w_mem_inst__abc_21203_new_n2185_; 
wire w_mem_inst__abc_21203_new_n2186_; 
wire w_mem_inst__abc_21203_new_n2187_; 
wire w_mem_inst__abc_21203_new_n2188_; 
wire w_mem_inst__abc_21203_new_n2189_; 
wire w_mem_inst__abc_21203_new_n2190_; 
wire w_mem_inst__abc_21203_new_n2192_; 
wire w_mem_inst__abc_21203_new_n2193_; 
wire w_mem_inst__abc_21203_new_n2194_; 
wire w_mem_inst__abc_21203_new_n2195_; 
wire w_mem_inst__abc_21203_new_n2196_; 
wire w_mem_inst__abc_21203_new_n2197_; 
wire w_mem_inst__abc_21203_new_n2198_; 
wire w_mem_inst__abc_21203_new_n2199_; 
wire w_mem_inst__abc_21203_new_n2200_; 
wire w_mem_inst__abc_21203_new_n2201_; 
wire w_mem_inst__abc_21203_new_n2202_; 
wire w_mem_inst__abc_21203_new_n2203_; 
wire w_mem_inst__abc_21203_new_n2204_; 
wire w_mem_inst__abc_21203_new_n2205_; 
wire w_mem_inst__abc_21203_new_n2206_; 
wire w_mem_inst__abc_21203_new_n2207_; 
wire w_mem_inst__abc_21203_new_n2208_; 
wire w_mem_inst__abc_21203_new_n2209_; 
wire w_mem_inst__abc_21203_new_n2210_; 
wire w_mem_inst__abc_21203_new_n2211_; 
wire w_mem_inst__abc_21203_new_n2212_; 
wire w_mem_inst__abc_21203_new_n2213_; 
wire w_mem_inst__abc_21203_new_n2214_; 
wire w_mem_inst__abc_21203_new_n2215_; 
wire w_mem_inst__abc_21203_new_n2216_; 
wire w_mem_inst__abc_21203_new_n2217_; 
wire w_mem_inst__abc_21203_new_n2218_; 
wire w_mem_inst__abc_21203_new_n2219_; 
wire w_mem_inst__abc_21203_new_n2220_; 
wire w_mem_inst__abc_21203_new_n2221_; 
wire w_mem_inst__abc_21203_new_n2222_; 
wire w_mem_inst__abc_21203_new_n2223_; 
wire w_mem_inst__abc_21203_new_n2224_; 
wire w_mem_inst__abc_21203_new_n2225_; 
wire w_mem_inst__abc_21203_new_n2226_; 
wire w_mem_inst__abc_21203_new_n2227_; 
wire w_mem_inst__abc_21203_new_n2228_; 
wire w_mem_inst__abc_21203_new_n2229_; 
wire w_mem_inst__abc_21203_new_n2230_; 
wire w_mem_inst__abc_21203_new_n2231_; 
wire w_mem_inst__abc_21203_new_n2232_; 
wire w_mem_inst__abc_21203_new_n2233_; 
wire w_mem_inst__abc_21203_new_n2234_; 
wire w_mem_inst__abc_21203_new_n2235_; 
wire w_mem_inst__abc_21203_new_n2236_; 
wire w_mem_inst__abc_21203_new_n2237_; 
wire w_mem_inst__abc_21203_new_n2238_; 
wire w_mem_inst__abc_21203_new_n2240_; 
wire w_mem_inst__abc_21203_new_n2241_; 
wire w_mem_inst__abc_21203_new_n2242_; 
wire w_mem_inst__abc_21203_new_n2243_; 
wire w_mem_inst__abc_21203_new_n2244_; 
wire w_mem_inst__abc_21203_new_n2245_; 
wire w_mem_inst__abc_21203_new_n2246_; 
wire w_mem_inst__abc_21203_new_n2247_; 
wire w_mem_inst__abc_21203_new_n2248_; 
wire w_mem_inst__abc_21203_new_n2249_; 
wire w_mem_inst__abc_21203_new_n2250_; 
wire w_mem_inst__abc_21203_new_n2251_; 
wire w_mem_inst__abc_21203_new_n2252_; 
wire w_mem_inst__abc_21203_new_n2253_; 
wire w_mem_inst__abc_21203_new_n2254_; 
wire w_mem_inst__abc_21203_new_n2255_; 
wire w_mem_inst__abc_21203_new_n2256_; 
wire w_mem_inst__abc_21203_new_n2257_; 
wire w_mem_inst__abc_21203_new_n2258_; 
wire w_mem_inst__abc_21203_new_n2259_; 
wire w_mem_inst__abc_21203_new_n2260_; 
wire w_mem_inst__abc_21203_new_n2261_; 
wire w_mem_inst__abc_21203_new_n2262_; 
wire w_mem_inst__abc_21203_new_n2263_; 
wire w_mem_inst__abc_21203_new_n2264_; 
wire w_mem_inst__abc_21203_new_n2265_; 
wire w_mem_inst__abc_21203_new_n2266_; 
wire w_mem_inst__abc_21203_new_n2267_; 
wire w_mem_inst__abc_21203_new_n2268_; 
wire w_mem_inst__abc_21203_new_n2269_; 
wire w_mem_inst__abc_21203_new_n2270_; 
wire w_mem_inst__abc_21203_new_n2271_; 
wire w_mem_inst__abc_21203_new_n2272_; 
wire w_mem_inst__abc_21203_new_n2273_; 
wire w_mem_inst__abc_21203_new_n2274_; 
wire w_mem_inst__abc_21203_new_n2275_; 
wire w_mem_inst__abc_21203_new_n2276_; 
wire w_mem_inst__abc_21203_new_n2277_; 
wire w_mem_inst__abc_21203_new_n2278_; 
wire w_mem_inst__abc_21203_new_n2279_; 
wire w_mem_inst__abc_21203_new_n2280_; 
wire w_mem_inst__abc_21203_new_n2281_; 
wire w_mem_inst__abc_21203_new_n2282_; 
wire w_mem_inst__abc_21203_new_n2283_; 
wire w_mem_inst__abc_21203_new_n2284_; 
wire w_mem_inst__abc_21203_new_n2285_; 
wire w_mem_inst__abc_21203_new_n2286_; 
wire w_mem_inst__abc_21203_new_n2288_; 
wire w_mem_inst__abc_21203_new_n2289_; 
wire w_mem_inst__abc_21203_new_n2290_; 
wire w_mem_inst__abc_21203_new_n2291_; 
wire w_mem_inst__abc_21203_new_n2292_; 
wire w_mem_inst__abc_21203_new_n2293_; 
wire w_mem_inst__abc_21203_new_n2294_; 
wire w_mem_inst__abc_21203_new_n2295_; 
wire w_mem_inst__abc_21203_new_n2296_; 
wire w_mem_inst__abc_21203_new_n2297_; 
wire w_mem_inst__abc_21203_new_n2298_; 
wire w_mem_inst__abc_21203_new_n2299_; 
wire w_mem_inst__abc_21203_new_n2300_; 
wire w_mem_inst__abc_21203_new_n2301_; 
wire w_mem_inst__abc_21203_new_n2302_; 
wire w_mem_inst__abc_21203_new_n2303_; 
wire w_mem_inst__abc_21203_new_n2304_; 
wire w_mem_inst__abc_21203_new_n2305_; 
wire w_mem_inst__abc_21203_new_n2306_; 
wire w_mem_inst__abc_21203_new_n2307_; 
wire w_mem_inst__abc_21203_new_n2308_; 
wire w_mem_inst__abc_21203_new_n2309_; 
wire w_mem_inst__abc_21203_new_n2310_; 
wire w_mem_inst__abc_21203_new_n2311_; 
wire w_mem_inst__abc_21203_new_n2312_; 
wire w_mem_inst__abc_21203_new_n2313_; 
wire w_mem_inst__abc_21203_new_n2314_; 
wire w_mem_inst__abc_21203_new_n2315_; 
wire w_mem_inst__abc_21203_new_n2316_; 
wire w_mem_inst__abc_21203_new_n2317_; 
wire w_mem_inst__abc_21203_new_n2318_; 
wire w_mem_inst__abc_21203_new_n2319_; 
wire w_mem_inst__abc_21203_new_n2320_; 
wire w_mem_inst__abc_21203_new_n2321_; 
wire w_mem_inst__abc_21203_new_n2322_; 
wire w_mem_inst__abc_21203_new_n2323_; 
wire w_mem_inst__abc_21203_new_n2324_; 
wire w_mem_inst__abc_21203_new_n2325_; 
wire w_mem_inst__abc_21203_new_n2326_; 
wire w_mem_inst__abc_21203_new_n2327_; 
wire w_mem_inst__abc_21203_new_n2328_; 
wire w_mem_inst__abc_21203_new_n2329_; 
wire w_mem_inst__abc_21203_new_n2330_; 
wire w_mem_inst__abc_21203_new_n2331_; 
wire w_mem_inst__abc_21203_new_n2332_; 
wire w_mem_inst__abc_21203_new_n2333_; 
wire w_mem_inst__abc_21203_new_n2334_; 
wire w_mem_inst__abc_21203_new_n2336_; 
wire w_mem_inst__abc_21203_new_n2337_; 
wire w_mem_inst__abc_21203_new_n2338_; 
wire w_mem_inst__abc_21203_new_n2339_; 
wire w_mem_inst__abc_21203_new_n2340_; 
wire w_mem_inst__abc_21203_new_n2341_; 
wire w_mem_inst__abc_21203_new_n2342_; 
wire w_mem_inst__abc_21203_new_n2343_; 
wire w_mem_inst__abc_21203_new_n2344_; 
wire w_mem_inst__abc_21203_new_n2345_; 
wire w_mem_inst__abc_21203_new_n2346_; 
wire w_mem_inst__abc_21203_new_n2347_; 
wire w_mem_inst__abc_21203_new_n2348_; 
wire w_mem_inst__abc_21203_new_n2349_; 
wire w_mem_inst__abc_21203_new_n2350_; 
wire w_mem_inst__abc_21203_new_n2351_; 
wire w_mem_inst__abc_21203_new_n2352_; 
wire w_mem_inst__abc_21203_new_n2353_; 
wire w_mem_inst__abc_21203_new_n2354_; 
wire w_mem_inst__abc_21203_new_n2355_; 
wire w_mem_inst__abc_21203_new_n2356_; 
wire w_mem_inst__abc_21203_new_n2357_; 
wire w_mem_inst__abc_21203_new_n2358_; 
wire w_mem_inst__abc_21203_new_n2359_; 
wire w_mem_inst__abc_21203_new_n2360_; 
wire w_mem_inst__abc_21203_new_n2361_; 
wire w_mem_inst__abc_21203_new_n2362_; 
wire w_mem_inst__abc_21203_new_n2363_; 
wire w_mem_inst__abc_21203_new_n2364_; 
wire w_mem_inst__abc_21203_new_n2365_; 
wire w_mem_inst__abc_21203_new_n2366_; 
wire w_mem_inst__abc_21203_new_n2367_; 
wire w_mem_inst__abc_21203_new_n2368_; 
wire w_mem_inst__abc_21203_new_n2369_; 
wire w_mem_inst__abc_21203_new_n2370_; 
wire w_mem_inst__abc_21203_new_n2371_; 
wire w_mem_inst__abc_21203_new_n2372_; 
wire w_mem_inst__abc_21203_new_n2373_; 
wire w_mem_inst__abc_21203_new_n2374_; 
wire w_mem_inst__abc_21203_new_n2375_; 
wire w_mem_inst__abc_21203_new_n2376_; 
wire w_mem_inst__abc_21203_new_n2377_; 
wire w_mem_inst__abc_21203_new_n2378_; 
wire w_mem_inst__abc_21203_new_n2379_; 
wire w_mem_inst__abc_21203_new_n2380_; 
wire w_mem_inst__abc_21203_new_n2381_; 
wire w_mem_inst__abc_21203_new_n2382_; 
wire w_mem_inst__abc_21203_new_n2384_; 
wire w_mem_inst__abc_21203_new_n2385_; 
wire w_mem_inst__abc_21203_new_n2386_; 
wire w_mem_inst__abc_21203_new_n2387_; 
wire w_mem_inst__abc_21203_new_n2388_; 
wire w_mem_inst__abc_21203_new_n2389_; 
wire w_mem_inst__abc_21203_new_n2390_; 
wire w_mem_inst__abc_21203_new_n2391_; 
wire w_mem_inst__abc_21203_new_n2392_; 
wire w_mem_inst__abc_21203_new_n2393_; 
wire w_mem_inst__abc_21203_new_n2394_; 
wire w_mem_inst__abc_21203_new_n2395_; 
wire w_mem_inst__abc_21203_new_n2396_; 
wire w_mem_inst__abc_21203_new_n2397_; 
wire w_mem_inst__abc_21203_new_n2398_; 
wire w_mem_inst__abc_21203_new_n2399_; 
wire w_mem_inst__abc_21203_new_n2400_; 
wire w_mem_inst__abc_21203_new_n2401_; 
wire w_mem_inst__abc_21203_new_n2402_; 
wire w_mem_inst__abc_21203_new_n2403_; 
wire w_mem_inst__abc_21203_new_n2404_; 
wire w_mem_inst__abc_21203_new_n2405_; 
wire w_mem_inst__abc_21203_new_n2406_; 
wire w_mem_inst__abc_21203_new_n2407_; 
wire w_mem_inst__abc_21203_new_n2408_; 
wire w_mem_inst__abc_21203_new_n2409_; 
wire w_mem_inst__abc_21203_new_n2410_; 
wire w_mem_inst__abc_21203_new_n2411_; 
wire w_mem_inst__abc_21203_new_n2412_; 
wire w_mem_inst__abc_21203_new_n2413_; 
wire w_mem_inst__abc_21203_new_n2414_; 
wire w_mem_inst__abc_21203_new_n2415_; 
wire w_mem_inst__abc_21203_new_n2416_; 
wire w_mem_inst__abc_21203_new_n2417_; 
wire w_mem_inst__abc_21203_new_n2418_; 
wire w_mem_inst__abc_21203_new_n2419_; 
wire w_mem_inst__abc_21203_new_n2420_; 
wire w_mem_inst__abc_21203_new_n2421_; 
wire w_mem_inst__abc_21203_new_n2422_; 
wire w_mem_inst__abc_21203_new_n2423_; 
wire w_mem_inst__abc_21203_new_n2424_; 
wire w_mem_inst__abc_21203_new_n2425_; 
wire w_mem_inst__abc_21203_new_n2426_; 
wire w_mem_inst__abc_21203_new_n2427_; 
wire w_mem_inst__abc_21203_new_n2428_; 
wire w_mem_inst__abc_21203_new_n2429_; 
wire w_mem_inst__abc_21203_new_n2430_; 
wire w_mem_inst__abc_21203_new_n2432_; 
wire w_mem_inst__abc_21203_new_n2433_; 
wire w_mem_inst__abc_21203_new_n2434_; 
wire w_mem_inst__abc_21203_new_n2435_; 
wire w_mem_inst__abc_21203_new_n2436_; 
wire w_mem_inst__abc_21203_new_n2437_; 
wire w_mem_inst__abc_21203_new_n2438_; 
wire w_mem_inst__abc_21203_new_n2439_; 
wire w_mem_inst__abc_21203_new_n2440_; 
wire w_mem_inst__abc_21203_new_n2441_; 
wire w_mem_inst__abc_21203_new_n2442_; 
wire w_mem_inst__abc_21203_new_n2443_; 
wire w_mem_inst__abc_21203_new_n2444_; 
wire w_mem_inst__abc_21203_new_n2445_; 
wire w_mem_inst__abc_21203_new_n2446_; 
wire w_mem_inst__abc_21203_new_n2447_; 
wire w_mem_inst__abc_21203_new_n2448_; 
wire w_mem_inst__abc_21203_new_n2449_; 
wire w_mem_inst__abc_21203_new_n2450_; 
wire w_mem_inst__abc_21203_new_n2451_; 
wire w_mem_inst__abc_21203_new_n2452_; 
wire w_mem_inst__abc_21203_new_n2453_; 
wire w_mem_inst__abc_21203_new_n2454_; 
wire w_mem_inst__abc_21203_new_n2455_; 
wire w_mem_inst__abc_21203_new_n2456_; 
wire w_mem_inst__abc_21203_new_n2457_; 
wire w_mem_inst__abc_21203_new_n2458_; 
wire w_mem_inst__abc_21203_new_n2459_; 
wire w_mem_inst__abc_21203_new_n2460_; 
wire w_mem_inst__abc_21203_new_n2461_; 
wire w_mem_inst__abc_21203_new_n2462_; 
wire w_mem_inst__abc_21203_new_n2463_; 
wire w_mem_inst__abc_21203_new_n2464_; 
wire w_mem_inst__abc_21203_new_n2465_; 
wire w_mem_inst__abc_21203_new_n2466_; 
wire w_mem_inst__abc_21203_new_n2467_; 
wire w_mem_inst__abc_21203_new_n2468_; 
wire w_mem_inst__abc_21203_new_n2469_; 
wire w_mem_inst__abc_21203_new_n2470_; 
wire w_mem_inst__abc_21203_new_n2471_; 
wire w_mem_inst__abc_21203_new_n2472_; 
wire w_mem_inst__abc_21203_new_n2473_; 
wire w_mem_inst__abc_21203_new_n2474_; 
wire w_mem_inst__abc_21203_new_n2475_; 
wire w_mem_inst__abc_21203_new_n2476_; 
wire w_mem_inst__abc_21203_new_n2477_; 
wire w_mem_inst__abc_21203_new_n2478_; 
wire w_mem_inst__abc_21203_new_n2480_; 
wire w_mem_inst__abc_21203_new_n2481_; 
wire w_mem_inst__abc_21203_new_n2482_; 
wire w_mem_inst__abc_21203_new_n2483_; 
wire w_mem_inst__abc_21203_new_n2484_; 
wire w_mem_inst__abc_21203_new_n2485_; 
wire w_mem_inst__abc_21203_new_n2486_; 
wire w_mem_inst__abc_21203_new_n2487_; 
wire w_mem_inst__abc_21203_new_n2488_; 
wire w_mem_inst__abc_21203_new_n2489_; 
wire w_mem_inst__abc_21203_new_n2490_; 
wire w_mem_inst__abc_21203_new_n2491_; 
wire w_mem_inst__abc_21203_new_n2492_; 
wire w_mem_inst__abc_21203_new_n2493_; 
wire w_mem_inst__abc_21203_new_n2494_; 
wire w_mem_inst__abc_21203_new_n2495_; 
wire w_mem_inst__abc_21203_new_n2496_; 
wire w_mem_inst__abc_21203_new_n2497_; 
wire w_mem_inst__abc_21203_new_n2498_; 
wire w_mem_inst__abc_21203_new_n2499_; 
wire w_mem_inst__abc_21203_new_n2500_; 
wire w_mem_inst__abc_21203_new_n2501_; 
wire w_mem_inst__abc_21203_new_n2502_; 
wire w_mem_inst__abc_21203_new_n2503_; 
wire w_mem_inst__abc_21203_new_n2504_; 
wire w_mem_inst__abc_21203_new_n2505_; 
wire w_mem_inst__abc_21203_new_n2506_; 
wire w_mem_inst__abc_21203_new_n2507_; 
wire w_mem_inst__abc_21203_new_n2508_; 
wire w_mem_inst__abc_21203_new_n2509_; 
wire w_mem_inst__abc_21203_new_n2510_; 
wire w_mem_inst__abc_21203_new_n2511_; 
wire w_mem_inst__abc_21203_new_n2512_; 
wire w_mem_inst__abc_21203_new_n2513_; 
wire w_mem_inst__abc_21203_new_n2514_; 
wire w_mem_inst__abc_21203_new_n2515_; 
wire w_mem_inst__abc_21203_new_n2516_; 
wire w_mem_inst__abc_21203_new_n2517_; 
wire w_mem_inst__abc_21203_new_n2518_; 
wire w_mem_inst__abc_21203_new_n2519_; 
wire w_mem_inst__abc_21203_new_n2520_; 
wire w_mem_inst__abc_21203_new_n2521_; 
wire w_mem_inst__abc_21203_new_n2522_; 
wire w_mem_inst__abc_21203_new_n2523_; 
wire w_mem_inst__abc_21203_new_n2524_; 
wire w_mem_inst__abc_21203_new_n2525_; 
wire w_mem_inst__abc_21203_new_n2526_; 
wire w_mem_inst__abc_21203_new_n2528_; 
wire w_mem_inst__abc_21203_new_n2529_; 
wire w_mem_inst__abc_21203_new_n2530_; 
wire w_mem_inst__abc_21203_new_n2531_; 
wire w_mem_inst__abc_21203_new_n2532_; 
wire w_mem_inst__abc_21203_new_n2533_; 
wire w_mem_inst__abc_21203_new_n2534_; 
wire w_mem_inst__abc_21203_new_n2535_; 
wire w_mem_inst__abc_21203_new_n2536_; 
wire w_mem_inst__abc_21203_new_n2537_; 
wire w_mem_inst__abc_21203_new_n2538_; 
wire w_mem_inst__abc_21203_new_n2539_; 
wire w_mem_inst__abc_21203_new_n2540_; 
wire w_mem_inst__abc_21203_new_n2541_; 
wire w_mem_inst__abc_21203_new_n2542_; 
wire w_mem_inst__abc_21203_new_n2543_; 
wire w_mem_inst__abc_21203_new_n2544_; 
wire w_mem_inst__abc_21203_new_n2545_; 
wire w_mem_inst__abc_21203_new_n2546_; 
wire w_mem_inst__abc_21203_new_n2547_; 
wire w_mem_inst__abc_21203_new_n2548_; 
wire w_mem_inst__abc_21203_new_n2549_; 
wire w_mem_inst__abc_21203_new_n2550_; 
wire w_mem_inst__abc_21203_new_n2551_; 
wire w_mem_inst__abc_21203_new_n2552_; 
wire w_mem_inst__abc_21203_new_n2553_; 
wire w_mem_inst__abc_21203_new_n2554_; 
wire w_mem_inst__abc_21203_new_n2555_; 
wire w_mem_inst__abc_21203_new_n2556_; 
wire w_mem_inst__abc_21203_new_n2557_; 
wire w_mem_inst__abc_21203_new_n2558_; 
wire w_mem_inst__abc_21203_new_n2559_; 
wire w_mem_inst__abc_21203_new_n2560_; 
wire w_mem_inst__abc_21203_new_n2561_; 
wire w_mem_inst__abc_21203_new_n2562_; 
wire w_mem_inst__abc_21203_new_n2563_; 
wire w_mem_inst__abc_21203_new_n2564_; 
wire w_mem_inst__abc_21203_new_n2565_; 
wire w_mem_inst__abc_21203_new_n2566_; 
wire w_mem_inst__abc_21203_new_n2567_; 
wire w_mem_inst__abc_21203_new_n2568_; 
wire w_mem_inst__abc_21203_new_n2569_; 
wire w_mem_inst__abc_21203_new_n2570_; 
wire w_mem_inst__abc_21203_new_n2571_; 
wire w_mem_inst__abc_21203_new_n2572_; 
wire w_mem_inst__abc_21203_new_n2573_; 
wire w_mem_inst__abc_21203_new_n2574_; 
wire w_mem_inst__abc_21203_new_n2576_; 
wire w_mem_inst__abc_21203_new_n2577_; 
wire w_mem_inst__abc_21203_new_n2578_; 
wire w_mem_inst__abc_21203_new_n2579_; 
wire w_mem_inst__abc_21203_new_n2580_; 
wire w_mem_inst__abc_21203_new_n2581_; 
wire w_mem_inst__abc_21203_new_n2582_; 
wire w_mem_inst__abc_21203_new_n2583_; 
wire w_mem_inst__abc_21203_new_n2584_; 
wire w_mem_inst__abc_21203_new_n2585_; 
wire w_mem_inst__abc_21203_new_n2586_; 
wire w_mem_inst__abc_21203_new_n2587_; 
wire w_mem_inst__abc_21203_new_n2588_; 
wire w_mem_inst__abc_21203_new_n2589_; 
wire w_mem_inst__abc_21203_new_n2590_; 
wire w_mem_inst__abc_21203_new_n2591_; 
wire w_mem_inst__abc_21203_new_n2592_; 
wire w_mem_inst__abc_21203_new_n2593_; 
wire w_mem_inst__abc_21203_new_n2594_; 
wire w_mem_inst__abc_21203_new_n2595_; 
wire w_mem_inst__abc_21203_new_n2596_; 
wire w_mem_inst__abc_21203_new_n2597_; 
wire w_mem_inst__abc_21203_new_n2598_; 
wire w_mem_inst__abc_21203_new_n2599_; 
wire w_mem_inst__abc_21203_new_n2600_; 
wire w_mem_inst__abc_21203_new_n2601_; 
wire w_mem_inst__abc_21203_new_n2602_; 
wire w_mem_inst__abc_21203_new_n2603_; 
wire w_mem_inst__abc_21203_new_n2604_; 
wire w_mem_inst__abc_21203_new_n2605_; 
wire w_mem_inst__abc_21203_new_n2606_; 
wire w_mem_inst__abc_21203_new_n2607_; 
wire w_mem_inst__abc_21203_new_n2608_; 
wire w_mem_inst__abc_21203_new_n2609_; 
wire w_mem_inst__abc_21203_new_n2610_; 
wire w_mem_inst__abc_21203_new_n2611_; 
wire w_mem_inst__abc_21203_new_n2612_; 
wire w_mem_inst__abc_21203_new_n2613_; 
wire w_mem_inst__abc_21203_new_n2614_; 
wire w_mem_inst__abc_21203_new_n2615_; 
wire w_mem_inst__abc_21203_new_n2616_; 
wire w_mem_inst__abc_21203_new_n2617_; 
wire w_mem_inst__abc_21203_new_n2618_; 
wire w_mem_inst__abc_21203_new_n2619_; 
wire w_mem_inst__abc_21203_new_n2620_; 
wire w_mem_inst__abc_21203_new_n2621_; 
wire w_mem_inst__abc_21203_new_n2622_; 
wire w_mem_inst__abc_21203_new_n2624_; 
wire w_mem_inst__abc_21203_new_n2625_; 
wire w_mem_inst__abc_21203_new_n2626_; 
wire w_mem_inst__abc_21203_new_n2627_; 
wire w_mem_inst__abc_21203_new_n2628_; 
wire w_mem_inst__abc_21203_new_n2629_; 
wire w_mem_inst__abc_21203_new_n2630_; 
wire w_mem_inst__abc_21203_new_n2631_; 
wire w_mem_inst__abc_21203_new_n2632_; 
wire w_mem_inst__abc_21203_new_n2633_; 
wire w_mem_inst__abc_21203_new_n2634_; 
wire w_mem_inst__abc_21203_new_n2635_; 
wire w_mem_inst__abc_21203_new_n2636_; 
wire w_mem_inst__abc_21203_new_n2637_; 
wire w_mem_inst__abc_21203_new_n2638_; 
wire w_mem_inst__abc_21203_new_n2639_; 
wire w_mem_inst__abc_21203_new_n2640_; 
wire w_mem_inst__abc_21203_new_n2641_; 
wire w_mem_inst__abc_21203_new_n2642_; 
wire w_mem_inst__abc_21203_new_n2643_; 
wire w_mem_inst__abc_21203_new_n2644_; 
wire w_mem_inst__abc_21203_new_n2645_; 
wire w_mem_inst__abc_21203_new_n2646_; 
wire w_mem_inst__abc_21203_new_n2647_; 
wire w_mem_inst__abc_21203_new_n2648_; 
wire w_mem_inst__abc_21203_new_n2649_; 
wire w_mem_inst__abc_21203_new_n2650_; 
wire w_mem_inst__abc_21203_new_n2651_; 
wire w_mem_inst__abc_21203_new_n2652_; 
wire w_mem_inst__abc_21203_new_n2653_; 
wire w_mem_inst__abc_21203_new_n2654_; 
wire w_mem_inst__abc_21203_new_n2655_; 
wire w_mem_inst__abc_21203_new_n2656_; 
wire w_mem_inst__abc_21203_new_n2657_; 
wire w_mem_inst__abc_21203_new_n2658_; 
wire w_mem_inst__abc_21203_new_n2659_; 
wire w_mem_inst__abc_21203_new_n2660_; 
wire w_mem_inst__abc_21203_new_n2661_; 
wire w_mem_inst__abc_21203_new_n2662_; 
wire w_mem_inst__abc_21203_new_n2663_; 
wire w_mem_inst__abc_21203_new_n2664_; 
wire w_mem_inst__abc_21203_new_n2665_; 
wire w_mem_inst__abc_21203_new_n2666_; 
wire w_mem_inst__abc_21203_new_n2667_; 
wire w_mem_inst__abc_21203_new_n2668_; 
wire w_mem_inst__abc_21203_new_n2669_; 
wire w_mem_inst__abc_21203_new_n2670_; 
wire w_mem_inst__abc_21203_new_n2672_; 
wire w_mem_inst__abc_21203_new_n2673_; 
wire w_mem_inst__abc_21203_new_n2674_; 
wire w_mem_inst__abc_21203_new_n2675_; 
wire w_mem_inst__abc_21203_new_n2676_; 
wire w_mem_inst__abc_21203_new_n2677_; 
wire w_mem_inst__abc_21203_new_n2678_; 
wire w_mem_inst__abc_21203_new_n2679_; 
wire w_mem_inst__abc_21203_new_n2680_; 
wire w_mem_inst__abc_21203_new_n2681_; 
wire w_mem_inst__abc_21203_new_n2682_; 
wire w_mem_inst__abc_21203_new_n2683_; 
wire w_mem_inst__abc_21203_new_n2684_; 
wire w_mem_inst__abc_21203_new_n2685_; 
wire w_mem_inst__abc_21203_new_n2686_; 
wire w_mem_inst__abc_21203_new_n2687_; 
wire w_mem_inst__abc_21203_new_n2688_; 
wire w_mem_inst__abc_21203_new_n2689_; 
wire w_mem_inst__abc_21203_new_n2690_; 
wire w_mem_inst__abc_21203_new_n2691_; 
wire w_mem_inst__abc_21203_new_n2692_; 
wire w_mem_inst__abc_21203_new_n2693_; 
wire w_mem_inst__abc_21203_new_n2694_; 
wire w_mem_inst__abc_21203_new_n2695_; 
wire w_mem_inst__abc_21203_new_n2696_; 
wire w_mem_inst__abc_21203_new_n2697_; 
wire w_mem_inst__abc_21203_new_n2698_; 
wire w_mem_inst__abc_21203_new_n2699_; 
wire w_mem_inst__abc_21203_new_n2700_; 
wire w_mem_inst__abc_21203_new_n2701_; 
wire w_mem_inst__abc_21203_new_n2702_; 
wire w_mem_inst__abc_21203_new_n2703_; 
wire w_mem_inst__abc_21203_new_n2704_; 
wire w_mem_inst__abc_21203_new_n2705_; 
wire w_mem_inst__abc_21203_new_n2706_; 
wire w_mem_inst__abc_21203_new_n2707_; 
wire w_mem_inst__abc_21203_new_n2708_; 
wire w_mem_inst__abc_21203_new_n2709_; 
wire w_mem_inst__abc_21203_new_n2710_; 
wire w_mem_inst__abc_21203_new_n2711_; 
wire w_mem_inst__abc_21203_new_n2712_; 
wire w_mem_inst__abc_21203_new_n2713_; 
wire w_mem_inst__abc_21203_new_n2714_; 
wire w_mem_inst__abc_21203_new_n2715_; 
wire w_mem_inst__abc_21203_new_n2716_; 
wire w_mem_inst__abc_21203_new_n2717_; 
wire w_mem_inst__abc_21203_new_n2718_; 
wire w_mem_inst__abc_21203_new_n2720_; 
wire w_mem_inst__abc_21203_new_n2721_; 
wire w_mem_inst__abc_21203_new_n2722_; 
wire w_mem_inst__abc_21203_new_n2723_; 
wire w_mem_inst__abc_21203_new_n2724_; 
wire w_mem_inst__abc_21203_new_n2725_; 
wire w_mem_inst__abc_21203_new_n2726_; 
wire w_mem_inst__abc_21203_new_n2727_; 
wire w_mem_inst__abc_21203_new_n2728_; 
wire w_mem_inst__abc_21203_new_n2729_; 
wire w_mem_inst__abc_21203_new_n2730_; 
wire w_mem_inst__abc_21203_new_n2731_; 
wire w_mem_inst__abc_21203_new_n2732_; 
wire w_mem_inst__abc_21203_new_n2733_; 
wire w_mem_inst__abc_21203_new_n2734_; 
wire w_mem_inst__abc_21203_new_n2735_; 
wire w_mem_inst__abc_21203_new_n2736_; 
wire w_mem_inst__abc_21203_new_n2737_; 
wire w_mem_inst__abc_21203_new_n2738_; 
wire w_mem_inst__abc_21203_new_n2739_; 
wire w_mem_inst__abc_21203_new_n2740_; 
wire w_mem_inst__abc_21203_new_n2741_; 
wire w_mem_inst__abc_21203_new_n2742_; 
wire w_mem_inst__abc_21203_new_n2743_; 
wire w_mem_inst__abc_21203_new_n2744_; 
wire w_mem_inst__abc_21203_new_n2745_; 
wire w_mem_inst__abc_21203_new_n2746_; 
wire w_mem_inst__abc_21203_new_n2747_; 
wire w_mem_inst__abc_21203_new_n2748_; 
wire w_mem_inst__abc_21203_new_n2749_; 
wire w_mem_inst__abc_21203_new_n2750_; 
wire w_mem_inst__abc_21203_new_n2751_; 
wire w_mem_inst__abc_21203_new_n2752_; 
wire w_mem_inst__abc_21203_new_n2753_; 
wire w_mem_inst__abc_21203_new_n2754_; 
wire w_mem_inst__abc_21203_new_n2755_; 
wire w_mem_inst__abc_21203_new_n2756_; 
wire w_mem_inst__abc_21203_new_n2757_; 
wire w_mem_inst__abc_21203_new_n2758_; 
wire w_mem_inst__abc_21203_new_n2759_; 
wire w_mem_inst__abc_21203_new_n2760_; 
wire w_mem_inst__abc_21203_new_n2761_; 
wire w_mem_inst__abc_21203_new_n2762_; 
wire w_mem_inst__abc_21203_new_n2763_; 
wire w_mem_inst__abc_21203_new_n2764_; 
wire w_mem_inst__abc_21203_new_n2765_; 
wire w_mem_inst__abc_21203_new_n2766_; 
wire w_mem_inst__abc_21203_new_n2768_; 
wire w_mem_inst__abc_21203_new_n2769_; 
wire w_mem_inst__abc_21203_new_n2770_; 
wire w_mem_inst__abc_21203_new_n2771_; 
wire w_mem_inst__abc_21203_new_n2772_; 
wire w_mem_inst__abc_21203_new_n2773_; 
wire w_mem_inst__abc_21203_new_n2774_; 
wire w_mem_inst__abc_21203_new_n2775_; 
wire w_mem_inst__abc_21203_new_n2776_; 
wire w_mem_inst__abc_21203_new_n2777_; 
wire w_mem_inst__abc_21203_new_n2778_; 
wire w_mem_inst__abc_21203_new_n2779_; 
wire w_mem_inst__abc_21203_new_n2780_; 
wire w_mem_inst__abc_21203_new_n2781_; 
wire w_mem_inst__abc_21203_new_n2782_; 
wire w_mem_inst__abc_21203_new_n2783_; 
wire w_mem_inst__abc_21203_new_n2784_; 
wire w_mem_inst__abc_21203_new_n2785_; 
wire w_mem_inst__abc_21203_new_n2786_; 
wire w_mem_inst__abc_21203_new_n2787_; 
wire w_mem_inst__abc_21203_new_n2788_; 
wire w_mem_inst__abc_21203_new_n2789_; 
wire w_mem_inst__abc_21203_new_n2790_; 
wire w_mem_inst__abc_21203_new_n2791_; 
wire w_mem_inst__abc_21203_new_n2792_; 
wire w_mem_inst__abc_21203_new_n2793_; 
wire w_mem_inst__abc_21203_new_n2794_; 
wire w_mem_inst__abc_21203_new_n2795_; 
wire w_mem_inst__abc_21203_new_n2796_; 
wire w_mem_inst__abc_21203_new_n2797_; 
wire w_mem_inst__abc_21203_new_n2798_; 
wire w_mem_inst__abc_21203_new_n2799_; 
wire w_mem_inst__abc_21203_new_n2800_; 
wire w_mem_inst__abc_21203_new_n2801_; 
wire w_mem_inst__abc_21203_new_n2802_; 
wire w_mem_inst__abc_21203_new_n2803_; 
wire w_mem_inst__abc_21203_new_n2804_; 
wire w_mem_inst__abc_21203_new_n2805_; 
wire w_mem_inst__abc_21203_new_n2806_; 
wire w_mem_inst__abc_21203_new_n2807_; 
wire w_mem_inst__abc_21203_new_n2808_; 
wire w_mem_inst__abc_21203_new_n2809_; 
wire w_mem_inst__abc_21203_new_n2810_; 
wire w_mem_inst__abc_21203_new_n2811_; 
wire w_mem_inst__abc_21203_new_n2812_; 
wire w_mem_inst__abc_21203_new_n2813_; 
wire w_mem_inst__abc_21203_new_n2814_; 
wire w_mem_inst__abc_21203_new_n2816_; 
wire w_mem_inst__abc_21203_new_n2817_; 
wire w_mem_inst__abc_21203_new_n2818_; 
wire w_mem_inst__abc_21203_new_n2819_; 
wire w_mem_inst__abc_21203_new_n2820_; 
wire w_mem_inst__abc_21203_new_n2821_; 
wire w_mem_inst__abc_21203_new_n2822_; 
wire w_mem_inst__abc_21203_new_n2823_; 
wire w_mem_inst__abc_21203_new_n2824_; 
wire w_mem_inst__abc_21203_new_n2825_; 
wire w_mem_inst__abc_21203_new_n2826_; 
wire w_mem_inst__abc_21203_new_n2827_; 
wire w_mem_inst__abc_21203_new_n2828_; 
wire w_mem_inst__abc_21203_new_n2829_; 
wire w_mem_inst__abc_21203_new_n2830_; 
wire w_mem_inst__abc_21203_new_n2831_; 
wire w_mem_inst__abc_21203_new_n2832_; 
wire w_mem_inst__abc_21203_new_n2833_; 
wire w_mem_inst__abc_21203_new_n2834_; 
wire w_mem_inst__abc_21203_new_n2835_; 
wire w_mem_inst__abc_21203_new_n2836_; 
wire w_mem_inst__abc_21203_new_n2837_; 
wire w_mem_inst__abc_21203_new_n2838_; 
wire w_mem_inst__abc_21203_new_n2839_; 
wire w_mem_inst__abc_21203_new_n2840_; 
wire w_mem_inst__abc_21203_new_n2841_; 
wire w_mem_inst__abc_21203_new_n2842_; 
wire w_mem_inst__abc_21203_new_n2843_; 
wire w_mem_inst__abc_21203_new_n2844_; 
wire w_mem_inst__abc_21203_new_n2845_; 
wire w_mem_inst__abc_21203_new_n2846_; 
wire w_mem_inst__abc_21203_new_n2847_; 
wire w_mem_inst__abc_21203_new_n2848_; 
wire w_mem_inst__abc_21203_new_n2849_; 
wire w_mem_inst__abc_21203_new_n2850_; 
wire w_mem_inst__abc_21203_new_n2851_; 
wire w_mem_inst__abc_21203_new_n2852_; 
wire w_mem_inst__abc_21203_new_n2853_; 
wire w_mem_inst__abc_21203_new_n2854_; 
wire w_mem_inst__abc_21203_new_n2855_; 
wire w_mem_inst__abc_21203_new_n2856_; 
wire w_mem_inst__abc_21203_new_n2857_; 
wire w_mem_inst__abc_21203_new_n2858_; 
wire w_mem_inst__abc_21203_new_n2859_; 
wire w_mem_inst__abc_21203_new_n2860_; 
wire w_mem_inst__abc_21203_new_n2861_; 
wire w_mem_inst__abc_21203_new_n2862_; 
wire w_mem_inst__abc_21203_new_n2864_; 
wire w_mem_inst__abc_21203_new_n2865_; 
wire w_mem_inst__abc_21203_new_n2866_; 
wire w_mem_inst__abc_21203_new_n2867_; 
wire w_mem_inst__abc_21203_new_n2868_; 
wire w_mem_inst__abc_21203_new_n2869_; 
wire w_mem_inst__abc_21203_new_n2870_; 
wire w_mem_inst__abc_21203_new_n2871_; 
wire w_mem_inst__abc_21203_new_n2872_; 
wire w_mem_inst__abc_21203_new_n2873_; 
wire w_mem_inst__abc_21203_new_n2874_; 
wire w_mem_inst__abc_21203_new_n2875_; 
wire w_mem_inst__abc_21203_new_n2876_; 
wire w_mem_inst__abc_21203_new_n2877_; 
wire w_mem_inst__abc_21203_new_n2878_; 
wire w_mem_inst__abc_21203_new_n2879_; 
wire w_mem_inst__abc_21203_new_n2880_; 
wire w_mem_inst__abc_21203_new_n2881_; 
wire w_mem_inst__abc_21203_new_n2882_; 
wire w_mem_inst__abc_21203_new_n2883_; 
wire w_mem_inst__abc_21203_new_n2884_; 
wire w_mem_inst__abc_21203_new_n2885_; 
wire w_mem_inst__abc_21203_new_n2886_; 
wire w_mem_inst__abc_21203_new_n2887_; 
wire w_mem_inst__abc_21203_new_n2888_; 
wire w_mem_inst__abc_21203_new_n2889_; 
wire w_mem_inst__abc_21203_new_n2890_; 
wire w_mem_inst__abc_21203_new_n2891_; 
wire w_mem_inst__abc_21203_new_n2892_; 
wire w_mem_inst__abc_21203_new_n2893_; 
wire w_mem_inst__abc_21203_new_n2894_; 
wire w_mem_inst__abc_21203_new_n2895_; 
wire w_mem_inst__abc_21203_new_n2896_; 
wire w_mem_inst__abc_21203_new_n2897_; 
wire w_mem_inst__abc_21203_new_n2898_; 
wire w_mem_inst__abc_21203_new_n2899_; 
wire w_mem_inst__abc_21203_new_n2900_; 
wire w_mem_inst__abc_21203_new_n2901_; 
wire w_mem_inst__abc_21203_new_n2902_; 
wire w_mem_inst__abc_21203_new_n2903_; 
wire w_mem_inst__abc_21203_new_n2904_; 
wire w_mem_inst__abc_21203_new_n2905_; 
wire w_mem_inst__abc_21203_new_n2906_; 
wire w_mem_inst__abc_21203_new_n2907_; 
wire w_mem_inst__abc_21203_new_n2908_; 
wire w_mem_inst__abc_21203_new_n2909_; 
wire w_mem_inst__abc_21203_new_n2910_; 
wire w_mem_inst__abc_21203_new_n2912_; 
wire w_mem_inst__abc_21203_new_n2913_; 
wire w_mem_inst__abc_21203_new_n2914_; 
wire w_mem_inst__abc_21203_new_n2915_; 
wire w_mem_inst__abc_21203_new_n2916_; 
wire w_mem_inst__abc_21203_new_n2917_; 
wire w_mem_inst__abc_21203_new_n2918_; 
wire w_mem_inst__abc_21203_new_n2919_; 
wire w_mem_inst__abc_21203_new_n2920_; 
wire w_mem_inst__abc_21203_new_n2921_; 
wire w_mem_inst__abc_21203_new_n2922_; 
wire w_mem_inst__abc_21203_new_n2923_; 
wire w_mem_inst__abc_21203_new_n2924_; 
wire w_mem_inst__abc_21203_new_n2925_; 
wire w_mem_inst__abc_21203_new_n2926_; 
wire w_mem_inst__abc_21203_new_n2927_; 
wire w_mem_inst__abc_21203_new_n2928_; 
wire w_mem_inst__abc_21203_new_n2929_; 
wire w_mem_inst__abc_21203_new_n2930_; 
wire w_mem_inst__abc_21203_new_n2931_; 
wire w_mem_inst__abc_21203_new_n2932_; 
wire w_mem_inst__abc_21203_new_n2933_; 
wire w_mem_inst__abc_21203_new_n2934_; 
wire w_mem_inst__abc_21203_new_n2935_; 
wire w_mem_inst__abc_21203_new_n2936_; 
wire w_mem_inst__abc_21203_new_n2937_; 
wire w_mem_inst__abc_21203_new_n2938_; 
wire w_mem_inst__abc_21203_new_n2939_; 
wire w_mem_inst__abc_21203_new_n2940_; 
wire w_mem_inst__abc_21203_new_n2941_; 
wire w_mem_inst__abc_21203_new_n2942_; 
wire w_mem_inst__abc_21203_new_n2943_; 
wire w_mem_inst__abc_21203_new_n2944_; 
wire w_mem_inst__abc_21203_new_n2945_; 
wire w_mem_inst__abc_21203_new_n2946_; 
wire w_mem_inst__abc_21203_new_n2947_; 
wire w_mem_inst__abc_21203_new_n2948_; 
wire w_mem_inst__abc_21203_new_n2949_; 
wire w_mem_inst__abc_21203_new_n2950_; 
wire w_mem_inst__abc_21203_new_n2951_; 
wire w_mem_inst__abc_21203_new_n2952_; 
wire w_mem_inst__abc_21203_new_n2953_; 
wire w_mem_inst__abc_21203_new_n2954_; 
wire w_mem_inst__abc_21203_new_n2955_; 
wire w_mem_inst__abc_21203_new_n2956_; 
wire w_mem_inst__abc_21203_new_n2957_; 
wire w_mem_inst__abc_21203_new_n2958_; 
wire w_mem_inst__abc_21203_new_n2960_; 
wire w_mem_inst__abc_21203_new_n2961_; 
wire w_mem_inst__abc_21203_new_n2962_; 
wire w_mem_inst__abc_21203_new_n2963_; 
wire w_mem_inst__abc_21203_new_n2964_; 
wire w_mem_inst__abc_21203_new_n2965_; 
wire w_mem_inst__abc_21203_new_n2966_; 
wire w_mem_inst__abc_21203_new_n2967_; 
wire w_mem_inst__abc_21203_new_n2968_; 
wire w_mem_inst__abc_21203_new_n2969_; 
wire w_mem_inst__abc_21203_new_n2970_; 
wire w_mem_inst__abc_21203_new_n2971_; 
wire w_mem_inst__abc_21203_new_n2972_; 
wire w_mem_inst__abc_21203_new_n2973_; 
wire w_mem_inst__abc_21203_new_n2974_; 
wire w_mem_inst__abc_21203_new_n2975_; 
wire w_mem_inst__abc_21203_new_n2976_; 
wire w_mem_inst__abc_21203_new_n2977_; 
wire w_mem_inst__abc_21203_new_n2978_; 
wire w_mem_inst__abc_21203_new_n2979_; 
wire w_mem_inst__abc_21203_new_n2980_; 
wire w_mem_inst__abc_21203_new_n2981_; 
wire w_mem_inst__abc_21203_new_n2982_; 
wire w_mem_inst__abc_21203_new_n2983_; 
wire w_mem_inst__abc_21203_new_n2984_; 
wire w_mem_inst__abc_21203_new_n2985_; 
wire w_mem_inst__abc_21203_new_n2986_; 
wire w_mem_inst__abc_21203_new_n2987_; 
wire w_mem_inst__abc_21203_new_n2988_; 
wire w_mem_inst__abc_21203_new_n2989_; 
wire w_mem_inst__abc_21203_new_n2990_; 
wire w_mem_inst__abc_21203_new_n2991_; 
wire w_mem_inst__abc_21203_new_n2992_; 
wire w_mem_inst__abc_21203_new_n2993_; 
wire w_mem_inst__abc_21203_new_n2994_; 
wire w_mem_inst__abc_21203_new_n2995_; 
wire w_mem_inst__abc_21203_new_n2996_; 
wire w_mem_inst__abc_21203_new_n2997_; 
wire w_mem_inst__abc_21203_new_n2998_; 
wire w_mem_inst__abc_21203_new_n2999_; 
wire w_mem_inst__abc_21203_new_n3000_; 
wire w_mem_inst__abc_21203_new_n3001_; 
wire w_mem_inst__abc_21203_new_n3002_; 
wire w_mem_inst__abc_21203_new_n3003_; 
wire w_mem_inst__abc_21203_new_n3004_; 
wire w_mem_inst__abc_21203_new_n3005_; 
wire w_mem_inst__abc_21203_new_n3006_; 
wire w_mem_inst__abc_21203_new_n3008_; 
wire w_mem_inst__abc_21203_new_n3009_; 
wire w_mem_inst__abc_21203_new_n3010_; 
wire w_mem_inst__abc_21203_new_n3011_; 
wire w_mem_inst__abc_21203_new_n3012_; 
wire w_mem_inst__abc_21203_new_n3013_; 
wire w_mem_inst__abc_21203_new_n3014_; 
wire w_mem_inst__abc_21203_new_n3015_; 
wire w_mem_inst__abc_21203_new_n3016_; 
wire w_mem_inst__abc_21203_new_n3017_; 
wire w_mem_inst__abc_21203_new_n3018_; 
wire w_mem_inst__abc_21203_new_n3019_; 
wire w_mem_inst__abc_21203_new_n3020_; 
wire w_mem_inst__abc_21203_new_n3021_; 
wire w_mem_inst__abc_21203_new_n3022_; 
wire w_mem_inst__abc_21203_new_n3023_; 
wire w_mem_inst__abc_21203_new_n3024_; 
wire w_mem_inst__abc_21203_new_n3025_; 
wire w_mem_inst__abc_21203_new_n3026_; 
wire w_mem_inst__abc_21203_new_n3027_; 
wire w_mem_inst__abc_21203_new_n3028_; 
wire w_mem_inst__abc_21203_new_n3029_; 
wire w_mem_inst__abc_21203_new_n3030_; 
wire w_mem_inst__abc_21203_new_n3031_; 
wire w_mem_inst__abc_21203_new_n3032_; 
wire w_mem_inst__abc_21203_new_n3033_; 
wire w_mem_inst__abc_21203_new_n3034_; 
wire w_mem_inst__abc_21203_new_n3035_; 
wire w_mem_inst__abc_21203_new_n3036_; 
wire w_mem_inst__abc_21203_new_n3037_; 
wire w_mem_inst__abc_21203_new_n3038_; 
wire w_mem_inst__abc_21203_new_n3039_; 
wire w_mem_inst__abc_21203_new_n3040_; 
wire w_mem_inst__abc_21203_new_n3041_; 
wire w_mem_inst__abc_21203_new_n3042_; 
wire w_mem_inst__abc_21203_new_n3043_; 
wire w_mem_inst__abc_21203_new_n3044_; 
wire w_mem_inst__abc_21203_new_n3045_; 
wire w_mem_inst__abc_21203_new_n3046_; 
wire w_mem_inst__abc_21203_new_n3047_; 
wire w_mem_inst__abc_21203_new_n3048_; 
wire w_mem_inst__abc_21203_new_n3049_; 
wire w_mem_inst__abc_21203_new_n3050_; 
wire w_mem_inst__abc_21203_new_n3051_; 
wire w_mem_inst__abc_21203_new_n3052_; 
wire w_mem_inst__abc_21203_new_n3053_; 
wire w_mem_inst__abc_21203_new_n3054_; 
wire w_mem_inst__abc_21203_new_n3056_; 
wire w_mem_inst__abc_21203_new_n3057_; 
wire w_mem_inst__abc_21203_new_n3058_; 
wire w_mem_inst__abc_21203_new_n3059_; 
wire w_mem_inst__abc_21203_new_n3060_; 
wire w_mem_inst__abc_21203_new_n3061_; 
wire w_mem_inst__abc_21203_new_n3062_; 
wire w_mem_inst__abc_21203_new_n3063_; 
wire w_mem_inst__abc_21203_new_n3064_; 
wire w_mem_inst__abc_21203_new_n3065_; 
wire w_mem_inst__abc_21203_new_n3066_; 
wire w_mem_inst__abc_21203_new_n3067_; 
wire w_mem_inst__abc_21203_new_n3068_; 
wire w_mem_inst__abc_21203_new_n3069_; 
wire w_mem_inst__abc_21203_new_n3070_; 
wire w_mem_inst__abc_21203_new_n3071_; 
wire w_mem_inst__abc_21203_new_n3072_; 
wire w_mem_inst__abc_21203_new_n3073_; 
wire w_mem_inst__abc_21203_new_n3074_; 
wire w_mem_inst__abc_21203_new_n3075_; 
wire w_mem_inst__abc_21203_new_n3076_; 
wire w_mem_inst__abc_21203_new_n3077_; 
wire w_mem_inst__abc_21203_new_n3078_; 
wire w_mem_inst__abc_21203_new_n3079_; 
wire w_mem_inst__abc_21203_new_n3080_; 
wire w_mem_inst__abc_21203_new_n3081_; 
wire w_mem_inst__abc_21203_new_n3082_; 
wire w_mem_inst__abc_21203_new_n3083_; 
wire w_mem_inst__abc_21203_new_n3084_; 
wire w_mem_inst__abc_21203_new_n3085_; 
wire w_mem_inst__abc_21203_new_n3086_; 
wire w_mem_inst__abc_21203_new_n3087_; 
wire w_mem_inst__abc_21203_new_n3088_; 
wire w_mem_inst__abc_21203_new_n3089_; 
wire w_mem_inst__abc_21203_new_n3090_; 
wire w_mem_inst__abc_21203_new_n3091_; 
wire w_mem_inst__abc_21203_new_n3092_; 
wire w_mem_inst__abc_21203_new_n3093_; 
wire w_mem_inst__abc_21203_new_n3094_; 
wire w_mem_inst__abc_21203_new_n3095_; 
wire w_mem_inst__abc_21203_new_n3096_; 
wire w_mem_inst__abc_21203_new_n3097_; 
wire w_mem_inst__abc_21203_new_n3098_; 
wire w_mem_inst__abc_21203_new_n3099_; 
wire w_mem_inst__abc_21203_new_n3100_; 
wire w_mem_inst__abc_21203_new_n3101_; 
wire w_mem_inst__abc_21203_new_n3102_; 
wire w_mem_inst__abc_21203_new_n3104_; 
wire w_mem_inst__abc_21203_new_n3105_; 
wire w_mem_inst__abc_21203_new_n3106_; 
wire w_mem_inst__abc_21203_new_n3107_; 
wire w_mem_inst__abc_21203_new_n3108_; 
wire w_mem_inst__abc_21203_new_n3109_; 
wire w_mem_inst__abc_21203_new_n3110_; 
wire w_mem_inst__abc_21203_new_n3111_; 
wire w_mem_inst__abc_21203_new_n3112_; 
wire w_mem_inst__abc_21203_new_n3113_; 
wire w_mem_inst__abc_21203_new_n3114_; 
wire w_mem_inst__abc_21203_new_n3115_; 
wire w_mem_inst__abc_21203_new_n3116_; 
wire w_mem_inst__abc_21203_new_n3117_; 
wire w_mem_inst__abc_21203_new_n3118_; 
wire w_mem_inst__abc_21203_new_n3119_; 
wire w_mem_inst__abc_21203_new_n3120_; 
wire w_mem_inst__abc_21203_new_n3121_; 
wire w_mem_inst__abc_21203_new_n3122_; 
wire w_mem_inst__abc_21203_new_n3123_; 
wire w_mem_inst__abc_21203_new_n3124_; 
wire w_mem_inst__abc_21203_new_n3125_; 
wire w_mem_inst__abc_21203_new_n3126_; 
wire w_mem_inst__abc_21203_new_n3127_; 
wire w_mem_inst__abc_21203_new_n3128_; 
wire w_mem_inst__abc_21203_new_n3129_; 
wire w_mem_inst__abc_21203_new_n3130_; 
wire w_mem_inst__abc_21203_new_n3131_; 
wire w_mem_inst__abc_21203_new_n3132_; 
wire w_mem_inst__abc_21203_new_n3133_; 
wire w_mem_inst__abc_21203_new_n3134_; 
wire w_mem_inst__abc_21203_new_n3135_; 
wire w_mem_inst__abc_21203_new_n3136_; 
wire w_mem_inst__abc_21203_new_n3137_; 
wire w_mem_inst__abc_21203_new_n3138_; 
wire w_mem_inst__abc_21203_new_n3139_; 
wire w_mem_inst__abc_21203_new_n3140_; 
wire w_mem_inst__abc_21203_new_n3141_; 
wire w_mem_inst__abc_21203_new_n3142_; 
wire w_mem_inst__abc_21203_new_n3143_; 
wire w_mem_inst__abc_21203_new_n3144_; 
wire w_mem_inst__abc_21203_new_n3145_; 
wire w_mem_inst__abc_21203_new_n3146_; 
wire w_mem_inst__abc_21203_new_n3147_; 
wire w_mem_inst__abc_21203_new_n3148_; 
wire w_mem_inst__abc_21203_new_n3149_; 
wire w_mem_inst__abc_21203_new_n3150_; 
wire w_mem_inst__abc_21203_new_n3152_; 
wire w_mem_inst__abc_21203_new_n3153_; 
wire w_mem_inst__abc_21203_new_n3154_; 
wire w_mem_inst__abc_21203_new_n3155_; 
wire w_mem_inst__abc_21203_new_n3156_; 
wire w_mem_inst__abc_21203_new_n3157_; 
wire w_mem_inst__abc_21203_new_n3158_; 
wire w_mem_inst__abc_21203_new_n3159_; 
wire w_mem_inst__abc_21203_new_n3160_; 
wire w_mem_inst__abc_21203_new_n3162_; 
wire w_mem_inst__abc_21203_new_n3163_; 
wire w_mem_inst__abc_21203_new_n3164_; 
wire w_mem_inst__abc_21203_new_n3165_; 
wire w_mem_inst__abc_21203_new_n3166_; 
wire w_mem_inst__abc_21203_new_n3168_; 
wire w_mem_inst__abc_21203_new_n3169_; 
wire w_mem_inst__abc_21203_new_n3170_; 
wire w_mem_inst__abc_21203_new_n3171_; 
wire w_mem_inst__abc_21203_new_n3172_; 
wire w_mem_inst__abc_21203_new_n3174_; 
wire w_mem_inst__abc_21203_new_n3175_; 
wire w_mem_inst__abc_21203_new_n3176_; 
wire w_mem_inst__abc_21203_new_n3177_; 
wire w_mem_inst__abc_21203_new_n3178_; 
wire w_mem_inst__abc_21203_new_n3180_; 
wire w_mem_inst__abc_21203_new_n3181_; 
wire w_mem_inst__abc_21203_new_n3182_; 
wire w_mem_inst__abc_21203_new_n3183_; 
wire w_mem_inst__abc_21203_new_n3184_; 
wire w_mem_inst__abc_21203_new_n3186_; 
wire w_mem_inst__abc_21203_new_n3187_; 
wire w_mem_inst__abc_21203_new_n3188_; 
wire w_mem_inst__abc_21203_new_n3189_; 
wire w_mem_inst__abc_21203_new_n3190_; 
wire w_mem_inst__abc_21203_new_n3192_; 
wire w_mem_inst__abc_21203_new_n3193_; 
wire w_mem_inst__abc_21203_new_n3194_; 
wire w_mem_inst__abc_21203_new_n3195_; 
wire w_mem_inst__abc_21203_new_n3196_; 
wire w_mem_inst__abc_21203_new_n3198_; 
wire w_mem_inst__abc_21203_new_n3199_; 
wire w_mem_inst__abc_21203_new_n3200_; 
wire w_mem_inst__abc_21203_new_n3201_; 
wire w_mem_inst__abc_21203_new_n3202_; 
wire w_mem_inst__abc_21203_new_n3204_; 
wire w_mem_inst__abc_21203_new_n3205_; 
wire w_mem_inst__abc_21203_new_n3206_; 
wire w_mem_inst__abc_21203_new_n3207_; 
wire w_mem_inst__abc_21203_new_n3208_; 
wire w_mem_inst__abc_21203_new_n3210_; 
wire w_mem_inst__abc_21203_new_n3211_; 
wire w_mem_inst__abc_21203_new_n3212_; 
wire w_mem_inst__abc_21203_new_n3213_; 
wire w_mem_inst__abc_21203_new_n3214_; 
wire w_mem_inst__abc_21203_new_n3216_; 
wire w_mem_inst__abc_21203_new_n3217_; 
wire w_mem_inst__abc_21203_new_n3218_; 
wire w_mem_inst__abc_21203_new_n3219_; 
wire w_mem_inst__abc_21203_new_n3220_; 
wire w_mem_inst__abc_21203_new_n3222_; 
wire w_mem_inst__abc_21203_new_n3223_; 
wire w_mem_inst__abc_21203_new_n3224_; 
wire w_mem_inst__abc_21203_new_n3225_; 
wire w_mem_inst__abc_21203_new_n3226_; 
wire w_mem_inst__abc_21203_new_n3228_; 
wire w_mem_inst__abc_21203_new_n3229_; 
wire w_mem_inst__abc_21203_new_n3230_; 
wire w_mem_inst__abc_21203_new_n3231_; 
wire w_mem_inst__abc_21203_new_n3232_; 
wire w_mem_inst__abc_21203_new_n3234_; 
wire w_mem_inst__abc_21203_new_n3235_; 
wire w_mem_inst__abc_21203_new_n3236_; 
wire w_mem_inst__abc_21203_new_n3237_; 
wire w_mem_inst__abc_21203_new_n3238_; 
wire w_mem_inst__abc_21203_new_n3240_; 
wire w_mem_inst__abc_21203_new_n3241_; 
wire w_mem_inst__abc_21203_new_n3242_; 
wire w_mem_inst__abc_21203_new_n3243_; 
wire w_mem_inst__abc_21203_new_n3244_; 
wire w_mem_inst__abc_21203_new_n3246_; 
wire w_mem_inst__abc_21203_new_n3247_; 
wire w_mem_inst__abc_21203_new_n3248_; 
wire w_mem_inst__abc_21203_new_n3249_; 
wire w_mem_inst__abc_21203_new_n3250_; 
wire w_mem_inst__abc_21203_new_n3252_; 
wire w_mem_inst__abc_21203_new_n3253_; 
wire w_mem_inst__abc_21203_new_n3254_; 
wire w_mem_inst__abc_21203_new_n3255_; 
wire w_mem_inst__abc_21203_new_n3256_; 
wire w_mem_inst__abc_21203_new_n3258_; 
wire w_mem_inst__abc_21203_new_n3259_; 
wire w_mem_inst__abc_21203_new_n3260_; 
wire w_mem_inst__abc_21203_new_n3261_; 
wire w_mem_inst__abc_21203_new_n3262_; 
wire w_mem_inst__abc_21203_new_n3264_; 
wire w_mem_inst__abc_21203_new_n3265_; 
wire w_mem_inst__abc_21203_new_n3266_; 
wire w_mem_inst__abc_21203_new_n3267_; 
wire w_mem_inst__abc_21203_new_n3268_; 
wire w_mem_inst__abc_21203_new_n3270_; 
wire w_mem_inst__abc_21203_new_n3271_; 
wire w_mem_inst__abc_21203_new_n3272_; 
wire w_mem_inst__abc_21203_new_n3273_; 
wire w_mem_inst__abc_21203_new_n3274_; 
wire w_mem_inst__abc_21203_new_n3276_; 
wire w_mem_inst__abc_21203_new_n3277_; 
wire w_mem_inst__abc_21203_new_n3278_; 
wire w_mem_inst__abc_21203_new_n3279_; 
wire w_mem_inst__abc_21203_new_n3280_; 
wire w_mem_inst__abc_21203_new_n3282_; 
wire w_mem_inst__abc_21203_new_n3283_; 
wire w_mem_inst__abc_21203_new_n3284_; 
wire w_mem_inst__abc_21203_new_n3285_; 
wire w_mem_inst__abc_21203_new_n3286_; 
wire w_mem_inst__abc_21203_new_n3288_; 
wire w_mem_inst__abc_21203_new_n3289_; 
wire w_mem_inst__abc_21203_new_n3290_; 
wire w_mem_inst__abc_21203_new_n3291_; 
wire w_mem_inst__abc_21203_new_n3292_; 
wire w_mem_inst__abc_21203_new_n3294_; 
wire w_mem_inst__abc_21203_new_n3295_; 
wire w_mem_inst__abc_21203_new_n3296_; 
wire w_mem_inst__abc_21203_new_n3297_; 
wire w_mem_inst__abc_21203_new_n3298_; 
wire w_mem_inst__abc_21203_new_n3300_; 
wire w_mem_inst__abc_21203_new_n3301_; 
wire w_mem_inst__abc_21203_new_n3302_; 
wire w_mem_inst__abc_21203_new_n3303_; 
wire w_mem_inst__abc_21203_new_n3304_; 
wire w_mem_inst__abc_21203_new_n3306_; 
wire w_mem_inst__abc_21203_new_n3307_; 
wire w_mem_inst__abc_21203_new_n3308_; 
wire w_mem_inst__abc_21203_new_n3309_; 
wire w_mem_inst__abc_21203_new_n3310_; 
wire w_mem_inst__abc_21203_new_n3312_; 
wire w_mem_inst__abc_21203_new_n3313_; 
wire w_mem_inst__abc_21203_new_n3314_; 
wire w_mem_inst__abc_21203_new_n3315_; 
wire w_mem_inst__abc_21203_new_n3316_; 
wire w_mem_inst__abc_21203_new_n3318_; 
wire w_mem_inst__abc_21203_new_n3319_; 
wire w_mem_inst__abc_21203_new_n3320_; 
wire w_mem_inst__abc_21203_new_n3321_; 
wire w_mem_inst__abc_21203_new_n3322_; 
wire w_mem_inst__abc_21203_new_n3324_; 
wire w_mem_inst__abc_21203_new_n3325_; 
wire w_mem_inst__abc_21203_new_n3326_; 
wire w_mem_inst__abc_21203_new_n3327_; 
wire w_mem_inst__abc_21203_new_n3328_; 
wire w_mem_inst__abc_21203_new_n3330_; 
wire w_mem_inst__abc_21203_new_n3331_; 
wire w_mem_inst__abc_21203_new_n3332_; 
wire w_mem_inst__abc_21203_new_n3333_; 
wire w_mem_inst__abc_21203_new_n3334_; 
wire w_mem_inst__abc_21203_new_n3336_; 
wire w_mem_inst__abc_21203_new_n3337_; 
wire w_mem_inst__abc_21203_new_n3338_; 
wire w_mem_inst__abc_21203_new_n3339_; 
wire w_mem_inst__abc_21203_new_n3340_; 
wire w_mem_inst__abc_21203_new_n3342_; 
wire w_mem_inst__abc_21203_new_n3343_; 
wire w_mem_inst__abc_21203_new_n3344_; 
wire w_mem_inst__abc_21203_new_n3345_; 
wire w_mem_inst__abc_21203_new_n3346_; 
wire w_mem_inst__abc_21203_new_n3348_; 
wire w_mem_inst__abc_21203_new_n3349_; 
wire w_mem_inst__abc_21203_new_n3350_; 
wire w_mem_inst__abc_21203_new_n3351_; 
wire w_mem_inst__abc_21203_new_n3352_; 
wire w_mem_inst__abc_21203_new_n3354_; 
wire w_mem_inst__abc_21203_new_n3355_; 
wire w_mem_inst__abc_21203_new_n3356_; 
wire w_mem_inst__abc_21203_new_n3357_; 
wire w_mem_inst__abc_21203_new_n3358_; 
wire w_mem_inst__abc_21203_new_n3360_; 
wire w_mem_inst__abc_21203_new_n3361_; 
wire w_mem_inst__abc_21203_new_n3362_; 
wire w_mem_inst__abc_21203_new_n3363_; 
wire w_mem_inst__abc_21203_new_n3364_; 
wire w_mem_inst__abc_21203_new_n3366_; 
wire w_mem_inst__abc_21203_new_n3367_; 
wire w_mem_inst__abc_21203_new_n3368_; 
wire w_mem_inst__abc_21203_new_n3369_; 
wire w_mem_inst__abc_21203_new_n3370_; 
wire w_mem_inst__abc_21203_new_n3372_; 
wire w_mem_inst__abc_21203_new_n3373_; 
wire w_mem_inst__abc_21203_new_n3374_; 
wire w_mem_inst__abc_21203_new_n3375_; 
wire w_mem_inst__abc_21203_new_n3376_; 
wire w_mem_inst__abc_21203_new_n3378_; 
wire w_mem_inst__abc_21203_new_n3379_; 
wire w_mem_inst__abc_21203_new_n3380_; 
wire w_mem_inst__abc_21203_new_n3381_; 
wire w_mem_inst__abc_21203_new_n3382_; 
wire w_mem_inst__abc_21203_new_n3384_; 
wire w_mem_inst__abc_21203_new_n3385_; 
wire w_mem_inst__abc_21203_new_n3386_; 
wire w_mem_inst__abc_21203_new_n3387_; 
wire w_mem_inst__abc_21203_new_n3388_; 
wire w_mem_inst__abc_21203_new_n3390_; 
wire w_mem_inst__abc_21203_new_n3391_; 
wire w_mem_inst__abc_21203_new_n3392_; 
wire w_mem_inst__abc_21203_new_n3393_; 
wire w_mem_inst__abc_21203_new_n3394_; 
wire w_mem_inst__abc_21203_new_n3396_; 
wire w_mem_inst__abc_21203_new_n3397_; 
wire w_mem_inst__abc_21203_new_n3398_; 
wire w_mem_inst__abc_21203_new_n3399_; 
wire w_mem_inst__abc_21203_new_n3400_; 
wire w_mem_inst__abc_21203_new_n3402_; 
wire w_mem_inst__abc_21203_new_n3403_; 
wire w_mem_inst__abc_21203_new_n3404_; 
wire w_mem_inst__abc_21203_new_n3405_; 
wire w_mem_inst__abc_21203_new_n3406_; 
wire w_mem_inst__abc_21203_new_n3408_; 
wire w_mem_inst__abc_21203_new_n3409_; 
wire w_mem_inst__abc_21203_new_n3410_; 
wire w_mem_inst__abc_21203_new_n3411_; 
wire w_mem_inst__abc_21203_new_n3412_; 
wire w_mem_inst__abc_21203_new_n3414_; 
wire w_mem_inst__abc_21203_new_n3415_; 
wire w_mem_inst__abc_21203_new_n3416_; 
wire w_mem_inst__abc_21203_new_n3417_; 
wire w_mem_inst__abc_21203_new_n3418_; 
wire w_mem_inst__abc_21203_new_n3420_; 
wire w_mem_inst__abc_21203_new_n3421_; 
wire w_mem_inst__abc_21203_new_n3422_; 
wire w_mem_inst__abc_21203_new_n3423_; 
wire w_mem_inst__abc_21203_new_n3424_; 
wire w_mem_inst__abc_21203_new_n3426_; 
wire w_mem_inst__abc_21203_new_n3427_; 
wire w_mem_inst__abc_21203_new_n3428_; 
wire w_mem_inst__abc_21203_new_n3429_; 
wire w_mem_inst__abc_21203_new_n3430_; 
wire w_mem_inst__abc_21203_new_n3432_; 
wire w_mem_inst__abc_21203_new_n3433_; 
wire w_mem_inst__abc_21203_new_n3434_; 
wire w_mem_inst__abc_21203_new_n3435_; 
wire w_mem_inst__abc_21203_new_n3436_; 
wire w_mem_inst__abc_21203_new_n3438_; 
wire w_mem_inst__abc_21203_new_n3439_; 
wire w_mem_inst__abc_21203_new_n3440_; 
wire w_mem_inst__abc_21203_new_n3441_; 
wire w_mem_inst__abc_21203_new_n3442_; 
wire w_mem_inst__abc_21203_new_n3444_; 
wire w_mem_inst__abc_21203_new_n3445_; 
wire w_mem_inst__abc_21203_new_n3446_; 
wire w_mem_inst__abc_21203_new_n3447_; 
wire w_mem_inst__abc_21203_new_n3448_; 
wire w_mem_inst__abc_21203_new_n3450_; 
wire w_mem_inst__abc_21203_new_n3451_; 
wire w_mem_inst__abc_21203_new_n3452_; 
wire w_mem_inst__abc_21203_new_n3453_; 
wire w_mem_inst__abc_21203_new_n3454_; 
wire w_mem_inst__abc_21203_new_n3456_; 
wire w_mem_inst__abc_21203_new_n3457_; 
wire w_mem_inst__abc_21203_new_n3458_; 
wire w_mem_inst__abc_21203_new_n3459_; 
wire w_mem_inst__abc_21203_new_n3460_; 
wire w_mem_inst__abc_21203_new_n3462_; 
wire w_mem_inst__abc_21203_new_n3463_; 
wire w_mem_inst__abc_21203_new_n3464_; 
wire w_mem_inst__abc_21203_new_n3465_; 
wire w_mem_inst__abc_21203_new_n3466_; 
wire w_mem_inst__abc_21203_new_n3468_; 
wire w_mem_inst__abc_21203_new_n3469_; 
wire w_mem_inst__abc_21203_new_n3470_; 
wire w_mem_inst__abc_21203_new_n3471_; 
wire w_mem_inst__abc_21203_new_n3472_; 
wire w_mem_inst__abc_21203_new_n3474_; 
wire w_mem_inst__abc_21203_new_n3475_; 
wire w_mem_inst__abc_21203_new_n3476_; 
wire w_mem_inst__abc_21203_new_n3477_; 
wire w_mem_inst__abc_21203_new_n3478_; 
wire w_mem_inst__abc_21203_new_n3480_; 
wire w_mem_inst__abc_21203_new_n3481_; 
wire w_mem_inst__abc_21203_new_n3482_; 
wire w_mem_inst__abc_21203_new_n3483_; 
wire w_mem_inst__abc_21203_new_n3484_; 
wire w_mem_inst__abc_21203_new_n3486_; 
wire w_mem_inst__abc_21203_new_n3487_; 
wire w_mem_inst__abc_21203_new_n3488_; 
wire w_mem_inst__abc_21203_new_n3489_; 
wire w_mem_inst__abc_21203_new_n3490_; 
wire w_mem_inst__abc_21203_new_n3492_; 
wire w_mem_inst__abc_21203_new_n3493_; 
wire w_mem_inst__abc_21203_new_n3494_; 
wire w_mem_inst__abc_21203_new_n3495_; 
wire w_mem_inst__abc_21203_new_n3496_; 
wire w_mem_inst__abc_21203_new_n3498_; 
wire w_mem_inst__abc_21203_new_n3499_; 
wire w_mem_inst__abc_21203_new_n3500_; 
wire w_mem_inst__abc_21203_new_n3501_; 
wire w_mem_inst__abc_21203_new_n3502_; 
wire w_mem_inst__abc_21203_new_n3504_; 
wire w_mem_inst__abc_21203_new_n3505_; 
wire w_mem_inst__abc_21203_new_n3506_; 
wire w_mem_inst__abc_21203_new_n3507_; 
wire w_mem_inst__abc_21203_new_n3508_; 
wire w_mem_inst__abc_21203_new_n3510_; 
wire w_mem_inst__abc_21203_new_n3511_; 
wire w_mem_inst__abc_21203_new_n3512_; 
wire w_mem_inst__abc_21203_new_n3513_; 
wire w_mem_inst__abc_21203_new_n3514_; 
wire w_mem_inst__abc_21203_new_n3516_; 
wire w_mem_inst__abc_21203_new_n3517_; 
wire w_mem_inst__abc_21203_new_n3518_; 
wire w_mem_inst__abc_21203_new_n3519_; 
wire w_mem_inst__abc_21203_new_n3520_; 
wire w_mem_inst__abc_21203_new_n3522_; 
wire w_mem_inst__abc_21203_new_n3523_; 
wire w_mem_inst__abc_21203_new_n3524_; 
wire w_mem_inst__abc_21203_new_n3525_; 
wire w_mem_inst__abc_21203_new_n3526_; 
wire w_mem_inst__abc_21203_new_n3528_; 
wire w_mem_inst__abc_21203_new_n3529_; 
wire w_mem_inst__abc_21203_new_n3530_; 
wire w_mem_inst__abc_21203_new_n3531_; 
wire w_mem_inst__abc_21203_new_n3532_; 
wire w_mem_inst__abc_21203_new_n3534_; 
wire w_mem_inst__abc_21203_new_n3535_; 
wire w_mem_inst__abc_21203_new_n3536_; 
wire w_mem_inst__abc_21203_new_n3537_; 
wire w_mem_inst__abc_21203_new_n3538_; 
wire w_mem_inst__abc_21203_new_n3540_; 
wire w_mem_inst__abc_21203_new_n3541_; 
wire w_mem_inst__abc_21203_new_n3542_; 
wire w_mem_inst__abc_21203_new_n3543_; 
wire w_mem_inst__abc_21203_new_n3544_; 
wire w_mem_inst__abc_21203_new_n3546_; 
wire w_mem_inst__abc_21203_new_n3547_; 
wire w_mem_inst__abc_21203_new_n3548_; 
wire w_mem_inst__abc_21203_new_n3549_; 
wire w_mem_inst__abc_21203_new_n3550_; 
wire w_mem_inst__abc_21203_new_n3552_; 
wire w_mem_inst__abc_21203_new_n3553_; 
wire w_mem_inst__abc_21203_new_n3554_; 
wire w_mem_inst__abc_21203_new_n3555_; 
wire w_mem_inst__abc_21203_new_n3556_; 
wire w_mem_inst__abc_21203_new_n3558_; 
wire w_mem_inst__abc_21203_new_n3559_; 
wire w_mem_inst__abc_21203_new_n3560_; 
wire w_mem_inst__abc_21203_new_n3561_; 
wire w_mem_inst__abc_21203_new_n3562_; 
wire w_mem_inst__abc_21203_new_n3564_; 
wire w_mem_inst__abc_21203_new_n3565_; 
wire w_mem_inst__abc_21203_new_n3566_; 
wire w_mem_inst__abc_21203_new_n3567_; 
wire w_mem_inst__abc_21203_new_n3568_; 
wire w_mem_inst__abc_21203_new_n3570_; 
wire w_mem_inst__abc_21203_new_n3571_; 
wire w_mem_inst__abc_21203_new_n3572_; 
wire w_mem_inst__abc_21203_new_n3573_; 
wire w_mem_inst__abc_21203_new_n3574_; 
wire w_mem_inst__abc_21203_new_n3576_; 
wire w_mem_inst__abc_21203_new_n3577_; 
wire w_mem_inst__abc_21203_new_n3578_; 
wire w_mem_inst__abc_21203_new_n3579_; 
wire w_mem_inst__abc_21203_new_n3580_; 
wire w_mem_inst__abc_21203_new_n3582_; 
wire w_mem_inst__abc_21203_new_n3583_; 
wire w_mem_inst__abc_21203_new_n3584_; 
wire w_mem_inst__abc_21203_new_n3585_; 
wire w_mem_inst__abc_21203_new_n3586_; 
wire w_mem_inst__abc_21203_new_n3588_; 
wire w_mem_inst__abc_21203_new_n3589_; 
wire w_mem_inst__abc_21203_new_n3590_; 
wire w_mem_inst__abc_21203_new_n3591_; 
wire w_mem_inst__abc_21203_new_n3592_; 
wire w_mem_inst__abc_21203_new_n3594_; 
wire w_mem_inst__abc_21203_new_n3595_; 
wire w_mem_inst__abc_21203_new_n3596_; 
wire w_mem_inst__abc_21203_new_n3597_; 
wire w_mem_inst__abc_21203_new_n3598_; 
wire w_mem_inst__abc_21203_new_n3600_; 
wire w_mem_inst__abc_21203_new_n3601_; 
wire w_mem_inst__abc_21203_new_n3602_; 
wire w_mem_inst__abc_21203_new_n3603_; 
wire w_mem_inst__abc_21203_new_n3604_; 
wire w_mem_inst__abc_21203_new_n3606_; 
wire w_mem_inst__abc_21203_new_n3607_; 
wire w_mem_inst__abc_21203_new_n3608_; 
wire w_mem_inst__abc_21203_new_n3609_; 
wire w_mem_inst__abc_21203_new_n3610_; 
wire w_mem_inst__abc_21203_new_n3612_; 
wire w_mem_inst__abc_21203_new_n3613_; 
wire w_mem_inst__abc_21203_new_n3614_; 
wire w_mem_inst__abc_21203_new_n3615_; 
wire w_mem_inst__abc_21203_new_n3616_; 
wire w_mem_inst__abc_21203_new_n3618_; 
wire w_mem_inst__abc_21203_new_n3619_; 
wire w_mem_inst__abc_21203_new_n3620_; 
wire w_mem_inst__abc_21203_new_n3621_; 
wire w_mem_inst__abc_21203_new_n3622_; 
wire w_mem_inst__abc_21203_new_n3624_; 
wire w_mem_inst__abc_21203_new_n3625_; 
wire w_mem_inst__abc_21203_new_n3626_; 
wire w_mem_inst__abc_21203_new_n3627_; 
wire w_mem_inst__abc_21203_new_n3628_; 
wire w_mem_inst__abc_21203_new_n3630_; 
wire w_mem_inst__abc_21203_new_n3631_; 
wire w_mem_inst__abc_21203_new_n3632_; 
wire w_mem_inst__abc_21203_new_n3633_; 
wire w_mem_inst__abc_21203_new_n3634_; 
wire w_mem_inst__abc_21203_new_n3636_; 
wire w_mem_inst__abc_21203_new_n3637_; 
wire w_mem_inst__abc_21203_new_n3638_; 
wire w_mem_inst__abc_21203_new_n3639_; 
wire w_mem_inst__abc_21203_new_n3640_; 
wire w_mem_inst__abc_21203_new_n3642_; 
wire w_mem_inst__abc_21203_new_n3643_; 
wire w_mem_inst__abc_21203_new_n3644_; 
wire w_mem_inst__abc_21203_new_n3645_; 
wire w_mem_inst__abc_21203_new_n3646_; 
wire w_mem_inst__abc_21203_new_n3648_; 
wire w_mem_inst__abc_21203_new_n3649_; 
wire w_mem_inst__abc_21203_new_n3650_; 
wire w_mem_inst__abc_21203_new_n3651_; 
wire w_mem_inst__abc_21203_new_n3652_; 
wire w_mem_inst__abc_21203_new_n3654_; 
wire w_mem_inst__abc_21203_new_n3655_; 
wire w_mem_inst__abc_21203_new_n3656_; 
wire w_mem_inst__abc_21203_new_n3657_; 
wire w_mem_inst__abc_21203_new_n3658_; 
wire w_mem_inst__abc_21203_new_n3660_; 
wire w_mem_inst__abc_21203_new_n3661_; 
wire w_mem_inst__abc_21203_new_n3662_; 
wire w_mem_inst__abc_21203_new_n3663_; 
wire w_mem_inst__abc_21203_new_n3664_; 
wire w_mem_inst__abc_21203_new_n3666_; 
wire w_mem_inst__abc_21203_new_n3667_; 
wire w_mem_inst__abc_21203_new_n3668_; 
wire w_mem_inst__abc_21203_new_n3669_; 
wire w_mem_inst__abc_21203_new_n3670_; 
wire w_mem_inst__abc_21203_new_n3672_; 
wire w_mem_inst__abc_21203_new_n3673_; 
wire w_mem_inst__abc_21203_new_n3674_; 
wire w_mem_inst__abc_21203_new_n3675_; 
wire w_mem_inst__abc_21203_new_n3676_; 
wire w_mem_inst__abc_21203_new_n3678_; 
wire w_mem_inst__abc_21203_new_n3679_; 
wire w_mem_inst__abc_21203_new_n3680_; 
wire w_mem_inst__abc_21203_new_n3681_; 
wire w_mem_inst__abc_21203_new_n3682_; 
wire w_mem_inst__abc_21203_new_n3684_; 
wire w_mem_inst__abc_21203_new_n3685_; 
wire w_mem_inst__abc_21203_new_n3686_; 
wire w_mem_inst__abc_21203_new_n3687_; 
wire w_mem_inst__abc_21203_new_n3688_; 
wire w_mem_inst__abc_21203_new_n3690_; 
wire w_mem_inst__abc_21203_new_n3691_; 
wire w_mem_inst__abc_21203_new_n3692_; 
wire w_mem_inst__abc_21203_new_n3693_; 
wire w_mem_inst__abc_21203_new_n3694_; 
wire w_mem_inst__abc_21203_new_n3696_; 
wire w_mem_inst__abc_21203_new_n3697_; 
wire w_mem_inst__abc_21203_new_n3698_; 
wire w_mem_inst__abc_21203_new_n3699_; 
wire w_mem_inst__abc_21203_new_n3700_; 
wire w_mem_inst__abc_21203_new_n3702_; 
wire w_mem_inst__abc_21203_new_n3703_; 
wire w_mem_inst__abc_21203_new_n3704_; 
wire w_mem_inst__abc_21203_new_n3705_; 
wire w_mem_inst__abc_21203_new_n3706_; 
wire w_mem_inst__abc_21203_new_n3708_; 
wire w_mem_inst__abc_21203_new_n3709_; 
wire w_mem_inst__abc_21203_new_n3710_; 
wire w_mem_inst__abc_21203_new_n3711_; 
wire w_mem_inst__abc_21203_new_n3712_; 
wire w_mem_inst__abc_21203_new_n3714_; 
wire w_mem_inst__abc_21203_new_n3715_; 
wire w_mem_inst__abc_21203_new_n3716_; 
wire w_mem_inst__abc_21203_new_n3717_; 
wire w_mem_inst__abc_21203_new_n3718_; 
wire w_mem_inst__abc_21203_new_n3720_; 
wire w_mem_inst__abc_21203_new_n3721_; 
wire w_mem_inst__abc_21203_new_n3722_; 
wire w_mem_inst__abc_21203_new_n3723_; 
wire w_mem_inst__abc_21203_new_n3724_; 
wire w_mem_inst__abc_21203_new_n3726_; 
wire w_mem_inst__abc_21203_new_n3727_; 
wire w_mem_inst__abc_21203_new_n3728_; 
wire w_mem_inst__abc_21203_new_n3729_; 
wire w_mem_inst__abc_21203_new_n3730_; 
wire w_mem_inst__abc_21203_new_n3732_; 
wire w_mem_inst__abc_21203_new_n3733_; 
wire w_mem_inst__abc_21203_new_n3734_; 
wire w_mem_inst__abc_21203_new_n3735_; 
wire w_mem_inst__abc_21203_new_n3736_; 
wire w_mem_inst__abc_21203_new_n3738_; 
wire w_mem_inst__abc_21203_new_n3739_; 
wire w_mem_inst__abc_21203_new_n3740_; 
wire w_mem_inst__abc_21203_new_n3741_; 
wire w_mem_inst__abc_21203_new_n3742_; 
wire w_mem_inst__abc_21203_new_n3744_; 
wire w_mem_inst__abc_21203_new_n3745_; 
wire w_mem_inst__abc_21203_new_n3746_; 
wire w_mem_inst__abc_21203_new_n3747_; 
wire w_mem_inst__abc_21203_new_n3748_; 
wire w_mem_inst__abc_21203_new_n3750_; 
wire w_mem_inst__abc_21203_new_n3751_; 
wire w_mem_inst__abc_21203_new_n3752_; 
wire w_mem_inst__abc_21203_new_n3753_; 
wire w_mem_inst__abc_21203_new_n3754_; 
wire w_mem_inst__abc_21203_new_n3756_; 
wire w_mem_inst__abc_21203_new_n3757_; 
wire w_mem_inst__abc_21203_new_n3758_; 
wire w_mem_inst__abc_21203_new_n3759_; 
wire w_mem_inst__abc_21203_new_n3760_; 
wire w_mem_inst__abc_21203_new_n3762_; 
wire w_mem_inst__abc_21203_new_n3763_; 
wire w_mem_inst__abc_21203_new_n3764_; 
wire w_mem_inst__abc_21203_new_n3765_; 
wire w_mem_inst__abc_21203_new_n3766_; 
wire w_mem_inst__abc_21203_new_n3768_; 
wire w_mem_inst__abc_21203_new_n3769_; 
wire w_mem_inst__abc_21203_new_n3770_; 
wire w_mem_inst__abc_21203_new_n3771_; 
wire w_mem_inst__abc_21203_new_n3772_; 
wire w_mem_inst__abc_21203_new_n3774_; 
wire w_mem_inst__abc_21203_new_n3775_; 
wire w_mem_inst__abc_21203_new_n3776_; 
wire w_mem_inst__abc_21203_new_n3777_; 
wire w_mem_inst__abc_21203_new_n3778_; 
wire w_mem_inst__abc_21203_new_n3780_; 
wire w_mem_inst__abc_21203_new_n3781_; 
wire w_mem_inst__abc_21203_new_n3782_; 
wire w_mem_inst__abc_21203_new_n3783_; 
wire w_mem_inst__abc_21203_new_n3784_; 
wire w_mem_inst__abc_21203_new_n3786_; 
wire w_mem_inst__abc_21203_new_n3787_; 
wire w_mem_inst__abc_21203_new_n3788_; 
wire w_mem_inst__abc_21203_new_n3789_; 
wire w_mem_inst__abc_21203_new_n3790_; 
wire w_mem_inst__abc_21203_new_n3792_; 
wire w_mem_inst__abc_21203_new_n3793_; 
wire w_mem_inst__abc_21203_new_n3794_; 
wire w_mem_inst__abc_21203_new_n3795_; 
wire w_mem_inst__abc_21203_new_n3796_; 
wire w_mem_inst__abc_21203_new_n3798_; 
wire w_mem_inst__abc_21203_new_n3799_; 
wire w_mem_inst__abc_21203_new_n3800_; 
wire w_mem_inst__abc_21203_new_n3801_; 
wire w_mem_inst__abc_21203_new_n3802_; 
wire w_mem_inst__abc_21203_new_n3804_; 
wire w_mem_inst__abc_21203_new_n3805_; 
wire w_mem_inst__abc_21203_new_n3806_; 
wire w_mem_inst__abc_21203_new_n3807_; 
wire w_mem_inst__abc_21203_new_n3808_; 
wire w_mem_inst__abc_21203_new_n3810_; 
wire w_mem_inst__abc_21203_new_n3811_; 
wire w_mem_inst__abc_21203_new_n3812_; 
wire w_mem_inst__abc_21203_new_n3813_; 
wire w_mem_inst__abc_21203_new_n3814_; 
wire w_mem_inst__abc_21203_new_n3816_; 
wire w_mem_inst__abc_21203_new_n3817_; 
wire w_mem_inst__abc_21203_new_n3818_; 
wire w_mem_inst__abc_21203_new_n3819_; 
wire w_mem_inst__abc_21203_new_n3820_; 
wire w_mem_inst__abc_21203_new_n3822_; 
wire w_mem_inst__abc_21203_new_n3823_; 
wire w_mem_inst__abc_21203_new_n3824_; 
wire w_mem_inst__abc_21203_new_n3825_; 
wire w_mem_inst__abc_21203_new_n3826_; 
wire w_mem_inst__abc_21203_new_n3828_; 
wire w_mem_inst__abc_21203_new_n3829_; 
wire w_mem_inst__abc_21203_new_n3830_; 
wire w_mem_inst__abc_21203_new_n3831_; 
wire w_mem_inst__abc_21203_new_n3832_; 
wire w_mem_inst__abc_21203_new_n3834_; 
wire w_mem_inst__abc_21203_new_n3835_; 
wire w_mem_inst__abc_21203_new_n3836_; 
wire w_mem_inst__abc_21203_new_n3837_; 
wire w_mem_inst__abc_21203_new_n3838_; 
wire w_mem_inst__abc_21203_new_n3840_; 
wire w_mem_inst__abc_21203_new_n3841_; 
wire w_mem_inst__abc_21203_new_n3842_; 
wire w_mem_inst__abc_21203_new_n3843_; 
wire w_mem_inst__abc_21203_new_n3844_; 
wire w_mem_inst__abc_21203_new_n3846_; 
wire w_mem_inst__abc_21203_new_n3847_; 
wire w_mem_inst__abc_21203_new_n3848_; 
wire w_mem_inst__abc_21203_new_n3849_; 
wire w_mem_inst__abc_21203_new_n3850_; 
wire w_mem_inst__abc_21203_new_n3852_; 
wire w_mem_inst__abc_21203_new_n3853_; 
wire w_mem_inst__abc_21203_new_n3854_; 
wire w_mem_inst__abc_21203_new_n3855_; 
wire w_mem_inst__abc_21203_new_n3856_; 
wire w_mem_inst__abc_21203_new_n3858_; 
wire w_mem_inst__abc_21203_new_n3859_; 
wire w_mem_inst__abc_21203_new_n3860_; 
wire w_mem_inst__abc_21203_new_n3861_; 
wire w_mem_inst__abc_21203_new_n3862_; 
wire w_mem_inst__abc_21203_new_n3864_; 
wire w_mem_inst__abc_21203_new_n3865_; 
wire w_mem_inst__abc_21203_new_n3866_; 
wire w_mem_inst__abc_21203_new_n3867_; 
wire w_mem_inst__abc_21203_new_n3868_; 
wire w_mem_inst__abc_21203_new_n3870_; 
wire w_mem_inst__abc_21203_new_n3871_; 
wire w_mem_inst__abc_21203_new_n3872_; 
wire w_mem_inst__abc_21203_new_n3873_; 
wire w_mem_inst__abc_21203_new_n3874_; 
wire w_mem_inst__abc_21203_new_n3876_; 
wire w_mem_inst__abc_21203_new_n3877_; 
wire w_mem_inst__abc_21203_new_n3878_; 
wire w_mem_inst__abc_21203_new_n3879_; 
wire w_mem_inst__abc_21203_new_n3880_; 
wire w_mem_inst__abc_21203_new_n3882_; 
wire w_mem_inst__abc_21203_new_n3883_; 
wire w_mem_inst__abc_21203_new_n3884_; 
wire w_mem_inst__abc_21203_new_n3885_; 
wire w_mem_inst__abc_21203_new_n3886_; 
wire w_mem_inst__abc_21203_new_n3888_; 
wire w_mem_inst__abc_21203_new_n3889_; 
wire w_mem_inst__abc_21203_new_n3890_; 
wire w_mem_inst__abc_21203_new_n3891_; 
wire w_mem_inst__abc_21203_new_n3892_; 
wire w_mem_inst__abc_21203_new_n3894_; 
wire w_mem_inst__abc_21203_new_n3895_; 
wire w_mem_inst__abc_21203_new_n3896_; 
wire w_mem_inst__abc_21203_new_n3897_; 
wire w_mem_inst__abc_21203_new_n3898_; 
wire w_mem_inst__abc_21203_new_n3900_; 
wire w_mem_inst__abc_21203_new_n3901_; 
wire w_mem_inst__abc_21203_new_n3902_; 
wire w_mem_inst__abc_21203_new_n3903_; 
wire w_mem_inst__abc_21203_new_n3904_; 
wire w_mem_inst__abc_21203_new_n3906_; 
wire w_mem_inst__abc_21203_new_n3907_; 
wire w_mem_inst__abc_21203_new_n3908_; 
wire w_mem_inst__abc_21203_new_n3909_; 
wire w_mem_inst__abc_21203_new_n3910_; 
wire w_mem_inst__abc_21203_new_n3912_; 
wire w_mem_inst__abc_21203_new_n3913_; 
wire w_mem_inst__abc_21203_new_n3914_; 
wire w_mem_inst__abc_21203_new_n3915_; 
wire w_mem_inst__abc_21203_new_n3916_; 
wire w_mem_inst__abc_21203_new_n3918_; 
wire w_mem_inst__abc_21203_new_n3919_; 
wire w_mem_inst__abc_21203_new_n3920_; 
wire w_mem_inst__abc_21203_new_n3921_; 
wire w_mem_inst__abc_21203_new_n3922_; 
wire w_mem_inst__abc_21203_new_n3924_; 
wire w_mem_inst__abc_21203_new_n3925_; 
wire w_mem_inst__abc_21203_new_n3926_; 
wire w_mem_inst__abc_21203_new_n3927_; 
wire w_mem_inst__abc_21203_new_n3928_; 
wire w_mem_inst__abc_21203_new_n3930_; 
wire w_mem_inst__abc_21203_new_n3931_; 
wire w_mem_inst__abc_21203_new_n3932_; 
wire w_mem_inst__abc_21203_new_n3933_; 
wire w_mem_inst__abc_21203_new_n3934_; 
wire w_mem_inst__abc_21203_new_n3936_; 
wire w_mem_inst__abc_21203_new_n3937_; 
wire w_mem_inst__abc_21203_new_n3938_; 
wire w_mem_inst__abc_21203_new_n3939_; 
wire w_mem_inst__abc_21203_new_n3940_; 
wire w_mem_inst__abc_21203_new_n3942_; 
wire w_mem_inst__abc_21203_new_n3943_; 
wire w_mem_inst__abc_21203_new_n3944_; 
wire w_mem_inst__abc_21203_new_n3945_; 
wire w_mem_inst__abc_21203_new_n3946_; 
wire w_mem_inst__abc_21203_new_n3948_; 
wire w_mem_inst__abc_21203_new_n3949_; 
wire w_mem_inst__abc_21203_new_n3950_; 
wire w_mem_inst__abc_21203_new_n3951_; 
wire w_mem_inst__abc_21203_new_n3952_; 
wire w_mem_inst__abc_21203_new_n3954_; 
wire w_mem_inst__abc_21203_new_n3955_; 
wire w_mem_inst__abc_21203_new_n3956_; 
wire w_mem_inst__abc_21203_new_n3957_; 
wire w_mem_inst__abc_21203_new_n3958_; 
wire w_mem_inst__abc_21203_new_n3960_; 
wire w_mem_inst__abc_21203_new_n3961_; 
wire w_mem_inst__abc_21203_new_n3962_; 
wire w_mem_inst__abc_21203_new_n3963_; 
wire w_mem_inst__abc_21203_new_n3964_; 
wire w_mem_inst__abc_21203_new_n3966_; 
wire w_mem_inst__abc_21203_new_n3967_; 
wire w_mem_inst__abc_21203_new_n3968_; 
wire w_mem_inst__abc_21203_new_n3969_; 
wire w_mem_inst__abc_21203_new_n3970_; 
wire w_mem_inst__abc_21203_new_n3972_; 
wire w_mem_inst__abc_21203_new_n3973_; 
wire w_mem_inst__abc_21203_new_n3974_; 
wire w_mem_inst__abc_21203_new_n3975_; 
wire w_mem_inst__abc_21203_new_n3976_; 
wire w_mem_inst__abc_21203_new_n3978_; 
wire w_mem_inst__abc_21203_new_n3979_; 
wire w_mem_inst__abc_21203_new_n3980_; 
wire w_mem_inst__abc_21203_new_n3981_; 
wire w_mem_inst__abc_21203_new_n3982_; 
wire w_mem_inst__abc_21203_new_n3984_; 
wire w_mem_inst__abc_21203_new_n3985_; 
wire w_mem_inst__abc_21203_new_n3986_; 
wire w_mem_inst__abc_21203_new_n3987_; 
wire w_mem_inst__abc_21203_new_n3988_; 
wire w_mem_inst__abc_21203_new_n3990_; 
wire w_mem_inst__abc_21203_new_n3991_; 
wire w_mem_inst__abc_21203_new_n3992_; 
wire w_mem_inst__abc_21203_new_n3993_; 
wire w_mem_inst__abc_21203_new_n3994_; 
wire w_mem_inst__abc_21203_new_n3996_; 
wire w_mem_inst__abc_21203_new_n3997_; 
wire w_mem_inst__abc_21203_new_n3998_; 
wire w_mem_inst__abc_21203_new_n3999_; 
wire w_mem_inst__abc_21203_new_n4000_; 
wire w_mem_inst__abc_21203_new_n4002_; 
wire w_mem_inst__abc_21203_new_n4003_; 
wire w_mem_inst__abc_21203_new_n4004_; 
wire w_mem_inst__abc_21203_new_n4005_; 
wire w_mem_inst__abc_21203_new_n4006_; 
wire w_mem_inst__abc_21203_new_n4008_; 
wire w_mem_inst__abc_21203_new_n4009_; 
wire w_mem_inst__abc_21203_new_n4010_; 
wire w_mem_inst__abc_21203_new_n4011_; 
wire w_mem_inst__abc_21203_new_n4012_; 
wire w_mem_inst__abc_21203_new_n4014_; 
wire w_mem_inst__abc_21203_new_n4015_; 
wire w_mem_inst__abc_21203_new_n4016_; 
wire w_mem_inst__abc_21203_new_n4017_; 
wire w_mem_inst__abc_21203_new_n4018_; 
wire w_mem_inst__abc_21203_new_n4020_; 
wire w_mem_inst__abc_21203_new_n4021_; 
wire w_mem_inst__abc_21203_new_n4022_; 
wire w_mem_inst__abc_21203_new_n4023_; 
wire w_mem_inst__abc_21203_new_n4024_; 
wire w_mem_inst__abc_21203_new_n4026_; 
wire w_mem_inst__abc_21203_new_n4027_; 
wire w_mem_inst__abc_21203_new_n4028_; 
wire w_mem_inst__abc_21203_new_n4029_; 
wire w_mem_inst__abc_21203_new_n4030_; 
wire w_mem_inst__abc_21203_new_n4032_; 
wire w_mem_inst__abc_21203_new_n4033_; 
wire w_mem_inst__abc_21203_new_n4034_; 
wire w_mem_inst__abc_21203_new_n4035_; 
wire w_mem_inst__abc_21203_new_n4036_; 
wire w_mem_inst__abc_21203_new_n4038_; 
wire w_mem_inst__abc_21203_new_n4039_; 
wire w_mem_inst__abc_21203_new_n4040_; 
wire w_mem_inst__abc_21203_new_n4041_; 
wire w_mem_inst__abc_21203_new_n4042_; 
wire w_mem_inst__abc_21203_new_n4044_; 
wire w_mem_inst__abc_21203_new_n4045_; 
wire w_mem_inst__abc_21203_new_n4046_; 
wire w_mem_inst__abc_21203_new_n4047_; 
wire w_mem_inst__abc_21203_new_n4048_; 
wire w_mem_inst__abc_21203_new_n4050_; 
wire w_mem_inst__abc_21203_new_n4051_; 
wire w_mem_inst__abc_21203_new_n4052_; 
wire w_mem_inst__abc_21203_new_n4053_; 
wire w_mem_inst__abc_21203_new_n4054_; 
wire w_mem_inst__abc_21203_new_n4056_; 
wire w_mem_inst__abc_21203_new_n4057_; 
wire w_mem_inst__abc_21203_new_n4058_; 
wire w_mem_inst__abc_21203_new_n4059_; 
wire w_mem_inst__abc_21203_new_n4060_; 
wire w_mem_inst__abc_21203_new_n4062_; 
wire w_mem_inst__abc_21203_new_n4063_; 
wire w_mem_inst__abc_21203_new_n4064_; 
wire w_mem_inst__abc_21203_new_n4065_; 
wire w_mem_inst__abc_21203_new_n4066_; 
wire w_mem_inst__abc_21203_new_n4068_; 
wire w_mem_inst__abc_21203_new_n4069_; 
wire w_mem_inst__abc_21203_new_n4070_; 
wire w_mem_inst__abc_21203_new_n4071_; 
wire w_mem_inst__abc_21203_new_n4072_; 
wire w_mem_inst__abc_21203_new_n4074_; 
wire w_mem_inst__abc_21203_new_n4075_; 
wire w_mem_inst__abc_21203_new_n4076_; 
wire w_mem_inst__abc_21203_new_n4077_; 
wire w_mem_inst__abc_21203_new_n4078_; 
wire w_mem_inst__abc_21203_new_n4080_; 
wire w_mem_inst__abc_21203_new_n4081_; 
wire w_mem_inst__abc_21203_new_n4082_; 
wire w_mem_inst__abc_21203_new_n4083_; 
wire w_mem_inst__abc_21203_new_n4084_; 
wire w_mem_inst__abc_21203_new_n4086_; 
wire w_mem_inst__abc_21203_new_n4087_; 
wire w_mem_inst__abc_21203_new_n4088_; 
wire w_mem_inst__abc_21203_new_n4089_; 
wire w_mem_inst__abc_21203_new_n4090_; 
wire w_mem_inst__abc_21203_new_n4092_; 
wire w_mem_inst__abc_21203_new_n4093_; 
wire w_mem_inst__abc_21203_new_n4094_; 
wire w_mem_inst__abc_21203_new_n4095_; 
wire w_mem_inst__abc_21203_new_n4096_; 
wire w_mem_inst__abc_21203_new_n4098_; 
wire w_mem_inst__abc_21203_new_n4099_; 
wire w_mem_inst__abc_21203_new_n4100_; 
wire w_mem_inst__abc_21203_new_n4101_; 
wire w_mem_inst__abc_21203_new_n4102_; 
wire w_mem_inst__abc_21203_new_n4104_; 
wire w_mem_inst__abc_21203_new_n4105_; 
wire w_mem_inst__abc_21203_new_n4106_; 
wire w_mem_inst__abc_21203_new_n4107_; 
wire w_mem_inst__abc_21203_new_n4108_; 
wire w_mem_inst__abc_21203_new_n4110_; 
wire w_mem_inst__abc_21203_new_n4111_; 
wire w_mem_inst__abc_21203_new_n4112_; 
wire w_mem_inst__abc_21203_new_n4113_; 
wire w_mem_inst__abc_21203_new_n4114_; 
wire w_mem_inst__abc_21203_new_n4116_; 
wire w_mem_inst__abc_21203_new_n4117_; 
wire w_mem_inst__abc_21203_new_n4118_; 
wire w_mem_inst__abc_21203_new_n4119_; 
wire w_mem_inst__abc_21203_new_n4120_; 
wire w_mem_inst__abc_21203_new_n4122_; 
wire w_mem_inst__abc_21203_new_n4123_; 
wire w_mem_inst__abc_21203_new_n4124_; 
wire w_mem_inst__abc_21203_new_n4125_; 
wire w_mem_inst__abc_21203_new_n4126_; 
wire w_mem_inst__abc_21203_new_n4128_; 
wire w_mem_inst__abc_21203_new_n4129_; 
wire w_mem_inst__abc_21203_new_n4130_; 
wire w_mem_inst__abc_21203_new_n4131_; 
wire w_mem_inst__abc_21203_new_n4132_; 
wire w_mem_inst__abc_21203_new_n4134_; 
wire w_mem_inst__abc_21203_new_n4135_; 
wire w_mem_inst__abc_21203_new_n4136_; 
wire w_mem_inst__abc_21203_new_n4137_; 
wire w_mem_inst__abc_21203_new_n4138_; 
wire w_mem_inst__abc_21203_new_n4140_; 
wire w_mem_inst__abc_21203_new_n4141_; 
wire w_mem_inst__abc_21203_new_n4142_; 
wire w_mem_inst__abc_21203_new_n4143_; 
wire w_mem_inst__abc_21203_new_n4144_; 
wire w_mem_inst__abc_21203_new_n4146_; 
wire w_mem_inst__abc_21203_new_n4147_; 
wire w_mem_inst__abc_21203_new_n4148_; 
wire w_mem_inst__abc_21203_new_n4149_; 
wire w_mem_inst__abc_21203_new_n4150_; 
wire w_mem_inst__abc_21203_new_n4152_; 
wire w_mem_inst__abc_21203_new_n4153_; 
wire w_mem_inst__abc_21203_new_n4154_; 
wire w_mem_inst__abc_21203_new_n4155_; 
wire w_mem_inst__abc_21203_new_n4156_; 
wire w_mem_inst__abc_21203_new_n4158_; 
wire w_mem_inst__abc_21203_new_n4159_; 
wire w_mem_inst__abc_21203_new_n4160_; 
wire w_mem_inst__abc_21203_new_n4161_; 
wire w_mem_inst__abc_21203_new_n4162_; 
wire w_mem_inst__abc_21203_new_n4164_; 
wire w_mem_inst__abc_21203_new_n4165_; 
wire w_mem_inst__abc_21203_new_n4166_; 
wire w_mem_inst__abc_21203_new_n4167_; 
wire w_mem_inst__abc_21203_new_n4168_; 
wire w_mem_inst__abc_21203_new_n4170_; 
wire w_mem_inst__abc_21203_new_n4171_; 
wire w_mem_inst__abc_21203_new_n4172_; 
wire w_mem_inst__abc_21203_new_n4173_; 
wire w_mem_inst__abc_21203_new_n4174_; 
wire w_mem_inst__abc_21203_new_n4176_; 
wire w_mem_inst__abc_21203_new_n4177_; 
wire w_mem_inst__abc_21203_new_n4178_; 
wire w_mem_inst__abc_21203_new_n4179_; 
wire w_mem_inst__abc_21203_new_n4180_; 
wire w_mem_inst__abc_21203_new_n4182_; 
wire w_mem_inst__abc_21203_new_n4183_; 
wire w_mem_inst__abc_21203_new_n4184_; 
wire w_mem_inst__abc_21203_new_n4185_; 
wire w_mem_inst__abc_21203_new_n4186_; 
wire w_mem_inst__abc_21203_new_n4188_; 
wire w_mem_inst__abc_21203_new_n4189_; 
wire w_mem_inst__abc_21203_new_n4190_; 
wire w_mem_inst__abc_21203_new_n4191_; 
wire w_mem_inst__abc_21203_new_n4192_; 
wire w_mem_inst__abc_21203_new_n4194_; 
wire w_mem_inst__abc_21203_new_n4195_; 
wire w_mem_inst__abc_21203_new_n4196_; 
wire w_mem_inst__abc_21203_new_n4197_; 
wire w_mem_inst__abc_21203_new_n4198_; 
wire w_mem_inst__abc_21203_new_n4200_; 
wire w_mem_inst__abc_21203_new_n4201_; 
wire w_mem_inst__abc_21203_new_n4202_; 
wire w_mem_inst__abc_21203_new_n4203_; 
wire w_mem_inst__abc_21203_new_n4204_; 
wire w_mem_inst__abc_21203_new_n4206_; 
wire w_mem_inst__abc_21203_new_n4207_; 
wire w_mem_inst__abc_21203_new_n4208_; 
wire w_mem_inst__abc_21203_new_n4209_; 
wire w_mem_inst__abc_21203_new_n4210_; 
wire w_mem_inst__abc_21203_new_n4212_; 
wire w_mem_inst__abc_21203_new_n4213_; 
wire w_mem_inst__abc_21203_new_n4214_; 
wire w_mem_inst__abc_21203_new_n4215_; 
wire w_mem_inst__abc_21203_new_n4216_; 
wire w_mem_inst__abc_21203_new_n4218_; 
wire w_mem_inst__abc_21203_new_n4219_; 
wire w_mem_inst__abc_21203_new_n4220_; 
wire w_mem_inst__abc_21203_new_n4221_; 
wire w_mem_inst__abc_21203_new_n4222_; 
wire w_mem_inst__abc_21203_new_n4224_; 
wire w_mem_inst__abc_21203_new_n4225_; 
wire w_mem_inst__abc_21203_new_n4226_; 
wire w_mem_inst__abc_21203_new_n4227_; 
wire w_mem_inst__abc_21203_new_n4228_; 
wire w_mem_inst__abc_21203_new_n4230_; 
wire w_mem_inst__abc_21203_new_n4231_; 
wire w_mem_inst__abc_21203_new_n4232_; 
wire w_mem_inst__abc_21203_new_n4233_; 
wire w_mem_inst__abc_21203_new_n4234_; 
wire w_mem_inst__abc_21203_new_n4236_; 
wire w_mem_inst__abc_21203_new_n4237_; 
wire w_mem_inst__abc_21203_new_n4238_; 
wire w_mem_inst__abc_21203_new_n4239_; 
wire w_mem_inst__abc_21203_new_n4240_; 
wire w_mem_inst__abc_21203_new_n4242_; 
wire w_mem_inst__abc_21203_new_n4243_; 
wire w_mem_inst__abc_21203_new_n4244_; 
wire w_mem_inst__abc_21203_new_n4245_; 
wire w_mem_inst__abc_21203_new_n4246_; 
wire w_mem_inst__abc_21203_new_n4248_; 
wire w_mem_inst__abc_21203_new_n4249_; 
wire w_mem_inst__abc_21203_new_n4250_; 
wire w_mem_inst__abc_21203_new_n4251_; 
wire w_mem_inst__abc_21203_new_n4252_; 
wire w_mem_inst__abc_21203_new_n4254_; 
wire w_mem_inst__abc_21203_new_n4255_; 
wire w_mem_inst__abc_21203_new_n4256_; 
wire w_mem_inst__abc_21203_new_n4257_; 
wire w_mem_inst__abc_21203_new_n4258_; 
wire w_mem_inst__abc_21203_new_n4260_; 
wire w_mem_inst__abc_21203_new_n4261_; 
wire w_mem_inst__abc_21203_new_n4262_; 
wire w_mem_inst__abc_21203_new_n4263_; 
wire w_mem_inst__abc_21203_new_n4264_; 
wire w_mem_inst__abc_21203_new_n4266_; 
wire w_mem_inst__abc_21203_new_n4267_; 
wire w_mem_inst__abc_21203_new_n4268_; 
wire w_mem_inst__abc_21203_new_n4269_; 
wire w_mem_inst__abc_21203_new_n4270_; 
wire w_mem_inst__abc_21203_new_n4272_; 
wire w_mem_inst__abc_21203_new_n4273_; 
wire w_mem_inst__abc_21203_new_n4274_; 
wire w_mem_inst__abc_21203_new_n4275_; 
wire w_mem_inst__abc_21203_new_n4276_; 
wire w_mem_inst__abc_21203_new_n4278_; 
wire w_mem_inst__abc_21203_new_n4279_; 
wire w_mem_inst__abc_21203_new_n4280_; 
wire w_mem_inst__abc_21203_new_n4281_; 
wire w_mem_inst__abc_21203_new_n4282_; 
wire w_mem_inst__abc_21203_new_n4284_; 
wire w_mem_inst__abc_21203_new_n4285_; 
wire w_mem_inst__abc_21203_new_n4286_; 
wire w_mem_inst__abc_21203_new_n4287_; 
wire w_mem_inst__abc_21203_new_n4288_; 
wire w_mem_inst__abc_21203_new_n4290_; 
wire w_mem_inst__abc_21203_new_n4291_; 
wire w_mem_inst__abc_21203_new_n4292_; 
wire w_mem_inst__abc_21203_new_n4293_; 
wire w_mem_inst__abc_21203_new_n4294_; 
wire w_mem_inst__abc_21203_new_n4296_; 
wire w_mem_inst__abc_21203_new_n4297_; 
wire w_mem_inst__abc_21203_new_n4298_; 
wire w_mem_inst__abc_21203_new_n4299_; 
wire w_mem_inst__abc_21203_new_n4300_; 
wire w_mem_inst__abc_21203_new_n4302_; 
wire w_mem_inst__abc_21203_new_n4303_; 
wire w_mem_inst__abc_21203_new_n4304_; 
wire w_mem_inst__abc_21203_new_n4305_; 
wire w_mem_inst__abc_21203_new_n4306_; 
wire w_mem_inst__abc_21203_new_n4308_; 
wire w_mem_inst__abc_21203_new_n4309_; 
wire w_mem_inst__abc_21203_new_n4310_; 
wire w_mem_inst__abc_21203_new_n4311_; 
wire w_mem_inst__abc_21203_new_n4312_; 
wire w_mem_inst__abc_21203_new_n4314_; 
wire w_mem_inst__abc_21203_new_n4315_; 
wire w_mem_inst__abc_21203_new_n4316_; 
wire w_mem_inst__abc_21203_new_n4317_; 
wire w_mem_inst__abc_21203_new_n4318_; 
wire w_mem_inst__abc_21203_new_n4320_; 
wire w_mem_inst__abc_21203_new_n4321_; 
wire w_mem_inst__abc_21203_new_n4322_; 
wire w_mem_inst__abc_21203_new_n4323_; 
wire w_mem_inst__abc_21203_new_n4324_; 
wire w_mem_inst__abc_21203_new_n4326_; 
wire w_mem_inst__abc_21203_new_n4327_; 
wire w_mem_inst__abc_21203_new_n4328_; 
wire w_mem_inst__abc_21203_new_n4329_; 
wire w_mem_inst__abc_21203_new_n4330_; 
wire w_mem_inst__abc_21203_new_n4332_; 
wire w_mem_inst__abc_21203_new_n4333_; 
wire w_mem_inst__abc_21203_new_n4334_; 
wire w_mem_inst__abc_21203_new_n4335_; 
wire w_mem_inst__abc_21203_new_n4336_; 
wire w_mem_inst__abc_21203_new_n4338_; 
wire w_mem_inst__abc_21203_new_n4339_; 
wire w_mem_inst__abc_21203_new_n4340_; 
wire w_mem_inst__abc_21203_new_n4341_; 
wire w_mem_inst__abc_21203_new_n4342_; 
wire w_mem_inst__abc_21203_new_n4344_; 
wire w_mem_inst__abc_21203_new_n4345_; 
wire w_mem_inst__abc_21203_new_n4346_; 
wire w_mem_inst__abc_21203_new_n4347_; 
wire w_mem_inst__abc_21203_new_n4348_; 
wire w_mem_inst__abc_21203_new_n4350_; 
wire w_mem_inst__abc_21203_new_n4351_; 
wire w_mem_inst__abc_21203_new_n4352_; 
wire w_mem_inst__abc_21203_new_n4353_; 
wire w_mem_inst__abc_21203_new_n4354_; 
wire w_mem_inst__abc_21203_new_n4356_; 
wire w_mem_inst__abc_21203_new_n4357_; 
wire w_mem_inst__abc_21203_new_n4358_; 
wire w_mem_inst__abc_21203_new_n4359_; 
wire w_mem_inst__abc_21203_new_n4360_; 
wire w_mem_inst__abc_21203_new_n4362_; 
wire w_mem_inst__abc_21203_new_n4363_; 
wire w_mem_inst__abc_21203_new_n4364_; 
wire w_mem_inst__abc_21203_new_n4365_; 
wire w_mem_inst__abc_21203_new_n4366_; 
wire w_mem_inst__abc_21203_new_n4368_; 
wire w_mem_inst__abc_21203_new_n4369_; 
wire w_mem_inst__abc_21203_new_n4370_; 
wire w_mem_inst__abc_21203_new_n4371_; 
wire w_mem_inst__abc_21203_new_n4372_; 
wire w_mem_inst__abc_21203_new_n4374_; 
wire w_mem_inst__abc_21203_new_n4375_; 
wire w_mem_inst__abc_21203_new_n4376_; 
wire w_mem_inst__abc_21203_new_n4377_; 
wire w_mem_inst__abc_21203_new_n4378_; 
wire w_mem_inst__abc_21203_new_n4380_; 
wire w_mem_inst__abc_21203_new_n4381_; 
wire w_mem_inst__abc_21203_new_n4382_; 
wire w_mem_inst__abc_21203_new_n4383_; 
wire w_mem_inst__abc_21203_new_n4384_; 
wire w_mem_inst__abc_21203_new_n4386_; 
wire w_mem_inst__abc_21203_new_n4387_; 
wire w_mem_inst__abc_21203_new_n4388_; 
wire w_mem_inst__abc_21203_new_n4389_; 
wire w_mem_inst__abc_21203_new_n4390_; 
wire w_mem_inst__abc_21203_new_n4392_; 
wire w_mem_inst__abc_21203_new_n4393_; 
wire w_mem_inst__abc_21203_new_n4394_; 
wire w_mem_inst__abc_21203_new_n4395_; 
wire w_mem_inst__abc_21203_new_n4396_; 
wire w_mem_inst__abc_21203_new_n4398_; 
wire w_mem_inst__abc_21203_new_n4399_; 
wire w_mem_inst__abc_21203_new_n4400_; 
wire w_mem_inst__abc_21203_new_n4401_; 
wire w_mem_inst__abc_21203_new_n4402_; 
wire w_mem_inst__abc_21203_new_n4404_; 
wire w_mem_inst__abc_21203_new_n4405_; 
wire w_mem_inst__abc_21203_new_n4406_; 
wire w_mem_inst__abc_21203_new_n4407_; 
wire w_mem_inst__abc_21203_new_n4408_; 
wire w_mem_inst__abc_21203_new_n4410_; 
wire w_mem_inst__abc_21203_new_n4411_; 
wire w_mem_inst__abc_21203_new_n4412_; 
wire w_mem_inst__abc_21203_new_n4413_; 
wire w_mem_inst__abc_21203_new_n4414_; 
wire w_mem_inst__abc_21203_new_n4416_; 
wire w_mem_inst__abc_21203_new_n4417_; 
wire w_mem_inst__abc_21203_new_n4418_; 
wire w_mem_inst__abc_21203_new_n4419_; 
wire w_mem_inst__abc_21203_new_n4420_; 
wire w_mem_inst__abc_21203_new_n4422_; 
wire w_mem_inst__abc_21203_new_n4423_; 
wire w_mem_inst__abc_21203_new_n4424_; 
wire w_mem_inst__abc_21203_new_n4425_; 
wire w_mem_inst__abc_21203_new_n4426_; 
wire w_mem_inst__abc_21203_new_n4428_; 
wire w_mem_inst__abc_21203_new_n4429_; 
wire w_mem_inst__abc_21203_new_n4430_; 
wire w_mem_inst__abc_21203_new_n4431_; 
wire w_mem_inst__abc_21203_new_n4432_; 
wire w_mem_inst__abc_21203_new_n4434_; 
wire w_mem_inst__abc_21203_new_n4435_; 
wire w_mem_inst__abc_21203_new_n4436_; 
wire w_mem_inst__abc_21203_new_n4437_; 
wire w_mem_inst__abc_21203_new_n4438_; 
wire w_mem_inst__abc_21203_new_n4440_; 
wire w_mem_inst__abc_21203_new_n4441_; 
wire w_mem_inst__abc_21203_new_n4442_; 
wire w_mem_inst__abc_21203_new_n4443_; 
wire w_mem_inst__abc_21203_new_n4444_; 
wire w_mem_inst__abc_21203_new_n4446_; 
wire w_mem_inst__abc_21203_new_n4447_; 
wire w_mem_inst__abc_21203_new_n4448_; 
wire w_mem_inst__abc_21203_new_n4449_; 
wire w_mem_inst__abc_21203_new_n4450_; 
wire w_mem_inst__abc_21203_new_n4452_; 
wire w_mem_inst__abc_21203_new_n4453_; 
wire w_mem_inst__abc_21203_new_n4454_; 
wire w_mem_inst__abc_21203_new_n4455_; 
wire w_mem_inst__abc_21203_new_n4456_; 
wire w_mem_inst__abc_21203_new_n4458_; 
wire w_mem_inst__abc_21203_new_n4459_; 
wire w_mem_inst__abc_21203_new_n4460_; 
wire w_mem_inst__abc_21203_new_n4461_; 
wire w_mem_inst__abc_21203_new_n4462_; 
wire w_mem_inst__abc_21203_new_n4464_; 
wire w_mem_inst__abc_21203_new_n4465_; 
wire w_mem_inst__abc_21203_new_n4466_; 
wire w_mem_inst__abc_21203_new_n4467_; 
wire w_mem_inst__abc_21203_new_n4468_; 
wire w_mem_inst__abc_21203_new_n4470_; 
wire w_mem_inst__abc_21203_new_n4471_; 
wire w_mem_inst__abc_21203_new_n4472_; 
wire w_mem_inst__abc_21203_new_n4473_; 
wire w_mem_inst__abc_21203_new_n4474_; 
wire w_mem_inst__abc_21203_new_n4476_; 
wire w_mem_inst__abc_21203_new_n4477_; 
wire w_mem_inst__abc_21203_new_n4478_; 
wire w_mem_inst__abc_21203_new_n4479_; 
wire w_mem_inst__abc_21203_new_n4480_; 
wire w_mem_inst__abc_21203_new_n4482_; 
wire w_mem_inst__abc_21203_new_n4483_; 
wire w_mem_inst__abc_21203_new_n4484_; 
wire w_mem_inst__abc_21203_new_n4485_; 
wire w_mem_inst__abc_21203_new_n4486_; 
wire w_mem_inst__abc_21203_new_n4488_; 
wire w_mem_inst__abc_21203_new_n4489_; 
wire w_mem_inst__abc_21203_new_n4490_; 
wire w_mem_inst__abc_21203_new_n4491_; 
wire w_mem_inst__abc_21203_new_n4492_; 
wire w_mem_inst__abc_21203_new_n4494_; 
wire w_mem_inst__abc_21203_new_n4495_; 
wire w_mem_inst__abc_21203_new_n4496_; 
wire w_mem_inst__abc_21203_new_n4497_; 
wire w_mem_inst__abc_21203_new_n4498_; 
wire w_mem_inst__abc_21203_new_n4500_; 
wire w_mem_inst__abc_21203_new_n4501_; 
wire w_mem_inst__abc_21203_new_n4502_; 
wire w_mem_inst__abc_21203_new_n4503_; 
wire w_mem_inst__abc_21203_new_n4504_; 
wire w_mem_inst__abc_21203_new_n4506_; 
wire w_mem_inst__abc_21203_new_n4507_; 
wire w_mem_inst__abc_21203_new_n4508_; 
wire w_mem_inst__abc_21203_new_n4509_; 
wire w_mem_inst__abc_21203_new_n4510_; 
wire w_mem_inst__abc_21203_new_n4512_; 
wire w_mem_inst__abc_21203_new_n4513_; 
wire w_mem_inst__abc_21203_new_n4514_; 
wire w_mem_inst__abc_21203_new_n4515_; 
wire w_mem_inst__abc_21203_new_n4516_; 
wire w_mem_inst__abc_21203_new_n4518_; 
wire w_mem_inst__abc_21203_new_n4519_; 
wire w_mem_inst__abc_21203_new_n4520_; 
wire w_mem_inst__abc_21203_new_n4521_; 
wire w_mem_inst__abc_21203_new_n4522_; 
wire w_mem_inst__abc_21203_new_n4524_; 
wire w_mem_inst__abc_21203_new_n4525_; 
wire w_mem_inst__abc_21203_new_n4526_; 
wire w_mem_inst__abc_21203_new_n4527_; 
wire w_mem_inst__abc_21203_new_n4528_; 
wire w_mem_inst__abc_21203_new_n4530_; 
wire w_mem_inst__abc_21203_new_n4531_; 
wire w_mem_inst__abc_21203_new_n4532_; 
wire w_mem_inst__abc_21203_new_n4533_; 
wire w_mem_inst__abc_21203_new_n4534_; 
wire w_mem_inst__abc_21203_new_n4536_; 
wire w_mem_inst__abc_21203_new_n4537_; 
wire w_mem_inst__abc_21203_new_n4538_; 
wire w_mem_inst__abc_21203_new_n4539_; 
wire w_mem_inst__abc_21203_new_n4540_; 
wire w_mem_inst__abc_21203_new_n4542_; 
wire w_mem_inst__abc_21203_new_n4543_; 
wire w_mem_inst__abc_21203_new_n4544_; 
wire w_mem_inst__abc_21203_new_n4545_; 
wire w_mem_inst__abc_21203_new_n4546_; 
wire w_mem_inst__abc_21203_new_n4548_; 
wire w_mem_inst__abc_21203_new_n4549_; 
wire w_mem_inst__abc_21203_new_n4550_; 
wire w_mem_inst__abc_21203_new_n4551_; 
wire w_mem_inst__abc_21203_new_n4552_; 
wire w_mem_inst__abc_21203_new_n4554_; 
wire w_mem_inst__abc_21203_new_n4555_; 
wire w_mem_inst__abc_21203_new_n4556_; 
wire w_mem_inst__abc_21203_new_n4557_; 
wire w_mem_inst__abc_21203_new_n4558_; 
wire w_mem_inst__abc_21203_new_n4560_; 
wire w_mem_inst__abc_21203_new_n4561_; 
wire w_mem_inst__abc_21203_new_n4562_; 
wire w_mem_inst__abc_21203_new_n4563_; 
wire w_mem_inst__abc_21203_new_n4564_; 
wire w_mem_inst__abc_21203_new_n4566_; 
wire w_mem_inst__abc_21203_new_n4567_; 
wire w_mem_inst__abc_21203_new_n4568_; 
wire w_mem_inst__abc_21203_new_n4569_; 
wire w_mem_inst__abc_21203_new_n4570_; 
wire w_mem_inst__abc_21203_new_n4572_; 
wire w_mem_inst__abc_21203_new_n4573_; 
wire w_mem_inst__abc_21203_new_n4574_; 
wire w_mem_inst__abc_21203_new_n4575_; 
wire w_mem_inst__abc_21203_new_n4576_; 
wire w_mem_inst__abc_21203_new_n4578_; 
wire w_mem_inst__abc_21203_new_n4579_; 
wire w_mem_inst__abc_21203_new_n4580_; 
wire w_mem_inst__abc_21203_new_n4581_; 
wire w_mem_inst__abc_21203_new_n4582_; 
wire w_mem_inst__abc_21203_new_n4584_; 
wire w_mem_inst__abc_21203_new_n4585_; 
wire w_mem_inst__abc_21203_new_n4586_; 
wire w_mem_inst__abc_21203_new_n4587_; 
wire w_mem_inst__abc_21203_new_n4588_; 
wire w_mem_inst__abc_21203_new_n4590_; 
wire w_mem_inst__abc_21203_new_n4591_; 
wire w_mem_inst__abc_21203_new_n4592_; 
wire w_mem_inst__abc_21203_new_n4593_; 
wire w_mem_inst__abc_21203_new_n4594_; 
wire w_mem_inst__abc_21203_new_n4596_; 
wire w_mem_inst__abc_21203_new_n4597_; 
wire w_mem_inst__abc_21203_new_n4598_; 
wire w_mem_inst__abc_21203_new_n4599_; 
wire w_mem_inst__abc_21203_new_n4600_; 
wire w_mem_inst__abc_21203_new_n4602_; 
wire w_mem_inst__abc_21203_new_n4603_; 
wire w_mem_inst__abc_21203_new_n4604_; 
wire w_mem_inst__abc_21203_new_n4605_; 
wire w_mem_inst__abc_21203_new_n4606_; 
wire w_mem_inst__abc_21203_new_n4608_; 
wire w_mem_inst__abc_21203_new_n4609_; 
wire w_mem_inst__abc_21203_new_n4610_; 
wire w_mem_inst__abc_21203_new_n4611_; 
wire w_mem_inst__abc_21203_new_n4612_; 
wire w_mem_inst__abc_21203_new_n4614_; 
wire w_mem_inst__abc_21203_new_n4615_; 
wire w_mem_inst__abc_21203_new_n4616_; 
wire w_mem_inst__abc_21203_new_n4617_; 
wire w_mem_inst__abc_21203_new_n4618_; 
wire w_mem_inst__abc_21203_new_n4620_; 
wire w_mem_inst__abc_21203_new_n4621_; 
wire w_mem_inst__abc_21203_new_n4622_; 
wire w_mem_inst__abc_21203_new_n4623_; 
wire w_mem_inst__abc_21203_new_n4624_; 
wire w_mem_inst__abc_21203_new_n4626_; 
wire w_mem_inst__abc_21203_new_n4627_; 
wire w_mem_inst__abc_21203_new_n4628_; 
wire w_mem_inst__abc_21203_new_n4629_; 
wire w_mem_inst__abc_21203_new_n4630_; 
wire w_mem_inst__abc_21203_new_n4632_; 
wire w_mem_inst__abc_21203_new_n4633_; 
wire w_mem_inst__abc_21203_new_n4634_; 
wire w_mem_inst__abc_21203_new_n4635_; 
wire w_mem_inst__abc_21203_new_n4636_; 
wire w_mem_inst__abc_21203_new_n4638_; 
wire w_mem_inst__abc_21203_new_n4639_; 
wire w_mem_inst__abc_21203_new_n4640_; 
wire w_mem_inst__abc_21203_new_n4641_; 
wire w_mem_inst__abc_21203_new_n4642_; 
wire w_mem_inst__abc_21203_new_n4644_; 
wire w_mem_inst__abc_21203_new_n4645_; 
wire w_mem_inst__abc_21203_new_n4646_; 
wire w_mem_inst__abc_21203_new_n4647_; 
wire w_mem_inst__abc_21203_new_n4648_; 
wire w_mem_inst__abc_21203_new_n4650_; 
wire w_mem_inst__abc_21203_new_n4651_; 
wire w_mem_inst__abc_21203_new_n4652_; 
wire w_mem_inst__abc_21203_new_n4653_; 
wire w_mem_inst__abc_21203_new_n4654_; 
wire w_mem_inst__abc_21203_new_n4656_; 
wire w_mem_inst__abc_21203_new_n4657_; 
wire w_mem_inst__abc_21203_new_n4658_; 
wire w_mem_inst__abc_21203_new_n4659_; 
wire w_mem_inst__abc_21203_new_n4660_; 
wire w_mem_inst__abc_21203_new_n4662_; 
wire w_mem_inst__abc_21203_new_n4663_; 
wire w_mem_inst__abc_21203_new_n4664_; 
wire w_mem_inst__abc_21203_new_n4665_; 
wire w_mem_inst__abc_21203_new_n4666_; 
wire w_mem_inst__abc_21203_new_n4668_; 
wire w_mem_inst__abc_21203_new_n4669_; 
wire w_mem_inst__abc_21203_new_n4670_; 
wire w_mem_inst__abc_21203_new_n4671_; 
wire w_mem_inst__abc_21203_new_n4672_; 
wire w_mem_inst__abc_21203_new_n4674_; 
wire w_mem_inst__abc_21203_new_n4675_; 
wire w_mem_inst__abc_21203_new_n4676_; 
wire w_mem_inst__abc_21203_new_n4677_; 
wire w_mem_inst__abc_21203_new_n4678_; 
wire w_mem_inst__abc_21203_new_n4680_; 
wire w_mem_inst__abc_21203_new_n4681_; 
wire w_mem_inst__abc_21203_new_n4682_; 
wire w_mem_inst__abc_21203_new_n4683_; 
wire w_mem_inst__abc_21203_new_n4684_; 
wire w_mem_inst__abc_21203_new_n4686_; 
wire w_mem_inst__abc_21203_new_n4687_; 
wire w_mem_inst__abc_21203_new_n4688_; 
wire w_mem_inst__abc_21203_new_n4689_; 
wire w_mem_inst__abc_21203_new_n4690_; 
wire w_mem_inst__abc_21203_new_n4692_; 
wire w_mem_inst__abc_21203_new_n4693_; 
wire w_mem_inst__abc_21203_new_n4694_; 
wire w_mem_inst__abc_21203_new_n4695_; 
wire w_mem_inst__abc_21203_new_n4696_; 
wire w_mem_inst__abc_21203_new_n4698_; 
wire w_mem_inst__abc_21203_new_n4699_; 
wire w_mem_inst__abc_21203_new_n4700_; 
wire w_mem_inst__abc_21203_new_n4701_; 
wire w_mem_inst__abc_21203_new_n4702_; 
wire w_mem_inst__abc_21203_new_n4704_; 
wire w_mem_inst__abc_21203_new_n4705_; 
wire w_mem_inst__abc_21203_new_n4706_; 
wire w_mem_inst__abc_21203_new_n4707_; 
wire w_mem_inst__abc_21203_new_n4708_; 
wire w_mem_inst__abc_21203_new_n4710_; 
wire w_mem_inst__abc_21203_new_n4711_; 
wire w_mem_inst__abc_21203_new_n4712_; 
wire w_mem_inst__abc_21203_new_n4713_; 
wire w_mem_inst__abc_21203_new_n4714_; 
wire w_mem_inst__abc_21203_new_n4716_; 
wire w_mem_inst__abc_21203_new_n4717_; 
wire w_mem_inst__abc_21203_new_n4718_; 
wire w_mem_inst__abc_21203_new_n4719_; 
wire w_mem_inst__abc_21203_new_n4720_; 
wire w_mem_inst__abc_21203_new_n4722_; 
wire w_mem_inst__abc_21203_new_n4723_; 
wire w_mem_inst__abc_21203_new_n4724_; 
wire w_mem_inst__abc_21203_new_n4725_; 
wire w_mem_inst__abc_21203_new_n4726_; 
wire w_mem_inst__abc_21203_new_n4728_; 
wire w_mem_inst__abc_21203_new_n4729_; 
wire w_mem_inst__abc_21203_new_n4730_; 
wire w_mem_inst__abc_21203_new_n4731_; 
wire w_mem_inst__abc_21203_new_n4732_; 
wire w_mem_inst__abc_21203_new_n4734_; 
wire w_mem_inst__abc_21203_new_n4735_; 
wire w_mem_inst__abc_21203_new_n4736_; 
wire w_mem_inst__abc_21203_new_n4737_; 
wire w_mem_inst__abc_21203_new_n4738_; 
wire w_mem_inst__abc_21203_new_n4740_; 
wire w_mem_inst__abc_21203_new_n4741_; 
wire w_mem_inst__abc_21203_new_n4742_; 
wire w_mem_inst__abc_21203_new_n4743_; 
wire w_mem_inst__abc_21203_new_n4744_; 
wire w_mem_inst__abc_21203_new_n4746_; 
wire w_mem_inst__abc_21203_new_n4747_; 
wire w_mem_inst__abc_21203_new_n4748_; 
wire w_mem_inst__abc_21203_new_n4749_; 
wire w_mem_inst__abc_21203_new_n4750_; 
wire w_mem_inst__abc_21203_new_n4752_; 
wire w_mem_inst__abc_21203_new_n4753_; 
wire w_mem_inst__abc_21203_new_n4754_; 
wire w_mem_inst__abc_21203_new_n4755_; 
wire w_mem_inst__abc_21203_new_n4756_; 
wire w_mem_inst__abc_21203_new_n4758_; 
wire w_mem_inst__abc_21203_new_n4759_; 
wire w_mem_inst__abc_21203_new_n4760_; 
wire w_mem_inst__abc_21203_new_n4761_; 
wire w_mem_inst__abc_21203_new_n4762_; 
wire w_mem_inst__abc_21203_new_n4764_; 
wire w_mem_inst__abc_21203_new_n4765_; 
wire w_mem_inst__abc_21203_new_n4766_; 
wire w_mem_inst__abc_21203_new_n4767_; 
wire w_mem_inst__abc_21203_new_n4768_; 
wire w_mem_inst__abc_21203_new_n4770_; 
wire w_mem_inst__abc_21203_new_n4771_; 
wire w_mem_inst__abc_21203_new_n4772_; 
wire w_mem_inst__abc_21203_new_n4773_; 
wire w_mem_inst__abc_21203_new_n4774_; 
wire w_mem_inst__abc_21203_new_n4776_; 
wire w_mem_inst__abc_21203_new_n4777_; 
wire w_mem_inst__abc_21203_new_n4778_; 
wire w_mem_inst__abc_21203_new_n4779_; 
wire w_mem_inst__abc_21203_new_n4780_; 
wire w_mem_inst__abc_21203_new_n4782_; 
wire w_mem_inst__abc_21203_new_n4783_; 
wire w_mem_inst__abc_21203_new_n4784_; 
wire w_mem_inst__abc_21203_new_n4785_; 
wire w_mem_inst__abc_21203_new_n4786_; 
wire w_mem_inst__abc_21203_new_n4788_; 
wire w_mem_inst__abc_21203_new_n4789_; 
wire w_mem_inst__abc_21203_new_n4790_; 
wire w_mem_inst__abc_21203_new_n4791_; 
wire w_mem_inst__abc_21203_new_n4792_; 
wire w_mem_inst__abc_21203_new_n4794_; 
wire w_mem_inst__abc_21203_new_n4795_; 
wire w_mem_inst__abc_21203_new_n4796_; 
wire w_mem_inst__abc_21203_new_n4797_; 
wire w_mem_inst__abc_21203_new_n4798_; 
wire w_mem_inst__abc_21203_new_n4800_; 
wire w_mem_inst__abc_21203_new_n4801_; 
wire w_mem_inst__abc_21203_new_n4802_; 
wire w_mem_inst__abc_21203_new_n4803_; 
wire w_mem_inst__abc_21203_new_n4804_; 
wire w_mem_inst__abc_21203_new_n4806_; 
wire w_mem_inst__abc_21203_new_n4807_; 
wire w_mem_inst__abc_21203_new_n4808_; 
wire w_mem_inst__abc_21203_new_n4809_; 
wire w_mem_inst__abc_21203_new_n4810_; 
wire w_mem_inst__abc_21203_new_n4812_; 
wire w_mem_inst__abc_21203_new_n4813_; 
wire w_mem_inst__abc_21203_new_n4814_; 
wire w_mem_inst__abc_21203_new_n4815_; 
wire w_mem_inst__abc_21203_new_n4816_; 
wire w_mem_inst__abc_21203_new_n4818_; 
wire w_mem_inst__abc_21203_new_n4819_; 
wire w_mem_inst__abc_21203_new_n4820_; 
wire w_mem_inst__abc_21203_new_n4821_; 
wire w_mem_inst__abc_21203_new_n4822_; 
wire w_mem_inst__abc_21203_new_n4824_; 
wire w_mem_inst__abc_21203_new_n4825_; 
wire w_mem_inst__abc_21203_new_n4826_; 
wire w_mem_inst__abc_21203_new_n4827_; 
wire w_mem_inst__abc_21203_new_n4828_; 
wire w_mem_inst__abc_21203_new_n4830_; 
wire w_mem_inst__abc_21203_new_n4831_; 
wire w_mem_inst__abc_21203_new_n4832_; 
wire w_mem_inst__abc_21203_new_n4833_; 
wire w_mem_inst__abc_21203_new_n4834_; 
wire w_mem_inst__abc_21203_new_n4836_; 
wire w_mem_inst__abc_21203_new_n4837_; 
wire w_mem_inst__abc_21203_new_n4838_; 
wire w_mem_inst__abc_21203_new_n4839_; 
wire w_mem_inst__abc_21203_new_n4840_; 
wire w_mem_inst__abc_21203_new_n4842_; 
wire w_mem_inst__abc_21203_new_n4843_; 
wire w_mem_inst__abc_21203_new_n4844_; 
wire w_mem_inst__abc_21203_new_n4845_; 
wire w_mem_inst__abc_21203_new_n4846_; 
wire w_mem_inst__abc_21203_new_n4848_; 
wire w_mem_inst__abc_21203_new_n4849_; 
wire w_mem_inst__abc_21203_new_n4850_; 
wire w_mem_inst__abc_21203_new_n4851_; 
wire w_mem_inst__abc_21203_new_n4852_; 
wire w_mem_inst__abc_21203_new_n4854_; 
wire w_mem_inst__abc_21203_new_n4855_; 
wire w_mem_inst__abc_21203_new_n4856_; 
wire w_mem_inst__abc_21203_new_n4857_; 
wire w_mem_inst__abc_21203_new_n4858_; 
wire w_mem_inst__abc_21203_new_n4860_; 
wire w_mem_inst__abc_21203_new_n4861_; 
wire w_mem_inst__abc_21203_new_n4862_; 
wire w_mem_inst__abc_21203_new_n4863_; 
wire w_mem_inst__abc_21203_new_n4864_; 
wire w_mem_inst__abc_21203_new_n4866_; 
wire w_mem_inst__abc_21203_new_n4867_; 
wire w_mem_inst__abc_21203_new_n4868_; 
wire w_mem_inst__abc_21203_new_n4869_; 
wire w_mem_inst__abc_21203_new_n4870_; 
wire w_mem_inst__abc_21203_new_n4872_; 
wire w_mem_inst__abc_21203_new_n4873_; 
wire w_mem_inst__abc_21203_new_n4874_; 
wire w_mem_inst__abc_21203_new_n4875_; 
wire w_mem_inst__abc_21203_new_n4876_; 
wire w_mem_inst__abc_21203_new_n4878_; 
wire w_mem_inst__abc_21203_new_n4879_; 
wire w_mem_inst__abc_21203_new_n4880_; 
wire w_mem_inst__abc_21203_new_n4881_; 
wire w_mem_inst__abc_21203_new_n4882_; 
wire w_mem_inst__abc_21203_new_n4884_; 
wire w_mem_inst__abc_21203_new_n4885_; 
wire w_mem_inst__abc_21203_new_n4886_; 
wire w_mem_inst__abc_21203_new_n4887_; 
wire w_mem_inst__abc_21203_new_n4888_; 
wire w_mem_inst__abc_21203_new_n4890_; 
wire w_mem_inst__abc_21203_new_n4891_; 
wire w_mem_inst__abc_21203_new_n4892_; 
wire w_mem_inst__abc_21203_new_n4893_; 
wire w_mem_inst__abc_21203_new_n4894_; 
wire w_mem_inst__abc_21203_new_n4896_; 
wire w_mem_inst__abc_21203_new_n4897_; 
wire w_mem_inst__abc_21203_new_n4898_; 
wire w_mem_inst__abc_21203_new_n4899_; 
wire w_mem_inst__abc_21203_new_n4900_; 
wire w_mem_inst__abc_21203_new_n4902_; 
wire w_mem_inst__abc_21203_new_n4903_; 
wire w_mem_inst__abc_21203_new_n4904_; 
wire w_mem_inst__abc_21203_new_n4905_; 
wire w_mem_inst__abc_21203_new_n4906_; 
wire w_mem_inst__abc_21203_new_n4908_; 
wire w_mem_inst__abc_21203_new_n4909_; 
wire w_mem_inst__abc_21203_new_n4910_; 
wire w_mem_inst__abc_21203_new_n4911_; 
wire w_mem_inst__abc_21203_new_n4912_; 
wire w_mem_inst__abc_21203_new_n4914_; 
wire w_mem_inst__abc_21203_new_n4915_; 
wire w_mem_inst__abc_21203_new_n4916_; 
wire w_mem_inst__abc_21203_new_n4917_; 
wire w_mem_inst__abc_21203_new_n4918_; 
wire w_mem_inst__abc_21203_new_n4920_; 
wire w_mem_inst__abc_21203_new_n4921_; 
wire w_mem_inst__abc_21203_new_n4922_; 
wire w_mem_inst__abc_21203_new_n4923_; 
wire w_mem_inst__abc_21203_new_n4924_; 
wire w_mem_inst__abc_21203_new_n4926_; 
wire w_mem_inst__abc_21203_new_n4927_; 
wire w_mem_inst__abc_21203_new_n4928_; 
wire w_mem_inst__abc_21203_new_n4929_; 
wire w_mem_inst__abc_21203_new_n4930_; 
wire w_mem_inst__abc_21203_new_n4932_; 
wire w_mem_inst__abc_21203_new_n4933_; 
wire w_mem_inst__abc_21203_new_n4934_; 
wire w_mem_inst__abc_21203_new_n4935_; 
wire w_mem_inst__abc_21203_new_n4936_; 
wire w_mem_inst__abc_21203_new_n4938_; 
wire w_mem_inst__abc_21203_new_n4939_; 
wire w_mem_inst__abc_21203_new_n4940_; 
wire w_mem_inst__abc_21203_new_n4941_; 
wire w_mem_inst__abc_21203_new_n4942_; 
wire w_mem_inst__abc_21203_new_n4944_; 
wire w_mem_inst__abc_21203_new_n4945_; 
wire w_mem_inst__abc_21203_new_n4946_; 
wire w_mem_inst__abc_21203_new_n4947_; 
wire w_mem_inst__abc_21203_new_n4948_; 
wire w_mem_inst__abc_21203_new_n4950_; 
wire w_mem_inst__abc_21203_new_n4951_; 
wire w_mem_inst__abc_21203_new_n4952_; 
wire w_mem_inst__abc_21203_new_n4953_; 
wire w_mem_inst__abc_21203_new_n4954_; 
wire w_mem_inst__abc_21203_new_n4956_; 
wire w_mem_inst__abc_21203_new_n4957_; 
wire w_mem_inst__abc_21203_new_n4958_; 
wire w_mem_inst__abc_21203_new_n4959_; 
wire w_mem_inst__abc_21203_new_n4960_; 
wire w_mem_inst__abc_21203_new_n4962_; 
wire w_mem_inst__abc_21203_new_n4963_; 
wire w_mem_inst__abc_21203_new_n4964_; 
wire w_mem_inst__abc_21203_new_n4965_; 
wire w_mem_inst__abc_21203_new_n4966_; 
wire w_mem_inst__abc_21203_new_n4968_; 
wire w_mem_inst__abc_21203_new_n4969_; 
wire w_mem_inst__abc_21203_new_n4970_; 
wire w_mem_inst__abc_21203_new_n4971_; 
wire w_mem_inst__abc_21203_new_n4972_; 
wire w_mem_inst__abc_21203_new_n4974_; 
wire w_mem_inst__abc_21203_new_n4975_; 
wire w_mem_inst__abc_21203_new_n4976_; 
wire w_mem_inst__abc_21203_new_n4977_; 
wire w_mem_inst__abc_21203_new_n4978_; 
wire w_mem_inst__abc_21203_new_n4980_; 
wire w_mem_inst__abc_21203_new_n4981_; 
wire w_mem_inst__abc_21203_new_n4982_; 
wire w_mem_inst__abc_21203_new_n4983_; 
wire w_mem_inst__abc_21203_new_n4984_; 
wire w_mem_inst__abc_21203_new_n4986_; 
wire w_mem_inst__abc_21203_new_n4987_; 
wire w_mem_inst__abc_21203_new_n4988_; 
wire w_mem_inst__abc_21203_new_n4989_; 
wire w_mem_inst__abc_21203_new_n4990_; 
wire w_mem_inst__abc_21203_new_n4992_; 
wire w_mem_inst__abc_21203_new_n4993_; 
wire w_mem_inst__abc_21203_new_n4994_; 
wire w_mem_inst__abc_21203_new_n4995_; 
wire w_mem_inst__abc_21203_new_n4996_; 
wire w_mem_inst__abc_21203_new_n4998_; 
wire w_mem_inst__abc_21203_new_n4999_; 
wire w_mem_inst__abc_21203_new_n5000_; 
wire w_mem_inst__abc_21203_new_n5001_; 
wire w_mem_inst__abc_21203_new_n5002_; 
wire w_mem_inst__abc_21203_new_n5004_; 
wire w_mem_inst__abc_21203_new_n5005_; 
wire w_mem_inst__abc_21203_new_n5006_; 
wire w_mem_inst__abc_21203_new_n5007_; 
wire w_mem_inst__abc_21203_new_n5008_; 
wire w_mem_inst__abc_21203_new_n5010_; 
wire w_mem_inst__abc_21203_new_n5011_; 
wire w_mem_inst__abc_21203_new_n5012_; 
wire w_mem_inst__abc_21203_new_n5013_; 
wire w_mem_inst__abc_21203_new_n5014_; 
wire w_mem_inst__abc_21203_new_n5016_; 
wire w_mem_inst__abc_21203_new_n5017_; 
wire w_mem_inst__abc_21203_new_n5018_; 
wire w_mem_inst__abc_21203_new_n5019_; 
wire w_mem_inst__abc_21203_new_n5020_; 
wire w_mem_inst__abc_21203_new_n5022_; 
wire w_mem_inst__abc_21203_new_n5023_; 
wire w_mem_inst__abc_21203_new_n5024_; 
wire w_mem_inst__abc_21203_new_n5025_; 
wire w_mem_inst__abc_21203_new_n5026_; 
wire w_mem_inst__abc_21203_new_n5028_; 
wire w_mem_inst__abc_21203_new_n5029_; 
wire w_mem_inst__abc_21203_new_n5030_; 
wire w_mem_inst__abc_21203_new_n5031_; 
wire w_mem_inst__abc_21203_new_n5032_; 
wire w_mem_inst__abc_21203_new_n5034_; 
wire w_mem_inst__abc_21203_new_n5035_; 
wire w_mem_inst__abc_21203_new_n5036_; 
wire w_mem_inst__abc_21203_new_n5037_; 
wire w_mem_inst__abc_21203_new_n5038_; 
wire w_mem_inst__abc_21203_new_n5040_; 
wire w_mem_inst__abc_21203_new_n5041_; 
wire w_mem_inst__abc_21203_new_n5042_; 
wire w_mem_inst__abc_21203_new_n5043_; 
wire w_mem_inst__abc_21203_new_n5044_; 
wire w_mem_inst__abc_21203_new_n5046_; 
wire w_mem_inst__abc_21203_new_n5047_; 
wire w_mem_inst__abc_21203_new_n5048_; 
wire w_mem_inst__abc_21203_new_n5049_; 
wire w_mem_inst__abc_21203_new_n5050_; 
wire w_mem_inst__abc_21203_new_n5052_; 
wire w_mem_inst__abc_21203_new_n5053_; 
wire w_mem_inst__abc_21203_new_n5054_; 
wire w_mem_inst__abc_21203_new_n5055_; 
wire w_mem_inst__abc_21203_new_n5056_; 
wire w_mem_inst__abc_21203_new_n5058_; 
wire w_mem_inst__abc_21203_new_n5059_; 
wire w_mem_inst__abc_21203_new_n5060_; 
wire w_mem_inst__abc_21203_new_n5061_; 
wire w_mem_inst__abc_21203_new_n5062_; 
wire w_mem_inst__abc_21203_new_n5064_; 
wire w_mem_inst__abc_21203_new_n5065_; 
wire w_mem_inst__abc_21203_new_n5066_; 
wire w_mem_inst__abc_21203_new_n5067_; 
wire w_mem_inst__abc_21203_new_n5068_; 
wire w_mem_inst__abc_21203_new_n5070_; 
wire w_mem_inst__abc_21203_new_n5071_; 
wire w_mem_inst__abc_21203_new_n5072_; 
wire w_mem_inst__abc_21203_new_n5073_; 
wire w_mem_inst__abc_21203_new_n5074_; 
wire w_mem_inst__abc_21203_new_n5076_; 
wire w_mem_inst__abc_21203_new_n5077_; 
wire w_mem_inst__abc_21203_new_n5078_; 
wire w_mem_inst__abc_21203_new_n5079_; 
wire w_mem_inst__abc_21203_new_n5080_; 
wire w_mem_inst__abc_21203_new_n5082_; 
wire w_mem_inst__abc_21203_new_n5083_; 
wire w_mem_inst__abc_21203_new_n5084_; 
wire w_mem_inst__abc_21203_new_n5085_; 
wire w_mem_inst__abc_21203_new_n5086_; 
wire w_mem_inst__abc_21203_new_n5088_; 
wire w_mem_inst__abc_21203_new_n5089_; 
wire w_mem_inst__abc_21203_new_n5090_; 
wire w_mem_inst__abc_21203_new_n5091_; 
wire w_mem_inst__abc_21203_new_n5092_; 
wire w_mem_inst__abc_21203_new_n5094_; 
wire w_mem_inst__abc_21203_new_n5095_; 
wire w_mem_inst__abc_21203_new_n5096_; 
wire w_mem_inst__abc_21203_new_n5097_; 
wire w_mem_inst__abc_21203_new_n5098_; 
wire w_mem_inst__abc_21203_new_n5100_; 
wire w_mem_inst__abc_21203_new_n5101_; 
wire w_mem_inst__abc_21203_new_n5102_; 
wire w_mem_inst__abc_21203_new_n5103_; 
wire w_mem_inst__abc_21203_new_n5104_; 
wire w_mem_inst__abc_21203_new_n5106_; 
wire w_mem_inst__abc_21203_new_n5107_; 
wire w_mem_inst__abc_21203_new_n5108_; 
wire w_mem_inst__abc_21203_new_n5109_; 
wire w_mem_inst__abc_21203_new_n5110_; 
wire w_mem_inst__abc_21203_new_n5112_; 
wire w_mem_inst__abc_21203_new_n5113_; 
wire w_mem_inst__abc_21203_new_n5114_; 
wire w_mem_inst__abc_21203_new_n5115_; 
wire w_mem_inst__abc_21203_new_n5116_; 
wire w_mem_inst__abc_21203_new_n5118_; 
wire w_mem_inst__abc_21203_new_n5119_; 
wire w_mem_inst__abc_21203_new_n5120_; 
wire w_mem_inst__abc_21203_new_n5121_; 
wire w_mem_inst__abc_21203_new_n5122_; 
wire w_mem_inst__abc_21203_new_n5124_; 
wire w_mem_inst__abc_21203_new_n5125_; 
wire w_mem_inst__abc_21203_new_n5126_; 
wire w_mem_inst__abc_21203_new_n5127_; 
wire w_mem_inst__abc_21203_new_n5128_; 
wire w_mem_inst__abc_21203_new_n5130_; 
wire w_mem_inst__abc_21203_new_n5131_; 
wire w_mem_inst__abc_21203_new_n5132_; 
wire w_mem_inst__abc_21203_new_n5133_; 
wire w_mem_inst__abc_21203_new_n5134_; 
wire w_mem_inst__abc_21203_new_n5136_; 
wire w_mem_inst__abc_21203_new_n5137_; 
wire w_mem_inst__abc_21203_new_n5138_; 
wire w_mem_inst__abc_21203_new_n5139_; 
wire w_mem_inst__abc_21203_new_n5140_; 
wire w_mem_inst__abc_21203_new_n5142_; 
wire w_mem_inst__abc_21203_new_n5143_; 
wire w_mem_inst__abc_21203_new_n5144_; 
wire w_mem_inst__abc_21203_new_n5145_; 
wire w_mem_inst__abc_21203_new_n5146_; 
wire w_mem_inst__abc_21203_new_n5148_; 
wire w_mem_inst__abc_21203_new_n5149_; 
wire w_mem_inst__abc_21203_new_n5150_; 
wire w_mem_inst__abc_21203_new_n5151_; 
wire w_mem_inst__abc_21203_new_n5152_; 
wire w_mem_inst__abc_21203_new_n5154_; 
wire w_mem_inst__abc_21203_new_n5155_; 
wire w_mem_inst__abc_21203_new_n5156_; 
wire w_mem_inst__abc_21203_new_n5157_; 
wire w_mem_inst__abc_21203_new_n5158_; 
wire w_mem_inst__abc_21203_new_n5160_; 
wire w_mem_inst__abc_21203_new_n5161_; 
wire w_mem_inst__abc_21203_new_n5162_; 
wire w_mem_inst__abc_21203_new_n5163_; 
wire w_mem_inst__abc_21203_new_n5164_; 
wire w_mem_inst__abc_21203_new_n5166_; 
wire w_mem_inst__abc_21203_new_n5167_; 
wire w_mem_inst__abc_21203_new_n5168_; 
wire w_mem_inst__abc_21203_new_n5169_; 
wire w_mem_inst__abc_21203_new_n5170_; 
wire w_mem_inst__abc_21203_new_n5172_; 
wire w_mem_inst__abc_21203_new_n5173_; 
wire w_mem_inst__abc_21203_new_n5174_; 
wire w_mem_inst__abc_21203_new_n5175_; 
wire w_mem_inst__abc_21203_new_n5176_; 
wire w_mem_inst__abc_21203_new_n5178_; 
wire w_mem_inst__abc_21203_new_n5179_; 
wire w_mem_inst__abc_21203_new_n5180_; 
wire w_mem_inst__abc_21203_new_n5181_; 
wire w_mem_inst__abc_21203_new_n5182_; 
wire w_mem_inst__abc_21203_new_n5184_; 
wire w_mem_inst__abc_21203_new_n5185_; 
wire w_mem_inst__abc_21203_new_n5186_; 
wire w_mem_inst__abc_21203_new_n5187_; 
wire w_mem_inst__abc_21203_new_n5188_; 
wire w_mem_inst__abc_21203_new_n5190_; 
wire w_mem_inst__abc_21203_new_n5191_; 
wire w_mem_inst__abc_21203_new_n5192_; 
wire w_mem_inst__abc_21203_new_n5193_; 
wire w_mem_inst__abc_21203_new_n5194_; 
wire w_mem_inst__abc_21203_new_n5196_; 
wire w_mem_inst__abc_21203_new_n5197_; 
wire w_mem_inst__abc_21203_new_n5198_; 
wire w_mem_inst__abc_21203_new_n5199_; 
wire w_mem_inst__abc_21203_new_n5200_; 
wire w_mem_inst__abc_21203_new_n5202_; 
wire w_mem_inst__abc_21203_new_n5203_; 
wire w_mem_inst__abc_21203_new_n5204_; 
wire w_mem_inst__abc_21203_new_n5205_; 
wire w_mem_inst__abc_21203_new_n5206_; 
wire w_mem_inst__abc_21203_new_n5208_; 
wire w_mem_inst__abc_21203_new_n5209_; 
wire w_mem_inst__abc_21203_new_n5210_; 
wire w_mem_inst__abc_21203_new_n5211_; 
wire w_mem_inst__abc_21203_new_n5212_; 
wire w_mem_inst__abc_21203_new_n5214_; 
wire w_mem_inst__abc_21203_new_n5215_; 
wire w_mem_inst__abc_21203_new_n5216_; 
wire w_mem_inst__abc_21203_new_n5217_; 
wire w_mem_inst__abc_21203_new_n5218_; 
wire w_mem_inst__abc_21203_new_n5220_; 
wire w_mem_inst__abc_21203_new_n5221_; 
wire w_mem_inst__abc_21203_new_n5222_; 
wire w_mem_inst__abc_21203_new_n5223_; 
wire w_mem_inst__abc_21203_new_n5224_; 
wire w_mem_inst__abc_21203_new_n5226_; 
wire w_mem_inst__abc_21203_new_n5227_; 
wire w_mem_inst__abc_21203_new_n5228_; 
wire w_mem_inst__abc_21203_new_n5229_; 
wire w_mem_inst__abc_21203_new_n5230_; 
wire w_mem_inst__abc_21203_new_n5232_; 
wire w_mem_inst__abc_21203_new_n5233_; 
wire w_mem_inst__abc_21203_new_n5234_; 
wire w_mem_inst__abc_21203_new_n5235_; 
wire w_mem_inst__abc_21203_new_n5236_; 
wire w_mem_inst__abc_21203_new_n5238_; 
wire w_mem_inst__abc_21203_new_n5239_; 
wire w_mem_inst__abc_21203_new_n5240_; 
wire w_mem_inst__abc_21203_new_n5241_; 
wire w_mem_inst__abc_21203_new_n5242_; 
wire w_mem_inst__abc_21203_new_n5244_; 
wire w_mem_inst__abc_21203_new_n5245_; 
wire w_mem_inst__abc_21203_new_n5246_; 
wire w_mem_inst__abc_21203_new_n5247_; 
wire w_mem_inst__abc_21203_new_n5248_; 
wire w_mem_inst__abc_21203_new_n5250_; 
wire w_mem_inst__abc_21203_new_n5251_; 
wire w_mem_inst__abc_21203_new_n5252_; 
wire w_mem_inst__abc_21203_new_n5253_; 
wire w_mem_inst__abc_21203_new_n5254_; 
wire w_mem_inst__abc_21203_new_n5256_; 
wire w_mem_inst__abc_21203_new_n5257_; 
wire w_mem_inst__abc_21203_new_n5258_; 
wire w_mem_inst__abc_21203_new_n5259_; 
wire w_mem_inst__abc_21203_new_n5260_; 
wire w_mem_inst__abc_21203_new_n5262_; 
wire w_mem_inst__abc_21203_new_n5263_; 
wire w_mem_inst__abc_21203_new_n5264_; 
wire w_mem_inst__abc_21203_new_n5265_; 
wire w_mem_inst__abc_21203_new_n5266_; 
wire w_mem_inst__abc_21203_new_n5268_; 
wire w_mem_inst__abc_21203_new_n5269_; 
wire w_mem_inst__abc_21203_new_n5270_; 
wire w_mem_inst__abc_21203_new_n5271_; 
wire w_mem_inst__abc_21203_new_n5272_; 
wire w_mem_inst__abc_21203_new_n5274_; 
wire w_mem_inst__abc_21203_new_n5275_; 
wire w_mem_inst__abc_21203_new_n5276_; 
wire w_mem_inst__abc_21203_new_n5277_; 
wire w_mem_inst__abc_21203_new_n5278_; 
wire w_mem_inst__abc_21203_new_n5280_; 
wire w_mem_inst__abc_21203_new_n5281_; 
wire w_mem_inst__abc_21203_new_n5282_; 
wire w_mem_inst__abc_21203_new_n5283_; 
wire w_mem_inst__abc_21203_new_n5284_; 
wire w_mem_inst__abc_21203_new_n5286_; 
wire w_mem_inst__abc_21203_new_n5287_; 
wire w_mem_inst__abc_21203_new_n5288_; 
wire w_mem_inst__abc_21203_new_n5289_; 
wire w_mem_inst__abc_21203_new_n5290_; 
wire w_mem_inst__abc_21203_new_n5292_; 
wire w_mem_inst__abc_21203_new_n5293_; 
wire w_mem_inst__abc_21203_new_n5294_; 
wire w_mem_inst__abc_21203_new_n5295_; 
wire w_mem_inst__abc_21203_new_n5296_; 
wire w_mem_inst__abc_21203_new_n5298_; 
wire w_mem_inst__abc_21203_new_n5299_; 
wire w_mem_inst__abc_21203_new_n5300_; 
wire w_mem_inst__abc_21203_new_n5301_; 
wire w_mem_inst__abc_21203_new_n5302_; 
wire w_mem_inst__abc_21203_new_n5304_; 
wire w_mem_inst__abc_21203_new_n5305_; 
wire w_mem_inst__abc_21203_new_n5306_; 
wire w_mem_inst__abc_21203_new_n5307_; 
wire w_mem_inst__abc_21203_new_n5308_; 
wire w_mem_inst__abc_21203_new_n5310_; 
wire w_mem_inst__abc_21203_new_n5311_; 
wire w_mem_inst__abc_21203_new_n5312_; 
wire w_mem_inst__abc_21203_new_n5313_; 
wire w_mem_inst__abc_21203_new_n5314_; 
wire w_mem_inst__abc_21203_new_n5316_; 
wire w_mem_inst__abc_21203_new_n5317_; 
wire w_mem_inst__abc_21203_new_n5318_; 
wire w_mem_inst__abc_21203_new_n5319_; 
wire w_mem_inst__abc_21203_new_n5320_; 
wire w_mem_inst__abc_21203_new_n5322_; 
wire w_mem_inst__abc_21203_new_n5323_; 
wire w_mem_inst__abc_21203_new_n5324_; 
wire w_mem_inst__abc_21203_new_n5325_; 
wire w_mem_inst__abc_21203_new_n5326_; 
wire w_mem_inst__abc_21203_new_n5328_; 
wire w_mem_inst__abc_21203_new_n5329_; 
wire w_mem_inst__abc_21203_new_n5330_; 
wire w_mem_inst__abc_21203_new_n5331_; 
wire w_mem_inst__abc_21203_new_n5332_; 
wire w_mem_inst__abc_21203_new_n5334_; 
wire w_mem_inst__abc_21203_new_n5335_; 
wire w_mem_inst__abc_21203_new_n5336_; 
wire w_mem_inst__abc_21203_new_n5337_; 
wire w_mem_inst__abc_21203_new_n5338_; 
wire w_mem_inst__abc_21203_new_n5340_; 
wire w_mem_inst__abc_21203_new_n5341_; 
wire w_mem_inst__abc_21203_new_n5342_; 
wire w_mem_inst__abc_21203_new_n5343_; 
wire w_mem_inst__abc_21203_new_n5344_; 
wire w_mem_inst__abc_21203_new_n5346_; 
wire w_mem_inst__abc_21203_new_n5347_; 
wire w_mem_inst__abc_21203_new_n5348_; 
wire w_mem_inst__abc_21203_new_n5349_; 
wire w_mem_inst__abc_21203_new_n5350_; 
wire w_mem_inst__abc_21203_new_n5352_; 
wire w_mem_inst__abc_21203_new_n5353_; 
wire w_mem_inst__abc_21203_new_n5354_; 
wire w_mem_inst__abc_21203_new_n5355_; 
wire w_mem_inst__abc_21203_new_n5356_; 
wire w_mem_inst__abc_21203_new_n5358_; 
wire w_mem_inst__abc_21203_new_n5359_; 
wire w_mem_inst__abc_21203_new_n5360_; 
wire w_mem_inst__abc_21203_new_n5361_; 
wire w_mem_inst__abc_21203_new_n5362_; 
wire w_mem_inst__abc_21203_new_n5364_; 
wire w_mem_inst__abc_21203_new_n5365_; 
wire w_mem_inst__abc_21203_new_n5366_; 
wire w_mem_inst__abc_21203_new_n5367_; 
wire w_mem_inst__abc_21203_new_n5368_; 
wire w_mem_inst__abc_21203_new_n5370_; 
wire w_mem_inst__abc_21203_new_n5371_; 
wire w_mem_inst__abc_21203_new_n5372_; 
wire w_mem_inst__abc_21203_new_n5373_; 
wire w_mem_inst__abc_21203_new_n5374_; 
wire w_mem_inst__abc_21203_new_n5376_; 
wire w_mem_inst__abc_21203_new_n5377_; 
wire w_mem_inst__abc_21203_new_n5378_; 
wire w_mem_inst__abc_21203_new_n5379_; 
wire w_mem_inst__abc_21203_new_n5380_; 
wire w_mem_inst__abc_21203_new_n5382_; 
wire w_mem_inst__abc_21203_new_n5383_; 
wire w_mem_inst__abc_21203_new_n5384_; 
wire w_mem_inst__abc_21203_new_n5385_; 
wire w_mem_inst__abc_21203_new_n5386_; 
wire w_mem_inst__abc_21203_new_n5388_; 
wire w_mem_inst__abc_21203_new_n5389_; 
wire w_mem_inst__abc_21203_new_n5390_; 
wire w_mem_inst__abc_21203_new_n5391_; 
wire w_mem_inst__abc_21203_new_n5392_; 
wire w_mem_inst__abc_21203_new_n5394_; 
wire w_mem_inst__abc_21203_new_n5395_; 
wire w_mem_inst__abc_21203_new_n5396_; 
wire w_mem_inst__abc_21203_new_n5397_; 
wire w_mem_inst__abc_21203_new_n5398_; 
wire w_mem_inst__abc_21203_new_n5400_; 
wire w_mem_inst__abc_21203_new_n5401_; 
wire w_mem_inst__abc_21203_new_n5402_; 
wire w_mem_inst__abc_21203_new_n5403_; 
wire w_mem_inst__abc_21203_new_n5404_; 
wire w_mem_inst__abc_21203_new_n5406_; 
wire w_mem_inst__abc_21203_new_n5407_; 
wire w_mem_inst__abc_21203_new_n5408_; 
wire w_mem_inst__abc_21203_new_n5409_; 
wire w_mem_inst__abc_21203_new_n5410_; 
wire w_mem_inst__abc_21203_new_n5412_; 
wire w_mem_inst__abc_21203_new_n5413_; 
wire w_mem_inst__abc_21203_new_n5414_; 
wire w_mem_inst__abc_21203_new_n5415_; 
wire w_mem_inst__abc_21203_new_n5416_; 
wire w_mem_inst__abc_21203_new_n5418_; 
wire w_mem_inst__abc_21203_new_n5419_; 
wire w_mem_inst__abc_21203_new_n5420_; 
wire w_mem_inst__abc_21203_new_n5421_; 
wire w_mem_inst__abc_21203_new_n5422_; 
wire w_mem_inst__abc_21203_new_n5424_; 
wire w_mem_inst__abc_21203_new_n5425_; 
wire w_mem_inst__abc_21203_new_n5426_; 
wire w_mem_inst__abc_21203_new_n5427_; 
wire w_mem_inst__abc_21203_new_n5428_; 
wire w_mem_inst__abc_21203_new_n5430_; 
wire w_mem_inst__abc_21203_new_n5431_; 
wire w_mem_inst__abc_21203_new_n5432_; 
wire w_mem_inst__abc_21203_new_n5433_; 
wire w_mem_inst__abc_21203_new_n5434_; 
wire w_mem_inst__abc_21203_new_n5436_; 
wire w_mem_inst__abc_21203_new_n5437_; 
wire w_mem_inst__abc_21203_new_n5438_; 
wire w_mem_inst__abc_21203_new_n5439_; 
wire w_mem_inst__abc_21203_new_n5440_; 
wire w_mem_inst__abc_21203_new_n5442_; 
wire w_mem_inst__abc_21203_new_n5443_; 
wire w_mem_inst__abc_21203_new_n5444_; 
wire w_mem_inst__abc_21203_new_n5445_; 
wire w_mem_inst__abc_21203_new_n5446_; 
wire w_mem_inst__abc_21203_new_n5448_; 
wire w_mem_inst__abc_21203_new_n5449_; 
wire w_mem_inst__abc_21203_new_n5450_; 
wire w_mem_inst__abc_21203_new_n5451_; 
wire w_mem_inst__abc_21203_new_n5452_; 
wire w_mem_inst__abc_21203_new_n5454_; 
wire w_mem_inst__abc_21203_new_n5455_; 
wire w_mem_inst__abc_21203_new_n5456_; 
wire w_mem_inst__abc_21203_new_n5457_; 
wire w_mem_inst__abc_21203_new_n5458_; 
wire w_mem_inst__abc_21203_new_n5460_; 
wire w_mem_inst__abc_21203_new_n5461_; 
wire w_mem_inst__abc_21203_new_n5462_; 
wire w_mem_inst__abc_21203_new_n5463_; 
wire w_mem_inst__abc_21203_new_n5464_; 
wire w_mem_inst__abc_21203_new_n5466_; 
wire w_mem_inst__abc_21203_new_n5467_; 
wire w_mem_inst__abc_21203_new_n5468_; 
wire w_mem_inst__abc_21203_new_n5469_; 
wire w_mem_inst__abc_21203_new_n5470_; 
wire w_mem_inst__abc_21203_new_n5472_; 
wire w_mem_inst__abc_21203_new_n5473_; 
wire w_mem_inst__abc_21203_new_n5474_; 
wire w_mem_inst__abc_21203_new_n5475_; 
wire w_mem_inst__abc_21203_new_n5476_; 
wire w_mem_inst__abc_21203_new_n5478_; 
wire w_mem_inst__abc_21203_new_n5479_; 
wire w_mem_inst__abc_21203_new_n5480_; 
wire w_mem_inst__abc_21203_new_n5481_; 
wire w_mem_inst__abc_21203_new_n5482_; 
wire w_mem_inst__abc_21203_new_n5484_; 
wire w_mem_inst__abc_21203_new_n5485_; 
wire w_mem_inst__abc_21203_new_n5486_; 
wire w_mem_inst__abc_21203_new_n5487_; 
wire w_mem_inst__abc_21203_new_n5488_; 
wire w_mem_inst__abc_21203_new_n5490_; 
wire w_mem_inst__abc_21203_new_n5491_; 
wire w_mem_inst__abc_21203_new_n5492_; 
wire w_mem_inst__abc_21203_new_n5493_; 
wire w_mem_inst__abc_21203_new_n5494_; 
wire w_mem_inst__abc_21203_new_n5496_; 
wire w_mem_inst__abc_21203_new_n5497_; 
wire w_mem_inst__abc_21203_new_n5498_; 
wire w_mem_inst__abc_21203_new_n5499_; 
wire w_mem_inst__abc_21203_new_n5500_; 
wire w_mem_inst__abc_21203_new_n5502_; 
wire w_mem_inst__abc_21203_new_n5503_; 
wire w_mem_inst__abc_21203_new_n5504_; 
wire w_mem_inst__abc_21203_new_n5505_; 
wire w_mem_inst__abc_21203_new_n5506_; 
wire w_mem_inst__abc_21203_new_n5508_; 
wire w_mem_inst__abc_21203_new_n5509_; 
wire w_mem_inst__abc_21203_new_n5510_; 
wire w_mem_inst__abc_21203_new_n5511_; 
wire w_mem_inst__abc_21203_new_n5512_; 
wire w_mem_inst__abc_21203_new_n5514_; 
wire w_mem_inst__abc_21203_new_n5515_; 
wire w_mem_inst__abc_21203_new_n5516_; 
wire w_mem_inst__abc_21203_new_n5517_; 
wire w_mem_inst__abc_21203_new_n5518_; 
wire w_mem_inst__abc_21203_new_n5520_; 
wire w_mem_inst__abc_21203_new_n5521_; 
wire w_mem_inst__abc_21203_new_n5522_; 
wire w_mem_inst__abc_21203_new_n5523_; 
wire w_mem_inst__abc_21203_new_n5524_; 
wire w_mem_inst__abc_21203_new_n5526_; 
wire w_mem_inst__abc_21203_new_n5527_; 
wire w_mem_inst__abc_21203_new_n5528_; 
wire w_mem_inst__abc_21203_new_n5529_; 
wire w_mem_inst__abc_21203_new_n5530_; 
wire w_mem_inst__abc_21203_new_n5532_; 
wire w_mem_inst__abc_21203_new_n5533_; 
wire w_mem_inst__abc_21203_new_n5534_; 
wire w_mem_inst__abc_21203_new_n5535_; 
wire w_mem_inst__abc_21203_new_n5536_; 
wire w_mem_inst__abc_21203_new_n5538_; 
wire w_mem_inst__abc_21203_new_n5539_; 
wire w_mem_inst__abc_21203_new_n5540_; 
wire w_mem_inst__abc_21203_new_n5541_; 
wire w_mem_inst__abc_21203_new_n5542_; 
wire w_mem_inst__abc_21203_new_n5544_; 
wire w_mem_inst__abc_21203_new_n5545_; 
wire w_mem_inst__abc_21203_new_n5546_; 
wire w_mem_inst__abc_21203_new_n5547_; 
wire w_mem_inst__abc_21203_new_n5548_; 
wire w_mem_inst__abc_21203_new_n5550_; 
wire w_mem_inst__abc_21203_new_n5551_; 
wire w_mem_inst__abc_21203_new_n5552_; 
wire w_mem_inst__abc_21203_new_n5553_; 
wire w_mem_inst__abc_21203_new_n5554_; 
wire w_mem_inst__abc_21203_new_n5556_; 
wire w_mem_inst__abc_21203_new_n5557_; 
wire w_mem_inst__abc_21203_new_n5558_; 
wire w_mem_inst__abc_21203_new_n5559_; 
wire w_mem_inst__abc_21203_new_n5560_; 
wire w_mem_inst__abc_21203_new_n5562_; 
wire w_mem_inst__abc_21203_new_n5563_; 
wire w_mem_inst__abc_21203_new_n5564_; 
wire w_mem_inst__abc_21203_new_n5565_; 
wire w_mem_inst__abc_21203_new_n5566_; 
wire w_mem_inst__abc_21203_new_n5568_; 
wire w_mem_inst__abc_21203_new_n5569_; 
wire w_mem_inst__abc_21203_new_n5570_; 
wire w_mem_inst__abc_21203_new_n5571_; 
wire w_mem_inst__abc_21203_new_n5572_; 
wire w_mem_inst__abc_21203_new_n5574_; 
wire w_mem_inst__abc_21203_new_n5575_; 
wire w_mem_inst__abc_21203_new_n5576_; 
wire w_mem_inst__abc_21203_new_n5577_; 
wire w_mem_inst__abc_21203_new_n5578_; 
wire w_mem_inst__abc_21203_new_n5580_; 
wire w_mem_inst__abc_21203_new_n5581_; 
wire w_mem_inst__abc_21203_new_n5582_; 
wire w_mem_inst__abc_21203_new_n5583_; 
wire w_mem_inst__abc_21203_new_n5584_; 
wire w_mem_inst__abc_21203_new_n5586_; 
wire w_mem_inst__abc_21203_new_n5587_; 
wire w_mem_inst__abc_21203_new_n5588_; 
wire w_mem_inst__abc_21203_new_n5589_; 
wire w_mem_inst__abc_21203_new_n5590_; 
wire w_mem_inst__abc_21203_new_n5592_; 
wire w_mem_inst__abc_21203_new_n5593_; 
wire w_mem_inst__abc_21203_new_n5594_; 
wire w_mem_inst__abc_21203_new_n5595_; 
wire w_mem_inst__abc_21203_new_n5596_; 
wire w_mem_inst__abc_21203_new_n5598_; 
wire w_mem_inst__abc_21203_new_n5599_; 
wire w_mem_inst__abc_21203_new_n5600_; 
wire w_mem_inst__abc_21203_new_n5601_; 
wire w_mem_inst__abc_21203_new_n5602_; 
wire w_mem_inst__abc_21203_new_n5604_; 
wire w_mem_inst__abc_21203_new_n5605_; 
wire w_mem_inst__abc_21203_new_n5606_; 
wire w_mem_inst__abc_21203_new_n5607_; 
wire w_mem_inst__abc_21203_new_n5608_; 
wire w_mem_inst__abc_21203_new_n5610_; 
wire w_mem_inst__abc_21203_new_n5611_; 
wire w_mem_inst__abc_21203_new_n5612_; 
wire w_mem_inst__abc_21203_new_n5613_; 
wire w_mem_inst__abc_21203_new_n5614_; 
wire w_mem_inst__abc_21203_new_n5616_; 
wire w_mem_inst__abc_21203_new_n5617_; 
wire w_mem_inst__abc_21203_new_n5618_; 
wire w_mem_inst__abc_21203_new_n5619_; 
wire w_mem_inst__abc_21203_new_n5620_; 
wire w_mem_inst__abc_21203_new_n5622_; 
wire w_mem_inst__abc_21203_new_n5623_; 
wire w_mem_inst__abc_21203_new_n5624_; 
wire w_mem_inst__abc_21203_new_n5625_; 
wire w_mem_inst__abc_21203_new_n5626_; 
wire w_mem_inst__abc_21203_new_n5628_; 
wire w_mem_inst__abc_21203_new_n5629_; 
wire w_mem_inst__abc_21203_new_n5630_; 
wire w_mem_inst__abc_21203_new_n5631_; 
wire w_mem_inst__abc_21203_new_n5632_; 
wire w_mem_inst__abc_21203_new_n5634_; 
wire w_mem_inst__abc_21203_new_n5635_; 
wire w_mem_inst__abc_21203_new_n5636_; 
wire w_mem_inst__abc_21203_new_n5637_; 
wire w_mem_inst__abc_21203_new_n5638_; 
wire w_mem_inst__abc_21203_new_n5640_; 
wire w_mem_inst__abc_21203_new_n5641_; 
wire w_mem_inst__abc_21203_new_n5642_; 
wire w_mem_inst__abc_21203_new_n5643_; 
wire w_mem_inst__abc_21203_new_n5644_; 
wire w_mem_inst__abc_21203_new_n5646_; 
wire w_mem_inst__abc_21203_new_n5647_; 
wire w_mem_inst__abc_21203_new_n5648_; 
wire w_mem_inst__abc_21203_new_n5649_; 
wire w_mem_inst__abc_21203_new_n5650_; 
wire w_mem_inst__abc_21203_new_n5652_; 
wire w_mem_inst__abc_21203_new_n5653_; 
wire w_mem_inst__abc_21203_new_n5654_; 
wire w_mem_inst__abc_21203_new_n5655_; 
wire w_mem_inst__abc_21203_new_n5656_; 
wire w_mem_inst__abc_21203_new_n5658_; 
wire w_mem_inst__abc_21203_new_n5659_; 
wire w_mem_inst__abc_21203_new_n5660_; 
wire w_mem_inst__abc_21203_new_n5661_; 
wire w_mem_inst__abc_21203_new_n5662_; 
wire w_mem_inst__abc_21203_new_n5664_; 
wire w_mem_inst__abc_21203_new_n5665_; 
wire w_mem_inst__abc_21203_new_n5666_; 
wire w_mem_inst__abc_21203_new_n5667_; 
wire w_mem_inst__abc_21203_new_n5668_; 
wire w_mem_inst__abc_21203_new_n5670_; 
wire w_mem_inst__abc_21203_new_n5671_; 
wire w_mem_inst__abc_21203_new_n5672_; 
wire w_mem_inst__abc_21203_new_n5673_; 
wire w_mem_inst__abc_21203_new_n5674_; 
wire w_mem_inst__abc_21203_new_n5676_; 
wire w_mem_inst__abc_21203_new_n5677_; 
wire w_mem_inst__abc_21203_new_n5678_; 
wire w_mem_inst__abc_21203_new_n5679_; 
wire w_mem_inst__abc_21203_new_n5680_; 
wire w_mem_inst__abc_21203_new_n5682_; 
wire w_mem_inst__abc_21203_new_n5683_; 
wire w_mem_inst__abc_21203_new_n5684_; 
wire w_mem_inst__abc_21203_new_n5685_; 
wire w_mem_inst__abc_21203_new_n5686_; 
wire w_mem_inst__abc_21203_new_n5688_; 
wire w_mem_inst__abc_21203_new_n5689_; 
wire w_mem_inst__abc_21203_new_n5690_; 
wire w_mem_inst__abc_21203_new_n5691_; 
wire w_mem_inst__abc_21203_new_n5692_; 
wire w_mem_inst__abc_21203_new_n5694_; 
wire w_mem_inst__abc_21203_new_n5695_; 
wire w_mem_inst__abc_21203_new_n5696_; 
wire w_mem_inst__abc_21203_new_n5697_; 
wire w_mem_inst__abc_21203_new_n5698_; 
wire w_mem_inst__abc_21203_new_n5700_; 
wire w_mem_inst__abc_21203_new_n5701_; 
wire w_mem_inst__abc_21203_new_n5702_; 
wire w_mem_inst__abc_21203_new_n5703_; 
wire w_mem_inst__abc_21203_new_n5704_; 
wire w_mem_inst__abc_21203_new_n5706_; 
wire w_mem_inst__abc_21203_new_n5707_; 
wire w_mem_inst__abc_21203_new_n5708_; 
wire w_mem_inst__abc_21203_new_n5709_; 
wire w_mem_inst__abc_21203_new_n5710_; 
wire w_mem_inst__abc_21203_new_n5712_; 
wire w_mem_inst__abc_21203_new_n5713_; 
wire w_mem_inst__abc_21203_new_n5714_; 
wire w_mem_inst__abc_21203_new_n5715_; 
wire w_mem_inst__abc_21203_new_n5716_; 
wire w_mem_inst__abc_21203_new_n5718_; 
wire w_mem_inst__abc_21203_new_n5719_; 
wire w_mem_inst__abc_21203_new_n5720_; 
wire w_mem_inst__abc_21203_new_n5721_; 
wire w_mem_inst__abc_21203_new_n5722_; 
wire w_mem_inst__abc_21203_new_n5724_; 
wire w_mem_inst__abc_21203_new_n5725_; 
wire w_mem_inst__abc_21203_new_n5726_; 
wire w_mem_inst__abc_21203_new_n5727_; 
wire w_mem_inst__abc_21203_new_n5728_; 
wire w_mem_inst__abc_21203_new_n5730_; 
wire w_mem_inst__abc_21203_new_n5731_; 
wire w_mem_inst__abc_21203_new_n5732_; 
wire w_mem_inst__abc_21203_new_n5733_; 
wire w_mem_inst__abc_21203_new_n5734_; 
wire w_mem_inst__abc_21203_new_n5736_; 
wire w_mem_inst__abc_21203_new_n5737_; 
wire w_mem_inst__abc_21203_new_n5738_; 
wire w_mem_inst__abc_21203_new_n5739_; 
wire w_mem_inst__abc_21203_new_n5740_; 
wire w_mem_inst__abc_21203_new_n5742_; 
wire w_mem_inst__abc_21203_new_n5743_; 
wire w_mem_inst__abc_21203_new_n5744_; 
wire w_mem_inst__abc_21203_new_n5745_; 
wire w_mem_inst__abc_21203_new_n5746_; 
wire w_mem_inst__abc_21203_new_n5748_; 
wire w_mem_inst__abc_21203_new_n5749_; 
wire w_mem_inst__abc_21203_new_n5750_; 
wire w_mem_inst__abc_21203_new_n5751_; 
wire w_mem_inst__abc_21203_new_n5752_; 
wire w_mem_inst__abc_21203_new_n5754_; 
wire w_mem_inst__abc_21203_new_n5755_; 
wire w_mem_inst__abc_21203_new_n5756_; 
wire w_mem_inst__abc_21203_new_n5757_; 
wire w_mem_inst__abc_21203_new_n5758_; 
wire w_mem_inst__abc_21203_new_n5760_; 
wire w_mem_inst__abc_21203_new_n5761_; 
wire w_mem_inst__abc_21203_new_n5762_; 
wire w_mem_inst__abc_21203_new_n5763_; 
wire w_mem_inst__abc_21203_new_n5764_; 
wire w_mem_inst__abc_21203_new_n5766_; 
wire w_mem_inst__abc_21203_new_n5767_; 
wire w_mem_inst__abc_21203_new_n5768_; 
wire w_mem_inst__abc_21203_new_n5769_; 
wire w_mem_inst__abc_21203_new_n5770_; 
wire w_mem_inst__abc_21203_new_n5772_; 
wire w_mem_inst__abc_21203_new_n5773_; 
wire w_mem_inst__abc_21203_new_n5774_; 
wire w_mem_inst__abc_21203_new_n5775_; 
wire w_mem_inst__abc_21203_new_n5776_; 
wire w_mem_inst__abc_21203_new_n5778_; 
wire w_mem_inst__abc_21203_new_n5779_; 
wire w_mem_inst__abc_21203_new_n5780_; 
wire w_mem_inst__abc_21203_new_n5781_; 
wire w_mem_inst__abc_21203_new_n5782_; 
wire w_mem_inst__abc_21203_new_n5784_; 
wire w_mem_inst__abc_21203_new_n5785_; 
wire w_mem_inst__abc_21203_new_n5786_; 
wire w_mem_inst__abc_21203_new_n5787_; 
wire w_mem_inst__abc_21203_new_n5788_; 
wire w_mem_inst__abc_21203_new_n5790_; 
wire w_mem_inst__abc_21203_new_n5791_; 
wire w_mem_inst__abc_21203_new_n5792_; 
wire w_mem_inst__abc_21203_new_n5793_; 
wire w_mem_inst__abc_21203_new_n5794_; 
wire w_mem_inst__abc_21203_new_n5796_; 
wire w_mem_inst__abc_21203_new_n5797_; 
wire w_mem_inst__abc_21203_new_n5798_; 
wire w_mem_inst__abc_21203_new_n5799_; 
wire w_mem_inst__abc_21203_new_n5800_; 
wire w_mem_inst__abc_21203_new_n5802_; 
wire w_mem_inst__abc_21203_new_n5803_; 
wire w_mem_inst__abc_21203_new_n5804_; 
wire w_mem_inst__abc_21203_new_n5805_; 
wire w_mem_inst__abc_21203_new_n5806_; 
wire w_mem_inst__abc_21203_new_n5808_; 
wire w_mem_inst__abc_21203_new_n5809_; 
wire w_mem_inst__abc_21203_new_n5810_; 
wire w_mem_inst__abc_21203_new_n5811_; 
wire w_mem_inst__abc_21203_new_n5812_; 
wire w_mem_inst__abc_21203_new_n5814_; 
wire w_mem_inst__abc_21203_new_n5815_; 
wire w_mem_inst__abc_21203_new_n5816_; 
wire w_mem_inst__abc_21203_new_n5817_; 
wire w_mem_inst__abc_21203_new_n5818_; 
wire w_mem_inst__abc_21203_new_n5820_; 
wire w_mem_inst__abc_21203_new_n5821_; 
wire w_mem_inst__abc_21203_new_n5822_; 
wire w_mem_inst__abc_21203_new_n5823_; 
wire w_mem_inst__abc_21203_new_n5824_; 
wire w_mem_inst__abc_21203_new_n5826_; 
wire w_mem_inst__abc_21203_new_n5827_; 
wire w_mem_inst__abc_21203_new_n5828_; 
wire w_mem_inst__abc_21203_new_n5829_; 
wire w_mem_inst__abc_21203_new_n5830_; 
wire w_mem_inst__abc_21203_new_n5832_; 
wire w_mem_inst__abc_21203_new_n5833_; 
wire w_mem_inst__abc_21203_new_n5834_; 
wire w_mem_inst__abc_21203_new_n5835_; 
wire w_mem_inst__abc_21203_new_n5836_; 
wire w_mem_inst__abc_21203_new_n5838_; 
wire w_mem_inst__abc_21203_new_n5839_; 
wire w_mem_inst__abc_21203_new_n5840_; 
wire w_mem_inst__abc_21203_new_n5841_; 
wire w_mem_inst__abc_21203_new_n5842_; 
wire w_mem_inst__abc_21203_new_n5844_; 
wire w_mem_inst__abc_21203_new_n5845_; 
wire w_mem_inst__abc_21203_new_n5846_; 
wire w_mem_inst__abc_21203_new_n5847_; 
wire w_mem_inst__abc_21203_new_n5848_; 
wire w_mem_inst__abc_21203_new_n5850_; 
wire w_mem_inst__abc_21203_new_n5851_; 
wire w_mem_inst__abc_21203_new_n5852_; 
wire w_mem_inst__abc_21203_new_n5853_; 
wire w_mem_inst__abc_21203_new_n5854_; 
wire w_mem_inst__abc_21203_new_n5856_; 
wire w_mem_inst__abc_21203_new_n5857_; 
wire w_mem_inst__abc_21203_new_n5858_; 
wire w_mem_inst__abc_21203_new_n5859_; 
wire w_mem_inst__abc_21203_new_n5860_; 
wire w_mem_inst__abc_21203_new_n5862_; 
wire w_mem_inst__abc_21203_new_n5863_; 
wire w_mem_inst__abc_21203_new_n5864_; 
wire w_mem_inst__abc_21203_new_n5865_; 
wire w_mem_inst__abc_21203_new_n5866_; 
wire w_mem_inst__abc_21203_new_n5868_; 
wire w_mem_inst__abc_21203_new_n5869_; 
wire w_mem_inst__abc_21203_new_n5870_; 
wire w_mem_inst__abc_21203_new_n5871_; 
wire w_mem_inst__abc_21203_new_n5872_; 
wire w_mem_inst__abc_21203_new_n5874_; 
wire w_mem_inst__abc_21203_new_n5875_; 
wire w_mem_inst__abc_21203_new_n5876_; 
wire w_mem_inst__abc_21203_new_n5877_; 
wire w_mem_inst__abc_21203_new_n5878_; 
wire w_mem_inst__abc_21203_new_n5880_; 
wire w_mem_inst__abc_21203_new_n5881_; 
wire w_mem_inst__abc_21203_new_n5882_; 
wire w_mem_inst__abc_21203_new_n5883_; 
wire w_mem_inst__abc_21203_new_n5884_; 
wire w_mem_inst__abc_21203_new_n5886_; 
wire w_mem_inst__abc_21203_new_n5887_; 
wire w_mem_inst__abc_21203_new_n5888_; 
wire w_mem_inst__abc_21203_new_n5889_; 
wire w_mem_inst__abc_21203_new_n5890_; 
wire w_mem_inst__abc_21203_new_n5892_; 
wire w_mem_inst__abc_21203_new_n5893_; 
wire w_mem_inst__abc_21203_new_n5894_; 
wire w_mem_inst__abc_21203_new_n5895_; 
wire w_mem_inst__abc_21203_new_n5896_; 
wire w_mem_inst__abc_21203_new_n5898_; 
wire w_mem_inst__abc_21203_new_n5899_; 
wire w_mem_inst__abc_21203_new_n5900_; 
wire w_mem_inst__abc_21203_new_n5901_; 
wire w_mem_inst__abc_21203_new_n5902_; 
wire w_mem_inst__abc_21203_new_n5904_; 
wire w_mem_inst__abc_21203_new_n5905_; 
wire w_mem_inst__abc_21203_new_n5906_; 
wire w_mem_inst__abc_21203_new_n5907_; 
wire w_mem_inst__abc_21203_new_n5908_; 
wire w_mem_inst__abc_21203_new_n5910_; 
wire w_mem_inst__abc_21203_new_n5911_; 
wire w_mem_inst__abc_21203_new_n5912_; 
wire w_mem_inst__abc_21203_new_n5913_; 
wire w_mem_inst__abc_21203_new_n5914_; 
wire w_mem_inst__abc_21203_new_n5916_; 
wire w_mem_inst__abc_21203_new_n5917_; 
wire w_mem_inst__abc_21203_new_n5918_; 
wire w_mem_inst__abc_21203_new_n5919_; 
wire w_mem_inst__abc_21203_new_n5920_; 
wire w_mem_inst__abc_21203_new_n5922_; 
wire w_mem_inst__abc_21203_new_n5923_; 
wire w_mem_inst__abc_21203_new_n5924_; 
wire w_mem_inst__abc_21203_new_n5925_; 
wire w_mem_inst__abc_21203_new_n5926_; 
wire w_mem_inst__abc_21203_new_n5928_; 
wire w_mem_inst__abc_21203_new_n5929_; 
wire w_mem_inst__abc_21203_new_n5930_; 
wire w_mem_inst__abc_21203_new_n5931_; 
wire w_mem_inst__abc_21203_new_n5932_; 
wire w_mem_inst__abc_21203_new_n5934_; 
wire w_mem_inst__abc_21203_new_n5935_; 
wire w_mem_inst__abc_21203_new_n5936_; 
wire w_mem_inst__abc_21203_new_n5937_; 
wire w_mem_inst__abc_21203_new_n5938_; 
wire w_mem_inst__abc_21203_new_n5940_; 
wire w_mem_inst__abc_21203_new_n5941_; 
wire w_mem_inst__abc_21203_new_n5942_; 
wire w_mem_inst__abc_21203_new_n5943_; 
wire w_mem_inst__abc_21203_new_n5944_; 
wire w_mem_inst__abc_21203_new_n5946_; 
wire w_mem_inst__abc_21203_new_n5947_; 
wire w_mem_inst__abc_21203_new_n5948_; 
wire w_mem_inst__abc_21203_new_n5949_; 
wire w_mem_inst__abc_21203_new_n5950_; 
wire w_mem_inst__abc_21203_new_n5952_; 
wire w_mem_inst__abc_21203_new_n5953_; 
wire w_mem_inst__abc_21203_new_n5954_; 
wire w_mem_inst__abc_21203_new_n5955_; 
wire w_mem_inst__abc_21203_new_n5956_; 
wire w_mem_inst__abc_21203_new_n5958_; 
wire w_mem_inst__abc_21203_new_n5959_; 
wire w_mem_inst__abc_21203_new_n5960_; 
wire w_mem_inst__abc_21203_new_n5961_; 
wire w_mem_inst__abc_21203_new_n5962_; 
wire w_mem_inst__abc_21203_new_n5964_; 
wire w_mem_inst__abc_21203_new_n5965_; 
wire w_mem_inst__abc_21203_new_n5966_; 
wire w_mem_inst__abc_21203_new_n5967_; 
wire w_mem_inst__abc_21203_new_n5968_; 
wire w_mem_inst__abc_21203_new_n5970_; 
wire w_mem_inst__abc_21203_new_n5971_; 
wire w_mem_inst__abc_21203_new_n5972_; 
wire w_mem_inst__abc_21203_new_n5973_; 
wire w_mem_inst__abc_21203_new_n5974_; 
wire w_mem_inst__abc_21203_new_n5976_; 
wire w_mem_inst__abc_21203_new_n5977_; 
wire w_mem_inst__abc_21203_new_n5978_; 
wire w_mem_inst__abc_21203_new_n5979_; 
wire w_mem_inst__abc_21203_new_n5980_; 
wire w_mem_inst__abc_21203_new_n5982_; 
wire w_mem_inst__abc_21203_new_n5983_; 
wire w_mem_inst__abc_21203_new_n5984_; 
wire w_mem_inst__abc_21203_new_n5985_; 
wire w_mem_inst__abc_21203_new_n5986_; 
wire w_mem_inst__abc_21203_new_n5988_; 
wire w_mem_inst__abc_21203_new_n5989_; 
wire w_mem_inst__abc_21203_new_n5990_; 
wire w_mem_inst__abc_21203_new_n5991_; 
wire w_mem_inst__abc_21203_new_n5992_; 
wire w_mem_inst__abc_21203_new_n5994_; 
wire w_mem_inst__abc_21203_new_n5995_; 
wire w_mem_inst__abc_21203_new_n5996_; 
wire w_mem_inst__abc_21203_new_n5997_; 
wire w_mem_inst__abc_21203_new_n5998_; 
wire w_mem_inst__abc_21203_new_n6000_; 
wire w_mem_inst__abc_21203_new_n6001_; 
wire w_mem_inst__abc_21203_new_n6002_; 
wire w_mem_inst__abc_21203_new_n6003_; 
wire w_mem_inst__abc_21203_new_n6004_; 
wire w_mem_inst__abc_21203_new_n6006_; 
wire w_mem_inst__abc_21203_new_n6007_; 
wire w_mem_inst__abc_21203_new_n6008_; 
wire w_mem_inst__abc_21203_new_n6009_; 
wire w_mem_inst__abc_21203_new_n6010_; 
wire w_mem_inst__abc_21203_new_n6012_; 
wire w_mem_inst__abc_21203_new_n6013_; 
wire w_mem_inst__abc_21203_new_n6014_; 
wire w_mem_inst__abc_21203_new_n6015_; 
wire w_mem_inst__abc_21203_new_n6016_; 
wire w_mem_inst__abc_21203_new_n6018_; 
wire w_mem_inst__abc_21203_new_n6019_; 
wire w_mem_inst__abc_21203_new_n6020_; 
wire w_mem_inst__abc_21203_new_n6021_; 
wire w_mem_inst__abc_21203_new_n6022_; 
wire w_mem_inst__abc_21203_new_n6024_; 
wire w_mem_inst__abc_21203_new_n6025_; 
wire w_mem_inst__abc_21203_new_n6026_; 
wire w_mem_inst__abc_21203_new_n6027_; 
wire w_mem_inst__abc_21203_new_n6028_; 
wire w_mem_inst__abc_21203_new_n6030_; 
wire w_mem_inst__abc_21203_new_n6031_; 
wire w_mem_inst__abc_21203_new_n6032_; 
wire w_mem_inst__abc_21203_new_n6033_; 
wire w_mem_inst__abc_21203_new_n6034_; 
wire w_mem_inst__abc_21203_new_n6036_; 
wire w_mem_inst__abc_21203_new_n6037_; 
wire w_mem_inst__abc_21203_new_n6038_; 
wire w_mem_inst__abc_21203_new_n6039_; 
wire w_mem_inst__abc_21203_new_n6040_; 
wire w_mem_inst__abc_21203_new_n6042_; 
wire w_mem_inst__abc_21203_new_n6043_; 
wire w_mem_inst__abc_21203_new_n6044_; 
wire w_mem_inst__abc_21203_new_n6045_; 
wire w_mem_inst__abc_21203_new_n6046_; 
wire w_mem_inst__abc_21203_new_n6048_; 
wire w_mem_inst__abc_21203_new_n6049_; 
wire w_mem_inst__abc_21203_new_n6050_; 
wire w_mem_inst__abc_21203_new_n6051_; 
wire w_mem_inst__abc_21203_new_n6052_; 
wire w_mem_inst__abc_21203_new_n6054_; 
wire w_mem_inst__abc_21203_new_n6055_; 
wire w_mem_inst__abc_21203_new_n6056_; 
wire w_mem_inst__abc_21203_new_n6057_; 
wire w_mem_inst__abc_21203_new_n6058_; 
wire w_mem_inst__abc_21203_new_n6060_; 
wire w_mem_inst__abc_21203_new_n6061_; 
wire w_mem_inst__abc_21203_new_n6062_; 
wire w_mem_inst__abc_21203_new_n6063_; 
wire w_mem_inst__abc_21203_new_n6064_; 
wire w_mem_inst__abc_21203_new_n6066_; 
wire w_mem_inst__abc_21203_new_n6067_; 
wire w_mem_inst__abc_21203_new_n6068_; 
wire w_mem_inst__abc_21203_new_n6069_; 
wire w_mem_inst__abc_21203_new_n6070_; 
wire w_mem_inst__abc_21203_new_n6072_; 
wire w_mem_inst__abc_21203_new_n6073_; 
wire w_mem_inst__abc_21203_new_n6074_; 
wire w_mem_inst__abc_21203_new_n6075_; 
wire w_mem_inst__abc_21203_new_n6076_; 
wire w_mem_inst__abc_21203_new_n6078_; 
wire w_mem_inst__abc_21203_new_n6079_; 
wire w_mem_inst__abc_21203_new_n6080_; 
wire w_mem_inst__abc_21203_new_n6081_; 
wire w_mem_inst__abc_21203_new_n6082_; 
wire w_mem_inst__abc_21203_new_n6084_; 
wire w_mem_inst__abc_21203_new_n6085_; 
wire w_mem_inst__abc_21203_new_n6086_; 
wire w_mem_inst__abc_21203_new_n6087_; 
wire w_mem_inst__abc_21203_new_n6088_; 
wire w_mem_inst__abc_21203_new_n6090_; 
wire w_mem_inst__abc_21203_new_n6091_; 
wire w_mem_inst__abc_21203_new_n6092_; 
wire w_mem_inst__abc_21203_new_n6093_; 
wire w_mem_inst__abc_21203_new_n6094_; 
wire w_mem_inst__abc_21203_new_n6096_; 
wire w_mem_inst__abc_21203_new_n6097_; 
wire w_mem_inst__abc_21203_new_n6098_; 
wire w_mem_inst__abc_21203_new_n6099_; 
wire w_mem_inst__abc_21203_new_n6100_; 
wire w_mem_inst__abc_21203_new_n6102_; 
wire w_mem_inst__abc_21203_new_n6103_; 
wire w_mem_inst__abc_21203_new_n6104_; 
wire w_mem_inst__abc_21203_new_n6105_; 
wire w_mem_inst__abc_21203_new_n6106_; 
wire w_mem_inst__abc_21203_new_n6108_; 
wire w_mem_inst__abc_21203_new_n6109_; 
wire w_mem_inst__abc_21203_new_n6110_; 
wire w_mem_inst__abc_21203_new_n6111_; 
wire w_mem_inst__abc_21203_new_n6112_; 
wire w_mem_inst__abc_21203_new_n6114_; 
wire w_mem_inst__abc_21203_new_n6115_; 
wire w_mem_inst__abc_21203_new_n6116_; 
wire w_mem_inst__abc_21203_new_n6117_; 
wire w_mem_inst__abc_21203_new_n6118_; 
wire w_mem_inst__abc_21203_new_n6120_; 
wire w_mem_inst__abc_21203_new_n6121_; 
wire w_mem_inst__abc_21203_new_n6122_; 
wire w_mem_inst__abc_21203_new_n6123_; 
wire w_mem_inst__abc_21203_new_n6124_; 
wire w_mem_inst__abc_21203_new_n6126_; 
wire w_mem_inst__abc_21203_new_n6127_; 
wire w_mem_inst__abc_21203_new_n6128_; 
wire w_mem_inst__abc_21203_new_n6129_; 
wire w_mem_inst__abc_21203_new_n6130_; 
wire w_mem_inst__abc_21203_new_n6132_; 
wire w_mem_inst__abc_21203_new_n6133_; 
wire w_mem_inst__abc_21203_new_n6134_; 
wire w_mem_inst__abc_21203_new_n6135_; 
wire w_mem_inst__abc_21203_new_n6136_; 
wire w_mem_inst__abc_21203_new_n6138_; 
wire w_mem_inst__abc_21203_new_n6139_; 
wire w_mem_inst__abc_21203_new_n6140_; 
wire w_mem_inst__abc_21203_new_n6141_; 
wire w_mem_inst__abc_21203_new_n6142_; 
wire w_mem_inst__abc_21203_new_n6144_; 
wire w_mem_inst__abc_21203_new_n6145_; 
wire w_mem_inst__abc_21203_new_n6146_; 
wire w_mem_inst__abc_21203_new_n6147_; 
wire w_mem_inst__abc_21203_new_n6148_; 
wire w_mem_inst__abc_21203_new_n6150_; 
wire w_mem_inst__abc_21203_new_n6151_; 
wire w_mem_inst__abc_21203_new_n6152_; 
wire w_mem_inst__abc_21203_new_n6153_; 
wire w_mem_inst__abc_21203_new_n6154_; 
wire w_mem_inst__abc_21203_new_n6156_; 
wire w_mem_inst__abc_21203_new_n6157_; 
wire w_mem_inst__abc_21203_new_n6158_; 
wire w_mem_inst__abc_21203_new_n6159_; 
wire w_mem_inst__abc_21203_new_n6160_; 
wire w_mem_inst__abc_21203_new_n6162_; 
wire w_mem_inst__abc_21203_new_n6163_; 
wire w_mem_inst__abc_21203_new_n6164_; 
wire w_mem_inst__abc_21203_new_n6165_; 
wire w_mem_inst__abc_21203_new_n6166_; 
wire w_mem_inst__abc_21203_new_n6168_; 
wire w_mem_inst__abc_21203_new_n6169_; 
wire w_mem_inst__abc_21203_new_n6170_; 
wire w_mem_inst__abc_21203_new_n6171_; 
wire w_mem_inst__abc_21203_new_n6172_; 
wire w_mem_inst__abc_21203_new_n6174_; 
wire w_mem_inst__abc_21203_new_n6175_; 
wire w_mem_inst__abc_21203_new_n6176_; 
wire w_mem_inst__abc_21203_new_n6177_; 
wire w_mem_inst__abc_21203_new_n6178_; 
wire w_mem_inst__abc_21203_new_n6180_; 
wire w_mem_inst__abc_21203_new_n6181_; 
wire w_mem_inst__abc_21203_new_n6182_; 
wire w_mem_inst__abc_21203_new_n6183_; 
wire w_mem_inst__abc_21203_new_n6184_; 
wire w_mem_inst__abc_21203_new_n6186_; 
wire w_mem_inst__abc_21203_new_n6187_; 
wire w_mem_inst__abc_21203_new_n6188_; 
wire w_mem_inst__abc_21203_new_n6189_; 
wire w_mem_inst__abc_21203_new_n6190_; 
wire w_mem_inst__abc_21203_new_n6192_; 
wire w_mem_inst__abc_21203_new_n6193_; 
wire w_mem_inst__abc_21203_new_n6194_; 
wire w_mem_inst__abc_21203_new_n6195_; 
wire w_mem_inst__abc_21203_new_n6196_; 
wire w_mem_inst__abc_21203_new_n6198_; 
wire w_mem_inst__abc_21203_new_n6199_; 
wire w_mem_inst__abc_21203_new_n6200_; 
wire w_mem_inst__abc_21203_new_n6201_; 
wire w_mem_inst__abc_21203_new_n6202_; 
wire w_mem_inst__abc_21203_new_n6204_; 
wire w_mem_inst__abc_21203_new_n6205_; 
wire w_mem_inst__abc_21203_new_n6206_; 
wire w_mem_inst__abc_21203_new_n6207_; 
wire w_mem_inst__abc_21203_new_n6208_; 
wire w_mem_inst__abc_21203_new_n6210_; 
wire w_mem_inst__abc_21203_new_n6211_; 
wire w_mem_inst__abc_21203_new_n6212_; 
wire w_mem_inst__abc_21203_new_n6213_; 
wire w_mem_inst__abc_21203_new_n6214_; 
wire w_mem_inst__abc_21203_new_n6216_; 
wire w_mem_inst__abc_21203_new_n6217_; 
wire w_mem_inst__abc_21203_new_n6218_; 
wire w_mem_inst__abc_21203_new_n6219_; 
wire w_mem_inst__abc_21203_new_n6220_; 
wire w_mem_inst__abc_21203_new_n6222_; 
wire w_mem_inst__abc_21203_new_n6223_; 
wire w_mem_inst__abc_21203_new_n6224_; 
wire w_mem_inst__abc_21203_new_n6225_; 
wire w_mem_inst__abc_21203_new_n6226_; 
wire w_mem_inst__abc_21203_new_n6228_; 
wire w_mem_inst__abc_21203_new_n6229_; 
wire w_mem_inst__abc_21203_new_n6230_; 
wire w_mem_inst__abc_21203_new_n6231_; 
wire w_mem_inst__abc_21203_new_n6233_; 
wire w_mem_inst__abc_21203_new_n6234_; 
wire w_mem_inst__abc_21203_new_n6235_; 
wire w_mem_inst__abc_21203_new_n6237_; 
wire w_mem_inst__abc_21203_new_n6238_; 
wire w_mem_inst__abc_21203_new_n6239_; 
wire w_mem_inst__abc_21203_new_n6240_; 
wire w_mem_inst__abc_21203_new_n6241_; 
wire w_mem_inst__abc_21203_new_n6242_; 
wire w_mem_inst__abc_21203_new_n6243_; 
wire w_mem_inst__abc_21203_new_n6245_; 
wire w_mem_inst__abc_21203_new_n6246_; 
wire w_mem_inst__abc_21203_new_n6247_; 
wire w_mem_inst__abc_21203_new_n6248_; 
wire w_mem_inst__abc_21203_new_n6250_; 
wire w_mem_inst__abc_21203_new_n6251_; 
wire w_mem_inst__abc_21203_new_n6252_; 
wire w_mem_inst__abc_21203_new_n6253_; 
wire w_mem_inst__abc_21203_new_n6255_; 
wire w_mem_inst__abc_21203_new_n6256_; 
wire w_mem_inst__abc_21203_new_n6257_; 
wire w_mem_inst__abc_21203_new_n6258_; 
wire w_mem_inst__abc_21203_new_n6260_; 
wire w_mem_inst__abc_21203_new_n6261_; 
wire w_mem_inst__abc_21203_new_n6262_; 
wire w_mem_inst__abc_21203_new_n6263_; 
wire w_mem_inst_w_ctr_reg_0_; 
wire w_mem_inst_w_ctr_reg_1_; 
wire w_mem_inst_w_ctr_reg_2_; 
wire w_mem_inst_w_ctr_reg_3_; 
wire w_mem_inst_w_ctr_reg_4_; 
wire w_mem_inst_w_ctr_reg_5_; 
wire w_mem_inst_w_ctr_reg_6_; 
wire w_mem_inst_w_mem_0__0_; 
wire w_mem_inst_w_mem_0__10_; 
wire w_mem_inst_w_mem_0__11_; 
wire w_mem_inst_w_mem_0__12_; 
wire w_mem_inst_w_mem_0__13_; 
wire w_mem_inst_w_mem_0__14_; 
wire w_mem_inst_w_mem_0__15_; 
wire w_mem_inst_w_mem_0__16_; 
wire w_mem_inst_w_mem_0__17_; 
wire w_mem_inst_w_mem_0__18_; 
wire w_mem_inst_w_mem_0__19_; 
wire w_mem_inst_w_mem_0__1_; 
wire w_mem_inst_w_mem_0__20_; 
wire w_mem_inst_w_mem_0__21_; 
wire w_mem_inst_w_mem_0__22_; 
wire w_mem_inst_w_mem_0__23_; 
wire w_mem_inst_w_mem_0__24_; 
wire w_mem_inst_w_mem_0__25_; 
wire w_mem_inst_w_mem_0__26_; 
wire w_mem_inst_w_mem_0__27_; 
wire w_mem_inst_w_mem_0__28_; 
wire w_mem_inst_w_mem_0__29_; 
wire w_mem_inst_w_mem_0__2_; 
wire w_mem_inst_w_mem_0__30_; 
wire w_mem_inst_w_mem_0__31_; 
wire w_mem_inst_w_mem_0__3_; 
wire w_mem_inst_w_mem_0__4_; 
wire w_mem_inst_w_mem_0__5_; 
wire w_mem_inst_w_mem_0__6_; 
wire w_mem_inst_w_mem_0__7_; 
wire w_mem_inst_w_mem_0__8_; 
wire w_mem_inst_w_mem_0__9_; 
wire w_mem_inst_w_mem_10__0_; 
wire w_mem_inst_w_mem_10__10_; 
wire w_mem_inst_w_mem_10__11_; 
wire w_mem_inst_w_mem_10__12_; 
wire w_mem_inst_w_mem_10__13_; 
wire w_mem_inst_w_mem_10__14_; 
wire w_mem_inst_w_mem_10__15_; 
wire w_mem_inst_w_mem_10__16_; 
wire w_mem_inst_w_mem_10__17_; 
wire w_mem_inst_w_mem_10__18_; 
wire w_mem_inst_w_mem_10__19_; 
wire w_mem_inst_w_mem_10__1_; 
wire w_mem_inst_w_mem_10__20_; 
wire w_mem_inst_w_mem_10__21_; 
wire w_mem_inst_w_mem_10__22_; 
wire w_mem_inst_w_mem_10__23_; 
wire w_mem_inst_w_mem_10__24_; 
wire w_mem_inst_w_mem_10__25_; 
wire w_mem_inst_w_mem_10__26_; 
wire w_mem_inst_w_mem_10__27_; 
wire w_mem_inst_w_mem_10__28_; 
wire w_mem_inst_w_mem_10__29_; 
wire w_mem_inst_w_mem_10__2_; 
wire w_mem_inst_w_mem_10__30_; 
wire w_mem_inst_w_mem_10__31_; 
wire w_mem_inst_w_mem_10__3_; 
wire w_mem_inst_w_mem_10__4_; 
wire w_mem_inst_w_mem_10__5_; 
wire w_mem_inst_w_mem_10__6_; 
wire w_mem_inst_w_mem_10__7_; 
wire w_mem_inst_w_mem_10__8_; 
wire w_mem_inst_w_mem_10__9_; 
wire w_mem_inst_w_mem_11__0_; 
wire w_mem_inst_w_mem_11__10_; 
wire w_mem_inst_w_mem_11__11_; 
wire w_mem_inst_w_mem_11__12_; 
wire w_mem_inst_w_mem_11__13_; 
wire w_mem_inst_w_mem_11__14_; 
wire w_mem_inst_w_mem_11__15_; 
wire w_mem_inst_w_mem_11__16_; 
wire w_mem_inst_w_mem_11__17_; 
wire w_mem_inst_w_mem_11__18_; 
wire w_mem_inst_w_mem_11__19_; 
wire w_mem_inst_w_mem_11__1_; 
wire w_mem_inst_w_mem_11__20_; 
wire w_mem_inst_w_mem_11__21_; 
wire w_mem_inst_w_mem_11__22_; 
wire w_mem_inst_w_mem_11__23_; 
wire w_mem_inst_w_mem_11__24_; 
wire w_mem_inst_w_mem_11__25_; 
wire w_mem_inst_w_mem_11__26_; 
wire w_mem_inst_w_mem_11__27_; 
wire w_mem_inst_w_mem_11__28_; 
wire w_mem_inst_w_mem_11__29_; 
wire w_mem_inst_w_mem_11__2_; 
wire w_mem_inst_w_mem_11__30_; 
wire w_mem_inst_w_mem_11__31_; 
wire w_mem_inst_w_mem_11__3_; 
wire w_mem_inst_w_mem_11__4_; 
wire w_mem_inst_w_mem_11__5_; 
wire w_mem_inst_w_mem_11__6_; 
wire w_mem_inst_w_mem_11__7_; 
wire w_mem_inst_w_mem_11__8_; 
wire w_mem_inst_w_mem_11__9_; 
wire w_mem_inst_w_mem_12__0_; 
wire w_mem_inst_w_mem_12__10_; 
wire w_mem_inst_w_mem_12__11_; 
wire w_mem_inst_w_mem_12__12_; 
wire w_mem_inst_w_mem_12__13_; 
wire w_mem_inst_w_mem_12__14_; 
wire w_mem_inst_w_mem_12__15_; 
wire w_mem_inst_w_mem_12__16_; 
wire w_mem_inst_w_mem_12__17_; 
wire w_mem_inst_w_mem_12__18_; 
wire w_mem_inst_w_mem_12__19_; 
wire w_mem_inst_w_mem_12__1_; 
wire w_mem_inst_w_mem_12__20_; 
wire w_mem_inst_w_mem_12__21_; 
wire w_mem_inst_w_mem_12__22_; 
wire w_mem_inst_w_mem_12__23_; 
wire w_mem_inst_w_mem_12__24_; 
wire w_mem_inst_w_mem_12__25_; 
wire w_mem_inst_w_mem_12__26_; 
wire w_mem_inst_w_mem_12__27_; 
wire w_mem_inst_w_mem_12__28_; 
wire w_mem_inst_w_mem_12__29_; 
wire w_mem_inst_w_mem_12__2_; 
wire w_mem_inst_w_mem_12__30_; 
wire w_mem_inst_w_mem_12__31_; 
wire w_mem_inst_w_mem_12__3_; 
wire w_mem_inst_w_mem_12__4_; 
wire w_mem_inst_w_mem_12__5_; 
wire w_mem_inst_w_mem_12__6_; 
wire w_mem_inst_w_mem_12__7_; 
wire w_mem_inst_w_mem_12__8_; 
wire w_mem_inst_w_mem_12__9_; 
wire w_mem_inst_w_mem_13__0_; 
wire w_mem_inst_w_mem_13__10_; 
wire w_mem_inst_w_mem_13__11_; 
wire w_mem_inst_w_mem_13__12_; 
wire w_mem_inst_w_mem_13__13_; 
wire w_mem_inst_w_mem_13__14_; 
wire w_mem_inst_w_mem_13__15_; 
wire w_mem_inst_w_mem_13__16_; 
wire w_mem_inst_w_mem_13__17_; 
wire w_mem_inst_w_mem_13__18_; 
wire w_mem_inst_w_mem_13__19_; 
wire w_mem_inst_w_mem_13__1_; 
wire w_mem_inst_w_mem_13__20_; 
wire w_mem_inst_w_mem_13__21_; 
wire w_mem_inst_w_mem_13__22_; 
wire w_mem_inst_w_mem_13__23_; 
wire w_mem_inst_w_mem_13__24_; 
wire w_mem_inst_w_mem_13__25_; 
wire w_mem_inst_w_mem_13__26_; 
wire w_mem_inst_w_mem_13__27_; 
wire w_mem_inst_w_mem_13__28_; 
wire w_mem_inst_w_mem_13__29_; 
wire w_mem_inst_w_mem_13__2_; 
wire w_mem_inst_w_mem_13__30_; 
wire w_mem_inst_w_mem_13__31_; 
wire w_mem_inst_w_mem_13__3_; 
wire w_mem_inst_w_mem_13__4_; 
wire w_mem_inst_w_mem_13__5_; 
wire w_mem_inst_w_mem_13__6_; 
wire w_mem_inst_w_mem_13__7_; 
wire w_mem_inst_w_mem_13__8_; 
wire w_mem_inst_w_mem_13__9_; 
wire w_mem_inst_w_mem_14__0_; 
wire w_mem_inst_w_mem_14__10_; 
wire w_mem_inst_w_mem_14__11_; 
wire w_mem_inst_w_mem_14__12_; 
wire w_mem_inst_w_mem_14__13_; 
wire w_mem_inst_w_mem_14__14_; 
wire w_mem_inst_w_mem_14__15_; 
wire w_mem_inst_w_mem_14__16_; 
wire w_mem_inst_w_mem_14__17_; 
wire w_mem_inst_w_mem_14__18_; 
wire w_mem_inst_w_mem_14__19_; 
wire w_mem_inst_w_mem_14__1_; 
wire w_mem_inst_w_mem_14__20_; 
wire w_mem_inst_w_mem_14__21_; 
wire w_mem_inst_w_mem_14__22_; 
wire w_mem_inst_w_mem_14__23_; 
wire w_mem_inst_w_mem_14__24_; 
wire w_mem_inst_w_mem_14__25_; 
wire w_mem_inst_w_mem_14__26_; 
wire w_mem_inst_w_mem_14__27_; 
wire w_mem_inst_w_mem_14__28_; 
wire w_mem_inst_w_mem_14__29_; 
wire w_mem_inst_w_mem_14__2_; 
wire w_mem_inst_w_mem_14__30_; 
wire w_mem_inst_w_mem_14__31_; 
wire w_mem_inst_w_mem_14__3_; 
wire w_mem_inst_w_mem_14__4_; 
wire w_mem_inst_w_mem_14__5_; 
wire w_mem_inst_w_mem_14__6_; 
wire w_mem_inst_w_mem_14__7_; 
wire w_mem_inst_w_mem_14__8_; 
wire w_mem_inst_w_mem_14__9_; 
wire w_mem_inst_w_mem_15__0_; 
wire w_mem_inst_w_mem_15__10_; 
wire w_mem_inst_w_mem_15__11_; 
wire w_mem_inst_w_mem_15__12_; 
wire w_mem_inst_w_mem_15__13_; 
wire w_mem_inst_w_mem_15__14_; 
wire w_mem_inst_w_mem_15__15_; 
wire w_mem_inst_w_mem_15__16_; 
wire w_mem_inst_w_mem_15__17_; 
wire w_mem_inst_w_mem_15__18_; 
wire w_mem_inst_w_mem_15__19_; 
wire w_mem_inst_w_mem_15__1_; 
wire w_mem_inst_w_mem_15__20_; 
wire w_mem_inst_w_mem_15__21_; 
wire w_mem_inst_w_mem_15__22_; 
wire w_mem_inst_w_mem_15__23_; 
wire w_mem_inst_w_mem_15__24_; 
wire w_mem_inst_w_mem_15__25_; 
wire w_mem_inst_w_mem_15__26_; 
wire w_mem_inst_w_mem_15__27_; 
wire w_mem_inst_w_mem_15__28_; 
wire w_mem_inst_w_mem_15__29_; 
wire w_mem_inst_w_mem_15__2_; 
wire w_mem_inst_w_mem_15__30_; 
wire w_mem_inst_w_mem_15__31_; 
wire w_mem_inst_w_mem_15__3_; 
wire w_mem_inst_w_mem_15__4_; 
wire w_mem_inst_w_mem_15__5_; 
wire w_mem_inst_w_mem_15__6_; 
wire w_mem_inst_w_mem_15__7_; 
wire w_mem_inst_w_mem_15__8_; 
wire w_mem_inst_w_mem_15__9_; 
wire w_mem_inst_w_mem_1__0_; 
wire w_mem_inst_w_mem_1__10_; 
wire w_mem_inst_w_mem_1__11_; 
wire w_mem_inst_w_mem_1__12_; 
wire w_mem_inst_w_mem_1__13_; 
wire w_mem_inst_w_mem_1__14_; 
wire w_mem_inst_w_mem_1__15_; 
wire w_mem_inst_w_mem_1__16_; 
wire w_mem_inst_w_mem_1__17_; 
wire w_mem_inst_w_mem_1__18_; 
wire w_mem_inst_w_mem_1__19_; 
wire w_mem_inst_w_mem_1__1_; 
wire w_mem_inst_w_mem_1__20_; 
wire w_mem_inst_w_mem_1__21_; 
wire w_mem_inst_w_mem_1__22_; 
wire w_mem_inst_w_mem_1__23_; 
wire w_mem_inst_w_mem_1__24_; 
wire w_mem_inst_w_mem_1__25_; 
wire w_mem_inst_w_mem_1__26_; 
wire w_mem_inst_w_mem_1__27_; 
wire w_mem_inst_w_mem_1__28_; 
wire w_mem_inst_w_mem_1__29_; 
wire w_mem_inst_w_mem_1__2_; 
wire w_mem_inst_w_mem_1__30_; 
wire w_mem_inst_w_mem_1__31_; 
wire w_mem_inst_w_mem_1__3_; 
wire w_mem_inst_w_mem_1__4_; 
wire w_mem_inst_w_mem_1__5_; 
wire w_mem_inst_w_mem_1__6_; 
wire w_mem_inst_w_mem_1__7_; 
wire w_mem_inst_w_mem_1__8_; 
wire w_mem_inst_w_mem_1__9_; 
wire w_mem_inst_w_mem_2__0_; 
wire w_mem_inst_w_mem_2__10_; 
wire w_mem_inst_w_mem_2__11_; 
wire w_mem_inst_w_mem_2__12_; 
wire w_mem_inst_w_mem_2__13_; 
wire w_mem_inst_w_mem_2__14_; 
wire w_mem_inst_w_mem_2__15_; 
wire w_mem_inst_w_mem_2__16_; 
wire w_mem_inst_w_mem_2__17_; 
wire w_mem_inst_w_mem_2__18_; 
wire w_mem_inst_w_mem_2__19_; 
wire w_mem_inst_w_mem_2__1_; 
wire w_mem_inst_w_mem_2__20_; 
wire w_mem_inst_w_mem_2__21_; 
wire w_mem_inst_w_mem_2__22_; 
wire w_mem_inst_w_mem_2__23_; 
wire w_mem_inst_w_mem_2__24_; 
wire w_mem_inst_w_mem_2__25_; 
wire w_mem_inst_w_mem_2__26_; 
wire w_mem_inst_w_mem_2__27_; 
wire w_mem_inst_w_mem_2__28_; 
wire w_mem_inst_w_mem_2__29_; 
wire w_mem_inst_w_mem_2__2_; 
wire w_mem_inst_w_mem_2__30_; 
wire w_mem_inst_w_mem_2__31_; 
wire w_mem_inst_w_mem_2__3_; 
wire w_mem_inst_w_mem_2__4_; 
wire w_mem_inst_w_mem_2__5_; 
wire w_mem_inst_w_mem_2__6_; 
wire w_mem_inst_w_mem_2__7_; 
wire w_mem_inst_w_mem_2__8_; 
wire w_mem_inst_w_mem_2__9_; 
wire w_mem_inst_w_mem_3__0_; 
wire w_mem_inst_w_mem_3__10_; 
wire w_mem_inst_w_mem_3__11_; 
wire w_mem_inst_w_mem_3__12_; 
wire w_mem_inst_w_mem_3__13_; 
wire w_mem_inst_w_mem_3__14_; 
wire w_mem_inst_w_mem_3__15_; 
wire w_mem_inst_w_mem_3__16_; 
wire w_mem_inst_w_mem_3__17_; 
wire w_mem_inst_w_mem_3__18_; 
wire w_mem_inst_w_mem_3__19_; 
wire w_mem_inst_w_mem_3__1_; 
wire w_mem_inst_w_mem_3__20_; 
wire w_mem_inst_w_mem_3__21_; 
wire w_mem_inst_w_mem_3__22_; 
wire w_mem_inst_w_mem_3__23_; 
wire w_mem_inst_w_mem_3__24_; 
wire w_mem_inst_w_mem_3__25_; 
wire w_mem_inst_w_mem_3__26_; 
wire w_mem_inst_w_mem_3__27_; 
wire w_mem_inst_w_mem_3__28_; 
wire w_mem_inst_w_mem_3__29_; 
wire w_mem_inst_w_mem_3__2_; 
wire w_mem_inst_w_mem_3__30_; 
wire w_mem_inst_w_mem_3__31_; 
wire w_mem_inst_w_mem_3__3_; 
wire w_mem_inst_w_mem_3__4_; 
wire w_mem_inst_w_mem_3__5_; 
wire w_mem_inst_w_mem_3__6_; 
wire w_mem_inst_w_mem_3__7_; 
wire w_mem_inst_w_mem_3__8_; 
wire w_mem_inst_w_mem_3__9_; 
wire w_mem_inst_w_mem_4__0_; 
wire w_mem_inst_w_mem_4__10_; 
wire w_mem_inst_w_mem_4__11_; 
wire w_mem_inst_w_mem_4__12_; 
wire w_mem_inst_w_mem_4__13_; 
wire w_mem_inst_w_mem_4__14_; 
wire w_mem_inst_w_mem_4__15_; 
wire w_mem_inst_w_mem_4__16_; 
wire w_mem_inst_w_mem_4__17_; 
wire w_mem_inst_w_mem_4__18_; 
wire w_mem_inst_w_mem_4__19_; 
wire w_mem_inst_w_mem_4__1_; 
wire w_mem_inst_w_mem_4__20_; 
wire w_mem_inst_w_mem_4__21_; 
wire w_mem_inst_w_mem_4__22_; 
wire w_mem_inst_w_mem_4__23_; 
wire w_mem_inst_w_mem_4__24_; 
wire w_mem_inst_w_mem_4__25_; 
wire w_mem_inst_w_mem_4__26_; 
wire w_mem_inst_w_mem_4__27_; 
wire w_mem_inst_w_mem_4__28_; 
wire w_mem_inst_w_mem_4__29_; 
wire w_mem_inst_w_mem_4__2_; 
wire w_mem_inst_w_mem_4__30_; 
wire w_mem_inst_w_mem_4__31_; 
wire w_mem_inst_w_mem_4__3_; 
wire w_mem_inst_w_mem_4__4_; 
wire w_mem_inst_w_mem_4__5_; 
wire w_mem_inst_w_mem_4__6_; 
wire w_mem_inst_w_mem_4__7_; 
wire w_mem_inst_w_mem_4__8_; 
wire w_mem_inst_w_mem_4__9_; 
wire w_mem_inst_w_mem_5__0_; 
wire w_mem_inst_w_mem_5__10_; 
wire w_mem_inst_w_mem_5__11_; 
wire w_mem_inst_w_mem_5__12_; 
wire w_mem_inst_w_mem_5__13_; 
wire w_mem_inst_w_mem_5__14_; 
wire w_mem_inst_w_mem_5__15_; 
wire w_mem_inst_w_mem_5__16_; 
wire w_mem_inst_w_mem_5__17_; 
wire w_mem_inst_w_mem_5__18_; 
wire w_mem_inst_w_mem_5__19_; 
wire w_mem_inst_w_mem_5__1_; 
wire w_mem_inst_w_mem_5__20_; 
wire w_mem_inst_w_mem_5__21_; 
wire w_mem_inst_w_mem_5__22_; 
wire w_mem_inst_w_mem_5__23_; 
wire w_mem_inst_w_mem_5__24_; 
wire w_mem_inst_w_mem_5__25_; 
wire w_mem_inst_w_mem_5__26_; 
wire w_mem_inst_w_mem_5__27_; 
wire w_mem_inst_w_mem_5__28_; 
wire w_mem_inst_w_mem_5__29_; 
wire w_mem_inst_w_mem_5__2_; 
wire w_mem_inst_w_mem_5__30_; 
wire w_mem_inst_w_mem_5__31_; 
wire w_mem_inst_w_mem_5__3_; 
wire w_mem_inst_w_mem_5__4_; 
wire w_mem_inst_w_mem_5__5_; 
wire w_mem_inst_w_mem_5__6_; 
wire w_mem_inst_w_mem_5__7_; 
wire w_mem_inst_w_mem_5__8_; 
wire w_mem_inst_w_mem_5__9_; 
wire w_mem_inst_w_mem_6__0_; 
wire w_mem_inst_w_mem_6__10_; 
wire w_mem_inst_w_mem_6__11_; 
wire w_mem_inst_w_mem_6__12_; 
wire w_mem_inst_w_mem_6__13_; 
wire w_mem_inst_w_mem_6__14_; 
wire w_mem_inst_w_mem_6__15_; 
wire w_mem_inst_w_mem_6__16_; 
wire w_mem_inst_w_mem_6__17_; 
wire w_mem_inst_w_mem_6__18_; 
wire w_mem_inst_w_mem_6__19_; 
wire w_mem_inst_w_mem_6__1_; 
wire w_mem_inst_w_mem_6__20_; 
wire w_mem_inst_w_mem_6__21_; 
wire w_mem_inst_w_mem_6__22_; 
wire w_mem_inst_w_mem_6__23_; 
wire w_mem_inst_w_mem_6__24_; 
wire w_mem_inst_w_mem_6__25_; 
wire w_mem_inst_w_mem_6__26_; 
wire w_mem_inst_w_mem_6__27_; 
wire w_mem_inst_w_mem_6__28_; 
wire w_mem_inst_w_mem_6__29_; 
wire w_mem_inst_w_mem_6__2_; 
wire w_mem_inst_w_mem_6__30_; 
wire w_mem_inst_w_mem_6__31_; 
wire w_mem_inst_w_mem_6__3_; 
wire w_mem_inst_w_mem_6__4_; 
wire w_mem_inst_w_mem_6__5_; 
wire w_mem_inst_w_mem_6__6_; 
wire w_mem_inst_w_mem_6__7_; 
wire w_mem_inst_w_mem_6__8_; 
wire w_mem_inst_w_mem_6__9_; 
wire w_mem_inst_w_mem_7__0_; 
wire w_mem_inst_w_mem_7__10_; 
wire w_mem_inst_w_mem_7__11_; 
wire w_mem_inst_w_mem_7__12_; 
wire w_mem_inst_w_mem_7__13_; 
wire w_mem_inst_w_mem_7__14_; 
wire w_mem_inst_w_mem_7__15_; 
wire w_mem_inst_w_mem_7__16_; 
wire w_mem_inst_w_mem_7__17_; 
wire w_mem_inst_w_mem_7__18_; 
wire w_mem_inst_w_mem_7__19_; 
wire w_mem_inst_w_mem_7__1_; 
wire w_mem_inst_w_mem_7__20_; 
wire w_mem_inst_w_mem_7__21_; 
wire w_mem_inst_w_mem_7__22_; 
wire w_mem_inst_w_mem_7__23_; 
wire w_mem_inst_w_mem_7__24_; 
wire w_mem_inst_w_mem_7__25_; 
wire w_mem_inst_w_mem_7__26_; 
wire w_mem_inst_w_mem_7__27_; 
wire w_mem_inst_w_mem_7__28_; 
wire w_mem_inst_w_mem_7__29_; 
wire w_mem_inst_w_mem_7__2_; 
wire w_mem_inst_w_mem_7__30_; 
wire w_mem_inst_w_mem_7__31_; 
wire w_mem_inst_w_mem_7__3_; 
wire w_mem_inst_w_mem_7__4_; 
wire w_mem_inst_w_mem_7__5_; 
wire w_mem_inst_w_mem_7__6_; 
wire w_mem_inst_w_mem_7__7_; 
wire w_mem_inst_w_mem_7__8_; 
wire w_mem_inst_w_mem_7__9_; 
wire w_mem_inst_w_mem_8__0_; 
wire w_mem_inst_w_mem_8__10_; 
wire w_mem_inst_w_mem_8__11_; 
wire w_mem_inst_w_mem_8__12_; 
wire w_mem_inst_w_mem_8__13_; 
wire w_mem_inst_w_mem_8__14_; 
wire w_mem_inst_w_mem_8__15_; 
wire w_mem_inst_w_mem_8__16_; 
wire w_mem_inst_w_mem_8__17_; 
wire w_mem_inst_w_mem_8__18_; 
wire w_mem_inst_w_mem_8__19_; 
wire w_mem_inst_w_mem_8__1_; 
wire w_mem_inst_w_mem_8__20_; 
wire w_mem_inst_w_mem_8__21_; 
wire w_mem_inst_w_mem_8__22_; 
wire w_mem_inst_w_mem_8__23_; 
wire w_mem_inst_w_mem_8__24_; 
wire w_mem_inst_w_mem_8__25_; 
wire w_mem_inst_w_mem_8__26_; 
wire w_mem_inst_w_mem_8__27_; 
wire w_mem_inst_w_mem_8__28_; 
wire w_mem_inst_w_mem_8__29_; 
wire w_mem_inst_w_mem_8__2_; 
wire w_mem_inst_w_mem_8__30_; 
wire w_mem_inst_w_mem_8__31_; 
wire w_mem_inst_w_mem_8__3_; 
wire w_mem_inst_w_mem_8__4_; 
wire w_mem_inst_w_mem_8__5_; 
wire w_mem_inst_w_mem_8__6_; 
wire w_mem_inst_w_mem_8__7_; 
wire w_mem_inst_w_mem_8__8_; 
wire w_mem_inst_w_mem_8__9_; 
wire w_mem_inst_w_mem_9__0_; 
wire w_mem_inst_w_mem_9__10_; 
wire w_mem_inst_w_mem_9__11_; 
wire w_mem_inst_w_mem_9__12_; 
wire w_mem_inst_w_mem_9__13_; 
wire w_mem_inst_w_mem_9__14_; 
wire w_mem_inst_w_mem_9__15_; 
wire w_mem_inst_w_mem_9__16_; 
wire w_mem_inst_w_mem_9__17_; 
wire w_mem_inst_w_mem_9__18_; 
wire w_mem_inst_w_mem_9__19_; 
wire w_mem_inst_w_mem_9__1_; 
wire w_mem_inst_w_mem_9__20_; 
wire w_mem_inst_w_mem_9__21_; 
wire w_mem_inst_w_mem_9__22_; 
wire w_mem_inst_w_mem_9__23_; 
wire w_mem_inst_w_mem_9__24_; 
wire w_mem_inst_w_mem_9__25_; 
wire w_mem_inst_w_mem_9__26_; 
wire w_mem_inst_w_mem_9__27_; 
wire w_mem_inst_w_mem_9__28_; 
wire w_mem_inst_w_mem_9__29_; 
wire w_mem_inst_w_mem_9__2_; 
wire w_mem_inst_w_mem_9__30_; 
wire w_mem_inst_w_mem_9__31_; 
wire w_mem_inst_w_mem_9__3_; 
wire w_mem_inst_w_mem_9__4_; 
wire w_mem_inst_w_mem_9__5_; 
wire w_mem_inst_w_mem_9__6_; 
wire w_mem_inst_w_mem_9__7_; 
wire w_mem_inst_w_mem_9__8_; 
wire w_mem_inst_w_mem_9__9_; 
AND2X2 AND2X2_1 ( .A(ready), .B(init), .Y(_abc_15497_new_n699_));
AND2X2 AND2X2_10 ( .A(c_reg_20_), .B(\digest[84] ), .Y(_abc_15497_new_n715_));
AND2X2 AND2X2_100 ( .A(_abc_15497_new_n887_), .B(_abc_15497_new_n885_), .Y(_abc_15497_new_n888_));
AND2X2 AND2X2_1000 ( .A(\digest[129] ), .B(a_reg_1_), .Y(_abc_15497_new_n2719_));
AND2X2 AND2X2_1001 ( .A(_abc_15497_new_n2720_), .B(_abc_15497_new_n2718_), .Y(_abc_15497_new_n2721_));
AND2X2 AND2X2_1002 ( .A(_abc_15497_new_n2721_), .B(_abc_15497_new_n2711_), .Y(_abc_15497_new_n2722_));
AND2X2 AND2X2_1003 ( .A(_abc_15497_new_n2724_), .B(digest_update), .Y(_abc_15497_new_n2725_));
AND2X2 AND2X2_1004 ( .A(_abc_15497_new_n2725_), .B(_abc_15497_new_n2723_), .Y(_abc_15497_new_n2726_));
AND2X2 AND2X2_1005 ( .A(_abc_15497_new_n701_), .B(\digest[129] ), .Y(_abc_15497_new_n2727_));
AND2X2 AND2X2_1006 ( .A(_abc_15497_new_n2723_), .B(_abc_15497_new_n2720_), .Y(_abc_15497_new_n2729_));
AND2X2 AND2X2_1007 ( .A(\digest[130] ), .B(a_reg_2_), .Y(_abc_15497_new_n2732_));
AND2X2 AND2X2_1008 ( .A(_abc_15497_new_n2733_), .B(_abc_15497_new_n2731_), .Y(_abc_15497_new_n2734_));
AND2X2 AND2X2_1009 ( .A(_abc_15497_new_n2737_), .B(digest_update), .Y(_abc_15497_new_n2738_));
AND2X2 AND2X2_101 ( .A(_abc_15497_new_n889_), .B(_abc_15497_new_n891_), .Y(_abc_15497_new_n892_));
AND2X2 AND2X2_1010 ( .A(_abc_15497_new_n2738_), .B(_abc_15497_new_n2735_), .Y(_abc_15497_new_n2739_));
AND2X2 AND2X2_1011 ( .A(_abc_15497_new_n701_), .B(\digest[130] ), .Y(_abc_15497_new_n2740_));
AND2X2 AND2X2_1012 ( .A(_abc_15497_new_n701_), .B(\digest[131] ), .Y(_abc_15497_new_n2742_));
AND2X2 AND2X2_1013 ( .A(_abc_15497_new_n2737_), .B(_abc_15497_new_n2733_), .Y(_abc_15497_new_n2743_));
AND2X2 AND2X2_1014 ( .A(\digest[131] ), .B(a_reg_3_), .Y(_abc_15497_new_n2746_));
AND2X2 AND2X2_1015 ( .A(_abc_15497_new_n2747_), .B(_abc_15497_new_n2745_), .Y(_abc_15497_new_n2748_));
AND2X2 AND2X2_1016 ( .A(_abc_15497_new_n2751_), .B(digest_update), .Y(_abc_15497_new_n2752_));
AND2X2 AND2X2_1017 ( .A(_abc_15497_new_n2752_), .B(_abc_15497_new_n2749_), .Y(_abc_15497_new_n2753_));
AND2X2 AND2X2_1018 ( .A(\digest[132] ), .B(a_reg_4_), .Y(_abc_15497_new_n2756_));
AND2X2 AND2X2_1019 ( .A(_abc_15497_new_n2757_), .B(_abc_15497_new_n2755_), .Y(_abc_15497_new_n2758_));
AND2X2 AND2X2_102 ( .A(_abc_15497_new_n892_), .B(digest_update), .Y(_abc_15497_new_n893_));
AND2X2 AND2X2_1020 ( .A(_abc_15497_new_n2760_), .B(_abc_15497_new_n2747_), .Y(_abc_15497_new_n2761_));
AND2X2 AND2X2_1021 ( .A(_abc_15497_new_n2765_), .B(digest_update), .Y(_abc_15497_new_n2766_));
AND2X2 AND2X2_1022 ( .A(_abc_15497_new_n2766_), .B(_abc_15497_new_n2763_), .Y(_abc_15497_new_n2767_));
AND2X2 AND2X2_1023 ( .A(_abc_15497_new_n701_), .B(\digest[132] ), .Y(_abc_15497_new_n2768_));
AND2X2 AND2X2_1024 ( .A(_abc_15497_new_n701_), .B(\digest[133] ), .Y(_abc_15497_new_n2770_));
AND2X2 AND2X2_1025 ( .A(_abc_15497_new_n2765_), .B(_abc_15497_new_n2757_), .Y(_abc_15497_new_n2771_));
AND2X2 AND2X2_1026 ( .A(\digest[133] ), .B(a_reg_5_), .Y(_abc_15497_new_n2774_));
AND2X2 AND2X2_1027 ( .A(_abc_15497_new_n2775_), .B(_abc_15497_new_n2773_), .Y(_abc_15497_new_n2776_));
AND2X2 AND2X2_1028 ( .A(_abc_15497_new_n2779_), .B(digest_update), .Y(_abc_15497_new_n2780_));
AND2X2 AND2X2_1029 ( .A(_abc_15497_new_n2780_), .B(_abc_15497_new_n2777_), .Y(_abc_15497_new_n2781_));
AND2X2 AND2X2_103 ( .A(_abc_15497_new_n894_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n895_));
AND2X2 AND2X2_1030 ( .A(_abc_15497_new_n701_), .B(\digest[134] ), .Y(_abc_15497_new_n2783_));
AND2X2 AND2X2_1031 ( .A(_abc_15497_new_n2779_), .B(_abc_15497_new_n2775_), .Y(_abc_15497_new_n2784_));
AND2X2 AND2X2_1032 ( .A(\digest[134] ), .B(a_reg_6_), .Y(_abc_15497_new_n2787_));
AND2X2 AND2X2_1033 ( .A(_abc_15497_new_n2788_), .B(_abc_15497_new_n2786_), .Y(_abc_15497_new_n2789_));
AND2X2 AND2X2_1034 ( .A(_abc_15497_new_n2792_), .B(digest_update), .Y(_abc_15497_new_n2793_));
AND2X2 AND2X2_1035 ( .A(_abc_15497_new_n2793_), .B(_abc_15497_new_n2790_), .Y(_abc_15497_new_n2794_));
AND2X2 AND2X2_1036 ( .A(_abc_15497_new_n701_), .B(\digest[135] ), .Y(_abc_15497_new_n2796_));
AND2X2 AND2X2_1037 ( .A(\digest[135] ), .B(a_reg_7_), .Y(_abc_15497_new_n2799_));
AND2X2 AND2X2_1038 ( .A(_abc_15497_new_n2800_), .B(_abc_15497_new_n2798_), .Y(_abc_15497_new_n2801_));
AND2X2 AND2X2_1039 ( .A(_abc_15497_new_n2801_), .B(_abc_15497_new_n2787_), .Y(_abc_15497_new_n2806_));
AND2X2 AND2X2_104 ( .A(_abc_15497_new_n885_), .B(_abc_15497_new_n874_), .Y(_abc_15497_new_n897_));
AND2X2 AND2X2_1040 ( .A(_abc_15497_new_n2805_), .B(_abc_15497_new_n2807_), .Y(_abc_15497_new_n2808_));
AND2X2 AND2X2_1041 ( .A(_abc_15497_new_n2808_), .B(_abc_15497_new_n2803_), .Y(_abc_15497_new_n2809_));
AND2X2 AND2X2_1042 ( .A(_abc_15497_new_n2809_), .B(digest_update), .Y(_abc_15497_new_n2810_));
AND2X2 AND2X2_1043 ( .A(\digest[136] ), .B(a_reg_8_), .Y(_abc_15497_new_n2816_));
AND2X2 AND2X2_1044 ( .A(_abc_15497_new_n2817_), .B(_abc_15497_new_n2815_), .Y(_abc_15497_new_n2818_));
AND2X2 AND2X2_1045 ( .A(_abc_15497_new_n2814_), .B(_abc_15497_new_n2818_), .Y(_abc_15497_new_n2820_));
AND2X2 AND2X2_1046 ( .A(_abc_15497_new_n2821_), .B(_abc_15497_new_n2819_), .Y(_abc_15497_new_n2822_));
AND2X2 AND2X2_1047 ( .A(_abc_15497_new_n2822_), .B(digest_update), .Y(_abc_15497_new_n2823_));
AND2X2 AND2X2_1048 ( .A(_abc_15497_new_n2824_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n2825_));
AND2X2 AND2X2_1049 ( .A(_abc_15497_new_n2821_), .B(_abc_15497_new_n2817_), .Y(_abc_15497_new_n2827_));
AND2X2 AND2X2_105 ( .A(_abc_15497_new_n876_), .B(_abc_15497_new_n888_), .Y(_abc_15497_new_n899_));
AND2X2 AND2X2_1050 ( .A(\digest[137] ), .B(a_reg_9_), .Y(_abc_15497_new_n2830_));
AND2X2 AND2X2_1051 ( .A(_abc_15497_new_n2831_), .B(_abc_15497_new_n2829_), .Y(_abc_15497_new_n2832_));
AND2X2 AND2X2_1052 ( .A(_abc_15497_new_n2833_), .B(_abc_15497_new_n2835_), .Y(_abc_15497_new_n2836_));
AND2X2 AND2X2_1053 ( .A(_abc_15497_new_n2836_), .B(digest_update), .Y(_abc_15497_new_n2837_));
AND2X2 AND2X2_1054 ( .A(_abc_15497_new_n2838_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n2839_));
AND2X2 AND2X2_1055 ( .A(_abc_15497_new_n701_), .B(\digest[138] ), .Y(_abc_15497_new_n2841_));
AND2X2 AND2X2_1056 ( .A(\digest[138] ), .B(a_reg_10_), .Y(_abc_15497_new_n2843_));
AND2X2 AND2X2_1057 ( .A(_abc_15497_new_n2844_), .B(_abc_15497_new_n2842_), .Y(_abc_15497_new_n2845_));
AND2X2 AND2X2_1058 ( .A(_abc_15497_new_n2846_), .B(_abc_15497_new_n2831_), .Y(_abc_15497_new_n2847_));
AND2X2 AND2X2_1059 ( .A(_abc_15497_new_n2818_), .B(_abc_15497_new_n2832_), .Y(_abc_15497_new_n2849_));
AND2X2 AND2X2_106 ( .A(_abc_15497_new_n872_), .B(_abc_15497_new_n899_), .Y(_abc_15497_new_n900_));
AND2X2 AND2X2_1060 ( .A(_abc_15497_new_n2814_), .B(_abc_15497_new_n2849_), .Y(_abc_15497_new_n2850_));
AND2X2 AND2X2_1061 ( .A(_abc_15497_new_n2851_), .B(_abc_15497_new_n2845_), .Y(_abc_15497_new_n2853_));
AND2X2 AND2X2_1062 ( .A(_abc_15497_new_n2854_), .B(_abc_15497_new_n2852_), .Y(_abc_15497_new_n2855_));
AND2X2 AND2X2_1063 ( .A(_abc_15497_new_n2855_), .B(digest_update), .Y(_abc_15497_new_n2856_));
AND2X2 AND2X2_1064 ( .A(_abc_15497_new_n701_), .B(\digest[139] ), .Y(_abc_15497_new_n2858_));
AND2X2 AND2X2_1065 ( .A(_abc_15497_new_n2854_), .B(_abc_15497_new_n2844_), .Y(_abc_15497_new_n2859_));
AND2X2 AND2X2_1066 ( .A(\digest[139] ), .B(a_reg_11_), .Y(_abc_15497_new_n2862_));
AND2X2 AND2X2_1067 ( .A(_abc_15497_new_n2863_), .B(_abc_15497_new_n2861_), .Y(_abc_15497_new_n2864_));
AND2X2 AND2X2_1068 ( .A(_abc_15497_new_n2867_), .B(digest_update), .Y(_abc_15497_new_n2868_));
AND2X2 AND2X2_1069 ( .A(_abc_15497_new_n2868_), .B(_abc_15497_new_n2865_), .Y(_abc_15497_new_n2869_));
AND2X2 AND2X2_107 ( .A(\digest[92] ), .B(c_reg_28_), .Y(_abc_15497_new_n903_));
AND2X2 AND2X2_1070 ( .A(_abc_15497_new_n701_), .B(\digest[140] ), .Y(_abc_15497_new_n2871_));
AND2X2 AND2X2_1071 ( .A(_abc_15497_new_n2845_), .B(_abc_15497_new_n2864_), .Y(_abc_15497_new_n2872_));
AND2X2 AND2X2_1072 ( .A(_abc_15497_new_n2849_), .B(_abc_15497_new_n2872_), .Y(_abc_15497_new_n2873_));
AND2X2 AND2X2_1073 ( .A(_abc_15497_new_n2814_), .B(_abc_15497_new_n2873_), .Y(_abc_15497_new_n2874_));
AND2X2 AND2X2_1074 ( .A(_abc_15497_new_n2848_), .B(_abc_15497_new_n2872_), .Y(_abc_15497_new_n2875_));
AND2X2 AND2X2_1075 ( .A(_abc_15497_new_n2877_), .B(_abc_15497_new_n2863_), .Y(_abc_15497_new_n2878_));
AND2X2 AND2X2_1076 ( .A(_abc_15497_new_n2876_), .B(_abc_15497_new_n2878_), .Y(_abc_15497_new_n2879_));
AND2X2 AND2X2_1077 ( .A(\digest[140] ), .B(a_reg_12_), .Y(_abc_15497_new_n2883_));
AND2X2 AND2X2_1078 ( .A(_abc_15497_new_n2884_), .B(_abc_15497_new_n2882_), .Y(_abc_15497_new_n2885_));
AND2X2 AND2X2_1079 ( .A(_abc_15497_new_n2881_), .B(_abc_15497_new_n2885_), .Y(_abc_15497_new_n2887_));
AND2X2 AND2X2_108 ( .A(_abc_15497_new_n904_), .B(_abc_15497_new_n902_), .Y(_abc_15497_new_n905_));
AND2X2 AND2X2_1080 ( .A(_abc_15497_new_n2888_), .B(_abc_15497_new_n2886_), .Y(_abc_15497_new_n2889_));
AND2X2 AND2X2_1081 ( .A(_abc_15497_new_n2889_), .B(digest_update), .Y(_abc_15497_new_n2890_));
AND2X2 AND2X2_1082 ( .A(_abc_15497_new_n2888_), .B(_abc_15497_new_n2884_), .Y(_abc_15497_new_n2892_));
AND2X2 AND2X2_1083 ( .A(\digest[141] ), .B(a_reg_13_), .Y(_abc_15497_new_n2895_));
AND2X2 AND2X2_1084 ( .A(_abc_15497_new_n2896_), .B(_abc_15497_new_n2894_), .Y(_abc_15497_new_n2897_));
AND2X2 AND2X2_1085 ( .A(_abc_15497_new_n2898_), .B(_abc_15497_new_n2900_), .Y(_abc_15497_new_n2901_));
AND2X2 AND2X2_1086 ( .A(_abc_15497_new_n2901_), .B(digest_update), .Y(_abc_15497_new_n2902_));
AND2X2 AND2X2_1087 ( .A(_abc_15497_new_n2903_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n2904_));
AND2X2 AND2X2_1088 ( .A(_abc_15497_new_n701_), .B(\digest[142] ), .Y(_abc_15497_new_n2906_));
AND2X2 AND2X2_1089 ( .A(\digest[142] ), .B(a_reg_14_), .Y(_abc_15497_new_n2908_));
AND2X2 AND2X2_109 ( .A(_abc_15497_new_n901_), .B(_abc_15497_new_n905_), .Y(_abc_15497_new_n907_));
AND2X2 AND2X2_1090 ( .A(_abc_15497_new_n2909_), .B(_abc_15497_new_n2907_), .Y(_abc_15497_new_n2910_));
AND2X2 AND2X2_1091 ( .A(_abc_15497_new_n2884_), .B(_abc_15497_new_n2896_), .Y(_abc_15497_new_n2912_));
AND2X2 AND2X2_1092 ( .A(_abc_15497_new_n2888_), .B(_abc_15497_new_n2912_), .Y(_abc_15497_new_n2913_));
AND2X2 AND2X2_1093 ( .A(_abc_15497_new_n2915_), .B(_abc_15497_new_n2910_), .Y(_abc_15497_new_n2917_));
AND2X2 AND2X2_1094 ( .A(_abc_15497_new_n2918_), .B(_abc_15497_new_n2916_), .Y(_abc_15497_new_n2919_));
AND2X2 AND2X2_1095 ( .A(_abc_15497_new_n2919_), .B(digest_update), .Y(_abc_15497_new_n2920_));
AND2X2 AND2X2_1096 ( .A(_abc_15497_new_n701_), .B(\digest[143] ), .Y(_abc_15497_new_n2922_));
AND2X2 AND2X2_1097 ( .A(_abc_15497_new_n2918_), .B(_abc_15497_new_n2909_), .Y(_abc_15497_new_n2923_));
AND2X2 AND2X2_1098 ( .A(\digest[143] ), .B(a_reg_15_), .Y(_abc_15497_new_n2926_));
AND2X2 AND2X2_1099 ( .A(_abc_15497_new_n2927_), .B(_abc_15497_new_n2925_), .Y(_abc_15497_new_n2928_));
AND2X2 AND2X2_11 ( .A(_abc_15497_new_n714_), .B(_abc_15497_new_n717_), .Y(_abc_15497_new_n718_));
AND2X2 AND2X2_110 ( .A(_abc_15497_new_n908_), .B(_abc_15497_new_n906_), .Y(_abc_15497_new_n909_));
AND2X2 AND2X2_1100 ( .A(_abc_15497_new_n2931_), .B(digest_update), .Y(_abc_15497_new_n2932_));
AND2X2 AND2X2_1101 ( .A(_abc_15497_new_n2932_), .B(_abc_15497_new_n2929_), .Y(_abc_15497_new_n2933_));
AND2X2 AND2X2_1102 ( .A(_abc_15497_new_n2928_), .B(_abc_15497_new_n2908_), .Y(_abc_15497_new_n2935_));
AND2X2 AND2X2_1103 ( .A(_abc_15497_new_n2910_), .B(_abc_15497_new_n2928_), .Y(_abc_15497_new_n2939_));
AND2X2 AND2X2_1104 ( .A(_abc_15497_new_n2941_), .B(_abc_15497_new_n2937_), .Y(_abc_15497_new_n2942_));
AND2X2 AND2X2_1105 ( .A(_abc_15497_new_n2885_), .B(_abc_15497_new_n2897_), .Y(_abc_15497_new_n2944_));
AND2X2 AND2X2_1106 ( .A(_abc_15497_new_n2944_), .B(_abc_15497_new_n2939_), .Y(_abc_15497_new_n2945_));
AND2X2 AND2X2_1107 ( .A(_abc_15497_new_n2881_), .B(_abc_15497_new_n2945_), .Y(_abc_15497_new_n2946_));
AND2X2 AND2X2_1108 ( .A(\digest[144] ), .B(a_reg_16_), .Y(_abc_15497_new_n2949_));
AND2X2 AND2X2_1109 ( .A(_abc_15497_new_n2950_), .B(_abc_15497_new_n2948_), .Y(_abc_15497_new_n2951_));
AND2X2 AND2X2_111 ( .A(_abc_15497_new_n909_), .B(digest_update), .Y(_abc_15497_new_n910_));
AND2X2 AND2X2_1110 ( .A(_abc_15497_new_n2947_), .B(_abc_15497_new_n2951_), .Y(_abc_15497_new_n2953_));
AND2X2 AND2X2_1111 ( .A(_abc_15497_new_n2954_), .B(_abc_15497_new_n2952_), .Y(_abc_15497_new_n2955_));
AND2X2 AND2X2_1112 ( .A(_abc_15497_new_n2955_), .B(digest_update), .Y(_abc_15497_new_n2956_));
AND2X2 AND2X2_1113 ( .A(_abc_15497_new_n2957_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n2958_));
AND2X2 AND2X2_1114 ( .A(_abc_15497_new_n701_), .B(\digest[145] ), .Y(_abc_15497_new_n2960_));
AND2X2 AND2X2_1115 ( .A(\digest[145] ), .B(a_reg_17_), .Y(_abc_15497_new_n2962_));
AND2X2 AND2X2_1116 ( .A(_abc_15497_new_n2963_), .B(_abc_15497_new_n2961_), .Y(_abc_15497_new_n2964_));
AND2X2 AND2X2_1117 ( .A(_abc_15497_new_n2951_), .B(_abc_15497_new_n2964_), .Y(_abc_15497_new_n2967_));
AND2X2 AND2X2_1118 ( .A(_abc_15497_new_n2947_), .B(_abc_15497_new_n2967_), .Y(_abc_15497_new_n2968_));
AND2X2 AND2X2_1119 ( .A(_abc_15497_new_n2964_), .B(_abc_15497_new_n2949_), .Y(_abc_15497_new_n2970_));
AND2X2 AND2X2_112 ( .A(_abc_15497_new_n911_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n912_));
AND2X2 AND2X2_1120 ( .A(_abc_15497_new_n2971_), .B(digest_update), .Y(_abc_15497_new_n2972_));
AND2X2 AND2X2_1121 ( .A(_abc_15497_new_n2969_), .B(_abc_15497_new_n2972_), .Y(_abc_15497_new_n2973_));
AND2X2 AND2X2_1122 ( .A(_abc_15497_new_n2973_), .B(_abc_15497_new_n2966_), .Y(_abc_15497_new_n2974_));
AND2X2 AND2X2_1123 ( .A(_abc_15497_new_n2971_), .B(_abc_15497_new_n2963_), .Y(_abc_15497_new_n2976_));
AND2X2 AND2X2_1124 ( .A(_abc_15497_new_n2969_), .B(_abc_15497_new_n2976_), .Y(_abc_15497_new_n2977_));
AND2X2 AND2X2_1125 ( .A(\digest[146] ), .B(a_reg_18_), .Y(_abc_15497_new_n2980_));
AND2X2 AND2X2_1126 ( .A(_abc_15497_new_n2981_), .B(_abc_15497_new_n2979_), .Y(_abc_15497_new_n2982_));
AND2X2 AND2X2_1127 ( .A(_abc_15497_new_n2978_), .B(_abc_15497_new_n2982_), .Y(_abc_15497_new_n2984_));
AND2X2 AND2X2_1128 ( .A(_abc_15497_new_n2985_), .B(_abc_15497_new_n2983_), .Y(_abc_15497_new_n2986_));
AND2X2 AND2X2_1129 ( .A(_abc_15497_new_n2986_), .B(digest_update), .Y(_abc_15497_new_n2987_));
AND2X2 AND2X2_113 ( .A(_abc_15497_new_n701_), .B(\digest[93] ), .Y(_abc_15497_new_n914_));
AND2X2 AND2X2_1130 ( .A(_abc_15497_new_n2988_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n2989_));
AND2X2 AND2X2_1131 ( .A(_abc_15497_new_n701_), .B(\digest[147] ), .Y(_abc_15497_new_n2991_));
AND2X2 AND2X2_1132 ( .A(_abc_15497_new_n2985_), .B(_abc_15497_new_n2981_), .Y(_abc_15497_new_n2992_));
AND2X2 AND2X2_1133 ( .A(\digest[147] ), .B(a_reg_19_), .Y(_abc_15497_new_n2995_));
AND2X2 AND2X2_1134 ( .A(_abc_15497_new_n2996_), .B(_abc_15497_new_n2994_), .Y(_abc_15497_new_n2997_));
AND2X2 AND2X2_1135 ( .A(_abc_15497_new_n3000_), .B(digest_update), .Y(_abc_15497_new_n3001_));
AND2X2 AND2X2_1136 ( .A(_abc_15497_new_n3001_), .B(_abc_15497_new_n2998_), .Y(_abc_15497_new_n3002_));
AND2X2 AND2X2_1137 ( .A(_abc_15497_new_n701_), .B(\digest[148] ), .Y(_abc_15497_new_n3004_));
AND2X2 AND2X2_1138 ( .A(_abc_15497_new_n2982_), .B(_abc_15497_new_n2997_), .Y(_abc_15497_new_n3005_));
AND2X2 AND2X2_1139 ( .A(_abc_15497_new_n2967_), .B(_abc_15497_new_n3005_), .Y(_abc_15497_new_n3006_));
AND2X2 AND2X2_114 ( .A(_abc_15497_new_n908_), .B(_abc_15497_new_n904_), .Y(_abc_15497_new_n915_));
AND2X2 AND2X2_1140 ( .A(_abc_15497_new_n2947_), .B(_abc_15497_new_n3006_), .Y(_abc_15497_new_n3007_));
AND2X2 AND2X2_1141 ( .A(_abc_15497_new_n3008_), .B(_abc_15497_new_n3005_), .Y(_abc_15497_new_n3009_));
AND2X2 AND2X2_1142 ( .A(_abc_15497_new_n2994_), .B(_abc_15497_new_n2980_), .Y(_abc_15497_new_n3010_));
AND2X2 AND2X2_1143 ( .A(\digest[148] ), .B(a_reg_20_), .Y(_abc_15497_new_n3015_));
AND2X2 AND2X2_1144 ( .A(_abc_15497_new_n3016_), .B(_abc_15497_new_n3014_), .Y(_abc_15497_new_n3017_));
AND2X2 AND2X2_1145 ( .A(_abc_15497_new_n3013_), .B(_abc_15497_new_n3017_), .Y(_abc_15497_new_n3019_));
AND2X2 AND2X2_1146 ( .A(_abc_15497_new_n3020_), .B(_abc_15497_new_n3018_), .Y(_abc_15497_new_n3021_));
AND2X2 AND2X2_1147 ( .A(_abc_15497_new_n3021_), .B(digest_update), .Y(_abc_15497_new_n3022_));
AND2X2 AND2X2_1148 ( .A(_abc_15497_new_n701_), .B(\digest[149] ), .Y(_abc_15497_new_n3024_));
AND2X2 AND2X2_1149 ( .A(\digest[149] ), .B(a_reg_21_), .Y(_abc_15497_new_n3026_));
AND2X2 AND2X2_115 ( .A(\digest[93] ), .B(c_reg_29_), .Y(_abc_15497_new_n918_));
AND2X2 AND2X2_1150 ( .A(_abc_15497_new_n3027_), .B(_abc_15497_new_n3025_), .Y(_abc_15497_new_n3028_));
AND2X2 AND2X2_1151 ( .A(_abc_15497_new_n3017_), .B(_abc_15497_new_n3028_), .Y(_abc_15497_new_n3031_));
AND2X2 AND2X2_1152 ( .A(_abc_15497_new_n3013_), .B(_abc_15497_new_n3031_), .Y(_abc_15497_new_n3032_));
AND2X2 AND2X2_1153 ( .A(_abc_15497_new_n3028_), .B(_abc_15497_new_n3015_), .Y(_abc_15497_new_n3033_));
AND2X2 AND2X2_1154 ( .A(_abc_15497_new_n3035_), .B(digest_update), .Y(_abc_15497_new_n3036_));
AND2X2 AND2X2_1155 ( .A(_abc_15497_new_n3036_), .B(_abc_15497_new_n3030_), .Y(_abc_15497_new_n3037_));
AND2X2 AND2X2_1156 ( .A(_abc_15497_new_n3035_), .B(_abc_15497_new_n3027_), .Y(_abc_15497_new_n3039_));
AND2X2 AND2X2_1157 ( .A(\digest[150] ), .B(a_reg_22_), .Y(_abc_15497_new_n3042_));
AND2X2 AND2X2_1158 ( .A(_abc_15497_new_n3043_), .B(_abc_15497_new_n3041_), .Y(_abc_15497_new_n3044_));
AND2X2 AND2X2_1159 ( .A(_abc_15497_new_n3040_), .B(_abc_15497_new_n3044_), .Y(_abc_15497_new_n3046_));
AND2X2 AND2X2_116 ( .A(_abc_15497_new_n919_), .B(_abc_15497_new_n917_), .Y(_abc_15497_new_n920_));
AND2X2 AND2X2_1160 ( .A(_abc_15497_new_n3047_), .B(_abc_15497_new_n3045_), .Y(_abc_15497_new_n3048_));
AND2X2 AND2X2_1161 ( .A(_abc_15497_new_n3048_), .B(digest_update), .Y(_abc_15497_new_n3049_));
AND2X2 AND2X2_1162 ( .A(_abc_15497_new_n3050_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n3051_));
AND2X2 AND2X2_1163 ( .A(_abc_15497_new_n701_), .B(\digest[151] ), .Y(_abc_15497_new_n3053_));
AND2X2 AND2X2_1164 ( .A(_abc_15497_new_n3047_), .B(_abc_15497_new_n3043_), .Y(_abc_15497_new_n3054_));
AND2X2 AND2X2_1165 ( .A(\digest[151] ), .B(a_reg_23_), .Y(_abc_15497_new_n3057_));
AND2X2 AND2X2_1166 ( .A(_abc_15497_new_n3058_), .B(_abc_15497_new_n3056_), .Y(_abc_15497_new_n3059_));
AND2X2 AND2X2_1167 ( .A(_abc_15497_new_n3062_), .B(digest_update), .Y(_abc_15497_new_n3063_));
AND2X2 AND2X2_1168 ( .A(_abc_15497_new_n3063_), .B(_abc_15497_new_n3060_), .Y(_abc_15497_new_n3064_));
AND2X2 AND2X2_1169 ( .A(_abc_15497_new_n3044_), .B(_abc_15497_new_n3059_), .Y(_abc_15497_new_n3067_));
AND2X2 AND2X2_117 ( .A(_abc_15497_new_n923_), .B(digest_update), .Y(_abc_15497_new_n924_));
AND2X2 AND2X2_1170 ( .A(_abc_15497_new_n3066_), .B(_abc_15497_new_n3067_), .Y(_abc_15497_new_n3068_));
AND2X2 AND2X2_1171 ( .A(_abc_15497_new_n3056_), .B(_abc_15497_new_n3042_), .Y(_abc_15497_new_n3069_));
AND2X2 AND2X2_1172 ( .A(_abc_15497_new_n3031_), .B(_abc_15497_new_n3067_), .Y(_abc_15497_new_n3072_));
AND2X2 AND2X2_1173 ( .A(_abc_15497_new_n3013_), .B(_abc_15497_new_n3072_), .Y(_abc_15497_new_n3073_));
AND2X2 AND2X2_1174 ( .A(\digest[152] ), .B(a_reg_24_), .Y(_abc_15497_new_n3076_));
AND2X2 AND2X2_1175 ( .A(_abc_15497_new_n3077_), .B(_abc_15497_new_n3075_), .Y(_abc_15497_new_n3078_));
AND2X2 AND2X2_1176 ( .A(_abc_15497_new_n3074_), .B(_abc_15497_new_n3078_), .Y(_abc_15497_new_n3080_));
AND2X2 AND2X2_1177 ( .A(_abc_15497_new_n3081_), .B(_abc_15497_new_n3079_), .Y(_abc_15497_new_n3082_));
AND2X2 AND2X2_1178 ( .A(_abc_15497_new_n3082_), .B(digest_update), .Y(_abc_15497_new_n3083_));
AND2X2 AND2X2_1179 ( .A(_abc_15497_new_n3084_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n3085_));
AND2X2 AND2X2_118 ( .A(_abc_15497_new_n924_), .B(_abc_15497_new_n921_), .Y(_abc_15497_new_n925_));
AND2X2 AND2X2_1180 ( .A(_abc_15497_new_n3081_), .B(_abc_15497_new_n3077_), .Y(_abc_15497_new_n3087_));
AND2X2 AND2X2_1181 ( .A(\digest[153] ), .B(a_reg_25_), .Y(_abc_15497_new_n3090_));
AND2X2 AND2X2_1182 ( .A(_abc_15497_new_n3091_), .B(_abc_15497_new_n3089_), .Y(_abc_15497_new_n3092_));
AND2X2 AND2X2_1183 ( .A(_abc_15497_new_n3093_), .B(_abc_15497_new_n3095_), .Y(_abc_15497_new_n3096_));
AND2X2 AND2X2_1184 ( .A(_abc_15497_new_n3096_), .B(digest_update), .Y(_abc_15497_new_n3097_));
AND2X2 AND2X2_1185 ( .A(_abc_15497_new_n3098_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n3099_));
AND2X2 AND2X2_1186 ( .A(_abc_15497_new_n3078_), .B(_abc_15497_new_n3092_), .Y(_abc_15497_new_n3101_));
AND2X2 AND2X2_1187 ( .A(_abc_15497_new_n3074_), .B(_abc_15497_new_n3101_), .Y(_abc_15497_new_n3102_));
AND2X2 AND2X2_1188 ( .A(_abc_15497_new_n3089_), .B(_abc_15497_new_n3076_), .Y(_abc_15497_new_n3103_));
AND2X2 AND2X2_1189 ( .A(\digest[154] ), .B(a_reg_26_), .Y(_abc_15497_new_n3107_));
AND2X2 AND2X2_119 ( .A(_abc_15497_new_n701_), .B(\digest[94] ), .Y(_abc_15497_new_n927_));
AND2X2 AND2X2_1190 ( .A(_abc_15497_new_n3108_), .B(_abc_15497_new_n3106_), .Y(_abc_15497_new_n3109_));
AND2X2 AND2X2_1191 ( .A(_abc_15497_new_n3105_), .B(_abc_15497_new_n3109_), .Y(_abc_15497_new_n3111_));
AND2X2 AND2X2_1192 ( .A(_abc_15497_new_n3112_), .B(_abc_15497_new_n3110_), .Y(_abc_15497_new_n3113_));
AND2X2 AND2X2_1193 ( .A(_abc_15497_new_n3113_), .B(digest_update), .Y(_abc_15497_new_n3114_));
AND2X2 AND2X2_1194 ( .A(_abc_15497_new_n3115_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n3116_));
AND2X2 AND2X2_1195 ( .A(_abc_15497_new_n701_), .B(\digest[155] ), .Y(_abc_15497_new_n3118_));
AND2X2 AND2X2_1196 ( .A(\digest[155] ), .B(a_reg_27_), .Y(_abc_15497_new_n3120_));
AND2X2 AND2X2_1197 ( .A(_abc_15497_new_n3121_), .B(_abc_15497_new_n3119_), .Y(_abc_15497_new_n3122_));
AND2X2 AND2X2_1198 ( .A(_abc_15497_new_n3112_), .B(_abc_15497_new_n3108_), .Y(_abc_15497_new_n3126_));
AND2X2 AND2X2_1199 ( .A(_abc_15497_new_n3127_), .B(_abc_15497_new_n3124_), .Y(_abc_15497_new_n3128_));
AND2X2 AND2X2_12 ( .A(_abc_15497_new_n720_), .B(_abc_15497_new_n714_), .Y(_abc_15497_new_n721_));
AND2X2 AND2X2_120 ( .A(\digest[94] ), .B(c_reg_30_), .Y(_abc_15497_new_n928_));
AND2X2 AND2X2_1200 ( .A(_abc_15497_new_n3128_), .B(digest_update), .Y(_abc_15497_new_n3129_));
AND2X2 AND2X2_1201 ( .A(_abc_15497_new_n701_), .B(\digest[156] ), .Y(_abc_15497_new_n3131_));
AND2X2 AND2X2_1202 ( .A(_abc_15497_new_n3109_), .B(_abc_15497_new_n3122_), .Y(_abc_15497_new_n3132_));
AND2X2 AND2X2_1203 ( .A(_abc_15497_new_n3101_), .B(_abc_15497_new_n3132_), .Y(_abc_15497_new_n3133_));
AND2X2 AND2X2_1204 ( .A(_abc_15497_new_n3074_), .B(_abc_15497_new_n3133_), .Y(_abc_15497_new_n3134_));
AND2X2 AND2X2_1205 ( .A(_abc_15497_new_n3122_), .B(_abc_15497_new_n3107_), .Y(_abc_15497_new_n3135_));
AND2X2 AND2X2_1206 ( .A(_abc_15497_new_n3136_), .B(_abc_15497_new_n3121_), .Y(_abc_15497_new_n3137_));
AND2X2 AND2X2_1207 ( .A(_abc_15497_new_n3132_), .B(_abc_15497_new_n3104_), .Y(_abc_15497_new_n3138_));
AND2X2 AND2X2_1208 ( .A(_abc_15497_new_n3139_), .B(_abc_15497_new_n3137_), .Y(_abc_15497_new_n3140_));
AND2X2 AND2X2_1209 ( .A(\digest[156] ), .B(a_reg_28_), .Y(_abc_15497_new_n3144_));
AND2X2 AND2X2_121 ( .A(_abc_15497_new_n929_), .B(_abc_15497_new_n930_), .Y(_abc_15497_new_n931_));
AND2X2 AND2X2_1210 ( .A(_abc_15497_new_n3145_), .B(_abc_15497_new_n3143_), .Y(_abc_15497_new_n3146_));
AND2X2 AND2X2_1211 ( .A(_abc_15497_new_n3142_), .B(_abc_15497_new_n3146_), .Y(_abc_15497_new_n3148_));
AND2X2 AND2X2_1212 ( .A(_abc_15497_new_n3149_), .B(_abc_15497_new_n3147_), .Y(_abc_15497_new_n3150_));
AND2X2 AND2X2_1213 ( .A(_abc_15497_new_n3150_), .B(digest_update), .Y(_abc_15497_new_n3151_));
AND2X2 AND2X2_1214 ( .A(_abc_15497_new_n3149_), .B(_abc_15497_new_n3145_), .Y(_abc_15497_new_n3153_));
AND2X2 AND2X2_1215 ( .A(\digest[157] ), .B(a_reg_29_), .Y(_abc_15497_new_n3155_));
AND2X2 AND2X2_1216 ( .A(_abc_15497_new_n3156_), .B(_abc_15497_new_n3154_), .Y(_abc_15497_new_n3157_));
AND2X2 AND2X2_1217 ( .A(_abc_15497_new_n3161_), .B(digest_update), .Y(_abc_15497_new_n3162_));
AND2X2 AND2X2_1218 ( .A(_abc_15497_new_n3162_), .B(_abc_15497_new_n3159_), .Y(_abc_15497_new_n3163_));
AND2X2 AND2X2_1219 ( .A(_abc_15497_new_n3164_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n3165_));
AND2X2 AND2X2_122 ( .A(_abc_15497_new_n920_), .B(_abc_15497_new_n903_), .Y(_abc_15497_new_n933_));
AND2X2 AND2X2_1220 ( .A(\digest[158] ), .B(a_reg_30_), .Y(_abc_15497_new_n3168_));
AND2X2 AND2X2_1221 ( .A(_abc_15497_new_n3169_), .B(_abc_15497_new_n3167_), .Y(_abc_15497_new_n3170_));
AND2X2 AND2X2_1222 ( .A(_abc_15497_new_n3157_), .B(_abc_15497_new_n3144_), .Y(_abc_15497_new_n3171_));
AND2X2 AND2X2_1223 ( .A(_abc_15497_new_n3146_), .B(_abc_15497_new_n3157_), .Y(_abc_15497_new_n3173_));
AND2X2 AND2X2_1224 ( .A(_abc_15497_new_n3142_), .B(_abc_15497_new_n3173_), .Y(_abc_15497_new_n3174_));
AND2X2 AND2X2_1225 ( .A(_abc_15497_new_n3175_), .B(_abc_15497_new_n3170_), .Y(_abc_15497_new_n3177_));
AND2X2 AND2X2_1226 ( .A(_abc_15497_new_n3178_), .B(_abc_15497_new_n3176_), .Y(_abc_15497_new_n3179_));
AND2X2 AND2X2_1227 ( .A(_abc_15497_new_n3179_), .B(digest_update), .Y(_abc_15497_new_n3180_));
AND2X2 AND2X2_1228 ( .A(_abc_15497_new_n3181_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n3182_));
AND2X2 AND2X2_1229 ( .A(_abc_15497_new_n701_), .B(\digest[159] ), .Y(_abc_15497_new_n3184_));
AND2X2 AND2X2_123 ( .A(_abc_15497_new_n951_), .B(_abc_15497_new_n820_), .Y(_abc_15497_new_n952_));
AND2X2 AND2X2_1230 ( .A(\digest[159] ), .B(a_reg_31_), .Y(_abc_15497_new_n3188_));
AND2X2 AND2X2_1231 ( .A(_abc_15497_new_n3189_), .B(_abc_15497_new_n3187_), .Y(_abc_15497_new_n3190_));
AND2X2 AND2X2_1232 ( .A(_abc_15497_new_n3193_), .B(digest_update), .Y(_abc_15497_new_n3194_));
AND2X2 AND2X2_1233 ( .A(_abc_15497_new_n3194_), .B(_abc_15497_new_n3192_), .Y(_abc_15497_new_n3195_));
AND2X2 AND2X2_1234 ( .A(_abc_15497_new_n2010_), .B(b_reg_0_), .Y(_abc_15497_new_n3197_));
AND2X2 AND2X2_1235 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n2192_), .Y(_abc_15497_new_n3198_));
AND2X2 AND2X2_1236 ( .A(round_ctr_inc), .B(a_reg_0_), .Y(_abc_15497_new_n3199_));
AND2X2 AND2X2_1237 ( .A(_abc_15497_new_n2010_), .B(b_reg_1_), .Y(_abc_15497_new_n3202_));
AND2X2 AND2X2_1238 ( .A(_abc_15497_new_n700_), .B(\digest[97] ), .Y(_abc_15497_new_n3203_));
AND2X2 AND2X2_1239 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3203_), .Y(_abc_15497_new_n3204_));
AND2X2 AND2X2_124 ( .A(_abc_15497_new_n954_), .B(_abc_15497_new_n825_), .Y(_abc_15497_new_n955_));
AND2X2 AND2X2_1240 ( .A(round_ctr_inc), .B(a_reg_1_), .Y(_abc_15497_new_n3205_));
AND2X2 AND2X2_1241 ( .A(_abc_15497_new_n2010_), .B(b_reg_2_), .Y(_abc_15497_new_n3208_));
AND2X2 AND2X2_1242 ( .A(_abc_15497_new_n700_), .B(\digest[98] ), .Y(_abc_15497_new_n3209_));
AND2X2 AND2X2_1243 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3209_), .Y(_abc_15497_new_n3210_));
AND2X2 AND2X2_1244 ( .A(round_ctr_inc), .B(a_reg_2_), .Y(_abc_15497_new_n3211_));
AND2X2 AND2X2_1245 ( .A(_abc_15497_new_n2010_), .B(b_reg_3_), .Y(_abc_15497_new_n3214_));
AND2X2 AND2X2_1246 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n2233_), .Y(_abc_15497_new_n3215_));
AND2X2 AND2X2_1247 ( .A(round_ctr_inc), .B(a_reg_3_), .Y(_abc_15497_new_n3216_));
AND2X2 AND2X2_1248 ( .A(_abc_15497_new_n2010_), .B(b_reg_4_), .Y(_abc_15497_new_n3219_));
AND2X2 AND2X2_1249 ( .A(_abc_15497_new_n700_), .B(\digest[100] ), .Y(_abc_15497_new_n3220_));
AND2X2 AND2X2_125 ( .A(_abc_15497_new_n956_), .B(_abc_15497_new_n946_), .Y(_abc_15497_new_n957_));
AND2X2 AND2X2_1250 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3220_), .Y(_abc_15497_new_n3221_));
AND2X2 AND2X2_1251 ( .A(round_ctr_inc), .B(a_reg_4_), .Y(_abc_15497_new_n3222_));
AND2X2 AND2X2_1252 ( .A(_abc_15497_new_n2010_), .B(b_reg_5_), .Y(_abc_15497_new_n3225_));
AND2X2 AND2X2_1253 ( .A(_abc_15497_new_n700_), .B(\digest[101] ), .Y(_abc_15497_new_n3226_));
AND2X2 AND2X2_1254 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3226_), .Y(_abc_15497_new_n3227_));
AND2X2 AND2X2_1255 ( .A(round_ctr_inc), .B(a_reg_5_), .Y(_abc_15497_new_n3228_));
AND2X2 AND2X2_1256 ( .A(_abc_15497_new_n2010_), .B(b_reg_6_), .Y(_abc_15497_new_n3231_));
AND2X2 AND2X2_1257 ( .A(_abc_15497_new_n700_), .B(\digest[102] ), .Y(_abc_15497_new_n3232_));
AND2X2 AND2X2_1258 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3232_), .Y(_abc_15497_new_n3233_));
AND2X2 AND2X2_1259 ( .A(round_ctr_inc), .B(a_reg_6_), .Y(_abc_15497_new_n3234_));
AND2X2 AND2X2_126 ( .A(_abc_15497_new_n959_), .B(_abc_15497_new_n832_), .Y(_abc_15497_new_n960_));
AND2X2 AND2X2_1260 ( .A(_abc_15497_new_n2010_), .B(b_reg_7_), .Y(_abc_15497_new_n3237_));
AND2X2 AND2X2_1261 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n2280_), .Y(_abc_15497_new_n3238_));
AND2X2 AND2X2_1262 ( .A(round_ctr_inc), .B(a_reg_7_), .Y(_abc_15497_new_n3239_));
AND2X2 AND2X2_1263 ( .A(_abc_15497_new_n2010_), .B(b_reg_8_), .Y(_abc_15497_new_n3242_));
AND2X2 AND2X2_1264 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n2306_), .Y(_abc_15497_new_n3243_));
AND2X2 AND2X2_1265 ( .A(round_ctr_inc), .B(a_reg_8_), .Y(_abc_15497_new_n3244_));
AND2X2 AND2X2_1266 ( .A(_abc_15497_new_n2010_), .B(b_reg_9_), .Y(_abc_15497_new_n3247_));
AND2X2 AND2X2_1267 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n2320_), .Y(_abc_15497_new_n3248_));
AND2X2 AND2X2_1268 ( .A(round_ctr_inc), .B(a_reg_9_), .Y(_abc_15497_new_n3249_));
AND2X2 AND2X2_1269 ( .A(_abc_15497_new_n2010_), .B(b_reg_10_), .Y(_abc_15497_new_n3252_));
AND2X2 AND2X2_127 ( .A(_abc_15497_new_n961_), .B(_abc_15497_new_n944_), .Y(_abc_15497_new_n962_));
AND2X2 AND2X2_1270 ( .A(_abc_15497_new_n700_), .B(\digest[106] ), .Y(_abc_15497_new_n3253_));
AND2X2 AND2X2_1271 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3253_), .Y(_abc_15497_new_n3254_));
AND2X2 AND2X2_1272 ( .A(round_ctr_inc), .B(a_reg_10_), .Y(_abc_15497_new_n3255_));
AND2X2 AND2X2_1273 ( .A(_abc_15497_new_n2010_), .B(b_reg_11_), .Y(_abc_15497_new_n3258_));
AND2X2 AND2X2_1274 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n2351_), .Y(_abc_15497_new_n3259_));
AND2X2 AND2X2_1275 ( .A(round_ctr_inc), .B(a_reg_11_), .Y(_abc_15497_new_n3260_));
AND2X2 AND2X2_1276 ( .A(_abc_15497_new_n2010_), .B(b_reg_12_), .Y(_abc_15497_new_n3263_));
AND2X2 AND2X2_1277 ( .A(_abc_15497_new_n700_), .B(\digest[108] ), .Y(_abc_15497_new_n3264_));
AND2X2 AND2X2_1278 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3264_), .Y(_abc_15497_new_n3265_));
AND2X2 AND2X2_1279 ( .A(round_ctr_inc), .B(a_reg_12_), .Y(_abc_15497_new_n3266_));
AND2X2 AND2X2_128 ( .A(_abc_15497_new_n963_), .B(_abc_15497_new_n942_), .Y(_abc_15497_new_n964_));
AND2X2 AND2X2_1280 ( .A(_abc_15497_new_n2010_), .B(b_reg_13_), .Y(_abc_15497_new_n3269_));
AND2X2 AND2X2_1281 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n2384_), .Y(_abc_15497_new_n3270_));
AND2X2 AND2X2_1282 ( .A(round_ctr_inc), .B(a_reg_13_), .Y(_abc_15497_new_n3271_));
AND2X2 AND2X2_1283 ( .A(_abc_15497_new_n2010_), .B(b_reg_14_), .Y(_abc_15497_new_n3274_));
AND2X2 AND2X2_1284 ( .A(_abc_15497_new_n700_), .B(\digest[110] ), .Y(_abc_15497_new_n3275_));
AND2X2 AND2X2_1285 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3275_), .Y(_abc_15497_new_n3276_));
AND2X2 AND2X2_1286 ( .A(round_ctr_inc), .B(a_reg_14_), .Y(_abc_15497_new_n3277_));
AND2X2 AND2X2_1287 ( .A(_abc_15497_new_n2010_), .B(b_reg_15_), .Y(_abc_15497_new_n3280_));
AND2X2 AND2X2_1288 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n2414_), .Y(_abc_15497_new_n3281_));
AND2X2 AND2X2_1289 ( .A(round_ctr_inc), .B(a_reg_15_), .Y(_abc_15497_new_n3282_));
AND2X2 AND2X2_129 ( .A(_abc_15497_new_n966_), .B(_abc_15497_new_n941_), .Y(_abc_15497_new_n967_));
AND2X2 AND2X2_1290 ( .A(_abc_15497_new_n2010_), .B(b_reg_16_), .Y(_abc_15497_new_n3285_));
AND2X2 AND2X2_1291 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n2439_), .Y(_abc_15497_new_n3286_));
AND2X2 AND2X2_1292 ( .A(round_ctr_inc), .B(a_reg_16_), .Y(_abc_15497_new_n3287_));
AND2X2 AND2X2_1293 ( .A(_abc_15497_new_n2010_), .B(b_reg_17_), .Y(_abc_15497_new_n3290_));
AND2X2 AND2X2_1294 ( .A(_abc_15497_new_n700_), .B(\digest[113] ), .Y(_abc_15497_new_n3291_));
AND2X2 AND2X2_1295 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3291_), .Y(_abc_15497_new_n3292_));
AND2X2 AND2X2_1296 ( .A(round_ctr_inc), .B(a_reg_17_), .Y(_abc_15497_new_n3293_));
AND2X2 AND2X2_1297 ( .A(_abc_15497_new_n2010_), .B(b_reg_18_), .Y(_abc_15497_new_n3296_));
AND2X2 AND2X2_1298 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n2470_), .Y(_abc_15497_new_n3297_));
AND2X2 AND2X2_1299 ( .A(round_ctr_inc), .B(a_reg_18_), .Y(_abc_15497_new_n3298_));
AND2X2 AND2X2_13 ( .A(_abc_15497_new_n703_), .B(_abc_15497_new_n707_), .Y(_abc_15497_new_n723_));
AND2X2 AND2X2_130 ( .A(_abc_15497_new_n968_), .B(_abc_15497_new_n939_), .Y(_abc_15497_new_n969_));
AND2X2 AND2X2_1300 ( .A(_abc_15497_new_n2010_), .B(b_reg_19_), .Y(_abc_15497_new_n3301_));
AND2X2 AND2X2_1301 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n2484_), .Y(_abc_15497_new_n3302_));
AND2X2 AND2X2_1302 ( .A(round_ctr_inc), .B(a_reg_19_), .Y(_abc_15497_new_n3303_));
AND2X2 AND2X2_1303 ( .A(_abc_15497_new_n2010_), .B(b_reg_20_), .Y(_abc_15497_new_n3306_));
AND2X2 AND2X2_1304 ( .A(_abc_15497_new_n700_), .B(\digest[116] ), .Y(_abc_15497_new_n3307_));
AND2X2 AND2X2_1305 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3307_), .Y(_abc_15497_new_n3308_));
AND2X2 AND2X2_1306 ( .A(round_ctr_inc), .B(a_reg_20_), .Y(_abc_15497_new_n3309_));
AND2X2 AND2X2_1307 ( .A(_abc_15497_new_n2010_), .B(b_reg_21_), .Y(_abc_15497_new_n3312_));
AND2X2 AND2X2_1308 ( .A(_abc_15497_new_n700_), .B(\digest[117] ), .Y(_abc_15497_new_n3313_));
AND2X2 AND2X2_1309 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3313_), .Y(_abc_15497_new_n3314_));
AND2X2 AND2X2_131 ( .A(_abc_15497_new_n970_), .B(_abc_15497_new_n937_), .Y(_abc_15497_new_n971_));
AND2X2 AND2X2_1310 ( .A(round_ctr_inc), .B(a_reg_21_), .Y(_abc_15497_new_n3315_));
AND2X2 AND2X2_1311 ( .A(_abc_15497_new_n2010_), .B(b_reg_22_), .Y(_abc_15497_new_n3318_));
AND2X2 AND2X2_1312 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n2535_), .Y(_abc_15497_new_n3319_));
AND2X2 AND2X2_1313 ( .A(round_ctr_inc), .B(a_reg_22_), .Y(_abc_15497_new_n3320_));
AND2X2 AND2X2_1314 ( .A(_abc_15497_new_n2010_), .B(b_reg_23_), .Y(_abc_15497_new_n3323_));
AND2X2 AND2X2_1315 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n2549_), .Y(_abc_15497_new_n3324_));
AND2X2 AND2X2_1316 ( .A(round_ctr_inc), .B(a_reg_23_), .Y(_abc_15497_new_n3325_));
AND2X2 AND2X2_1317 ( .A(_abc_15497_new_n2010_), .B(b_reg_24_), .Y(_abc_15497_new_n3328_));
AND2X2 AND2X2_1318 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n2573_), .Y(_abc_15497_new_n3329_));
AND2X2 AND2X2_1319 ( .A(round_ctr_inc), .B(a_reg_24_), .Y(_abc_15497_new_n3330_));
AND2X2 AND2X2_132 ( .A(_abc_15497_new_n973_), .B(_abc_15497_new_n756_), .Y(_abc_15497_new_n974_));
AND2X2 AND2X2_1320 ( .A(_abc_15497_new_n2010_), .B(b_reg_25_), .Y(_abc_15497_new_n3333_));
AND2X2 AND2X2_1321 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n2587_), .Y(_abc_15497_new_n3334_));
AND2X2 AND2X2_1322 ( .A(round_ctr_inc), .B(a_reg_25_), .Y(_abc_15497_new_n3335_));
AND2X2 AND2X2_1323 ( .A(_abc_15497_new_n2010_), .B(b_reg_26_), .Y(_abc_15497_new_n3338_));
AND2X2 AND2X2_1324 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n2604_), .Y(_abc_15497_new_n3339_));
AND2X2 AND2X2_1325 ( .A(round_ctr_inc), .B(a_reg_26_), .Y(_abc_15497_new_n3340_));
AND2X2 AND2X2_1326 ( .A(_abc_15497_new_n2010_), .B(b_reg_27_), .Y(_abc_15497_new_n3343_));
AND2X2 AND2X2_1327 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n2618_), .Y(_abc_15497_new_n3344_));
AND2X2 AND2X2_1328 ( .A(round_ctr_inc), .B(a_reg_27_), .Y(_abc_15497_new_n3345_));
AND2X2 AND2X2_1329 ( .A(_abc_15497_new_n2010_), .B(b_reg_28_), .Y(_abc_15497_new_n3348_));
AND2X2 AND2X2_133 ( .A(_abc_15497_new_n976_), .B(_abc_15497_new_n977_), .Y(_abc_15497_new_n978_));
AND2X2 AND2X2_1330 ( .A(_abc_15497_new_n700_), .B(\digest[124] ), .Y(_abc_15497_new_n3349_));
AND2X2 AND2X2_1331 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3349_), .Y(_abc_15497_new_n3350_));
AND2X2 AND2X2_1332 ( .A(round_ctr_inc), .B(a_reg_28_), .Y(_abc_15497_new_n3351_));
AND2X2 AND2X2_1333 ( .A(_abc_15497_new_n2010_), .B(b_reg_29_), .Y(_abc_15497_new_n3354_));
AND2X2 AND2X2_1334 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n2637_), .Y(_abc_15497_new_n3355_));
AND2X2 AND2X2_1335 ( .A(round_ctr_inc), .B(a_reg_29_), .Y(_abc_15497_new_n3356_));
AND2X2 AND2X2_1336 ( .A(_abc_15497_new_n2010_), .B(b_reg_30_), .Y(_abc_15497_new_n3359_));
AND2X2 AND2X2_1337 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n2691_), .Y(_abc_15497_new_n3360_));
AND2X2 AND2X2_1338 ( .A(round_ctr_inc), .B(a_reg_30_), .Y(_abc_15497_new_n3361_));
AND2X2 AND2X2_1339 ( .A(_abc_15497_new_n2010_), .B(b_reg_31_), .Y(_abc_15497_new_n3364_));
AND2X2 AND2X2_134 ( .A(_abc_15497_new_n980_), .B(_abc_15497_new_n936_), .Y(_abc_15497_new_n981_));
AND2X2 AND2X2_1340 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n2707_), .Y(_abc_15497_new_n3365_));
AND2X2 AND2X2_1341 ( .A(round_ctr_inc), .B(a_reg_31_), .Y(_abc_15497_new_n3366_));
AND2X2 AND2X2_1342 ( .A(_abc_15497_new_n2010_), .B(d_reg_0_), .Y(_abc_15497_new_n3369_));
AND2X2 AND2X2_1343 ( .A(_abc_15497_new_n700_), .B(\digest[32] ), .Y(_abc_15497_new_n3370_));
AND2X2 AND2X2_1344 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3370_), .Y(_abc_15497_new_n3371_));
AND2X2 AND2X2_1345 ( .A(round_ctr_inc), .B(c_reg_0_), .Y(_abc_15497_new_n3372_));
AND2X2 AND2X2_1346 ( .A(_abc_15497_new_n2010_), .B(d_reg_1_), .Y(_abc_15497_new_n3375_));
AND2X2 AND2X2_1347 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n1545_), .Y(_abc_15497_new_n3376_));
AND2X2 AND2X2_1348 ( .A(round_ctr_inc), .B(c_reg_1_), .Y(_abc_15497_new_n3377_));
AND2X2 AND2X2_1349 ( .A(_abc_15497_new_n2010_), .B(d_reg_2_), .Y(_abc_15497_new_n3380_));
AND2X2 AND2X2_135 ( .A(_abc_15497_new_n905_), .B(_abc_15497_new_n920_), .Y(_abc_15497_new_n982_));
AND2X2 AND2X2_1350 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n1558_), .Y(_abc_15497_new_n3381_));
AND2X2 AND2X2_1351 ( .A(round_ctr_inc), .B(c_reg_2_), .Y(_abc_15497_new_n3382_));
AND2X2 AND2X2_1352 ( .A(_abc_15497_new_n2010_), .B(d_reg_3_), .Y(_abc_15497_new_n3385_));
AND2X2 AND2X2_1353 ( .A(_abc_15497_new_n700_), .B(\digest[35] ), .Y(_abc_15497_new_n3386_));
AND2X2 AND2X2_1354 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3386_), .Y(_abc_15497_new_n3387_));
AND2X2 AND2X2_1355 ( .A(round_ctr_inc), .B(c_reg_3_), .Y(_abc_15497_new_n3388_));
AND2X2 AND2X2_1356 ( .A(_abc_15497_new_n2010_), .B(d_reg_4_), .Y(_abc_15497_new_n3391_));
AND2X2 AND2X2_1357 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n1585_), .Y(_abc_15497_new_n3392_));
AND2X2 AND2X2_1358 ( .A(round_ctr_inc), .B(c_reg_4_), .Y(_abc_15497_new_n3393_));
AND2X2 AND2X2_1359 ( .A(_abc_15497_new_n2010_), .B(d_reg_5_), .Y(_abc_15497_new_n3396_));
AND2X2 AND2X2_136 ( .A(_abc_15497_new_n984_), .B(_abc_15497_new_n935_), .Y(_abc_15497_new_n985_));
AND2X2 AND2X2_1360 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n1598_), .Y(_abc_15497_new_n3397_));
AND2X2 AND2X2_1361 ( .A(round_ctr_inc), .B(c_reg_5_), .Y(_abc_15497_new_n3398_));
AND2X2 AND2X2_1362 ( .A(_abc_15497_new_n2010_), .B(d_reg_6_), .Y(_abc_15497_new_n3401_));
AND2X2 AND2X2_1363 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n1611_), .Y(_abc_15497_new_n3402_));
AND2X2 AND2X2_1364 ( .A(round_ctr_inc), .B(c_reg_6_), .Y(_abc_15497_new_n3403_));
AND2X2 AND2X2_1365 ( .A(_abc_15497_new_n2010_), .B(d_reg_7_), .Y(_abc_15497_new_n3406_));
AND2X2 AND2X2_1366 ( .A(_abc_15497_new_n700_), .B(\digest[39] ), .Y(_abc_15497_new_n3407_));
AND2X2 AND2X2_1367 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3407_), .Y(_abc_15497_new_n3408_));
AND2X2 AND2X2_1368 ( .A(round_ctr_inc), .B(c_reg_7_), .Y(_abc_15497_new_n3409_));
AND2X2 AND2X2_1369 ( .A(_abc_15497_new_n2010_), .B(d_reg_8_), .Y(_abc_15497_new_n3412_));
AND2X2 AND2X2_137 ( .A(_abc_15497_new_n901_), .B(_abc_15497_new_n982_), .Y(_abc_15497_new_n987_));
AND2X2 AND2X2_1370 ( .A(_abc_15497_new_n700_), .B(\digest[40] ), .Y(_abc_15497_new_n3413_));
AND2X2 AND2X2_1371 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3413_), .Y(_abc_15497_new_n3414_));
AND2X2 AND2X2_1372 ( .A(round_ctr_inc), .B(c_reg_8_), .Y(_abc_15497_new_n3415_));
AND2X2 AND2X2_1373 ( .A(_abc_15497_new_n2010_), .B(d_reg_9_), .Y(_abc_15497_new_n3418_));
AND2X2 AND2X2_1374 ( .A(_abc_15497_new_n700_), .B(\digest[41] ), .Y(_abc_15497_new_n3419_));
AND2X2 AND2X2_1375 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3419_), .Y(_abc_15497_new_n3420_));
AND2X2 AND2X2_1376 ( .A(round_ctr_inc), .B(c_reg_9_), .Y(_abc_15497_new_n3421_));
AND2X2 AND2X2_1377 ( .A(_abc_15497_new_n2010_), .B(d_reg_10_), .Y(_abc_15497_new_n3424_));
AND2X2 AND2X2_1378 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n1666_), .Y(_abc_15497_new_n3425_));
AND2X2 AND2X2_1379 ( .A(round_ctr_inc), .B(c_reg_10_), .Y(_abc_15497_new_n3426_));
AND2X2 AND2X2_138 ( .A(_abc_15497_new_n989_), .B(digest_update), .Y(_abc_15497_new_n990_));
AND2X2 AND2X2_1380 ( .A(_abc_15497_new_n2010_), .B(d_reg_11_), .Y(_abc_15497_new_n3429_));
AND2X2 AND2X2_1381 ( .A(_abc_15497_new_n700_), .B(\digest[43] ), .Y(_abc_15497_new_n3430_));
AND2X2 AND2X2_1382 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3430_), .Y(_abc_15497_new_n3431_));
AND2X2 AND2X2_1383 ( .A(round_ctr_inc), .B(c_reg_11_), .Y(_abc_15497_new_n3432_));
AND2X2 AND2X2_1384 ( .A(_abc_15497_new_n2010_), .B(d_reg_12_), .Y(_abc_15497_new_n3435_));
AND2X2 AND2X2_1385 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n1700_), .Y(_abc_15497_new_n3436_));
AND2X2 AND2X2_1386 ( .A(round_ctr_inc), .B(c_reg_12_), .Y(_abc_15497_new_n3437_));
AND2X2 AND2X2_1387 ( .A(_abc_15497_new_n2010_), .B(d_reg_13_), .Y(_abc_15497_new_n3440_));
AND2X2 AND2X2_1388 ( .A(_abc_15497_new_n700_), .B(\digest[45] ), .Y(_abc_15497_new_n3441_));
AND2X2 AND2X2_1389 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3441_), .Y(_abc_15497_new_n3442_));
AND2X2 AND2X2_139 ( .A(_abc_15497_new_n990_), .B(_abc_15497_new_n986_), .Y(_abc_15497_new_n991_));
AND2X2 AND2X2_1390 ( .A(round_ctr_inc), .B(c_reg_13_), .Y(_abc_15497_new_n3443_));
AND2X2 AND2X2_1391 ( .A(_abc_15497_new_n2010_), .B(d_reg_14_), .Y(_abc_15497_new_n3446_));
AND2X2 AND2X2_1392 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n1731_), .Y(_abc_15497_new_n3447_));
AND2X2 AND2X2_1393 ( .A(round_ctr_inc), .B(c_reg_14_), .Y(_abc_15497_new_n3448_));
AND2X2 AND2X2_1394 ( .A(_abc_15497_new_n2010_), .B(d_reg_15_), .Y(_abc_15497_new_n3451_));
AND2X2 AND2X2_1395 ( .A(_abc_15497_new_n700_), .B(\digest[47] ), .Y(_abc_15497_new_n3452_));
AND2X2 AND2X2_1396 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3452_), .Y(_abc_15497_new_n3453_));
AND2X2 AND2X2_1397 ( .A(round_ctr_inc), .B(c_reg_15_), .Y(_abc_15497_new_n3454_));
AND2X2 AND2X2_1398 ( .A(_abc_15497_new_n2010_), .B(d_reg_16_), .Y(_abc_15497_new_n3457_));
AND2X2 AND2X2_1399 ( .A(_abc_15497_new_n700_), .B(\digest[48] ), .Y(_abc_15497_new_n3458_));
AND2X2 AND2X2_14 ( .A(_abc_15497_new_n722_), .B(_abc_15497_new_n725_), .Y(_abc_15497_new_n726_));
AND2X2 AND2X2_140 ( .A(_abc_15497_new_n988_), .B(_abc_15497_new_n931_), .Y(_abc_15497_new_n993_));
AND2X2 AND2X2_1400 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3458_), .Y(_abc_15497_new_n3459_));
AND2X2 AND2X2_1401 ( .A(round_ctr_inc), .B(c_reg_16_), .Y(_abc_15497_new_n3460_));
AND2X2 AND2X2_1402 ( .A(_abc_15497_new_n2010_), .B(d_reg_17_), .Y(_abc_15497_new_n3463_));
AND2X2 AND2X2_1403 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n1780_), .Y(_abc_15497_new_n3464_));
AND2X2 AND2X2_1404 ( .A(round_ctr_inc), .B(c_reg_17_), .Y(_abc_15497_new_n3465_));
AND2X2 AND2X2_1405 ( .A(_abc_15497_new_n2010_), .B(d_reg_18_), .Y(_abc_15497_new_n3468_));
AND2X2 AND2X2_1406 ( .A(_abc_15497_new_n700_), .B(\digest[50] ), .Y(_abc_15497_new_n3469_));
AND2X2 AND2X2_1407 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3469_), .Y(_abc_15497_new_n3470_));
AND2X2 AND2X2_1408 ( .A(round_ctr_inc), .B(c_reg_18_), .Y(_abc_15497_new_n3471_));
AND2X2 AND2X2_1409 ( .A(_abc_15497_new_n2010_), .B(d_reg_19_), .Y(_abc_15497_new_n3474_));
AND2X2 AND2X2_141 ( .A(_abc_15497_new_n996_), .B(_abc_15497_new_n998_), .Y(_abc_15497_new_n999_));
AND2X2 AND2X2_1410 ( .A(_abc_15497_new_n700_), .B(\digest[51] ), .Y(_abc_15497_new_n3475_));
AND2X2 AND2X2_1411 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3475_), .Y(_abc_15497_new_n3476_));
AND2X2 AND2X2_1412 ( .A(round_ctr_inc), .B(c_reg_19_), .Y(_abc_15497_new_n3477_));
AND2X2 AND2X2_1413 ( .A(_abc_15497_new_n2010_), .B(d_reg_20_), .Y(_abc_15497_new_n3480_));
AND2X2 AND2X2_1414 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n1829_), .Y(_abc_15497_new_n3481_));
AND2X2 AND2X2_1415 ( .A(round_ctr_inc), .B(c_reg_20_), .Y(_abc_15497_new_n3482_));
AND2X2 AND2X2_1416 ( .A(_abc_15497_new_n2010_), .B(d_reg_21_), .Y(_abc_15497_new_n3485_));
AND2X2 AND2X2_1417 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n1843_), .Y(_abc_15497_new_n3486_));
AND2X2 AND2X2_1418 ( .A(round_ctr_inc), .B(c_reg_21_), .Y(_abc_15497_new_n3487_));
AND2X2 AND2X2_1419 ( .A(_abc_15497_new_n2010_), .B(d_reg_22_), .Y(_abc_15497_new_n3490_));
AND2X2 AND2X2_142 ( .A(_abc_15497_new_n986_), .B(_abc_15497_new_n929_), .Y(_abc_15497_new_n1002_));
AND2X2 AND2X2_1420 ( .A(_abc_15497_new_n700_), .B(\digest[54] ), .Y(_abc_15497_new_n3491_));
AND2X2 AND2X2_1421 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3491_), .Y(_abc_15497_new_n3492_));
AND2X2 AND2X2_1422 ( .A(round_ctr_inc), .B(c_reg_22_), .Y(_abc_15497_new_n3493_));
AND2X2 AND2X2_1423 ( .A(_abc_15497_new_n2010_), .B(d_reg_23_), .Y(_abc_15497_new_n3496_));
AND2X2 AND2X2_1424 ( .A(_abc_15497_new_n700_), .B(\digest[55] ), .Y(_abc_15497_new_n3497_));
AND2X2 AND2X2_1425 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3497_), .Y(_abc_15497_new_n3498_));
AND2X2 AND2X2_1426 ( .A(round_ctr_inc), .B(c_reg_23_), .Y(_abc_15497_new_n3499_));
AND2X2 AND2X2_1427 ( .A(_abc_15497_new_n2010_), .B(d_reg_24_), .Y(_abc_15497_new_n3502_));
AND2X2 AND2X2_1428 ( .A(_abc_15497_new_n700_), .B(\digest[56] ), .Y(_abc_15497_new_n3503_));
AND2X2 AND2X2_1429 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3503_), .Y(_abc_15497_new_n3504_));
AND2X2 AND2X2_143 ( .A(_abc_15497_new_n1003_), .B(_abc_15497_new_n1001_), .Y(_abc_15497_new_n1004_));
AND2X2 AND2X2_1430 ( .A(round_ctr_inc), .B(c_reg_24_), .Y(_abc_15497_new_n3505_));
AND2X2 AND2X2_1431 ( .A(_abc_15497_new_n2010_), .B(d_reg_25_), .Y(_abc_15497_new_n3508_));
AND2X2 AND2X2_1432 ( .A(_abc_15497_new_n700_), .B(\digest[57] ), .Y(_abc_15497_new_n3509_));
AND2X2 AND2X2_1433 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3509_), .Y(_abc_15497_new_n3510_));
AND2X2 AND2X2_1434 ( .A(round_ctr_inc), .B(c_reg_25_), .Y(_abc_15497_new_n3511_));
AND2X2 AND2X2_1435 ( .A(_abc_15497_new_n2010_), .B(d_reg_26_), .Y(_abc_15497_new_n3514_));
AND2X2 AND2X2_1436 ( .A(_abc_15497_new_n700_), .B(\digest[58] ), .Y(_abc_15497_new_n3515_));
AND2X2 AND2X2_1437 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3515_), .Y(_abc_15497_new_n3516_));
AND2X2 AND2X2_1438 ( .A(c_reg_26_), .B(round_ctr_inc), .Y(_abc_15497_new_n3517_));
AND2X2 AND2X2_1439 ( .A(_abc_15497_new_n2010_), .B(d_reg_27_), .Y(_abc_15497_new_n3520_));
AND2X2 AND2X2_144 ( .A(_abc_15497_new_n1004_), .B(digest_update), .Y(_abc_15497_new_n1005_));
AND2X2 AND2X2_1440 ( .A(_abc_15497_new_n700_), .B(\digest[59] ), .Y(_abc_15497_new_n3521_));
AND2X2 AND2X2_1441 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3521_), .Y(_abc_15497_new_n3522_));
AND2X2 AND2X2_1442 ( .A(c_reg_27_), .B(round_ctr_inc), .Y(_abc_15497_new_n3523_));
AND2X2 AND2X2_1443 ( .A(_abc_15497_new_n2010_), .B(d_reg_28_), .Y(_abc_15497_new_n3526_));
AND2X2 AND2X2_1444 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n1961_), .Y(_abc_15497_new_n3527_));
AND2X2 AND2X2_1445 ( .A(c_reg_28_), .B(round_ctr_inc), .Y(_abc_15497_new_n3528_));
AND2X2 AND2X2_1446 ( .A(_abc_15497_new_n2010_), .B(d_reg_29_), .Y(_abc_15497_new_n3531_));
AND2X2 AND2X2_1447 ( .A(_abc_15497_new_n700_), .B(\digest[61] ), .Y(_abc_15497_new_n3532_));
AND2X2 AND2X2_1448 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3532_), .Y(_abc_15497_new_n3533_));
AND2X2 AND2X2_1449 ( .A(c_reg_29_), .B(round_ctr_inc), .Y(_abc_15497_new_n3534_));
AND2X2 AND2X2_145 ( .A(_abc_15497_new_n1006_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n1007_));
AND2X2 AND2X2_1450 ( .A(_abc_15497_new_n2010_), .B(d_reg_30_), .Y(_abc_15497_new_n3537_));
AND2X2 AND2X2_1451 ( .A(_abc_15497_new_n700_), .B(\digest[62] ), .Y(_abc_15497_new_n3538_));
AND2X2 AND2X2_1452 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3538_), .Y(_abc_15497_new_n3539_));
AND2X2 AND2X2_1453 ( .A(c_reg_30_), .B(round_ctr_inc), .Y(_abc_15497_new_n3540_));
AND2X2 AND2X2_1454 ( .A(_abc_15497_new_n2010_), .B(d_reg_31_), .Y(_abc_15497_new_n3543_));
AND2X2 AND2X2_1455 ( .A(_abc_15497_new_n700_), .B(\digest[63] ), .Y(_abc_15497_new_n3544_));
AND2X2 AND2X2_1456 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3544_), .Y(_abc_15497_new_n3545_));
AND2X2 AND2X2_1457 ( .A(c_reg_31_), .B(round_ctr_inc), .Y(_abc_15497_new_n3546_));
AND2X2 AND2X2_1458 ( .A(_abc_15497_new_n2010_), .B(c_reg_0_), .Y(_abc_15497_new_n3549_));
AND2X2 AND2X2_1459 ( .A(_abc_15497_new_n700_), .B(\digest[64] ), .Y(_abc_15497_new_n3550_));
AND2X2 AND2X2_146 ( .A(e_reg_0_), .B(\digest[0] ), .Y(_abc_15497_new_n1009_));
AND2X2 AND2X2_1460 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3550_), .Y(_abc_15497_new_n3551_));
AND2X2 AND2X2_1461 ( .A(round_ctr_inc), .B(b_reg_2_), .Y(_abc_15497_new_n3552_));
AND2X2 AND2X2_1462 ( .A(_abc_15497_new_n2010_), .B(c_reg_1_), .Y(_abc_15497_new_n3555_));
AND2X2 AND2X2_1463 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3556_), .Y(_abc_15497_new_n3557_));
AND2X2 AND2X2_1464 ( .A(round_ctr_inc), .B(b_reg_3_), .Y(_abc_15497_new_n3558_));
AND2X2 AND2X2_1465 ( .A(_abc_15497_new_n2010_), .B(c_reg_2_), .Y(_abc_15497_new_n3561_));
AND2X2 AND2X2_1466 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3562_), .Y(_abc_15497_new_n3563_));
AND2X2 AND2X2_1467 ( .A(round_ctr_inc), .B(b_reg_4_), .Y(_abc_15497_new_n3564_));
AND2X2 AND2X2_1468 ( .A(_abc_15497_new_n2010_), .B(c_reg_3_), .Y(_abc_15497_new_n3567_));
AND2X2 AND2X2_1469 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3568_), .Y(_abc_15497_new_n3569_));
AND2X2 AND2X2_147 ( .A(_abc_15497_new_n1011_), .B(digest_update), .Y(_abc_15497_new_n1012_));
AND2X2 AND2X2_1470 ( .A(round_ctr_inc), .B(b_reg_5_), .Y(_abc_15497_new_n3570_));
AND2X2 AND2X2_1471 ( .A(_abc_15497_new_n2010_), .B(c_reg_4_), .Y(_abc_15497_new_n3573_));
AND2X2 AND2X2_1472 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3574_), .Y(_abc_15497_new_n3575_));
AND2X2 AND2X2_1473 ( .A(round_ctr_inc), .B(b_reg_6_), .Y(_abc_15497_new_n3576_));
AND2X2 AND2X2_1474 ( .A(_abc_15497_new_n2010_), .B(c_reg_5_), .Y(_abc_15497_new_n3579_));
AND2X2 AND2X2_1475 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3580_), .Y(_abc_15497_new_n3581_));
AND2X2 AND2X2_1476 ( .A(round_ctr_inc), .B(b_reg_7_), .Y(_abc_15497_new_n3582_));
AND2X2 AND2X2_1477 ( .A(_abc_15497_new_n2010_), .B(c_reg_6_), .Y(_abc_15497_new_n3585_));
AND2X2 AND2X2_1478 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3586_), .Y(_abc_15497_new_n3587_));
AND2X2 AND2X2_1479 ( .A(round_ctr_inc), .B(b_reg_8_), .Y(_abc_15497_new_n3588_));
AND2X2 AND2X2_148 ( .A(_abc_15497_new_n1012_), .B(_abc_15497_new_n1010_), .Y(_abc_15497_new_n1013_));
AND2X2 AND2X2_1480 ( .A(_abc_15497_new_n2010_), .B(c_reg_7_), .Y(_abc_15497_new_n3591_));
AND2X2 AND2X2_1481 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3592_), .Y(_abc_15497_new_n3593_));
AND2X2 AND2X2_1482 ( .A(round_ctr_inc), .B(b_reg_9_), .Y(_abc_15497_new_n3594_));
AND2X2 AND2X2_1483 ( .A(_abc_15497_new_n2010_), .B(c_reg_8_), .Y(_abc_15497_new_n3597_));
AND2X2 AND2X2_1484 ( .A(_abc_15497_new_n700_), .B(\digest[72] ), .Y(_abc_15497_new_n3598_));
AND2X2 AND2X2_1485 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3598_), .Y(_abc_15497_new_n3599_));
AND2X2 AND2X2_1486 ( .A(round_ctr_inc), .B(b_reg_10_), .Y(_abc_15497_new_n3600_));
AND2X2 AND2X2_1487 ( .A(_abc_15497_new_n2010_), .B(c_reg_9_), .Y(_abc_15497_new_n3603_));
AND2X2 AND2X2_1488 ( .A(_abc_15497_new_n700_), .B(\digest[73] ), .Y(_abc_15497_new_n3604_));
AND2X2 AND2X2_1489 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3604_), .Y(_abc_15497_new_n3605_));
AND2X2 AND2X2_149 ( .A(_abc_15497_new_n701_), .B(\digest[0] ), .Y(_abc_15497_new_n1014_));
AND2X2 AND2X2_1490 ( .A(round_ctr_inc), .B(b_reg_11_), .Y(_abc_15497_new_n3606_));
AND2X2 AND2X2_1491 ( .A(_abc_15497_new_n2010_), .B(c_reg_10_), .Y(_abc_15497_new_n3609_));
AND2X2 AND2X2_1492 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3610_), .Y(_abc_15497_new_n3611_));
AND2X2 AND2X2_1493 ( .A(round_ctr_inc), .B(b_reg_12_), .Y(_abc_15497_new_n3612_));
AND2X2 AND2X2_1494 ( .A(_abc_15497_new_n2010_), .B(c_reg_11_), .Y(_abc_15497_new_n3615_));
AND2X2 AND2X2_1495 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3616_), .Y(_abc_15497_new_n3617_));
AND2X2 AND2X2_1496 ( .A(round_ctr_inc), .B(b_reg_13_), .Y(_abc_15497_new_n3618_));
AND2X2 AND2X2_1497 ( .A(_abc_15497_new_n2010_), .B(c_reg_12_), .Y(_abc_15497_new_n3621_));
AND2X2 AND2X2_1498 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3622_), .Y(_abc_15497_new_n3623_));
AND2X2 AND2X2_1499 ( .A(round_ctr_inc), .B(b_reg_14_), .Y(_abc_15497_new_n3624_));
AND2X2 AND2X2_15 ( .A(_abc_15497_new_n716_), .B(_abc_15497_new_n727_), .Y(_abc_15497_new_n728_));
AND2X2 AND2X2_150 ( .A(e_reg_1_), .B(\digest[1] ), .Y(_abc_15497_new_n1018_));
AND2X2 AND2X2_1500 ( .A(_abc_15497_new_n2010_), .B(c_reg_13_), .Y(_abc_15497_new_n3627_));
AND2X2 AND2X2_1501 ( .A(_abc_15497_new_n700_), .B(\digest[77] ), .Y(_abc_15497_new_n3628_));
AND2X2 AND2X2_1502 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3628_), .Y(_abc_15497_new_n3629_));
AND2X2 AND2X2_1503 ( .A(round_ctr_inc), .B(b_reg_15_), .Y(_abc_15497_new_n3630_));
AND2X2 AND2X2_1504 ( .A(_abc_15497_new_n2010_), .B(c_reg_14_), .Y(_abc_15497_new_n3633_));
AND2X2 AND2X2_1505 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3634_), .Y(_abc_15497_new_n3635_));
AND2X2 AND2X2_1506 ( .A(round_ctr_inc), .B(b_reg_16_), .Y(_abc_15497_new_n3636_));
AND2X2 AND2X2_1507 ( .A(_abc_15497_new_n2010_), .B(c_reg_15_), .Y(_abc_15497_new_n3639_));
AND2X2 AND2X2_1508 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3640_), .Y(_abc_15497_new_n3641_));
AND2X2 AND2X2_1509 ( .A(round_ctr_inc), .B(b_reg_17_), .Y(_abc_15497_new_n3642_));
AND2X2 AND2X2_151 ( .A(_abc_15497_new_n1021_), .B(_abc_15497_new_n1016_), .Y(_abc_15497_new_n1022_));
AND2X2 AND2X2_1510 ( .A(_abc_15497_new_n2010_), .B(c_reg_16_), .Y(_abc_15497_new_n3645_));
AND2X2 AND2X2_1511 ( .A(_abc_15497_new_n700_), .B(\digest[80] ), .Y(_abc_15497_new_n3646_));
AND2X2 AND2X2_1512 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3646_), .Y(_abc_15497_new_n3647_));
AND2X2 AND2X2_1513 ( .A(round_ctr_inc), .B(b_reg_18_), .Y(_abc_15497_new_n3648_));
AND2X2 AND2X2_1514 ( .A(_abc_15497_new_n2010_), .B(c_reg_17_), .Y(_abc_15497_new_n3651_));
AND2X2 AND2X2_1515 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3652_), .Y(_abc_15497_new_n3653_));
AND2X2 AND2X2_1516 ( .A(round_ctr_inc), .B(b_reg_19_), .Y(_abc_15497_new_n3654_));
AND2X2 AND2X2_1517 ( .A(_abc_15497_new_n2010_), .B(c_reg_18_), .Y(_abc_15497_new_n3657_));
AND2X2 AND2X2_1518 ( .A(_abc_15497_new_n700_), .B(\digest[82] ), .Y(_abc_15497_new_n3658_));
AND2X2 AND2X2_1519 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3658_), .Y(_abc_15497_new_n3659_));
AND2X2 AND2X2_152 ( .A(_abc_15497_new_n1023_), .B(digest_update), .Y(_abc_15497_new_n1024_));
AND2X2 AND2X2_1520 ( .A(round_ctr_inc), .B(b_reg_20_), .Y(_abc_15497_new_n3660_));
AND2X2 AND2X2_1521 ( .A(_abc_15497_new_n2010_), .B(c_reg_19_), .Y(_abc_15497_new_n3663_));
AND2X2 AND2X2_1522 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3664_), .Y(_abc_15497_new_n3665_));
AND2X2 AND2X2_1523 ( .A(round_ctr_inc), .B(b_reg_21_), .Y(_abc_15497_new_n3666_));
AND2X2 AND2X2_1524 ( .A(_abc_15497_new_n2010_), .B(c_reg_20_), .Y(_abc_15497_new_n3669_));
AND2X2 AND2X2_1525 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3670_), .Y(_abc_15497_new_n3671_));
AND2X2 AND2X2_1526 ( .A(round_ctr_inc), .B(b_reg_22_), .Y(_abc_15497_new_n3672_));
AND2X2 AND2X2_1527 ( .A(_abc_15497_new_n2010_), .B(c_reg_21_), .Y(_abc_15497_new_n3675_));
AND2X2 AND2X2_1528 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3676_), .Y(_abc_15497_new_n3677_));
AND2X2 AND2X2_1529 ( .A(round_ctr_inc), .B(b_reg_23_), .Y(_abc_15497_new_n3678_));
AND2X2 AND2X2_153 ( .A(_abc_15497_new_n1024_), .B(_abc_15497_new_n1020_), .Y(_abc_15497_new_n1025_));
AND2X2 AND2X2_1530 ( .A(_abc_15497_new_n2010_), .B(c_reg_22_), .Y(_abc_15497_new_n3681_));
AND2X2 AND2X2_1531 ( .A(_abc_15497_new_n700_), .B(\digest[86] ), .Y(_abc_15497_new_n3682_));
AND2X2 AND2X2_1532 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3682_), .Y(_abc_15497_new_n3683_));
AND2X2 AND2X2_1533 ( .A(round_ctr_inc), .B(b_reg_24_), .Y(_abc_15497_new_n3684_));
AND2X2 AND2X2_1534 ( .A(_abc_15497_new_n2010_), .B(c_reg_23_), .Y(_abc_15497_new_n3687_));
AND2X2 AND2X2_1535 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3688_), .Y(_abc_15497_new_n3689_));
AND2X2 AND2X2_1536 ( .A(round_ctr_inc), .B(b_reg_25_), .Y(_abc_15497_new_n3690_));
AND2X2 AND2X2_1537 ( .A(_abc_15497_new_n2010_), .B(c_reg_24_), .Y(_abc_15497_new_n3693_));
AND2X2 AND2X2_1538 ( .A(_abc_15497_new_n700_), .B(\digest[88] ), .Y(_abc_15497_new_n3694_));
AND2X2 AND2X2_1539 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3694_), .Y(_abc_15497_new_n3695_));
AND2X2 AND2X2_154 ( .A(_abc_15497_new_n701_), .B(\digest[1] ), .Y(_abc_15497_new_n1026_));
AND2X2 AND2X2_1540 ( .A(round_ctr_inc), .B(b_reg_26_), .Y(_abc_15497_new_n3696_));
AND2X2 AND2X2_1541 ( .A(_abc_15497_new_n2010_), .B(c_reg_25_), .Y(_abc_15497_new_n3699_));
AND2X2 AND2X2_1542 ( .A(_abc_15497_new_n700_), .B(\digest[89] ), .Y(_abc_15497_new_n3700_));
AND2X2 AND2X2_1543 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3700_), .Y(_abc_15497_new_n3701_));
AND2X2 AND2X2_1544 ( .A(round_ctr_inc), .B(b_reg_27_), .Y(_abc_15497_new_n3702_));
AND2X2 AND2X2_1545 ( .A(_abc_15497_new_n2010_), .B(c_reg_26_), .Y(_abc_15497_new_n3705_));
AND2X2 AND2X2_1546 ( .A(_abc_15497_new_n700_), .B(\digest[90] ), .Y(_abc_15497_new_n3706_));
AND2X2 AND2X2_1547 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3706_), .Y(_abc_15497_new_n3707_));
AND2X2 AND2X2_1548 ( .A(round_ctr_inc), .B(b_reg_28_), .Y(_abc_15497_new_n3708_));
AND2X2 AND2X2_1549 ( .A(_abc_15497_new_n2010_), .B(c_reg_27_), .Y(_abc_15497_new_n3711_));
AND2X2 AND2X2_155 ( .A(_abc_15497_new_n1020_), .B(_abc_15497_new_n1021_), .Y(_abc_15497_new_n1028_));
AND2X2 AND2X2_1550 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n894_), .Y(_abc_15497_new_n3712_));
AND2X2 AND2X2_1551 ( .A(round_ctr_inc), .B(b_reg_29_), .Y(_abc_15497_new_n3713_));
AND2X2 AND2X2_1552 ( .A(_abc_15497_new_n2010_), .B(c_reg_28_), .Y(_abc_15497_new_n3716_));
AND2X2 AND2X2_1553 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n911_), .Y(_abc_15497_new_n3717_));
AND2X2 AND2X2_1554 ( .A(round_ctr_inc), .B(b_reg_30_), .Y(_abc_15497_new_n3718_));
AND2X2 AND2X2_1555 ( .A(_abc_15497_new_n2010_), .B(c_reg_29_), .Y(_abc_15497_new_n3721_));
AND2X2 AND2X2_1556 ( .A(_abc_15497_new_n700_), .B(\digest[93] ), .Y(_abc_15497_new_n3722_));
AND2X2 AND2X2_1557 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3722_), .Y(_abc_15497_new_n3723_));
AND2X2 AND2X2_1558 ( .A(round_ctr_inc), .B(b_reg_31_), .Y(_abc_15497_new_n3724_));
AND2X2 AND2X2_1559 ( .A(_abc_15497_new_n2010_), .B(c_reg_30_), .Y(_abc_15497_new_n3727_));
AND2X2 AND2X2_156 ( .A(e_reg_2_), .B(\digest[2] ), .Y(_abc_15497_new_n1030_));
AND2X2 AND2X2_1560 ( .A(_abc_15497_new_n700_), .B(\digest[94] ), .Y(_abc_15497_new_n3728_));
AND2X2 AND2X2_1561 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3728_), .Y(_abc_15497_new_n3729_));
AND2X2 AND2X2_1562 ( .A(round_ctr_inc), .B(b_reg_0_), .Y(_abc_15497_new_n3730_));
AND2X2 AND2X2_1563 ( .A(_abc_15497_new_n2010_), .B(c_reg_31_), .Y(_abc_15497_new_n3733_));
AND2X2 AND2X2_1564 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n1006_), .Y(_abc_15497_new_n3734_));
AND2X2 AND2X2_1565 ( .A(round_ctr_inc), .B(b_reg_1_), .Y(_abc_15497_new_n3735_));
AND2X2 AND2X2_1566 ( .A(round_ctr_reg_5_), .B(round_ctr_reg_4_), .Y(_abc_15497_new_n3738_));
AND2X2 AND2X2_1567 ( .A(round_ctr_reg_5_), .B(round_ctr_reg_3_), .Y(_abc_15497_new_n3741_));
AND2X2 AND2X2_1568 ( .A(_abc_15497_new_n3742_), .B(_abc_15497_new_n3740_), .Y(_abc_15497_new_n3743_));
AND2X2 AND2X2_1569 ( .A(_abc_15497_new_n3743_), .B(_abc_15497_new_n3739_), .Y(_abc_15497_new_n3744_));
AND2X2 AND2X2_157 ( .A(_abc_15497_new_n1031_), .B(_abc_15497_new_n1029_), .Y(_abc_15497_new_n1032_));
AND2X2 AND2X2_1570 ( .A(_abc_15497_new_n3745_), .B(_abc_15497_new_n3746_), .Y(_abc_15497_new_n3747_));
AND2X2 AND2X2_1571 ( .A(_abc_15497_new_n3745_), .B(_abc_15497_new_n3749_), .Y(_abc_15497_new_n3750_));
AND2X2 AND2X2_1572 ( .A(_abc_15497_new_n3750_), .B(_abc_15497_new_n3748_), .Y(_abc_15497_new_n3751_));
AND2X2 AND2X2_1573 ( .A(_abc_15497_new_n3752_), .B(_abc_15497_new_n3740_), .Y(_abc_15497_new_n3753_));
AND2X2 AND2X2_1574 ( .A(_abc_15497_new_n3754_), .B(b_reg_0_), .Y(_abc_15497_new_n3755_));
AND2X2 AND2X2_1575 ( .A(b_reg_0_), .B(c_reg_0_), .Y(_abc_15497_new_n3757_));
AND2X2 AND2X2_1576 ( .A(_abc_15497_new_n3758_), .B(_abc_15497_new_n3756_), .Y(_abc_15497_new_n3759_));
AND2X2 AND2X2_1577 ( .A(_abc_15497_new_n3753_), .B(_abc_15497_new_n3760_), .Y(_abc_15497_new_n3761_));
AND2X2 AND2X2_1578 ( .A(_abc_15497_new_n3758_), .B(_abc_15497_new_n3762_), .Y(_abc_15497_new_n3763_));
AND2X2 AND2X2_1579 ( .A(_abc_15497_new_n3764_), .B(_abc_15497_new_n3756_), .Y(_abc_15497_new_n3765_));
AND2X2 AND2X2_158 ( .A(_abc_15497_new_n1022_), .B(_abc_15497_new_n1009_), .Y(_abc_15497_new_n1035_));
AND2X2 AND2X2_1580 ( .A(_abc_15497_new_n3763_), .B(d_reg_0_), .Y(_abc_15497_new_n3766_));
AND2X2 AND2X2_1581 ( .A(round_ctr_reg_3_), .B(round_ctr_reg_2_), .Y(_abc_15497_new_n3770_));
AND2X2 AND2X2_1582 ( .A(_abc_15497_new_n3738_), .B(_abc_15497_new_n3770_), .Y(_abc_15497_new_n3771_));
AND2X2 AND2X2_1583 ( .A(_abc_15497_new_n3772_), .B(_abc_15497_new_n3740_), .Y(_abc_15497_new_n3773_));
AND2X2 AND2X2_1584 ( .A(_abc_15497_new_n3773_), .B(_abc_15497_new_n3769_), .Y(_abc_15497_new_n3774_));
AND2X2 AND2X2_1585 ( .A(_abc_15497_new_n3777_), .B(round_ctr_reg_4_), .Y(_abc_15497_new_n3778_));
AND2X2 AND2X2_1586 ( .A(_abc_15497_new_n3785_), .B(_abc_15497_new_n3780_), .Y(_abc_15497_new_n3786_));
AND2X2 AND2X2_1587 ( .A(_abc_15497_new_n3776_), .B(_abc_15497_new_n3786_), .Y(_abc_15497_new_n3787_));
AND2X2 AND2X2_1588 ( .A(e_reg_0_), .B(a_reg_27_), .Y(_abc_15497_new_n3790_));
AND2X2 AND2X2_1589 ( .A(_abc_15497_new_n3791_), .B(_abc_15497_new_n3789_), .Y(_abc_15497_new_n3792_));
AND2X2 AND2X2_159 ( .A(_abc_15497_new_n1037_), .B(digest_update), .Y(_abc_15497_new_n1038_));
AND2X2 AND2X2_1590 ( .A(_abc_15497_new_n3792_), .B(w_0_), .Y(_abc_15497_new_n3793_));
AND2X2 AND2X2_1591 ( .A(_abc_15497_new_n3795_), .B(_abc_15497_new_n3794_), .Y(_abc_15497_new_n3796_));
AND2X2 AND2X2_1592 ( .A(_abc_15497_new_n3788_), .B(_abc_15497_new_n3797_), .Y(_abc_15497_new_n3798_));
AND2X2 AND2X2_1593 ( .A(_abc_15497_new_n3800_), .B(_abc_15497_new_n3801_), .Y(_abc_15497_new_n3802_));
AND2X2 AND2X2_1594 ( .A(_abc_15497_new_n3784_), .B(_abc_15497_new_n3780_), .Y(_abc_15497_new_n3803_));
AND2X2 AND2X2_1595 ( .A(_abc_15497_new_n3802_), .B(_abc_15497_new_n3803_), .Y(_abc_15497_new_n3804_));
AND2X2 AND2X2_1596 ( .A(_abc_15497_new_n3774_), .B(_abc_15497_new_n3805_), .Y(_abc_15497_new_n3806_));
AND2X2 AND2X2_1597 ( .A(_abc_15497_new_n3808_), .B(_abc_15497_new_n3799_), .Y(_abc_15497_new_n3809_));
AND2X2 AND2X2_1598 ( .A(_abc_15497_new_n3809_), .B(_abc_15497_new_n3810_), .Y(_abc_15497_new_n3811_));
AND2X2 AND2X2_1599 ( .A(_abc_15497_new_n3813_), .B(_abc_15497_new_n3744_), .Y(_abc_15497_new_n3815_));
AND2X2 AND2X2_16 ( .A(_abc_15497_new_n718_), .B(_abc_15497_new_n728_), .Y(_abc_15497_new_n729_));
AND2X2 AND2X2_160 ( .A(_abc_15497_new_n1038_), .B(_abc_15497_new_n1034_), .Y(_abc_15497_new_n1039_));
AND2X2 AND2X2_1600 ( .A(_abc_15497_new_n3816_), .B(round_ctr_inc), .Y(_abc_15497_new_n3817_));
AND2X2 AND2X2_1601 ( .A(_abc_15497_new_n3817_), .B(_abc_15497_new_n3814_), .Y(_abc_15497_new_n3818_));
AND2X2 AND2X2_1602 ( .A(_abc_15497_new_n2010_), .B(a_reg_0_), .Y(_abc_15497_new_n3819_));
AND2X2 AND2X2_1603 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n2715_), .Y(_abc_15497_new_n3820_));
AND2X2 AND2X2_1604 ( .A(b_reg_1_), .B(c_reg_1_), .Y(_abc_15497_new_n3825_));
AND2X2 AND2X2_1605 ( .A(_abc_15497_new_n3826_), .B(_abc_15497_new_n3824_), .Y(_abc_15497_new_n3827_));
AND2X2 AND2X2_1606 ( .A(_abc_15497_new_n3827_), .B(d_reg_1_), .Y(_abc_15497_new_n3830_));
AND2X2 AND2X2_1607 ( .A(_abc_15497_new_n3834_), .B(_abc_15497_new_n3826_), .Y(_abc_15497_new_n3835_));
AND2X2 AND2X2_1608 ( .A(_abc_15497_new_n3826_), .B(_abc_15497_new_n3833_), .Y(_abc_15497_new_n3838_));
AND2X2 AND2X2_1609 ( .A(_abc_15497_new_n3840_), .B(_abc_15497_new_n3836_), .Y(_abc_15497_new_n3841_));
AND2X2 AND2X2_161 ( .A(_abc_15497_new_n701_), .B(\digest[2] ), .Y(_abc_15497_new_n1040_));
AND2X2 AND2X2_1610 ( .A(_abc_15497_new_n3832_), .B(_abc_15497_new_n3841_), .Y(_abc_15497_new_n3842_));
AND2X2 AND2X2_1611 ( .A(e_reg_1_), .B(a_reg_28_), .Y(_abc_15497_new_n3845_));
AND2X2 AND2X2_1612 ( .A(_abc_15497_new_n3846_), .B(_abc_15497_new_n3844_), .Y(_abc_15497_new_n3847_));
AND2X2 AND2X2_1613 ( .A(_abc_15497_new_n3847_), .B(w_1_), .Y(_abc_15497_new_n3849_));
AND2X2 AND2X2_1614 ( .A(_abc_15497_new_n3850_), .B(_abc_15497_new_n3848_), .Y(_abc_15497_new_n3851_));
AND2X2 AND2X2_1615 ( .A(_abc_15497_new_n3851_), .B(_abc_15497_new_n3843_), .Y(_abc_15497_new_n3852_));
AND2X2 AND2X2_1616 ( .A(_abc_15497_new_n3853_), .B(_abc_15497_new_n3854_), .Y(_abc_15497_new_n3855_));
AND2X2 AND2X2_1617 ( .A(_abc_15497_new_n3857_), .B(_abc_15497_new_n3828_), .Y(_abc_15497_new_n3858_));
AND2X2 AND2X2_1618 ( .A(_abc_15497_new_n3803_), .B(_abc_15497_new_n3858_), .Y(_abc_15497_new_n3859_));
AND2X2 AND2X2_1619 ( .A(_abc_15497_new_n3753_), .B(_abc_15497_new_n3860_), .Y(_abc_15497_new_n3861_));
AND2X2 AND2X2_162 ( .A(_abc_15497_new_n701_), .B(\digest[3] ), .Y(_abc_15497_new_n1042_));
AND2X2 AND2X2_1620 ( .A(_abc_15497_new_n3774_), .B(_abc_15497_new_n3862_), .Y(_abc_15497_new_n3863_));
AND2X2 AND2X2_1621 ( .A(_abc_15497_new_n3868_), .B(_abc_15497_new_n3866_), .Y(_abc_15497_new_n3869_));
AND2X2 AND2X2_1622 ( .A(_abc_15497_new_n3856_), .B(_abc_15497_new_n3871_), .Y(_abc_15497_new_n3872_));
AND2X2 AND2X2_1623 ( .A(_abc_15497_new_n3874_), .B(_abc_15497_new_n3875_), .Y(_abc_15497_new_n3876_));
AND2X2 AND2X2_1624 ( .A(_abc_15497_new_n3873_), .B(_abc_15497_new_n3877_), .Y(_abc_15497_new_n3878_));
AND2X2 AND2X2_1625 ( .A(_abc_15497_new_n3878_), .B(_abc_15497_new_n3783_), .Y(_abc_15497_new_n3879_));
AND2X2 AND2X2_1626 ( .A(_abc_15497_new_n3876_), .B(_abc_15497_new_n3811_), .Y(_abc_15497_new_n3880_));
AND2X2 AND2X2_1627 ( .A(_abc_15497_new_n3823_), .B(_abc_15497_new_n3872_), .Y(_abc_15497_new_n3881_));
AND2X2 AND2X2_1628 ( .A(_abc_15497_new_n3882_), .B(_abc_15497_new_n3773_), .Y(_abc_15497_new_n3883_));
AND2X2 AND2X2_1629 ( .A(_abc_15497_new_n3887_), .B(round_ctr_inc), .Y(_abc_15497_new_n3888_));
AND2X2 AND2X2_163 ( .A(_abc_15497_new_n1036_), .B(_abc_15497_new_n1032_), .Y(_abc_15497_new_n1043_));
AND2X2 AND2X2_1630 ( .A(_abc_15497_new_n3888_), .B(_abc_15497_new_n3886_), .Y(_abc_15497_new_n3889_));
AND2X2 AND2X2_1631 ( .A(_abc_15497_new_n2010_), .B(a_reg_1_), .Y(_abc_15497_new_n3890_));
AND2X2 AND2X2_1632 ( .A(_abc_15497_new_n700_), .B(\digest[129] ), .Y(_abc_15497_new_n3891_));
AND2X2 AND2X2_1633 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3891_), .Y(_abc_15497_new_n3892_));
AND2X2 AND2X2_1634 ( .A(_abc_15497_new_n3896_), .B(_abc_15497_new_n3873_), .Y(_abc_15497_new_n3897_));
AND2X2 AND2X2_1635 ( .A(_abc_15497_new_n3865_), .B(_abc_15497_new_n3855_), .Y(_abc_15497_new_n3898_));
AND2X2 AND2X2_1636 ( .A(b_reg_2_), .B(c_reg_2_), .Y(_abc_15497_new_n3901_));
AND2X2 AND2X2_1637 ( .A(_abc_15497_new_n3902_), .B(_abc_15497_new_n3900_), .Y(_abc_15497_new_n3903_));
AND2X2 AND2X2_1638 ( .A(_abc_15497_new_n3903_), .B(d_reg_2_), .Y(_abc_15497_new_n3905_));
AND2X2 AND2X2_1639 ( .A(_abc_15497_new_n3906_), .B(_abc_15497_new_n3904_), .Y(_abc_15497_new_n3907_));
AND2X2 AND2X2_164 ( .A(e_reg_3_), .B(\digest[3] ), .Y(_abc_15497_new_n1046_));
AND2X2 AND2X2_1640 ( .A(_abc_15497_new_n3911_), .B(_abc_15497_new_n3902_), .Y(_abc_15497_new_n3912_));
AND2X2 AND2X2_1641 ( .A(_abc_15497_new_n3902_), .B(_abc_15497_new_n3910_), .Y(_abc_15497_new_n3915_));
AND2X2 AND2X2_1642 ( .A(_abc_15497_new_n3917_), .B(_abc_15497_new_n3913_), .Y(_abc_15497_new_n3918_));
AND2X2 AND2X2_1643 ( .A(_abc_15497_new_n3909_), .B(_abc_15497_new_n3918_), .Y(_abc_15497_new_n3919_));
AND2X2 AND2X2_1644 ( .A(e_reg_2_), .B(a_reg_29_), .Y(_abc_15497_new_n3922_));
AND2X2 AND2X2_1645 ( .A(_abc_15497_new_n3923_), .B(_abc_15497_new_n3921_), .Y(_abc_15497_new_n3924_));
AND2X2 AND2X2_1646 ( .A(_abc_15497_new_n3924_), .B(w_2_), .Y(_abc_15497_new_n3926_));
AND2X2 AND2X2_1647 ( .A(_abc_15497_new_n3927_), .B(_abc_15497_new_n3925_), .Y(_abc_15497_new_n3928_));
AND2X2 AND2X2_1648 ( .A(_abc_15497_new_n3928_), .B(_abc_15497_new_n3920_), .Y(_abc_15497_new_n3929_));
AND2X2 AND2X2_1649 ( .A(_abc_15497_new_n3932_), .B(_abc_15497_new_n3930_), .Y(_abc_15497_new_n3933_));
AND2X2 AND2X2_165 ( .A(_abc_15497_new_n1047_), .B(_abc_15497_new_n1045_), .Y(_abc_15497_new_n1048_));
AND2X2 AND2X2_1650 ( .A(_abc_15497_new_n3803_), .B(_abc_15497_new_n3907_), .Y(_abc_15497_new_n3936_));
AND2X2 AND2X2_1651 ( .A(_abc_15497_new_n3753_), .B(_abc_15497_new_n3937_), .Y(_abc_15497_new_n3938_));
AND2X2 AND2X2_1652 ( .A(_abc_15497_new_n3774_), .B(_abc_15497_new_n3939_), .Y(_abc_15497_new_n3940_));
AND2X2 AND2X2_1653 ( .A(_abc_15497_new_n3943_), .B(_abc_15497_new_n3944_), .Y(_abc_15497_new_n3945_));
AND2X2 AND2X2_1654 ( .A(_abc_15497_new_n3935_), .B(_abc_15497_new_n3946_), .Y(_abc_15497_new_n3947_));
AND2X2 AND2X2_1655 ( .A(_abc_15497_new_n3947_), .B(_abc_15497_new_n3899_), .Y(_abc_15497_new_n3948_));
AND2X2 AND2X2_1656 ( .A(_abc_15497_new_n3874_), .B(_abc_15497_new_n3853_), .Y(_abc_15497_new_n3949_));
AND2X2 AND2X2_1657 ( .A(_abc_15497_new_n3950_), .B(_abc_15497_new_n3951_), .Y(_abc_15497_new_n3952_));
AND2X2 AND2X2_1658 ( .A(_abc_15497_new_n3952_), .B(_abc_15497_new_n3949_), .Y(_abc_15497_new_n3953_));
AND2X2 AND2X2_1659 ( .A(_abc_15497_new_n3954_), .B(_abc_15497_new_n3744_), .Y(_abc_15497_new_n3955_));
AND2X2 AND2X2_166 ( .A(_abc_15497_new_n1034_), .B(_abc_15497_new_n1031_), .Y(_abc_15497_new_n1050_));
AND2X2 AND2X2_1660 ( .A(_abc_15497_new_n3956_), .B(_abc_15497_new_n3957_), .Y(_abc_15497_new_n3958_));
AND2X2 AND2X2_1661 ( .A(_abc_15497_new_n3958_), .B(_abc_15497_new_n3769_), .Y(_abc_15497_new_n3959_));
AND2X2 AND2X2_1662 ( .A(_abc_15497_new_n3963_), .B(_abc_15497_new_n3964_), .Y(_abc_15497_new_n3965_));
AND2X2 AND2X2_1663 ( .A(_abc_15497_new_n3961_), .B(_abc_15497_new_n3966_), .Y(_abc_15497_new_n3967_));
AND2X2 AND2X2_1664 ( .A(_abc_15497_new_n3965_), .B(_abc_15497_new_n3962_), .Y(_abc_15497_new_n3969_));
AND2X2 AND2X2_1665 ( .A(_abc_15497_new_n3960_), .B(_abc_15497_new_n3897_), .Y(_abc_15497_new_n3970_));
AND2X2 AND2X2_1666 ( .A(_abc_15497_new_n3972_), .B(round_ctr_inc), .Y(_abc_15497_new_n3973_));
AND2X2 AND2X2_1667 ( .A(_abc_15497_new_n3973_), .B(_abc_15497_new_n3968_), .Y(_abc_15497_new_n3974_));
AND2X2 AND2X2_1668 ( .A(_abc_15497_new_n2010_), .B(a_reg_2_), .Y(_abc_15497_new_n3975_));
AND2X2 AND2X2_1669 ( .A(_abc_15497_new_n700_), .B(\digest[130] ), .Y(_abc_15497_new_n3976_));
AND2X2 AND2X2_167 ( .A(_abc_15497_new_n1052_), .B(_abc_15497_new_n1049_), .Y(_abc_15497_new_n1053_));
AND2X2 AND2X2_1670 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3976_), .Y(_abc_15497_new_n3977_));
AND2X2 AND2X2_1671 ( .A(_abc_15497_new_n3972_), .B(_abc_15497_new_n3961_), .Y(_abc_15497_new_n3980_));
AND2X2 AND2X2_1672 ( .A(_abc_15497_new_n3964_), .B(_abc_15497_new_n3956_), .Y(_abc_15497_new_n3981_));
AND2X2 AND2X2_1673 ( .A(_abc_15497_new_n3935_), .B(_abc_15497_new_n3943_), .Y(_abc_15497_new_n3983_));
AND2X2 AND2X2_1674 ( .A(b_reg_3_), .B(c_reg_3_), .Y(_abc_15497_new_n3986_));
AND2X2 AND2X2_1675 ( .A(_abc_15497_new_n3987_), .B(_abc_15497_new_n3985_), .Y(_abc_15497_new_n3988_));
AND2X2 AND2X2_1676 ( .A(_abc_15497_new_n3989_), .B(_abc_15497_new_n3984_), .Y(_abc_15497_new_n3990_));
AND2X2 AND2X2_1677 ( .A(_abc_15497_new_n3988_), .B(d_reg_3_), .Y(_abc_15497_new_n3991_));
AND2X2 AND2X2_1678 ( .A(_abc_15497_new_n3994_), .B(_abc_15497_new_n3987_), .Y(_abc_15497_new_n3995_));
AND2X2 AND2X2_1679 ( .A(_abc_15497_new_n3987_), .B(_abc_15497_new_n3984_), .Y(_abc_15497_new_n3998_));
AND2X2 AND2X2_168 ( .A(_abc_15497_new_n1053_), .B(digest_update), .Y(_abc_15497_new_n1054_));
AND2X2 AND2X2_1680 ( .A(_abc_15497_new_n4000_), .B(_abc_15497_new_n3996_), .Y(_abc_15497_new_n4001_));
AND2X2 AND2X2_1681 ( .A(_abc_15497_new_n3993_), .B(_abc_15497_new_n4001_), .Y(_abc_15497_new_n4002_));
AND2X2 AND2X2_1682 ( .A(_abc_15497_new_n3927_), .B(_abc_15497_new_n3923_), .Y(_abc_15497_new_n4003_));
AND2X2 AND2X2_1683 ( .A(e_reg_3_), .B(a_reg_30_), .Y(_abc_15497_new_n4007_));
AND2X2 AND2X2_1684 ( .A(_abc_15497_new_n4008_), .B(_abc_15497_new_n4006_), .Y(_abc_15497_new_n4009_));
AND2X2 AND2X2_1685 ( .A(_abc_15497_new_n4010_), .B(_abc_15497_new_n4005_), .Y(_abc_15497_new_n4011_));
AND2X2 AND2X2_1686 ( .A(_abc_15497_new_n4009_), .B(w_3_), .Y(_abc_15497_new_n4012_));
AND2X2 AND2X2_1687 ( .A(_abc_15497_new_n4014_), .B(_abc_15497_new_n4004_), .Y(_abc_15497_new_n4015_));
AND2X2 AND2X2_1688 ( .A(_abc_15497_new_n4013_), .B(_abc_15497_new_n4003_), .Y(_abc_15497_new_n4016_));
AND2X2 AND2X2_1689 ( .A(_abc_15497_new_n4017_), .B(_abc_15497_new_n4002_), .Y(_abc_15497_new_n4020_));
AND2X2 AND2X2_169 ( .A(e_reg_4_), .B(\digest[4] ), .Y(_abc_15497_new_n1057_));
AND2X2 AND2X2_1690 ( .A(_abc_15497_new_n4024_), .B(_abc_15497_new_n4018_), .Y(_abc_15497_new_n4025_));
AND2X2 AND2X2_1691 ( .A(_abc_15497_new_n4022_), .B(_abc_15497_new_n4026_), .Y(_abc_15497_new_n4027_));
AND2X2 AND2X2_1692 ( .A(_abc_15497_new_n4023_), .B(_abc_15497_new_n4025_), .Y(_abc_15497_new_n4029_));
AND2X2 AND2X2_1693 ( .A(_abc_15497_new_n4021_), .B(_abc_15497_new_n3983_), .Y(_abc_15497_new_n4030_));
AND2X2 AND2X2_1694 ( .A(_abc_15497_new_n4032_), .B(_abc_15497_new_n4028_), .Y(_abc_15497_new_n4033_));
AND2X2 AND2X2_1695 ( .A(_abc_15497_new_n4033_), .B(_abc_15497_new_n3982_), .Y(_abc_15497_new_n4034_));
AND2X2 AND2X2_1696 ( .A(_abc_15497_new_n4031_), .B(_abc_15497_new_n3803_), .Y(_abc_15497_new_n4035_));
AND2X2 AND2X2_1697 ( .A(_abc_15497_new_n4027_), .B(_abc_15497_new_n3775_), .Y(_abc_15497_new_n4036_));
AND2X2 AND2X2_1698 ( .A(_abc_15497_new_n4037_), .B(_abc_15497_new_n3981_), .Y(_abc_15497_new_n4038_));
AND2X2 AND2X2_1699 ( .A(_abc_15497_new_n4042_), .B(_abc_15497_new_n4043_), .Y(_abc_15497_new_n4044_));
AND2X2 AND2X2_17 ( .A(_abc_15497_new_n711_), .B(_abc_15497_new_n729_), .Y(_abc_15497_new_n730_));
AND2X2 AND2X2_170 ( .A(_abc_15497_new_n1058_), .B(_abc_15497_new_n1056_), .Y(_abc_15497_new_n1059_));
AND2X2 AND2X2_1700 ( .A(_abc_15497_new_n4045_), .B(round_ctr_inc), .Y(_abc_15497_new_n4046_));
AND2X2 AND2X2_1701 ( .A(_abc_15497_new_n4046_), .B(_abc_15497_new_n4040_), .Y(_abc_15497_new_n4047_));
AND2X2 AND2X2_1702 ( .A(_abc_15497_new_n2010_), .B(a_reg_3_), .Y(_abc_15497_new_n4048_));
AND2X2 AND2X2_1703 ( .A(_abc_15497_new_n700_), .B(\digest[131] ), .Y(_abc_15497_new_n4049_));
AND2X2 AND2X2_1704 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n4049_), .Y(_abc_15497_new_n4050_));
AND2X2 AND2X2_1705 ( .A(_abc_15497_new_n3967_), .B(_abc_15497_new_n3895_), .Y(_abc_15497_new_n4053_));
AND2X2 AND2X2_1706 ( .A(_abc_15497_new_n4053_), .B(_abc_15497_new_n4044_), .Y(_abc_15497_new_n4054_));
AND2X2 AND2X2_1707 ( .A(_abc_15497_new_n4043_), .B(_abc_15497_new_n3969_), .Y(_abc_15497_new_n4055_));
AND2X2 AND2X2_1708 ( .A(_abc_15497_new_n4032_), .B(_abc_15497_new_n4022_), .Y(_abc_15497_new_n4058_));
AND2X2 AND2X2_1709 ( .A(_abc_15497_new_n3744_), .B(_abc_15497_new_n3779_), .Y(_abc_15497_new_n4059_));
AND2X2 AND2X2_171 ( .A(_abc_15497_new_n1062_), .B(_abc_15497_new_n1047_), .Y(_abc_15497_new_n1063_));
AND2X2 AND2X2_1710 ( .A(_abc_15497_new_n4018_), .B(_abc_15497_new_n4061_), .Y(_abc_15497_new_n4062_));
AND2X2 AND2X2_1711 ( .A(b_reg_4_), .B(c_reg_4_), .Y(_abc_15497_new_n4065_));
AND2X2 AND2X2_1712 ( .A(_abc_15497_new_n4066_), .B(_abc_15497_new_n4064_), .Y(_abc_15497_new_n4067_));
AND2X2 AND2X2_1713 ( .A(_abc_15497_new_n4068_), .B(_abc_15497_new_n4063_), .Y(_abc_15497_new_n4069_));
AND2X2 AND2X2_1714 ( .A(_abc_15497_new_n4067_), .B(d_reg_4_), .Y(_abc_15497_new_n4070_));
AND2X2 AND2X2_1715 ( .A(_abc_15497_new_n4072_), .B(_abc_15497_new_n3803_), .Y(_abc_15497_new_n4073_));
AND2X2 AND2X2_1716 ( .A(_abc_15497_new_n4074_), .B(d_reg_4_), .Y(_abc_15497_new_n4075_));
AND2X2 AND2X2_1717 ( .A(_abc_15497_new_n3753_), .B(_abc_15497_new_n4076_), .Y(_abc_15497_new_n4077_));
AND2X2 AND2X2_1718 ( .A(_abc_15497_new_n4066_), .B(_abc_15497_new_n4063_), .Y(_abc_15497_new_n4079_));
AND2X2 AND2X2_1719 ( .A(_abc_15497_new_n3774_), .B(_abc_15497_new_n4081_), .Y(_abc_15497_new_n4082_));
AND2X2 AND2X2_172 ( .A(_abc_15497_new_n1044_), .B(_abc_15497_new_n1045_), .Y(_abc_15497_new_n1065_));
AND2X2 AND2X2_1720 ( .A(e_reg_4_), .B(a_reg_31_), .Y(_abc_15497_new_n4088_));
AND2X2 AND2X2_1721 ( .A(_abc_15497_new_n4089_), .B(_abc_15497_new_n4087_), .Y(_abc_15497_new_n4090_));
AND2X2 AND2X2_1722 ( .A(_abc_15497_new_n4091_), .B(_abc_15497_new_n4086_), .Y(_abc_15497_new_n4092_));
AND2X2 AND2X2_1723 ( .A(_abc_15497_new_n4090_), .B(w_4_), .Y(_abc_15497_new_n4093_));
AND2X2 AND2X2_1724 ( .A(_abc_15497_new_n4095_), .B(_abc_15497_new_n4085_), .Y(_abc_15497_new_n4096_));
AND2X2 AND2X2_1725 ( .A(_abc_15497_new_n4097_), .B(_abc_15497_new_n4094_), .Y(_abc_15497_new_n4098_));
AND2X2 AND2X2_1726 ( .A(_abc_15497_new_n4100_), .B(_abc_15497_new_n4084_), .Y(_abc_15497_new_n4101_));
AND2X2 AND2X2_1727 ( .A(_abc_15497_new_n4102_), .B(_abc_15497_new_n4099_), .Y(_abc_15497_new_n4103_));
AND2X2 AND2X2_1728 ( .A(_abc_15497_new_n4107_), .B(_abc_15497_new_n4108_), .Y(_abc_15497_new_n4109_));
AND2X2 AND2X2_1729 ( .A(_abc_15497_new_n4110_), .B(_abc_15497_new_n4105_), .Y(_abc_15497_new_n4111_));
AND2X2 AND2X2_173 ( .A(_abc_15497_new_n1064_), .B(_abc_15497_new_n1067_), .Y(_abc_15497_new_n1068_));
AND2X2 AND2X2_1730 ( .A(_abc_15497_new_n4111_), .B(_abc_15497_new_n4060_), .Y(_abc_15497_new_n4112_));
AND2X2 AND2X2_1731 ( .A(_abc_15497_new_n4109_), .B(_abc_15497_new_n4106_), .Y(_abc_15497_new_n4113_));
AND2X2 AND2X2_1732 ( .A(_abc_15497_new_n4104_), .B(_abc_15497_new_n4062_), .Y(_abc_15497_new_n4114_));
AND2X2 AND2X2_1733 ( .A(_abc_15497_new_n4115_), .B(_abc_15497_new_n4059_), .Y(_abc_15497_new_n4116_));
AND2X2 AND2X2_1734 ( .A(_abc_15497_new_n4117_), .B(_abc_15497_new_n4058_), .Y(_abc_15497_new_n4118_));
AND2X2 AND2X2_1735 ( .A(_abc_15497_new_n4120_), .B(_abc_15497_new_n4121_), .Y(_abc_15497_new_n4122_));
AND2X2 AND2X2_1736 ( .A(_abc_15497_new_n4122_), .B(_abc_15497_new_n4119_), .Y(_abc_15497_new_n4123_));
AND2X2 AND2X2_1737 ( .A(_abc_15497_new_n4057_), .B(_abc_15497_new_n4125_), .Y(_abc_15497_new_n4127_));
AND2X2 AND2X2_1738 ( .A(_abc_15497_new_n4128_), .B(round_ctr_inc), .Y(_abc_15497_new_n4129_));
AND2X2 AND2X2_1739 ( .A(_abc_15497_new_n4129_), .B(_abc_15497_new_n4126_), .Y(_abc_15497_new_n4130_));
AND2X2 AND2X2_174 ( .A(_abc_15497_new_n1069_), .B(_abc_15497_new_n1071_), .Y(_0H4_reg_31_0__4_));
AND2X2 AND2X2_1740 ( .A(_abc_15497_new_n2010_), .B(a_reg_4_), .Y(_abc_15497_new_n4131_));
AND2X2 AND2X2_1741 ( .A(_abc_15497_new_n700_), .B(\digest[132] ), .Y(_abc_15497_new_n4132_));
AND2X2 AND2X2_1742 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n4132_), .Y(_abc_15497_new_n4133_));
AND2X2 AND2X2_1743 ( .A(_abc_15497_new_n4128_), .B(_abc_15497_new_n4136_), .Y(_abc_15497_new_n4137_));
AND2X2 AND2X2_1744 ( .A(b_reg_5_), .B(c_reg_5_), .Y(_abc_15497_new_n4143_));
AND2X2 AND2X2_1745 ( .A(_abc_15497_new_n4144_), .B(_abc_15497_new_n4142_), .Y(_abc_15497_new_n4145_));
AND2X2 AND2X2_1746 ( .A(_abc_15497_new_n4146_), .B(_abc_15497_new_n4141_), .Y(_abc_15497_new_n4147_));
AND2X2 AND2X2_1747 ( .A(_abc_15497_new_n4145_), .B(d_reg_5_), .Y(_abc_15497_new_n4148_));
AND2X2 AND2X2_1748 ( .A(_abc_15497_new_n4150_), .B(_abc_15497_new_n3803_), .Y(_abc_15497_new_n4151_));
AND2X2 AND2X2_1749 ( .A(_abc_15497_new_n4152_), .B(d_reg_5_), .Y(_abc_15497_new_n4153_));
AND2X2 AND2X2_175 ( .A(_abc_15497_new_n1066_), .B(_abc_15497_new_n1059_), .Y(_abc_15497_new_n1073_));
AND2X2 AND2X2_1750 ( .A(_abc_15497_new_n3753_), .B(_abc_15497_new_n4154_), .Y(_abc_15497_new_n4155_));
AND2X2 AND2X2_1751 ( .A(_abc_15497_new_n4144_), .B(_abc_15497_new_n4141_), .Y(_abc_15497_new_n4157_));
AND2X2 AND2X2_1752 ( .A(_abc_15497_new_n3774_), .B(_abc_15497_new_n4159_), .Y(_abc_15497_new_n4160_));
AND2X2 AND2X2_1753 ( .A(e_reg_5_), .B(a_reg_0_), .Y(_abc_15497_new_n4167_));
AND2X2 AND2X2_1754 ( .A(_abc_15497_new_n4168_), .B(_abc_15497_new_n4166_), .Y(_abc_15497_new_n4169_));
AND2X2 AND2X2_1755 ( .A(_abc_15497_new_n4170_), .B(_abc_15497_new_n4165_), .Y(_abc_15497_new_n4171_));
AND2X2 AND2X2_1756 ( .A(_abc_15497_new_n4169_), .B(w_5_), .Y(_abc_15497_new_n4172_));
AND2X2 AND2X2_1757 ( .A(_abc_15497_new_n4174_), .B(_abc_15497_new_n4164_), .Y(_abc_15497_new_n4175_));
AND2X2 AND2X2_1758 ( .A(_abc_15497_new_n4176_), .B(_abc_15497_new_n4173_), .Y(_abc_15497_new_n4177_));
AND2X2 AND2X2_1759 ( .A(_abc_15497_new_n4179_), .B(_abc_15497_new_n4181_), .Y(_abc_15497_new_n4182_));
AND2X2 AND2X2_176 ( .A(e_reg_5_), .B(\digest[5] ), .Y(_abc_15497_new_n1076_));
AND2X2 AND2X2_1760 ( .A(_abc_15497_new_n4107_), .B(_abc_15497_new_n4184_), .Y(_abc_15497_new_n4185_));
AND2X2 AND2X2_1761 ( .A(_abc_15497_new_n4180_), .B(_abc_15497_new_n4162_), .Y(_abc_15497_new_n4186_));
AND2X2 AND2X2_1762 ( .A(_abc_15497_new_n4163_), .B(_abc_15497_new_n4178_), .Y(_abc_15497_new_n4187_));
AND2X2 AND2X2_1763 ( .A(_abc_15497_new_n4189_), .B(_abc_15497_new_n4183_), .Y(_abc_15497_new_n4190_));
AND2X2 AND2X2_1764 ( .A(_abc_15497_new_n4188_), .B(_abc_15497_new_n4185_), .Y(_abc_15497_new_n4192_));
AND2X2 AND2X2_1765 ( .A(_abc_15497_new_n4182_), .B(_abc_15497_new_n4140_), .Y(_abc_15497_new_n4193_));
AND2X2 AND2X2_1766 ( .A(_abc_15497_new_n4191_), .B(_abc_15497_new_n4195_), .Y(_abc_15497_new_n4196_));
AND2X2 AND2X2_1767 ( .A(_abc_15497_new_n4196_), .B(_abc_15497_new_n4139_), .Y(_abc_15497_new_n4197_));
AND2X2 AND2X2_1768 ( .A(_abc_15497_new_n4120_), .B(_abc_15497_new_n4105_), .Y(_abc_15497_new_n4198_));
AND2X2 AND2X2_1769 ( .A(_abc_15497_new_n4194_), .B(_abc_15497_new_n4060_), .Y(_abc_15497_new_n4199_));
AND2X2 AND2X2_177 ( .A(_abc_15497_new_n1077_), .B(_abc_15497_new_n1075_), .Y(_abc_15497_new_n1078_));
AND2X2 AND2X2_1770 ( .A(_abc_15497_new_n4190_), .B(_abc_15497_new_n4059_), .Y(_abc_15497_new_n4200_));
AND2X2 AND2X2_1771 ( .A(_abc_15497_new_n4201_), .B(_abc_15497_new_n4198_), .Y(_abc_15497_new_n4202_));
AND2X2 AND2X2_1772 ( .A(_abc_15497_new_n4206_), .B(round_ctr_inc), .Y(_abc_15497_new_n4207_));
AND2X2 AND2X2_1773 ( .A(_abc_15497_new_n4207_), .B(_abc_15497_new_n4205_), .Y(_abc_15497_new_n4208_));
AND2X2 AND2X2_1774 ( .A(_abc_15497_new_n2010_), .B(a_reg_5_), .Y(_abc_15497_new_n4209_));
AND2X2 AND2X2_1775 ( .A(_abc_15497_new_n700_), .B(\digest[133] ), .Y(_abc_15497_new_n4210_));
AND2X2 AND2X2_1776 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n4210_), .Y(_abc_15497_new_n4211_));
AND2X2 AND2X2_1777 ( .A(_abc_15497_new_n4057_), .B(_abc_15497_new_n4215_), .Y(_abc_15497_new_n4216_));
AND2X2 AND2X2_1778 ( .A(_abc_15497_new_n4218_), .B(_abc_15497_new_n4217_), .Y(_abc_15497_new_n4219_));
AND2X2 AND2X2_1779 ( .A(b_reg_6_), .B(c_reg_6_), .Y(_abc_15497_new_n4226_));
AND2X2 AND2X2_178 ( .A(_abc_15497_new_n1064_), .B(_abc_15497_new_n1058_), .Y(_abc_15497_new_n1080_));
AND2X2 AND2X2_1780 ( .A(_abc_15497_new_n4227_), .B(_abc_15497_new_n4225_), .Y(_abc_15497_new_n4228_));
AND2X2 AND2X2_1781 ( .A(_abc_15497_new_n4229_), .B(_abc_15497_new_n4224_), .Y(_abc_15497_new_n4230_));
AND2X2 AND2X2_1782 ( .A(_abc_15497_new_n4228_), .B(d_reg_6_), .Y(_abc_15497_new_n4231_));
AND2X2 AND2X2_1783 ( .A(_abc_15497_new_n4233_), .B(_abc_15497_new_n3803_), .Y(_abc_15497_new_n4234_));
AND2X2 AND2X2_1784 ( .A(_abc_15497_new_n4235_), .B(d_reg_6_), .Y(_abc_15497_new_n4236_));
AND2X2 AND2X2_1785 ( .A(_abc_15497_new_n3753_), .B(_abc_15497_new_n4237_), .Y(_abc_15497_new_n4238_));
AND2X2 AND2X2_1786 ( .A(_abc_15497_new_n4227_), .B(_abc_15497_new_n4224_), .Y(_abc_15497_new_n4240_));
AND2X2 AND2X2_1787 ( .A(_abc_15497_new_n3774_), .B(_abc_15497_new_n4242_), .Y(_abc_15497_new_n4243_));
AND2X2 AND2X2_1788 ( .A(e_reg_6_), .B(a_reg_1_), .Y(_abc_15497_new_n4250_));
AND2X2 AND2X2_1789 ( .A(_abc_15497_new_n4251_), .B(_abc_15497_new_n4249_), .Y(_abc_15497_new_n4252_));
AND2X2 AND2X2_179 ( .A(_abc_15497_new_n1082_), .B(_abc_15497_new_n1079_), .Y(_abc_15497_new_n1083_));
AND2X2 AND2X2_1790 ( .A(_abc_15497_new_n4253_), .B(_abc_15497_new_n4248_), .Y(_abc_15497_new_n4254_));
AND2X2 AND2X2_1791 ( .A(_abc_15497_new_n4252_), .B(w_6_), .Y(_abc_15497_new_n4255_));
AND2X2 AND2X2_1792 ( .A(_abc_15497_new_n4257_), .B(_abc_15497_new_n4247_), .Y(_abc_15497_new_n4258_));
AND2X2 AND2X2_1793 ( .A(_abc_15497_new_n4259_), .B(_abc_15497_new_n4256_), .Y(_abc_15497_new_n4260_));
AND2X2 AND2X2_1794 ( .A(_abc_15497_new_n4262_), .B(_abc_15497_new_n4264_), .Y(_abc_15497_new_n4265_));
AND2X2 AND2X2_1795 ( .A(_abc_15497_new_n4179_), .B(_abc_15497_new_n4267_), .Y(_abc_15497_new_n4268_));
AND2X2 AND2X2_1796 ( .A(_abc_15497_new_n4263_), .B(_abc_15497_new_n4245_), .Y(_abc_15497_new_n4269_));
AND2X2 AND2X2_1797 ( .A(_abc_15497_new_n4246_), .B(_abc_15497_new_n4261_), .Y(_abc_15497_new_n4270_));
AND2X2 AND2X2_1798 ( .A(_abc_15497_new_n4272_), .B(_abc_15497_new_n4266_), .Y(_abc_15497_new_n4273_));
AND2X2 AND2X2_1799 ( .A(_abc_15497_new_n4271_), .B(_abc_15497_new_n4268_), .Y(_abc_15497_new_n4275_));
AND2X2 AND2X2_18 ( .A(c_reg_19_), .B(\digest[83] ), .Y(_abc_15497_new_n731_));
AND2X2 AND2X2_180 ( .A(_abc_15497_new_n1083_), .B(digest_update), .Y(_abc_15497_new_n1084_));
AND2X2 AND2X2_1800 ( .A(_abc_15497_new_n4265_), .B(_abc_15497_new_n4223_), .Y(_abc_15497_new_n4276_));
AND2X2 AND2X2_1801 ( .A(_abc_15497_new_n4274_), .B(_abc_15497_new_n4278_), .Y(_abc_15497_new_n4279_));
AND2X2 AND2X2_1802 ( .A(_abc_15497_new_n4279_), .B(_abc_15497_new_n4222_), .Y(_abc_15497_new_n4280_));
AND2X2 AND2X2_1803 ( .A(_abc_15497_new_n4195_), .B(_abc_15497_new_n4189_), .Y(_abc_15497_new_n4281_));
AND2X2 AND2X2_1804 ( .A(_abc_15497_new_n4277_), .B(_abc_15497_new_n3744_), .Y(_abc_15497_new_n4282_));
AND2X2 AND2X2_1805 ( .A(_abc_15497_new_n4273_), .B(_abc_15497_new_n3769_), .Y(_abc_15497_new_n4283_));
AND2X2 AND2X2_1806 ( .A(_abc_15497_new_n4284_), .B(_abc_15497_new_n4281_), .Y(_abc_15497_new_n4285_));
AND2X2 AND2X2_1807 ( .A(_abc_15497_new_n4221_), .B(_abc_15497_new_n4287_), .Y(_abc_15497_new_n4289_));
AND2X2 AND2X2_1808 ( .A(_abc_15497_new_n4290_), .B(round_ctr_inc), .Y(_abc_15497_new_n4291_));
AND2X2 AND2X2_1809 ( .A(_abc_15497_new_n4291_), .B(_abc_15497_new_n4288_), .Y(_abc_15497_new_n4292_));
AND2X2 AND2X2_181 ( .A(_abc_15497_new_n1085_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n1086_));
AND2X2 AND2X2_1810 ( .A(_abc_15497_new_n2010_), .B(a_reg_6_), .Y(_abc_15497_new_n4293_));
AND2X2 AND2X2_1811 ( .A(_abc_15497_new_n700_), .B(\digest[134] ), .Y(_abc_15497_new_n4294_));
AND2X2 AND2X2_1812 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n4294_), .Y(_abc_15497_new_n4295_));
AND2X2 AND2X2_1813 ( .A(_abc_15497_new_n4290_), .B(_abc_15497_new_n4298_), .Y(_abc_15497_new_n4299_));
AND2X2 AND2X2_1814 ( .A(_abc_15497_new_n4262_), .B(_abc_15497_new_n4301_), .Y(_abc_15497_new_n4302_));
AND2X2 AND2X2_1815 ( .A(b_reg_7_), .B(c_reg_7_), .Y(_abc_15497_new_n4306_));
AND2X2 AND2X2_1816 ( .A(_abc_15497_new_n4307_), .B(_abc_15497_new_n4305_), .Y(_abc_15497_new_n4308_));
AND2X2 AND2X2_1817 ( .A(_abc_15497_new_n4309_), .B(_abc_15497_new_n4304_), .Y(_abc_15497_new_n4310_));
AND2X2 AND2X2_1818 ( .A(_abc_15497_new_n4308_), .B(d_reg_7_), .Y(_abc_15497_new_n4311_));
AND2X2 AND2X2_1819 ( .A(_abc_15497_new_n4314_), .B(d_reg_7_), .Y(_abc_15497_new_n4315_));
AND2X2 AND2X2_182 ( .A(_abc_15497_new_n1074_), .B(_abc_15497_new_n1078_), .Y(_abc_15497_new_n1088_));
AND2X2 AND2X2_1820 ( .A(_abc_15497_new_n3753_), .B(_abc_15497_new_n4316_), .Y(_abc_15497_new_n4317_));
AND2X2 AND2X2_1821 ( .A(_abc_15497_new_n4307_), .B(_abc_15497_new_n4304_), .Y(_abc_15497_new_n4320_));
AND2X2 AND2X2_1822 ( .A(_abc_15497_new_n4318_), .B(_abc_15497_new_n4322_), .Y(_abc_15497_new_n4323_));
AND2X2 AND2X2_1823 ( .A(_abc_15497_new_n4323_), .B(_abc_15497_new_n4313_), .Y(_abc_15497_new_n4324_));
AND2X2 AND2X2_1824 ( .A(e_reg_7_), .B(a_reg_2_), .Y(_abc_15497_new_n4329_));
AND2X2 AND2X2_1825 ( .A(_abc_15497_new_n4330_), .B(_abc_15497_new_n4328_), .Y(_abc_15497_new_n4331_));
AND2X2 AND2X2_1826 ( .A(_abc_15497_new_n4332_), .B(_abc_15497_new_n4327_), .Y(_abc_15497_new_n4333_));
AND2X2 AND2X2_1827 ( .A(_abc_15497_new_n4331_), .B(w_7_), .Y(_abc_15497_new_n4334_));
AND2X2 AND2X2_1828 ( .A(_abc_15497_new_n4336_), .B(_abc_15497_new_n4326_), .Y(_abc_15497_new_n4337_));
AND2X2 AND2X2_1829 ( .A(_abc_15497_new_n4338_), .B(_abc_15497_new_n4339_), .Y(_abc_15497_new_n4340_));
AND2X2 AND2X2_183 ( .A(e_reg_6_), .B(\digest[6] ), .Y(_abc_15497_new_n1091_));
AND2X2 AND2X2_1830 ( .A(_abc_15497_new_n4325_), .B(_abc_15497_new_n4340_), .Y(_abc_15497_new_n4341_));
AND2X2 AND2X2_1831 ( .A(_abc_15497_new_n4343_), .B(_abc_15497_new_n4324_), .Y(_abc_15497_new_n4344_));
AND2X2 AND2X2_1832 ( .A(_abc_15497_new_n4346_), .B(_abc_15497_new_n4303_), .Y(_abc_15497_new_n4347_));
AND2X2 AND2X2_1833 ( .A(_abc_15497_new_n4345_), .B(_abc_15497_new_n4302_), .Y(_abc_15497_new_n4348_));
AND2X2 AND2X2_1834 ( .A(_abc_15497_new_n4300_), .B(_abc_15497_new_n4349_), .Y(_abc_15497_new_n4350_));
AND2X2 AND2X2_1835 ( .A(_abc_15497_new_n4278_), .B(_abc_15497_new_n4272_), .Y(_abc_15497_new_n4351_));
AND2X2 AND2X2_1836 ( .A(_abc_15497_new_n4351_), .B(_abc_15497_new_n4352_), .Y(_abc_15497_new_n4353_));
AND2X2 AND2X2_1837 ( .A(_abc_15497_new_n4358_), .B(round_ctr_inc), .Y(_abc_15497_new_n4359_));
AND2X2 AND2X2_1838 ( .A(_abc_15497_new_n4359_), .B(_abc_15497_new_n4355_), .Y(_abc_15497_new_n4360_));
AND2X2 AND2X2_1839 ( .A(_abc_15497_new_n2010_), .B(a_reg_7_), .Y(_abc_15497_new_n4361_));
AND2X2 AND2X2_184 ( .A(_abc_15497_new_n1092_), .B(_abc_15497_new_n1090_), .Y(_abc_15497_new_n1093_));
AND2X2 AND2X2_1840 ( .A(_abc_15497_new_n700_), .B(\digest[135] ), .Y(_abc_15497_new_n4362_));
AND2X2 AND2X2_1841 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n4362_), .Y(_abc_15497_new_n4363_));
AND2X2 AND2X2_1842 ( .A(b_reg_8_), .B(c_reg_8_), .Y(_abc_15497_new_n4370_));
AND2X2 AND2X2_1843 ( .A(_abc_15497_new_n4371_), .B(_abc_15497_new_n4369_), .Y(_abc_15497_new_n4372_));
AND2X2 AND2X2_1844 ( .A(_abc_15497_new_n4373_), .B(_abc_15497_new_n4368_), .Y(_abc_15497_new_n4374_));
AND2X2 AND2X2_1845 ( .A(_abc_15497_new_n4372_), .B(d_reg_8_), .Y(_abc_15497_new_n4375_));
AND2X2 AND2X2_1846 ( .A(_abc_15497_new_n4378_), .B(d_reg_8_), .Y(_abc_15497_new_n4379_));
AND2X2 AND2X2_1847 ( .A(_abc_15497_new_n3753_), .B(_abc_15497_new_n4380_), .Y(_abc_15497_new_n4381_));
AND2X2 AND2X2_1848 ( .A(_abc_15497_new_n4371_), .B(_abc_15497_new_n4368_), .Y(_abc_15497_new_n4384_));
AND2X2 AND2X2_1849 ( .A(_abc_15497_new_n4382_), .B(_abc_15497_new_n4386_), .Y(_abc_15497_new_n4387_));
AND2X2 AND2X2_185 ( .A(_abc_15497_new_n1082_), .B(_abc_15497_new_n1077_), .Y(_abc_15497_new_n1095_));
AND2X2 AND2X2_1850 ( .A(_abc_15497_new_n4387_), .B(_abc_15497_new_n4377_), .Y(_abc_15497_new_n4388_));
AND2X2 AND2X2_1851 ( .A(e_reg_8_), .B(a_reg_3_), .Y(_abc_15497_new_n4392_));
AND2X2 AND2X2_1852 ( .A(_abc_15497_new_n4393_), .B(_abc_15497_new_n4391_), .Y(_abc_15497_new_n4394_));
AND2X2 AND2X2_1853 ( .A(_abc_15497_new_n4395_), .B(_abc_15497_new_n4390_), .Y(_abc_15497_new_n4396_));
AND2X2 AND2X2_1854 ( .A(_abc_15497_new_n4394_), .B(w_8_), .Y(_abc_15497_new_n4397_));
AND2X2 AND2X2_1855 ( .A(_abc_15497_new_n4399_), .B(_abc_15497_new_n4389_), .Y(_abc_15497_new_n4400_));
AND2X2 AND2X2_1856 ( .A(_abc_15497_new_n4406_), .B(_abc_15497_new_n4401_), .Y(_abc_15497_new_n4407_));
AND2X2 AND2X2_1857 ( .A(_abc_15497_new_n4408_), .B(_abc_15497_new_n4404_), .Y(_abc_15497_new_n4409_));
AND2X2 AND2X2_1858 ( .A(_abc_15497_new_n4409_), .B(_abc_15497_new_n4367_), .Y(_abc_15497_new_n4410_));
AND2X2 AND2X2_1859 ( .A(_abc_15497_new_n4411_), .B(_abc_15497_new_n4338_), .Y(_abc_15497_new_n4412_));
AND2X2 AND2X2_186 ( .A(_abc_15497_new_n1097_), .B(_abc_15497_new_n1094_), .Y(_abc_15497_new_n1098_));
AND2X2 AND2X2_1860 ( .A(_abc_15497_new_n4405_), .B(_abc_15497_new_n4407_), .Y(_abc_15497_new_n4413_));
AND2X2 AND2X2_1861 ( .A(_abc_15497_new_n4403_), .B(_abc_15497_new_n4388_), .Y(_abc_15497_new_n4414_));
AND2X2 AND2X2_1862 ( .A(_abc_15497_new_n4415_), .B(_abc_15497_new_n4412_), .Y(_abc_15497_new_n4416_));
AND2X2 AND2X2_1863 ( .A(_abc_15497_new_n4417_), .B(_abc_15497_new_n3774_), .Y(_abc_15497_new_n4418_));
AND2X2 AND2X2_1864 ( .A(_abc_15497_new_n4420_), .B(_abc_15497_new_n4419_), .Y(_abc_15497_new_n4421_));
AND2X2 AND2X2_1865 ( .A(_abc_15497_new_n4421_), .B(_abc_15497_new_n3784_), .Y(_abc_15497_new_n4422_));
AND2X2 AND2X2_1866 ( .A(_abc_15497_new_n4424_), .B(_abc_15497_new_n4366_), .Y(_abc_15497_new_n4425_));
AND2X2 AND2X2_1867 ( .A(_abc_15497_new_n4423_), .B(_abc_15497_new_n4348_), .Y(_abc_15497_new_n4426_));
AND2X2 AND2X2_1868 ( .A(_abc_15497_new_n4430_), .B(_abc_15497_new_n4042_), .Y(_abc_15497_new_n4431_));
AND2X2 AND2X2_1869 ( .A(_abc_15497_new_n4429_), .B(_abc_15497_new_n4431_), .Y(_abc_15497_new_n4432_));
AND2X2 AND2X2_187 ( .A(_abc_15497_new_n1098_), .B(digest_update), .Y(_abc_15497_new_n1099_));
AND2X2 AND2X2_1870 ( .A(_abc_15497_new_n4298_), .B(_abc_15497_new_n4436_), .Y(_abc_15497_new_n4437_));
AND2X2 AND2X2_1871 ( .A(_abc_15497_new_n4439_), .B(_abc_15497_new_n4438_), .Y(_abc_15497_new_n4440_));
AND2X2 AND2X2_1872 ( .A(_abc_15497_new_n4435_), .B(_abc_15497_new_n4440_), .Y(_abc_15497_new_n4441_));
AND2X2 AND2X2_1873 ( .A(_abc_15497_new_n4442_), .B(_abc_15497_new_n4428_), .Y(_abc_15497_new_n4444_));
AND2X2 AND2X2_1874 ( .A(_abc_15497_new_n4445_), .B(round_ctr_inc), .Y(_abc_15497_new_n4446_));
AND2X2 AND2X2_1875 ( .A(_abc_15497_new_n4446_), .B(_abc_15497_new_n4443_), .Y(_abc_15497_new_n4447_));
AND2X2 AND2X2_1876 ( .A(_abc_15497_new_n2010_), .B(a_reg_8_), .Y(_abc_15497_new_n4448_));
AND2X2 AND2X2_1877 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n2824_), .Y(_abc_15497_new_n4449_));
AND2X2 AND2X2_1878 ( .A(_abc_15497_new_n4445_), .B(_abc_15497_new_n4452_), .Y(_abc_15497_new_n4453_));
AND2X2 AND2X2_1879 ( .A(_abc_15497_new_n4454_), .B(_abc_15497_new_n4419_), .Y(_abc_15497_new_n4455_));
AND2X2 AND2X2_188 ( .A(_abc_15497_new_n1100_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n1101_));
AND2X2 AND2X2_1880 ( .A(_abc_15497_new_n4404_), .B(_abc_15497_new_n4406_), .Y(_abc_15497_new_n4457_));
AND2X2 AND2X2_1881 ( .A(b_reg_9_), .B(c_reg_9_), .Y(_abc_15497_new_n4460_));
AND2X2 AND2X2_1882 ( .A(_abc_15497_new_n4461_), .B(_abc_15497_new_n4459_), .Y(_abc_15497_new_n4462_));
AND2X2 AND2X2_1883 ( .A(_abc_15497_new_n4463_), .B(_abc_15497_new_n4458_), .Y(_abc_15497_new_n4464_));
AND2X2 AND2X2_1884 ( .A(_abc_15497_new_n4462_), .B(d_reg_9_), .Y(_abc_15497_new_n4465_));
AND2X2 AND2X2_1885 ( .A(_abc_15497_new_n4468_), .B(d_reg_9_), .Y(_abc_15497_new_n4469_));
AND2X2 AND2X2_1886 ( .A(_abc_15497_new_n3753_), .B(_abc_15497_new_n4470_), .Y(_abc_15497_new_n4471_));
AND2X2 AND2X2_1887 ( .A(_abc_15497_new_n4461_), .B(_abc_15497_new_n4458_), .Y(_abc_15497_new_n4474_));
AND2X2 AND2X2_1888 ( .A(_abc_15497_new_n4472_), .B(_abc_15497_new_n4476_), .Y(_abc_15497_new_n4477_));
AND2X2 AND2X2_1889 ( .A(_abc_15497_new_n4477_), .B(_abc_15497_new_n4467_), .Y(_abc_15497_new_n4478_));
AND2X2 AND2X2_189 ( .A(_abc_15497_new_n1097_), .B(_abc_15497_new_n1092_), .Y(_abc_15497_new_n1105_));
AND2X2 AND2X2_1890 ( .A(e_reg_9_), .B(a_reg_4_), .Y(_abc_15497_new_n4483_));
AND2X2 AND2X2_1891 ( .A(_abc_15497_new_n4484_), .B(_abc_15497_new_n4482_), .Y(_abc_15497_new_n4485_));
AND2X2 AND2X2_1892 ( .A(_abc_15497_new_n4486_), .B(_abc_15497_new_n4481_), .Y(_abc_15497_new_n4487_));
AND2X2 AND2X2_1893 ( .A(_abc_15497_new_n4485_), .B(w_9_), .Y(_abc_15497_new_n4488_));
AND2X2 AND2X2_1894 ( .A(_abc_15497_new_n4490_), .B(_abc_15497_new_n4480_), .Y(_abc_15497_new_n4491_));
AND2X2 AND2X2_1895 ( .A(_abc_15497_new_n4492_), .B(_abc_15497_new_n4493_), .Y(_abc_15497_new_n4494_));
AND2X2 AND2X2_1896 ( .A(_abc_15497_new_n4479_), .B(_abc_15497_new_n4494_), .Y(_abc_15497_new_n4495_));
AND2X2 AND2X2_1897 ( .A(_abc_15497_new_n4497_), .B(_abc_15497_new_n4478_), .Y(_abc_15497_new_n4498_));
AND2X2 AND2X2_1898 ( .A(_abc_15497_new_n4499_), .B(_abc_15497_new_n4457_), .Y(_abc_15497_new_n4500_));
AND2X2 AND2X2_1899 ( .A(_abc_15497_new_n4503_), .B(_abc_15497_new_n4502_), .Y(_abc_15497_new_n4504_));
AND2X2 AND2X2_19 ( .A(_abc_15497_new_n732_), .B(_abc_15497_new_n733_), .Y(_abc_15497_new_n734_));
AND2X2 AND2X2_190 ( .A(e_reg_7_), .B(\digest[7] ), .Y(_abc_15497_new_n1107_));
AND2X2 AND2X2_1900 ( .A(_abc_15497_new_n4504_), .B(_abc_15497_new_n4501_), .Y(_abc_15497_new_n4505_));
AND2X2 AND2X2_1901 ( .A(_abc_15497_new_n4506_), .B(_abc_15497_new_n4060_), .Y(_abc_15497_new_n4507_));
AND2X2 AND2X2_1902 ( .A(_abc_15497_new_n4508_), .B(_abc_15497_new_n4509_), .Y(_abc_15497_new_n4510_));
AND2X2 AND2X2_1903 ( .A(_abc_15497_new_n4510_), .B(_abc_15497_new_n4059_), .Y(_abc_15497_new_n4511_));
AND2X2 AND2X2_1904 ( .A(_abc_15497_new_n4513_), .B(_abc_15497_new_n4456_), .Y(_abc_15497_new_n4514_));
AND2X2 AND2X2_1905 ( .A(_abc_15497_new_n4512_), .B(_abc_15497_new_n4455_), .Y(_abc_15497_new_n4515_));
AND2X2 AND2X2_1906 ( .A(_abc_15497_new_n4520_), .B(round_ctr_inc), .Y(_abc_15497_new_n4521_));
AND2X2 AND2X2_1907 ( .A(_abc_15497_new_n4521_), .B(_abc_15497_new_n4517_), .Y(_abc_15497_new_n4522_));
AND2X2 AND2X2_1908 ( .A(_abc_15497_new_n2010_), .B(a_reg_9_), .Y(_abc_15497_new_n4523_));
AND2X2 AND2X2_1909 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n2838_), .Y(_abc_15497_new_n4524_));
AND2X2 AND2X2_191 ( .A(_abc_15497_new_n1108_), .B(_abc_15497_new_n1106_), .Y(_abc_15497_new_n1109_));
AND2X2 AND2X2_1910 ( .A(_abc_15497_new_n4528_), .B(_abc_15497_new_n4527_), .Y(_abc_15497_new_n4529_));
AND2X2 AND2X2_1911 ( .A(_abc_15497_new_n4442_), .B(_abc_15497_new_n4532_), .Y(_abc_15497_new_n4533_));
AND2X2 AND2X2_1912 ( .A(b_reg_10_), .B(c_reg_10_), .Y(_abc_15497_new_n4539_));
AND2X2 AND2X2_1913 ( .A(_abc_15497_new_n4540_), .B(_abc_15497_new_n4538_), .Y(_abc_15497_new_n4541_));
AND2X2 AND2X2_1914 ( .A(_abc_15497_new_n4542_), .B(_abc_15497_new_n4537_), .Y(_abc_15497_new_n4543_));
AND2X2 AND2X2_1915 ( .A(_abc_15497_new_n4541_), .B(d_reg_10_), .Y(_abc_15497_new_n4544_));
AND2X2 AND2X2_1916 ( .A(_abc_15497_new_n4547_), .B(d_reg_10_), .Y(_abc_15497_new_n4548_));
AND2X2 AND2X2_1917 ( .A(_abc_15497_new_n3753_), .B(_abc_15497_new_n4549_), .Y(_abc_15497_new_n4550_));
AND2X2 AND2X2_1918 ( .A(_abc_15497_new_n4540_), .B(_abc_15497_new_n4537_), .Y(_abc_15497_new_n4553_));
AND2X2 AND2X2_1919 ( .A(_abc_15497_new_n4551_), .B(_abc_15497_new_n4555_), .Y(_abc_15497_new_n4556_));
AND2X2 AND2X2_192 ( .A(_abc_15497_new_n1105_), .B(_abc_15497_new_n1109_), .Y(_abc_15497_new_n1110_));
AND2X2 AND2X2_1920 ( .A(_abc_15497_new_n4556_), .B(_abc_15497_new_n4546_), .Y(_abc_15497_new_n4557_));
AND2X2 AND2X2_1921 ( .A(e_reg_10_), .B(a_reg_5_), .Y(_abc_15497_new_n4561_));
AND2X2 AND2X2_1922 ( .A(_abc_15497_new_n4562_), .B(_abc_15497_new_n4560_), .Y(_abc_15497_new_n4563_));
AND2X2 AND2X2_1923 ( .A(_abc_15497_new_n4564_), .B(_abc_15497_new_n4559_), .Y(_abc_15497_new_n4565_));
AND2X2 AND2X2_1924 ( .A(_abc_15497_new_n4563_), .B(w_10_), .Y(_abc_15497_new_n4566_));
AND2X2 AND2X2_1925 ( .A(_abc_15497_new_n4568_), .B(_abc_15497_new_n4558_), .Y(_abc_15497_new_n4569_));
AND2X2 AND2X2_1926 ( .A(_abc_15497_new_n4575_), .B(_abc_15497_new_n4570_), .Y(_abc_15497_new_n4576_));
AND2X2 AND2X2_1927 ( .A(_abc_15497_new_n4577_), .B(_abc_15497_new_n4573_), .Y(_abc_15497_new_n4578_));
AND2X2 AND2X2_1928 ( .A(_abc_15497_new_n4502_), .B(_abc_15497_new_n4492_), .Y(_abc_15497_new_n4580_));
AND2X2 AND2X2_1929 ( .A(_abc_15497_new_n4574_), .B(_abc_15497_new_n4576_), .Y(_abc_15497_new_n4581_));
AND2X2 AND2X2_193 ( .A(_abc_15497_new_n1089_), .B(_abc_15497_new_n1093_), .Y(_abc_15497_new_n1111_));
AND2X2 AND2X2_1930 ( .A(_abc_15497_new_n4572_), .B(_abc_15497_new_n4557_), .Y(_abc_15497_new_n4582_));
AND2X2 AND2X2_1931 ( .A(_abc_15497_new_n4579_), .B(_abc_15497_new_n4584_), .Y(_abc_15497_new_n4585_));
AND2X2 AND2X2_1932 ( .A(_abc_15497_new_n4583_), .B(_abc_15497_new_n4580_), .Y(_abc_15497_new_n4587_));
AND2X2 AND2X2_1933 ( .A(_abc_15497_new_n4578_), .B(_abc_15497_new_n4536_), .Y(_abc_15497_new_n4588_));
AND2X2 AND2X2_1934 ( .A(_abc_15497_new_n4590_), .B(_abc_15497_new_n4586_), .Y(_abc_15497_new_n4591_));
AND2X2 AND2X2_1935 ( .A(_abc_15497_new_n4591_), .B(_abc_15497_new_n4535_), .Y(_abc_15497_new_n4592_));
AND2X2 AND2X2_1936 ( .A(_abc_15497_new_n4593_), .B(_abc_15497_new_n4509_), .Y(_abc_15497_new_n4594_));
AND2X2 AND2X2_1937 ( .A(_abc_15497_new_n4589_), .B(_abc_15497_new_n3784_), .Y(_abc_15497_new_n4595_));
AND2X2 AND2X2_1938 ( .A(_abc_15497_new_n4585_), .B(_abc_15497_new_n3774_), .Y(_abc_15497_new_n4596_));
AND2X2 AND2X2_1939 ( .A(_abc_15497_new_n4597_), .B(_abc_15497_new_n4594_), .Y(_abc_15497_new_n4598_));
AND2X2 AND2X2_194 ( .A(_abc_15497_new_n1112_), .B(_abc_15497_new_n1113_), .Y(_abc_15497_new_n1114_));
AND2X2 AND2X2_1940 ( .A(_abc_15497_new_n4534_), .B(_abc_15497_new_n4600_), .Y(_abc_15497_new_n4602_));
AND2X2 AND2X2_1941 ( .A(_abc_15497_new_n4603_), .B(round_ctr_inc), .Y(_abc_15497_new_n4604_));
AND2X2 AND2X2_1942 ( .A(_abc_15497_new_n4604_), .B(_abc_15497_new_n4601_), .Y(_abc_15497_new_n4605_));
AND2X2 AND2X2_1943 ( .A(_abc_15497_new_n2010_), .B(a_reg_10_), .Y(_abc_15497_new_n4606_));
AND2X2 AND2X2_1944 ( .A(_abc_15497_new_n700_), .B(\digest[138] ), .Y(_abc_15497_new_n4607_));
AND2X2 AND2X2_1945 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n4607_), .Y(_abc_15497_new_n4608_));
AND2X2 AND2X2_1946 ( .A(_abc_15497_new_n4603_), .B(_abc_15497_new_n4611_), .Y(_abc_15497_new_n4612_));
AND2X2 AND2X2_1947 ( .A(_abc_15497_new_n4573_), .B(_abc_15497_new_n4575_), .Y(_abc_15497_new_n4614_));
AND2X2 AND2X2_1948 ( .A(b_reg_11_), .B(c_reg_11_), .Y(_abc_15497_new_n4617_));
AND2X2 AND2X2_1949 ( .A(_abc_15497_new_n4618_), .B(_abc_15497_new_n4616_), .Y(_abc_15497_new_n4619_));
AND2X2 AND2X2_195 ( .A(_abc_15497_new_n1116_), .B(_abc_15497_new_n1104_), .Y(_0H4_reg_31_0__7_));
AND2X2 AND2X2_1950 ( .A(_abc_15497_new_n4620_), .B(_abc_15497_new_n4615_), .Y(_abc_15497_new_n4621_));
AND2X2 AND2X2_1951 ( .A(_abc_15497_new_n4619_), .B(d_reg_11_), .Y(_abc_15497_new_n4622_));
AND2X2 AND2X2_1952 ( .A(_abc_15497_new_n4625_), .B(d_reg_11_), .Y(_abc_15497_new_n4626_));
AND2X2 AND2X2_1953 ( .A(_abc_15497_new_n3753_), .B(_abc_15497_new_n4627_), .Y(_abc_15497_new_n4628_));
AND2X2 AND2X2_1954 ( .A(_abc_15497_new_n4618_), .B(_abc_15497_new_n4615_), .Y(_abc_15497_new_n4631_));
AND2X2 AND2X2_1955 ( .A(_abc_15497_new_n4629_), .B(_abc_15497_new_n4633_), .Y(_abc_15497_new_n4634_));
AND2X2 AND2X2_1956 ( .A(_abc_15497_new_n4634_), .B(_abc_15497_new_n4624_), .Y(_abc_15497_new_n4635_));
AND2X2 AND2X2_1957 ( .A(e_reg_11_), .B(a_reg_6_), .Y(_abc_15497_new_n4640_));
AND2X2 AND2X2_1958 ( .A(_abc_15497_new_n4641_), .B(_abc_15497_new_n4639_), .Y(_abc_15497_new_n4642_));
AND2X2 AND2X2_1959 ( .A(_abc_15497_new_n4643_), .B(_abc_15497_new_n4638_), .Y(_abc_15497_new_n4644_));
AND2X2 AND2X2_196 ( .A(e_reg_8_), .B(\digest[8] ), .Y(_abc_15497_new_n1119_));
AND2X2 AND2X2_1960 ( .A(_abc_15497_new_n4642_), .B(w_11_), .Y(_abc_15497_new_n4645_));
AND2X2 AND2X2_1961 ( .A(_abc_15497_new_n4647_), .B(_abc_15497_new_n4637_), .Y(_abc_15497_new_n4648_));
AND2X2 AND2X2_1962 ( .A(_abc_15497_new_n4649_), .B(_abc_15497_new_n4650_), .Y(_abc_15497_new_n4651_));
AND2X2 AND2X2_1963 ( .A(_abc_15497_new_n4636_), .B(_abc_15497_new_n4651_), .Y(_abc_15497_new_n4652_));
AND2X2 AND2X2_1964 ( .A(_abc_15497_new_n4654_), .B(_abc_15497_new_n4635_), .Y(_abc_15497_new_n4655_));
AND2X2 AND2X2_1965 ( .A(_abc_15497_new_n4660_), .B(_abc_15497_new_n4659_), .Y(_abc_15497_new_n4661_));
AND2X2 AND2X2_1966 ( .A(_abc_15497_new_n4662_), .B(_abc_15497_new_n4657_), .Y(_abc_15497_new_n4663_));
AND2X2 AND2X2_1967 ( .A(_abc_15497_new_n4661_), .B(_abc_15497_new_n4658_), .Y(_abc_15497_new_n4665_));
AND2X2 AND2X2_1968 ( .A(_abc_15497_new_n4656_), .B(_abc_15497_new_n4614_), .Y(_abc_15497_new_n4666_));
AND2X2 AND2X2_1969 ( .A(_abc_15497_new_n4664_), .B(_abc_15497_new_n4668_), .Y(_abc_15497_new_n4669_));
AND2X2 AND2X2_197 ( .A(_abc_15497_new_n1120_), .B(_abc_15497_new_n1118_), .Y(_abc_15497_new_n1121_));
AND2X2 AND2X2_1970 ( .A(_abc_15497_new_n4669_), .B(_abc_15497_new_n4613_), .Y(_abc_15497_new_n4670_));
AND2X2 AND2X2_1971 ( .A(_abc_15497_new_n4590_), .B(_abc_15497_new_n4584_), .Y(_abc_15497_new_n4671_));
AND2X2 AND2X2_1972 ( .A(_abc_15497_new_n4667_), .B(_abc_15497_new_n3783_), .Y(_abc_15497_new_n4672_));
AND2X2 AND2X2_1973 ( .A(_abc_15497_new_n4663_), .B(_abc_15497_new_n3773_), .Y(_abc_15497_new_n4673_));
AND2X2 AND2X2_1974 ( .A(_abc_15497_new_n4674_), .B(_abc_15497_new_n4671_), .Y(_abc_15497_new_n4675_));
AND2X2 AND2X2_1975 ( .A(_abc_15497_new_n4680_), .B(round_ctr_inc), .Y(_abc_15497_new_n4681_));
AND2X2 AND2X2_1976 ( .A(_abc_15497_new_n4681_), .B(_abc_15497_new_n4677_), .Y(_abc_15497_new_n4682_));
AND2X2 AND2X2_1977 ( .A(_abc_15497_new_n2010_), .B(a_reg_11_), .Y(_abc_15497_new_n4683_));
AND2X2 AND2X2_1978 ( .A(_abc_15497_new_n700_), .B(\digest[139] ), .Y(_abc_15497_new_n4684_));
AND2X2 AND2X2_1979 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n4684_), .Y(_abc_15497_new_n4685_));
AND2X2 AND2X2_198 ( .A(_abc_15497_new_n1112_), .B(_abc_15497_new_n1106_), .Y(_abc_15497_new_n1122_));
AND2X2 AND2X2_1980 ( .A(_abc_15497_new_n4691_), .B(_abc_15497_new_n4690_), .Y(_abc_15497_new_n4692_));
AND2X2 AND2X2_1981 ( .A(_abc_15497_new_n4689_), .B(_abc_15497_new_n4692_), .Y(_abc_15497_new_n4693_));
AND2X2 AND2X2_1982 ( .A(_abc_15497_new_n4442_), .B(_abc_15497_new_n4696_), .Y(_abc_15497_new_n4697_));
AND2X2 AND2X2_1983 ( .A(_abc_15497_new_n4668_), .B(_abc_15497_new_n4657_), .Y(_abc_15497_new_n4699_));
AND2X2 AND2X2_1984 ( .A(_abc_15497_new_n4659_), .B(_abc_15497_new_n4649_), .Y(_abc_15497_new_n4700_));
AND2X2 AND2X2_1985 ( .A(b_reg_12_), .B(c_reg_12_), .Y(_abc_15497_new_n4703_));
AND2X2 AND2X2_1986 ( .A(_abc_15497_new_n4704_), .B(_abc_15497_new_n4702_), .Y(_abc_15497_new_n4705_));
AND2X2 AND2X2_1987 ( .A(_abc_15497_new_n4705_), .B(d_reg_12_), .Y(_abc_15497_new_n4707_));
AND2X2 AND2X2_1988 ( .A(_abc_15497_new_n4708_), .B(_abc_15497_new_n4706_), .Y(_abc_15497_new_n4709_));
AND2X2 AND2X2_1989 ( .A(_abc_15497_new_n3803_), .B(_abc_15497_new_n4709_), .Y(_abc_15497_new_n4710_));
AND2X2 AND2X2_199 ( .A(_abc_15497_new_n1123_), .B(_abc_15497_new_n1121_), .Y(_abc_15497_new_n1125_));
AND2X2 AND2X2_1990 ( .A(_abc_15497_new_n4713_), .B(_abc_15497_new_n4704_), .Y(_abc_15497_new_n4714_));
AND2X2 AND2X2_1991 ( .A(_abc_15497_new_n4704_), .B(_abc_15497_new_n4712_), .Y(_abc_15497_new_n4717_));
AND2X2 AND2X2_1992 ( .A(_abc_15497_new_n4719_), .B(_abc_15497_new_n4715_), .Y(_abc_15497_new_n4720_));
AND2X2 AND2X2_1993 ( .A(_abc_15497_new_n4711_), .B(_abc_15497_new_n4720_), .Y(_abc_15497_new_n4721_));
AND2X2 AND2X2_1994 ( .A(e_reg_12_), .B(a_reg_7_), .Y(_abc_15497_new_n4726_));
AND2X2 AND2X2_1995 ( .A(_abc_15497_new_n4727_), .B(_abc_15497_new_n4725_), .Y(_abc_15497_new_n4728_));
AND2X2 AND2X2_1996 ( .A(_abc_15497_new_n4729_), .B(_abc_15497_new_n4724_), .Y(_abc_15497_new_n4730_));
AND2X2 AND2X2_1997 ( .A(_abc_15497_new_n4728_), .B(w_12_), .Y(_abc_15497_new_n4731_));
AND2X2 AND2X2_1998 ( .A(_abc_15497_new_n4733_), .B(_abc_15497_new_n4723_), .Y(_abc_15497_new_n4734_));
AND2X2 AND2X2_1999 ( .A(_abc_15497_new_n4735_), .B(_abc_15497_new_n4736_), .Y(_abc_15497_new_n4737_));
AND2X2 AND2X2_2 ( .A(_abc_15497_new_n700_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n701_));
AND2X2 AND2X2_20 ( .A(c_reg_18_), .B(\digest[82] ), .Y(_abc_15497_new_n735_));
AND2X2 AND2X2_200 ( .A(_abc_15497_new_n1126_), .B(_abc_15497_new_n1124_), .Y(_abc_15497_new_n1127_));
AND2X2 AND2X2_2000 ( .A(_abc_15497_new_n4722_), .B(_abc_15497_new_n4737_), .Y(_abc_15497_new_n4738_));
AND2X2 AND2X2_2001 ( .A(_abc_15497_new_n4739_), .B(_abc_15497_new_n4740_), .Y(_abc_15497_new_n4741_));
AND2X2 AND2X2_2002 ( .A(_abc_15497_new_n4701_), .B(_abc_15497_new_n4741_), .Y(_abc_15497_new_n4743_));
AND2X2 AND2X2_2003 ( .A(_abc_15497_new_n4744_), .B(_abc_15497_new_n4742_), .Y(_abc_15497_new_n4745_));
AND2X2 AND2X2_2004 ( .A(_abc_15497_new_n4745_), .B(_abc_15497_new_n3775_), .Y(_abc_15497_new_n4746_));
AND2X2 AND2X2_2005 ( .A(_abc_15497_new_n4748_), .B(_abc_15497_new_n4700_), .Y(_abc_15497_new_n4749_));
AND2X2 AND2X2_2006 ( .A(_abc_15497_new_n4750_), .B(_abc_15497_new_n3803_), .Y(_abc_15497_new_n4751_));
AND2X2 AND2X2_2007 ( .A(_abc_15497_new_n4752_), .B(_abc_15497_new_n4699_), .Y(_abc_15497_new_n4753_));
AND2X2 AND2X2_2008 ( .A(_abc_15497_new_n4756_), .B(_abc_15497_new_n4755_), .Y(_abc_15497_new_n4757_));
AND2X2 AND2X2_2009 ( .A(_abc_15497_new_n4757_), .B(_abc_15497_new_n4754_), .Y(_abc_15497_new_n4758_));
AND2X2 AND2X2_201 ( .A(_abc_15497_new_n1127_), .B(digest_update), .Y(_abc_15497_new_n1128_));
AND2X2 AND2X2_2010 ( .A(_abc_15497_new_n4698_), .B(_abc_15497_new_n4760_), .Y(_abc_15497_new_n4762_));
AND2X2 AND2X2_2011 ( .A(_abc_15497_new_n4763_), .B(round_ctr_inc), .Y(_abc_15497_new_n4764_));
AND2X2 AND2X2_2012 ( .A(_abc_15497_new_n4764_), .B(_abc_15497_new_n4761_), .Y(_abc_15497_new_n4765_));
AND2X2 AND2X2_2013 ( .A(_abc_15497_new_n2010_), .B(a_reg_12_), .Y(_abc_15497_new_n4766_));
AND2X2 AND2X2_2014 ( .A(_abc_15497_new_n700_), .B(\digest[140] ), .Y(_abc_15497_new_n4767_));
AND2X2 AND2X2_2015 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n4767_), .Y(_abc_15497_new_n4768_));
AND2X2 AND2X2_2016 ( .A(_abc_15497_new_n4763_), .B(_abc_15497_new_n4771_), .Y(_abc_15497_new_n4772_));
AND2X2 AND2X2_2017 ( .A(b_reg_13_), .B(c_reg_13_), .Y(_abc_15497_new_n4776_));
AND2X2 AND2X2_2018 ( .A(_abc_15497_new_n4777_), .B(_abc_15497_new_n4775_), .Y(_abc_15497_new_n4778_));
AND2X2 AND2X2_2019 ( .A(_abc_15497_new_n4778_), .B(d_reg_13_), .Y(_abc_15497_new_n4780_));
AND2X2 AND2X2_202 ( .A(_abc_15497_new_n1129_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n1130_));
AND2X2 AND2X2_2020 ( .A(_abc_15497_new_n4781_), .B(_abc_15497_new_n4779_), .Y(_abc_15497_new_n4782_));
AND2X2 AND2X2_2021 ( .A(_abc_15497_new_n3803_), .B(_abc_15497_new_n4782_), .Y(_abc_15497_new_n4783_));
AND2X2 AND2X2_2022 ( .A(_abc_15497_new_n4786_), .B(_abc_15497_new_n4777_), .Y(_abc_15497_new_n4787_));
AND2X2 AND2X2_2023 ( .A(_abc_15497_new_n4777_), .B(_abc_15497_new_n4785_), .Y(_abc_15497_new_n4790_));
AND2X2 AND2X2_2024 ( .A(_abc_15497_new_n4792_), .B(_abc_15497_new_n4788_), .Y(_abc_15497_new_n4793_));
AND2X2 AND2X2_2025 ( .A(_abc_15497_new_n4784_), .B(_abc_15497_new_n4793_), .Y(_abc_15497_new_n4794_));
AND2X2 AND2X2_2026 ( .A(e_reg_13_), .B(a_reg_8_), .Y(_abc_15497_new_n4799_));
AND2X2 AND2X2_2027 ( .A(_abc_15497_new_n4800_), .B(_abc_15497_new_n4798_), .Y(_abc_15497_new_n4801_));
AND2X2 AND2X2_2028 ( .A(_abc_15497_new_n4802_), .B(_abc_15497_new_n4797_), .Y(_abc_15497_new_n4803_));
AND2X2 AND2X2_2029 ( .A(_abc_15497_new_n4801_), .B(w_13_), .Y(_abc_15497_new_n4804_));
AND2X2 AND2X2_203 ( .A(_abc_15497_new_n701_), .B(\digest[9] ), .Y(_abc_15497_new_n1132_));
AND2X2 AND2X2_2030 ( .A(_abc_15497_new_n4806_), .B(_abc_15497_new_n4796_), .Y(_abc_15497_new_n4807_));
AND2X2 AND2X2_2031 ( .A(_abc_15497_new_n4808_), .B(_abc_15497_new_n4809_), .Y(_abc_15497_new_n4810_));
AND2X2 AND2X2_2032 ( .A(_abc_15497_new_n4795_), .B(_abc_15497_new_n4810_), .Y(_abc_15497_new_n4811_));
AND2X2 AND2X2_2033 ( .A(_abc_15497_new_n4812_), .B(_abc_15497_new_n4813_), .Y(_abc_15497_new_n4814_));
AND2X2 AND2X2_2034 ( .A(_abc_15497_new_n4814_), .B(_abc_15497_new_n4774_), .Y(_abc_15497_new_n4816_));
AND2X2 AND2X2_2035 ( .A(_abc_15497_new_n4817_), .B(_abc_15497_new_n4815_), .Y(_abc_15497_new_n4818_));
AND2X2 AND2X2_2036 ( .A(_abc_15497_new_n4822_), .B(_abc_15497_new_n4820_), .Y(_abc_15497_new_n4823_));
AND2X2 AND2X2_2037 ( .A(_abc_15497_new_n4819_), .B(_abc_15497_new_n4825_), .Y(_abc_15497_new_n4826_));
AND2X2 AND2X2_2038 ( .A(_abc_15497_new_n4773_), .B(_abc_15497_new_n4826_), .Y(_abc_15497_new_n4827_));
AND2X2 AND2X2_2039 ( .A(_abc_15497_new_n4755_), .B(_abc_15497_new_n4744_), .Y(_abc_15497_new_n4828_));
AND2X2 AND2X2_204 ( .A(e_reg_9_), .B(\digest[9] ), .Y(_abc_15497_new_n1134_));
AND2X2 AND2X2_2040 ( .A(_abc_15497_new_n4824_), .B(_abc_15497_new_n3783_), .Y(_abc_15497_new_n4829_));
AND2X2 AND2X2_2041 ( .A(_abc_15497_new_n4818_), .B(_abc_15497_new_n3773_), .Y(_abc_15497_new_n4830_));
AND2X2 AND2X2_2042 ( .A(_abc_15497_new_n4831_), .B(_abc_15497_new_n4828_), .Y(_abc_15497_new_n4832_));
AND2X2 AND2X2_2043 ( .A(_abc_15497_new_n4837_), .B(round_ctr_inc), .Y(_abc_15497_new_n4838_));
AND2X2 AND2X2_2044 ( .A(_abc_15497_new_n4838_), .B(_abc_15497_new_n4834_), .Y(_abc_15497_new_n4839_));
AND2X2 AND2X2_2045 ( .A(_abc_15497_new_n2010_), .B(a_reg_13_), .Y(_abc_15497_new_n4840_));
AND2X2 AND2X2_2046 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n2903_), .Y(_abc_15497_new_n4841_));
AND2X2 AND2X2_2047 ( .A(_abc_15497_new_n4845_), .B(_abc_15497_new_n4844_), .Y(_abc_15497_new_n4846_));
AND2X2 AND2X2_2048 ( .A(_abc_15497_new_n4698_), .B(_abc_15497_new_n4849_), .Y(_abc_15497_new_n4850_));
AND2X2 AND2X2_2049 ( .A(b_reg_14_), .B(c_reg_14_), .Y(_abc_15497_new_n4855_));
AND2X2 AND2X2_205 ( .A(_abc_15497_new_n1135_), .B(_abc_15497_new_n1133_), .Y(_abc_15497_new_n1136_));
AND2X2 AND2X2_2050 ( .A(_abc_15497_new_n4856_), .B(_abc_15497_new_n4854_), .Y(_abc_15497_new_n4857_));
AND2X2 AND2X2_2051 ( .A(_abc_15497_new_n4857_), .B(d_reg_14_), .Y(_abc_15497_new_n4859_));
AND2X2 AND2X2_2052 ( .A(_abc_15497_new_n4860_), .B(_abc_15497_new_n4858_), .Y(_abc_15497_new_n4861_));
AND2X2 AND2X2_2053 ( .A(_abc_15497_new_n3803_), .B(_abc_15497_new_n4861_), .Y(_abc_15497_new_n4862_));
AND2X2 AND2X2_2054 ( .A(_abc_15497_new_n4865_), .B(_abc_15497_new_n4856_), .Y(_abc_15497_new_n4866_));
AND2X2 AND2X2_2055 ( .A(_abc_15497_new_n4856_), .B(_abc_15497_new_n4864_), .Y(_abc_15497_new_n4868_));
AND2X2 AND2X2_2056 ( .A(_abc_15497_new_n4869_), .B(_abc_15497_new_n4854_), .Y(_abc_15497_new_n4870_));
AND2X2 AND2X2_2057 ( .A(_abc_15497_new_n3774_), .B(_abc_15497_new_n4870_), .Y(_abc_15497_new_n4871_));
AND2X2 AND2X2_2058 ( .A(_abc_15497_new_n4872_), .B(_abc_15497_new_n4867_), .Y(_abc_15497_new_n4873_));
AND2X2 AND2X2_2059 ( .A(_abc_15497_new_n4863_), .B(_abc_15497_new_n4873_), .Y(_abc_15497_new_n4874_));
AND2X2 AND2X2_206 ( .A(_abc_15497_new_n1121_), .B(_abc_15497_new_n1136_), .Y(_abc_15497_new_n1137_));
AND2X2 AND2X2_2060 ( .A(e_reg_14_), .B(a_reg_9_), .Y(_abc_15497_new_n4878_));
AND2X2 AND2X2_2061 ( .A(_abc_15497_new_n4879_), .B(_abc_15497_new_n4877_), .Y(_abc_15497_new_n4880_));
AND2X2 AND2X2_2062 ( .A(_abc_15497_new_n4880_), .B(w_14_), .Y(_abc_15497_new_n4882_));
AND2X2 AND2X2_2063 ( .A(_abc_15497_new_n4883_), .B(_abc_15497_new_n4881_), .Y(_abc_15497_new_n4884_));
AND2X2 AND2X2_2064 ( .A(_abc_15497_new_n4884_), .B(_abc_15497_new_n4876_), .Y(_abc_15497_new_n4885_));
AND2X2 AND2X2_2065 ( .A(_abc_15497_new_n4886_), .B(_abc_15497_new_n4887_), .Y(_abc_15497_new_n4888_));
AND2X2 AND2X2_2066 ( .A(_abc_15497_new_n4875_), .B(_abc_15497_new_n4888_), .Y(_abc_15497_new_n4889_));
AND2X2 AND2X2_2067 ( .A(_abc_15497_new_n4890_), .B(_abc_15497_new_n4891_), .Y(_abc_15497_new_n4892_));
AND2X2 AND2X2_2068 ( .A(_abc_15497_new_n4897_), .B(_abc_15497_new_n4893_), .Y(_abc_15497_new_n4898_));
AND2X2 AND2X2_2069 ( .A(_abc_15497_new_n4896_), .B(_abc_15497_new_n4894_), .Y(_abc_15497_new_n4900_));
AND2X2 AND2X2_207 ( .A(_abc_15497_new_n1123_), .B(_abc_15497_new_n1137_), .Y(_abc_15497_new_n1138_));
AND2X2 AND2X2_2070 ( .A(_abc_15497_new_n4892_), .B(_abc_15497_new_n4853_), .Y(_abc_15497_new_n4901_));
AND2X2 AND2X2_2071 ( .A(_abc_15497_new_n4899_), .B(_abc_15497_new_n4903_), .Y(_abc_15497_new_n4904_));
AND2X2 AND2X2_2072 ( .A(_abc_15497_new_n4852_), .B(_abc_15497_new_n4904_), .Y(_abc_15497_new_n4905_));
AND2X2 AND2X2_2073 ( .A(_abc_15497_new_n4825_), .B(_abc_15497_new_n4817_), .Y(_abc_15497_new_n4906_));
AND2X2 AND2X2_2074 ( .A(_abc_15497_new_n4902_), .B(_abc_15497_new_n3774_), .Y(_abc_15497_new_n4907_));
AND2X2 AND2X2_2075 ( .A(_abc_15497_new_n4898_), .B(_abc_15497_new_n3784_), .Y(_abc_15497_new_n4908_));
AND2X2 AND2X2_2076 ( .A(_abc_15497_new_n4909_), .B(_abc_15497_new_n4906_), .Y(_abc_15497_new_n4910_));
AND2X2 AND2X2_2077 ( .A(_abc_15497_new_n4851_), .B(_abc_15497_new_n4912_), .Y(_abc_15497_new_n4914_));
AND2X2 AND2X2_2078 ( .A(_abc_15497_new_n4915_), .B(round_ctr_inc), .Y(_abc_15497_new_n4916_));
AND2X2 AND2X2_2079 ( .A(_abc_15497_new_n4916_), .B(_abc_15497_new_n4913_), .Y(_abc_15497_new_n4917_));
AND2X2 AND2X2_208 ( .A(_abc_15497_new_n1136_), .B(_abc_15497_new_n1119_), .Y(_abc_15497_new_n1142_));
AND2X2 AND2X2_2080 ( .A(_abc_15497_new_n2010_), .B(a_reg_14_), .Y(_abc_15497_new_n4918_));
AND2X2 AND2X2_2081 ( .A(_abc_15497_new_n700_), .B(\digest[142] ), .Y(_abc_15497_new_n4919_));
AND2X2 AND2X2_2082 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n4919_), .Y(_abc_15497_new_n4920_));
AND2X2 AND2X2_2083 ( .A(_abc_15497_new_n4915_), .B(_abc_15497_new_n4923_), .Y(_abc_15497_new_n4924_));
AND2X2 AND2X2_2084 ( .A(b_reg_15_), .B(c_reg_15_), .Y(_abc_15497_new_n4928_));
AND2X2 AND2X2_2085 ( .A(_abc_15497_new_n4929_), .B(_abc_15497_new_n4927_), .Y(_abc_15497_new_n4930_));
AND2X2 AND2X2_2086 ( .A(_abc_15497_new_n4930_), .B(d_reg_15_), .Y(_abc_15497_new_n4932_));
AND2X2 AND2X2_2087 ( .A(_abc_15497_new_n4933_), .B(_abc_15497_new_n4931_), .Y(_abc_15497_new_n4934_));
AND2X2 AND2X2_2088 ( .A(_abc_15497_new_n3803_), .B(_abc_15497_new_n4934_), .Y(_abc_15497_new_n4935_));
AND2X2 AND2X2_2089 ( .A(_abc_15497_new_n4938_), .B(_abc_15497_new_n4929_), .Y(_abc_15497_new_n4939_));
AND2X2 AND2X2_209 ( .A(_abc_15497_new_n1143_), .B(digest_update), .Y(_abc_15497_new_n1144_));
AND2X2 AND2X2_2090 ( .A(_abc_15497_new_n4929_), .B(_abc_15497_new_n4937_), .Y(_abc_15497_new_n4941_));
AND2X2 AND2X2_2091 ( .A(_abc_15497_new_n4942_), .B(_abc_15497_new_n4927_), .Y(_abc_15497_new_n4943_));
AND2X2 AND2X2_2092 ( .A(_abc_15497_new_n3774_), .B(_abc_15497_new_n4943_), .Y(_abc_15497_new_n4944_));
AND2X2 AND2X2_2093 ( .A(_abc_15497_new_n4945_), .B(_abc_15497_new_n4940_), .Y(_abc_15497_new_n4946_));
AND2X2 AND2X2_2094 ( .A(_abc_15497_new_n4936_), .B(_abc_15497_new_n4946_), .Y(_abc_15497_new_n4947_));
AND2X2 AND2X2_2095 ( .A(e_reg_15_), .B(a_reg_10_), .Y(_abc_15497_new_n4951_));
AND2X2 AND2X2_2096 ( .A(_abc_15497_new_n4952_), .B(_abc_15497_new_n4950_), .Y(_abc_15497_new_n4953_));
AND2X2 AND2X2_2097 ( .A(_abc_15497_new_n4953_), .B(w_15_), .Y(_abc_15497_new_n4955_));
AND2X2 AND2X2_2098 ( .A(_abc_15497_new_n4956_), .B(_abc_15497_new_n4954_), .Y(_abc_15497_new_n4957_));
AND2X2 AND2X2_2099 ( .A(_abc_15497_new_n4957_), .B(_abc_15497_new_n4949_), .Y(_abc_15497_new_n4958_));
AND2X2 AND2X2_21 ( .A(_abc_15497_new_n736_), .B(_abc_15497_new_n737_), .Y(_abc_15497_new_n738_));
AND2X2 AND2X2_210 ( .A(_abc_15497_new_n1141_), .B(_abc_15497_new_n1144_), .Y(_abc_15497_new_n1145_));
AND2X2 AND2X2_2100 ( .A(_abc_15497_new_n4959_), .B(_abc_15497_new_n4960_), .Y(_abc_15497_new_n4961_));
AND2X2 AND2X2_2101 ( .A(_abc_15497_new_n4948_), .B(_abc_15497_new_n4961_), .Y(_abc_15497_new_n4962_));
AND2X2 AND2X2_2102 ( .A(_abc_15497_new_n4963_), .B(_abc_15497_new_n4964_), .Y(_abc_15497_new_n4965_));
AND2X2 AND2X2_2103 ( .A(_abc_15497_new_n4965_), .B(_abc_15497_new_n4926_), .Y(_abc_15497_new_n4967_));
AND2X2 AND2X2_2104 ( .A(_abc_15497_new_n4968_), .B(_abc_15497_new_n4966_), .Y(_abc_15497_new_n4969_));
AND2X2 AND2X2_2105 ( .A(_abc_15497_new_n4973_), .B(_abc_15497_new_n4971_), .Y(_abc_15497_new_n4974_));
AND2X2 AND2X2_2106 ( .A(_abc_15497_new_n4970_), .B(_abc_15497_new_n4976_), .Y(_abc_15497_new_n4977_));
AND2X2 AND2X2_2107 ( .A(_abc_15497_new_n4977_), .B(_abc_15497_new_n4925_), .Y(_abc_15497_new_n4978_));
AND2X2 AND2X2_2108 ( .A(_abc_15497_new_n4903_), .B(_abc_15497_new_n4897_), .Y(_abc_15497_new_n4979_));
AND2X2 AND2X2_2109 ( .A(_abc_15497_new_n4975_), .B(_abc_15497_new_n3753_), .Y(_abc_15497_new_n4980_));
AND2X2 AND2X2_211 ( .A(_abc_15497_new_n1145_), .B(_abc_15497_new_n1139_), .Y(_abc_15497_new_n1146_));
AND2X2 AND2X2_2110 ( .A(_abc_15497_new_n4969_), .B(_abc_15497_new_n3780_), .Y(_abc_15497_new_n4981_));
AND2X2 AND2X2_2111 ( .A(_abc_15497_new_n4982_), .B(_abc_15497_new_n4979_), .Y(_abc_15497_new_n4983_));
AND2X2 AND2X2_2112 ( .A(_abc_15497_new_n4988_), .B(round_ctr_inc), .Y(_abc_15497_new_n4989_));
AND2X2 AND2X2_2113 ( .A(_abc_15497_new_n4989_), .B(_abc_15497_new_n4985_), .Y(_abc_15497_new_n4990_));
AND2X2 AND2X2_2114 ( .A(_abc_15497_new_n2010_), .B(a_reg_15_), .Y(_abc_15497_new_n4991_));
AND2X2 AND2X2_2115 ( .A(_abc_15497_new_n700_), .B(\digest[143] ), .Y(_abc_15497_new_n4992_));
AND2X2 AND2X2_2116 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n4992_), .Y(_abc_15497_new_n4993_));
AND2X2 AND2X2_2117 ( .A(_abc_15497_new_n5001_), .B(_abc_15497_new_n5000_), .Y(_abc_15497_new_n5002_));
AND2X2 AND2X2_2118 ( .A(_abc_15497_new_n4999_), .B(_abc_15497_new_n5002_), .Y(_abc_15497_new_n5003_));
AND2X2 AND2X2_2119 ( .A(_abc_15497_new_n4998_), .B(_abc_15497_new_n5003_), .Y(_abc_15497_new_n5004_));
AND2X2 AND2X2_212 ( .A(_abc_15497_new_n701_), .B(\digest[10] ), .Y(_abc_15497_new_n1148_));
AND2X2 AND2X2_2120 ( .A(_abc_15497_new_n5006_), .B(_abc_15497_new_n5004_), .Y(_abc_15497_new_n5007_));
AND2X2 AND2X2_2121 ( .A(_abc_15497_new_n4976_), .B(_abc_15497_new_n4968_), .Y(_abc_15497_new_n5009_));
AND2X2 AND2X2_2122 ( .A(_abc_15497_new_n4060_), .B(_abc_15497_new_n3784_), .Y(_abc_15497_new_n5010_));
AND2X2 AND2X2_2123 ( .A(_abc_15497_new_n4963_), .B(_abc_15497_new_n4959_), .Y(_abc_15497_new_n5012_));
AND2X2 AND2X2_2124 ( .A(d_reg_16_), .B(b_reg_16_), .Y(_abc_15497_new_n5015_));
AND2X2 AND2X2_2125 ( .A(_abc_15497_new_n5016_), .B(_abc_15497_new_n5014_), .Y(_abc_15497_new_n5017_));
AND2X2 AND2X2_2126 ( .A(_abc_15497_new_n5017_), .B(c_reg_16_), .Y(_abc_15497_new_n5018_));
AND2X2 AND2X2_2127 ( .A(_abc_15497_new_n5019_), .B(_abc_15497_new_n5020_), .Y(_abc_15497_new_n5021_));
AND2X2 AND2X2_2128 ( .A(_abc_15497_new_n3803_), .B(_abc_15497_new_n5021_), .Y(_abc_15497_new_n5022_));
AND2X2 AND2X2_2129 ( .A(_abc_15497_new_n5025_), .B(b_reg_16_), .Y(_abc_15497_new_n5026_));
AND2X2 AND2X2_213 ( .A(_abc_15497_new_n1143_), .B(_abc_15497_new_n1135_), .Y(_abc_15497_new_n1149_));
AND2X2 AND2X2_2130 ( .A(_abc_15497_new_n5014_), .B(c_reg_16_), .Y(_abc_15497_new_n5029_));
AND2X2 AND2X2_2131 ( .A(_abc_15497_new_n3774_), .B(_abc_15497_new_n5030_), .Y(_abc_15497_new_n5031_));
AND2X2 AND2X2_2132 ( .A(_abc_15497_new_n5032_), .B(_abc_15497_new_n5028_), .Y(_abc_15497_new_n5033_));
AND2X2 AND2X2_2133 ( .A(_abc_15497_new_n5023_), .B(_abc_15497_new_n5033_), .Y(_abc_15497_new_n5034_));
AND2X2 AND2X2_2134 ( .A(_abc_15497_new_n4956_), .B(_abc_15497_new_n4952_), .Y(_abc_15497_new_n5035_));
AND2X2 AND2X2_2135 ( .A(e_reg_16_), .B(a_reg_11_), .Y(_abc_15497_new_n5039_));
AND2X2 AND2X2_2136 ( .A(_abc_15497_new_n5040_), .B(_abc_15497_new_n5038_), .Y(_abc_15497_new_n5041_));
AND2X2 AND2X2_2137 ( .A(_abc_15497_new_n5042_), .B(_abc_15497_new_n5037_), .Y(_abc_15497_new_n5043_));
AND2X2 AND2X2_2138 ( .A(_abc_15497_new_n5041_), .B(w_16_), .Y(_abc_15497_new_n5044_));
AND2X2 AND2X2_2139 ( .A(_abc_15497_new_n5046_), .B(_abc_15497_new_n5036_), .Y(_abc_15497_new_n5047_));
AND2X2 AND2X2_214 ( .A(_abc_15497_new_n1139_), .B(_abc_15497_new_n1149_), .Y(_abc_15497_new_n1150_));
AND2X2 AND2X2_2140 ( .A(_abc_15497_new_n5045_), .B(_abc_15497_new_n5035_), .Y(_abc_15497_new_n5048_));
AND2X2 AND2X2_2141 ( .A(_abc_15497_new_n5034_), .B(_abc_15497_new_n5049_), .Y(_abc_15497_new_n5051_));
AND2X2 AND2X2_2142 ( .A(_abc_15497_new_n5052_), .B(_abc_15497_new_n5050_), .Y(_abc_15497_new_n5053_));
AND2X2 AND2X2_2143 ( .A(_abc_15497_new_n5013_), .B(_abc_15497_new_n5053_), .Y(_abc_15497_new_n5055_));
AND2X2 AND2X2_2144 ( .A(_abc_15497_new_n5056_), .B(_abc_15497_new_n5054_), .Y(_abc_15497_new_n5057_));
AND2X2 AND2X2_2145 ( .A(_abc_15497_new_n5057_), .B(_abc_15497_new_n5011_), .Y(_abc_15497_new_n5058_));
AND2X2 AND2X2_2146 ( .A(_abc_15497_new_n5059_), .B(_abc_15497_new_n5010_), .Y(_abc_15497_new_n5060_));
AND2X2 AND2X2_2147 ( .A(_abc_15497_new_n5061_), .B(_abc_15497_new_n5009_), .Y(_abc_15497_new_n5062_));
AND2X2 AND2X2_2148 ( .A(_abc_15497_new_n5008_), .B(_abc_15497_new_n5066_), .Y(_abc_15497_new_n5068_));
AND2X2 AND2X2_2149 ( .A(_abc_15497_new_n5069_), .B(round_ctr_inc), .Y(_abc_15497_new_n5070_));
AND2X2 AND2X2_215 ( .A(e_reg_10_), .B(\digest[10] ), .Y(_abc_15497_new_n1153_));
AND2X2 AND2X2_2150 ( .A(_abc_15497_new_n5070_), .B(_abc_15497_new_n5067_), .Y(_abc_15497_new_n5071_));
AND2X2 AND2X2_2151 ( .A(_abc_15497_new_n2010_), .B(a_reg_16_), .Y(_abc_15497_new_n5072_));
AND2X2 AND2X2_2152 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n2957_), .Y(_abc_15497_new_n5073_));
AND2X2 AND2X2_2153 ( .A(_abc_15497_new_n5069_), .B(_abc_15497_new_n5063_), .Y(_abc_15497_new_n5076_));
AND2X2 AND2X2_2154 ( .A(_abc_15497_new_n5078_), .B(_abc_15497_new_n5056_), .Y(_abc_15497_new_n5079_));
AND2X2 AND2X2_2155 ( .A(_abc_15497_new_n5050_), .B(_abc_15497_new_n5081_), .Y(_abc_15497_new_n5082_));
AND2X2 AND2X2_2156 ( .A(b_reg_17_), .B(c_reg_17_), .Y(_abc_15497_new_n5084_));
AND2X2 AND2X2_2157 ( .A(_abc_15497_new_n5085_), .B(_abc_15497_new_n5083_), .Y(_abc_15497_new_n5086_));
AND2X2 AND2X2_2158 ( .A(_abc_15497_new_n5086_), .B(d_reg_17_), .Y(_abc_15497_new_n5088_));
AND2X2 AND2X2_2159 ( .A(_abc_15497_new_n5089_), .B(_abc_15497_new_n5087_), .Y(_abc_15497_new_n5090_));
AND2X2 AND2X2_216 ( .A(_abc_15497_new_n1154_), .B(_abc_15497_new_n1152_), .Y(_abc_15497_new_n1155_));
AND2X2 AND2X2_2160 ( .A(_abc_15497_new_n3803_), .B(_abc_15497_new_n5090_), .Y(_abc_15497_new_n5091_));
AND2X2 AND2X2_2161 ( .A(_abc_15497_new_n5094_), .B(_abc_15497_new_n5085_), .Y(_abc_15497_new_n5095_));
AND2X2 AND2X2_2162 ( .A(_abc_15497_new_n5085_), .B(_abc_15497_new_n5093_), .Y(_abc_15497_new_n5098_));
AND2X2 AND2X2_2163 ( .A(_abc_15497_new_n5100_), .B(_abc_15497_new_n5096_), .Y(_abc_15497_new_n5101_));
AND2X2 AND2X2_2164 ( .A(_abc_15497_new_n5092_), .B(_abc_15497_new_n5101_), .Y(_abc_15497_new_n5102_));
AND2X2 AND2X2_2165 ( .A(e_reg_17_), .B(a_reg_12_), .Y(_abc_15497_new_n5107_));
AND2X2 AND2X2_2166 ( .A(_abc_15497_new_n5108_), .B(_abc_15497_new_n5106_), .Y(_abc_15497_new_n5109_));
AND2X2 AND2X2_2167 ( .A(_abc_15497_new_n5110_), .B(_abc_15497_new_n5105_), .Y(_abc_15497_new_n5111_));
AND2X2 AND2X2_2168 ( .A(_abc_15497_new_n5109_), .B(w_17_), .Y(_abc_15497_new_n5112_));
AND2X2 AND2X2_2169 ( .A(_abc_15497_new_n5114_), .B(_abc_15497_new_n5104_), .Y(_abc_15497_new_n5115_));
AND2X2 AND2X2_217 ( .A(_abc_15497_new_n1151_), .B(_abc_15497_new_n1155_), .Y(_abc_15497_new_n1157_));
AND2X2 AND2X2_2170 ( .A(_abc_15497_new_n5116_), .B(_abc_15497_new_n5117_), .Y(_abc_15497_new_n5118_));
AND2X2 AND2X2_2171 ( .A(_abc_15497_new_n5103_), .B(_abc_15497_new_n5118_), .Y(_abc_15497_new_n5119_));
AND2X2 AND2X2_2172 ( .A(_abc_15497_new_n5120_), .B(_abc_15497_new_n5121_), .Y(_abc_15497_new_n5122_));
AND2X2 AND2X2_2173 ( .A(_abc_15497_new_n5123_), .B(_abc_15497_new_n5082_), .Y(_abc_15497_new_n5124_));
AND2X2 AND2X2_2174 ( .A(_abc_15497_new_n5127_), .B(_abc_15497_new_n4059_), .Y(_abc_15497_new_n5130_));
AND2X2 AND2X2_2175 ( .A(_abc_15497_new_n5132_), .B(_abc_15497_new_n5080_), .Y(_abc_15497_new_n5133_));
AND2X2 AND2X2_2176 ( .A(_abc_15497_new_n5131_), .B(_abc_15497_new_n5079_), .Y(_abc_15497_new_n5134_));
AND2X2 AND2X2_2177 ( .A(_abc_15497_new_n5138_), .B(round_ctr_inc), .Y(_abc_15497_new_n5139_));
AND2X2 AND2X2_2178 ( .A(_abc_15497_new_n5139_), .B(_abc_15497_new_n5137_), .Y(_abc_15497_new_n5140_));
AND2X2 AND2X2_2179 ( .A(_abc_15497_new_n2010_), .B(a_reg_17_), .Y(_abc_15497_new_n5141_));
AND2X2 AND2X2_218 ( .A(_abc_15497_new_n1158_), .B(_abc_15497_new_n1156_), .Y(_abc_15497_new_n1159_));
AND2X2 AND2X2_2180 ( .A(_abc_15497_new_n700_), .B(\digest[145] ), .Y(_abc_15497_new_n5142_));
AND2X2 AND2X2_2181 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n5142_), .Y(_abc_15497_new_n5143_));
AND2X2 AND2X2_2182 ( .A(_abc_15497_new_n5068_), .B(_abc_15497_new_n5136_), .Y(_abc_15497_new_n5146_));
AND2X2 AND2X2_2183 ( .A(_abc_15497_new_n5147_), .B(_abc_15497_new_n5148_), .Y(_abc_15497_new_n5149_));
AND2X2 AND2X2_2184 ( .A(_abc_15497_new_n5128_), .B(_abc_15497_new_n5125_), .Y(_abc_15497_new_n5152_));
AND2X2 AND2X2_2185 ( .A(_abc_15497_new_n5120_), .B(_abc_15497_new_n5116_), .Y(_abc_15497_new_n5154_));
AND2X2 AND2X2_2186 ( .A(d_reg_18_), .B(b_reg_18_), .Y(_abc_15497_new_n5157_));
AND2X2 AND2X2_2187 ( .A(_abc_15497_new_n5158_), .B(_abc_15497_new_n5156_), .Y(_abc_15497_new_n5159_));
AND2X2 AND2X2_2188 ( .A(_abc_15497_new_n5159_), .B(c_reg_18_), .Y(_abc_15497_new_n5160_));
AND2X2 AND2X2_2189 ( .A(_abc_15497_new_n5161_), .B(_abc_15497_new_n5162_), .Y(_abc_15497_new_n5163_));
AND2X2 AND2X2_219 ( .A(_abc_15497_new_n1159_), .B(digest_update), .Y(_abc_15497_new_n1160_));
AND2X2 AND2X2_2190 ( .A(_abc_15497_new_n3803_), .B(_abc_15497_new_n5163_), .Y(_abc_15497_new_n5164_));
AND2X2 AND2X2_2191 ( .A(_abc_15497_new_n5167_), .B(b_reg_18_), .Y(_abc_15497_new_n5168_));
AND2X2 AND2X2_2192 ( .A(_abc_15497_new_n5156_), .B(c_reg_18_), .Y(_abc_15497_new_n5171_));
AND2X2 AND2X2_2193 ( .A(_abc_15497_new_n3774_), .B(_abc_15497_new_n5172_), .Y(_abc_15497_new_n5173_));
AND2X2 AND2X2_2194 ( .A(_abc_15497_new_n5174_), .B(_abc_15497_new_n5170_), .Y(_abc_15497_new_n5175_));
AND2X2 AND2X2_2195 ( .A(_abc_15497_new_n5165_), .B(_abc_15497_new_n5175_), .Y(_abc_15497_new_n5176_));
AND2X2 AND2X2_2196 ( .A(e_reg_18_), .B(a_reg_13_), .Y(_abc_15497_new_n5180_));
AND2X2 AND2X2_2197 ( .A(_abc_15497_new_n5181_), .B(_abc_15497_new_n5179_), .Y(_abc_15497_new_n5182_));
AND2X2 AND2X2_2198 ( .A(_abc_15497_new_n5183_), .B(_abc_15497_new_n5178_), .Y(_abc_15497_new_n5184_));
AND2X2 AND2X2_2199 ( .A(_abc_15497_new_n5182_), .B(w_18_), .Y(_abc_15497_new_n5185_));
AND2X2 AND2X2_22 ( .A(_abc_15497_new_n734_), .B(_abc_15497_new_n738_), .Y(_abc_15497_new_n739_));
AND2X2 AND2X2_220 ( .A(_abc_15497_new_n701_), .B(\digest[11] ), .Y(_abc_15497_new_n1162_));
AND2X2 AND2X2_2200 ( .A(_abc_15497_new_n5187_), .B(_abc_15497_new_n5177_), .Y(_abc_15497_new_n5188_));
AND2X2 AND2X2_2201 ( .A(_abc_15497_new_n5189_), .B(_abc_15497_new_n5190_), .Y(_abc_15497_new_n5191_));
AND2X2 AND2X2_2202 ( .A(_abc_15497_new_n5192_), .B(_abc_15497_new_n5176_), .Y(_abc_15497_new_n5193_));
AND2X2 AND2X2_2203 ( .A(_abc_15497_new_n5194_), .B(_abc_15497_new_n5191_), .Y(_abc_15497_new_n5195_));
AND2X2 AND2X2_2204 ( .A(_abc_15497_new_n5155_), .B(_abc_15497_new_n5197_), .Y(_abc_15497_new_n5198_));
AND2X2 AND2X2_2205 ( .A(_abc_15497_new_n5154_), .B(_abc_15497_new_n5196_), .Y(_abc_15497_new_n5199_));
AND2X2 AND2X2_2206 ( .A(_abc_15497_new_n5153_), .B(_abc_15497_new_n5201_), .Y(_abc_15497_new_n5202_));
AND2X2 AND2X2_2207 ( .A(_abc_15497_new_n5152_), .B(_abc_15497_new_n5200_), .Y(_abc_15497_new_n5203_));
AND2X2 AND2X2_2208 ( .A(_abc_15497_new_n5151_), .B(_abc_15497_new_n5205_), .Y(_abc_15497_new_n5207_));
AND2X2 AND2X2_2209 ( .A(_abc_15497_new_n5208_), .B(round_ctr_inc), .Y(_abc_15497_new_n5209_));
AND2X2 AND2X2_221 ( .A(_abc_15497_new_n1158_), .B(_abc_15497_new_n1154_), .Y(_abc_15497_new_n1163_));
AND2X2 AND2X2_2210 ( .A(_abc_15497_new_n5209_), .B(_abc_15497_new_n5206_), .Y(_abc_15497_new_n5210_));
AND2X2 AND2X2_2211 ( .A(_abc_15497_new_n2010_), .B(a_reg_18_), .Y(_abc_15497_new_n5211_));
AND2X2 AND2X2_2212 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n2988_), .Y(_abc_15497_new_n5212_));
AND2X2 AND2X2_2213 ( .A(_abc_15497_new_n5208_), .B(_abc_15497_new_n5215_), .Y(_abc_15497_new_n5216_));
AND2X2 AND2X2_2214 ( .A(d_reg_19_), .B(b_reg_19_), .Y(_abc_15497_new_n5220_));
AND2X2 AND2X2_2215 ( .A(_abc_15497_new_n5221_), .B(_abc_15497_new_n5219_), .Y(_abc_15497_new_n5222_));
AND2X2 AND2X2_2216 ( .A(_abc_15497_new_n5222_), .B(c_reg_19_), .Y(_abc_15497_new_n5223_));
AND2X2 AND2X2_2217 ( .A(_abc_15497_new_n5224_), .B(_abc_15497_new_n5225_), .Y(_abc_15497_new_n5226_));
AND2X2 AND2X2_2218 ( .A(_abc_15497_new_n3803_), .B(_abc_15497_new_n5226_), .Y(_abc_15497_new_n5227_));
AND2X2 AND2X2_2219 ( .A(_abc_15497_new_n5230_), .B(b_reg_19_), .Y(_abc_15497_new_n5231_));
AND2X2 AND2X2_222 ( .A(e_reg_11_), .B(\digest[11] ), .Y(_abc_15497_new_n1166_));
AND2X2 AND2X2_2220 ( .A(_abc_15497_new_n5219_), .B(c_reg_19_), .Y(_abc_15497_new_n5234_));
AND2X2 AND2X2_2221 ( .A(_abc_15497_new_n3774_), .B(_abc_15497_new_n5235_), .Y(_abc_15497_new_n5236_));
AND2X2 AND2X2_2222 ( .A(_abc_15497_new_n5237_), .B(_abc_15497_new_n5233_), .Y(_abc_15497_new_n5238_));
AND2X2 AND2X2_2223 ( .A(_abc_15497_new_n5228_), .B(_abc_15497_new_n5238_), .Y(_abc_15497_new_n5239_));
AND2X2 AND2X2_2224 ( .A(e_reg_19_), .B(a_reg_14_), .Y(_abc_15497_new_n5244_));
AND2X2 AND2X2_2225 ( .A(_abc_15497_new_n5245_), .B(_abc_15497_new_n5243_), .Y(_abc_15497_new_n5246_));
AND2X2 AND2X2_2226 ( .A(_abc_15497_new_n5247_), .B(_abc_15497_new_n5242_), .Y(_abc_15497_new_n5248_));
AND2X2 AND2X2_2227 ( .A(_abc_15497_new_n5246_), .B(w_19_), .Y(_abc_15497_new_n5249_));
AND2X2 AND2X2_2228 ( .A(_abc_15497_new_n5251_), .B(_abc_15497_new_n5241_), .Y(_abc_15497_new_n5252_));
AND2X2 AND2X2_2229 ( .A(_abc_15497_new_n5253_), .B(_abc_15497_new_n5254_), .Y(_abc_15497_new_n5255_));
AND2X2 AND2X2_223 ( .A(_abc_15497_new_n1167_), .B(_abc_15497_new_n1165_), .Y(_abc_15497_new_n1168_));
AND2X2 AND2X2_2230 ( .A(_abc_15497_new_n5240_), .B(_abc_15497_new_n5255_), .Y(_abc_15497_new_n5256_));
AND2X2 AND2X2_2231 ( .A(_abc_15497_new_n5257_), .B(_abc_15497_new_n5258_), .Y(_abc_15497_new_n5259_));
AND2X2 AND2X2_2232 ( .A(_abc_15497_new_n5260_), .B(_abc_15497_new_n5218_), .Y(_abc_15497_new_n5261_));
AND2X2 AND2X2_2233 ( .A(_abc_15497_new_n5259_), .B(_abc_15497_new_n5217_), .Y(_abc_15497_new_n5262_));
AND2X2 AND2X2_2234 ( .A(_abc_15497_new_n5264_), .B(_abc_15497_new_n5011_), .Y(_abc_15497_new_n5265_));
AND2X2 AND2X2_2235 ( .A(_abc_15497_new_n5263_), .B(_abc_15497_new_n5010_), .Y(_abc_15497_new_n5266_));
AND2X2 AND2X2_2236 ( .A(_abc_15497_new_n5268_), .B(_abc_15497_new_n5198_), .Y(_abc_15497_new_n5269_));
AND2X2 AND2X2_2237 ( .A(_abc_15497_new_n5267_), .B(_abc_15497_new_n5270_), .Y(_abc_15497_new_n5271_));
AND2X2 AND2X2_2238 ( .A(_abc_15497_new_n5276_), .B(round_ctr_inc), .Y(_abc_15497_new_n5277_));
AND2X2 AND2X2_2239 ( .A(_abc_15497_new_n5277_), .B(_abc_15497_new_n5273_), .Y(_abc_15497_new_n5278_));
AND2X2 AND2X2_224 ( .A(_abc_15497_new_n1171_), .B(digest_update), .Y(_abc_15497_new_n1172_));
AND2X2 AND2X2_2240 ( .A(_abc_15497_new_n2010_), .B(a_reg_19_), .Y(_abc_15497_new_n5279_));
AND2X2 AND2X2_2241 ( .A(_abc_15497_new_n700_), .B(\digest[147] ), .Y(_abc_15497_new_n5280_));
AND2X2 AND2X2_2242 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n5280_), .Y(_abc_15497_new_n5281_));
AND2X2 AND2X2_2243 ( .A(_abc_15497_new_n5287_), .B(_abc_15497_new_n5286_), .Y(_abc_15497_new_n5288_));
AND2X2 AND2X2_2244 ( .A(_abc_15497_new_n5285_), .B(_abc_15497_new_n5289_), .Y(_abc_15497_new_n5290_));
AND2X2 AND2X2_2245 ( .A(_abc_15497_new_n5293_), .B(_abc_15497_new_n5290_), .Y(_abc_15497_new_n5294_));
AND2X2 AND2X2_2246 ( .A(_abc_15497_new_n5297_), .B(_abc_15497_new_n5296_), .Y(_abc_15497_new_n5298_));
AND2X2 AND2X2_2247 ( .A(d_reg_20_), .B(b_reg_20_), .Y(_abc_15497_new_n5303_));
AND2X2 AND2X2_2248 ( .A(_abc_15497_new_n5304_), .B(_abc_15497_new_n5302_), .Y(_abc_15497_new_n5305_));
AND2X2 AND2X2_2249 ( .A(_abc_15497_new_n5305_), .B(c_reg_20_), .Y(_abc_15497_new_n5306_));
AND2X2 AND2X2_225 ( .A(_abc_15497_new_n1172_), .B(_abc_15497_new_n1169_), .Y(_abc_15497_new_n1173_));
AND2X2 AND2X2_2250 ( .A(_abc_15497_new_n5307_), .B(_abc_15497_new_n5308_), .Y(_abc_15497_new_n5309_));
AND2X2 AND2X2_2251 ( .A(_abc_15497_new_n3803_), .B(_abc_15497_new_n5309_), .Y(_abc_15497_new_n5310_));
AND2X2 AND2X2_2252 ( .A(_abc_15497_new_n5313_), .B(b_reg_20_), .Y(_abc_15497_new_n5314_));
AND2X2 AND2X2_2253 ( .A(_abc_15497_new_n5302_), .B(c_reg_20_), .Y(_abc_15497_new_n5317_));
AND2X2 AND2X2_2254 ( .A(_abc_15497_new_n3774_), .B(_abc_15497_new_n5318_), .Y(_abc_15497_new_n5319_));
AND2X2 AND2X2_2255 ( .A(_abc_15497_new_n5320_), .B(_abc_15497_new_n5316_), .Y(_abc_15497_new_n5321_));
AND2X2 AND2X2_2256 ( .A(_abc_15497_new_n5311_), .B(_abc_15497_new_n5321_), .Y(_abc_15497_new_n5322_));
AND2X2 AND2X2_2257 ( .A(e_reg_20_), .B(a_reg_15_), .Y(_abc_15497_new_n5327_));
AND2X2 AND2X2_2258 ( .A(_abc_15497_new_n5328_), .B(_abc_15497_new_n5326_), .Y(_abc_15497_new_n5329_));
AND2X2 AND2X2_2259 ( .A(_abc_15497_new_n5330_), .B(_abc_15497_new_n5325_), .Y(_abc_15497_new_n5331_));
AND2X2 AND2X2_226 ( .A(_abc_15497_new_n701_), .B(\digest[12] ), .Y(_abc_15497_new_n1175_));
AND2X2 AND2X2_2260 ( .A(_abc_15497_new_n5329_), .B(w_20_), .Y(_abc_15497_new_n5332_));
AND2X2 AND2X2_2261 ( .A(_abc_15497_new_n5334_), .B(_abc_15497_new_n5324_), .Y(_abc_15497_new_n5335_));
AND2X2 AND2X2_2262 ( .A(_abc_15497_new_n5336_), .B(_abc_15497_new_n5337_), .Y(_abc_15497_new_n5338_));
AND2X2 AND2X2_2263 ( .A(_abc_15497_new_n5323_), .B(_abc_15497_new_n5338_), .Y(_abc_15497_new_n5339_));
AND2X2 AND2X2_2264 ( .A(_abc_15497_new_n5340_), .B(_abc_15497_new_n5341_), .Y(_abc_15497_new_n5342_));
AND2X2 AND2X2_2265 ( .A(_abc_15497_new_n5343_), .B(_abc_15497_new_n5301_), .Y(_abc_15497_new_n5344_));
AND2X2 AND2X2_2266 ( .A(_abc_15497_new_n5342_), .B(_abc_15497_new_n5300_), .Y(_abc_15497_new_n5345_));
AND2X2 AND2X2_2267 ( .A(_abc_15497_new_n5346_), .B(_abc_15497_new_n5010_), .Y(_abc_15497_new_n5349_));
AND2X2 AND2X2_2268 ( .A(_abc_15497_new_n5299_), .B(_abc_15497_new_n5351_), .Y(_abc_15497_new_n5352_));
AND2X2 AND2X2_2269 ( .A(_abc_15497_new_n5298_), .B(_abc_15497_new_n5350_), .Y(_abc_15497_new_n5353_));
AND2X2 AND2X2_227 ( .A(_abc_15497_new_n1155_), .B(_abc_15497_new_n1168_), .Y(_abc_15497_new_n1176_));
AND2X2 AND2X2_2270 ( .A(_abc_15497_new_n5357_), .B(round_ctr_inc), .Y(_abc_15497_new_n5358_));
AND2X2 AND2X2_2271 ( .A(_abc_15497_new_n5358_), .B(_abc_15497_new_n5356_), .Y(_abc_15497_new_n5359_));
AND2X2 AND2X2_2272 ( .A(_abc_15497_new_n2010_), .B(a_reg_20_), .Y(_abc_15497_new_n5360_));
AND2X2 AND2X2_2273 ( .A(_abc_15497_new_n700_), .B(\digest[148] ), .Y(_abc_15497_new_n5361_));
AND2X2 AND2X2_2274 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n5361_), .Y(_abc_15497_new_n5362_));
AND2X2 AND2X2_2275 ( .A(_abc_15497_new_n5357_), .B(_abc_15497_new_n5365_), .Y(_abc_15497_new_n5366_));
AND2X2 AND2X2_2276 ( .A(d_reg_21_), .B(b_reg_21_), .Y(_abc_15497_new_n5372_));
AND2X2 AND2X2_2277 ( .A(_abc_15497_new_n5373_), .B(_abc_15497_new_n5371_), .Y(_abc_15497_new_n5374_));
AND2X2 AND2X2_2278 ( .A(_abc_15497_new_n5374_), .B(c_reg_21_), .Y(_abc_15497_new_n5375_));
AND2X2 AND2X2_2279 ( .A(_abc_15497_new_n5376_), .B(_abc_15497_new_n5377_), .Y(_abc_15497_new_n5378_));
AND2X2 AND2X2_228 ( .A(_abc_15497_new_n1165_), .B(_abc_15497_new_n1153_), .Y(_abc_15497_new_n1179_));
AND2X2 AND2X2_2280 ( .A(_abc_15497_new_n3803_), .B(_abc_15497_new_n5378_), .Y(_abc_15497_new_n5379_));
AND2X2 AND2X2_2281 ( .A(_abc_15497_new_n5382_), .B(b_reg_21_), .Y(_abc_15497_new_n5383_));
AND2X2 AND2X2_2282 ( .A(_abc_15497_new_n5371_), .B(c_reg_21_), .Y(_abc_15497_new_n5386_));
AND2X2 AND2X2_2283 ( .A(_abc_15497_new_n3774_), .B(_abc_15497_new_n5387_), .Y(_abc_15497_new_n5388_));
AND2X2 AND2X2_2284 ( .A(_abc_15497_new_n5389_), .B(_abc_15497_new_n5385_), .Y(_abc_15497_new_n5390_));
AND2X2 AND2X2_2285 ( .A(_abc_15497_new_n5380_), .B(_abc_15497_new_n5390_), .Y(_abc_15497_new_n5391_));
AND2X2 AND2X2_2286 ( .A(e_reg_21_), .B(a_reg_16_), .Y(_abc_15497_new_n5396_));
AND2X2 AND2X2_2287 ( .A(_abc_15497_new_n5397_), .B(_abc_15497_new_n5395_), .Y(_abc_15497_new_n5398_));
AND2X2 AND2X2_2288 ( .A(_abc_15497_new_n5399_), .B(_abc_15497_new_n5394_), .Y(_abc_15497_new_n5400_));
AND2X2 AND2X2_2289 ( .A(_abc_15497_new_n5398_), .B(w_21_), .Y(_abc_15497_new_n5401_));
AND2X2 AND2X2_229 ( .A(_abc_15497_new_n1178_), .B(_abc_15497_new_n1181_), .Y(_abc_15497_new_n1182_));
AND2X2 AND2X2_2290 ( .A(_abc_15497_new_n5403_), .B(_abc_15497_new_n5393_), .Y(_abc_15497_new_n5404_));
AND2X2 AND2X2_2291 ( .A(_abc_15497_new_n5405_), .B(_abc_15497_new_n5406_), .Y(_abc_15497_new_n5407_));
AND2X2 AND2X2_2292 ( .A(_abc_15497_new_n5392_), .B(_abc_15497_new_n5407_), .Y(_abc_15497_new_n5408_));
AND2X2 AND2X2_2293 ( .A(_abc_15497_new_n5409_), .B(_abc_15497_new_n5410_), .Y(_abc_15497_new_n5411_));
AND2X2 AND2X2_2294 ( .A(_abc_15497_new_n5412_), .B(_abc_15497_new_n5370_), .Y(_abc_15497_new_n5413_));
AND2X2 AND2X2_2295 ( .A(_abc_15497_new_n5411_), .B(_abc_15497_new_n5369_), .Y(_abc_15497_new_n5414_));
AND2X2 AND2X2_2296 ( .A(_abc_15497_new_n5416_), .B(_abc_15497_new_n3783_), .Y(_abc_15497_new_n5417_));
AND2X2 AND2X2_2297 ( .A(_abc_15497_new_n5415_), .B(_abc_15497_new_n3773_), .Y(_abc_15497_new_n5418_));
AND2X2 AND2X2_2298 ( .A(_abc_15497_new_n5420_), .B(_abc_15497_new_n5368_), .Y(_abc_15497_new_n5421_));
AND2X2 AND2X2_2299 ( .A(_abc_15497_new_n5422_), .B(_abc_15497_new_n5419_), .Y(_abc_15497_new_n5423_));
AND2X2 AND2X2_23 ( .A(c_reg_17_), .B(\digest[81] ), .Y(_abc_15497_new_n740_));
AND2X2 AND2X2_230 ( .A(_abc_15497_new_n1137_), .B(_abc_15497_new_n1176_), .Y(_abc_15497_new_n1184_));
AND2X2 AND2X2_2300 ( .A(_abc_15497_new_n5427_), .B(round_ctr_inc), .Y(_abc_15497_new_n5428_));
AND2X2 AND2X2_2301 ( .A(_abc_15497_new_n5428_), .B(_abc_15497_new_n5426_), .Y(_abc_15497_new_n5429_));
AND2X2 AND2X2_2302 ( .A(_abc_15497_new_n2010_), .B(a_reg_21_), .Y(_abc_15497_new_n5430_));
AND2X2 AND2X2_2303 ( .A(_abc_15497_new_n700_), .B(\digest[149] ), .Y(_abc_15497_new_n5431_));
AND2X2 AND2X2_2304 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n5431_), .Y(_abc_15497_new_n5432_));
AND2X2 AND2X2_2305 ( .A(_abc_15497_new_n5438_), .B(_abc_15497_new_n5437_), .Y(_abc_15497_new_n5439_));
AND2X2 AND2X2_2306 ( .A(_abc_15497_new_n5436_), .B(_abc_15497_new_n5439_), .Y(_abc_15497_new_n5440_));
AND2X2 AND2X2_2307 ( .A(_abc_15497_new_n5443_), .B(_abc_15497_new_n5442_), .Y(_abc_15497_new_n5444_));
AND2X2 AND2X2_2308 ( .A(_abc_15497_new_n5409_), .B(_abc_15497_new_n5405_), .Y(_abc_15497_new_n5446_));
AND2X2 AND2X2_2309 ( .A(d_reg_22_), .B(b_reg_22_), .Y(_abc_15497_new_n5448_));
AND2X2 AND2X2_231 ( .A(_abc_15497_new_n1123_), .B(_abc_15497_new_n1184_), .Y(_abc_15497_new_n1185_));
AND2X2 AND2X2_2310 ( .A(_abc_15497_new_n5449_), .B(_abc_15497_new_n5447_), .Y(_abc_15497_new_n5450_));
AND2X2 AND2X2_2311 ( .A(_abc_15497_new_n5450_), .B(c_reg_22_), .Y(_abc_15497_new_n5451_));
AND2X2 AND2X2_2312 ( .A(_abc_15497_new_n5452_), .B(_abc_15497_new_n5453_), .Y(_abc_15497_new_n5454_));
AND2X2 AND2X2_2313 ( .A(_abc_15497_new_n3803_), .B(_abc_15497_new_n5454_), .Y(_abc_15497_new_n5455_));
AND2X2 AND2X2_2314 ( .A(_abc_15497_new_n5458_), .B(b_reg_22_), .Y(_abc_15497_new_n5459_));
AND2X2 AND2X2_2315 ( .A(_abc_15497_new_n5447_), .B(c_reg_22_), .Y(_abc_15497_new_n5462_));
AND2X2 AND2X2_2316 ( .A(_abc_15497_new_n3774_), .B(_abc_15497_new_n5463_), .Y(_abc_15497_new_n5464_));
AND2X2 AND2X2_2317 ( .A(_abc_15497_new_n5465_), .B(_abc_15497_new_n5461_), .Y(_abc_15497_new_n5466_));
AND2X2 AND2X2_2318 ( .A(_abc_15497_new_n5456_), .B(_abc_15497_new_n5466_), .Y(_abc_15497_new_n5467_));
AND2X2 AND2X2_2319 ( .A(e_reg_22_), .B(a_reg_17_), .Y(_abc_15497_new_n5472_));
AND2X2 AND2X2_232 ( .A(e_reg_12_), .B(\digest[12] ), .Y(_abc_15497_new_n1188_));
AND2X2 AND2X2_2320 ( .A(_abc_15497_new_n5473_), .B(_abc_15497_new_n5471_), .Y(_abc_15497_new_n5474_));
AND2X2 AND2X2_2321 ( .A(_abc_15497_new_n5475_), .B(_abc_15497_new_n5470_), .Y(_abc_15497_new_n5476_));
AND2X2 AND2X2_2322 ( .A(_abc_15497_new_n5474_), .B(w_22_), .Y(_abc_15497_new_n5477_));
AND2X2 AND2X2_2323 ( .A(_abc_15497_new_n5479_), .B(_abc_15497_new_n5469_), .Y(_abc_15497_new_n5480_));
AND2X2 AND2X2_2324 ( .A(_abc_15497_new_n5481_), .B(_abc_15497_new_n5482_), .Y(_abc_15497_new_n5483_));
AND2X2 AND2X2_2325 ( .A(_abc_15497_new_n5468_), .B(_abc_15497_new_n5483_), .Y(_abc_15497_new_n5484_));
AND2X2 AND2X2_2326 ( .A(_abc_15497_new_n5485_), .B(_abc_15497_new_n5486_), .Y(_abc_15497_new_n5487_));
AND2X2 AND2X2_2327 ( .A(_abc_15497_new_n5488_), .B(_abc_15497_new_n5446_), .Y(_abc_15497_new_n5489_));
AND2X2 AND2X2_2328 ( .A(_abc_15497_new_n5493_), .B(_abc_15497_new_n3803_), .Y(_abc_15497_new_n5494_));
AND2X2 AND2X2_2329 ( .A(_abc_15497_new_n5492_), .B(_abc_15497_new_n3775_), .Y(_abc_15497_new_n5495_));
AND2X2 AND2X2_233 ( .A(_abc_15497_new_n1189_), .B(_abc_15497_new_n1187_), .Y(_abc_15497_new_n1190_));
AND2X2 AND2X2_2330 ( .A(_abc_15497_new_n5497_), .B(_abc_15497_new_n5445_), .Y(_abc_15497_new_n5498_));
AND2X2 AND2X2_2331 ( .A(_abc_15497_new_n5496_), .B(_abc_15497_new_n5444_), .Y(_abc_15497_new_n5499_));
AND2X2 AND2X2_2332 ( .A(_abc_15497_new_n5503_), .B(round_ctr_inc), .Y(_abc_15497_new_n5504_));
AND2X2 AND2X2_2333 ( .A(_abc_15497_new_n5504_), .B(_abc_15497_new_n5502_), .Y(_abc_15497_new_n5505_));
AND2X2 AND2X2_2334 ( .A(_abc_15497_new_n2010_), .B(a_reg_22_), .Y(_abc_15497_new_n5506_));
AND2X2 AND2X2_2335 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3050_), .Y(_abc_15497_new_n5507_));
AND2X2 AND2X2_2336 ( .A(_abc_15497_new_n5503_), .B(_abc_15497_new_n5510_), .Y(_abc_15497_new_n5511_));
AND2X2 AND2X2_2337 ( .A(_abc_15497_new_n5485_), .B(_abc_15497_new_n5481_), .Y(_abc_15497_new_n5514_));
AND2X2 AND2X2_2338 ( .A(b_reg_23_), .B(c_reg_23_), .Y(_abc_15497_new_n5516_));
AND2X2 AND2X2_2339 ( .A(_abc_15497_new_n5517_), .B(_abc_15497_new_n5515_), .Y(_abc_15497_new_n5518_));
AND2X2 AND2X2_234 ( .A(_abc_15497_new_n1186_), .B(_abc_15497_new_n1190_), .Y(_abc_15497_new_n1192_));
AND2X2 AND2X2_2340 ( .A(_abc_15497_new_n5518_), .B(d_reg_23_), .Y(_abc_15497_new_n5520_));
AND2X2 AND2X2_2341 ( .A(_abc_15497_new_n5521_), .B(_abc_15497_new_n5519_), .Y(_abc_15497_new_n5522_));
AND2X2 AND2X2_2342 ( .A(_abc_15497_new_n3803_), .B(_abc_15497_new_n5522_), .Y(_abc_15497_new_n5523_));
AND2X2 AND2X2_2343 ( .A(_abc_15497_new_n5526_), .B(_abc_15497_new_n5517_), .Y(_abc_15497_new_n5527_));
AND2X2 AND2X2_2344 ( .A(_abc_15497_new_n5517_), .B(_abc_15497_new_n5525_), .Y(_abc_15497_new_n5530_));
AND2X2 AND2X2_2345 ( .A(_abc_15497_new_n5532_), .B(_abc_15497_new_n5528_), .Y(_abc_15497_new_n5533_));
AND2X2 AND2X2_2346 ( .A(_abc_15497_new_n5524_), .B(_abc_15497_new_n5533_), .Y(_abc_15497_new_n5534_));
AND2X2 AND2X2_2347 ( .A(e_reg_23_), .B(a_reg_18_), .Y(_abc_15497_new_n5539_));
AND2X2 AND2X2_2348 ( .A(_abc_15497_new_n5540_), .B(_abc_15497_new_n5538_), .Y(_abc_15497_new_n5541_));
AND2X2 AND2X2_2349 ( .A(_abc_15497_new_n5542_), .B(_abc_15497_new_n5537_), .Y(_abc_15497_new_n5543_));
AND2X2 AND2X2_235 ( .A(_abc_15497_new_n1193_), .B(_abc_15497_new_n1191_), .Y(_abc_15497_new_n1194_));
AND2X2 AND2X2_2350 ( .A(_abc_15497_new_n5541_), .B(w_23_), .Y(_abc_15497_new_n5544_));
AND2X2 AND2X2_2351 ( .A(_abc_15497_new_n5546_), .B(_abc_15497_new_n5536_), .Y(_abc_15497_new_n5547_));
AND2X2 AND2X2_2352 ( .A(_abc_15497_new_n5548_), .B(_abc_15497_new_n5549_), .Y(_abc_15497_new_n5550_));
AND2X2 AND2X2_2353 ( .A(_abc_15497_new_n5535_), .B(_abc_15497_new_n5550_), .Y(_abc_15497_new_n5551_));
AND2X2 AND2X2_2354 ( .A(_abc_15497_new_n5552_), .B(_abc_15497_new_n5553_), .Y(_abc_15497_new_n5554_));
AND2X2 AND2X2_2355 ( .A(_abc_15497_new_n5555_), .B(_abc_15497_new_n5514_), .Y(_abc_15497_new_n5556_));
AND2X2 AND2X2_2356 ( .A(_abc_15497_new_n5557_), .B(_abc_15497_new_n5558_), .Y(_abc_15497_new_n5559_));
AND2X2 AND2X2_2357 ( .A(_abc_15497_new_n5559_), .B(_abc_15497_new_n3744_), .Y(_abc_15497_new_n5560_));
AND2X2 AND2X2_2358 ( .A(_abc_15497_new_n5561_), .B(_abc_15497_new_n5562_), .Y(_abc_15497_new_n5563_));
AND2X2 AND2X2_2359 ( .A(_abc_15497_new_n5513_), .B(_abc_15497_new_n5563_), .Y(_abc_15497_new_n5564_));
AND2X2 AND2X2_236 ( .A(_abc_15497_new_n1194_), .B(digest_update), .Y(_abc_15497_new_n1195_));
AND2X2 AND2X2_2360 ( .A(_abc_15497_new_n5565_), .B(_abc_15497_new_n5566_), .Y(_abc_15497_new_n5567_));
AND2X2 AND2X2_2361 ( .A(_abc_15497_new_n5571_), .B(round_ctr_inc), .Y(_abc_15497_new_n5572_));
AND2X2 AND2X2_2362 ( .A(_abc_15497_new_n5572_), .B(_abc_15497_new_n5570_), .Y(_abc_15497_new_n5573_));
AND2X2 AND2X2_2363 ( .A(_abc_15497_new_n2010_), .B(a_reg_23_), .Y(_abc_15497_new_n5574_));
AND2X2 AND2X2_2364 ( .A(_abc_15497_new_n700_), .B(\digest[151] ), .Y(_abc_15497_new_n5575_));
AND2X2 AND2X2_2365 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n5575_), .Y(_abc_15497_new_n5576_));
AND2X2 AND2X2_2366 ( .A(_abc_15497_new_n5584_), .B(_abc_15497_new_n5583_), .Y(_abc_15497_new_n5585_));
AND2X2 AND2X2_2367 ( .A(_abc_15497_new_n5582_), .B(_abc_15497_new_n5585_), .Y(_abc_15497_new_n5586_));
AND2X2 AND2X2_2368 ( .A(_abc_15497_new_n5581_), .B(_abc_15497_new_n5586_), .Y(_abc_15497_new_n5587_));
AND2X2 AND2X2_2369 ( .A(_abc_15497_new_n5589_), .B(_abc_15497_new_n5587_), .Y(_abc_15497_new_n5590_));
AND2X2 AND2X2_237 ( .A(_abc_15497_new_n1193_), .B(_abc_15497_new_n1189_), .Y(_abc_15497_new_n1197_));
AND2X2 AND2X2_2370 ( .A(_abc_15497_new_n5561_), .B(_abc_15497_new_n5558_), .Y(_abc_15497_new_n5592_));
AND2X2 AND2X2_2371 ( .A(_abc_15497_new_n5552_), .B(_abc_15497_new_n5548_), .Y(_abc_15497_new_n5594_));
AND2X2 AND2X2_2372 ( .A(b_reg_24_), .B(c_reg_24_), .Y(_abc_15497_new_n5596_));
AND2X2 AND2X2_2373 ( .A(_abc_15497_new_n5597_), .B(_abc_15497_new_n5595_), .Y(_abc_15497_new_n5598_));
AND2X2 AND2X2_2374 ( .A(_abc_15497_new_n5598_), .B(d_reg_24_), .Y(_abc_15497_new_n5600_));
AND2X2 AND2X2_2375 ( .A(_abc_15497_new_n5601_), .B(_abc_15497_new_n5599_), .Y(_abc_15497_new_n5602_));
AND2X2 AND2X2_2376 ( .A(_abc_15497_new_n3803_), .B(_abc_15497_new_n5602_), .Y(_abc_15497_new_n5603_));
AND2X2 AND2X2_2377 ( .A(_abc_15497_new_n5606_), .B(_abc_15497_new_n5597_), .Y(_abc_15497_new_n5607_));
AND2X2 AND2X2_2378 ( .A(_abc_15497_new_n5597_), .B(_abc_15497_new_n5605_), .Y(_abc_15497_new_n5610_));
AND2X2 AND2X2_2379 ( .A(_abc_15497_new_n5612_), .B(_abc_15497_new_n5608_), .Y(_abc_15497_new_n5613_));
AND2X2 AND2X2_238 ( .A(e_reg_13_), .B(\digest[13] ), .Y(_abc_15497_new_n1199_));
AND2X2 AND2X2_2380 ( .A(_abc_15497_new_n5604_), .B(_abc_15497_new_n5613_), .Y(_abc_15497_new_n5614_));
AND2X2 AND2X2_2381 ( .A(e_reg_24_), .B(a_reg_19_), .Y(_abc_15497_new_n5619_));
AND2X2 AND2X2_2382 ( .A(_abc_15497_new_n5620_), .B(_abc_15497_new_n5618_), .Y(_abc_15497_new_n5621_));
AND2X2 AND2X2_2383 ( .A(_abc_15497_new_n5622_), .B(_abc_15497_new_n5617_), .Y(_abc_15497_new_n5623_));
AND2X2 AND2X2_2384 ( .A(_abc_15497_new_n5621_), .B(w_24_), .Y(_abc_15497_new_n5624_));
AND2X2 AND2X2_2385 ( .A(_abc_15497_new_n5626_), .B(_abc_15497_new_n5616_), .Y(_abc_15497_new_n5627_));
AND2X2 AND2X2_2386 ( .A(_abc_15497_new_n5628_), .B(_abc_15497_new_n5629_), .Y(_abc_15497_new_n5630_));
AND2X2 AND2X2_2387 ( .A(_abc_15497_new_n5615_), .B(_abc_15497_new_n5630_), .Y(_abc_15497_new_n5631_));
AND2X2 AND2X2_2388 ( .A(_abc_15497_new_n5632_), .B(_abc_15497_new_n5633_), .Y(_abc_15497_new_n5634_));
AND2X2 AND2X2_2389 ( .A(_abc_15497_new_n5635_), .B(_abc_15497_new_n5594_), .Y(_abc_15497_new_n5636_));
AND2X2 AND2X2_239 ( .A(_abc_15497_new_n1200_), .B(_abc_15497_new_n1198_), .Y(_abc_15497_new_n1201_));
AND2X2 AND2X2_2390 ( .A(_abc_15497_new_n5640_), .B(_abc_15497_new_n3774_), .Y(_abc_15497_new_n5641_));
AND2X2 AND2X2_2391 ( .A(_abc_15497_new_n5639_), .B(_abc_15497_new_n3784_), .Y(_abc_15497_new_n5642_));
AND2X2 AND2X2_2392 ( .A(_abc_15497_new_n5644_), .B(_abc_15497_new_n5593_), .Y(_abc_15497_new_n5645_));
AND2X2 AND2X2_2393 ( .A(_abc_15497_new_n5643_), .B(_abc_15497_new_n5592_), .Y(_abc_15497_new_n5646_));
AND2X2 AND2X2_2394 ( .A(_abc_15497_new_n5591_), .B(_abc_15497_new_n5648_), .Y(_abc_15497_new_n5650_));
AND2X2 AND2X2_2395 ( .A(_abc_15497_new_n5651_), .B(round_ctr_inc), .Y(_abc_15497_new_n5652_));
AND2X2 AND2X2_2396 ( .A(_abc_15497_new_n5652_), .B(_abc_15497_new_n5649_), .Y(_abc_15497_new_n5653_));
AND2X2 AND2X2_2397 ( .A(_abc_15497_new_n2010_), .B(a_reg_24_), .Y(_abc_15497_new_n5654_));
AND2X2 AND2X2_2398 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3084_), .Y(_abc_15497_new_n5655_));
AND2X2 AND2X2_2399 ( .A(_abc_15497_new_n5651_), .B(_abc_15497_new_n5658_), .Y(_abc_15497_new_n5659_));
AND2X2 AND2X2_24 ( .A(_abc_15497_new_n741_), .B(_abc_15497_new_n742_), .Y(_abc_15497_new_n743_));
AND2X2 AND2X2_240 ( .A(_abc_15497_new_n1197_), .B(_abc_15497_new_n1201_), .Y(_abc_15497_new_n1202_));
AND2X2 AND2X2_2400 ( .A(_abc_15497_new_n5632_), .B(_abc_15497_new_n5628_), .Y(_abc_15497_new_n5662_));
AND2X2 AND2X2_2401 ( .A(b_reg_25_), .B(c_reg_25_), .Y(_abc_15497_new_n5664_));
AND2X2 AND2X2_2402 ( .A(_abc_15497_new_n5665_), .B(_abc_15497_new_n5663_), .Y(_abc_15497_new_n5666_));
AND2X2 AND2X2_2403 ( .A(_abc_15497_new_n5666_), .B(d_reg_25_), .Y(_abc_15497_new_n5668_));
AND2X2 AND2X2_2404 ( .A(_abc_15497_new_n5669_), .B(_abc_15497_new_n5667_), .Y(_abc_15497_new_n5670_));
AND2X2 AND2X2_2405 ( .A(_abc_15497_new_n3803_), .B(_abc_15497_new_n5670_), .Y(_abc_15497_new_n5671_));
AND2X2 AND2X2_2406 ( .A(_abc_15497_new_n5674_), .B(_abc_15497_new_n5665_), .Y(_abc_15497_new_n5675_));
AND2X2 AND2X2_2407 ( .A(_abc_15497_new_n5665_), .B(_abc_15497_new_n5673_), .Y(_abc_15497_new_n5678_));
AND2X2 AND2X2_2408 ( .A(_abc_15497_new_n5680_), .B(_abc_15497_new_n5676_), .Y(_abc_15497_new_n5681_));
AND2X2 AND2X2_2409 ( .A(_abc_15497_new_n5672_), .B(_abc_15497_new_n5681_), .Y(_abc_15497_new_n5682_));
AND2X2 AND2X2_241 ( .A(_abc_15497_new_n1203_), .B(_abc_15497_new_n1204_), .Y(_abc_15497_new_n1205_));
AND2X2 AND2X2_2410 ( .A(e_reg_25_), .B(a_reg_20_), .Y(_abc_15497_new_n5687_));
AND2X2 AND2X2_2411 ( .A(_abc_15497_new_n5688_), .B(_abc_15497_new_n5686_), .Y(_abc_15497_new_n5689_));
AND2X2 AND2X2_2412 ( .A(_abc_15497_new_n5690_), .B(_abc_15497_new_n5685_), .Y(_abc_15497_new_n5691_));
AND2X2 AND2X2_2413 ( .A(_abc_15497_new_n5689_), .B(w_25_), .Y(_abc_15497_new_n5692_));
AND2X2 AND2X2_2414 ( .A(_abc_15497_new_n5694_), .B(_abc_15497_new_n5684_), .Y(_abc_15497_new_n5695_));
AND2X2 AND2X2_2415 ( .A(_abc_15497_new_n5696_), .B(_abc_15497_new_n5697_), .Y(_abc_15497_new_n5698_));
AND2X2 AND2X2_2416 ( .A(_abc_15497_new_n5683_), .B(_abc_15497_new_n5698_), .Y(_abc_15497_new_n5699_));
AND2X2 AND2X2_2417 ( .A(_abc_15497_new_n5700_), .B(_abc_15497_new_n5701_), .Y(_abc_15497_new_n5702_));
AND2X2 AND2X2_2418 ( .A(_abc_15497_new_n5703_), .B(_abc_15497_new_n5662_), .Y(_abc_15497_new_n5704_));
AND2X2 AND2X2_2419 ( .A(_abc_15497_new_n5705_), .B(_abc_15497_new_n5706_), .Y(_abc_15497_new_n5707_));
AND2X2 AND2X2_242 ( .A(_abc_15497_new_n1206_), .B(digest_update), .Y(_abc_15497_new_n1207_));
AND2X2 AND2X2_2420 ( .A(_abc_15497_new_n5661_), .B(_abc_15497_new_n5707_), .Y(_abc_15497_new_n5708_));
AND2X2 AND2X2_2421 ( .A(_abc_15497_new_n5715_), .B(round_ctr_inc), .Y(_abc_15497_new_n5716_));
AND2X2 AND2X2_2422 ( .A(_abc_15497_new_n5716_), .B(_abc_15497_new_n5712_), .Y(_abc_15497_new_n5717_));
AND2X2 AND2X2_2423 ( .A(_abc_15497_new_n2010_), .B(a_reg_25_), .Y(_abc_15497_new_n5718_));
AND2X2 AND2X2_2424 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3098_), .Y(_abc_15497_new_n5719_));
AND2X2 AND2X2_2425 ( .A(_abc_15497_new_n5722_), .B(_abc_15497_new_n5709_), .Y(_abc_15497_new_n5723_));
AND2X2 AND2X2_2426 ( .A(_abc_15497_new_n5591_), .B(_abc_15497_new_n5725_), .Y(_abc_15497_new_n5726_));
AND2X2 AND2X2_2427 ( .A(_abc_15497_new_n5727_), .B(_abc_15497_new_n5723_), .Y(_abc_15497_new_n5728_));
AND2X2 AND2X2_2428 ( .A(_abc_15497_new_n5700_), .B(_abc_15497_new_n5696_), .Y(_abc_15497_new_n5730_));
AND2X2 AND2X2_2429 ( .A(c_reg_26_), .B(b_reg_26_), .Y(_abc_15497_new_n5731_));
AND2X2 AND2X2_243 ( .A(_abc_15497_new_n1208_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n1209_));
AND2X2 AND2X2_2430 ( .A(_abc_15497_new_n5732_), .B(_abc_15497_new_n5733_), .Y(_abc_15497_new_n5734_));
AND2X2 AND2X2_2431 ( .A(_abc_15497_new_n5734_), .B(d_reg_26_), .Y(_abc_15497_new_n5735_));
AND2X2 AND2X2_2432 ( .A(_abc_15497_new_n5736_), .B(_abc_15497_new_n5737_), .Y(_abc_15497_new_n5738_));
AND2X2 AND2X2_2433 ( .A(_abc_15497_new_n3803_), .B(_abc_15497_new_n5738_), .Y(_abc_15497_new_n5739_));
AND2X2 AND2X2_2434 ( .A(_abc_15497_new_n5742_), .B(_abc_15497_new_n5732_), .Y(_abc_15497_new_n5743_));
AND2X2 AND2X2_2435 ( .A(_abc_15497_new_n5732_), .B(_abc_15497_new_n5741_), .Y(_abc_15497_new_n5745_));
AND2X2 AND2X2_2436 ( .A(_abc_15497_new_n5746_), .B(_abc_15497_new_n5733_), .Y(_abc_15497_new_n5747_));
AND2X2 AND2X2_2437 ( .A(_abc_15497_new_n3774_), .B(_abc_15497_new_n5747_), .Y(_abc_15497_new_n5748_));
AND2X2 AND2X2_2438 ( .A(_abc_15497_new_n5749_), .B(_abc_15497_new_n5744_), .Y(_abc_15497_new_n5750_));
AND2X2 AND2X2_2439 ( .A(_abc_15497_new_n5740_), .B(_abc_15497_new_n5750_), .Y(_abc_15497_new_n5751_));
AND2X2 AND2X2_244 ( .A(e_reg_14_), .B(\digest[14] ), .Y(_abc_15497_new_n1212_));
AND2X2 AND2X2_2440 ( .A(e_reg_26_), .B(a_reg_21_), .Y(_abc_15497_new_n5756_));
AND2X2 AND2X2_2441 ( .A(_abc_15497_new_n5757_), .B(_abc_15497_new_n5755_), .Y(_abc_15497_new_n5758_));
AND2X2 AND2X2_2442 ( .A(_abc_15497_new_n5759_), .B(_abc_15497_new_n5754_), .Y(_abc_15497_new_n5760_));
AND2X2 AND2X2_2443 ( .A(_abc_15497_new_n5758_), .B(w_26_), .Y(_abc_15497_new_n5761_));
AND2X2 AND2X2_2444 ( .A(_abc_15497_new_n5763_), .B(_abc_15497_new_n5753_), .Y(_abc_15497_new_n5764_));
AND2X2 AND2X2_2445 ( .A(_abc_15497_new_n5765_), .B(_abc_15497_new_n5766_), .Y(_abc_15497_new_n5767_));
AND2X2 AND2X2_2446 ( .A(_abc_15497_new_n5752_), .B(_abc_15497_new_n5767_), .Y(_abc_15497_new_n5768_));
AND2X2 AND2X2_2447 ( .A(_abc_15497_new_n5769_), .B(_abc_15497_new_n5770_), .Y(_abc_15497_new_n5771_));
AND2X2 AND2X2_2448 ( .A(_abc_15497_new_n5772_), .B(_abc_15497_new_n5730_), .Y(_abc_15497_new_n5773_));
AND2X2 AND2X2_2449 ( .A(_abc_15497_new_n5777_), .B(_abc_15497_new_n5011_), .Y(_abc_15497_new_n5778_));
AND2X2 AND2X2_245 ( .A(_abc_15497_new_n1213_), .B(_abc_15497_new_n1211_), .Y(_abc_15497_new_n1214_));
AND2X2 AND2X2_2450 ( .A(_abc_15497_new_n5776_), .B(_abc_15497_new_n5010_), .Y(_abc_15497_new_n5779_));
AND2X2 AND2X2_2451 ( .A(_abc_15497_new_n5781_), .B(_abc_15497_new_n5705_), .Y(_abc_15497_new_n5782_));
AND2X2 AND2X2_2452 ( .A(_abc_15497_new_n5780_), .B(_abc_15497_new_n5704_), .Y(_abc_15497_new_n5783_));
AND2X2 AND2X2_2453 ( .A(_abc_15497_new_n5729_), .B(_abc_15497_new_n5785_), .Y(_abc_15497_new_n5787_));
AND2X2 AND2X2_2454 ( .A(_abc_15497_new_n5788_), .B(round_ctr_inc), .Y(_abc_15497_new_n5789_));
AND2X2 AND2X2_2455 ( .A(_abc_15497_new_n5789_), .B(_abc_15497_new_n5786_), .Y(_abc_15497_new_n5790_));
AND2X2 AND2X2_2456 ( .A(_abc_15497_new_n2010_), .B(a_reg_26_), .Y(_abc_15497_new_n5791_));
AND2X2 AND2X2_2457 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3115_), .Y(_abc_15497_new_n5792_));
AND2X2 AND2X2_2458 ( .A(_abc_15497_new_n5769_), .B(_abc_15497_new_n5765_), .Y(_abc_15497_new_n5799_));
AND2X2 AND2X2_2459 ( .A(c_reg_27_), .B(b_reg_27_), .Y(_abc_15497_new_n5800_));
AND2X2 AND2X2_246 ( .A(_abc_15497_new_n1189_), .B(_abc_15497_new_n1200_), .Y(_abc_15497_new_n1216_));
AND2X2 AND2X2_2460 ( .A(_abc_15497_new_n5801_), .B(_abc_15497_new_n5802_), .Y(_abc_15497_new_n5803_));
AND2X2 AND2X2_2461 ( .A(_abc_15497_new_n5803_), .B(d_reg_27_), .Y(_abc_15497_new_n5804_));
AND2X2 AND2X2_2462 ( .A(_abc_15497_new_n5805_), .B(_abc_15497_new_n5806_), .Y(_abc_15497_new_n5807_));
AND2X2 AND2X2_2463 ( .A(_abc_15497_new_n3803_), .B(_abc_15497_new_n5807_), .Y(_abc_15497_new_n5808_));
AND2X2 AND2X2_2464 ( .A(_abc_15497_new_n5811_), .B(_abc_15497_new_n5801_), .Y(_abc_15497_new_n5812_));
AND2X2 AND2X2_2465 ( .A(_abc_15497_new_n5801_), .B(_abc_15497_new_n5810_), .Y(_abc_15497_new_n5814_));
AND2X2 AND2X2_2466 ( .A(_abc_15497_new_n5815_), .B(_abc_15497_new_n5802_), .Y(_abc_15497_new_n5816_));
AND2X2 AND2X2_2467 ( .A(_abc_15497_new_n3774_), .B(_abc_15497_new_n5816_), .Y(_abc_15497_new_n5817_));
AND2X2 AND2X2_2468 ( .A(_abc_15497_new_n5818_), .B(_abc_15497_new_n5813_), .Y(_abc_15497_new_n5819_));
AND2X2 AND2X2_2469 ( .A(_abc_15497_new_n5809_), .B(_abc_15497_new_n5819_), .Y(_abc_15497_new_n5820_));
AND2X2 AND2X2_247 ( .A(_abc_15497_new_n1193_), .B(_abc_15497_new_n1216_), .Y(_abc_15497_new_n1217_));
AND2X2 AND2X2_2470 ( .A(e_reg_27_), .B(a_reg_22_), .Y(_abc_15497_new_n5825_));
AND2X2 AND2X2_2471 ( .A(_abc_15497_new_n5826_), .B(_abc_15497_new_n5824_), .Y(_abc_15497_new_n5827_));
AND2X2 AND2X2_2472 ( .A(_abc_15497_new_n5828_), .B(_abc_15497_new_n5823_), .Y(_abc_15497_new_n5829_));
AND2X2 AND2X2_2473 ( .A(_abc_15497_new_n5827_), .B(w_27_), .Y(_abc_15497_new_n5830_));
AND2X2 AND2X2_2474 ( .A(_abc_15497_new_n5832_), .B(_abc_15497_new_n5822_), .Y(_abc_15497_new_n5833_));
AND2X2 AND2X2_2475 ( .A(_abc_15497_new_n5834_), .B(_abc_15497_new_n5835_), .Y(_abc_15497_new_n5836_));
AND2X2 AND2X2_2476 ( .A(_abc_15497_new_n5821_), .B(_abc_15497_new_n5836_), .Y(_abc_15497_new_n5837_));
AND2X2 AND2X2_2477 ( .A(_abc_15497_new_n5838_), .B(_abc_15497_new_n5839_), .Y(_abc_15497_new_n5840_));
AND2X2 AND2X2_2478 ( .A(_abc_15497_new_n5841_), .B(_abc_15497_new_n5799_), .Y(_abc_15497_new_n5842_));
AND2X2 AND2X2_2479 ( .A(_abc_15497_new_n5843_), .B(_abc_15497_new_n5844_), .Y(_abc_15497_new_n5845_));
AND2X2 AND2X2_248 ( .A(_abc_15497_new_n1219_), .B(_abc_15497_new_n1214_), .Y(_abc_15497_new_n1221_));
AND2X2 AND2X2_2480 ( .A(_abc_15497_new_n5798_), .B(_abc_15497_new_n5845_), .Y(_abc_15497_new_n5846_));
AND2X2 AND2X2_2481 ( .A(_abc_15497_new_n5852_), .B(round_ctr_inc), .Y(_abc_15497_new_n5853_));
AND2X2 AND2X2_2482 ( .A(_abc_15497_new_n5853_), .B(_abc_15497_new_n5850_), .Y(_abc_15497_new_n5854_));
AND2X2 AND2X2_2483 ( .A(_abc_15497_new_n2010_), .B(a_reg_27_), .Y(_abc_15497_new_n5855_));
AND2X2 AND2X2_2484 ( .A(_abc_15497_new_n700_), .B(\digest[155] ), .Y(_abc_15497_new_n5856_));
AND2X2 AND2X2_2485 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n5856_), .Y(_abc_15497_new_n5857_));
AND2X2 AND2X2_2486 ( .A(_abc_15497_new_n5851_), .B(_abc_15497_new_n5785_), .Y(_abc_15497_new_n5860_));
AND2X2 AND2X2_2487 ( .A(_abc_15497_new_n5725_), .B(_abc_15497_new_n5860_), .Y(_abc_15497_new_n5861_));
AND2X2 AND2X2_2488 ( .A(_abc_15497_new_n5851_), .B(_abc_15497_new_n5782_), .Y(_abc_15497_new_n5866_));
AND2X2 AND2X2_2489 ( .A(_abc_15497_new_n5865_), .B(_abc_15497_new_n5868_), .Y(_abc_15497_new_n5869_));
AND2X2 AND2X2_249 ( .A(_abc_15497_new_n1222_), .B(_abc_15497_new_n1220_), .Y(_abc_15497_new_n1223_));
AND2X2 AND2X2_2490 ( .A(_abc_15497_new_n5863_), .B(_abc_15497_new_n5869_), .Y(_abc_15497_new_n5870_));
AND2X2 AND2X2_2491 ( .A(_abc_15497_new_n5838_), .B(_abc_15497_new_n5834_), .Y(_abc_15497_new_n5872_));
AND2X2 AND2X2_2492 ( .A(c_reg_28_), .B(b_reg_28_), .Y(_abc_15497_new_n5873_));
AND2X2 AND2X2_2493 ( .A(_abc_15497_new_n5874_), .B(_abc_15497_new_n5875_), .Y(_abc_15497_new_n5876_));
AND2X2 AND2X2_2494 ( .A(_abc_15497_new_n5876_), .B(d_reg_28_), .Y(_abc_15497_new_n5877_));
AND2X2 AND2X2_2495 ( .A(_abc_15497_new_n5878_), .B(_abc_15497_new_n5879_), .Y(_abc_15497_new_n5880_));
AND2X2 AND2X2_2496 ( .A(_abc_15497_new_n3803_), .B(_abc_15497_new_n5880_), .Y(_abc_15497_new_n5881_));
AND2X2 AND2X2_2497 ( .A(_abc_15497_new_n5884_), .B(_abc_15497_new_n5874_), .Y(_abc_15497_new_n5885_));
AND2X2 AND2X2_2498 ( .A(_abc_15497_new_n5874_), .B(_abc_15497_new_n5883_), .Y(_abc_15497_new_n5887_));
AND2X2 AND2X2_2499 ( .A(_abc_15497_new_n5888_), .B(_abc_15497_new_n5875_), .Y(_abc_15497_new_n5889_));
AND2X2 AND2X2_25 ( .A(c_reg_16_), .B(\digest[80] ), .Y(_abc_15497_new_n745_));
AND2X2 AND2X2_250 ( .A(_abc_15497_new_n1223_), .B(digest_update), .Y(_abc_15497_new_n1224_));
AND2X2 AND2X2_2500 ( .A(_abc_15497_new_n3774_), .B(_abc_15497_new_n5889_), .Y(_abc_15497_new_n5890_));
AND2X2 AND2X2_2501 ( .A(_abc_15497_new_n5891_), .B(_abc_15497_new_n5886_), .Y(_abc_15497_new_n5892_));
AND2X2 AND2X2_2502 ( .A(_abc_15497_new_n5882_), .B(_abc_15497_new_n5892_), .Y(_abc_15497_new_n5893_));
AND2X2 AND2X2_2503 ( .A(e_reg_28_), .B(a_reg_23_), .Y(_abc_15497_new_n5898_));
AND2X2 AND2X2_2504 ( .A(_abc_15497_new_n5899_), .B(_abc_15497_new_n5897_), .Y(_abc_15497_new_n5900_));
AND2X2 AND2X2_2505 ( .A(_abc_15497_new_n5901_), .B(_abc_15497_new_n5896_), .Y(_abc_15497_new_n5902_));
AND2X2 AND2X2_2506 ( .A(_abc_15497_new_n5900_), .B(w_28_), .Y(_abc_15497_new_n5903_));
AND2X2 AND2X2_2507 ( .A(_abc_15497_new_n5905_), .B(_abc_15497_new_n5895_), .Y(_abc_15497_new_n5906_));
AND2X2 AND2X2_2508 ( .A(_abc_15497_new_n5907_), .B(_abc_15497_new_n5908_), .Y(_abc_15497_new_n5909_));
AND2X2 AND2X2_2509 ( .A(_abc_15497_new_n5894_), .B(_abc_15497_new_n5909_), .Y(_abc_15497_new_n5910_));
AND2X2 AND2X2_251 ( .A(_abc_15497_new_n1225_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n1226_));
AND2X2 AND2X2_2510 ( .A(_abc_15497_new_n5911_), .B(_abc_15497_new_n5912_), .Y(_abc_15497_new_n5913_));
AND2X2 AND2X2_2511 ( .A(_abc_15497_new_n5914_), .B(_abc_15497_new_n5872_), .Y(_abc_15497_new_n5915_));
AND2X2 AND2X2_2512 ( .A(_abc_15497_new_n5919_), .B(_abc_15497_new_n3753_), .Y(_abc_15497_new_n5920_));
AND2X2 AND2X2_2513 ( .A(_abc_15497_new_n5918_), .B(_abc_15497_new_n3780_), .Y(_abc_15497_new_n5921_));
AND2X2 AND2X2_2514 ( .A(_abc_15497_new_n5922_), .B(_abc_15497_new_n5842_), .Y(_abc_15497_new_n5923_));
AND2X2 AND2X2_2515 ( .A(_abc_15497_new_n5871_), .B(_abc_15497_new_n5927_), .Y(_abc_15497_new_n5929_));
AND2X2 AND2X2_2516 ( .A(_abc_15497_new_n5930_), .B(round_ctr_inc), .Y(_abc_15497_new_n5931_));
AND2X2 AND2X2_2517 ( .A(_abc_15497_new_n5931_), .B(_abc_15497_new_n5928_), .Y(_abc_15497_new_n5932_));
AND2X2 AND2X2_2518 ( .A(_abc_15497_new_n2010_), .B(a_reg_28_), .Y(_abc_15497_new_n5933_));
AND2X2 AND2X2_2519 ( .A(_abc_15497_new_n700_), .B(\digest[156] ), .Y(_abc_15497_new_n5934_));
AND2X2 AND2X2_252 ( .A(_abc_15497_new_n1222_), .B(_abc_15497_new_n1213_), .Y(_abc_15497_new_n1228_));
AND2X2 AND2X2_2520 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n5934_), .Y(_abc_15497_new_n5935_));
AND2X2 AND2X2_2521 ( .A(_abc_15497_new_n5930_), .B(_abc_15497_new_n5924_), .Y(_abc_15497_new_n5938_));
AND2X2 AND2X2_2522 ( .A(_abc_15497_new_n5911_), .B(_abc_15497_new_n5907_), .Y(_abc_15497_new_n5941_));
AND2X2 AND2X2_2523 ( .A(c_reg_29_), .B(b_reg_29_), .Y(_abc_15497_new_n5942_));
AND2X2 AND2X2_2524 ( .A(_abc_15497_new_n5943_), .B(d_reg_29_), .Y(_abc_15497_new_n5944_));
AND2X2 AND2X2_2525 ( .A(_abc_15497_new_n5948_), .B(_abc_15497_new_n5949_), .Y(_abc_15497_new_n5950_));
AND2X2 AND2X2_2526 ( .A(_abc_15497_new_n5950_), .B(_abc_15497_new_n5947_), .Y(_abc_15497_new_n5951_));
AND2X2 AND2X2_2527 ( .A(_abc_15497_new_n5952_), .B(_abc_15497_new_n5953_), .Y(_abc_15497_new_n5954_));
AND2X2 AND2X2_2528 ( .A(_abc_15497_new_n5948_), .B(_abc_15497_new_n5947_), .Y(_abc_15497_new_n5956_));
AND2X2 AND2X2_2529 ( .A(_abc_15497_new_n5957_), .B(_abc_15497_new_n5949_), .Y(_abc_15497_new_n5958_));
AND2X2 AND2X2_253 ( .A(e_reg_15_), .B(\digest[15] ), .Y(_abc_15497_new_n1230_));
AND2X2 AND2X2_2530 ( .A(_abc_15497_new_n3774_), .B(_abc_15497_new_n5958_), .Y(_abc_15497_new_n5959_));
AND2X2 AND2X2_2531 ( .A(_abc_15497_new_n5961_), .B(_abc_15497_new_n5955_), .Y(_abc_15497_new_n5962_));
AND2X2 AND2X2_2532 ( .A(_abc_15497_new_n5963_), .B(_abc_15497_new_n5946_), .Y(_abc_15497_new_n5964_));
AND2X2 AND2X2_2533 ( .A(e_reg_29_), .B(a_reg_24_), .Y(_abc_15497_new_n5968_));
AND2X2 AND2X2_2534 ( .A(_abc_15497_new_n5969_), .B(_abc_15497_new_n5967_), .Y(_abc_15497_new_n5970_));
AND2X2 AND2X2_2535 ( .A(_abc_15497_new_n5971_), .B(_abc_15497_new_n5966_), .Y(_abc_15497_new_n5972_));
AND2X2 AND2X2_2536 ( .A(_abc_15497_new_n5970_), .B(w_29_), .Y(_abc_15497_new_n5973_));
AND2X2 AND2X2_2537 ( .A(_abc_15497_new_n5975_), .B(_abc_15497_new_n5965_), .Y(_abc_15497_new_n5976_));
AND2X2 AND2X2_2538 ( .A(_abc_15497_new_n5977_), .B(_abc_15497_new_n5978_), .Y(_abc_15497_new_n5979_));
AND2X2 AND2X2_2539 ( .A(_abc_15497_new_n5964_), .B(_abc_15497_new_n5979_), .Y(_abc_15497_new_n5980_));
AND2X2 AND2X2_254 ( .A(_abc_15497_new_n1231_), .B(_abc_15497_new_n1229_), .Y(_abc_15497_new_n1232_));
AND2X2 AND2X2_2540 ( .A(_abc_15497_new_n5981_), .B(_abc_15497_new_n5982_), .Y(_abc_15497_new_n5983_));
AND2X2 AND2X2_2541 ( .A(_abc_15497_new_n5984_), .B(_abc_15497_new_n5941_), .Y(_abc_15497_new_n5985_));
AND2X2 AND2X2_2542 ( .A(_abc_15497_new_n5988_), .B(_abc_15497_new_n4060_), .Y(_abc_15497_new_n5989_));
AND2X2 AND2X2_2543 ( .A(_abc_15497_new_n5992_), .B(_abc_15497_new_n5940_), .Y(_abc_15497_new_n5993_));
AND2X2 AND2X2_2544 ( .A(_abc_15497_new_n6000_), .B(round_ctr_inc), .Y(_abc_15497_new_n6001_));
AND2X2 AND2X2_2545 ( .A(_abc_15497_new_n6001_), .B(_abc_15497_new_n5997_), .Y(_abc_15497_new_n6002_));
AND2X2 AND2X2_2546 ( .A(_abc_15497_new_n2010_), .B(a_reg_29_), .Y(_abc_15497_new_n6003_));
AND2X2 AND2X2_2547 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3164_), .Y(_abc_15497_new_n6004_));
AND2X2 AND2X2_2548 ( .A(_abc_15497_new_n5999_), .B(_abc_15497_new_n5927_), .Y(_abc_15497_new_n6007_));
AND2X2 AND2X2_2549 ( .A(_abc_15497_new_n5999_), .B(_abc_15497_new_n5925_), .Y(_abc_15497_new_n6010_));
AND2X2 AND2X2_255 ( .A(_abc_15497_new_n1228_), .B(_abc_15497_new_n1232_), .Y(_abc_15497_new_n1233_));
AND2X2 AND2X2_2550 ( .A(_abc_15497_new_n6009_), .B(_abc_15497_new_n6012_), .Y(_abc_15497_new_n6013_));
AND2X2 AND2X2_2551 ( .A(_abc_15497_new_n5990_), .B(_abc_15497_new_n5986_), .Y(_abc_15497_new_n6015_));
AND2X2 AND2X2_2552 ( .A(_abc_15497_new_n5981_), .B(_abc_15497_new_n5977_), .Y(_abc_15497_new_n6016_));
AND2X2 AND2X2_2553 ( .A(c_reg_30_), .B(b_reg_30_), .Y(_abc_15497_new_n6017_));
AND2X2 AND2X2_2554 ( .A(_abc_15497_new_n6018_), .B(d_reg_30_), .Y(_abc_15497_new_n6019_));
AND2X2 AND2X2_2555 ( .A(_abc_15497_new_n6023_), .B(_abc_15497_new_n6024_), .Y(_abc_15497_new_n6025_));
AND2X2 AND2X2_2556 ( .A(_abc_15497_new_n6025_), .B(_abc_15497_new_n6022_), .Y(_abc_15497_new_n6026_));
AND2X2 AND2X2_2557 ( .A(_abc_15497_new_n6027_), .B(_abc_15497_new_n6028_), .Y(_abc_15497_new_n6029_));
AND2X2 AND2X2_2558 ( .A(_abc_15497_new_n6023_), .B(_abc_15497_new_n6022_), .Y(_abc_15497_new_n6031_));
AND2X2 AND2X2_2559 ( .A(_abc_15497_new_n6032_), .B(_abc_15497_new_n6024_), .Y(_abc_15497_new_n6033_));
AND2X2 AND2X2_256 ( .A(_abc_15497_new_n1234_), .B(_abc_15497_new_n1235_), .Y(_abc_15497_new_n1236_));
AND2X2 AND2X2_2560 ( .A(_abc_15497_new_n3774_), .B(_abc_15497_new_n6033_), .Y(_abc_15497_new_n6034_));
AND2X2 AND2X2_2561 ( .A(_abc_15497_new_n6036_), .B(_abc_15497_new_n6030_), .Y(_abc_15497_new_n6037_));
AND2X2 AND2X2_2562 ( .A(_abc_15497_new_n6038_), .B(_abc_15497_new_n6021_), .Y(_abc_15497_new_n6039_));
AND2X2 AND2X2_2563 ( .A(e_reg_30_), .B(a_reg_25_), .Y(_abc_15497_new_n6043_));
AND2X2 AND2X2_2564 ( .A(_abc_15497_new_n6044_), .B(_abc_15497_new_n6042_), .Y(_abc_15497_new_n6045_));
AND2X2 AND2X2_2565 ( .A(_abc_15497_new_n6046_), .B(_abc_15497_new_n6041_), .Y(_abc_15497_new_n6047_));
AND2X2 AND2X2_2566 ( .A(_abc_15497_new_n6045_), .B(w_30_), .Y(_abc_15497_new_n6048_));
AND2X2 AND2X2_2567 ( .A(_abc_15497_new_n6050_), .B(_abc_15497_new_n6040_), .Y(_abc_15497_new_n6051_));
AND2X2 AND2X2_2568 ( .A(_abc_15497_new_n6052_), .B(_abc_15497_new_n6053_), .Y(_abc_15497_new_n6054_));
AND2X2 AND2X2_2569 ( .A(_abc_15497_new_n6039_), .B(_abc_15497_new_n6054_), .Y(_abc_15497_new_n6055_));
AND2X2 AND2X2_257 ( .A(_abc_15497_new_n1237_), .B(digest_update), .Y(_abc_15497_new_n1238_));
AND2X2 AND2X2_2570 ( .A(_abc_15497_new_n6056_), .B(_abc_15497_new_n6057_), .Y(_abc_15497_new_n6058_));
AND2X2 AND2X2_2571 ( .A(_abc_15497_new_n6059_), .B(_abc_15497_new_n6016_), .Y(_abc_15497_new_n6060_));
AND2X2 AND2X2_2572 ( .A(_abc_15497_new_n6064_), .B(_abc_15497_new_n3784_), .Y(_abc_15497_new_n6065_));
AND2X2 AND2X2_2573 ( .A(_abc_15497_new_n6063_), .B(_abc_15497_new_n3774_), .Y(_abc_15497_new_n6066_));
AND2X2 AND2X2_2574 ( .A(_abc_15497_new_n6067_), .B(_abc_15497_new_n6015_), .Y(_abc_15497_new_n6068_));
AND2X2 AND2X2_2575 ( .A(_abc_15497_new_n6074_), .B(round_ctr_inc), .Y(_abc_15497_new_n6075_));
AND2X2 AND2X2_2576 ( .A(_abc_15497_new_n6075_), .B(_abc_15497_new_n6073_), .Y(_abc_15497_new_n6076_));
AND2X2 AND2X2_2577 ( .A(_abc_15497_new_n2010_), .B(a_reg_30_), .Y(_abc_15497_new_n6077_));
AND2X2 AND2X2_2578 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n3181_), .Y(_abc_15497_new_n6078_));
AND2X2 AND2X2_2579 ( .A(_abc_15497_new_n6074_), .B(_abc_15497_new_n6069_), .Y(_abc_15497_new_n6081_));
AND2X2 AND2X2_258 ( .A(_abc_15497_new_n1239_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n1240_));
AND2X2 AND2X2_2580 ( .A(_abc_15497_new_n6056_), .B(_abc_15497_new_n6052_), .Y(_abc_15497_new_n6085_));
AND2X2 AND2X2_2581 ( .A(c_reg_31_), .B(b_reg_31_), .Y(_abc_15497_new_n6087_));
AND2X2 AND2X2_2582 ( .A(_abc_15497_new_n6090_), .B(_abc_15497_new_n6088_), .Y(_abc_15497_new_n6091_));
AND2X2 AND2X2_2583 ( .A(_abc_15497_new_n3753_), .B(_abc_15497_new_n6091_), .Y(_abc_15497_new_n6092_));
AND2X2 AND2X2_2584 ( .A(_abc_15497_new_n997_), .B(_abc_15497_new_n2698_), .Y(_abc_15497_new_n6093_));
AND2X2 AND2X2_2585 ( .A(_abc_15497_new_n6094_), .B(_abc_15497_new_n6088_), .Y(_abc_15497_new_n6095_));
AND2X2 AND2X2_2586 ( .A(_abc_15497_new_n6095_), .B(_abc_15497_new_n6089_), .Y(_abc_15497_new_n6096_));
AND2X2 AND2X2_2587 ( .A(_abc_15497_new_n6097_), .B(_abc_15497_new_n6098_), .Y(_abc_15497_new_n6099_));
AND2X2 AND2X2_2588 ( .A(_abc_15497_new_n6088_), .B(_abc_15497_new_n6089_), .Y(_abc_15497_new_n6101_));
AND2X2 AND2X2_2589 ( .A(_abc_15497_new_n6103_), .B(_abc_15497_new_n3780_), .Y(_abc_15497_new_n6104_));
AND2X2 AND2X2_259 ( .A(_abc_15497_new_n701_), .B(\digest[16] ), .Y(_abc_15497_new_n1242_));
AND2X2 AND2X2_2590 ( .A(_abc_15497_new_n6100_), .B(_abc_15497_new_n6104_), .Y(_abc_15497_new_n6105_));
AND2X2 AND2X2_2591 ( .A(e_reg_31_), .B(w_31_), .Y(_abc_15497_new_n6111_));
AND2X2 AND2X2_2592 ( .A(_abc_15497_new_n6112_), .B(_abc_15497_new_n6110_), .Y(_abc_15497_new_n6113_));
AND2X2 AND2X2_2593 ( .A(_abc_15497_new_n6113_), .B(a_reg_26_), .Y(_abc_15497_new_n6114_));
AND2X2 AND2X2_2594 ( .A(_abc_15497_new_n6115_), .B(_abc_15497_new_n6116_), .Y(_abc_15497_new_n6117_));
AND2X2 AND2X2_2595 ( .A(_abc_15497_new_n6118_), .B(_abc_15497_new_n6109_), .Y(_abc_15497_new_n6119_));
AND2X2 AND2X2_2596 ( .A(_abc_15497_new_n6117_), .B(_abc_15497_new_n6108_), .Y(_abc_15497_new_n6120_));
AND2X2 AND2X2_2597 ( .A(_abc_15497_new_n6107_), .B(_abc_15497_new_n6122_), .Y(_abc_15497_new_n6123_));
AND2X2 AND2X2_2598 ( .A(_abc_15497_new_n6106_), .B(_abc_15497_new_n6121_), .Y(_abc_15497_new_n6124_));
AND2X2 AND2X2_2599 ( .A(_abc_15497_new_n6086_), .B(_abc_15497_new_n6125_), .Y(_abc_15497_new_n6126_));
AND2X2 AND2X2_26 ( .A(_abc_15497_new_n747_), .B(_abc_15497_new_n741_), .Y(_abc_15497_new_n748_));
AND2X2 AND2X2_260 ( .A(_abc_15497_new_n1190_), .B(_abc_15497_new_n1201_), .Y(_abc_15497_new_n1243_));
AND2X2 AND2X2_2600 ( .A(_abc_15497_new_n6127_), .B(_abc_15497_new_n6128_), .Y(_abc_15497_new_n6129_));
AND2X2 AND2X2_2601 ( .A(_abc_15497_new_n6132_), .B(_abc_15497_new_n6130_), .Y(_abc_15497_new_n6133_));
AND2X2 AND2X2_2602 ( .A(_abc_15497_new_n6084_), .B(_abc_15497_new_n6133_), .Y(_abc_15497_new_n6134_));
AND2X2 AND2X2_2603 ( .A(_abc_15497_new_n6135_), .B(_abc_15497_new_n6136_), .Y(_abc_15497_new_n6137_));
AND2X2 AND2X2_2604 ( .A(_abc_15497_new_n6140_), .B(round_ctr_inc), .Y(_abc_15497_new_n6141_));
AND2X2 AND2X2_2605 ( .A(_abc_15497_new_n6141_), .B(_abc_15497_new_n6138_), .Y(_abc_15497_new_n6142_));
AND2X2 AND2X2_2606 ( .A(_abc_15497_new_n2010_), .B(a_reg_31_), .Y(_abc_15497_new_n6143_));
AND2X2 AND2X2_2607 ( .A(_abc_15497_new_n700_), .B(\digest[159] ), .Y(_abc_15497_new_n6144_));
AND2X2 AND2X2_2608 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n6144_), .Y(_abc_15497_new_n6145_));
AND2X2 AND2X2_2609 ( .A(round_ctr_reg_1_), .B(round_ctr_reg_0_), .Y(_abc_15497_new_n6148_));
AND2X2 AND2X2_261 ( .A(_abc_15497_new_n1214_), .B(_abc_15497_new_n1232_), .Y(_abc_15497_new_n1244_));
AND2X2 AND2X2_2610 ( .A(_abc_15497_new_n3770_), .B(_abc_15497_new_n6148_), .Y(_abc_15497_new_n6149_));
AND2X2 AND2X2_2611 ( .A(_abc_15497_new_n3747_), .B(round_ctr_reg_6_), .Y(_abc_15497_new_n6150_));
AND2X2 AND2X2_2612 ( .A(_abc_15497_new_n6150_), .B(_abc_15497_new_n6149_), .Y(_abc_15497_new_n6151_));
AND2X2 AND2X2_2613 ( .A(_abc_15497_new_n6151_), .B(round_ctr_inc), .Y(_abc_15497_abc_9717_auto_fsm_map_cc_118_implement_pattern_cache_863));
AND2X2 AND2X2_2614 ( .A(_abc_15497_new_n6154_), .B(round_ctr_inc), .Y(_abc_15497_new_n6155_));
AND2X2 AND2X2_2615 ( .A(_abc_15497_new_n6156_), .B(ready), .Y(_abc_15497_new_n6157_));
AND2X2 AND2X2_2616 ( .A(_abc_15497_new_n6155_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n6159_));
AND2X2 AND2X2_2617 ( .A(_abc_15497_new_n6162_), .B(_abc_15497_new_n6163_), .Y(_0round_ctr_reg_6_0__0_));
AND2X2 AND2X2_2618 ( .A(_abc_15497_new_n2010_), .B(round_ctr_reg_1_), .Y(_abc_15497_new_n6165_));
AND2X2 AND2X2_2619 ( .A(_abc_15497_new_n6166_), .B(_abc_15497_new_n6167_), .Y(_abc_15497_new_n6168_));
AND2X2 AND2X2_262 ( .A(_abc_15497_new_n1243_), .B(_abc_15497_new_n1244_), .Y(_abc_15497_new_n1245_));
AND2X2 AND2X2_2620 ( .A(_abc_15497_new_n6168_), .B(round_ctr_inc), .Y(_abc_15497_new_n6169_));
AND2X2 AND2X2_2621 ( .A(_abc_15497_new_n2010_), .B(round_ctr_reg_2_), .Y(_abc_15497_new_n6171_));
AND2X2 AND2X2_2622 ( .A(_abc_15497_new_n6148_), .B(round_ctr_reg_2_), .Y(_abc_15497_new_n6172_));
AND2X2 AND2X2_2623 ( .A(_abc_15497_new_n6173_), .B(_abc_15497_new_n6174_), .Y(_abc_15497_new_n6175_));
AND2X2 AND2X2_2624 ( .A(_abc_15497_new_n6175_), .B(round_ctr_inc), .Y(_abc_15497_new_n6176_));
AND2X2 AND2X2_2625 ( .A(_abc_15497_new_n6178_), .B(round_ctr_reg_3_), .Y(_abc_15497_new_n6179_));
AND2X2 AND2X2_2626 ( .A(_abc_15497_new_n6172_), .B(round_ctr_inc), .Y(_abc_15497_new_n6180_));
AND2X2 AND2X2_2627 ( .A(_abc_15497_new_n6149_), .B(round_ctr_inc), .Y(_abc_15497_new_n6182_));
AND2X2 AND2X2_2628 ( .A(_abc_15497_new_n6181_), .B(_abc_15497_new_n6183_), .Y(_0round_ctr_reg_6_0__3_));
AND2X2 AND2X2_2629 ( .A(_abc_15497_new_n6178_), .B(round_ctr_reg_4_), .Y(_abc_15497_new_n6185_));
AND2X2 AND2X2_263 ( .A(_abc_15497_new_n1183_), .B(_abc_15497_new_n1245_), .Y(_abc_15497_new_n1246_));
AND2X2 AND2X2_2630 ( .A(_abc_15497_new_n6182_), .B(round_ctr_reg_4_), .Y(_abc_15497_new_n6187_));
AND2X2 AND2X2_2631 ( .A(_abc_15497_new_n6186_), .B(_abc_15497_new_n6188_), .Y(_0round_ctr_reg_6_0__4_));
AND2X2 AND2X2_2632 ( .A(_abc_15497_new_n6178_), .B(round_ctr_reg_5_), .Y(_abc_15497_new_n6190_));
AND2X2 AND2X2_2633 ( .A(_abc_15497_new_n6149_), .B(_abc_15497_new_n3738_), .Y(_abc_15497_new_n6192_));
AND2X2 AND2X2_2634 ( .A(_abc_15497_new_n6192_), .B(round_ctr_inc), .Y(_abc_15497_new_n6193_));
AND2X2 AND2X2_2635 ( .A(_abc_15497_new_n6191_), .B(_abc_15497_new_n6194_), .Y(_0round_ctr_reg_6_0__5_));
AND2X2 AND2X2_2636 ( .A(_abc_15497_new_n6194_), .B(_abc_15497_new_n6178_), .Y(_abc_15497_new_n6196_));
AND2X2 AND2X2_2637 ( .A(_abc_15497_new_n6197_), .B(_abc_15497_new_n6198_), .Y(_0round_ctr_reg_6_0__6_));
AND2X2 AND2X2_2638 ( .A(_abc_15497_new_n2009_), .B(digest_valid), .Y(_abc_15497_new_n6200_));
AND2X2 AND2X2_2639 ( .A(_abc_15497_new_n948_), .B(digest_update), .Y(_abc_15497_new_n6203_));
AND2X2 AND2X2_264 ( .A(_abc_15497_new_n1229_), .B(_abc_15497_new_n1212_), .Y(_abc_15497_new_n1247_));
AND2X2 AND2X2_2640 ( .A(_abc_15497_new_n6203_), .B(_abc_15497_new_n6202_), .Y(_abc_15497_new_n6204_));
AND2X2 AND2X2_2641 ( .A(_abc_15497_new_n701_), .B(\digest[64] ), .Y(_abc_15497_new_n6205_));
AND2X2 AND2X2_2642 ( .A(_abc_15497_new_n951_), .B(_abc_15497_new_n6207_), .Y(_abc_15497_new_n6208_));
AND2X2 AND2X2_2643 ( .A(_abc_15497_new_n6209_), .B(_abc_15497_new_n6210_), .Y(_0H2_reg_31_0__1_));
AND2X2 AND2X2_2644 ( .A(_abc_15497_new_n954_), .B(_abc_15497_new_n6212_), .Y(_abc_15497_new_n6213_));
AND2X2 AND2X2_2645 ( .A(_abc_15497_new_n6214_), .B(_abc_15497_new_n6215_), .Y(_0H2_reg_31_0__2_));
AND2X2 AND2X2_2646 ( .A(_abc_15497_new_n946_), .B(_abc_15497_new_n816_), .Y(_abc_15497_new_n6217_));
AND2X2 AND2X2_2647 ( .A(_abc_15497_new_n6220_), .B(_abc_15497_new_n6218_), .Y(_abc_15497_new_n6221_));
AND2X2 AND2X2_2648 ( .A(_abc_15497_new_n6221_), .B(digest_update), .Y(_abc_15497_new_n6222_));
AND2X2 AND2X2_2649 ( .A(_abc_15497_new_n3568_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n6223_));
AND2X2 AND2X2_265 ( .A(_abc_15497_new_n1250_), .B(_abc_15497_new_n1244_), .Y(_abc_15497_new_n1251_));
AND2X2 AND2X2_2650 ( .A(_abc_15497_new_n959_), .B(_abc_15497_new_n6225_), .Y(_abc_15497_new_n6226_));
AND2X2 AND2X2_2651 ( .A(_abc_15497_new_n6227_), .B(_abc_15497_new_n6228_), .Y(_0H2_reg_31_0__4_));
AND2X2 AND2X2_2652 ( .A(_abc_15497_new_n944_), .B(_abc_15497_new_n813_), .Y(_abc_15497_new_n6231_));
AND2X2 AND2X2_2653 ( .A(_abc_15497_new_n960_), .B(_abc_15497_new_n6231_), .Y(_abc_15497_new_n6232_));
AND2X2 AND2X2_2654 ( .A(_abc_15497_new_n836_), .B(_abc_15497_new_n6233_), .Y(_abc_15497_new_n6234_));
AND2X2 AND2X2_2655 ( .A(_abc_15497_new_n6236_), .B(_abc_15497_new_n6230_), .Y(_0H2_reg_31_0__5_));
AND2X2 AND2X2_2656 ( .A(_abc_15497_new_n838_), .B(_abc_15497_new_n810_), .Y(_abc_15497_new_n6239_));
AND2X2 AND2X2_2657 ( .A(_abc_15497_new_n6240_), .B(_abc_15497_new_n6238_), .Y(_abc_15497_new_n6241_));
AND2X2 AND2X2_2658 ( .A(_abc_15497_new_n6241_), .B(digest_update), .Y(_abc_15497_new_n6242_));
AND2X2 AND2X2_2659 ( .A(_abc_15497_new_n3586_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n6243_));
AND2X2 AND2X2_266 ( .A(_abc_15497_new_n1184_), .B(_abc_15497_new_n1245_), .Y(_abc_15497_new_n1254_));
AND2X2 AND2X2_2660 ( .A(_abc_15497_new_n6240_), .B(_abc_15497_new_n808_), .Y(_abc_15497_new_n6245_));
AND2X2 AND2X2_2661 ( .A(_abc_15497_new_n6247_), .B(_abc_15497_new_n6249_), .Y(_abc_15497_new_n6250_));
AND2X2 AND2X2_2662 ( .A(_abc_15497_new_n6250_), .B(digest_update), .Y(_abc_15497_new_n6251_));
AND2X2 AND2X2_2663 ( .A(_abc_15497_new_n3592_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n6252_));
AND2X2 AND2X2_2664 ( .A(_abc_15497_new_n701_), .B(\digest[72] ), .Y(_abc_15497_new_n6254_));
AND2X2 AND2X2_2665 ( .A(_abc_15497_new_n840_), .B(_abc_15497_new_n845_), .Y(_abc_15497_new_n6256_));
AND2X2 AND2X2_2666 ( .A(_abc_15497_new_n6257_), .B(_abc_15497_new_n6255_), .Y(_abc_15497_new_n6258_));
AND2X2 AND2X2_2667 ( .A(_abc_15497_new_n6258_), .B(digest_update), .Y(_abc_15497_new_n6259_));
AND2X2 AND2X2_2668 ( .A(_abc_15497_new_n701_), .B(\digest[73] ), .Y(_abc_15497_new_n6261_));
AND2X2 AND2X2_2669 ( .A(_abc_15497_new_n6257_), .B(_abc_15497_new_n843_), .Y(_abc_15497_new_n6262_));
AND2X2 AND2X2_267 ( .A(_abc_15497_new_n1123_), .B(_abc_15497_new_n1254_), .Y(_abc_15497_new_n1255_));
AND2X2 AND2X2_2670 ( .A(_abc_15497_new_n6266_), .B(digest_update), .Y(_abc_15497_new_n6267_));
AND2X2 AND2X2_2671 ( .A(_abc_15497_new_n6267_), .B(_abc_15497_new_n6264_), .Y(_abc_15497_new_n6268_));
AND2X2 AND2X2_2672 ( .A(_abc_15497_new_n848_), .B(_abc_15497_new_n794_), .Y(_abc_15497_new_n6271_));
AND2X2 AND2X2_2673 ( .A(_abc_15497_new_n6272_), .B(_abc_15497_new_n6270_), .Y(_abc_15497_new_n6273_));
AND2X2 AND2X2_2674 ( .A(_abc_15497_new_n6273_), .B(digest_update), .Y(_abc_15497_new_n6274_));
AND2X2 AND2X2_2675 ( .A(_abc_15497_new_n3610_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n6275_));
AND2X2 AND2X2_2676 ( .A(_abc_15497_new_n6272_), .B(_abc_15497_new_n792_), .Y(_abc_15497_new_n6277_));
AND2X2 AND2X2_2677 ( .A(_abc_15497_new_n6279_), .B(_abc_15497_new_n6281_), .Y(_abc_15497_new_n6282_));
AND2X2 AND2X2_2678 ( .A(_abc_15497_new_n6282_), .B(digest_update), .Y(_abc_15497_new_n6283_));
AND2X2 AND2X2_2679 ( .A(_abc_15497_new_n3616_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n6284_));
AND2X2 AND2X2_268 ( .A(e_reg_16_), .B(\digest[16] ), .Y(_abc_15497_new_n1258_));
AND2X2 AND2X2_2680 ( .A(_abc_15497_new_n850_), .B(_abc_15497_new_n782_), .Y(_abc_15497_new_n6287_));
AND2X2 AND2X2_2681 ( .A(_abc_15497_new_n6288_), .B(_abc_15497_new_n6286_), .Y(_abc_15497_new_n6289_));
AND2X2 AND2X2_2682 ( .A(_abc_15497_new_n6289_), .B(digest_update), .Y(_abc_15497_new_n6290_));
AND2X2 AND2X2_2683 ( .A(_abc_15497_new_n3622_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n6291_));
AND2X2 AND2X2_2684 ( .A(_abc_15497_new_n701_), .B(\digest[77] ), .Y(_abc_15497_new_n6293_));
AND2X2 AND2X2_2685 ( .A(_abc_15497_new_n6288_), .B(_abc_15497_new_n770_), .Y(_abc_15497_new_n6294_));
AND2X2 AND2X2_2686 ( .A(_abc_15497_new_n6297_), .B(digest_update), .Y(_abc_15497_new_n6298_));
AND2X2 AND2X2_2687 ( .A(_abc_15497_new_n6298_), .B(_abc_15497_new_n6296_), .Y(_abc_15497_new_n6299_));
AND2X2 AND2X2_2688 ( .A(_abc_15497_new_n850_), .B(_abc_15497_new_n783_), .Y(_abc_15497_new_n6301_));
AND2X2 AND2X2_2689 ( .A(_abc_15497_new_n6302_), .B(_abc_15497_new_n765_), .Y(_abc_15497_new_n6304_));
AND2X2 AND2X2_269 ( .A(_abc_15497_new_n1259_), .B(_abc_15497_new_n1257_), .Y(_abc_15497_new_n1260_));
AND2X2 AND2X2_2690 ( .A(_abc_15497_new_n6305_), .B(_abc_15497_new_n6303_), .Y(_abc_15497_new_n6306_));
AND2X2 AND2X2_2691 ( .A(_abc_15497_new_n6306_), .B(digest_update), .Y(_abc_15497_new_n6307_));
AND2X2 AND2X2_2692 ( .A(_abc_15497_new_n3634_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n6308_));
AND2X2 AND2X2_2693 ( .A(_abc_15497_new_n6305_), .B(_abc_15497_new_n763_), .Y(_abc_15497_new_n6310_));
AND2X2 AND2X2_2694 ( .A(_abc_15497_new_n6312_), .B(_abc_15497_new_n6314_), .Y(_abc_15497_new_n6315_));
AND2X2 AND2X2_2695 ( .A(_abc_15497_new_n6315_), .B(digest_update), .Y(_abc_15497_new_n6316_));
AND2X2 AND2X2_2696 ( .A(_abc_15497_new_n3640_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n6317_));
AND2X2 AND2X2_2697 ( .A(_abc_15497_new_n701_), .B(\digest[80] ), .Y(_abc_15497_new_n6319_));
AND2X2 AND2X2_2698 ( .A(_abc_15497_new_n852_), .B(_abc_15497_new_n854_), .Y(_abc_15497_new_n6321_));
AND2X2 AND2X2_2699 ( .A(_abc_15497_new_n6322_), .B(_abc_15497_new_n6320_), .Y(_abc_15497_new_n6323_));
AND2X2 AND2X2_27 ( .A(_abc_15497_new_n749_), .B(_abc_15497_new_n739_), .Y(_abc_15497_new_n750_));
AND2X2 AND2X2_270 ( .A(_abc_15497_new_n1256_), .B(_abc_15497_new_n1260_), .Y(_abc_15497_new_n1262_));
AND2X2 AND2X2_2700 ( .A(_abc_15497_new_n6323_), .B(digest_update), .Y(_abc_15497_new_n6324_));
AND2X2 AND2X2_2701 ( .A(_abc_15497_new_n6322_), .B(_abc_15497_new_n746_), .Y(_abc_15497_new_n6326_));
AND2X2 AND2X2_2702 ( .A(_abc_15497_new_n6328_), .B(_abc_15497_new_n6329_), .Y(_abc_15497_new_n6330_));
AND2X2 AND2X2_2703 ( .A(_abc_15497_new_n6330_), .B(digest_update), .Y(_abc_15497_new_n6331_));
AND2X2 AND2X2_2704 ( .A(_abc_15497_new_n3652_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n6332_));
AND2X2 AND2X2_2705 ( .A(_abc_15497_new_n701_), .B(\digest[82] ), .Y(_abc_15497_new_n6334_));
AND2X2 AND2X2_2706 ( .A(_abc_15497_new_n852_), .B(_abc_15497_new_n855_), .Y(_abc_15497_new_n6335_));
AND2X2 AND2X2_2707 ( .A(_abc_15497_new_n6336_), .B(_abc_15497_new_n738_), .Y(_abc_15497_new_n6338_));
AND2X2 AND2X2_2708 ( .A(_abc_15497_new_n6339_), .B(_abc_15497_new_n6337_), .Y(_abc_15497_new_n6340_));
AND2X2 AND2X2_2709 ( .A(_abc_15497_new_n6340_), .B(digest_update), .Y(_abc_15497_new_n6341_));
AND2X2 AND2X2_271 ( .A(_abc_15497_new_n1263_), .B(_abc_15497_new_n1261_), .Y(_abc_15497_new_n1264_));
AND2X2 AND2X2_2710 ( .A(_abc_15497_new_n6339_), .B(_abc_15497_new_n736_), .Y(_abc_15497_new_n6343_));
AND2X2 AND2X2_2711 ( .A(_abc_15497_new_n6343_), .B(_abc_15497_new_n734_), .Y(_abc_15497_new_n6344_));
AND2X2 AND2X2_2712 ( .A(_abc_15497_new_n6346_), .B(_abc_15497_new_n6345_), .Y(_abc_15497_new_n6347_));
AND2X2 AND2X2_2713 ( .A(_abc_15497_new_n6348_), .B(digest_update), .Y(_abc_15497_new_n6349_));
AND2X2 AND2X2_2714 ( .A(_abc_15497_new_n3664_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n6350_));
AND2X2 AND2X2_2715 ( .A(_abc_15497_new_n852_), .B(_abc_15497_new_n856_), .Y(_abc_15497_new_n6352_));
AND2X2 AND2X2_2716 ( .A(_abc_15497_new_n6353_), .B(_abc_15497_new_n728_), .Y(_abc_15497_new_n6355_));
AND2X2 AND2X2_2717 ( .A(_abc_15497_new_n6356_), .B(_abc_15497_new_n6354_), .Y(_abc_15497_new_n6357_));
AND2X2 AND2X2_2718 ( .A(_abc_15497_new_n6357_), .B(digest_update), .Y(_abc_15497_new_n6358_));
AND2X2 AND2X2_2719 ( .A(_abc_15497_new_n3670_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n6359_));
AND2X2 AND2X2_272 ( .A(_abc_15497_new_n1264_), .B(digest_update), .Y(_abc_15497_new_n1265_));
AND2X2 AND2X2_2720 ( .A(_abc_15497_new_n6363_), .B(_abc_15497_new_n718_), .Y(_abc_15497_new_n6364_));
AND2X2 AND2X2_2721 ( .A(_abc_15497_new_n6362_), .B(_abc_15497_new_n719_), .Y(_abc_15497_new_n6365_));
AND2X2 AND2X2_2722 ( .A(_abc_15497_new_n6367_), .B(_abc_15497_new_n6361_), .Y(_0H2_reg_31_0__21_));
AND2X2 AND2X2_2723 ( .A(_abc_15497_new_n701_), .B(\digest[86] ), .Y(_abc_15497_new_n6369_));
AND2X2 AND2X2_2724 ( .A(_abc_15497_new_n6362_), .B(_abc_15497_new_n717_), .Y(_abc_15497_new_n6370_));
AND2X2 AND2X2_2725 ( .A(_abc_15497_new_n6371_), .B(_abc_15497_new_n710_), .Y(_abc_15497_new_n6373_));
AND2X2 AND2X2_2726 ( .A(_abc_15497_new_n6374_), .B(_abc_15497_new_n6372_), .Y(_abc_15497_new_n6375_));
AND2X2 AND2X2_2727 ( .A(_abc_15497_new_n6375_), .B(digest_update), .Y(_abc_15497_new_n6376_));
AND2X2 AND2X2_2728 ( .A(_abc_15497_new_n6379_), .B(_abc_15497_new_n706_), .Y(_abc_15497_new_n6380_));
AND2X2 AND2X2_2729 ( .A(_abc_15497_new_n6378_), .B(_abc_15497_new_n6381_), .Y(_abc_15497_new_n6382_));
AND2X2 AND2X2_273 ( .A(_abc_15497_new_n1263_), .B(_abc_15497_new_n1259_), .Y(_abc_15497_new_n1267_));
AND2X2 AND2X2_2730 ( .A(_abc_15497_new_n6384_), .B(_abc_15497_new_n6385_), .Y(_0H2_reg_31_0__23_));
AND2X2 AND2X2_2731 ( .A(_abc_15497_new_n701_), .B(\digest[88] ), .Y(_abc_15497_new_n6387_));
AND2X2 AND2X2_2732 ( .A(_abc_15497_new_n859_), .B(_abc_15497_new_n867_), .Y(_abc_15497_new_n6389_));
AND2X2 AND2X2_2733 ( .A(_abc_15497_new_n6390_), .B(_abc_15497_new_n6388_), .Y(_abc_15497_new_n6391_));
AND2X2 AND2X2_2734 ( .A(_abc_15497_new_n6391_), .B(digest_update), .Y(_abc_15497_new_n6392_));
AND2X2 AND2X2_2735 ( .A(_abc_15497_new_n701_), .B(\digest[89] ), .Y(_abc_15497_new_n6394_));
AND2X2 AND2X2_2736 ( .A(_abc_15497_new_n6390_), .B(_abc_15497_new_n865_), .Y(_abc_15497_new_n6395_));
AND2X2 AND2X2_2737 ( .A(_abc_15497_new_n6399_), .B(digest_update), .Y(_abc_15497_new_n6400_));
AND2X2 AND2X2_2738 ( .A(_abc_15497_new_n6400_), .B(_abc_15497_new_n6397_), .Y(_abc_15497_new_n6401_));
AND2X2 AND2X2_2739 ( .A(w_mem_inst__abc_21203_new_n1589_), .B(w_mem_inst__abc_21203_new_n1591_), .Y(w_mem_inst__abc_21203_new_n1592_));
AND2X2 AND2X2_274 ( .A(e_reg_17_), .B(\digest[17] ), .Y(_abc_15497_new_n1270_));
AND2X2 AND2X2_2740 ( .A(w_mem_inst_w_mem_2__31_), .B(w_mem_inst_w_mem_0__31_), .Y(w_mem_inst__abc_21203_new_n1595_));
AND2X2 AND2X2_2741 ( .A(w_mem_inst__abc_21203_new_n1596_), .B(w_mem_inst__abc_21203_new_n1594_), .Y(w_mem_inst__abc_21203_new_n1597_));
AND2X2 AND2X2_2742 ( .A(w_mem_inst__abc_21203_new_n1598_), .B(w_mem_inst__abc_21203_new_n1600_), .Y(w_mem_inst__abc_21203_new_n1601_));
AND2X2 AND2X2_2743 ( .A(w_mem_inst__abc_21203_new_n1603_), .B(w_mem_inst_w_ctr_reg_0_), .Y(w_mem_inst__abc_21203_new_n1604_));
AND2X2 AND2X2_2744 ( .A(w_mem_inst__abc_21203_new_n1605_), .B(w_mem_inst_w_ctr_reg_2_), .Y(w_mem_inst__abc_21203_new_n1606_));
AND2X2 AND2X2_2745 ( .A(w_mem_inst__abc_21203_new_n1604_), .B(w_mem_inst__abc_21203_new_n1606_), .Y(w_mem_inst__abc_21203_new_n1607_));
AND2X2 AND2X2_2746 ( .A(w_mem_inst__abc_21203_new_n1607_), .B(w_mem_inst_w_mem_5__0_), .Y(w_mem_inst__abc_21203_new_n1608_));
AND2X2 AND2X2_2747 ( .A(w_mem_inst__abc_21203_new_n1603_), .B(w_mem_inst__abc_21203_new_n1610_), .Y(w_mem_inst__abc_21203_new_n1611_));
AND2X2 AND2X2_2748 ( .A(w_mem_inst__abc_21203_new_n1612_), .B(w_mem_inst_w_ctr_reg_3_), .Y(w_mem_inst__abc_21203_new_n1613_));
AND2X2 AND2X2_2749 ( .A(w_mem_inst__abc_21203_new_n1611_), .B(w_mem_inst__abc_21203_new_n1613_), .Y(w_mem_inst__abc_21203_new_n1614_));
AND2X2 AND2X2_275 ( .A(_abc_15497_new_n1271_), .B(_abc_15497_new_n1269_), .Y(_abc_15497_new_n1272_));
AND2X2 AND2X2_2750 ( .A(w_mem_inst__abc_21203_new_n1614_), .B(w_mem_inst_w_mem_8__0_), .Y(w_mem_inst__abc_21203_new_n1615_));
AND2X2 AND2X2_2751 ( .A(w_mem_inst_w_ctr_reg_1_), .B(w_mem_inst_w_ctr_reg_0_), .Y(w_mem_inst__abc_21203_new_n1616_));
AND2X2 AND2X2_2752 ( .A(w_mem_inst__abc_21203_new_n1613_), .B(w_mem_inst__abc_21203_new_n1616_), .Y(w_mem_inst__abc_21203_new_n1617_));
AND2X2 AND2X2_2753 ( .A(w_mem_inst__abc_21203_new_n1617_), .B(w_mem_inst_w_mem_11__0_), .Y(w_mem_inst__abc_21203_new_n1618_));
AND2X2 AND2X2_2754 ( .A(w_mem_inst__abc_21203_new_n1606_), .B(w_mem_inst__abc_21203_new_n1616_), .Y(w_mem_inst__abc_21203_new_n1621_));
AND2X2 AND2X2_2755 ( .A(w_mem_inst__abc_21203_new_n1621_), .B(w_mem_inst_w_mem_7__0_), .Y(w_mem_inst__abc_21203_new_n1622_));
AND2X2 AND2X2_2756 ( .A(w_mem_inst_w_ctr_reg_3_), .B(w_mem_inst_w_ctr_reg_2_), .Y(w_mem_inst__abc_21203_new_n1623_));
AND2X2 AND2X2_2757 ( .A(w_mem_inst__abc_21203_new_n1616_), .B(w_mem_inst__abc_21203_new_n1623_), .Y(w_mem_inst__abc_21203_new_n1624_));
AND2X2 AND2X2_2758 ( .A(w_mem_inst__abc_21203_new_n1624_), .B(w_mem_inst_w_mem_15__0_), .Y(w_mem_inst__abc_21203_new_n1625_));
AND2X2 AND2X2_2759 ( .A(w_mem_inst__abc_21203_new_n1604_), .B(w_mem_inst__abc_21203_new_n1623_), .Y(w_mem_inst__abc_21203_new_n1628_));
AND2X2 AND2X2_276 ( .A(_abc_15497_new_n1273_), .B(_abc_15497_new_n1275_), .Y(_abc_15497_new_n1276_));
AND2X2 AND2X2_2760 ( .A(w_mem_inst__abc_21203_new_n1628_), .B(w_mem_inst_w_mem_13__0_), .Y(w_mem_inst__abc_21203_new_n1629_));
AND2X2 AND2X2_2761 ( .A(w_mem_inst__abc_21203_new_n1605_), .B(w_mem_inst__abc_21203_new_n1612_), .Y(w_mem_inst__abc_21203_new_n1630_));
AND2X2 AND2X2_2762 ( .A(w_mem_inst__abc_21203_new_n1611_), .B(w_mem_inst__abc_21203_new_n1630_), .Y(w_mem_inst__abc_21203_new_n1631_));
AND2X2 AND2X2_2763 ( .A(w_mem_inst__abc_21203_new_n1631_), .B(w_mem_inst_w_mem_0__0_), .Y(w_mem_inst__abc_21203_new_n1632_));
AND2X2 AND2X2_2764 ( .A(w_mem_inst__abc_21203_new_n1611_), .B(w_mem_inst__abc_21203_new_n1623_), .Y(w_mem_inst__abc_21203_new_n1633_));
AND2X2 AND2X2_2765 ( .A(w_mem_inst__abc_21203_new_n1633_), .B(w_mem_inst_w_mem_12__0_), .Y(w_mem_inst__abc_21203_new_n1634_));
AND2X2 AND2X2_2766 ( .A(w_mem_inst__abc_21203_new_n1604_), .B(w_mem_inst__abc_21203_new_n1613_), .Y(w_mem_inst__abc_21203_new_n1637_));
AND2X2 AND2X2_2767 ( .A(w_mem_inst__abc_21203_new_n1637_), .B(w_mem_inst_w_mem_9__0_), .Y(w_mem_inst__abc_21203_new_n1638_));
AND2X2 AND2X2_2768 ( .A(w_mem_inst__abc_21203_new_n1610_), .B(w_mem_inst_w_ctr_reg_1_), .Y(w_mem_inst__abc_21203_new_n1639_));
AND2X2 AND2X2_2769 ( .A(w_mem_inst__abc_21203_new_n1613_), .B(w_mem_inst__abc_21203_new_n1639_), .Y(w_mem_inst__abc_21203_new_n1640_));
AND2X2 AND2X2_277 ( .A(_abc_15497_new_n1276_), .B(digest_update), .Y(_abc_15497_new_n1277_));
AND2X2 AND2X2_2770 ( .A(w_mem_inst__abc_21203_new_n1640_), .B(w_mem_inst_w_mem_10__0_), .Y(w_mem_inst__abc_21203_new_n1641_));
AND2X2 AND2X2_2771 ( .A(w_mem_inst__abc_21203_new_n1611_), .B(w_mem_inst__abc_21203_new_n1606_), .Y(w_mem_inst__abc_21203_new_n1643_));
AND2X2 AND2X2_2772 ( .A(w_mem_inst__abc_21203_new_n1643_), .B(w_mem_inst_w_mem_4__0_), .Y(w_mem_inst__abc_21203_new_n1644_));
AND2X2 AND2X2_2773 ( .A(w_mem_inst__abc_21203_new_n1606_), .B(w_mem_inst__abc_21203_new_n1639_), .Y(w_mem_inst__abc_21203_new_n1645_));
AND2X2 AND2X2_2774 ( .A(w_mem_inst__abc_21203_new_n1645_), .B(w_mem_inst_w_mem_6__0_), .Y(w_mem_inst__abc_21203_new_n1646_));
AND2X2 AND2X2_2775 ( .A(w_mem_inst__abc_21203_new_n1630_), .B(w_mem_inst__abc_21203_new_n1604_), .Y(w_mem_inst__abc_21203_new_n1649_));
AND2X2 AND2X2_2776 ( .A(w_mem_inst__abc_21203_new_n1649_), .B(w_mem_inst_w_mem_1__0_), .Y(w_mem_inst__abc_21203_new_n1650_));
AND2X2 AND2X2_2777 ( .A(w_mem_inst__abc_21203_new_n1630_), .B(w_mem_inst__abc_21203_new_n1639_), .Y(w_mem_inst__abc_21203_new_n1651_));
AND2X2 AND2X2_2778 ( .A(w_mem_inst__abc_21203_new_n1651_), .B(w_mem_inst_w_mem_2__0_), .Y(w_mem_inst__abc_21203_new_n1652_));
AND2X2 AND2X2_2779 ( .A(w_mem_inst__abc_21203_new_n1630_), .B(w_mem_inst__abc_21203_new_n1616_), .Y(w_mem_inst__abc_21203_new_n1654_));
AND2X2 AND2X2_278 ( .A(_abc_15497_new_n1278_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n1279_));
AND2X2 AND2X2_2780 ( .A(w_mem_inst__abc_21203_new_n1654_), .B(w_mem_inst_w_mem_3__0_), .Y(w_mem_inst__abc_21203_new_n1655_));
AND2X2 AND2X2_2781 ( .A(w_mem_inst__abc_21203_new_n1639_), .B(w_mem_inst__abc_21203_new_n1623_), .Y(w_mem_inst__abc_21203_new_n1656_));
AND2X2 AND2X2_2782 ( .A(w_mem_inst__abc_21203_new_n1656_), .B(w_mem_inst_w_mem_14__0_), .Y(w_mem_inst__abc_21203_new_n1657_));
AND2X2 AND2X2_2783 ( .A(w_mem_inst__abc_21203_new_n1662_), .B(w_mem_inst__abc_21203_new_n1602_), .Y(w_0_));
AND2X2 AND2X2_2784 ( .A(w_mem_inst__abc_21203_new_n1665_), .B(w_mem_inst__abc_21203_new_n1667_), .Y(w_mem_inst__abc_21203_new_n1668_));
AND2X2 AND2X2_2785 ( .A(w_mem_inst_w_mem_2__0_), .B(w_mem_inst_w_mem_0__0_), .Y(w_mem_inst__abc_21203_new_n1671_));
AND2X2 AND2X2_2786 ( .A(w_mem_inst__abc_21203_new_n1672_), .B(w_mem_inst__abc_21203_new_n1670_), .Y(w_mem_inst__abc_21203_new_n1673_));
AND2X2 AND2X2_2787 ( .A(w_mem_inst__abc_21203_new_n1674_), .B(w_mem_inst__abc_21203_new_n1676_), .Y(w_mem_inst__abc_21203_new_n1677_));
AND2X2 AND2X2_2788 ( .A(w_mem_inst__abc_21203_new_n1607_), .B(w_mem_inst_w_mem_5__1_), .Y(w_mem_inst__abc_21203_new_n1679_));
AND2X2 AND2X2_2789 ( .A(w_mem_inst__abc_21203_new_n1614_), .B(w_mem_inst_w_mem_8__1_), .Y(w_mem_inst__abc_21203_new_n1681_));
AND2X2 AND2X2_279 ( .A(_abc_15497_new_n701_), .B(\digest[18] ), .Y(_abc_15497_new_n1281_));
AND2X2 AND2X2_2790 ( .A(w_mem_inst__abc_21203_new_n1617_), .B(w_mem_inst_w_mem_11__1_), .Y(w_mem_inst__abc_21203_new_n1682_));
AND2X2 AND2X2_2791 ( .A(w_mem_inst__abc_21203_new_n1621_), .B(w_mem_inst_w_mem_7__1_), .Y(w_mem_inst__abc_21203_new_n1685_));
AND2X2 AND2X2_2792 ( .A(w_mem_inst__abc_21203_new_n1624_), .B(w_mem_inst_w_mem_15__1_), .Y(w_mem_inst__abc_21203_new_n1686_));
AND2X2 AND2X2_2793 ( .A(w_mem_inst__abc_21203_new_n1628_), .B(w_mem_inst_w_mem_13__1_), .Y(w_mem_inst__abc_21203_new_n1689_));
AND2X2 AND2X2_2794 ( .A(w_mem_inst__abc_21203_new_n1631_), .B(w_mem_inst_w_mem_0__1_), .Y(w_mem_inst__abc_21203_new_n1690_));
AND2X2 AND2X2_2795 ( .A(w_mem_inst__abc_21203_new_n1633_), .B(w_mem_inst_w_mem_12__1_), .Y(w_mem_inst__abc_21203_new_n1691_));
AND2X2 AND2X2_2796 ( .A(w_mem_inst__abc_21203_new_n1637_), .B(w_mem_inst_w_mem_9__1_), .Y(w_mem_inst__abc_21203_new_n1694_));
AND2X2 AND2X2_2797 ( .A(w_mem_inst__abc_21203_new_n1640_), .B(w_mem_inst_w_mem_10__1_), .Y(w_mem_inst__abc_21203_new_n1695_));
AND2X2 AND2X2_2798 ( .A(w_mem_inst__abc_21203_new_n1643_), .B(w_mem_inst_w_mem_4__1_), .Y(w_mem_inst__abc_21203_new_n1697_));
AND2X2 AND2X2_2799 ( .A(w_mem_inst__abc_21203_new_n1645_), .B(w_mem_inst_w_mem_6__1_), .Y(w_mem_inst__abc_21203_new_n1698_));
AND2X2 AND2X2_28 ( .A(_abc_15497_new_n733_), .B(_abc_15497_new_n735_), .Y(_abc_15497_new_n751_));
AND2X2 AND2X2_280 ( .A(e_reg_18_), .B(\digest[18] ), .Y(_abc_15497_new_n1283_));
AND2X2 AND2X2_2800 ( .A(w_mem_inst__abc_21203_new_n1649_), .B(w_mem_inst_w_mem_1__1_), .Y(w_mem_inst__abc_21203_new_n1701_));
AND2X2 AND2X2_2801 ( .A(w_mem_inst__abc_21203_new_n1651_), .B(w_mem_inst_w_mem_2__1_), .Y(w_mem_inst__abc_21203_new_n1702_));
AND2X2 AND2X2_2802 ( .A(w_mem_inst__abc_21203_new_n1654_), .B(w_mem_inst_w_mem_3__1_), .Y(w_mem_inst__abc_21203_new_n1704_));
AND2X2 AND2X2_2803 ( .A(w_mem_inst__abc_21203_new_n1656_), .B(w_mem_inst_w_mem_14__1_), .Y(w_mem_inst__abc_21203_new_n1705_));
AND2X2 AND2X2_2804 ( .A(w_mem_inst__abc_21203_new_n1710_), .B(w_mem_inst__abc_21203_new_n1678_), .Y(w_1_));
AND2X2 AND2X2_2805 ( .A(w_mem_inst__abc_21203_new_n1713_), .B(w_mem_inst__abc_21203_new_n1715_), .Y(w_mem_inst__abc_21203_new_n1716_));
AND2X2 AND2X2_2806 ( .A(w_mem_inst_w_mem_2__1_), .B(w_mem_inst_w_mem_0__1_), .Y(w_mem_inst__abc_21203_new_n1719_));
AND2X2 AND2X2_2807 ( .A(w_mem_inst__abc_21203_new_n1720_), .B(w_mem_inst__abc_21203_new_n1718_), .Y(w_mem_inst__abc_21203_new_n1721_));
AND2X2 AND2X2_2808 ( .A(w_mem_inst__abc_21203_new_n1722_), .B(w_mem_inst__abc_21203_new_n1724_), .Y(w_mem_inst__abc_21203_new_n1725_));
AND2X2 AND2X2_2809 ( .A(w_mem_inst__abc_21203_new_n1607_), .B(w_mem_inst_w_mem_5__2_), .Y(w_mem_inst__abc_21203_new_n1727_));
AND2X2 AND2X2_281 ( .A(_abc_15497_new_n1284_), .B(_abc_15497_new_n1282_), .Y(_abc_15497_new_n1285_));
AND2X2 AND2X2_2810 ( .A(w_mem_inst__abc_21203_new_n1614_), .B(w_mem_inst_w_mem_8__2_), .Y(w_mem_inst__abc_21203_new_n1729_));
AND2X2 AND2X2_2811 ( .A(w_mem_inst__abc_21203_new_n1617_), .B(w_mem_inst_w_mem_11__2_), .Y(w_mem_inst__abc_21203_new_n1730_));
AND2X2 AND2X2_2812 ( .A(w_mem_inst__abc_21203_new_n1621_), .B(w_mem_inst_w_mem_7__2_), .Y(w_mem_inst__abc_21203_new_n1733_));
AND2X2 AND2X2_2813 ( .A(w_mem_inst__abc_21203_new_n1624_), .B(w_mem_inst_w_mem_15__2_), .Y(w_mem_inst__abc_21203_new_n1734_));
AND2X2 AND2X2_2814 ( .A(w_mem_inst__abc_21203_new_n1628_), .B(w_mem_inst_w_mem_13__2_), .Y(w_mem_inst__abc_21203_new_n1737_));
AND2X2 AND2X2_2815 ( .A(w_mem_inst__abc_21203_new_n1631_), .B(w_mem_inst_w_mem_0__2_), .Y(w_mem_inst__abc_21203_new_n1738_));
AND2X2 AND2X2_2816 ( .A(w_mem_inst__abc_21203_new_n1633_), .B(w_mem_inst_w_mem_12__2_), .Y(w_mem_inst__abc_21203_new_n1739_));
AND2X2 AND2X2_2817 ( .A(w_mem_inst__abc_21203_new_n1637_), .B(w_mem_inst_w_mem_9__2_), .Y(w_mem_inst__abc_21203_new_n1742_));
AND2X2 AND2X2_2818 ( .A(w_mem_inst__abc_21203_new_n1640_), .B(w_mem_inst_w_mem_10__2_), .Y(w_mem_inst__abc_21203_new_n1743_));
AND2X2 AND2X2_2819 ( .A(w_mem_inst__abc_21203_new_n1643_), .B(w_mem_inst_w_mem_4__2_), .Y(w_mem_inst__abc_21203_new_n1745_));
AND2X2 AND2X2_282 ( .A(_abc_15497_new_n1259_), .B(_abc_15497_new_n1271_), .Y(_abc_15497_new_n1287_));
AND2X2 AND2X2_2820 ( .A(w_mem_inst__abc_21203_new_n1645_), .B(w_mem_inst_w_mem_6__2_), .Y(w_mem_inst__abc_21203_new_n1746_));
AND2X2 AND2X2_2821 ( .A(w_mem_inst__abc_21203_new_n1649_), .B(w_mem_inst_w_mem_1__2_), .Y(w_mem_inst__abc_21203_new_n1749_));
AND2X2 AND2X2_2822 ( .A(w_mem_inst__abc_21203_new_n1651_), .B(w_mem_inst_w_mem_2__2_), .Y(w_mem_inst__abc_21203_new_n1750_));
AND2X2 AND2X2_2823 ( .A(w_mem_inst__abc_21203_new_n1654_), .B(w_mem_inst_w_mem_3__2_), .Y(w_mem_inst__abc_21203_new_n1752_));
AND2X2 AND2X2_2824 ( .A(w_mem_inst__abc_21203_new_n1656_), .B(w_mem_inst_w_mem_14__2_), .Y(w_mem_inst__abc_21203_new_n1753_));
AND2X2 AND2X2_2825 ( .A(w_mem_inst__abc_21203_new_n1758_), .B(w_mem_inst__abc_21203_new_n1726_), .Y(w_2_));
AND2X2 AND2X2_2826 ( .A(w_mem_inst__abc_21203_new_n1761_), .B(w_mem_inst__abc_21203_new_n1763_), .Y(w_mem_inst__abc_21203_new_n1764_));
AND2X2 AND2X2_2827 ( .A(w_mem_inst_w_mem_2__2_), .B(w_mem_inst_w_mem_0__2_), .Y(w_mem_inst__abc_21203_new_n1767_));
AND2X2 AND2X2_2828 ( .A(w_mem_inst__abc_21203_new_n1768_), .B(w_mem_inst__abc_21203_new_n1766_), .Y(w_mem_inst__abc_21203_new_n1769_));
AND2X2 AND2X2_2829 ( .A(w_mem_inst__abc_21203_new_n1770_), .B(w_mem_inst__abc_21203_new_n1772_), .Y(w_mem_inst__abc_21203_new_n1773_));
AND2X2 AND2X2_283 ( .A(_abc_15497_new_n1263_), .B(_abc_15497_new_n1287_), .Y(_abc_15497_new_n1288_));
AND2X2 AND2X2_2830 ( .A(w_mem_inst__abc_21203_new_n1607_), .B(w_mem_inst_w_mem_5__3_), .Y(w_mem_inst__abc_21203_new_n1775_));
AND2X2 AND2X2_2831 ( .A(w_mem_inst__abc_21203_new_n1614_), .B(w_mem_inst_w_mem_8__3_), .Y(w_mem_inst__abc_21203_new_n1777_));
AND2X2 AND2X2_2832 ( .A(w_mem_inst__abc_21203_new_n1617_), .B(w_mem_inst_w_mem_11__3_), .Y(w_mem_inst__abc_21203_new_n1778_));
AND2X2 AND2X2_2833 ( .A(w_mem_inst__abc_21203_new_n1621_), .B(w_mem_inst_w_mem_7__3_), .Y(w_mem_inst__abc_21203_new_n1781_));
AND2X2 AND2X2_2834 ( .A(w_mem_inst__abc_21203_new_n1624_), .B(w_mem_inst_w_mem_15__3_), .Y(w_mem_inst__abc_21203_new_n1782_));
AND2X2 AND2X2_2835 ( .A(w_mem_inst__abc_21203_new_n1628_), .B(w_mem_inst_w_mem_13__3_), .Y(w_mem_inst__abc_21203_new_n1785_));
AND2X2 AND2X2_2836 ( .A(w_mem_inst__abc_21203_new_n1631_), .B(w_mem_inst_w_mem_0__3_), .Y(w_mem_inst__abc_21203_new_n1786_));
AND2X2 AND2X2_2837 ( .A(w_mem_inst__abc_21203_new_n1633_), .B(w_mem_inst_w_mem_12__3_), .Y(w_mem_inst__abc_21203_new_n1787_));
AND2X2 AND2X2_2838 ( .A(w_mem_inst__abc_21203_new_n1637_), .B(w_mem_inst_w_mem_9__3_), .Y(w_mem_inst__abc_21203_new_n1790_));
AND2X2 AND2X2_2839 ( .A(w_mem_inst__abc_21203_new_n1640_), .B(w_mem_inst_w_mem_10__3_), .Y(w_mem_inst__abc_21203_new_n1791_));
AND2X2 AND2X2_284 ( .A(_abc_15497_new_n1290_), .B(_abc_15497_new_n1285_), .Y(_abc_15497_new_n1292_));
AND2X2 AND2X2_2840 ( .A(w_mem_inst__abc_21203_new_n1643_), .B(w_mem_inst_w_mem_4__3_), .Y(w_mem_inst__abc_21203_new_n1793_));
AND2X2 AND2X2_2841 ( .A(w_mem_inst__abc_21203_new_n1645_), .B(w_mem_inst_w_mem_6__3_), .Y(w_mem_inst__abc_21203_new_n1794_));
AND2X2 AND2X2_2842 ( .A(w_mem_inst__abc_21203_new_n1649_), .B(w_mem_inst_w_mem_1__3_), .Y(w_mem_inst__abc_21203_new_n1797_));
AND2X2 AND2X2_2843 ( .A(w_mem_inst__abc_21203_new_n1651_), .B(w_mem_inst_w_mem_2__3_), .Y(w_mem_inst__abc_21203_new_n1798_));
AND2X2 AND2X2_2844 ( .A(w_mem_inst__abc_21203_new_n1654_), .B(w_mem_inst_w_mem_3__3_), .Y(w_mem_inst__abc_21203_new_n1800_));
AND2X2 AND2X2_2845 ( .A(w_mem_inst__abc_21203_new_n1656_), .B(w_mem_inst_w_mem_14__3_), .Y(w_mem_inst__abc_21203_new_n1801_));
AND2X2 AND2X2_2846 ( .A(w_mem_inst__abc_21203_new_n1806_), .B(w_mem_inst__abc_21203_new_n1774_), .Y(w_3_));
AND2X2 AND2X2_2847 ( .A(w_mem_inst__abc_21203_new_n1809_), .B(w_mem_inst__abc_21203_new_n1811_), .Y(w_mem_inst__abc_21203_new_n1812_));
AND2X2 AND2X2_2848 ( .A(w_mem_inst_w_mem_2__3_), .B(w_mem_inst_w_mem_0__3_), .Y(w_mem_inst__abc_21203_new_n1815_));
AND2X2 AND2X2_2849 ( .A(w_mem_inst__abc_21203_new_n1816_), .B(w_mem_inst__abc_21203_new_n1814_), .Y(w_mem_inst__abc_21203_new_n1817_));
AND2X2 AND2X2_285 ( .A(_abc_15497_new_n1293_), .B(_abc_15497_new_n1291_), .Y(_abc_15497_new_n1294_));
AND2X2 AND2X2_2850 ( .A(w_mem_inst__abc_21203_new_n1818_), .B(w_mem_inst__abc_21203_new_n1820_), .Y(w_mem_inst__abc_21203_new_n1821_));
AND2X2 AND2X2_2851 ( .A(w_mem_inst__abc_21203_new_n1607_), .B(w_mem_inst_w_mem_5__4_), .Y(w_mem_inst__abc_21203_new_n1823_));
AND2X2 AND2X2_2852 ( .A(w_mem_inst__abc_21203_new_n1614_), .B(w_mem_inst_w_mem_8__4_), .Y(w_mem_inst__abc_21203_new_n1825_));
AND2X2 AND2X2_2853 ( .A(w_mem_inst__abc_21203_new_n1617_), .B(w_mem_inst_w_mem_11__4_), .Y(w_mem_inst__abc_21203_new_n1826_));
AND2X2 AND2X2_2854 ( .A(w_mem_inst__abc_21203_new_n1621_), .B(w_mem_inst_w_mem_7__4_), .Y(w_mem_inst__abc_21203_new_n1829_));
AND2X2 AND2X2_2855 ( .A(w_mem_inst__abc_21203_new_n1624_), .B(w_mem_inst_w_mem_15__4_), .Y(w_mem_inst__abc_21203_new_n1830_));
AND2X2 AND2X2_2856 ( .A(w_mem_inst__abc_21203_new_n1628_), .B(w_mem_inst_w_mem_13__4_), .Y(w_mem_inst__abc_21203_new_n1833_));
AND2X2 AND2X2_2857 ( .A(w_mem_inst__abc_21203_new_n1631_), .B(w_mem_inst_w_mem_0__4_), .Y(w_mem_inst__abc_21203_new_n1834_));
AND2X2 AND2X2_2858 ( .A(w_mem_inst__abc_21203_new_n1633_), .B(w_mem_inst_w_mem_12__4_), .Y(w_mem_inst__abc_21203_new_n1835_));
AND2X2 AND2X2_2859 ( .A(w_mem_inst__abc_21203_new_n1637_), .B(w_mem_inst_w_mem_9__4_), .Y(w_mem_inst__abc_21203_new_n1838_));
AND2X2 AND2X2_286 ( .A(_abc_15497_new_n1294_), .B(digest_update), .Y(_abc_15497_new_n1295_));
AND2X2 AND2X2_2860 ( .A(w_mem_inst__abc_21203_new_n1640_), .B(w_mem_inst_w_mem_10__4_), .Y(w_mem_inst__abc_21203_new_n1839_));
AND2X2 AND2X2_2861 ( .A(w_mem_inst__abc_21203_new_n1643_), .B(w_mem_inst_w_mem_4__4_), .Y(w_mem_inst__abc_21203_new_n1841_));
AND2X2 AND2X2_2862 ( .A(w_mem_inst__abc_21203_new_n1645_), .B(w_mem_inst_w_mem_6__4_), .Y(w_mem_inst__abc_21203_new_n1842_));
AND2X2 AND2X2_2863 ( .A(w_mem_inst__abc_21203_new_n1649_), .B(w_mem_inst_w_mem_1__4_), .Y(w_mem_inst__abc_21203_new_n1845_));
AND2X2 AND2X2_2864 ( .A(w_mem_inst__abc_21203_new_n1651_), .B(w_mem_inst_w_mem_2__4_), .Y(w_mem_inst__abc_21203_new_n1846_));
AND2X2 AND2X2_2865 ( .A(w_mem_inst__abc_21203_new_n1654_), .B(w_mem_inst_w_mem_3__4_), .Y(w_mem_inst__abc_21203_new_n1848_));
AND2X2 AND2X2_2866 ( .A(w_mem_inst__abc_21203_new_n1656_), .B(w_mem_inst_w_mem_14__4_), .Y(w_mem_inst__abc_21203_new_n1849_));
AND2X2 AND2X2_2867 ( .A(w_mem_inst__abc_21203_new_n1854_), .B(w_mem_inst__abc_21203_new_n1822_), .Y(w_4_));
AND2X2 AND2X2_2868 ( .A(w_mem_inst__abc_21203_new_n1857_), .B(w_mem_inst__abc_21203_new_n1859_), .Y(w_mem_inst__abc_21203_new_n1860_));
AND2X2 AND2X2_2869 ( .A(w_mem_inst_w_mem_2__4_), .B(w_mem_inst_w_mem_0__4_), .Y(w_mem_inst__abc_21203_new_n1863_));
AND2X2 AND2X2_287 ( .A(_abc_15497_new_n701_), .B(\digest[19] ), .Y(_abc_15497_new_n1297_));
AND2X2 AND2X2_2870 ( .A(w_mem_inst__abc_21203_new_n1864_), .B(w_mem_inst__abc_21203_new_n1862_), .Y(w_mem_inst__abc_21203_new_n1865_));
AND2X2 AND2X2_2871 ( .A(w_mem_inst__abc_21203_new_n1866_), .B(w_mem_inst__abc_21203_new_n1868_), .Y(w_mem_inst__abc_21203_new_n1869_));
AND2X2 AND2X2_2872 ( .A(w_mem_inst__abc_21203_new_n1607_), .B(w_mem_inst_w_mem_5__5_), .Y(w_mem_inst__abc_21203_new_n1871_));
AND2X2 AND2X2_2873 ( .A(w_mem_inst__abc_21203_new_n1614_), .B(w_mem_inst_w_mem_8__5_), .Y(w_mem_inst__abc_21203_new_n1873_));
AND2X2 AND2X2_2874 ( .A(w_mem_inst__abc_21203_new_n1617_), .B(w_mem_inst_w_mem_11__5_), .Y(w_mem_inst__abc_21203_new_n1874_));
AND2X2 AND2X2_2875 ( .A(w_mem_inst__abc_21203_new_n1621_), .B(w_mem_inst_w_mem_7__5_), .Y(w_mem_inst__abc_21203_new_n1877_));
AND2X2 AND2X2_2876 ( .A(w_mem_inst__abc_21203_new_n1624_), .B(w_mem_inst_w_mem_15__5_), .Y(w_mem_inst__abc_21203_new_n1878_));
AND2X2 AND2X2_2877 ( .A(w_mem_inst__abc_21203_new_n1628_), .B(w_mem_inst_w_mem_13__5_), .Y(w_mem_inst__abc_21203_new_n1881_));
AND2X2 AND2X2_2878 ( .A(w_mem_inst__abc_21203_new_n1631_), .B(w_mem_inst_w_mem_0__5_), .Y(w_mem_inst__abc_21203_new_n1882_));
AND2X2 AND2X2_2879 ( .A(w_mem_inst__abc_21203_new_n1633_), .B(w_mem_inst_w_mem_12__5_), .Y(w_mem_inst__abc_21203_new_n1883_));
AND2X2 AND2X2_288 ( .A(_abc_15497_new_n1293_), .B(_abc_15497_new_n1284_), .Y(_abc_15497_new_n1298_));
AND2X2 AND2X2_2880 ( .A(w_mem_inst__abc_21203_new_n1637_), .B(w_mem_inst_w_mem_9__5_), .Y(w_mem_inst__abc_21203_new_n1886_));
AND2X2 AND2X2_2881 ( .A(w_mem_inst__abc_21203_new_n1640_), .B(w_mem_inst_w_mem_10__5_), .Y(w_mem_inst__abc_21203_new_n1887_));
AND2X2 AND2X2_2882 ( .A(w_mem_inst__abc_21203_new_n1643_), .B(w_mem_inst_w_mem_4__5_), .Y(w_mem_inst__abc_21203_new_n1889_));
AND2X2 AND2X2_2883 ( .A(w_mem_inst__abc_21203_new_n1645_), .B(w_mem_inst_w_mem_6__5_), .Y(w_mem_inst__abc_21203_new_n1890_));
AND2X2 AND2X2_2884 ( .A(w_mem_inst__abc_21203_new_n1649_), .B(w_mem_inst_w_mem_1__5_), .Y(w_mem_inst__abc_21203_new_n1893_));
AND2X2 AND2X2_2885 ( .A(w_mem_inst__abc_21203_new_n1651_), .B(w_mem_inst_w_mem_2__5_), .Y(w_mem_inst__abc_21203_new_n1894_));
AND2X2 AND2X2_2886 ( .A(w_mem_inst__abc_21203_new_n1654_), .B(w_mem_inst_w_mem_3__5_), .Y(w_mem_inst__abc_21203_new_n1896_));
AND2X2 AND2X2_2887 ( .A(w_mem_inst__abc_21203_new_n1656_), .B(w_mem_inst_w_mem_14__5_), .Y(w_mem_inst__abc_21203_new_n1897_));
AND2X2 AND2X2_2888 ( .A(w_mem_inst__abc_21203_new_n1902_), .B(w_mem_inst__abc_21203_new_n1870_), .Y(w_5_));
AND2X2 AND2X2_2889 ( .A(w_mem_inst__abc_21203_new_n1905_), .B(w_mem_inst__abc_21203_new_n1907_), .Y(w_mem_inst__abc_21203_new_n1908_));
AND2X2 AND2X2_289 ( .A(e_reg_19_), .B(\digest[19] ), .Y(_abc_15497_new_n1301_));
AND2X2 AND2X2_2890 ( .A(w_mem_inst_w_mem_2__5_), .B(w_mem_inst_w_mem_0__5_), .Y(w_mem_inst__abc_21203_new_n1911_));
AND2X2 AND2X2_2891 ( .A(w_mem_inst__abc_21203_new_n1912_), .B(w_mem_inst__abc_21203_new_n1910_), .Y(w_mem_inst__abc_21203_new_n1913_));
AND2X2 AND2X2_2892 ( .A(w_mem_inst__abc_21203_new_n1914_), .B(w_mem_inst__abc_21203_new_n1916_), .Y(w_mem_inst__abc_21203_new_n1917_));
AND2X2 AND2X2_2893 ( .A(w_mem_inst__abc_21203_new_n1607_), .B(w_mem_inst_w_mem_5__6_), .Y(w_mem_inst__abc_21203_new_n1919_));
AND2X2 AND2X2_2894 ( .A(w_mem_inst__abc_21203_new_n1614_), .B(w_mem_inst_w_mem_8__6_), .Y(w_mem_inst__abc_21203_new_n1921_));
AND2X2 AND2X2_2895 ( .A(w_mem_inst__abc_21203_new_n1617_), .B(w_mem_inst_w_mem_11__6_), .Y(w_mem_inst__abc_21203_new_n1922_));
AND2X2 AND2X2_2896 ( .A(w_mem_inst__abc_21203_new_n1621_), .B(w_mem_inst_w_mem_7__6_), .Y(w_mem_inst__abc_21203_new_n1925_));
AND2X2 AND2X2_2897 ( .A(w_mem_inst__abc_21203_new_n1624_), .B(w_mem_inst_w_mem_15__6_), .Y(w_mem_inst__abc_21203_new_n1926_));
AND2X2 AND2X2_2898 ( .A(w_mem_inst__abc_21203_new_n1628_), .B(w_mem_inst_w_mem_13__6_), .Y(w_mem_inst__abc_21203_new_n1929_));
AND2X2 AND2X2_2899 ( .A(w_mem_inst__abc_21203_new_n1631_), .B(w_mem_inst_w_mem_0__6_), .Y(w_mem_inst__abc_21203_new_n1930_));
AND2X2 AND2X2_29 ( .A(_abc_15497_new_n753_), .B(_abc_15497_new_n730_), .Y(_abc_15497_new_n754_));
AND2X2 AND2X2_290 ( .A(_abc_15497_new_n1302_), .B(_abc_15497_new_n1300_), .Y(_abc_15497_new_n1303_));
AND2X2 AND2X2_2900 ( .A(w_mem_inst__abc_21203_new_n1633_), .B(w_mem_inst_w_mem_12__6_), .Y(w_mem_inst__abc_21203_new_n1931_));
AND2X2 AND2X2_2901 ( .A(w_mem_inst__abc_21203_new_n1637_), .B(w_mem_inst_w_mem_9__6_), .Y(w_mem_inst__abc_21203_new_n1934_));
AND2X2 AND2X2_2902 ( .A(w_mem_inst__abc_21203_new_n1640_), .B(w_mem_inst_w_mem_10__6_), .Y(w_mem_inst__abc_21203_new_n1935_));
AND2X2 AND2X2_2903 ( .A(w_mem_inst__abc_21203_new_n1643_), .B(w_mem_inst_w_mem_4__6_), .Y(w_mem_inst__abc_21203_new_n1937_));
AND2X2 AND2X2_2904 ( .A(w_mem_inst__abc_21203_new_n1645_), .B(w_mem_inst_w_mem_6__6_), .Y(w_mem_inst__abc_21203_new_n1938_));
AND2X2 AND2X2_2905 ( .A(w_mem_inst__abc_21203_new_n1649_), .B(w_mem_inst_w_mem_1__6_), .Y(w_mem_inst__abc_21203_new_n1941_));
AND2X2 AND2X2_2906 ( .A(w_mem_inst__abc_21203_new_n1651_), .B(w_mem_inst_w_mem_2__6_), .Y(w_mem_inst__abc_21203_new_n1942_));
AND2X2 AND2X2_2907 ( .A(w_mem_inst__abc_21203_new_n1654_), .B(w_mem_inst_w_mem_3__6_), .Y(w_mem_inst__abc_21203_new_n1944_));
AND2X2 AND2X2_2908 ( .A(w_mem_inst__abc_21203_new_n1656_), .B(w_mem_inst_w_mem_14__6_), .Y(w_mem_inst__abc_21203_new_n1945_));
AND2X2 AND2X2_2909 ( .A(w_mem_inst__abc_21203_new_n1950_), .B(w_mem_inst__abc_21203_new_n1918_), .Y(w_6_));
AND2X2 AND2X2_291 ( .A(_abc_15497_new_n1306_), .B(digest_update), .Y(_abc_15497_new_n1307_));
AND2X2 AND2X2_2910 ( .A(w_mem_inst__abc_21203_new_n1953_), .B(w_mem_inst__abc_21203_new_n1955_), .Y(w_mem_inst__abc_21203_new_n1956_));
AND2X2 AND2X2_2911 ( .A(w_mem_inst_w_mem_2__6_), .B(w_mem_inst_w_mem_0__6_), .Y(w_mem_inst__abc_21203_new_n1959_));
AND2X2 AND2X2_2912 ( .A(w_mem_inst__abc_21203_new_n1960_), .B(w_mem_inst__abc_21203_new_n1958_), .Y(w_mem_inst__abc_21203_new_n1961_));
AND2X2 AND2X2_2913 ( .A(w_mem_inst__abc_21203_new_n1962_), .B(w_mem_inst__abc_21203_new_n1964_), .Y(w_mem_inst__abc_21203_new_n1965_));
AND2X2 AND2X2_2914 ( .A(w_mem_inst__abc_21203_new_n1607_), .B(w_mem_inst_w_mem_5__7_), .Y(w_mem_inst__abc_21203_new_n1967_));
AND2X2 AND2X2_2915 ( .A(w_mem_inst__abc_21203_new_n1614_), .B(w_mem_inst_w_mem_8__7_), .Y(w_mem_inst__abc_21203_new_n1969_));
AND2X2 AND2X2_2916 ( .A(w_mem_inst__abc_21203_new_n1617_), .B(w_mem_inst_w_mem_11__7_), .Y(w_mem_inst__abc_21203_new_n1970_));
AND2X2 AND2X2_2917 ( .A(w_mem_inst__abc_21203_new_n1621_), .B(w_mem_inst_w_mem_7__7_), .Y(w_mem_inst__abc_21203_new_n1973_));
AND2X2 AND2X2_2918 ( .A(w_mem_inst__abc_21203_new_n1624_), .B(w_mem_inst_w_mem_15__7_), .Y(w_mem_inst__abc_21203_new_n1974_));
AND2X2 AND2X2_2919 ( .A(w_mem_inst__abc_21203_new_n1628_), .B(w_mem_inst_w_mem_13__7_), .Y(w_mem_inst__abc_21203_new_n1977_));
AND2X2 AND2X2_292 ( .A(_abc_15497_new_n1307_), .B(_abc_15497_new_n1304_), .Y(_abc_15497_new_n1308_));
AND2X2 AND2X2_2920 ( .A(w_mem_inst__abc_21203_new_n1631_), .B(w_mem_inst_w_mem_0__7_), .Y(w_mem_inst__abc_21203_new_n1978_));
AND2X2 AND2X2_2921 ( .A(w_mem_inst__abc_21203_new_n1633_), .B(w_mem_inst_w_mem_12__7_), .Y(w_mem_inst__abc_21203_new_n1979_));
AND2X2 AND2X2_2922 ( .A(w_mem_inst__abc_21203_new_n1637_), .B(w_mem_inst_w_mem_9__7_), .Y(w_mem_inst__abc_21203_new_n1982_));
AND2X2 AND2X2_2923 ( .A(w_mem_inst__abc_21203_new_n1640_), .B(w_mem_inst_w_mem_10__7_), .Y(w_mem_inst__abc_21203_new_n1983_));
AND2X2 AND2X2_2924 ( .A(w_mem_inst__abc_21203_new_n1643_), .B(w_mem_inst_w_mem_4__7_), .Y(w_mem_inst__abc_21203_new_n1985_));
AND2X2 AND2X2_2925 ( .A(w_mem_inst__abc_21203_new_n1645_), .B(w_mem_inst_w_mem_6__7_), .Y(w_mem_inst__abc_21203_new_n1986_));
AND2X2 AND2X2_2926 ( .A(w_mem_inst__abc_21203_new_n1649_), .B(w_mem_inst_w_mem_1__7_), .Y(w_mem_inst__abc_21203_new_n1989_));
AND2X2 AND2X2_2927 ( .A(w_mem_inst__abc_21203_new_n1651_), .B(w_mem_inst_w_mem_2__7_), .Y(w_mem_inst__abc_21203_new_n1990_));
AND2X2 AND2X2_2928 ( .A(w_mem_inst__abc_21203_new_n1654_), .B(w_mem_inst_w_mem_3__7_), .Y(w_mem_inst__abc_21203_new_n1992_));
AND2X2 AND2X2_2929 ( .A(w_mem_inst__abc_21203_new_n1656_), .B(w_mem_inst_w_mem_14__7_), .Y(w_mem_inst__abc_21203_new_n1993_));
AND2X2 AND2X2_293 ( .A(_abc_15497_new_n1303_), .B(_abc_15497_new_n1283_), .Y(_abc_15497_new_n1310_));
AND2X2 AND2X2_2930 ( .A(w_mem_inst__abc_21203_new_n1998_), .B(w_mem_inst__abc_21203_new_n1966_), .Y(w_7_));
AND2X2 AND2X2_2931 ( .A(w_mem_inst__abc_21203_new_n2001_), .B(w_mem_inst__abc_21203_new_n2003_), .Y(w_mem_inst__abc_21203_new_n2004_));
AND2X2 AND2X2_2932 ( .A(w_mem_inst_w_mem_2__7_), .B(w_mem_inst_w_mem_0__7_), .Y(w_mem_inst__abc_21203_new_n2007_));
AND2X2 AND2X2_2933 ( .A(w_mem_inst__abc_21203_new_n2008_), .B(w_mem_inst__abc_21203_new_n2006_), .Y(w_mem_inst__abc_21203_new_n2009_));
AND2X2 AND2X2_2934 ( .A(w_mem_inst__abc_21203_new_n2010_), .B(w_mem_inst__abc_21203_new_n2012_), .Y(w_mem_inst__abc_21203_new_n2013_));
AND2X2 AND2X2_2935 ( .A(w_mem_inst__abc_21203_new_n1607_), .B(w_mem_inst_w_mem_5__8_), .Y(w_mem_inst__abc_21203_new_n2015_));
AND2X2 AND2X2_2936 ( .A(w_mem_inst__abc_21203_new_n1614_), .B(w_mem_inst_w_mem_8__8_), .Y(w_mem_inst__abc_21203_new_n2017_));
AND2X2 AND2X2_2937 ( .A(w_mem_inst__abc_21203_new_n1617_), .B(w_mem_inst_w_mem_11__8_), .Y(w_mem_inst__abc_21203_new_n2018_));
AND2X2 AND2X2_2938 ( .A(w_mem_inst__abc_21203_new_n1621_), .B(w_mem_inst_w_mem_7__8_), .Y(w_mem_inst__abc_21203_new_n2021_));
AND2X2 AND2X2_2939 ( .A(w_mem_inst__abc_21203_new_n1624_), .B(w_mem_inst_w_mem_15__8_), .Y(w_mem_inst__abc_21203_new_n2022_));
AND2X2 AND2X2_294 ( .A(_abc_15497_new_n1285_), .B(_abc_15497_new_n1303_), .Y(_abc_15497_new_n1314_));
AND2X2 AND2X2_2940 ( .A(w_mem_inst__abc_21203_new_n1628_), .B(w_mem_inst_w_mem_13__8_), .Y(w_mem_inst__abc_21203_new_n2025_));
AND2X2 AND2X2_2941 ( .A(w_mem_inst__abc_21203_new_n1631_), .B(w_mem_inst_w_mem_0__8_), .Y(w_mem_inst__abc_21203_new_n2026_));
AND2X2 AND2X2_2942 ( .A(w_mem_inst__abc_21203_new_n1633_), .B(w_mem_inst_w_mem_12__8_), .Y(w_mem_inst__abc_21203_new_n2027_));
AND2X2 AND2X2_2943 ( .A(w_mem_inst__abc_21203_new_n1637_), .B(w_mem_inst_w_mem_9__8_), .Y(w_mem_inst__abc_21203_new_n2030_));
AND2X2 AND2X2_2944 ( .A(w_mem_inst__abc_21203_new_n1640_), .B(w_mem_inst_w_mem_10__8_), .Y(w_mem_inst__abc_21203_new_n2031_));
AND2X2 AND2X2_2945 ( .A(w_mem_inst__abc_21203_new_n1643_), .B(w_mem_inst_w_mem_4__8_), .Y(w_mem_inst__abc_21203_new_n2033_));
AND2X2 AND2X2_2946 ( .A(w_mem_inst__abc_21203_new_n1645_), .B(w_mem_inst_w_mem_6__8_), .Y(w_mem_inst__abc_21203_new_n2034_));
AND2X2 AND2X2_2947 ( .A(w_mem_inst__abc_21203_new_n1649_), .B(w_mem_inst_w_mem_1__8_), .Y(w_mem_inst__abc_21203_new_n2037_));
AND2X2 AND2X2_2948 ( .A(w_mem_inst__abc_21203_new_n1651_), .B(w_mem_inst_w_mem_2__8_), .Y(w_mem_inst__abc_21203_new_n2038_));
AND2X2 AND2X2_2949 ( .A(w_mem_inst__abc_21203_new_n1654_), .B(w_mem_inst_w_mem_3__8_), .Y(w_mem_inst__abc_21203_new_n2040_));
AND2X2 AND2X2_295 ( .A(_abc_15497_new_n1316_), .B(_abc_15497_new_n1312_), .Y(_abc_15497_new_n1317_));
AND2X2 AND2X2_2950 ( .A(w_mem_inst__abc_21203_new_n1656_), .B(w_mem_inst_w_mem_14__8_), .Y(w_mem_inst__abc_21203_new_n2041_));
AND2X2 AND2X2_2951 ( .A(w_mem_inst__abc_21203_new_n2046_), .B(w_mem_inst__abc_21203_new_n2014_), .Y(w_8_));
AND2X2 AND2X2_2952 ( .A(w_mem_inst__abc_21203_new_n2049_), .B(w_mem_inst__abc_21203_new_n2051_), .Y(w_mem_inst__abc_21203_new_n2052_));
AND2X2 AND2X2_2953 ( .A(w_mem_inst_w_mem_2__8_), .B(w_mem_inst_w_mem_0__8_), .Y(w_mem_inst__abc_21203_new_n2055_));
AND2X2 AND2X2_2954 ( .A(w_mem_inst__abc_21203_new_n2056_), .B(w_mem_inst__abc_21203_new_n2054_), .Y(w_mem_inst__abc_21203_new_n2057_));
AND2X2 AND2X2_2955 ( .A(w_mem_inst__abc_21203_new_n2058_), .B(w_mem_inst__abc_21203_new_n2060_), .Y(w_mem_inst__abc_21203_new_n2061_));
AND2X2 AND2X2_2956 ( .A(w_mem_inst__abc_21203_new_n1607_), .B(w_mem_inst_w_mem_5__9_), .Y(w_mem_inst__abc_21203_new_n2063_));
AND2X2 AND2X2_2957 ( .A(w_mem_inst__abc_21203_new_n1614_), .B(w_mem_inst_w_mem_8__9_), .Y(w_mem_inst__abc_21203_new_n2065_));
AND2X2 AND2X2_2958 ( .A(w_mem_inst__abc_21203_new_n1617_), .B(w_mem_inst_w_mem_11__9_), .Y(w_mem_inst__abc_21203_new_n2066_));
AND2X2 AND2X2_2959 ( .A(w_mem_inst__abc_21203_new_n1621_), .B(w_mem_inst_w_mem_7__9_), .Y(w_mem_inst__abc_21203_new_n2069_));
AND2X2 AND2X2_296 ( .A(_abc_15497_new_n1260_), .B(_abc_15497_new_n1272_), .Y(_abc_15497_new_n1319_));
AND2X2 AND2X2_2960 ( .A(w_mem_inst__abc_21203_new_n1624_), .B(w_mem_inst_w_mem_15__9_), .Y(w_mem_inst__abc_21203_new_n2070_));
AND2X2 AND2X2_2961 ( .A(w_mem_inst__abc_21203_new_n1628_), .B(w_mem_inst_w_mem_13__9_), .Y(w_mem_inst__abc_21203_new_n2073_));
AND2X2 AND2X2_2962 ( .A(w_mem_inst__abc_21203_new_n1631_), .B(w_mem_inst_w_mem_0__9_), .Y(w_mem_inst__abc_21203_new_n2074_));
AND2X2 AND2X2_2963 ( .A(w_mem_inst__abc_21203_new_n1633_), .B(w_mem_inst_w_mem_12__9_), .Y(w_mem_inst__abc_21203_new_n2075_));
AND2X2 AND2X2_2964 ( .A(w_mem_inst__abc_21203_new_n1637_), .B(w_mem_inst_w_mem_9__9_), .Y(w_mem_inst__abc_21203_new_n2078_));
AND2X2 AND2X2_2965 ( .A(w_mem_inst__abc_21203_new_n1640_), .B(w_mem_inst_w_mem_10__9_), .Y(w_mem_inst__abc_21203_new_n2079_));
AND2X2 AND2X2_2966 ( .A(w_mem_inst__abc_21203_new_n1643_), .B(w_mem_inst_w_mem_4__9_), .Y(w_mem_inst__abc_21203_new_n2081_));
AND2X2 AND2X2_2967 ( .A(w_mem_inst__abc_21203_new_n1645_), .B(w_mem_inst_w_mem_6__9_), .Y(w_mem_inst__abc_21203_new_n2082_));
AND2X2 AND2X2_2968 ( .A(w_mem_inst__abc_21203_new_n1649_), .B(w_mem_inst_w_mem_1__9_), .Y(w_mem_inst__abc_21203_new_n2085_));
AND2X2 AND2X2_2969 ( .A(w_mem_inst__abc_21203_new_n1651_), .B(w_mem_inst_w_mem_2__9_), .Y(w_mem_inst__abc_21203_new_n2086_));
AND2X2 AND2X2_297 ( .A(_abc_15497_new_n1319_), .B(_abc_15497_new_n1314_), .Y(_abc_15497_new_n1320_));
AND2X2 AND2X2_2970 ( .A(w_mem_inst__abc_21203_new_n1654_), .B(w_mem_inst_w_mem_3__9_), .Y(w_mem_inst__abc_21203_new_n2088_));
AND2X2 AND2X2_2971 ( .A(w_mem_inst__abc_21203_new_n1656_), .B(w_mem_inst_w_mem_14__9_), .Y(w_mem_inst__abc_21203_new_n2089_));
AND2X2 AND2X2_2972 ( .A(w_mem_inst__abc_21203_new_n2094_), .B(w_mem_inst__abc_21203_new_n2062_), .Y(w_9_));
AND2X2 AND2X2_2973 ( .A(w_mem_inst__abc_21203_new_n2097_), .B(w_mem_inst__abc_21203_new_n2099_), .Y(w_mem_inst__abc_21203_new_n2100_));
AND2X2 AND2X2_2974 ( .A(w_mem_inst_w_mem_2__9_), .B(w_mem_inst_w_mem_0__9_), .Y(w_mem_inst__abc_21203_new_n2103_));
AND2X2 AND2X2_2975 ( .A(w_mem_inst__abc_21203_new_n2104_), .B(w_mem_inst__abc_21203_new_n2102_), .Y(w_mem_inst__abc_21203_new_n2105_));
AND2X2 AND2X2_2976 ( .A(w_mem_inst__abc_21203_new_n2106_), .B(w_mem_inst__abc_21203_new_n2108_), .Y(w_mem_inst__abc_21203_new_n2109_));
AND2X2 AND2X2_2977 ( .A(w_mem_inst__abc_21203_new_n1607_), .B(w_mem_inst_w_mem_5__10_), .Y(w_mem_inst__abc_21203_new_n2111_));
AND2X2 AND2X2_2978 ( .A(w_mem_inst__abc_21203_new_n1614_), .B(w_mem_inst_w_mem_8__10_), .Y(w_mem_inst__abc_21203_new_n2113_));
AND2X2 AND2X2_2979 ( .A(w_mem_inst__abc_21203_new_n1617_), .B(w_mem_inst_w_mem_11__10_), .Y(w_mem_inst__abc_21203_new_n2114_));
AND2X2 AND2X2_298 ( .A(_abc_15497_new_n1256_), .B(_abc_15497_new_n1320_), .Y(_abc_15497_new_n1321_));
AND2X2 AND2X2_2980 ( .A(w_mem_inst__abc_21203_new_n1621_), .B(w_mem_inst_w_mem_7__10_), .Y(w_mem_inst__abc_21203_new_n2117_));
AND2X2 AND2X2_2981 ( .A(w_mem_inst__abc_21203_new_n1624_), .B(w_mem_inst_w_mem_15__10_), .Y(w_mem_inst__abc_21203_new_n2118_));
AND2X2 AND2X2_2982 ( .A(w_mem_inst__abc_21203_new_n1628_), .B(w_mem_inst_w_mem_13__10_), .Y(w_mem_inst__abc_21203_new_n2121_));
AND2X2 AND2X2_2983 ( .A(w_mem_inst__abc_21203_new_n1631_), .B(w_mem_inst_w_mem_0__10_), .Y(w_mem_inst__abc_21203_new_n2122_));
AND2X2 AND2X2_2984 ( .A(w_mem_inst__abc_21203_new_n1633_), .B(w_mem_inst_w_mem_12__10_), .Y(w_mem_inst__abc_21203_new_n2123_));
AND2X2 AND2X2_2985 ( .A(w_mem_inst__abc_21203_new_n1637_), .B(w_mem_inst_w_mem_9__10_), .Y(w_mem_inst__abc_21203_new_n2126_));
AND2X2 AND2X2_2986 ( .A(w_mem_inst__abc_21203_new_n1640_), .B(w_mem_inst_w_mem_10__10_), .Y(w_mem_inst__abc_21203_new_n2127_));
AND2X2 AND2X2_2987 ( .A(w_mem_inst__abc_21203_new_n1643_), .B(w_mem_inst_w_mem_4__10_), .Y(w_mem_inst__abc_21203_new_n2129_));
AND2X2 AND2X2_2988 ( .A(w_mem_inst__abc_21203_new_n1645_), .B(w_mem_inst_w_mem_6__10_), .Y(w_mem_inst__abc_21203_new_n2130_));
AND2X2 AND2X2_2989 ( .A(w_mem_inst__abc_21203_new_n1649_), .B(w_mem_inst_w_mem_1__10_), .Y(w_mem_inst__abc_21203_new_n2133_));
AND2X2 AND2X2_299 ( .A(e_reg_20_), .B(\digest[20] ), .Y(_abc_15497_new_n1324_));
AND2X2 AND2X2_2990 ( .A(w_mem_inst__abc_21203_new_n1651_), .B(w_mem_inst_w_mem_2__10_), .Y(w_mem_inst__abc_21203_new_n2134_));
AND2X2 AND2X2_2991 ( .A(w_mem_inst__abc_21203_new_n1654_), .B(w_mem_inst_w_mem_3__10_), .Y(w_mem_inst__abc_21203_new_n2136_));
AND2X2 AND2X2_2992 ( .A(w_mem_inst__abc_21203_new_n1656_), .B(w_mem_inst_w_mem_14__10_), .Y(w_mem_inst__abc_21203_new_n2137_));
AND2X2 AND2X2_2993 ( .A(w_mem_inst__abc_21203_new_n2142_), .B(w_mem_inst__abc_21203_new_n2110_), .Y(w_10_));
AND2X2 AND2X2_2994 ( .A(w_mem_inst__abc_21203_new_n2145_), .B(w_mem_inst__abc_21203_new_n2147_), .Y(w_mem_inst__abc_21203_new_n2148_));
AND2X2 AND2X2_2995 ( .A(w_mem_inst_w_mem_2__10_), .B(w_mem_inst_w_mem_0__10_), .Y(w_mem_inst__abc_21203_new_n2151_));
AND2X2 AND2X2_2996 ( .A(w_mem_inst__abc_21203_new_n2152_), .B(w_mem_inst__abc_21203_new_n2150_), .Y(w_mem_inst__abc_21203_new_n2153_));
AND2X2 AND2X2_2997 ( .A(w_mem_inst__abc_21203_new_n2154_), .B(w_mem_inst__abc_21203_new_n2156_), .Y(w_mem_inst__abc_21203_new_n2157_));
AND2X2 AND2X2_2998 ( .A(w_mem_inst__abc_21203_new_n1607_), .B(w_mem_inst_w_mem_5__11_), .Y(w_mem_inst__abc_21203_new_n2159_));
AND2X2 AND2X2_2999 ( .A(w_mem_inst__abc_21203_new_n1614_), .B(w_mem_inst_w_mem_8__11_), .Y(w_mem_inst__abc_21203_new_n2161_));
AND2X2 AND2X2_3 ( .A(_abc_15497_new_n701_), .B(\digest[90] ), .Y(_abc_15497_new_n702_));
AND2X2 AND2X2_30 ( .A(_abc_15497_new_n755_), .B(_abc_15497_new_n726_), .Y(_abc_15497_new_n756_));
AND2X2 AND2X2_300 ( .A(_abc_15497_new_n1325_), .B(_abc_15497_new_n1323_), .Y(_abc_15497_new_n1326_));
AND2X2 AND2X2_3000 ( .A(w_mem_inst__abc_21203_new_n1617_), .B(w_mem_inst_w_mem_11__11_), .Y(w_mem_inst__abc_21203_new_n2162_));
AND2X2 AND2X2_3001 ( .A(w_mem_inst__abc_21203_new_n1621_), .B(w_mem_inst_w_mem_7__11_), .Y(w_mem_inst__abc_21203_new_n2165_));
AND2X2 AND2X2_3002 ( .A(w_mem_inst__abc_21203_new_n1624_), .B(w_mem_inst_w_mem_15__11_), .Y(w_mem_inst__abc_21203_new_n2166_));
AND2X2 AND2X2_3003 ( .A(w_mem_inst__abc_21203_new_n1628_), .B(w_mem_inst_w_mem_13__11_), .Y(w_mem_inst__abc_21203_new_n2169_));
AND2X2 AND2X2_3004 ( .A(w_mem_inst__abc_21203_new_n1631_), .B(w_mem_inst_w_mem_0__11_), .Y(w_mem_inst__abc_21203_new_n2170_));
AND2X2 AND2X2_3005 ( .A(w_mem_inst__abc_21203_new_n1633_), .B(w_mem_inst_w_mem_12__11_), .Y(w_mem_inst__abc_21203_new_n2171_));
AND2X2 AND2X2_3006 ( .A(w_mem_inst__abc_21203_new_n1637_), .B(w_mem_inst_w_mem_9__11_), .Y(w_mem_inst__abc_21203_new_n2174_));
AND2X2 AND2X2_3007 ( .A(w_mem_inst__abc_21203_new_n1640_), .B(w_mem_inst_w_mem_10__11_), .Y(w_mem_inst__abc_21203_new_n2175_));
AND2X2 AND2X2_3008 ( .A(w_mem_inst__abc_21203_new_n1643_), .B(w_mem_inst_w_mem_4__11_), .Y(w_mem_inst__abc_21203_new_n2177_));
AND2X2 AND2X2_3009 ( .A(w_mem_inst__abc_21203_new_n1645_), .B(w_mem_inst_w_mem_6__11_), .Y(w_mem_inst__abc_21203_new_n2178_));
AND2X2 AND2X2_301 ( .A(_abc_15497_new_n1322_), .B(_abc_15497_new_n1326_), .Y(_abc_15497_new_n1328_));
AND2X2 AND2X2_3010 ( .A(w_mem_inst__abc_21203_new_n1649_), .B(w_mem_inst_w_mem_1__11_), .Y(w_mem_inst__abc_21203_new_n2181_));
AND2X2 AND2X2_3011 ( .A(w_mem_inst__abc_21203_new_n1651_), .B(w_mem_inst_w_mem_2__11_), .Y(w_mem_inst__abc_21203_new_n2182_));
AND2X2 AND2X2_3012 ( .A(w_mem_inst__abc_21203_new_n1654_), .B(w_mem_inst_w_mem_3__11_), .Y(w_mem_inst__abc_21203_new_n2184_));
AND2X2 AND2X2_3013 ( .A(w_mem_inst__abc_21203_new_n1656_), .B(w_mem_inst_w_mem_14__11_), .Y(w_mem_inst__abc_21203_new_n2185_));
AND2X2 AND2X2_3014 ( .A(w_mem_inst__abc_21203_new_n2190_), .B(w_mem_inst__abc_21203_new_n2158_), .Y(w_11_));
AND2X2 AND2X2_3015 ( .A(w_mem_inst__abc_21203_new_n2193_), .B(w_mem_inst__abc_21203_new_n2195_), .Y(w_mem_inst__abc_21203_new_n2196_));
AND2X2 AND2X2_3016 ( .A(w_mem_inst_w_mem_2__11_), .B(w_mem_inst_w_mem_0__11_), .Y(w_mem_inst__abc_21203_new_n2199_));
AND2X2 AND2X2_3017 ( .A(w_mem_inst__abc_21203_new_n2200_), .B(w_mem_inst__abc_21203_new_n2198_), .Y(w_mem_inst__abc_21203_new_n2201_));
AND2X2 AND2X2_3018 ( .A(w_mem_inst__abc_21203_new_n2202_), .B(w_mem_inst__abc_21203_new_n2204_), .Y(w_mem_inst__abc_21203_new_n2205_));
AND2X2 AND2X2_3019 ( .A(w_mem_inst__abc_21203_new_n1607_), .B(w_mem_inst_w_mem_5__12_), .Y(w_mem_inst__abc_21203_new_n2207_));
AND2X2 AND2X2_302 ( .A(_abc_15497_new_n1329_), .B(_abc_15497_new_n1327_), .Y(_abc_15497_new_n1330_));
AND2X2 AND2X2_3020 ( .A(w_mem_inst__abc_21203_new_n1614_), .B(w_mem_inst_w_mem_8__12_), .Y(w_mem_inst__abc_21203_new_n2209_));
AND2X2 AND2X2_3021 ( .A(w_mem_inst__abc_21203_new_n1617_), .B(w_mem_inst_w_mem_11__12_), .Y(w_mem_inst__abc_21203_new_n2210_));
AND2X2 AND2X2_3022 ( .A(w_mem_inst__abc_21203_new_n1621_), .B(w_mem_inst_w_mem_7__12_), .Y(w_mem_inst__abc_21203_new_n2213_));
AND2X2 AND2X2_3023 ( .A(w_mem_inst__abc_21203_new_n1624_), .B(w_mem_inst_w_mem_15__12_), .Y(w_mem_inst__abc_21203_new_n2214_));
AND2X2 AND2X2_3024 ( .A(w_mem_inst__abc_21203_new_n1628_), .B(w_mem_inst_w_mem_13__12_), .Y(w_mem_inst__abc_21203_new_n2217_));
AND2X2 AND2X2_3025 ( .A(w_mem_inst__abc_21203_new_n1631_), .B(w_mem_inst_w_mem_0__12_), .Y(w_mem_inst__abc_21203_new_n2218_));
AND2X2 AND2X2_3026 ( .A(w_mem_inst__abc_21203_new_n1633_), .B(w_mem_inst_w_mem_12__12_), .Y(w_mem_inst__abc_21203_new_n2219_));
AND2X2 AND2X2_3027 ( .A(w_mem_inst__abc_21203_new_n1637_), .B(w_mem_inst_w_mem_9__12_), .Y(w_mem_inst__abc_21203_new_n2222_));
AND2X2 AND2X2_3028 ( .A(w_mem_inst__abc_21203_new_n1640_), .B(w_mem_inst_w_mem_10__12_), .Y(w_mem_inst__abc_21203_new_n2223_));
AND2X2 AND2X2_3029 ( .A(w_mem_inst__abc_21203_new_n1643_), .B(w_mem_inst_w_mem_4__12_), .Y(w_mem_inst__abc_21203_new_n2225_));
AND2X2 AND2X2_303 ( .A(_abc_15497_new_n1330_), .B(digest_update), .Y(_abc_15497_new_n1331_));
AND2X2 AND2X2_3030 ( .A(w_mem_inst__abc_21203_new_n1645_), .B(w_mem_inst_w_mem_6__12_), .Y(w_mem_inst__abc_21203_new_n2226_));
AND2X2 AND2X2_3031 ( .A(w_mem_inst__abc_21203_new_n1649_), .B(w_mem_inst_w_mem_1__12_), .Y(w_mem_inst__abc_21203_new_n2229_));
AND2X2 AND2X2_3032 ( .A(w_mem_inst__abc_21203_new_n1651_), .B(w_mem_inst_w_mem_2__12_), .Y(w_mem_inst__abc_21203_new_n2230_));
AND2X2 AND2X2_3033 ( .A(w_mem_inst__abc_21203_new_n1654_), .B(w_mem_inst_w_mem_3__12_), .Y(w_mem_inst__abc_21203_new_n2232_));
AND2X2 AND2X2_3034 ( .A(w_mem_inst__abc_21203_new_n1656_), .B(w_mem_inst_w_mem_14__12_), .Y(w_mem_inst__abc_21203_new_n2233_));
AND2X2 AND2X2_3035 ( .A(w_mem_inst__abc_21203_new_n2238_), .B(w_mem_inst__abc_21203_new_n2206_), .Y(w_12_));
AND2X2 AND2X2_3036 ( .A(w_mem_inst__abc_21203_new_n2241_), .B(w_mem_inst__abc_21203_new_n2243_), .Y(w_mem_inst__abc_21203_new_n2244_));
AND2X2 AND2X2_3037 ( .A(w_mem_inst_w_mem_2__12_), .B(w_mem_inst_w_mem_0__12_), .Y(w_mem_inst__abc_21203_new_n2247_));
AND2X2 AND2X2_3038 ( .A(w_mem_inst__abc_21203_new_n2248_), .B(w_mem_inst__abc_21203_new_n2246_), .Y(w_mem_inst__abc_21203_new_n2249_));
AND2X2 AND2X2_3039 ( .A(w_mem_inst__abc_21203_new_n2250_), .B(w_mem_inst__abc_21203_new_n2252_), .Y(w_mem_inst__abc_21203_new_n2253_));
AND2X2 AND2X2_304 ( .A(_abc_15497_new_n1332_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n1333_));
AND2X2 AND2X2_3040 ( .A(w_mem_inst__abc_21203_new_n1607_), .B(w_mem_inst_w_mem_5__13_), .Y(w_mem_inst__abc_21203_new_n2255_));
AND2X2 AND2X2_3041 ( .A(w_mem_inst__abc_21203_new_n1614_), .B(w_mem_inst_w_mem_8__13_), .Y(w_mem_inst__abc_21203_new_n2257_));
AND2X2 AND2X2_3042 ( .A(w_mem_inst__abc_21203_new_n1617_), .B(w_mem_inst_w_mem_11__13_), .Y(w_mem_inst__abc_21203_new_n2258_));
AND2X2 AND2X2_3043 ( .A(w_mem_inst__abc_21203_new_n1621_), .B(w_mem_inst_w_mem_7__13_), .Y(w_mem_inst__abc_21203_new_n2261_));
AND2X2 AND2X2_3044 ( .A(w_mem_inst__abc_21203_new_n1624_), .B(w_mem_inst_w_mem_15__13_), .Y(w_mem_inst__abc_21203_new_n2262_));
AND2X2 AND2X2_3045 ( .A(w_mem_inst__abc_21203_new_n1628_), .B(w_mem_inst_w_mem_13__13_), .Y(w_mem_inst__abc_21203_new_n2265_));
AND2X2 AND2X2_3046 ( .A(w_mem_inst__abc_21203_new_n1631_), .B(w_mem_inst_w_mem_0__13_), .Y(w_mem_inst__abc_21203_new_n2266_));
AND2X2 AND2X2_3047 ( .A(w_mem_inst__abc_21203_new_n1633_), .B(w_mem_inst_w_mem_12__13_), .Y(w_mem_inst__abc_21203_new_n2267_));
AND2X2 AND2X2_3048 ( .A(w_mem_inst__abc_21203_new_n1637_), .B(w_mem_inst_w_mem_9__13_), .Y(w_mem_inst__abc_21203_new_n2270_));
AND2X2 AND2X2_3049 ( .A(w_mem_inst__abc_21203_new_n1640_), .B(w_mem_inst_w_mem_10__13_), .Y(w_mem_inst__abc_21203_new_n2271_));
AND2X2 AND2X2_305 ( .A(_abc_15497_new_n701_), .B(\digest[21] ), .Y(_abc_15497_new_n1335_));
AND2X2 AND2X2_3050 ( .A(w_mem_inst__abc_21203_new_n1643_), .B(w_mem_inst_w_mem_4__13_), .Y(w_mem_inst__abc_21203_new_n2273_));
AND2X2 AND2X2_3051 ( .A(w_mem_inst__abc_21203_new_n1645_), .B(w_mem_inst_w_mem_6__13_), .Y(w_mem_inst__abc_21203_new_n2274_));
AND2X2 AND2X2_3052 ( .A(w_mem_inst__abc_21203_new_n1649_), .B(w_mem_inst_w_mem_1__13_), .Y(w_mem_inst__abc_21203_new_n2277_));
AND2X2 AND2X2_3053 ( .A(w_mem_inst__abc_21203_new_n1651_), .B(w_mem_inst_w_mem_2__13_), .Y(w_mem_inst__abc_21203_new_n2278_));
AND2X2 AND2X2_3054 ( .A(w_mem_inst__abc_21203_new_n1654_), .B(w_mem_inst_w_mem_3__13_), .Y(w_mem_inst__abc_21203_new_n2280_));
AND2X2 AND2X2_3055 ( .A(w_mem_inst__abc_21203_new_n1656_), .B(w_mem_inst_w_mem_14__13_), .Y(w_mem_inst__abc_21203_new_n2281_));
AND2X2 AND2X2_3056 ( .A(w_mem_inst__abc_21203_new_n2286_), .B(w_mem_inst__abc_21203_new_n2254_), .Y(w_13_));
AND2X2 AND2X2_3057 ( .A(w_mem_inst__abc_21203_new_n2289_), .B(w_mem_inst__abc_21203_new_n2291_), .Y(w_mem_inst__abc_21203_new_n2292_));
AND2X2 AND2X2_3058 ( .A(w_mem_inst_w_mem_2__13_), .B(w_mem_inst_w_mem_0__13_), .Y(w_mem_inst__abc_21203_new_n2295_));
AND2X2 AND2X2_3059 ( .A(w_mem_inst__abc_21203_new_n2296_), .B(w_mem_inst__abc_21203_new_n2294_), .Y(w_mem_inst__abc_21203_new_n2297_));
AND2X2 AND2X2_306 ( .A(e_reg_21_), .B(\digest[21] ), .Y(_abc_15497_new_n1337_));
AND2X2 AND2X2_3060 ( .A(w_mem_inst__abc_21203_new_n2298_), .B(w_mem_inst__abc_21203_new_n2300_), .Y(w_mem_inst__abc_21203_new_n2301_));
AND2X2 AND2X2_3061 ( .A(w_mem_inst__abc_21203_new_n1607_), .B(w_mem_inst_w_mem_5__14_), .Y(w_mem_inst__abc_21203_new_n2303_));
AND2X2 AND2X2_3062 ( .A(w_mem_inst__abc_21203_new_n1614_), .B(w_mem_inst_w_mem_8__14_), .Y(w_mem_inst__abc_21203_new_n2305_));
AND2X2 AND2X2_3063 ( .A(w_mem_inst__abc_21203_new_n1617_), .B(w_mem_inst_w_mem_11__14_), .Y(w_mem_inst__abc_21203_new_n2306_));
AND2X2 AND2X2_3064 ( .A(w_mem_inst__abc_21203_new_n1621_), .B(w_mem_inst_w_mem_7__14_), .Y(w_mem_inst__abc_21203_new_n2309_));
AND2X2 AND2X2_3065 ( .A(w_mem_inst__abc_21203_new_n1624_), .B(w_mem_inst_w_mem_15__14_), .Y(w_mem_inst__abc_21203_new_n2310_));
AND2X2 AND2X2_3066 ( .A(w_mem_inst__abc_21203_new_n1628_), .B(w_mem_inst_w_mem_13__14_), .Y(w_mem_inst__abc_21203_new_n2313_));
AND2X2 AND2X2_3067 ( .A(w_mem_inst__abc_21203_new_n1631_), .B(w_mem_inst_w_mem_0__14_), .Y(w_mem_inst__abc_21203_new_n2314_));
AND2X2 AND2X2_3068 ( .A(w_mem_inst__abc_21203_new_n1633_), .B(w_mem_inst_w_mem_12__14_), .Y(w_mem_inst__abc_21203_new_n2315_));
AND2X2 AND2X2_3069 ( .A(w_mem_inst__abc_21203_new_n1637_), .B(w_mem_inst_w_mem_9__14_), .Y(w_mem_inst__abc_21203_new_n2318_));
AND2X2 AND2X2_307 ( .A(_abc_15497_new_n1338_), .B(_abc_15497_new_n1336_), .Y(_abc_15497_new_n1339_));
AND2X2 AND2X2_3070 ( .A(w_mem_inst__abc_21203_new_n1640_), .B(w_mem_inst_w_mem_10__14_), .Y(w_mem_inst__abc_21203_new_n2319_));
AND2X2 AND2X2_3071 ( .A(w_mem_inst__abc_21203_new_n1643_), .B(w_mem_inst_w_mem_4__14_), .Y(w_mem_inst__abc_21203_new_n2321_));
AND2X2 AND2X2_3072 ( .A(w_mem_inst__abc_21203_new_n1645_), .B(w_mem_inst_w_mem_6__14_), .Y(w_mem_inst__abc_21203_new_n2322_));
AND2X2 AND2X2_3073 ( .A(w_mem_inst__abc_21203_new_n1649_), .B(w_mem_inst_w_mem_1__14_), .Y(w_mem_inst__abc_21203_new_n2325_));
AND2X2 AND2X2_3074 ( .A(w_mem_inst__abc_21203_new_n1651_), .B(w_mem_inst_w_mem_2__14_), .Y(w_mem_inst__abc_21203_new_n2326_));
AND2X2 AND2X2_3075 ( .A(w_mem_inst__abc_21203_new_n1654_), .B(w_mem_inst_w_mem_3__14_), .Y(w_mem_inst__abc_21203_new_n2328_));
AND2X2 AND2X2_3076 ( .A(w_mem_inst__abc_21203_new_n1656_), .B(w_mem_inst_w_mem_14__14_), .Y(w_mem_inst__abc_21203_new_n2329_));
AND2X2 AND2X2_3077 ( .A(w_mem_inst__abc_21203_new_n2334_), .B(w_mem_inst__abc_21203_new_n2302_), .Y(w_14_));
AND2X2 AND2X2_3078 ( .A(w_mem_inst__abc_21203_new_n2337_), .B(w_mem_inst__abc_21203_new_n2339_), .Y(w_mem_inst__abc_21203_new_n2340_));
AND2X2 AND2X2_3079 ( .A(w_mem_inst_w_mem_2__14_), .B(w_mem_inst_w_mem_0__14_), .Y(w_mem_inst__abc_21203_new_n2343_));
AND2X2 AND2X2_308 ( .A(_abc_15497_new_n1326_), .B(_abc_15497_new_n1339_), .Y(_abc_15497_new_n1342_));
AND2X2 AND2X2_3080 ( .A(w_mem_inst__abc_21203_new_n2344_), .B(w_mem_inst__abc_21203_new_n2342_), .Y(w_mem_inst__abc_21203_new_n2345_));
AND2X2 AND2X2_3081 ( .A(w_mem_inst__abc_21203_new_n2346_), .B(w_mem_inst__abc_21203_new_n2348_), .Y(w_mem_inst__abc_21203_new_n2349_));
AND2X2 AND2X2_3082 ( .A(w_mem_inst__abc_21203_new_n1607_), .B(w_mem_inst_w_mem_5__15_), .Y(w_mem_inst__abc_21203_new_n2351_));
AND2X2 AND2X2_3083 ( .A(w_mem_inst__abc_21203_new_n1614_), .B(w_mem_inst_w_mem_8__15_), .Y(w_mem_inst__abc_21203_new_n2353_));
AND2X2 AND2X2_3084 ( .A(w_mem_inst__abc_21203_new_n1617_), .B(w_mem_inst_w_mem_11__15_), .Y(w_mem_inst__abc_21203_new_n2354_));
AND2X2 AND2X2_3085 ( .A(w_mem_inst__abc_21203_new_n1621_), .B(w_mem_inst_w_mem_7__15_), .Y(w_mem_inst__abc_21203_new_n2357_));
AND2X2 AND2X2_3086 ( .A(w_mem_inst__abc_21203_new_n1624_), .B(w_mem_inst_w_mem_15__15_), .Y(w_mem_inst__abc_21203_new_n2358_));
AND2X2 AND2X2_3087 ( .A(w_mem_inst__abc_21203_new_n1628_), .B(w_mem_inst_w_mem_13__15_), .Y(w_mem_inst__abc_21203_new_n2361_));
AND2X2 AND2X2_3088 ( .A(w_mem_inst__abc_21203_new_n1631_), .B(w_mem_inst_w_mem_0__15_), .Y(w_mem_inst__abc_21203_new_n2362_));
AND2X2 AND2X2_3089 ( .A(w_mem_inst__abc_21203_new_n1633_), .B(w_mem_inst_w_mem_12__15_), .Y(w_mem_inst__abc_21203_new_n2363_));
AND2X2 AND2X2_309 ( .A(_abc_15497_new_n1322_), .B(_abc_15497_new_n1342_), .Y(_abc_15497_new_n1343_));
AND2X2 AND2X2_3090 ( .A(w_mem_inst__abc_21203_new_n1637_), .B(w_mem_inst_w_mem_9__15_), .Y(w_mem_inst__abc_21203_new_n2366_));
AND2X2 AND2X2_3091 ( .A(w_mem_inst__abc_21203_new_n1640_), .B(w_mem_inst_w_mem_10__15_), .Y(w_mem_inst__abc_21203_new_n2367_));
AND2X2 AND2X2_3092 ( .A(w_mem_inst__abc_21203_new_n1643_), .B(w_mem_inst_w_mem_4__15_), .Y(w_mem_inst__abc_21203_new_n2369_));
AND2X2 AND2X2_3093 ( .A(w_mem_inst__abc_21203_new_n1645_), .B(w_mem_inst_w_mem_6__15_), .Y(w_mem_inst__abc_21203_new_n2370_));
AND2X2 AND2X2_3094 ( .A(w_mem_inst__abc_21203_new_n1649_), .B(w_mem_inst_w_mem_1__15_), .Y(w_mem_inst__abc_21203_new_n2373_));
AND2X2 AND2X2_3095 ( .A(w_mem_inst__abc_21203_new_n1651_), .B(w_mem_inst_w_mem_2__15_), .Y(w_mem_inst__abc_21203_new_n2374_));
AND2X2 AND2X2_3096 ( .A(w_mem_inst__abc_21203_new_n1654_), .B(w_mem_inst_w_mem_3__15_), .Y(w_mem_inst__abc_21203_new_n2376_));
AND2X2 AND2X2_3097 ( .A(w_mem_inst__abc_21203_new_n1656_), .B(w_mem_inst_w_mem_14__15_), .Y(w_mem_inst__abc_21203_new_n2377_));
AND2X2 AND2X2_3098 ( .A(w_mem_inst__abc_21203_new_n2382_), .B(w_mem_inst__abc_21203_new_n2350_), .Y(w_15_));
AND2X2 AND2X2_3099 ( .A(w_mem_inst__abc_21203_new_n2385_), .B(w_mem_inst__abc_21203_new_n2387_), .Y(w_mem_inst__abc_21203_new_n2388_));
AND2X2 AND2X2_31 ( .A(c_reg_15_), .B(\digest[79] ), .Y(_abc_15497_new_n758_));
AND2X2 AND2X2_310 ( .A(_abc_15497_new_n1339_), .B(_abc_15497_new_n1324_), .Y(_abc_15497_new_n1345_));
AND2X2 AND2X2_3100 ( .A(w_mem_inst_w_mem_2__15_), .B(w_mem_inst_w_mem_0__15_), .Y(w_mem_inst__abc_21203_new_n2391_));
AND2X2 AND2X2_3101 ( .A(w_mem_inst__abc_21203_new_n2392_), .B(w_mem_inst__abc_21203_new_n2390_), .Y(w_mem_inst__abc_21203_new_n2393_));
AND2X2 AND2X2_3102 ( .A(w_mem_inst__abc_21203_new_n2394_), .B(w_mem_inst__abc_21203_new_n2396_), .Y(w_mem_inst__abc_21203_new_n2397_));
AND2X2 AND2X2_3103 ( .A(w_mem_inst__abc_21203_new_n1607_), .B(w_mem_inst_w_mem_5__16_), .Y(w_mem_inst__abc_21203_new_n2399_));
AND2X2 AND2X2_3104 ( .A(w_mem_inst__abc_21203_new_n1614_), .B(w_mem_inst_w_mem_8__16_), .Y(w_mem_inst__abc_21203_new_n2401_));
AND2X2 AND2X2_3105 ( .A(w_mem_inst__abc_21203_new_n1617_), .B(w_mem_inst_w_mem_11__16_), .Y(w_mem_inst__abc_21203_new_n2402_));
AND2X2 AND2X2_3106 ( .A(w_mem_inst__abc_21203_new_n1621_), .B(w_mem_inst_w_mem_7__16_), .Y(w_mem_inst__abc_21203_new_n2405_));
AND2X2 AND2X2_3107 ( .A(w_mem_inst__abc_21203_new_n1624_), .B(w_mem_inst_w_mem_15__16_), .Y(w_mem_inst__abc_21203_new_n2406_));
AND2X2 AND2X2_3108 ( .A(w_mem_inst__abc_21203_new_n1628_), .B(w_mem_inst_w_mem_13__16_), .Y(w_mem_inst__abc_21203_new_n2409_));
AND2X2 AND2X2_3109 ( .A(w_mem_inst__abc_21203_new_n1631_), .B(w_mem_inst_w_mem_0__16_), .Y(w_mem_inst__abc_21203_new_n2410_));
AND2X2 AND2X2_311 ( .A(_abc_15497_new_n1346_), .B(digest_update), .Y(_abc_15497_new_n1347_));
AND2X2 AND2X2_3110 ( .A(w_mem_inst__abc_21203_new_n1633_), .B(w_mem_inst_w_mem_12__16_), .Y(w_mem_inst__abc_21203_new_n2411_));
AND2X2 AND2X2_3111 ( .A(w_mem_inst__abc_21203_new_n1637_), .B(w_mem_inst_w_mem_9__16_), .Y(w_mem_inst__abc_21203_new_n2414_));
AND2X2 AND2X2_3112 ( .A(w_mem_inst__abc_21203_new_n1640_), .B(w_mem_inst_w_mem_10__16_), .Y(w_mem_inst__abc_21203_new_n2415_));
AND2X2 AND2X2_3113 ( .A(w_mem_inst__abc_21203_new_n1643_), .B(w_mem_inst_w_mem_4__16_), .Y(w_mem_inst__abc_21203_new_n2417_));
AND2X2 AND2X2_3114 ( .A(w_mem_inst__abc_21203_new_n1645_), .B(w_mem_inst_w_mem_6__16_), .Y(w_mem_inst__abc_21203_new_n2418_));
AND2X2 AND2X2_3115 ( .A(w_mem_inst__abc_21203_new_n1649_), .B(w_mem_inst_w_mem_1__16_), .Y(w_mem_inst__abc_21203_new_n2421_));
AND2X2 AND2X2_3116 ( .A(w_mem_inst__abc_21203_new_n1651_), .B(w_mem_inst_w_mem_2__16_), .Y(w_mem_inst__abc_21203_new_n2422_));
AND2X2 AND2X2_3117 ( .A(w_mem_inst__abc_21203_new_n1654_), .B(w_mem_inst_w_mem_3__16_), .Y(w_mem_inst__abc_21203_new_n2424_));
AND2X2 AND2X2_3118 ( .A(w_mem_inst__abc_21203_new_n1656_), .B(w_mem_inst_w_mem_14__16_), .Y(w_mem_inst__abc_21203_new_n2425_));
AND2X2 AND2X2_3119 ( .A(w_mem_inst__abc_21203_new_n2430_), .B(w_mem_inst__abc_21203_new_n2398_), .Y(w_16_));
AND2X2 AND2X2_312 ( .A(_abc_15497_new_n1344_), .B(_abc_15497_new_n1347_), .Y(_abc_15497_new_n1348_));
AND2X2 AND2X2_3120 ( .A(w_mem_inst__abc_21203_new_n2433_), .B(w_mem_inst__abc_21203_new_n2435_), .Y(w_mem_inst__abc_21203_new_n2436_));
AND2X2 AND2X2_3121 ( .A(w_mem_inst_w_mem_2__16_), .B(w_mem_inst_w_mem_0__16_), .Y(w_mem_inst__abc_21203_new_n2439_));
AND2X2 AND2X2_3122 ( .A(w_mem_inst__abc_21203_new_n2440_), .B(w_mem_inst__abc_21203_new_n2438_), .Y(w_mem_inst__abc_21203_new_n2441_));
AND2X2 AND2X2_3123 ( .A(w_mem_inst__abc_21203_new_n2442_), .B(w_mem_inst__abc_21203_new_n2444_), .Y(w_mem_inst__abc_21203_new_n2445_));
AND2X2 AND2X2_3124 ( .A(w_mem_inst__abc_21203_new_n1607_), .B(w_mem_inst_w_mem_5__17_), .Y(w_mem_inst__abc_21203_new_n2447_));
AND2X2 AND2X2_3125 ( .A(w_mem_inst__abc_21203_new_n1614_), .B(w_mem_inst_w_mem_8__17_), .Y(w_mem_inst__abc_21203_new_n2449_));
AND2X2 AND2X2_3126 ( .A(w_mem_inst__abc_21203_new_n1617_), .B(w_mem_inst_w_mem_11__17_), .Y(w_mem_inst__abc_21203_new_n2450_));
AND2X2 AND2X2_3127 ( .A(w_mem_inst__abc_21203_new_n1621_), .B(w_mem_inst_w_mem_7__17_), .Y(w_mem_inst__abc_21203_new_n2453_));
AND2X2 AND2X2_3128 ( .A(w_mem_inst__abc_21203_new_n1624_), .B(w_mem_inst_w_mem_15__17_), .Y(w_mem_inst__abc_21203_new_n2454_));
AND2X2 AND2X2_3129 ( .A(w_mem_inst__abc_21203_new_n1628_), .B(w_mem_inst_w_mem_13__17_), .Y(w_mem_inst__abc_21203_new_n2457_));
AND2X2 AND2X2_313 ( .A(_abc_15497_new_n1348_), .B(_abc_15497_new_n1341_), .Y(_abc_15497_new_n1349_));
AND2X2 AND2X2_3130 ( .A(w_mem_inst__abc_21203_new_n1631_), .B(w_mem_inst_w_mem_0__17_), .Y(w_mem_inst__abc_21203_new_n2458_));
AND2X2 AND2X2_3131 ( .A(w_mem_inst__abc_21203_new_n1633_), .B(w_mem_inst_w_mem_12__17_), .Y(w_mem_inst__abc_21203_new_n2459_));
AND2X2 AND2X2_3132 ( .A(w_mem_inst__abc_21203_new_n1637_), .B(w_mem_inst_w_mem_9__17_), .Y(w_mem_inst__abc_21203_new_n2462_));
AND2X2 AND2X2_3133 ( .A(w_mem_inst__abc_21203_new_n1640_), .B(w_mem_inst_w_mem_10__17_), .Y(w_mem_inst__abc_21203_new_n2463_));
AND2X2 AND2X2_3134 ( .A(w_mem_inst__abc_21203_new_n1643_), .B(w_mem_inst_w_mem_4__17_), .Y(w_mem_inst__abc_21203_new_n2465_));
AND2X2 AND2X2_3135 ( .A(w_mem_inst__abc_21203_new_n1645_), .B(w_mem_inst_w_mem_6__17_), .Y(w_mem_inst__abc_21203_new_n2466_));
AND2X2 AND2X2_3136 ( .A(w_mem_inst__abc_21203_new_n1649_), .B(w_mem_inst_w_mem_1__17_), .Y(w_mem_inst__abc_21203_new_n2469_));
AND2X2 AND2X2_3137 ( .A(w_mem_inst__abc_21203_new_n1651_), .B(w_mem_inst_w_mem_2__17_), .Y(w_mem_inst__abc_21203_new_n2470_));
AND2X2 AND2X2_3138 ( .A(w_mem_inst__abc_21203_new_n1654_), .B(w_mem_inst_w_mem_3__17_), .Y(w_mem_inst__abc_21203_new_n2472_));
AND2X2 AND2X2_3139 ( .A(w_mem_inst__abc_21203_new_n1656_), .B(w_mem_inst_w_mem_14__17_), .Y(w_mem_inst__abc_21203_new_n2473_));
AND2X2 AND2X2_314 ( .A(_abc_15497_new_n1346_), .B(_abc_15497_new_n1338_), .Y(_abc_15497_new_n1351_));
AND2X2 AND2X2_3140 ( .A(w_mem_inst__abc_21203_new_n2478_), .B(w_mem_inst__abc_21203_new_n2446_), .Y(w_17_));
AND2X2 AND2X2_3141 ( .A(w_mem_inst__abc_21203_new_n2481_), .B(w_mem_inst__abc_21203_new_n2483_), .Y(w_mem_inst__abc_21203_new_n2484_));
AND2X2 AND2X2_3142 ( .A(w_mem_inst_w_mem_2__17_), .B(w_mem_inst_w_mem_0__17_), .Y(w_mem_inst__abc_21203_new_n2487_));
AND2X2 AND2X2_3143 ( .A(w_mem_inst__abc_21203_new_n2488_), .B(w_mem_inst__abc_21203_new_n2486_), .Y(w_mem_inst__abc_21203_new_n2489_));
AND2X2 AND2X2_3144 ( .A(w_mem_inst__abc_21203_new_n2490_), .B(w_mem_inst__abc_21203_new_n2492_), .Y(w_mem_inst__abc_21203_new_n2493_));
AND2X2 AND2X2_3145 ( .A(w_mem_inst__abc_21203_new_n1607_), .B(w_mem_inst_w_mem_5__18_), .Y(w_mem_inst__abc_21203_new_n2495_));
AND2X2 AND2X2_3146 ( .A(w_mem_inst__abc_21203_new_n1614_), .B(w_mem_inst_w_mem_8__18_), .Y(w_mem_inst__abc_21203_new_n2497_));
AND2X2 AND2X2_3147 ( .A(w_mem_inst__abc_21203_new_n1617_), .B(w_mem_inst_w_mem_11__18_), .Y(w_mem_inst__abc_21203_new_n2498_));
AND2X2 AND2X2_3148 ( .A(w_mem_inst__abc_21203_new_n1621_), .B(w_mem_inst_w_mem_7__18_), .Y(w_mem_inst__abc_21203_new_n2501_));
AND2X2 AND2X2_3149 ( .A(w_mem_inst__abc_21203_new_n1624_), .B(w_mem_inst_w_mem_15__18_), .Y(w_mem_inst__abc_21203_new_n2502_));
AND2X2 AND2X2_315 ( .A(_abc_15497_new_n1344_), .B(_abc_15497_new_n1351_), .Y(_abc_15497_new_n1352_));
AND2X2 AND2X2_3150 ( .A(w_mem_inst__abc_21203_new_n1628_), .B(w_mem_inst_w_mem_13__18_), .Y(w_mem_inst__abc_21203_new_n2505_));
AND2X2 AND2X2_3151 ( .A(w_mem_inst__abc_21203_new_n1631_), .B(w_mem_inst_w_mem_0__18_), .Y(w_mem_inst__abc_21203_new_n2506_));
AND2X2 AND2X2_3152 ( .A(w_mem_inst__abc_21203_new_n1633_), .B(w_mem_inst_w_mem_12__18_), .Y(w_mem_inst__abc_21203_new_n2507_));
AND2X2 AND2X2_3153 ( .A(w_mem_inst__abc_21203_new_n1637_), .B(w_mem_inst_w_mem_9__18_), .Y(w_mem_inst__abc_21203_new_n2510_));
AND2X2 AND2X2_3154 ( .A(w_mem_inst__abc_21203_new_n1640_), .B(w_mem_inst_w_mem_10__18_), .Y(w_mem_inst__abc_21203_new_n2511_));
AND2X2 AND2X2_3155 ( .A(w_mem_inst__abc_21203_new_n1643_), .B(w_mem_inst_w_mem_4__18_), .Y(w_mem_inst__abc_21203_new_n2513_));
AND2X2 AND2X2_3156 ( .A(w_mem_inst__abc_21203_new_n1645_), .B(w_mem_inst_w_mem_6__18_), .Y(w_mem_inst__abc_21203_new_n2514_));
AND2X2 AND2X2_3157 ( .A(w_mem_inst__abc_21203_new_n1649_), .B(w_mem_inst_w_mem_1__18_), .Y(w_mem_inst__abc_21203_new_n2517_));
AND2X2 AND2X2_3158 ( .A(w_mem_inst__abc_21203_new_n1651_), .B(w_mem_inst_w_mem_2__18_), .Y(w_mem_inst__abc_21203_new_n2518_));
AND2X2 AND2X2_3159 ( .A(w_mem_inst__abc_21203_new_n1654_), .B(w_mem_inst_w_mem_3__18_), .Y(w_mem_inst__abc_21203_new_n2520_));
AND2X2 AND2X2_316 ( .A(e_reg_22_), .B(\digest[22] ), .Y(_abc_15497_new_n1355_));
AND2X2 AND2X2_3160 ( .A(w_mem_inst__abc_21203_new_n1656_), .B(w_mem_inst_w_mem_14__18_), .Y(w_mem_inst__abc_21203_new_n2521_));
AND2X2 AND2X2_3161 ( .A(w_mem_inst__abc_21203_new_n2526_), .B(w_mem_inst__abc_21203_new_n2494_), .Y(w_18_));
AND2X2 AND2X2_3162 ( .A(w_mem_inst__abc_21203_new_n2529_), .B(w_mem_inst__abc_21203_new_n2531_), .Y(w_mem_inst__abc_21203_new_n2532_));
AND2X2 AND2X2_3163 ( .A(w_mem_inst_w_mem_2__18_), .B(w_mem_inst_w_mem_0__18_), .Y(w_mem_inst__abc_21203_new_n2535_));
AND2X2 AND2X2_3164 ( .A(w_mem_inst__abc_21203_new_n2536_), .B(w_mem_inst__abc_21203_new_n2534_), .Y(w_mem_inst__abc_21203_new_n2537_));
AND2X2 AND2X2_3165 ( .A(w_mem_inst__abc_21203_new_n2538_), .B(w_mem_inst__abc_21203_new_n2540_), .Y(w_mem_inst__abc_21203_new_n2541_));
AND2X2 AND2X2_3166 ( .A(w_mem_inst__abc_21203_new_n1607_), .B(w_mem_inst_w_mem_5__19_), .Y(w_mem_inst__abc_21203_new_n2543_));
AND2X2 AND2X2_3167 ( .A(w_mem_inst__abc_21203_new_n1614_), .B(w_mem_inst_w_mem_8__19_), .Y(w_mem_inst__abc_21203_new_n2545_));
AND2X2 AND2X2_3168 ( .A(w_mem_inst__abc_21203_new_n1617_), .B(w_mem_inst_w_mem_11__19_), .Y(w_mem_inst__abc_21203_new_n2546_));
AND2X2 AND2X2_3169 ( .A(w_mem_inst__abc_21203_new_n1621_), .B(w_mem_inst_w_mem_7__19_), .Y(w_mem_inst__abc_21203_new_n2549_));
AND2X2 AND2X2_317 ( .A(_abc_15497_new_n1356_), .B(_abc_15497_new_n1354_), .Y(_abc_15497_new_n1357_));
AND2X2 AND2X2_3170 ( .A(w_mem_inst__abc_21203_new_n1624_), .B(w_mem_inst_w_mem_15__19_), .Y(w_mem_inst__abc_21203_new_n2550_));
AND2X2 AND2X2_3171 ( .A(w_mem_inst__abc_21203_new_n1628_), .B(w_mem_inst_w_mem_13__19_), .Y(w_mem_inst__abc_21203_new_n2553_));
AND2X2 AND2X2_3172 ( .A(w_mem_inst__abc_21203_new_n1631_), .B(w_mem_inst_w_mem_0__19_), .Y(w_mem_inst__abc_21203_new_n2554_));
AND2X2 AND2X2_3173 ( .A(w_mem_inst__abc_21203_new_n1633_), .B(w_mem_inst_w_mem_12__19_), .Y(w_mem_inst__abc_21203_new_n2555_));
AND2X2 AND2X2_3174 ( .A(w_mem_inst__abc_21203_new_n1637_), .B(w_mem_inst_w_mem_9__19_), .Y(w_mem_inst__abc_21203_new_n2558_));
AND2X2 AND2X2_3175 ( .A(w_mem_inst__abc_21203_new_n1640_), .B(w_mem_inst_w_mem_10__19_), .Y(w_mem_inst__abc_21203_new_n2559_));
AND2X2 AND2X2_3176 ( .A(w_mem_inst__abc_21203_new_n1643_), .B(w_mem_inst_w_mem_4__19_), .Y(w_mem_inst__abc_21203_new_n2561_));
AND2X2 AND2X2_3177 ( .A(w_mem_inst__abc_21203_new_n1645_), .B(w_mem_inst_w_mem_6__19_), .Y(w_mem_inst__abc_21203_new_n2562_));
AND2X2 AND2X2_3178 ( .A(w_mem_inst__abc_21203_new_n1649_), .B(w_mem_inst_w_mem_1__19_), .Y(w_mem_inst__abc_21203_new_n2565_));
AND2X2 AND2X2_3179 ( .A(w_mem_inst__abc_21203_new_n1651_), .B(w_mem_inst_w_mem_2__19_), .Y(w_mem_inst__abc_21203_new_n2566_));
AND2X2 AND2X2_318 ( .A(_abc_15497_new_n1353_), .B(_abc_15497_new_n1357_), .Y(_abc_15497_new_n1359_));
AND2X2 AND2X2_3180 ( .A(w_mem_inst__abc_21203_new_n1654_), .B(w_mem_inst_w_mem_3__19_), .Y(w_mem_inst__abc_21203_new_n2568_));
AND2X2 AND2X2_3181 ( .A(w_mem_inst__abc_21203_new_n1656_), .B(w_mem_inst_w_mem_14__19_), .Y(w_mem_inst__abc_21203_new_n2569_));
AND2X2 AND2X2_3182 ( .A(w_mem_inst__abc_21203_new_n2574_), .B(w_mem_inst__abc_21203_new_n2542_), .Y(w_19_));
AND2X2 AND2X2_3183 ( .A(w_mem_inst__abc_21203_new_n2577_), .B(w_mem_inst__abc_21203_new_n2579_), .Y(w_mem_inst__abc_21203_new_n2580_));
AND2X2 AND2X2_3184 ( .A(w_mem_inst_w_mem_2__19_), .B(w_mem_inst_w_mem_0__19_), .Y(w_mem_inst__abc_21203_new_n2583_));
AND2X2 AND2X2_3185 ( .A(w_mem_inst__abc_21203_new_n2584_), .B(w_mem_inst__abc_21203_new_n2582_), .Y(w_mem_inst__abc_21203_new_n2585_));
AND2X2 AND2X2_3186 ( .A(w_mem_inst__abc_21203_new_n2586_), .B(w_mem_inst__abc_21203_new_n2588_), .Y(w_mem_inst__abc_21203_new_n2589_));
AND2X2 AND2X2_3187 ( .A(w_mem_inst__abc_21203_new_n1607_), .B(w_mem_inst_w_mem_5__20_), .Y(w_mem_inst__abc_21203_new_n2591_));
AND2X2 AND2X2_3188 ( .A(w_mem_inst__abc_21203_new_n1614_), .B(w_mem_inst_w_mem_8__20_), .Y(w_mem_inst__abc_21203_new_n2593_));
AND2X2 AND2X2_3189 ( .A(w_mem_inst__abc_21203_new_n1617_), .B(w_mem_inst_w_mem_11__20_), .Y(w_mem_inst__abc_21203_new_n2594_));
AND2X2 AND2X2_319 ( .A(_abc_15497_new_n1360_), .B(_abc_15497_new_n1358_), .Y(_abc_15497_new_n1361_));
AND2X2 AND2X2_3190 ( .A(w_mem_inst__abc_21203_new_n1621_), .B(w_mem_inst_w_mem_7__20_), .Y(w_mem_inst__abc_21203_new_n2597_));
AND2X2 AND2X2_3191 ( .A(w_mem_inst__abc_21203_new_n1624_), .B(w_mem_inst_w_mem_15__20_), .Y(w_mem_inst__abc_21203_new_n2598_));
AND2X2 AND2X2_3192 ( .A(w_mem_inst__abc_21203_new_n1628_), .B(w_mem_inst_w_mem_13__20_), .Y(w_mem_inst__abc_21203_new_n2601_));
AND2X2 AND2X2_3193 ( .A(w_mem_inst__abc_21203_new_n1631_), .B(w_mem_inst_w_mem_0__20_), .Y(w_mem_inst__abc_21203_new_n2602_));
AND2X2 AND2X2_3194 ( .A(w_mem_inst__abc_21203_new_n1633_), .B(w_mem_inst_w_mem_12__20_), .Y(w_mem_inst__abc_21203_new_n2603_));
AND2X2 AND2X2_3195 ( .A(w_mem_inst__abc_21203_new_n1637_), .B(w_mem_inst_w_mem_9__20_), .Y(w_mem_inst__abc_21203_new_n2606_));
AND2X2 AND2X2_3196 ( .A(w_mem_inst__abc_21203_new_n1640_), .B(w_mem_inst_w_mem_10__20_), .Y(w_mem_inst__abc_21203_new_n2607_));
AND2X2 AND2X2_3197 ( .A(w_mem_inst__abc_21203_new_n1643_), .B(w_mem_inst_w_mem_4__20_), .Y(w_mem_inst__abc_21203_new_n2609_));
AND2X2 AND2X2_3198 ( .A(w_mem_inst__abc_21203_new_n1645_), .B(w_mem_inst_w_mem_6__20_), .Y(w_mem_inst__abc_21203_new_n2610_));
AND2X2 AND2X2_3199 ( .A(w_mem_inst__abc_21203_new_n1649_), .B(w_mem_inst_w_mem_1__20_), .Y(w_mem_inst__abc_21203_new_n2613_));
AND2X2 AND2X2_32 ( .A(_abc_15497_new_n759_), .B(_abc_15497_new_n760_), .Y(_abc_15497_new_n761_));
AND2X2 AND2X2_320 ( .A(_abc_15497_new_n1361_), .B(digest_update), .Y(_abc_15497_new_n1362_));
AND2X2 AND2X2_3200 ( .A(w_mem_inst__abc_21203_new_n1651_), .B(w_mem_inst_w_mem_2__20_), .Y(w_mem_inst__abc_21203_new_n2614_));
AND2X2 AND2X2_3201 ( .A(w_mem_inst__abc_21203_new_n1654_), .B(w_mem_inst_w_mem_3__20_), .Y(w_mem_inst__abc_21203_new_n2616_));
AND2X2 AND2X2_3202 ( .A(w_mem_inst__abc_21203_new_n1656_), .B(w_mem_inst_w_mem_14__20_), .Y(w_mem_inst__abc_21203_new_n2617_));
AND2X2 AND2X2_3203 ( .A(w_mem_inst__abc_21203_new_n2622_), .B(w_mem_inst__abc_21203_new_n2590_), .Y(w_20_));
AND2X2 AND2X2_3204 ( .A(w_mem_inst__abc_21203_new_n2625_), .B(w_mem_inst__abc_21203_new_n2627_), .Y(w_mem_inst__abc_21203_new_n2628_));
AND2X2 AND2X2_3205 ( .A(w_mem_inst_w_mem_2__20_), .B(w_mem_inst_w_mem_0__20_), .Y(w_mem_inst__abc_21203_new_n2631_));
AND2X2 AND2X2_3206 ( .A(w_mem_inst__abc_21203_new_n2632_), .B(w_mem_inst__abc_21203_new_n2630_), .Y(w_mem_inst__abc_21203_new_n2633_));
AND2X2 AND2X2_3207 ( .A(w_mem_inst__abc_21203_new_n2634_), .B(w_mem_inst__abc_21203_new_n2636_), .Y(w_mem_inst__abc_21203_new_n2637_));
AND2X2 AND2X2_3208 ( .A(w_mem_inst__abc_21203_new_n1607_), .B(w_mem_inst_w_mem_5__21_), .Y(w_mem_inst__abc_21203_new_n2639_));
AND2X2 AND2X2_3209 ( .A(w_mem_inst__abc_21203_new_n1614_), .B(w_mem_inst_w_mem_8__21_), .Y(w_mem_inst__abc_21203_new_n2641_));
AND2X2 AND2X2_321 ( .A(_abc_15497_new_n1363_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n1364_));
AND2X2 AND2X2_3210 ( .A(w_mem_inst__abc_21203_new_n1617_), .B(w_mem_inst_w_mem_11__21_), .Y(w_mem_inst__abc_21203_new_n2642_));
AND2X2 AND2X2_3211 ( .A(w_mem_inst__abc_21203_new_n1621_), .B(w_mem_inst_w_mem_7__21_), .Y(w_mem_inst__abc_21203_new_n2645_));
AND2X2 AND2X2_3212 ( .A(w_mem_inst__abc_21203_new_n1624_), .B(w_mem_inst_w_mem_15__21_), .Y(w_mem_inst__abc_21203_new_n2646_));
AND2X2 AND2X2_3213 ( .A(w_mem_inst__abc_21203_new_n1628_), .B(w_mem_inst_w_mem_13__21_), .Y(w_mem_inst__abc_21203_new_n2649_));
AND2X2 AND2X2_3214 ( .A(w_mem_inst__abc_21203_new_n1631_), .B(w_mem_inst_w_mem_0__21_), .Y(w_mem_inst__abc_21203_new_n2650_));
AND2X2 AND2X2_3215 ( .A(w_mem_inst__abc_21203_new_n1633_), .B(w_mem_inst_w_mem_12__21_), .Y(w_mem_inst__abc_21203_new_n2651_));
AND2X2 AND2X2_3216 ( .A(w_mem_inst__abc_21203_new_n1637_), .B(w_mem_inst_w_mem_9__21_), .Y(w_mem_inst__abc_21203_new_n2654_));
AND2X2 AND2X2_3217 ( .A(w_mem_inst__abc_21203_new_n1640_), .B(w_mem_inst_w_mem_10__21_), .Y(w_mem_inst__abc_21203_new_n2655_));
AND2X2 AND2X2_3218 ( .A(w_mem_inst__abc_21203_new_n1643_), .B(w_mem_inst_w_mem_4__21_), .Y(w_mem_inst__abc_21203_new_n2657_));
AND2X2 AND2X2_3219 ( .A(w_mem_inst__abc_21203_new_n1645_), .B(w_mem_inst_w_mem_6__21_), .Y(w_mem_inst__abc_21203_new_n2658_));
AND2X2 AND2X2_322 ( .A(_abc_15497_new_n1360_), .B(_abc_15497_new_n1356_), .Y(_abc_15497_new_n1366_));
AND2X2 AND2X2_3220 ( .A(w_mem_inst__abc_21203_new_n1649_), .B(w_mem_inst_w_mem_1__21_), .Y(w_mem_inst__abc_21203_new_n2661_));
AND2X2 AND2X2_3221 ( .A(w_mem_inst__abc_21203_new_n1651_), .B(w_mem_inst_w_mem_2__21_), .Y(w_mem_inst__abc_21203_new_n2662_));
AND2X2 AND2X2_3222 ( .A(w_mem_inst__abc_21203_new_n1654_), .B(w_mem_inst_w_mem_3__21_), .Y(w_mem_inst__abc_21203_new_n2664_));
AND2X2 AND2X2_3223 ( .A(w_mem_inst__abc_21203_new_n1656_), .B(w_mem_inst_w_mem_14__21_), .Y(w_mem_inst__abc_21203_new_n2665_));
AND2X2 AND2X2_3224 ( .A(w_mem_inst__abc_21203_new_n2670_), .B(w_mem_inst__abc_21203_new_n2638_), .Y(w_21_));
AND2X2 AND2X2_3225 ( .A(w_mem_inst__abc_21203_new_n2673_), .B(w_mem_inst__abc_21203_new_n2675_), .Y(w_mem_inst__abc_21203_new_n2676_));
AND2X2 AND2X2_3226 ( .A(w_mem_inst_w_mem_2__21_), .B(w_mem_inst_w_mem_0__21_), .Y(w_mem_inst__abc_21203_new_n2679_));
AND2X2 AND2X2_3227 ( .A(w_mem_inst__abc_21203_new_n2680_), .B(w_mem_inst__abc_21203_new_n2678_), .Y(w_mem_inst__abc_21203_new_n2681_));
AND2X2 AND2X2_3228 ( .A(w_mem_inst__abc_21203_new_n2682_), .B(w_mem_inst__abc_21203_new_n2684_), .Y(w_mem_inst__abc_21203_new_n2685_));
AND2X2 AND2X2_3229 ( .A(w_mem_inst__abc_21203_new_n1607_), .B(w_mem_inst_w_mem_5__22_), .Y(w_mem_inst__abc_21203_new_n2687_));
AND2X2 AND2X2_323 ( .A(e_reg_23_), .B(\digest[23] ), .Y(_abc_15497_new_n1368_));
AND2X2 AND2X2_3230 ( .A(w_mem_inst__abc_21203_new_n1614_), .B(w_mem_inst_w_mem_8__22_), .Y(w_mem_inst__abc_21203_new_n2689_));
AND2X2 AND2X2_3231 ( .A(w_mem_inst__abc_21203_new_n1617_), .B(w_mem_inst_w_mem_11__22_), .Y(w_mem_inst__abc_21203_new_n2690_));
AND2X2 AND2X2_3232 ( .A(w_mem_inst__abc_21203_new_n1621_), .B(w_mem_inst_w_mem_7__22_), .Y(w_mem_inst__abc_21203_new_n2693_));
AND2X2 AND2X2_3233 ( .A(w_mem_inst__abc_21203_new_n1624_), .B(w_mem_inst_w_mem_15__22_), .Y(w_mem_inst__abc_21203_new_n2694_));
AND2X2 AND2X2_3234 ( .A(w_mem_inst__abc_21203_new_n1628_), .B(w_mem_inst_w_mem_13__22_), .Y(w_mem_inst__abc_21203_new_n2697_));
AND2X2 AND2X2_3235 ( .A(w_mem_inst__abc_21203_new_n1631_), .B(w_mem_inst_w_mem_0__22_), .Y(w_mem_inst__abc_21203_new_n2698_));
AND2X2 AND2X2_3236 ( .A(w_mem_inst__abc_21203_new_n1633_), .B(w_mem_inst_w_mem_12__22_), .Y(w_mem_inst__abc_21203_new_n2699_));
AND2X2 AND2X2_3237 ( .A(w_mem_inst__abc_21203_new_n1637_), .B(w_mem_inst_w_mem_9__22_), .Y(w_mem_inst__abc_21203_new_n2702_));
AND2X2 AND2X2_3238 ( .A(w_mem_inst__abc_21203_new_n1640_), .B(w_mem_inst_w_mem_10__22_), .Y(w_mem_inst__abc_21203_new_n2703_));
AND2X2 AND2X2_3239 ( .A(w_mem_inst__abc_21203_new_n1643_), .B(w_mem_inst_w_mem_4__22_), .Y(w_mem_inst__abc_21203_new_n2705_));
AND2X2 AND2X2_324 ( .A(_abc_15497_new_n1369_), .B(_abc_15497_new_n1367_), .Y(_abc_15497_new_n1370_));
AND2X2 AND2X2_3240 ( .A(w_mem_inst__abc_21203_new_n1645_), .B(w_mem_inst_w_mem_6__22_), .Y(w_mem_inst__abc_21203_new_n2706_));
AND2X2 AND2X2_3241 ( .A(w_mem_inst__abc_21203_new_n1649_), .B(w_mem_inst_w_mem_1__22_), .Y(w_mem_inst__abc_21203_new_n2709_));
AND2X2 AND2X2_3242 ( .A(w_mem_inst__abc_21203_new_n1651_), .B(w_mem_inst_w_mem_2__22_), .Y(w_mem_inst__abc_21203_new_n2710_));
AND2X2 AND2X2_3243 ( .A(w_mem_inst__abc_21203_new_n1654_), .B(w_mem_inst_w_mem_3__22_), .Y(w_mem_inst__abc_21203_new_n2712_));
AND2X2 AND2X2_3244 ( .A(w_mem_inst__abc_21203_new_n1656_), .B(w_mem_inst_w_mem_14__22_), .Y(w_mem_inst__abc_21203_new_n2713_));
AND2X2 AND2X2_3245 ( .A(w_mem_inst__abc_21203_new_n2718_), .B(w_mem_inst__abc_21203_new_n2686_), .Y(w_22_));
AND2X2 AND2X2_3246 ( .A(w_mem_inst__abc_21203_new_n2721_), .B(w_mem_inst__abc_21203_new_n2723_), .Y(w_mem_inst__abc_21203_new_n2724_));
AND2X2 AND2X2_3247 ( .A(w_mem_inst_w_mem_2__22_), .B(w_mem_inst_w_mem_0__22_), .Y(w_mem_inst__abc_21203_new_n2727_));
AND2X2 AND2X2_3248 ( .A(w_mem_inst__abc_21203_new_n2728_), .B(w_mem_inst__abc_21203_new_n2726_), .Y(w_mem_inst__abc_21203_new_n2729_));
AND2X2 AND2X2_3249 ( .A(w_mem_inst__abc_21203_new_n2730_), .B(w_mem_inst__abc_21203_new_n2732_), .Y(w_mem_inst__abc_21203_new_n2733_));
AND2X2 AND2X2_325 ( .A(_abc_15497_new_n1366_), .B(_abc_15497_new_n1370_), .Y(_abc_15497_new_n1371_));
AND2X2 AND2X2_3250 ( .A(w_mem_inst__abc_21203_new_n1607_), .B(w_mem_inst_w_mem_5__23_), .Y(w_mem_inst__abc_21203_new_n2735_));
AND2X2 AND2X2_3251 ( .A(w_mem_inst__abc_21203_new_n1614_), .B(w_mem_inst_w_mem_8__23_), .Y(w_mem_inst__abc_21203_new_n2737_));
AND2X2 AND2X2_3252 ( .A(w_mem_inst__abc_21203_new_n1617_), .B(w_mem_inst_w_mem_11__23_), .Y(w_mem_inst__abc_21203_new_n2738_));
AND2X2 AND2X2_3253 ( .A(w_mem_inst__abc_21203_new_n1621_), .B(w_mem_inst_w_mem_7__23_), .Y(w_mem_inst__abc_21203_new_n2741_));
AND2X2 AND2X2_3254 ( .A(w_mem_inst__abc_21203_new_n1624_), .B(w_mem_inst_w_mem_15__23_), .Y(w_mem_inst__abc_21203_new_n2742_));
AND2X2 AND2X2_3255 ( .A(w_mem_inst__abc_21203_new_n1628_), .B(w_mem_inst_w_mem_13__23_), .Y(w_mem_inst__abc_21203_new_n2745_));
AND2X2 AND2X2_3256 ( .A(w_mem_inst__abc_21203_new_n1631_), .B(w_mem_inst_w_mem_0__23_), .Y(w_mem_inst__abc_21203_new_n2746_));
AND2X2 AND2X2_3257 ( .A(w_mem_inst__abc_21203_new_n1633_), .B(w_mem_inst_w_mem_12__23_), .Y(w_mem_inst__abc_21203_new_n2747_));
AND2X2 AND2X2_3258 ( .A(w_mem_inst__abc_21203_new_n1637_), .B(w_mem_inst_w_mem_9__23_), .Y(w_mem_inst__abc_21203_new_n2750_));
AND2X2 AND2X2_3259 ( .A(w_mem_inst__abc_21203_new_n1640_), .B(w_mem_inst_w_mem_10__23_), .Y(w_mem_inst__abc_21203_new_n2751_));
AND2X2 AND2X2_326 ( .A(_abc_15497_new_n1372_), .B(_abc_15497_new_n1373_), .Y(_abc_15497_new_n1374_));
AND2X2 AND2X2_3260 ( .A(w_mem_inst__abc_21203_new_n1643_), .B(w_mem_inst_w_mem_4__23_), .Y(w_mem_inst__abc_21203_new_n2753_));
AND2X2 AND2X2_3261 ( .A(w_mem_inst__abc_21203_new_n1645_), .B(w_mem_inst_w_mem_6__23_), .Y(w_mem_inst__abc_21203_new_n2754_));
AND2X2 AND2X2_3262 ( .A(w_mem_inst__abc_21203_new_n1649_), .B(w_mem_inst_w_mem_1__23_), .Y(w_mem_inst__abc_21203_new_n2757_));
AND2X2 AND2X2_3263 ( .A(w_mem_inst__abc_21203_new_n1651_), .B(w_mem_inst_w_mem_2__23_), .Y(w_mem_inst__abc_21203_new_n2758_));
AND2X2 AND2X2_3264 ( .A(w_mem_inst__abc_21203_new_n1654_), .B(w_mem_inst_w_mem_3__23_), .Y(w_mem_inst__abc_21203_new_n2760_));
AND2X2 AND2X2_3265 ( .A(w_mem_inst__abc_21203_new_n1656_), .B(w_mem_inst_w_mem_14__23_), .Y(w_mem_inst__abc_21203_new_n2761_));
AND2X2 AND2X2_3266 ( .A(w_mem_inst__abc_21203_new_n2766_), .B(w_mem_inst__abc_21203_new_n2734_), .Y(w_23_));
AND2X2 AND2X2_3267 ( .A(w_mem_inst__abc_21203_new_n2769_), .B(w_mem_inst__abc_21203_new_n2771_), .Y(w_mem_inst__abc_21203_new_n2772_));
AND2X2 AND2X2_3268 ( .A(w_mem_inst_w_mem_2__23_), .B(w_mem_inst_w_mem_0__23_), .Y(w_mem_inst__abc_21203_new_n2775_));
AND2X2 AND2X2_3269 ( .A(w_mem_inst__abc_21203_new_n2776_), .B(w_mem_inst__abc_21203_new_n2774_), .Y(w_mem_inst__abc_21203_new_n2777_));
AND2X2 AND2X2_327 ( .A(_abc_15497_new_n1375_), .B(digest_update), .Y(_abc_15497_new_n1376_));
AND2X2 AND2X2_3270 ( .A(w_mem_inst__abc_21203_new_n2778_), .B(w_mem_inst__abc_21203_new_n2780_), .Y(w_mem_inst__abc_21203_new_n2781_));
AND2X2 AND2X2_3271 ( .A(w_mem_inst__abc_21203_new_n1607_), .B(w_mem_inst_w_mem_5__24_), .Y(w_mem_inst__abc_21203_new_n2783_));
AND2X2 AND2X2_3272 ( .A(w_mem_inst__abc_21203_new_n1614_), .B(w_mem_inst_w_mem_8__24_), .Y(w_mem_inst__abc_21203_new_n2785_));
AND2X2 AND2X2_3273 ( .A(w_mem_inst__abc_21203_new_n1617_), .B(w_mem_inst_w_mem_11__24_), .Y(w_mem_inst__abc_21203_new_n2786_));
AND2X2 AND2X2_3274 ( .A(w_mem_inst__abc_21203_new_n1621_), .B(w_mem_inst_w_mem_7__24_), .Y(w_mem_inst__abc_21203_new_n2789_));
AND2X2 AND2X2_3275 ( .A(w_mem_inst__abc_21203_new_n1624_), .B(w_mem_inst_w_mem_15__24_), .Y(w_mem_inst__abc_21203_new_n2790_));
AND2X2 AND2X2_3276 ( .A(w_mem_inst__abc_21203_new_n1628_), .B(w_mem_inst_w_mem_13__24_), .Y(w_mem_inst__abc_21203_new_n2793_));
AND2X2 AND2X2_3277 ( .A(w_mem_inst__abc_21203_new_n1631_), .B(w_mem_inst_w_mem_0__24_), .Y(w_mem_inst__abc_21203_new_n2794_));
AND2X2 AND2X2_3278 ( .A(w_mem_inst__abc_21203_new_n1633_), .B(w_mem_inst_w_mem_12__24_), .Y(w_mem_inst__abc_21203_new_n2795_));
AND2X2 AND2X2_3279 ( .A(w_mem_inst__abc_21203_new_n1637_), .B(w_mem_inst_w_mem_9__24_), .Y(w_mem_inst__abc_21203_new_n2798_));
AND2X2 AND2X2_328 ( .A(_abc_15497_new_n1377_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n1378_));
AND2X2 AND2X2_3280 ( .A(w_mem_inst__abc_21203_new_n1640_), .B(w_mem_inst_w_mem_10__24_), .Y(w_mem_inst__abc_21203_new_n2799_));
AND2X2 AND2X2_3281 ( .A(w_mem_inst__abc_21203_new_n1643_), .B(w_mem_inst_w_mem_4__24_), .Y(w_mem_inst__abc_21203_new_n2801_));
AND2X2 AND2X2_3282 ( .A(w_mem_inst__abc_21203_new_n1645_), .B(w_mem_inst_w_mem_6__24_), .Y(w_mem_inst__abc_21203_new_n2802_));
AND2X2 AND2X2_3283 ( .A(w_mem_inst__abc_21203_new_n1649_), .B(w_mem_inst_w_mem_1__24_), .Y(w_mem_inst__abc_21203_new_n2805_));
AND2X2 AND2X2_3284 ( .A(w_mem_inst__abc_21203_new_n1651_), .B(w_mem_inst_w_mem_2__24_), .Y(w_mem_inst__abc_21203_new_n2806_));
AND2X2 AND2X2_3285 ( .A(w_mem_inst__abc_21203_new_n1654_), .B(w_mem_inst_w_mem_3__24_), .Y(w_mem_inst__abc_21203_new_n2808_));
AND2X2 AND2X2_3286 ( .A(w_mem_inst__abc_21203_new_n1656_), .B(w_mem_inst_w_mem_14__24_), .Y(w_mem_inst__abc_21203_new_n2809_));
AND2X2 AND2X2_3287 ( .A(w_mem_inst__abc_21203_new_n2814_), .B(w_mem_inst__abc_21203_new_n2782_), .Y(w_24_));
AND2X2 AND2X2_3288 ( .A(w_mem_inst__abc_21203_new_n2817_), .B(w_mem_inst__abc_21203_new_n2819_), .Y(w_mem_inst__abc_21203_new_n2820_));
AND2X2 AND2X2_3289 ( .A(w_mem_inst_w_mem_2__24_), .B(w_mem_inst_w_mem_0__24_), .Y(w_mem_inst__abc_21203_new_n2823_));
AND2X2 AND2X2_329 ( .A(_abc_15497_new_n1357_), .B(_abc_15497_new_n1370_), .Y(_abc_15497_new_n1380_));
AND2X2 AND2X2_3290 ( .A(w_mem_inst__abc_21203_new_n2824_), .B(w_mem_inst__abc_21203_new_n2822_), .Y(w_mem_inst__abc_21203_new_n2825_));
AND2X2 AND2X2_3291 ( .A(w_mem_inst__abc_21203_new_n2826_), .B(w_mem_inst__abc_21203_new_n2828_), .Y(w_mem_inst__abc_21203_new_n2829_));
AND2X2 AND2X2_3292 ( .A(w_mem_inst__abc_21203_new_n1607_), .B(w_mem_inst_w_mem_5__25_), .Y(w_mem_inst__abc_21203_new_n2831_));
AND2X2 AND2X2_3293 ( .A(w_mem_inst__abc_21203_new_n1614_), .B(w_mem_inst_w_mem_8__25_), .Y(w_mem_inst__abc_21203_new_n2833_));
AND2X2 AND2X2_3294 ( .A(w_mem_inst__abc_21203_new_n1617_), .B(w_mem_inst_w_mem_11__25_), .Y(w_mem_inst__abc_21203_new_n2834_));
AND2X2 AND2X2_3295 ( .A(w_mem_inst__abc_21203_new_n1621_), .B(w_mem_inst_w_mem_7__25_), .Y(w_mem_inst__abc_21203_new_n2837_));
AND2X2 AND2X2_3296 ( .A(w_mem_inst__abc_21203_new_n1624_), .B(w_mem_inst_w_mem_15__25_), .Y(w_mem_inst__abc_21203_new_n2838_));
AND2X2 AND2X2_3297 ( .A(w_mem_inst__abc_21203_new_n1628_), .B(w_mem_inst_w_mem_13__25_), .Y(w_mem_inst__abc_21203_new_n2841_));
AND2X2 AND2X2_3298 ( .A(w_mem_inst__abc_21203_new_n1631_), .B(w_mem_inst_w_mem_0__25_), .Y(w_mem_inst__abc_21203_new_n2842_));
AND2X2 AND2X2_3299 ( .A(w_mem_inst__abc_21203_new_n1633_), .B(w_mem_inst_w_mem_12__25_), .Y(w_mem_inst__abc_21203_new_n2843_));
AND2X2 AND2X2_33 ( .A(c_reg_14_), .B(\digest[78] ), .Y(_abc_15497_new_n762_));
AND2X2 AND2X2_330 ( .A(_abc_15497_new_n1342_), .B(_abc_15497_new_n1380_), .Y(_abc_15497_new_n1381_));
AND2X2 AND2X2_3300 ( .A(w_mem_inst__abc_21203_new_n1637_), .B(w_mem_inst_w_mem_9__25_), .Y(w_mem_inst__abc_21203_new_n2846_));
AND2X2 AND2X2_3301 ( .A(w_mem_inst__abc_21203_new_n1640_), .B(w_mem_inst_w_mem_10__25_), .Y(w_mem_inst__abc_21203_new_n2847_));
AND2X2 AND2X2_3302 ( .A(w_mem_inst__abc_21203_new_n1643_), .B(w_mem_inst_w_mem_4__25_), .Y(w_mem_inst__abc_21203_new_n2849_));
AND2X2 AND2X2_3303 ( .A(w_mem_inst__abc_21203_new_n1645_), .B(w_mem_inst_w_mem_6__25_), .Y(w_mem_inst__abc_21203_new_n2850_));
AND2X2 AND2X2_3304 ( .A(w_mem_inst__abc_21203_new_n1649_), .B(w_mem_inst_w_mem_1__25_), .Y(w_mem_inst__abc_21203_new_n2853_));
AND2X2 AND2X2_3305 ( .A(w_mem_inst__abc_21203_new_n1651_), .B(w_mem_inst_w_mem_2__25_), .Y(w_mem_inst__abc_21203_new_n2854_));
AND2X2 AND2X2_3306 ( .A(w_mem_inst__abc_21203_new_n1654_), .B(w_mem_inst_w_mem_3__25_), .Y(w_mem_inst__abc_21203_new_n2856_));
AND2X2 AND2X2_3307 ( .A(w_mem_inst__abc_21203_new_n1656_), .B(w_mem_inst_w_mem_14__25_), .Y(w_mem_inst__abc_21203_new_n2857_));
AND2X2 AND2X2_3308 ( .A(w_mem_inst__abc_21203_new_n2862_), .B(w_mem_inst__abc_21203_new_n2830_), .Y(w_25_));
AND2X2 AND2X2_3309 ( .A(w_mem_inst__abc_21203_new_n2865_), .B(w_mem_inst__abc_21203_new_n2867_), .Y(w_mem_inst__abc_21203_new_n2868_));
AND2X2 AND2X2_331 ( .A(_abc_15497_new_n1318_), .B(_abc_15497_new_n1381_), .Y(_abc_15497_new_n1382_));
AND2X2 AND2X2_3310 ( .A(w_mem_inst_w_mem_2__25_), .B(w_mem_inst_w_mem_0__25_), .Y(w_mem_inst__abc_21203_new_n2871_));
AND2X2 AND2X2_3311 ( .A(w_mem_inst__abc_21203_new_n2872_), .B(w_mem_inst__abc_21203_new_n2870_), .Y(w_mem_inst__abc_21203_new_n2873_));
AND2X2 AND2X2_3312 ( .A(w_mem_inst__abc_21203_new_n2874_), .B(w_mem_inst__abc_21203_new_n2876_), .Y(w_mem_inst__abc_21203_new_n2877_));
AND2X2 AND2X2_3313 ( .A(w_mem_inst__abc_21203_new_n1607_), .B(w_mem_inst_w_mem_5__26_), .Y(w_mem_inst__abc_21203_new_n2879_));
AND2X2 AND2X2_3314 ( .A(w_mem_inst__abc_21203_new_n1614_), .B(w_mem_inst_w_mem_8__26_), .Y(w_mem_inst__abc_21203_new_n2881_));
AND2X2 AND2X2_3315 ( .A(w_mem_inst__abc_21203_new_n1617_), .B(w_mem_inst_w_mem_11__26_), .Y(w_mem_inst__abc_21203_new_n2882_));
AND2X2 AND2X2_3316 ( .A(w_mem_inst__abc_21203_new_n1621_), .B(w_mem_inst_w_mem_7__26_), .Y(w_mem_inst__abc_21203_new_n2885_));
AND2X2 AND2X2_3317 ( .A(w_mem_inst__abc_21203_new_n1624_), .B(w_mem_inst_w_mem_15__26_), .Y(w_mem_inst__abc_21203_new_n2886_));
AND2X2 AND2X2_3318 ( .A(w_mem_inst__abc_21203_new_n1628_), .B(w_mem_inst_w_mem_13__26_), .Y(w_mem_inst__abc_21203_new_n2889_));
AND2X2 AND2X2_3319 ( .A(w_mem_inst__abc_21203_new_n1631_), .B(w_mem_inst_w_mem_0__26_), .Y(w_mem_inst__abc_21203_new_n2890_));
AND2X2 AND2X2_332 ( .A(_abc_15497_new_n1367_), .B(_abc_15497_new_n1355_), .Y(_abc_15497_new_n1383_));
AND2X2 AND2X2_3320 ( .A(w_mem_inst__abc_21203_new_n1633_), .B(w_mem_inst_w_mem_12__26_), .Y(w_mem_inst__abc_21203_new_n2891_));
AND2X2 AND2X2_3321 ( .A(w_mem_inst__abc_21203_new_n1637_), .B(w_mem_inst_w_mem_9__26_), .Y(w_mem_inst__abc_21203_new_n2894_));
AND2X2 AND2X2_3322 ( .A(w_mem_inst__abc_21203_new_n1640_), .B(w_mem_inst_w_mem_10__26_), .Y(w_mem_inst__abc_21203_new_n2895_));
AND2X2 AND2X2_3323 ( .A(w_mem_inst__abc_21203_new_n1643_), .B(w_mem_inst_w_mem_4__26_), .Y(w_mem_inst__abc_21203_new_n2897_));
AND2X2 AND2X2_3324 ( .A(w_mem_inst__abc_21203_new_n1645_), .B(w_mem_inst_w_mem_6__26_), .Y(w_mem_inst__abc_21203_new_n2898_));
AND2X2 AND2X2_3325 ( .A(w_mem_inst__abc_21203_new_n1649_), .B(w_mem_inst_w_mem_1__26_), .Y(w_mem_inst__abc_21203_new_n2901_));
AND2X2 AND2X2_3326 ( .A(w_mem_inst__abc_21203_new_n1651_), .B(w_mem_inst_w_mem_2__26_), .Y(w_mem_inst__abc_21203_new_n2902_));
AND2X2 AND2X2_3327 ( .A(w_mem_inst__abc_21203_new_n1654_), .B(w_mem_inst_w_mem_3__26_), .Y(w_mem_inst__abc_21203_new_n2904_));
AND2X2 AND2X2_3328 ( .A(w_mem_inst__abc_21203_new_n1656_), .B(w_mem_inst_w_mem_14__26_), .Y(w_mem_inst__abc_21203_new_n2905_));
AND2X2 AND2X2_3329 ( .A(w_mem_inst__abc_21203_new_n2910_), .B(w_mem_inst__abc_21203_new_n2878_), .Y(w_26_));
AND2X2 AND2X2_333 ( .A(_abc_15497_new_n1385_), .B(_abc_15497_new_n1380_), .Y(_abc_15497_new_n1386_));
AND2X2 AND2X2_3330 ( .A(w_mem_inst__abc_21203_new_n2913_), .B(w_mem_inst__abc_21203_new_n2915_), .Y(w_mem_inst__abc_21203_new_n2916_));
AND2X2 AND2X2_3331 ( .A(w_mem_inst_w_mem_2__26_), .B(w_mem_inst_w_mem_0__26_), .Y(w_mem_inst__abc_21203_new_n2919_));
AND2X2 AND2X2_3332 ( .A(w_mem_inst__abc_21203_new_n2920_), .B(w_mem_inst__abc_21203_new_n2918_), .Y(w_mem_inst__abc_21203_new_n2921_));
AND2X2 AND2X2_3333 ( .A(w_mem_inst__abc_21203_new_n2922_), .B(w_mem_inst__abc_21203_new_n2924_), .Y(w_mem_inst__abc_21203_new_n2925_));
AND2X2 AND2X2_3334 ( .A(w_mem_inst__abc_21203_new_n1607_), .B(w_mem_inst_w_mem_5__27_), .Y(w_mem_inst__abc_21203_new_n2927_));
AND2X2 AND2X2_3335 ( .A(w_mem_inst__abc_21203_new_n1614_), .B(w_mem_inst_w_mem_8__27_), .Y(w_mem_inst__abc_21203_new_n2929_));
AND2X2 AND2X2_3336 ( .A(w_mem_inst__abc_21203_new_n1617_), .B(w_mem_inst_w_mem_11__27_), .Y(w_mem_inst__abc_21203_new_n2930_));
AND2X2 AND2X2_3337 ( .A(w_mem_inst__abc_21203_new_n1621_), .B(w_mem_inst_w_mem_7__27_), .Y(w_mem_inst__abc_21203_new_n2933_));
AND2X2 AND2X2_3338 ( .A(w_mem_inst__abc_21203_new_n1624_), .B(w_mem_inst_w_mem_15__27_), .Y(w_mem_inst__abc_21203_new_n2934_));
AND2X2 AND2X2_3339 ( .A(w_mem_inst__abc_21203_new_n1628_), .B(w_mem_inst_w_mem_13__27_), .Y(w_mem_inst__abc_21203_new_n2937_));
AND2X2 AND2X2_334 ( .A(_abc_15497_new_n1320_), .B(_abc_15497_new_n1381_), .Y(_abc_15497_new_n1389_));
AND2X2 AND2X2_3340 ( .A(w_mem_inst__abc_21203_new_n1631_), .B(w_mem_inst_w_mem_0__27_), .Y(w_mem_inst__abc_21203_new_n2938_));
AND2X2 AND2X2_3341 ( .A(w_mem_inst__abc_21203_new_n1633_), .B(w_mem_inst_w_mem_12__27_), .Y(w_mem_inst__abc_21203_new_n2939_));
AND2X2 AND2X2_3342 ( .A(w_mem_inst__abc_21203_new_n1637_), .B(w_mem_inst_w_mem_9__27_), .Y(w_mem_inst__abc_21203_new_n2942_));
AND2X2 AND2X2_3343 ( .A(w_mem_inst__abc_21203_new_n1640_), .B(w_mem_inst_w_mem_10__27_), .Y(w_mem_inst__abc_21203_new_n2943_));
AND2X2 AND2X2_3344 ( .A(w_mem_inst__abc_21203_new_n1643_), .B(w_mem_inst_w_mem_4__27_), .Y(w_mem_inst__abc_21203_new_n2945_));
AND2X2 AND2X2_3345 ( .A(w_mem_inst__abc_21203_new_n1645_), .B(w_mem_inst_w_mem_6__27_), .Y(w_mem_inst__abc_21203_new_n2946_));
AND2X2 AND2X2_3346 ( .A(w_mem_inst__abc_21203_new_n1649_), .B(w_mem_inst_w_mem_1__27_), .Y(w_mem_inst__abc_21203_new_n2949_));
AND2X2 AND2X2_3347 ( .A(w_mem_inst__abc_21203_new_n1651_), .B(w_mem_inst_w_mem_2__27_), .Y(w_mem_inst__abc_21203_new_n2950_));
AND2X2 AND2X2_3348 ( .A(w_mem_inst__abc_21203_new_n1654_), .B(w_mem_inst_w_mem_3__27_), .Y(w_mem_inst__abc_21203_new_n2952_));
AND2X2 AND2X2_3349 ( .A(w_mem_inst__abc_21203_new_n1656_), .B(w_mem_inst_w_mem_14__27_), .Y(w_mem_inst__abc_21203_new_n2953_));
AND2X2 AND2X2_335 ( .A(_abc_15497_new_n1256_), .B(_abc_15497_new_n1389_), .Y(_abc_15497_new_n1390_));
AND2X2 AND2X2_3350 ( .A(w_mem_inst__abc_21203_new_n2958_), .B(w_mem_inst__abc_21203_new_n2926_), .Y(w_27_));
AND2X2 AND2X2_3351 ( .A(w_mem_inst__abc_21203_new_n2961_), .B(w_mem_inst__abc_21203_new_n2963_), .Y(w_mem_inst__abc_21203_new_n2964_));
AND2X2 AND2X2_3352 ( .A(w_mem_inst_w_mem_2__27_), .B(w_mem_inst_w_mem_0__27_), .Y(w_mem_inst__abc_21203_new_n2967_));
AND2X2 AND2X2_3353 ( .A(w_mem_inst__abc_21203_new_n2968_), .B(w_mem_inst__abc_21203_new_n2966_), .Y(w_mem_inst__abc_21203_new_n2969_));
AND2X2 AND2X2_3354 ( .A(w_mem_inst__abc_21203_new_n2970_), .B(w_mem_inst__abc_21203_new_n2972_), .Y(w_mem_inst__abc_21203_new_n2973_));
AND2X2 AND2X2_3355 ( .A(w_mem_inst__abc_21203_new_n1607_), .B(w_mem_inst_w_mem_5__28_), .Y(w_mem_inst__abc_21203_new_n2975_));
AND2X2 AND2X2_3356 ( .A(w_mem_inst__abc_21203_new_n1614_), .B(w_mem_inst_w_mem_8__28_), .Y(w_mem_inst__abc_21203_new_n2977_));
AND2X2 AND2X2_3357 ( .A(w_mem_inst__abc_21203_new_n1617_), .B(w_mem_inst_w_mem_11__28_), .Y(w_mem_inst__abc_21203_new_n2978_));
AND2X2 AND2X2_3358 ( .A(w_mem_inst__abc_21203_new_n1621_), .B(w_mem_inst_w_mem_7__28_), .Y(w_mem_inst__abc_21203_new_n2981_));
AND2X2 AND2X2_3359 ( .A(w_mem_inst__abc_21203_new_n1624_), .B(w_mem_inst_w_mem_15__28_), .Y(w_mem_inst__abc_21203_new_n2982_));
AND2X2 AND2X2_336 ( .A(e_reg_24_), .B(\digest[24] ), .Y(_abc_15497_new_n1393_));
AND2X2 AND2X2_3360 ( .A(w_mem_inst__abc_21203_new_n1628_), .B(w_mem_inst_w_mem_13__28_), .Y(w_mem_inst__abc_21203_new_n2985_));
AND2X2 AND2X2_3361 ( .A(w_mem_inst__abc_21203_new_n1631_), .B(w_mem_inst_w_mem_0__28_), .Y(w_mem_inst__abc_21203_new_n2986_));
AND2X2 AND2X2_3362 ( .A(w_mem_inst__abc_21203_new_n1633_), .B(w_mem_inst_w_mem_12__28_), .Y(w_mem_inst__abc_21203_new_n2987_));
AND2X2 AND2X2_3363 ( .A(w_mem_inst__abc_21203_new_n1637_), .B(w_mem_inst_w_mem_9__28_), .Y(w_mem_inst__abc_21203_new_n2990_));
AND2X2 AND2X2_3364 ( .A(w_mem_inst__abc_21203_new_n1640_), .B(w_mem_inst_w_mem_10__28_), .Y(w_mem_inst__abc_21203_new_n2991_));
AND2X2 AND2X2_3365 ( .A(w_mem_inst__abc_21203_new_n1643_), .B(w_mem_inst_w_mem_4__28_), .Y(w_mem_inst__abc_21203_new_n2993_));
AND2X2 AND2X2_3366 ( .A(w_mem_inst__abc_21203_new_n1645_), .B(w_mem_inst_w_mem_6__28_), .Y(w_mem_inst__abc_21203_new_n2994_));
AND2X2 AND2X2_3367 ( .A(w_mem_inst__abc_21203_new_n1649_), .B(w_mem_inst_w_mem_1__28_), .Y(w_mem_inst__abc_21203_new_n2997_));
AND2X2 AND2X2_3368 ( .A(w_mem_inst__abc_21203_new_n1651_), .B(w_mem_inst_w_mem_2__28_), .Y(w_mem_inst__abc_21203_new_n2998_));
AND2X2 AND2X2_3369 ( .A(w_mem_inst__abc_21203_new_n1654_), .B(w_mem_inst_w_mem_3__28_), .Y(w_mem_inst__abc_21203_new_n3000_));
AND2X2 AND2X2_337 ( .A(_abc_15497_new_n1394_), .B(_abc_15497_new_n1392_), .Y(_abc_15497_new_n1395_));
AND2X2 AND2X2_3370 ( .A(w_mem_inst__abc_21203_new_n1656_), .B(w_mem_inst_w_mem_14__28_), .Y(w_mem_inst__abc_21203_new_n3001_));
AND2X2 AND2X2_3371 ( .A(w_mem_inst__abc_21203_new_n3006_), .B(w_mem_inst__abc_21203_new_n2974_), .Y(w_28_));
AND2X2 AND2X2_3372 ( .A(w_mem_inst__abc_21203_new_n3009_), .B(w_mem_inst__abc_21203_new_n3011_), .Y(w_mem_inst__abc_21203_new_n3012_));
AND2X2 AND2X2_3373 ( .A(w_mem_inst_w_mem_2__28_), .B(w_mem_inst_w_mem_0__28_), .Y(w_mem_inst__abc_21203_new_n3015_));
AND2X2 AND2X2_3374 ( .A(w_mem_inst__abc_21203_new_n3016_), .B(w_mem_inst__abc_21203_new_n3014_), .Y(w_mem_inst__abc_21203_new_n3017_));
AND2X2 AND2X2_3375 ( .A(w_mem_inst__abc_21203_new_n3018_), .B(w_mem_inst__abc_21203_new_n3020_), .Y(w_mem_inst__abc_21203_new_n3021_));
AND2X2 AND2X2_3376 ( .A(w_mem_inst__abc_21203_new_n1607_), .B(w_mem_inst_w_mem_5__29_), .Y(w_mem_inst__abc_21203_new_n3023_));
AND2X2 AND2X2_3377 ( .A(w_mem_inst__abc_21203_new_n1614_), .B(w_mem_inst_w_mem_8__29_), .Y(w_mem_inst__abc_21203_new_n3025_));
AND2X2 AND2X2_3378 ( .A(w_mem_inst__abc_21203_new_n1617_), .B(w_mem_inst_w_mem_11__29_), .Y(w_mem_inst__abc_21203_new_n3026_));
AND2X2 AND2X2_3379 ( .A(w_mem_inst__abc_21203_new_n1621_), .B(w_mem_inst_w_mem_7__29_), .Y(w_mem_inst__abc_21203_new_n3029_));
AND2X2 AND2X2_338 ( .A(_abc_15497_new_n1391_), .B(_abc_15497_new_n1395_), .Y(_abc_15497_new_n1397_));
AND2X2 AND2X2_3380 ( .A(w_mem_inst__abc_21203_new_n1624_), .B(w_mem_inst_w_mem_15__29_), .Y(w_mem_inst__abc_21203_new_n3030_));
AND2X2 AND2X2_3381 ( .A(w_mem_inst__abc_21203_new_n1628_), .B(w_mem_inst_w_mem_13__29_), .Y(w_mem_inst__abc_21203_new_n3033_));
AND2X2 AND2X2_3382 ( .A(w_mem_inst__abc_21203_new_n1631_), .B(w_mem_inst_w_mem_0__29_), .Y(w_mem_inst__abc_21203_new_n3034_));
AND2X2 AND2X2_3383 ( .A(w_mem_inst__abc_21203_new_n1633_), .B(w_mem_inst_w_mem_12__29_), .Y(w_mem_inst__abc_21203_new_n3035_));
AND2X2 AND2X2_3384 ( .A(w_mem_inst__abc_21203_new_n1637_), .B(w_mem_inst_w_mem_9__29_), .Y(w_mem_inst__abc_21203_new_n3038_));
AND2X2 AND2X2_3385 ( .A(w_mem_inst__abc_21203_new_n1640_), .B(w_mem_inst_w_mem_10__29_), .Y(w_mem_inst__abc_21203_new_n3039_));
AND2X2 AND2X2_3386 ( .A(w_mem_inst__abc_21203_new_n1643_), .B(w_mem_inst_w_mem_4__29_), .Y(w_mem_inst__abc_21203_new_n3041_));
AND2X2 AND2X2_3387 ( .A(w_mem_inst__abc_21203_new_n1645_), .B(w_mem_inst_w_mem_6__29_), .Y(w_mem_inst__abc_21203_new_n3042_));
AND2X2 AND2X2_3388 ( .A(w_mem_inst__abc_21203_new_n1649_), .B(w_mem_inst_w_mem_1__29_), .Y(w_mem_inst__abc_21203_new_n3045_));
AND2X2 AND2X2_3389 ( .A(w_mem_inst__abc_21203_new_n1651_), .B(w_mem_inst_w_mem_2__29_), .Y(w_mem_inst__abc_21203_new_n3046_));
AND2X2 AND2X2_339 ( .A(_abc_15497_new_n1398_), .B(_abc_15497_new_n1396_), .Y(_abc_15497_new_n1399_));
AND2X2 AND2X2_3390 ( .A(w_mem_inst__abc_21203_new_n1654_), .B(w_mem_inst_w_mem_3__29_), .Y(w_mem_inst__abc_21203_new_n3048_));
AND2X2 AND2X2_3391 ( .A(w_mem_inst__abc_21203_new_n1656_), .B(w_mem_inst_w_mem_14__29_), .Y(w_mem_inst__abc_21203_new_n3049_));
AND2X2 AND2X2_3392 ( .A(w_mem_inst__abc_21203_new_n3054_), .B(w_mem_inst__abc_21203_new_n3022_), .Y(w_29_));
AND2X2 AND2X2_3393 ( .A(w_mem_inst__abc_21203_new_n3057_), .B(w_mem_inst__abc_21203_new_n3059_), .Y(w_mem_inst__abc_21203_new_n3060_));
AND2X2 AND2X2_3394 ( .A(w_mem_inst_w_mem_2__29_), .B(w_mem_inst_w_mem_0__29_), .Y(w_mem_inst__abc_21203_new_n3063_));
AND2X2 AND2X2_3395 ( .A(w_mem_inst__abc_21203_new_n3064_), .B(w_mem_inst__abc_21203_new_n3062_), .Y(w_mem_inst__abc_21203_new_n3065_));
AND2X2 AND2X2_3396 ( .A(w_mem_inst__abc_21203_new_n3066_), .B(w_mem_inst__abc_21203_new_n3068_), .Y(w_mem_inst__abc_21203_new_n3069_));
AND2X2 AND2X2_3397 ( .A(w_mem_inst__abc_21203_new_n1607_), .B(w_mem_inst_w_mem_5__30_), .Y(w_mem_inst__abc_21203_new_n3071_));
AND2X2 AND2X2_3398 ( .A(w_mem_inst__abc_21203_new_n1614_), .B(w_mem_inst_w_mem_8__30_), .Y(w_mem_inst__abc_21203_new_n3073_));
AND2X2 AND2X2_3399 ( .A(w_mem_inst__abc_21203_new_n1617_), .B(w_mem_inst_w_mem_11__30_), .Y(w_mem_inst__abc_21203_new_n3074_));
AND2X2 AND2X2_34 ( .A(_abc_15497_new_n763_), .B(_abc_15497_new_n764_), .Y(_abc_15497_new_n765_));
AND2X2 AND2X2_340 ( .A(_abc_15497_new_n1399_), .B(digest_update), .Y(_abc_15497_new_n1400_));
AND2X2 AND2X2_3400 ( .A(w_mem_inst__abc_21203_new_n1621_), .B(w_mem_inst_w_mem_7__30_), .Y(w_mem_inst__abc_21203_new_n3077_));
AND2X2 AND2X2_3401 ( .A(w_mem_inst__abc_21203_new_n1624_), .B(w_mem_inst_w_mem_15__30_), .Y(w_mem_inst__abc_21203_new_n3078_));
AND2X2 AND2X2_3402 ( .A(w_mem_inst__abc_21203_new_n1628_), .B(w_mem_inst_w_mem_13__30_), .Y(w_mem_inst__abc_21203_new_n3081_));
AND2X2 AND2X2_3403 ( .A(w_mem_inst__abc_21203_new_n1631_), .B(w_mem_inst_w_mem_0__30_), .Y(w_mem_inst__abc_21203_new_n3082_));
AND2X2 AND2X2_3404 ( .A(w_mem_inst__abc_21203_new_n1633_), .B(w_mem_inst_w_mem_12__30_), .Y(w_mem_inst__abc_21203_new_n3083_));
AND2X2 AND2X2_3405 ( .A(w_mem_inst__abc_21203_new_n1637_), .B(w_mem_inst_w_mem_9__30_), .Y(w_mem_inst__abc_21203_new_n3086_));
AND2X2 AND2X2_3406 ( .A(w_mem_inst__abc_21203_new_n1640_), .B(w_mem_inst_w_mem_10__30_), .Y(w_mem_inst__abc_21203_new_n3087_));
AND2X2 AND2X2_3407 ( .A(w_mem_inst__abc_21203_new_n1643_), .B(w_mem_inst_w_mem_4__30_), .Y(w_mem_inst__abc_21203_new_n3089_));
AND2X2 AND2X2_3408 ( .A(w_mem_inst__abc_21203_new_n1645_), .B(w_mem_inst_w_mem_6__30_), .Y(w_mem_inst__abc_21203_new_n3090_));
AND2X2 AND2X2_3409 ( .A(w_mem_inst__abc_21203_new_n1649_), .B(w_mem_inst_w_mem_1__30_), .Y(w_mem_inst__abc_21203_new_n3093_));
AND2X2 AND2X2_341 ( .A(_abc_15497_new_n1401_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n1402_));
AND2X2 AND2X2_3410 ( .A(w_mem_inst__abc_21203_new_n1651_), .B(w_mem_inst_w_mem_2__30_), .Y(w_mem_inst__abc_21203_new_n3094_));
AND2X2 AND2X2_3411 ( .A(w_mem_inst__abc_21203_new_n1654_), .B(w_mem_inst_w_mem_3__30_), .Y(w_mem_inst__abc_21203_new_n3096_));
AND2X2 AND2X2_3412 ( .A(w_mem_inst__abc_21203_new_n1656_), .B(w_mem_inst_w_mem_14__30_), .Y(w_mem_inst__abc_21203_new_n3097_));
AND2X2 AND2X2_3413 ( .A(w_mem_inst__abc_21203_new_n3102_), .B(w_mem_inst__abc_21203_new_n3070_), .Y(w_30_));
AND2X2 AND2X2_3414 ( .A(w_mem_inst__abc_21203_new_n3105_), .B(w_mem_inst__abc_21203_new_n3107_), .Y(w_mem_inst__abc_21203_new_n3108_));
AND2X2 AND2X2_3415 ( .A(w_mem_inst_w_mem_2__30_), .B(w_mem_inst_w_mem_0__30_), .Y(w_mem_inst__abc_21203_new_n3111_));
AND2X2 AND2X2_3416 ( .A(w_mem_inst__abc_21203_new_n3112_), .B(w_mem_inst__abc_21203_new_n3110_), .Y(w_mem_inst__abc_21203_new_n3113_));
AND2X2 AND2X2_3417 ( .A(w_mem_inst__abc_21203_new_n3114_), .B(w_mem_inst__abc_21203_new_n3116_), .Y(w_mem_inst__abc_21203_new_n3117_));
AND2X2 AND2X2_3418 ( .A(w_mem_inst__abc_21203_new_n1607_), .B(w_mem_inst_w_mem_5__31_), .Y(w_mem_inst__abc_21203_new_n3119_));
AND2X2 AND2X2_3419 ( .A(w_mem_inst__abc_21203_new_n1614_), .B(w_mem_inst_w_mem_8__31_), .Y(w_mem_inst__abc_21203_new_n3121_));
AND2X2 AND2X2_342 ( .A(_abc_15497_new_n1398_), .B(_abc_15497_new_n1394_), .Y(_abc_15497_new_n1404_));
AND2X2 AND2X2_3420 ( .A(w_mem_inst__abc_21203_new_n1617_), .B(w_mem_inst_w_mem_11__31_), .Y(w_mem_inst__abc_21203_new_n3122_));
AND2X2 AND2X2_3421 ( .A(w_mem_inst__abc_21203_new_n1621_), .B(w_mem_inst_w_mem_7__31_), .Y(w_mem_inst__abc_21203_new_n3125_));
AND2X2 AND2X2_3422 ( .A(w_mem_inst__abc_21203_new_n1624_), .B(w_mem_inst_w_mem_15__31_), .Y(w_mem_inst__abc_21203_new_n3126_));
AND2X2 AND2X2_3423 ( .A(w_mem_inst__abc_21203_new_n1628_), .B(w_mem_inst_w_mem_13__31_), .Y(w_mem_inst__abc_21203_new_n3129_));
AND2X2 AND2X2_3424 ( .A(w_mem_inst__abc_21203_new_n1631_), .B(w_mem_inst_w_mem_0__31_), .Y(w_mem_inst__abc_21203_new_n3130_));
AND2X2 AND2X2_3425 ( .A(w_mem_inst__abc_21203_new_n1633_), .B(w_mem_inst_w_mem_12__31_), .Y(w_mem_inst__abc_21203_new_n3131_));
AND2X2 AND2X2_3426 ( .A(w_mem_inst__abc_21203_new_n1637_), .B(w_mem_inst_w_mem_9__31_), .Y(w_mem_inst__abc_21203_new_n3134_));
AND2X2 AND2X2_3427 ( .A(w_mem_inst__abc_21203_new_n1640_), .B(w_mem_inst_w_mem_10__31_), .Y(w_mem_inst__abc_21203_new_n3135_));
AND2X2 AND2X2_3428 ( .A(w_mem_inst__abc_21203_new_n1643_), .B(w_mem_inst_w_mem_4__31_), .Y(w_mem_inst__abc_21203_new_n3137_));
AND2X2 AND2X2_3429 ( .A(w_mem_inst__abc_21203_new_n1645_), .B(w_mem_inst_w_mem_6__31_), .Y(w_mem_inst__abc_21203_new_n3138_));
AND2X2 AND2X2_343 ( .A(e_reg_25_), .B(\digest[25] ), .Y(_abc_15497_new_n1407_));
AND2X2 AND2X2_3430 ( .A(w_mem_inst__abc_21203_new_n1649_), .B(w_mem_inst_w_mem_1__31_), .Y(w_mem_inst__abc_21203_new_n3141_));
AND2X2 AND2X2_3431 ( .A(w_mem_inst__abc_21203_new_n1651_), .B(w_mem_inst_w_mem_2__31_), .Y(w_mem_inst__abc_21203_new_n3142_));
AND2X2 AND2X2_3432 ( .A(w_mem_inst__abc_21203_new_n1654_), .B(w_mem_inst_w_mem_3__31_), .Y(w_mem_inst__abc_21203_new_n3144_));
AND2X2 AND2X2_3433 ( .A(w_mem_inst__abc_21203_new_n1656_), .B(w_mem_inst_w_mem_14__31_), .Y(w_mem_inst__abc_21203_new_n3145_));
AND2X2 AND2X2_3434 ( .A(w_mem_inst__abc_21203_new_n3150_), .B(w_mem_inst__abc_21203_new_n3118_), .Y(w_31_));
AND2X2 AND2X2_3435 ( .A(w_mem_inst__abc_21203_new_n1586_), .B(round_ctr_inc), .Y(w_mem_inst__abc_21203_new_n3153_));
AND2X2 AND2X2_3436 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3152_), .Y(w_mem_inst__abc_21203_new_n3155_));
AND2X2 AND2X2_3437 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_13__0_), .Y(w_mem_inst__abc_21203_new_n3156_));
AND2X2 AND2X2_3438 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_14__0_), .Y(w_mem_inst__abc_21203_new_n3157_));
AND2X2 AND2X2_3439 ( .A(round_ctr_rst), .B(\block[64] ), .Y(w_mem_inst__abc_21203_new_n3158_));
AND2X2 AND2X2_344 ( .A(_abc_15497_new_n1408_), .B(_abc_15497_new_n1406_), .Y(_abc_15497_new_n1409_));
AND2X2 AND2X2_3440 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3158_), .Y(w_mem_inst__abc_21203_new_n3159_));
AND2X2 AND2X2_3441 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_13__1_), .Y(w_mem_inst__abc_21203_new_n3162_));
AND2X2 AND2X2_3442 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_14__1_), .Y(w_mem_inst__abc_21203_new_n3163_));
AND2X2 AND2X2_3443 ( .A(round_ctr_rst), .B(\block[65] ), .Y(w_mem_inst__abc_21203_new_n3164_));
AND2X2 AND2X2_3444 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3164_), .Y(w_mem_inst__abc_21203_new_n3165_));
AND2X2 AND2X2_3445 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_13__2_), .Y(w_mem_inst__abc_21203_new_n3168_));
AND2X2 AND2X2_3446 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_14__2_), .Y(w_mem_inst__abc_21203_new_n3169_));
AND2X2 AND2X2_3447 ( .A(round_ctr_rst), .B(\block[66] ), .Y(w_mem_inst__abc_21203_new_n3170_));
AND2X2 AND2X2_3448 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3170_), .Y(w_mem_inst__abc_21203_new_n3171_));
AND2X2 AND2X2_3449 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_13__3_), .Y(w_mem_inst__abc_21203_new_n3174_));
AND2X2 AND2X2_345 ( .A(_abc_15497_new_n1410_), .B(_abc_15497_new_n1412_), .Y(_abc_15497_new_n1413_));
AND2X2 AND2X2_3450 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_14__3_), .Y(w_mem_inst__abc_21203_new_n3175_));
AND2X2 AND2X2_3451 ( .A(round_ctr_rst), .B(\block[67] ), .Y(w_mem_inst__abc_21203_new_n3176_));
AND2X2 AND2X2_3452 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3176_), .Y(w_mem_inst__abc_21203_new_n3177_));
AND2X2 AND2X2_3453 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_13__4_), .Y(w_mem_inst__abc_21203_new_n3180_));
AND2X2 AND2X2_3454 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_14__4_), .Y(w_mem_inst__abc_21203_new_n3181_));
AND2X2 AND2X2_3455 ( .A(round_ctr_rst), .B(\block[68] ), .Y(w_mem_inst__abc_21203_new_n3182_));
AND2X2 AND2X2_3456 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3182_), .Y(w_mem_inst__abc_21203_new_n3183_));
AND2X2 AND2X2_3457 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_13__5_), .Y(w_mem_inst__abc_21203_new_n3186_));
AND2X2 AND2X2_3458 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_14__5_), .Y(w_mem_inst__abc_21203_new_n3187_));
AND2X2 AND2X2_3459 ( .A(round_ctr_rst), .B(\block[69] ), .Y(w_mem_inst__abc_21203_new_n3188_));
AND2X2 AND2X2_346 ( .A(_abc_15497_new_n1413_), .B(digest_update), .Y(_abc_15497_new_n1414_));
AND2X2 AND2X2_3460 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3188_), .Y(w_mem_inst__abc_21203_new_n3189_));
AND2X2 AND2X2_3461 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_13__6_), .Y(w_mem_inst__abc_21203_new_n3192_));
AND2X2 AND2X2_3462 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_14__6_), .Y(w_mem_inst__abc_21203_new_n3193_));
AND2X2 AND2X2_3463 ( .A(round_ctr_rst), .B(\block[70] ), .Y(w_mem_inst__abc_21203_new_n3194_));
AND2X2 AND2X2_3464 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3194_), .Y(w_mem_inst__abc_21203_new_n3195_));
AND2X2 AND2X2_3465 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_13__7_), .Y(w_mem_inst__abc_21203_new_n3198_));
AND2X2 AND2X2_3466 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_14__7_), .Y(w_mem_inst__abc_21203_new_n3199_));
AND2X2 AND2X2_3467 ( .A(round_ctr_rst), .B(\block[71] ), .Y(w_mem_inst__abc_21203_new_n3200_));
AND2X2 AND2X2_3468 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3200_), .Y(w_mem_inst__abc_21203_new_n3201_));
AND2X2 AND2X2_3469 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_13__8_), .Y(w_mem_inst__abc_21203_new_n3204_));
AND2X2 AND2X2_347 ( .A(_abc_15497_new_n1415_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n1416_));
AND2X2 AND2X2_3470 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_14__8_), .Y(w_mem_inst__abc_21203_new_n3205_));
AND2X2 AND2X2_3471 ( .A(round_ctr_rst), .B(\block[72] ), .Y(w_mem_inst__abc_21203_new_n3206_));
AND2X2 AND2X2_3472 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3206_), .Y(w_mem_inst__abc_21203_new_n3207_));
AND2X2 AND2X2_3473 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_13__9_), .Y(w_mem_inst__abc_21203_new_n3210_));
AND2X2 AND2X2_3474 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_14__9_), .Y(w_mem_inst__abc_21203_new_n3211_));
AND2X2 AND2X2_3475 ( .A(round_ctr_rst), .B(\block[73] ), .Y(w_mem_inst__abc_21203_new_n3212_));
AND2X2 AND2X2_3476 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3212_), .Y(w_mem_inst__abc_21203_new_n3213_));
AND2X2 AND2X2_3477 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_13__10_), .Y(w_mem_inst__abc_21203_new_n3216_));
AND2X2 AND2X2_3478 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_14__10_), .Y(w_mem_inst__abc_21203_new_n3217_));
AND2X2 AND2X2_3479 ( .A(round_ctr_rst), .B(\block[74] ), .Y(w_mem_inst__abc_21203_new_n3218_));
AND2X2 AND2X2_348 ( .A(_abc_15497_new_n701_), .B(\digest[26] ), .Y(_abc_15497_new_n1418_));
AND2X2 AND2X2_3480 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3218_), .Y(w_mem_inst__abc_21203_new_n3219_));
AND2X2 AND2X2_3481 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_13__11_), .Y(w_mem_inst__abc_21203_new_n3222_));
AND2X2 AND2X2_3482 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_14__11_), .Y(w_mem_inst__abc_21203_new_n3223_));
AND2X2 AND2X2_3483 ( .A(round_ctr_rst), .B(\block[75] ), .Y(w_mem_inst__abc_21203_new_n3224_));
AND2X2 AND2X2_3484 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3224_), .Y(w_mem_inst__abc_21203_new_n3225_));
AND2X2 AND2X2_3485 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_13__12_), .Y(w_mem_inst__abc_21203_new_n3228_));
AND2X2 AND2X2_3486 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_14__12_), .Y(w_mem_inst__abc_21203_new_n3229_));
AND2X2 AND2X2_3487 ( .A(round_ctr_rst), .B(\block[76] ), .Y(w_mem_inst__abc_21203_new_n3230_));
AND2X2 AND2X2_3488 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3230_), .Y(w_mem_inst__abc_21203_new_n3231_));
AND2X2 AND2X2_3489 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_13__13_), .Y(w_mem_inst__abc_21203_new_n3234_));
AND2X2 AND2X2_349 ( .A(_abc_15497_new_n1395_), .B(_abc_15497_new_n1409_), .Y(_abc_15497_new_n1419_));
AND2X2 AND2X2_3490 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_14__13_), .Y(w_mem_inst__abc_21203_new_n3235_));
AND2X2 AND2X2_3491 ( .A(round_ctr_rst), .B(\block[77] ), .Y(w_mem_inst__abc_21203_new_n3236_));
AND2X2 AND2X2_3492 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3236_), .Y(w_mem_inst__abc_21203_new_n3237_));
AND2X2 AND2X2_3493 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_13__14_), .Y(w_mem_inst__abc_21203_new_n3240_));
AND2X2 AND2X2_3494 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_14__14_), .Y(w_mem_inst__abc_21203_new_n3241_));
AND2X2 AND2X2_3495 ( .A(round_ctr_rst), .B(\block[78] ), .Y(w_mem_inst__abc_21203_new_n3242_));
AND2X2 AND2X2_3496 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3242_), .Y(w_mem_inst__abc_21203_new_n3243_));
AND2X2 AND2X2_3497 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_13__15_), .Y(w_mem_inst__abc_21203_new_n3246_));
AND2X2 AND2X2_3498 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_14__15_), .Y(w_mem_inst__abc_21203_new_n3247_));
AND2X2 AND2X2_3499 ( .A(round_ctr_rst), .B(\block[79] ), .Y(w_mem_inst__abc_21203_new_n3248_));
AND2X2 AND2X2_35 ( .A(_abc_15497_new_n761_), .B(_abc_15497_new_n765_), .Y(_abc_15497_new_n766_));
AND2X2 AND2X2_350 ( .A(_abc_15497_new_n1391_), .B(_abc_15497_new_n1419_), .Y(_abc_15497_new_n1420_));
AND2X2 AND2X2_3500 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3248_), .Y(w_mem_inst__abc_21203_new_n3249_));
AND2X2 AND2X2_3501 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_13__16_), .Y(w_mem_inst__abc_21203_new_n3252_));
AND2X2 AND2X2_3502 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_14__16_), .Y(w_mem_inst__abc_21203_new_n3253_));
AND2X2 AND2X2_3503 ( .A(round_ctr_rst), .B(\block[80] ), .Y(w_mem_inst__abc_21203_new_n3254_));
AND2X2 AND2X2_3504 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3254_), .Y(w_mem_inst__abc_21203_new_n3255_));
AND2X2 AND2X2_3505 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_13__17_), .Y(w_mem_inst__abc_21203_new_n3258_));
AND2X2 AND2X2_3506 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_14__17_), .Y(w_mem_inst__abc_21203_new_n3259_));
AND2X2 AND2X2_3507 ( .A(round_ctr_rst), .B(\block[81] ), .Y(w_mem_inst__abc_21203_new_n3260_));
AND2X2 AND2X2_3508 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3260_), .Y(w_mem_inst__abc_21203_new_n3261_));
AND2X2 AND2X2_3509 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_13__18_), .Y(w_mem_inst__abc_21203_new_n3264_));
AND2X2 AND2X2_351 ( .A(_abc_15497_new_n1406_), .B(_abc_15497_new_n1393_), .Y(_abc_15497_new_n1421_));
AND2X2 AND2X2_3510 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_14__18_), .Y(w_mem_inst__abc_21203_new_n3265_));
AND2X2 AND2X2_3511 ( .A(round_ctr_rst), .B(\block[82] ), .Y(w_mem_inst__abc_21203_new_n3266_));
AND2X2 AND2X2_3512 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3266_), .Y(w_mem_inst__abc_21203_new_n3267_));
AND2X2 AND2X2_3513 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_13__19_), .Y(w_mem_inst__abc_21203_new_n3270_));
AND2X2 AND2X2_3514 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_14__19_), .Y(w_mem_inst__abc_21203_new_n3271_));
AND2X2 AND2X2_3515 ( .A(round_ctr_rst), .B(\block[83] ), .Y(w_mem_inst__abc_21203_new_n3272_));
AND2X2 AND2X2_3516 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3272_), .Y(w_mem_inst__abc_21203_new_n3273_));
AND2X2 AND2X2_3517 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_13__20_), .Y(w_mem_inst__abc_21203_new_n3276_));
AND2X2 AND2X2_3518 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_14__20_), .Y(w_mem_inst__abc_21203_new_n3277_));
AND2X2 AND2X2_3519 ( .A(round_ctr_rst), .B(\block[84] ), .Y(w_mem_inst__abc_21203_new_n3278_));
AND2X2 AND2X2_352 ( .A(e_reg_26_), .B(\digest[26] ), .Y(_abc_15497_new_n1425_));
AND2X2 AND2X2_3520 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3278_), .Y(w_mem_inst__abc_21203_new_n3279_));
AND2X2 AND2X2_3521 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_13__21_), .Y(w_mem_inst__abc_21203_new_n3282_));
AND2X2 AND2X2_3522 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_14__21_), .Y(w_mem_inst__abc_21203_new_n3283_));
AND2X2 AND2X2_3523 ( .A(round_ctr_rst), .B(\block[85] ), .Y(w_mem_inst__abc_21203_new_n3284_));
AND2X2 AND2X2_3524 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3284_), .Y(w_mem_inst__abc_21203_new_n3285_));
AND2X2 AND2X2_3525 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_13__22_), .Y(w_mem_inst__abc_21203_new_n3288_));
AND2X2 AND2X2_3526 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_14__22_), .Y(w_mem_inst__abc_21203_new_n3289_));
AND2X2 AND2X2_3527 ( .A(round_ctr_rst), .B(\block[86] ), .Y(w_mem_inst__abc_21203_new_n3290_));
AND2X2 AND2X2_3528 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3290_), .Y(w_mem_inst__abc_21203_new_n3291_));
AND2X2 AND2X2_3529 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_13__23_), .Y(w_mem_inst__abc_21203_new_n3294_));
AND2X2 AND2X2_353 ( .A(_abc_15497_new_n1426_), .B(_abc_15497_new_n1424_), .Y(_abc_15497_new_n1427_));
AND2X2 AND2X2_3530 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_14__23_), .Y(w_mem_inst__abc_21203_new_n3295_));
AND2X2 AND2X2_3531 ( .A(round_ctr_rst), .B(\block[87] ), .Y(w_mem_inst__abc_21203_new_n3296_));
AND2X2 AND2X2_3532 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3296_), .Y(w_mem_inst__abc_21203_new_n3297_));
AND2X2 AND2X2_3533 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_13__24_), .Y(w_mem_inst__abc_21203_new_n3300_));
AND2X2 AND2X2_3534 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_14__24_), .Y(w_mem_inst__abc_21203_new_n3301_));
AND2X2 AND2X2_3535 ( .A(round_ctr_rst), .B(\block[88] ), .Y(w_mem_inst__abc_21203_new_n3302_));
AND2X2 AND2X2_3536 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3302_), .Y(w_mem_inst__abc_21203_new_n3303_));
AND2X2 AND2X2_3537 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_13__25_), .Y(w_mem_inst__abc_21203_new_n3306_));
AND2X2 AND2X2_3538 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_14__25_), .Y(w_mem_inst__abc_21203_new_n3307_));
AND2X2 AND2X2_3539 ( .A(round_ctr_rst), .B(\block[89] ), .Y(w_mem_inst__abc_21203_new_n3308_));
AND2X2 AND2X2_354 ( .A(_abc_15497_new_n1423_), .B(_abc_15497_new_n1427_), .Y(_abc_15497_new_n1429_));
AND2X2 AND2X2_3540 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3308_), .Y(w_mem_inst__abc_21203_new_n3309_));
AND2X2 AND2X2_3541 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_13__26_), .Y(w_mem_inst__abc_21203_new_n3312_));
AND2X2 AND2X2_3542 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_14__26_), .Y(w_mem_inst__abc_21203_new_n3313_));
AND2X2 AND2X2_3543 ( .A(round_ctr_rst), .B(\block[90] ), .Y(w_mem_inst__abc_21203_new_n3314_));
AND2X2 AND2X2_3544 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3314_), .Y(w_mem_inst__abc_21203_new_n3315_));
AND2X2 AND2X2_3545 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_13__27_), .Y(w_mem_inst__abc_21203_new_n3318_));
AND2X2 AND2X2_3546 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_14__27_), .Y(w_mem_inst__abc_21203_new_n3319_));
AND2X2 AND2X2_3547 ( .A(round_ctr_rst), .B(\block[91] ), .Y(w_mem_inst__abc_21203_new_n3320_));
AND2X2 AND2X2_3548 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3320_), .Y(w_mem_inst__abc_21203_new_n3321_));
AND2X2 AND2X2_3549 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_13__28_), .Y(w_mem_inst__abc_21203_new_n3324_));
AND2X2 AND2X2_355 ( .A(_abc_15497_new_n1430_), .B(_abc_15497_new_n1428_), .Y(_abc_15497_new_n1431_));
AND2X2 AND2X2_3550 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_14__28_), .Y(w_mem_inst__abc_21203_new_n3325_));
AND2X2 AND2X2_3551 ( .A(round_ctr_rst), .B(\block[92] ), .Y(w_mem_inst__abc_21203_new_n3326_));
AND2X2 AND2X2_3552 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3326_), .Y(w_mem_inst__abc_21203_new_n3327_));
AND2X2 AND2X2_3553 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_13__29_), .Y(w_mem_inst__abc_21203_new_n3330_));
AND2X2 AND2X2_3554 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_14__29_), .Y(w_mem_inst__abc_21203_new_n3331_));
AND2X2 AND2X2_3555 ( .A(round_ctr_rst), .B(\block[93] ), .Y(w_mem_inst__abc_21203_new_n3332_));
AND2X2 AND2X2_3556 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3332_), .Y(w_mem_inst__abc_21203_new_n3333_));
AND2X2 AND2X2_3557 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_13__30_), .Y(w_mem_inst__abc_21203_new_n3336_));
AND2X2 AND2X2_3558 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_14__30_), .Y(w_mem_inst__abc_21203_new_n3337_));
AND2X2 AND2X2_3559 ( .A(round_ctr_rst), .B(\block[94] ), .Y(w_mem_inst__abc_21203_new_n3338_));
AND2X2 AND2X2_356 ( .A(_abc_15497_new_n1431_), .B(digest_update), .Y(_abc_15497_new_n1432_));
AND2X2 AND2X2_3560 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3338_), .Y(w_mem_inst__abc_21203_new_n3339_));
AND2X2 AND2X2_3561 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_13__31_), .Y(w_mem_inst__abc_21203_new_n3342_));
AND2X2 AND2X2_3562 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_14__31_), .Y(w_mem_inst__abc_21203_new_n3343_));
AND2X2 AND2X2_3563 ( .A(round_ctr_rst), .B(\block[95] ), .Y(w_mem_inst__abc_21203_new_n3344_));
AND2X2 AND2X2_3564 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3344_), .Y(w_mem_inst__abc_21203_new_n3345_));
AND2X2 AND2X2_3565 ( .A(w_mem_inst__abc_21203_new_n1601_), .B(w_mem_inst__abc_21203_new_n3153_), .Y(w_mem_inst__abc_21203_new_n3348_));
AND2X2 AND2X2_3566 ( .A(round_ctr_rst), .B(\block[0] ), .Y(w_mem_inst__abc_21203_new_n3349_));
AND2X2 AND2X2_3567 ( .A(w_mem_inst__abc_21203_new_n3152_), .B(w_mem_inst_w_mem_15__0_), .Y(w_mem_inst__abc_21203_new_n3350_));
AND2X2 AND2X2_3568 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3351_), .Y(w_mem_inst__abc_21203_new_n3352_));
AND2X2 AND2X2_3569 ( .A(round_ctr_rst), .B(\block[1] ), .Y(w_mem_inst__abc_21203_new_n3354_));
AND2X2 AND2X2_357 ( .A(_abc_15497_new_n701_), .B(\digest[27] ), .Y(_abc_15497_new_n1434_));
AND2X2 AND2X2_3570 ( .A(w_mem_inst__abc_21203_new_n3152_), .B(w_mem_inst_w_mem_15__1_), .Y(w_mem_inst__abc_21203_new_n3355_));
AND2X2 AND2X2_3571 ( .A(w_mem_inst__abc_21203_new_n3358_), .B(w_mem_inst__abc_21203_new_n3357_), .Y(w_mem_inst__0w_mem_15__31_0__1_));
AND2X2 AND2X2_3572 ( .A(round_ctr_rst), .B(\block[2] ), .Y(w_mem_inst__abc_21203_new_n3360_));
AND2X2 AND2X2_3573 ( .A(w_mem_inst__abc_21203_new_n3152_), .B(w_mem_inst_w_mem_15__2_), .Y(w_mem_inst__abc_21203_new_n3361_));
AND2X2 AND2X2_3574 ( .A(w_mem_inst__abc_21203_new_n3364_), .B(w_mem_inst__abc_21203_new_n3363_), .Y(w_mem_inst__0w_mem_15__31_0__2_));
AND2X2 AND2X2_3575 ( .A(w_mem_inst__abc_21203_new_n1773_), .B(w_mem_inst__abc_21203_new_n3153_), .Y(w_mem_inst__abc_21203_new_n3366_));
AND2X2 AND2X2_3576 ( .A(round_ctr_rst), .B(\block[3] ), .Y(w_mem_inst__abc_21203_new_n3367_));
AND2X2 AND2X2_3577 ( .A(w_mem_inst__abc_21203_new_n3152_), .B(w_mem_inst_w_mem_15__3_), .Y(w_mem_inst__abc_21203_new_n3368_));
AND2X2 AND2X2_3578 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3369_), .Y(w_mem_inst__abc_21203_new_n3370_));
AND2X2 AND2X2_3579 ( .A(round_ctr_rst), .B(\block[4] ), .Y(w_mem_inst__abc_21203_new_n3372_));
AND2X2 AND2X2_358 ( .A(e_reg_27_), .B(\digest[27] ), .Y(_abc_15497_new_n1436_));
AND2X2 AND2X2_3580 ( .A(w_mem_inst__abc_21203_new_n3152_), .B(w_mem_inst_w_mem_15__4_), .Y(w_mem_inst__abc_21203_new_n3373_));
AND2X2 AND2X2_3581 ( .A(w_mem_inst__abc_21203_new_n3376_), .B(w_mem_inst__abc_21203_new_n3375_), .Y(w_mem_inst__0w_mem_15__31_0__4_));
AND2X2 AND2X2_3582 ( .A(w_mem_inst__abc_21203_new_n1869_), .B(w_mem_inst__abc_21203_new_n3153_), .Y(w_mem_inst__abc_21203_new_n3378_));
AND2X2 AND2X2_3583 ( .A(round_ctr_rst), .B(\block[5] ), .Y(w_mem_inst__abc_21203_new_n3379_));
AND2X2 AND2X2_3584 ( .A(w_mem_inst__abc_21203_new_n3152_), .B(w_mem_inst_w_mem_15__5_), .Y(w_mem_inst__abc_21203_new_n3380_));
AND2X2 AND2X2_3585 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3381_), .Y(w_mem_inst__abc_21203_new_n3382_));
AND2X2 AND2X2_3586 ( .A(w_mem_inst__abc_21203_new_n1917_), .B(w_mem_inst__abc_21203_new_n3153_), .Y(w_mem_inst__abc_21203_new_n3384_));
AND2X2 AND2X2_3587 ( .A(round_ctr_rst), .B(\block[6] ), .Y(w_mem_inst__abc_21203_new_n3385_));
AND2X2 AND2X2_3588 ( .A(w_mem_inst__abc_21203_new_n3152_), .B(w_mem_inst_w_mem_15__6_), .Y(w_mem_inst__abc_21203_new_n3386_));
AND2X2 AND2X2_3589 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3387_), .Y(w_mem_inst__abc_21203_new_n3388_));
AND2X2 AND2X2_359 ( .A(_abc_15497_new_n1437_), .B(_abc_15497_new_n1435_), .Y(_abc_15497_new_n1438_));
AND2X2 AND2X2_3590 ( .A(w_mem_inst__abc_21203_new_n1965_), .B(w_mem_inst__abc_21203_new_n3153_), .Y(w_mem_inst__abc_21203_new_n3390_));
AND2X2 AND2X2_3591 ( .A(round_ctr_rst), .B(\block[7] ), .Y(w_mem_inst__abc_21203_new_n3391_));
AND2X2 AND2X2_3592 ( .A(w_mem_inst__abc_21203_new_n3152_), .B(w_mem_inst_w_mem_15__7_), .Y(w_mem_inst__abc_21203_new_n3392_));
AND2X2 AND2X2_3593 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3393_), .Y(w_mem_inst__abc_21203_new_n3394_));
AND2X2 AND2X2_3594 ( .A(round_ctr_rst), .B(\block[8] ), .Y(w_mem_inst__abc_21203_new_n3396_));
AND2X2 AND2X2_3595 ( .A(w_mem_inst__abc_21203_new_n3152_), .B(w_mem_inst_w_mem_15__8_), .Y(w_mem_inst__abc_21203_new_n3397_));
AND2X2 AND2X2_3596 ( .A(w_mem_inst__abc_21203_new_n3400_), .B(w_mem_inst__abc_21203_new_n3399_), .Y(w_mem_inst__0w_mem_15__31_0__8_));
AND2X2 AND2X2_3597 ( .A(round_ctr_rst), .B(\block[9] ), .Y(w_mem_inst__abc_21203_new_n3402_));
AND2X2 AND2X2_3598 ( .A(w_mem_inst__abc_21203_new_n3152_), .B(w_mem_inst_w_mem_15__9_), .Y(w_mem_inst__abc_21203_new_n3403_));
AND2X2 AND2X2_3599 ( .A(w_mem_inst__abc_21203_new_n3406_), .B(w_mem_inst__abc_21203_new_n3405_), .Y(w_mem_inst__0w_mem_15__31_0__9_));
AND2X2 AND2X2_36 ( .A(c_reg_13_), .B(\digest[77] ), .Y(_abc_15497_new_n767_));
AND2X2 AND2X2_360 ( .A(_abc_15497_new_n1444_), .B(_abc_15497_new_n1108_), .Y(_abc_15497_new_n1445_));
AND2X2 AND2X2_3600 ( .A(w_mem_inst__abc_21203_new_n2109_), .B(w_mem_inst__abc_21203_new_n3153_), .Y(w_mem_inst__abc_21203_new_n3408_));
AND2X2 AND2X2_3601 ( .A(round_ctr_rst), .B(\block[10] ), .Y(w_mem_inst__abc_21203_new_n3409_));
AND2X2 AND2X2_3602 ( .A(w_mem_inst__abc_21203_new_n3152_), .B(w_mem_inst_w_mem_15__10_), .Y(w_mem_inst__abc_21203_new_n3410_));
AND2X2 AND2X2_3603 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3411_), .Y(w_mem_inst__abc_21203_new_n3412_));
AND2X2 AND2X2_3604 ( .A(w_mem_inst__abc_21203_new_n2157_), .B(w_mem_inst__abc_21203_new_n3153_), .Y(w_mem_inst__abc_21203_new_n3414_));
AND2X2 AND2X2_3605 ( .A(round_ctr_rst), .B(\block[11] ), .Y(w_mem_inst__abc_21203_new_n3415_));
AND2X2 AND2X2_3606 ( .A(w_mem_inst__abc_21203_new_n3152_), .B(w_mem_inst_w_mem_15__11_), .Y(w_mem_inst__abc_21203_new_n3416_));
AND2X2 AND2X2_3607 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3417_), .Y(w_mem_inst__abc_21203_new_n3418_));
AND2X2 AND2X2_3608 ( .A(round_ctr_rst), .B(\block[12] ), .Y(w_mem_inst__abc_21203_new_n3420_));
AND2X2 AND2X2_3609 ( .A(w_mem_inst__abc_21203_new_n3152_), .B(w_mem_inst_w_mem_15__12_), .Y(w_mem_inst__abc_21203_new_n3421_));
AND2X2 AND2X2_361 ( .A(_abc_15497_new_n1447_), .B(_abc_15497_new_n1442_), .Y(_abc_15497_new_n1448_));
AND2X2 AND2X2_3610 ( .A(w_mem_inst__abc_21203_new_n3424_), .B(w_mem_inst__abc_21203_new_n3423_), .Y(w_mem_inst__0w_mem_15__31_0__12_));
AND2X2 AND2X2_3611 ( .A(w_mem_inst__abc_21203_new_n2253_), .B(w_mem_inst__abc_21203_new_n3153_), .Y(w_mem_inst__abc_21203_new_n3426_));
AND2X2 AND2X2_3612 ( .A(round_ctr_rst), .B(\block[13] ), .Y(w_mem_inst__abc_21203_new_n3427_));
AND2X2 AND2X2_3613 ( .A(w_mem_inst__abc_21203_new_n3152_), .B(w_mem_inst_w_mem_15__13_), .Y(w_mem_inst__abc_21203_new_n3428_));
AND2X2 AND2X2_3614 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3429_), .Y(w_mem_inst__abc_21203_new_n3430_));
AND2X2 AND2X2_3615 ( .A(w_mem_inst__abc_21203_new_n2301_), .B(w_mem_inst__abc_21203_new_n3153_), .Y(w_mem_inst__abc_21203_new_n3432_));
AND2X2 AND2X2_3616 ( .A(round_ctr_rst), .B(\block[14] ), .Y(w_mem_inst__abc_21203_new_n3433_));
AND2X2 AND2X2_3617 ( .A(w_mem_inst__abc_21203_new_n3152_), .B(w_mem_inst_w_mem_15__14_), .Y(w_mem_inst__abc_21203_new_n3434_));
AND2X2 AND2X2_3618 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3435_), .Y(w_mem_inst__abc_21203_new_n3436_));
AND2X2 AND2X2_3619 ( .A(round_ctr_rst), .B(\block[15] ), .Y(w_mem_inst__abc_21203_new_n3438_));
AND2X2 AND2X2_362 ( .A(_abc_15497_new_n1450_), .B(_abc_15497_new_n1441_), .Y(_abc_15497_new_n1451_));
AND2X2 AND2X2_3620 ( .A(w_mem_inst__abc_21203_new_n3152_), .B(w_mem_inst_w_mem_15__15_), .Y(w_mem_inst__abc_21203_new_n3439_));
AND2X2 AND2X2_3621 ( .A(w_mem_inst__abc_21203_new_n3442_), .B(w_mem_inst__abc_21203_new_n3441_), .Y(w_mem_inst__0w_mem_15__31_0__15_));
AND2X2 AND2X2_3622 ( .A(w_mem_inst__abc_21203_new_n2397_), .B(w_mem_inst__abc_21203_new_n3153_), .Y(w_mem_inst__abc_21203_new_n3444_));
AND2X2 AND2X2_3623 ( .A(round_ctr_rst), .B(\block[16] ), .Y(w_mem_inst__abc_21203_new_n3445_));
AND2X2 AND2X2_3624 ( .A(w_mem_inst__abc_21203_new_n3152_), .B(w_mem_inst_w_mem_15__16_), .Y(w_mem_inst__abc_21203_new_n3446_));
AND2X2 AND2X2_3625 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3447_), .Y(w_mem_inst__abc_21203_new_n3448_));
AND2X2 AND2X2_3626 ( .A(w_mem_inst__abc_21203_new_n2445_), .B(w_mem_inst__abc_21203_new_n3153_), .Y(w_mem_inst__abc_21203_new_n3450_));
AND2X2 AND2X2_3627 ( .A(round_ctr_rst), .B(\block[17] ), .Y(w_mem_inst__abc_21203_new_n3451_));
AND2X2 AND2X2_3628 ( .A(w_mem_inst__abc_21203_new_n3152_), .B(w_mem_inst_w_mem_15__17_), .Y(w_mem_inst__abc_21203_new_n3452_));
AND2X2 AND2X2_3629 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3453_), .Y(w_mem_inst__abc_21203_new_n3454_));
AND2X2 AND2X2_363 ( .A(_abc_15497_new_n1453_), .B(_abc_15497_new_n1454_), .Y(_abc_15497_new_n1455_));
AND2X2 AND2X2_3630 ( .A(w_mem_inst__abc_21203_new_n2493_), .B(w_mem_inst__abc_21203_new_n3153_), .Y(w_mem_inst__abc_21203_new_n3456_));
AND2X2 AND2X2_3631 ( .A(round_ctr_rst), .B(\block[18] ), .Y(w_mem_inst__abc_21203_new_n3457_));
AND2X2 AND2X2_3632 ( .A(w_mem_inst__abc_21203_new_n3152_), .B(w_mem_inst_w_mem_15__18_), .Y(w_mem_inst__abc_21203_new_n3458_));
AND2X2 AND2X2_3633 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3459_), .Y(w_mem_inst__abc_21203_new_n3460_));
AND2X2 AND2X2_3634 ( .A(w_mem_inst__abc_21203_new_n2541_), .B(w_mem_inst__abc_21203_new_n3153_), .Y(w_mem_inst__abc_21203_new_n3462_));
AND2X2 AND2X2_3635 ( .A(round_ctr_rst), .B(\block[19] ), .Y(w_mem_inst__abc_21203_new_n3463_));
AND2X2 AND2X2_3636 ( .A(w_mem_inst__abc_21203_new_n3152_), .B(w_mem_inst_w_mem_15__19_), .Y(w_mem_inst__abc_21203_new_n3464_));
AND2X2 AND2X2_3637 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3465_), .Y(w_mem_inst__abc_21203_new_n3466_));
AND2X2 AND2X2_3638 ( .A(w_mem_inst__abc_21203_new_n2589_), .B(w_mem_inst__abc_21203_new_n3153_), .Y(w_mem_inst__abc_21203_new_n3468_));
AND2X2 AND2X2_3639 ( .A(round_ctr_rst), .B(\block[20] ), .Y(w_mem_inst__abc_21203_new_n3469_));
AND2X2 AND2X2_364 ( .A(_abc_15497_new_n1427_), .B(_abc_15497_new_n1438_), .Y(_abc_15497_new_n1456_));
AND2X2 AND2X2_3640 ( .A(w_mem_inst__abc_21203_new_n3152_), .B(w_mem_inst_w_mem_15__20_), .Y(w_mem_inst__abc_21203_new_n3470_));
AND2X2 AND2X2_3641 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3471_), .Y(w_mem_inst__abc_21203_new_n3472_));
AND2X2 AND2X2_3642 ( .A(w_mem_inst__abc_21203_new_n2637_), .B(w_mem_inst__abc_21203_new_n3153_), .Y(w_mem_inst__abc_21203_new_n3474_));
AND2X2 AND2X2_3643 ( .A(round_ctr_rst), .B(\block[21] ), .Y(w_mem_inst__abc_21203_new_n3475_));
AND2X2 AND2X2_3644 ( .A(w_mem_inst__abc_21203_new_n3152_), .B(w_mem_inst_w_mem_15__21_), .Y(w_mem_inst__abc_21203_new_n3476_));
AND2X2 AND2X2_3645 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3477_), .Y(w_mem_inst__abc_21203_new_n3478_));
AND2X2 AND2X2_3646 ( .A(w_mem_inst__abc_21203_new_n2685_), .B(w_mem_inst__abc_21203_new_n3153_), .Y(w_mem_inst__abc_21203_new_n3480_));
AND2X2 AND2X2_3647 ( .A(round_ctr_rst), .B(\block[22] ), .Y(w_mem_inst__abc_21203_new_n3481_));
AND2X2 AND2X2_3648 ( .A(w_mem_inst__abc_21203_new_n3152_), .B(w_mem_inst_w_mem_15__22_), .Y(w_mem_inst__abc_21203_new_n3482_));
AND2X2 AND2X2_3649 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3483_), .Y(w_mem_inst__abc_21203_new_n3484_));
AND2X2 AND2X2_365 ( .A(_abc_15497_new_n1438_), .B(_abc_15497_new_n1425_), .Y(_abc_15497_new_n1459_));
AND2X2 AND2X2_3650 ( .A(w_mem_inst__abc_21203_new_n2733_), .B(w_mem_inst__abc_21203_new_n3153_), .Y(w_mem_inst__abc_21203_new_n3486_));
AND2X2 AND2X2_3651 ( .A(round_ctr_rst), .B(\block[23] ), .Y(w_mem_inst__abc_21203_new_n3487_));
AND2X2 AND2X2_3652 ( .A(w_mem_inst__abc_21203_new_n3152_), .B(w_mem_inst_w_mem_15__23_), .Y(w_mem_inst__abc_21203_new_n3488_));
AND2X2 AND2X2_3653 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3489_), .Y(w_mem_inst__abc_21203_new_n3490_));
AND2X2 AND2X2_3654 ( .A(round_ctr_rst), .B(\block[24] ), .Y(w_mem_inst__abc_21203_new_n3492_));
AND2X2 AND2X2_3655 ( .A(w_mem_inst__abc_21203_new_n3152_), .B(w_mem_inst_w_mem_15__24_), .Y(w_mem_inst__abc_21203_new_n3493_));
AND2X2 AND2X2_3656 ( .A(w_mem_inst__abc_21203_new_n3496_), .B(w_mem_inst__abc_21203_new_n3495_), .Y(w_mem_inst__0w_mem_15__31_0__24_));
AND2X2 AND2X2_3657 ( .A(round_ctr_rst), .B(\block[25] ), .Y(w_mem_inst__abc_21203_new_n3498_));
AND2X2 AND2X2_3658 ( .A(w_mem_inst__abc_21203_new_n3152_), .B(w_mem_inst_w_mem_15__25_), .Y(w_mem_inst__abc_21203_new_n3499_));
AND2X2 AND2X2_3659 ( .A(w_mem_inst__abc_21203_new_n3502_), .B(w_mem_inst__abc_21203_new_n3501_), .Y(w_mem_inst__0w_mem_15__31_0__25_));
AND2X2 AND2X2_366 ( .A(_abc_15497_new_n1460_), .B(digest_update), .Y(_abc_15497_new_n1461_));
AND2X2 AND2X2_3660 ( .A(w_mem_inst__abc_21203_new_n2877_), .B(w_mem_inst__abc_21203_new_n3153_), .Y(w_mem_inst__abc_21203_new_n3504_));
AND2X2 AND2X2_3661 ( .A(round_ctr_rst), .B(\block[26] ), .Y(w_mem_inst__abc_21203_new_n3505_));
AND2X2 AND2X2_3662 ( .A(w_mem_inst__abc_21203_new_n3152_), .B(w_mem_inst_w_mem_15__26_), .Y(w_mem_inst__abc_21203_new_n3506_));
AND2X2 AND2X2_3663 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3507_), .Y(w_mem_inst__abc_21203_new_n3508_));
AND2X2 AND2X2_3664 ( .A(w_mem_inst__abc_21203_new_n2925_), .B(w_mem_inst__abc_21203_new_n3153_), .Y(w_mem_inst__abc_21203_new_n3510_));
AND2X2 AND2X2_3665 ( .A(round_ctr_rst), .B(\block[27] ), .Y(w_mem_inst__abc_21203_new_n3511_));
AND2X2 AND2X2_3666 ( .A(w_mem_inst__abc_21203_new_n3152_), .B(w_mem_inst_w_mem_15__27_), .Y(w_mem_inst__abc_21203_new_n3512_));
AND2X2 AND2X2_3667 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3513_), .Y(w_mem_inst__abc_21203_new_n3514_));
AND2X2 AND2X2_3668 ( .A(round_ctr_rst), .B(\block[28] ), .Y(w_mem_inst__abc_21203_new_n3516_));
AND2X2 AND2X2_3669 ( .A(w_mem_inst__abc_21203_new_n3152_), .B(w_mem_inst_w_mem_15__28_), .Y(w_mem_inst__abc_21203_new_n3517_));
AND2X2 AND2X2_367 ( .A(_abc_15497_new_n1458_), .B(_abc_15497_new_n1461_), .Y(_abc_15497_new_n1462_));
AND2X2 AND2X2_3670 ( .A(w_mem_inst__abc_21203_new_n3520_), .B(w_mem_inst__abc_21203_new_n3519_), .Y(w_mem_inst__0w_mem_15__31_0__28_));
AND2X2 AND2X2_3671 ( .A(w_mem_inst__abc_21203_new_n3021_), .B(w_mem_inst__abc_21203_new_n3153_), .Y(w_mem_inst__abc_21203_new_n3522_));
AND2X2 AND2X2_3672 ( .A(round_ctr_rst), .B(\block[29] ), .Y(w_mem_inst__abc_21203_new_n3523_));
AND2X2 AND2X2_3673 ( .A(w_mem_inst__abc_21203_new_n3152_), .B(w_mem_inst_w_mem_15__29_), .Y(w_mem_inst__abc_21203_new_n3524_));
AND2X2 AND2X2_3674 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3525_), .Y(w_mem_inst__abc_21203_new_n3526_));
AND2X2 AND2X2_3675 ( .A(w_mem_inst__abc_21203_new_n3069_), .B(w_mem_inst__abc_21203_new_n3153_), .Y(w_mem_inst__abc_21203_new_n3528_));
AND2X2 AND2X2_3676 ( .A(round_ctr_rst), .B(\block[30] ), .Y(w_mem_inst__abc_21203_new_n3529_));
AND2X2 AND2X2_3677 ( .A(w_mem_inst__abc_21203_new_n3152_), .B(w_mem_inst_w_mem_15__30_), .Y(w_mem_inst__abc_21203_new_n3530_));
AND2X2 AND2X2_3678 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3531_), .Y(w_mem_inst__abc_21203_new_n3532_));
AND2X2 AND2X2_3679 ( .A(round_ctr_rst), .B(\block[31] ), .Y(w_mem_inst__abc_21203_new_n3534_));
AND2X2 AND2X2_368 ( .A(_abc_15497_new_n1462_), .B(_abc_15497_new_n1440_), .Y(_abc_15497_new_n1463_));
AND2X2 AND2X2_3680 ( .A(w_mem_inst__abc_21203_new_n3152_), .B(w_mem_inst_w_mem_15__31_), .Y(w_mem_inst__abc_21203_new_n3535_));
AND2X2 AND2X2_3681 ( .A(w_mem_inst__abc_21203_new_n3538_), .B(w_mem_inst__abc_21203_new_n3537_), .Y(w_mem_inst__0w_mem_15__31_0__31_));
AND2X2 AND2X2_3682 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_14__0_), .Y(w_mem_inst__abc_21203_new_n3540_));
AND2X2 AND2X2_3683 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_15__0_), .Y(w_mem_inst__abc_21203_new_n3541_));
AND2X2 AND2X2_3684 ( .A(round_ctr_rst), .B(\block[32] ), .Y(w_mem_inst__abc_21203_new_n3542_));
AND2X2 AND2X2_3685 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3542_), .Y(w_mem_inst__abc_21203_new_n3543_));
AND2X2 AND2X2_3686 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_14__1_), .Y(w_mem_inst__abc_21203_new_n3546_));
AND2X2 AND2X2_3687 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_15__1_), .Y(w_mem_inst__abc_21203_new_n3547_));
AND2X2 AND2X2_3688 ( .A(round_ctr_rst), .B(\block[33] ), .Y(w_mem_inst__abc_21203_new_n3548_));
AND2X2 AND2X2_3689 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3548_), .Y(w_mem_inst__abc_21203_new_n3549_));
AND2X2 AND2X2_369 ( .A(_abc_15497_new_n701_), .B(\digest[28] ), .Y(_abc_15497_new_n1465_));
AND2X2 AND2X2_3690 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_14__2_), .Y(w_mem_inst__abc_21203_new_n3552_));
AND2X2 AND2X2_3691 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_15__2_), .Y(w_mem_inst__abc_21203_new_n3553_));
AND2X2 AND2X2_3692 ( .A(round_ctr_rst), .B(\block[34] ), .Y(w_mem_inst__abc_21203_new_n3554_));
AND2X2 AND2X2_3693 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3554_), .Y(w_mem_inst__abc_21203_new_n3555_));
AND2X2 AND2X2_3694 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_14__3_), .Y(w_mem_inst__abc_21203_new_n3558_));
AND2X2 AND2X2_3695 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_15__3_), .Y(w_mem_inst__abc_21203_new_n3559_));
AND2X2 AND2X2_3696 ( .A(round_ctr_rst), .B(\block[35] ), .Y(w_mem_inst__abc_21203_new_n3560_));
AND2X2 AND2X2_3697 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3560_), .Y(w_mem_inst__abc_21203_new_n3561_));
AND2X2 AND2X2_3698 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_14__4_), .Y(w_mem_inst__abc_21203_new_n3564_));
AND2X2 AND2X2_3699 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_15__4_), .Y(w_mem_inst__abc_21203_new_n3565_));
AND2X2 AND2X2_37 ( .A(c_reg_12_), .B(\digest[76] ), .Y(_abc_15497_new_n769_));
AND2X2 AND2X2_370 ( .A(_abc_15497_new_n1423_), .B(_abc_15497_new_n1456_), .Y(_abc_15497_new_n1466_));
AND2X2 AND2X2_3700 ( .A(round_ctr_rst), .B(\block[36] ), .Y(w_mem_inst__abc_21203_new_n3566_));
AND2X2 AND2X2_3701 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3566_), .Y(w_mem_inst__abc_21203_new_n3567_));
AND2X2 AND2X2_3702 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_14__5_), .Y(w_mem_inst__abc_21203_new_n3570_));
AND2X2 AND2X2_3703 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_15__5_), .Y(w_mem_inst__abc_21203_new_n3571_));
AND2X2 AND2X2_3704 ( .A(round_ctr_rst), .B(\block[37] ), .Y(w_mem_inst__abc_21203_new_n3572_));
AND2X2 AND2X2_3705 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3572_), .Y(w_mem_inst__abc_21203_new_n3573_));
AND2X2 AND2X2_3706 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_14__6_), .Y(w_mem_inst__abc_21203_new_n3576_));
AND2X2 AND2X2_3707 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_15__6_), .Y(w_mem_inst__abc_21203_new_n3577_));
AND2X2 AND2X2_3708 ( .A(round_ctr_rst), .B(\block[38] ), .Y(w_mem_inst__abc_21203_new_n3578_));
AND2X2 AND2X2_3709 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3578_), .Y(w_mem_inst__abc_21203_new_n3579_));
AND2X2 AND2X2_371 ( .A(_abc_15497_new_n1460_), .B(_abc_15497_new_n1437_), .Y(_abc_15497_new_n1467_));
AND2X2 AND2X2_3710 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_14__7_), .Y(w_mem_inst__abc_21203_new_n3582_));
AND2X2 AND2X2_3711 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_15__7_), .Y(w_mem_inst__abc_21203_new_n3583_));
AND2X2 AND2X2_3712 ( .A(round_ctr_rst), .B(\block[39] ), .Y(w_mem_inst__abc_21203_new_n3584_));
AND2X2 AND2X2_3713 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3584_), .Y(w_mem_inst__abc_21203_new_n3585_));
AND2X2 AND2X2_3714 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_14__8_), .Y(w_mem_inst__abc_21203_new_n3588_));
AND2X2 AND2X2_3715 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_15__8_), .Y(w_mem_inst__abc_21203_new_n3589_));
AND2X2 AND2X2_3716 ( .A(round_ctr_rst), .B(\block[40] ), .Y(w_mem_inst__abc_21203_new_n3590_));
AND2X2 AND2X2_3717 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3590_), .Y(w_mem_inst__abc_21203_new_n3591_));
AND2X2 AND2X2_3718 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_14__9_), .Y(w_mem_inst__abc_21203_new_n3594_));
AND2X2 AND2X2_3719 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_15__9_), .Y(w_mem_inst__abc_21203_new_n3595_));
AND2X2 AND2X2_372 ( .A(e_reg_28_), .B(\digest[28] ), .Y(_abc_15497_new_n1471_));
AND2X2 AND2X2_3720 ( .A(round_ctr_rst), .B(\block[41] ), .Y(w_mem_inst__abc_21203_new_n3596_));
AND2X2 AND2X2_3721 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3596_), .Y(w_mem_inst__abc_21203_new_n3597_));
AND2X2 AND2X2_3722 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_14__10_), .Y(w_mem_inst__abc_21203_new_n3600_));
AND2X2 AND2X2_3723 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_15__10_), .Y(w_mem_inst__abc_21203_new_n3601_));
AND2X2 AND2X2_3724 ( .A(round_ctr_rst), .B(\block[42] ), .Y(w_mem_inst__abc_21203_new_n3602_));
AND2X2 AND2X2_3725 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3602_), .Y(w_mem_inst__abc_21203_new_n3603_));
AND2X2 AND2X2_3726 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_14__11_), .Y(w_mem_inst__abc_21203_new_n3606_));
AND2X2 AND2X2_3727 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_15__11_), .Y(w_mem_inst__abc_21203_new_n3607_));
AND2X2 AND2X2_3728 ( .A(round_ctr_rst), .B(\block[43] ), .Y(w_mem_inst__abc_21203_new_n3608_));
AND2X2 AND2X2_3729 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3608_), .Y(w_mem_inst__abc_21203_new_n3609_));
AND2X2 AND2X2_373 ( .A(_abc_15497_new_n1472_), .B(_abc_15497_new_n1470_), .Y(_abc_15497_new_n1473_));
AND2X2 AND2X2_3730 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_14__12_), .Y(w_mem_inst__abc_21203_new_n3612_));
AND2X2 AND2X2_3731 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_15__12_), .Y(w_mem_inst__abc_21203_new_n3613_));
AND2X2 AND2X2_3732 ( .A(round_ctr_rst), .B(\block[44] ), .Y(w_mem_inst__abc_21203_new_n3614_));
AND2X2 AND2X2_3733 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3614_), .Y(w_mem_inst__abc_21203_new_n3615_));
AND2X2 AND2X2_3734 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_14__13_), .Y(w_mem_inst__abc_21203_new_n3618_));
AND2X2 AND2X2_3735 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_15__13_), .Y(w_mem_inst__abc_21203_new_n3619_));
AND2X2 AND2X2_3736 ( .A(round_ctr_rst), .B(\block[45] ), .Y(w_mem_inst__abc_21203_new_n3620_));
AND2X2 AND2X2_3737 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3620_), .Y(w_mem_inst__abc_21203_new_n3621_));
AND2X2 AND2X2_3738 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_14__14_), .Y(w_mem_inst__abc_21203_new_n3624_));
AND2X2 AND2X2_3739 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_15__14_), .Y(w_mem_inst__abc_21203_new_n3625_));
AND2X2 AND2X2_374 ( .A(_abc_15497_new_n1458_), .B(_abc_15497_new_n1467_), .Y(_abc_15497_new_n1475_));
AND2X2 AND2X2_3740 ( .A(round_ctr_rst), .B(\block[46] ), .Y(w_mem_inst__abc_21203_new_n3626_));
AND2X2 AND2X2_3741 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3626_), .Y(w_mem_inst__abc_21203_new_n3627_));
AND2X2 AND2X2_3742 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_14__15_), .Y(w_mem_inst__abc_21203_new_n3630_));
AND2X2 AND2X2_3743 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_15__15_), .Y(w_mem_inst__abc_21203_new_n3631_));
AND2X2 AND2X2_3744 ( .A(round_ctr_rst), .B(\block[47] ), .Y(w_mem_inst__abc_21203_new_n3632_));
AND2X2 AND2X2_3745 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3632_), .Y(w_mem_inst__abc_21203_new_n3633_));
AND2X2 AND2X2_3746 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_14__16_), .Y(w_mem_inst__abc_21203_new_n3636_));
AND2X2 AND2X2_3747 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_15__16_), .Y(w_mem_inst__abc_21203_new_n3637_));
AND2X2 AND2X2_3748 ( .A(round_ctr_rst), .B(\block[48] ), .Y(w_mem_inst__abc_21203_new_n3638_));
AND2X2 AND2X2_3749 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3638_), .Y(w_mem_inst__abc_21203_new_n3639_));
AND2X2 AND2X2_375 ( .A(_abc_15497_new_n1477_), .B(_abc_15497_new_n1474_), .Y(_abc_15497_new_n1478_));
AND2X2 AND2X2_3750 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_14__17_), .Y(w_mem_inst__abc_21203_new_n3642_));
AND2X2 AND2X2_3751 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_15__17_), .Y(w_mem_inst__abc_21203_new_n3643_));
AND2X2 AND2X2_3752 ( .A(round_ctr_rst), .B(\block[49] ), .Y(w_mem_inst__abc_21203_new_n3644_));
AND2X2 AND2X2_3753 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3644_), .Y(w_mem_inst__abc_21203_new_n3645_));
AND2X2 AND2X2_3754 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_14__18_), .Y(w_mem_inst__abc_21203_new_n3648_));
AND2X2 AND2X2_3755 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_15__18_), .Y(w_mem_inst__abc_21203_new_n3649_));
AND2X2 AND2X2_3756 ( .A(round_ctr_rst), .B(\block[50] ), .Y(w_mem_inst__abc_21203_new_n3650_));
AND2X2 AND2X2_3757 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3650_), .Y(w_mem_inst__abc_21203_new_n3651_));
AND2X2 AND2X2_3758 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_14__19_), .Y(w_mem_inst__abc_21203_new_n3654_));
AND2X2 AND2X2_3759 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_15__19_), .Y(w_mem_inst__abc_21203_new_n3655_));
AND2X2 AND2X2_376 ( .A(_abc_15497_new_n1478_), .B(digest_update), .Y(_abc_15497_new_n1479_));
AND2X2 AND2X2_3760 ( .A(round_ctr_rst), .B(\block[51] ), .Y(w_mem_inst__abc_21203_new_n3656_));
AND2X2 AND2X2_3761 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3656_), .Y(w_mem_inst__abc_21203_new_n3657_));
AND2X2 AND2X2_3762 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_14__20_), .Y(w_mem_inst__abc_21203_new_n3660_));
AND2X2 AND2X2_3763 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_15__20_), .Y(w_mem_inst__abc_21203_new_n3661_));
AND2X2 AND2X2_3764 ( .A(round_ctr_rst), .B(\block[52] ), .Y(w_mem_inst__abc_21203_new_n3662_));
AND2X2 AND2X2_3765 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3662_), .Y(w_mem_inst__abc_21203_new_n3663_));
AND2X2 AND2X2_3766 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_14__21_), .Y(w_mem_inst__abc_21203_new_n3666_));
AND2X2 AND2X2_3767 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_15__21_), .Y(w_mem_inst__abc_21203_new_n3667_));
AND2X2 AND2X2_3768 ( .A(round_ctr_rst), .B(\block[53] ), .Y(w_mem_inst__abc_21203_new_n3668_));
AND2X2 AND2X2_3769 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3668_), .Y(w_mem_inst__abc_21203_new_n3669_));
AND2X2 AND2X2_377 ( .A(_abc_15497_new_n700_), .B(\digest[29] ), .Y(_abc_15497_new_n1481_));
AND2X2 AND2X2_3770 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_14__22_), .Y(w_mem_inst__abc_21203_new_n3672_));
AND2X2 AND2X2_3771 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_15__22_), .Y(w_mem_inst__abc_21203_new_n3673_));
AND2X2 AND2X2_3772 ( .A(round_ctr_rst), .B(\block[54] ), .Y(w_mem_inst__abc_21203_new_n3674_));
AND2X2 AND2X2_3773 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3674_), .Y(w_mem_inst__abc_21203_new_n3675_));
AND2X2 AND2X2_3774 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_14__23_), .Y(w_mem_inst__abc_21203_new_n3678_));
AND2X2 AND2X2_3775 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_15__23_), .Y(w_mem_inst__abc_21203_new_n3679_));
AND2X2 AND2X2_3776 ( .A(round_ctr_rst), .B(\block[55] ), .Y(w_mem_inst__abc_21203_new_n3680_));
AND2X2 AND2X2_3777 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3680_), .Y(w_mem_inst__abc_21203_new_n3681_));
AND2X2 AND2X2_3778 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_14__24_), .Y(w_mem_inst__abc_21203_new_n3684_));
AND2X2 AND2X2_3779 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_15__24_), .Y(w_mem_inst__abc_21203_new_n3685_));
AND2X2 AND2X2_378 ( .A(_abc_15497_new_n1477_), .B(_abc_15497_new_n1472_), .Y(_abc_15497_new_n1483_));
AND2X2 AND2X2_3780 ( .A(round_ctr_rst), .B(\block[56] ), .Y(w_mem_inst__abc_21203_new_n3686_));
AND2X2 AND2X2_3781 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3686_), .Y(w_mem_inst__abc_21203_new_n3687_));
AND2X2 AND2X2_3782 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_14__25_), .Y(w_mem_inst__abc_21203_new_n3690_));
AND2X2 AND2X2_3783 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_15__25_), .Y(w_mem_inst__abc_21203_new_n3691_));
AND2X2 AND2X2_3784 ( .A(round_ctr_rst), .B(\block[57] ), .Y(w_mem_inst__abc_21203_new_n3692_));
AND2X2 AND2X2_3785 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3692_), .Y(w_mem_inst__abc_21203_new_n3693_));
AND2X2 AND2X2_3786 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_14__26_), .Y(w_mem_inst__abc_21203_new_n3696_));
AND2X2 AND2X2_3787 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_15__26_), .Y(w_mem_inst__abc_21203_new_n3697_));
AND2X2 AND2X2_3788 ( .A(round_ctr_rst), .B(\block[58] ), .Y(w_mem_inst__abc_21203_new_n3698_));
AND2X2 AND2X2_3789 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3698_), .Y(w_mem_inst__abc_21203_new_n3699_));
AND2X2 AND2X2_379 ( .A(e_reg_29_), .B(\digest[29] ), .Y(_abc_15497_new_n1485_));
AND2X2 AND2X2_3790 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_14__27_), .Y(w_mem_inst__abc_21203_new_n3702_));
AND2X2 AND2X2_3791 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_15__27_), .Y(w_mem_inst__abc_21203_new_n3703_));
AND2X2 AND2X2_3792 ( .A(round_ctr_rst), .B(\block[59] ), .Y(w_mem_inst__abc_21203_new_n3704_));
AND2X2 AND2X2_3793 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3704_), .Y(w_mem_inst__abc_21203_new_n3705_));
AND2X2 AND2X2_3794 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_14__28_), .Y(w_mem_inst__abc_21203_new_n3708_));
AND2X2 AND2X2_3795 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_15__28_), .Y(w_mem_inst__abc_21203_new_n3709_));
AND2X2 AND2X2_3796 ( .A(round_ctr_rst), .B(\block[60] ), .Y(w_mem_inst__abc_21203_new_n3710_));
AND2X2 AND2X2_3797 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3710_), .Y(w_mem_inst__abc_21203_new_n3711_));
AND2X2 AND2X2_3798 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_14__29_), .Y(w_mem_inst__abc_21203_new_n3714_));
AND2X2 AND2X2_3799 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_15__29_), .Y(w_mem_inst__abc_21203_new_n3715_));
AND2X2 AND2X2_38 ( .A(_abc_15497_new_n768_), .B(_abc_15497_new_n771_), .Y(_abc_15497_new_n772_));
AND2X2 AND2X2_380 ( .A(_abc_15497_new_n1486_), .B(_abc_15497_new_n1484_), .Y(_abc_15497_new_n1487_));
AND2X2 AND2X2_3800 ( .A(round_ctr_rst), .B(\block[61] ), .Y(w_mem_inst__abc_21203_new_n3716_));
AND2X2 AND2X2_3801 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3716_), .Y(w_mem_inst__abc_21203_new_n3717_));
AND2X2 AND2X2_3802 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_14__30_), .Y(w_mem_inst__abc_21203_new_n3720_));
AND2X2 AND2X2_3803 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_15__30_), .Y(w_mem_inst__abc_21203_new_n3721_));
AND2X2 AND2X2_3804 ( .A(round_ctr_rst), .B(\block[62] ), .Y(w_mem_inst__abc_21203_new_n3722_));
AND2X2 AND2X2_3805 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3722_), .Y(w_mem_inst__abc_21203_new_n3723_));
AND2X2 AND2X2_3806 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_14__31_), .Y(w_mem_inst__abc_21203_new_n3726_));
AND2X2 AND2X2_3807 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_15__31_), .Y(w_mem_inst__abc_21203_new_n3727_));
AND2X2 AND2X2_3808 ( .A(round_ctr_rst), .B(\block[63] ), .Y(w_mem_inst__abc_21203_new_n3728_));
AND2X2 AND2X2_3809 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3728_), .Y(w_mem_inst__abc_21203_new_n3729_));
AND2X2 AND2X2_381 ( .A(_abc_15497_new_n1483_), .B(_abc_15497_new_n1487_), .Y(_abc_15497_new_n1488_));
AND2X2 AND2X2_3810 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_10__0_), .Y(w_mem_inst__abc_21203_new_n3732_));
AND2X2 AND2X2_3811 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_11__0_), .Y(w_mem_inst__abc_21203_new_n3733_));
AND2X2 AND2X2_3812 ( .A(round_ctr_rst), .B(\block[160] ), .Y(w_mem_inst__abc_21203_new_n3734_));
AND2X2 AND2X2_3813 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3734_), .Y(w_mem_inst__abc_21203_new_n3735_));
AND2X2 AND2X2_3814 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_10__1_), .Y(w_mem_inst__abc_21203_new_n3738_));
AND2X2 AND2X2_3815 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_11__1_), .Y(w_mem_inst__abc_21203_new_n3739_));
AND2X2 AND2X2_3816 ( .A(round_ctr_rst), .B(\block[161] ), .Y(w_mem_inst__abc_21203_new_n3740_));
AND2X2 AND2X2_3817 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3740_), .Y(w_mem_inst__abc_21203_new_n3741_));
AND2X2 AND2X2_3818 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_10__2_), .Y(w_mem_inst__abc_21203_new_n3744_));
AND2X2 AND2X2_3819 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_11__2_), .Y(w_mem_inst__abc_21203_new_n3745_));
AND2X2 AND2X2_382 ( .A(_abc_15497_new_n1469_), .B(_abc_15497_new_n1473_), .Y(_abc_15497_new_n1489_));
AND2X2 AND2X2_3820 ( .A(round_ctr_rst), .B(\block[162] ), .Y(w_mem_inst__abc_21203_new_n3746_));
AND2X2 AND2X2_3821 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3746_), .Y(w_mem_inst__abc_21203_new_n3747_));
AND2X2 AND2X2_3822 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_10__3_), .Y(w_mem_inst__abc_21203_new_n3750_));
AND2X2 AND2X2_3823 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_11__3_), .Y(w_mem_inst__abc_21203_new_n3751_));
AND2X2 AND2X2_3824 ( .A(round_ctr_rst), .B(\block[163] ), .Y(w_mem_inst__abc_21203_new_n3752_));
AND2X2 AND2X2_3825 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3752_), .Y(w_mem_inst__abc_21203_new_n3753_));
AND2X2 AND2X2_3826 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_10__4_), .Y(w_mem_inst__abc_21203_new_n3756_));
AND2X2 AND2X2_3827 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_11__4_), .Y(w_mem_inst__abc_21203_new_n3757_));
AND2X2 AND2X2_3828 ( .A(round_ctr_rst), .B(\block[164] ), .Y(w_mem_inst__abc_21203_new_n3758_));
AND2X2 AND2X2_3829 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3758_), .Y(w_mem_inst__abc_21203_new_n3759_));
AND2X2 AND2X2_383 ( .A(_abc_15497_new_n1490_), .B(_abc_15497_new_n1491_), .Y(_abc_15497_new_n1492_));
AND2X2 AND2X2_3830 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_10__5_), .Y(w_mem_inst__abc_21203_new_n3762_));
AND2X2 AND2X2_3831 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_11__5_), .Y(w_mem_inst__abc_21203_new_n3763_));
AND2X2 AND2X2_3832 ( .A(round_ctr_rst), .B(\block[165] ), .Y(w_mem_inst__abc_21203_new_n3764_));
AND2X2 AND2X2_3833 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3764_), .Y(w_mem_inst__abc_21203_new_n3765_));
AND2X2 AND2X2_3834 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_10__6_), .Y(w_mem_inst__abc_21203_new_n3768_));
AND2X2 AND2X2_3835 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_11__6_), .Y(w_mem_inst__abc_21203_new_n3769_));
AND2X2 AND2X2_3836 ( .A(round_ctr_rst), .B(\block[166] ), .Y(w_mem_inst__abc_21203_new_n3770_));
AND2X2 AND2X2_3837 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3770_), .Y(w_mem_inst__abc_21203_new_n3771_));
AND2X2 AND2X2_3838 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_10__7_), .Y(w_mem_inst__abc_21203_new_n3774_));
AND2X2 AND2X2_3839 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_11__7_), .Y(w_mem_inst__abc_21203_new_n3775_));
AND2X2 AND2X2_384 ( .A(_abc_15497_new_n1494_), .B(_abc_15497_new_n1482_), .Y(_0H4_reg_31_0__29_));
AND2X2 AND2X2_3840 ( .A(round_ctr_rst), .B(\block[167] ), .Y(w_mem_inst__abc_21203_new_n3776_));
AND2X2 AND2X2_3841 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3776_), .Y(w_mem_inst__abc_21203_new_n3777_));
AND2X2 AND2X2_3842 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_10__8_), .Y(w_mem_inst__abc_21203_new_n3780_));
AND2X2 AND2X2_3843 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_11__8_), .Y(w_mem_inst__abc_21203_new_n3781_));
AND2X2 AND2X2_3844 ( .A(round_ctr_rst), .B(\block[168] ), .Y(w_mem_inst__abc_21203_new_n3782_));
AND2X2 AND2X2_3845 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3782_), .Y(w_mem_inst__abc_21203_new_n3783_));
AND2X2 AND2X2_3846 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_10__9_), .Y(w_mem_inst__abc_21203_new_n3786_));
AND2X2 AND2X2_3847 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_11__9_), .Y(w_mem_inst__abc_21203_new_n3787_));
AND2X2 AND2X2_3848 ( .A(round_ctr_rst), .B(\block[169] ), .Y(w_mem_inst__abc_21203_new_n3788_));
AND2X2 AND2X2_3849 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3788_), .Y(w_mem_inst__abc_21203_new_n3789_));
AND2X2 AND2X2_385 ( .A(e_reg_30_), .B(\digest[30] ), .Y(_abc_15497_new_n1497_));
AND2X2 AND2X2_3850 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_10__10_), .Y(w_mem_inst__abc_21203_new_n3792_));
AND2X2 AND2X2_3851 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_11__10_), .Y(w_mem_inst__abc_21203_new_n3793_));
AND2X2 AND2X2_3852 ( .A(round_ctr_rst), .B(\block[170] ), .Y(w_mem_inst__abc_21203_new_n3794_));
AND2X2 AND2X2_3853 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3794_), .Y(w_mem_inst__abc_21203_new_n3795_));
AND2X2 AND2X2_3854 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_10__11_), .Y(w_mem_inst__abc_21203_new_n3798_));
AND2X2 AND2X2_3855 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_11__11_), .Y(w_mem_inst__abc_21203_new_n3799_));
AND2X2 AND2X2_3856 ( .A(round_ctr_rst), .B(\block[171] ), .Y(w_mem_inst__abc_21203_new_n3800_));
AND2X2 AND2X2_3857 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3800_), .Y(w_mem_inst__abc_21203_new_n3801_));
AND2X2 AND2X2_3858 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_10__12_), .Y(w_mem_inst__abc_21203_new_n3804_));
AND2X2 AND2X2_3859 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_11__12_), .Y(w_mem_inst__abc_21203_new_n3805_));
AND2X2 AND2X2_386 ( .A(_abc_15497_new_n1498_), .B(_abc_15497_new_n1496_), .Y(_abc_15497_new_n1499_));
AND2X2 AND2X2_3860 ( .A(round_ctr_rst), .B(\block[172] ), .Y(w_mem_inst__abc_21203_new_n3806_));
AND2X2 AND2X2_3861 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3806_), .Y(w_mem_inst__abc_21203_new_n3807_));
AND2X2 AND2X2_3862 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_10__13_), .Y(w_mem_inst__abc_21203_new_n3810_));
AND2X2 AND2X2_3863 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_11__13_), .Y(w_mem_inst__abc_21203_new_n3811_));
AND2X2 AND2X2_3864 ( .A(round_ctr_rst), .B(\block[173] ), .Y(w_mem_inst__abc_21203_new_n3812_));
AND2X2 AND2X2_3865 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3812_), .Y(w_mem_inst__abc_21203_new_n3813_));
AND2X2 AND2X2_3866 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_10__14_), .Y(w_mem_inst__abc_21203_new_n3816_));
AND2X2 AND2X2_3867 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_11__14_), .Y(w_mem_inst__abc_21203_new_n3817_));
AND2X2 AND2X2_3868 ( .A(round_ctr_rst), .B(\block[174] ), .Y(w_mem_inst__abc_21203_new_n3818_));
AND2X2 AND2X2_3869 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3818_), .Y(w_mem_inst__abc_21203_new_n3819_));
AND2X2 AND2X2_387 ( .A(_abc_15497_new_n1490_), .B(_abc_15497_new_n1484_), .Y(_abc_15497_new_n1500_));
AND2X2 AND2X2_3870 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_10__15_), .Y(w_mem_inst__abc_21203_new_n3822_));
AND2X2 AND2X2_3871 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_11__15_), .Y(w_mem_inst__abc_21203_new_n3823_));
AND2X2 AND2X2_3872 ( .A(round_ctr_rst), .B(\block[175] ), .Y(w_mem_inst__abc_21203_new_n3824_));
AND2X2 AND2X2_3873 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3824_), .Y(w_mem_inst__abc_21203_new_n3825_));
AND2X2 AND2X2_3874 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_10__16_), .Y(w_mem_inst__abc_21203_new_n3828_));
AND2X2 AND2X2_3875 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_11__16_), .Y(w_mem_inst__abc_21203_new_n3829_));
AND2X2 AND2X2_3876 ( .A(round_ctr_rst), .B(\block[176] ), .Y(w_mem_inst__abc_21203_new_n3830_));
AND2X2 AND2X2_3877 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3830_), .Y(w_mem_inst__abc_21203_new_n3831_));
AND2X2 AND2X2_3878 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_10__17_), .Y(w_mem_inst__abc_21203_new_n3834_));
AND2X2 AND2X2_3879 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_11__17_), .Y(w_mem_inst__abc_21203_new_n3835_));
AND2X2 AND2X2_388 ( .A(_abc_15497_new_n1483_), .B(_abc_15497_new_n1486_), .Y(_abc_15497_new_n1505_));
AND2X2 AND2X2_3880 ( .A(round_ctr_rst), .B(\block[177] ), .Y(w_mem_inst__abc_21203_new_n3836_));
AND2X2 AND2X2_3881 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3836_), .Y(w_mem_inst__abc_21203_new_n3837_));
AND2X2 AND2X2_3882 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_10__18_), .Y(w_mem_inst__abc_21203_new_n3840_));
AND2X2 AND2X2_3883 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_11__18_), .Y(w_mem_inst__abc_21203_new_n3841_));
AND2X2 AND2X2_3884 ( .A(round_ctr_rst), .B(\block[178] ), .Y(w_mem_inst__abc_21203_new_n3842_));
AND2X2 AND2X2_3885 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3842_), .Y(w_mem_inst__abc_21203_new_n3843_));
AND2X2 AND2X2_3886 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_10__19_), .Y(w_mem_inst__abc_21203_new_n3846_));
AND2X2 AND2X2_3887 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_11__19_), .Y(w_mem_inst__abc_21203_new_n3847_));
AND2X2 AND2X2_3888 ( .A(round_ctr_rst), .B(\block[179] ), .Y(w_mem_inst__abc_21203_new_n3848_));
AND2X2 AND2X2_3889 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3848_), .Y(w_mem_inst__abc_21203_new_n3849_));
AND2X2 AND2X2_389 ( .A(_abc_15497_new_n1507_), .B(_abc_15497_new_n1502_), .Y(_abc_15497_new_n1508_));
AND2X2 AND2X2_3890 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_10__20_), .Y(w_mem_inst__abc_21203_new_n3852_));
AND2X2 AND2X2_3891 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_11__20_), .Y(w_mem_inst__abc_21203_new_n3853_));
AND2X2 AND2X2_3892 ( .A(round_ctr_rst), .B(\block[180] ), .Y(w_mem_inst__abc_21203_new_n3854_));
AND2X2 AND2X2_3893 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3854_), .Y(w_mem_inst__abc_21203_new_n3855_));
AND2X2 AND2X2_3894 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_10__21_), .Y(w_mem_inst__abc_21203_new_n3858_));
AND2X2 AND2X2_3895 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_11__21_), .Y(w_mem_inst__abc_21203_new_n3859_));
AND2X2 AND2X2_3896 ( .A(round_ctr_rst), .B(\block[181] ), .Y(w_mem_inst__abc_21203_new_n3860_));
AND2X2 AND2X2_3897 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3860_), .Y(w_mem_inst__abc_21203_new_n3861_));
AND2X2 AND2X2_3898 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_10__22_), .Y(w_mem_inst__abc_21203_new_n3864_));
AND2X2 AND2X2_3899 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_11__22_), .Y(w_mem_inst__abc_21203_new_n3865_));
AND2X2 AND2X2_39 ( .A(_abc_15497_new_n774_), .B(_abc_15497_new_n768_), .Y(_abc_15497_new_n775_));
AND2X2 AND2X2_390 ( .A(_abc_15497_new_n1508_), .B(digest_update), .Y(_abc_15497_new_n1509_));
AND2X2 AND2X2_3900 ( .A(round_ctr_rst), .B(\block[182] ), .Y(w_mem_inst__abc_21203_new_n3866_));
AND2X2 AND2X2_3901 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3866_), .Y(w_mem_inst__abc_21203_new_n3867_));
AND2X2 AND2X2_3902 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_10__23_), .Y(w_mem_inst__abc_21203_new_n3870_));
AND2X2 AND2X2_3903 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_11__23_), .Y(w_mem_inst__abc_21203_new_n3871_));
AND2X2 AND2X2_3904 ( .A(round_ctr_rst), .B(\block[183] ), .Y(w_mem_inst__abc_21203_new_n3872_));
AND2X2 AND2X2_3905 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3872_), .Y(w_mem_inst__abc_21203_new_n3873_));
AND2X2 AND2X2_3906 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_10__24_), .Y(w_mem_inst__abc_21203_new_n3876_));
AND2X2 AND2X2_3907 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_11__24_), .Y(w_mem_inst__abc_21203_new_n3877_));
AND2X2 AND2X2_3908 ( .A(round_ctr_rst), .B(\block[184] ), .Y(w_mem_inst__abc_21203_new_n3878_));
AND2X2 AND2X2_3909 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3878_), .Y(w_mem_inst__abc_21203_new_n3879_));
AND2X2 AND2X2_391 ( .A(_abc_15497_new_n1510_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n1511_));
AND2X2 AND2X2_3910 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_10__25_), .Y(w_mem_inst__abc_21203_new_n3882_));
AND2X2 AND2X2_3911 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_11__25_), .Y(w_mem_inst__abc_21203_new_n3883_));
AND2X2 AND2X2_3912 ( .A(round_ctr_rst), .B(\block[185] ), .Y(w_mem_inst__abc_21203_new_n3884_));
AND2X2 AND2X2_3913 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3884_), .Y(w_mem_inst__abc_21203_new_n3885_));
AND2X2 AND2X2_3914 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_10__26_), .Y(w_mem_inst__abc_21203_new_n3888_));
AND2X2 AND2X2_3915 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_11__26_), .Y(w_mem_inst__abc_21203_new_n3889_));
AND2X2 AND2X2_3916 ( .A(round_ctr_rst), .B(\block[186] ), .Y(w_mem_inst__abc_21203_new_n3890_));
AND2X2 AND2X2_3917 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3890_), .Y(w_mem_inst__abc_21203_new_n3891_));
AND2X2 AND2X2_3918 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_10__27_), .Y(w_mem_inst__abc_21203_new_n3894_));
AND2X2 AND2X2_3919 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_11__27_), .Y(w_mem_inst__abc_21203_new_n3895_));
AND2X2 AND2X2_392 ( .A(_abc_15497_new_n1501_), .B(_abc_15497_new_n1499_), .Y(_abc_15497_new_n1513_));
AND2X2 AND2X2_3920 ( .A(round_ctr_rst), .B(\block[187] ), .Y(w_mem_inst__abc_21203_new_n3896_));
AND2X2 AND2X2_3921 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3896_), .Y(w_mem_inst__abc_21203_new_n3897_));
AND2X2 AND2X2_3922 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_10__28_), .Y(w_mem_inst__abc_21203_new_n3900_));
AND2X2 AND2X2_3923 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_11__28_), .Y(w_mem_inst__abc_21203_new_n3901_));
AND2X2 AND2X2_3924 ( .A(round_ctr_rst), .B(\block[188] ), .Y(w_mem_inst__abc_21203_new_n3902_));
AND2X2 AND2X2_3925 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3902_), .Y(w_mem_inst__abc_21203_new_n3903_));
AND2X2 AND2X2_3926 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_10__29_), .Y(w_mem_inst__abc_21203_new_n3906_));
AND2X2 AND2X2_3927 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_11__29_), .Y(w_mem_inst__abc_21203_new_n3907_));
AND2X2 AND2X2_3928 ( .A(round_ctr_rst), .B(\block[189] ), .Y(w_mem_inst__abc_21203_new_n3908_));
AND2X2 AND2X2_3929 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3908_), .Y(w_mem_inst__abc_21203_new_n3909_));
AND2X2 AND2X2_393 ( .A(_abc_15497_new_n1516_), .B(_abc_15497_new_n1518_), .Y(_abc_15497_new_n1519_));
AND2X2 AND2X2_3930 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_10__30_), .Y(w_mem_inst__abc_21203_new_n3912_));
AND2X2 AND2X2_3931 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_11__30_), .Y(w_mem_inst__abc_21203_new_n3913_));
AND2X2 AND2X2_3932 ( .A(round_ctr_rst), .B(\block[190] ), .Y(w_mem_inst__abc_21203_new_n3914_));
AND2X2 AND2X2_3933 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3914_), .Y(w_mem_inst__abc_21203_new_n3915_));
AND2X2 AND2X2_3934 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_10__31_), .Y(w_mem_inst__abc_21203_new_n3918_));
AND2X2 AND2X2_3935 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_11__31_), .Y(w_mem_inst__abc_21203_new_n3919_));
AND2X2 AND2X2_3936 ( .A(round_ctr_rst), .B(\block[191] ), .Y(w_mem_inst__abc_21203_new_n3920_));
AND2X2 AND2X2_3937 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3920_), .Y(w_mem_inst__abc_21203_new_n3921_));
AND2X2 AND2X2_3938 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_12__0_), .Y(w_mem_inst__abc_21203_new_n3924_));
AND2X2 AND2X2_3939 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_13__0_), .Y(w_mem_inst__abc_21203_new_n3925_));
AND2X2 AND2X2_394 ( .A(_abc_15497_new_n1507_), .B(_abc_15497_new_n1498_), .Y(_abc_15497_new_n1522_));
AND2X2 AND2X2_3940 ( .A(round_ctr_rst), .B(\block[96] ), .Y(w_mem_inst__abc_21203_new_n3926_));
AND2X2 AND2X2_3941 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3926_), .Y(w_mem_inst__abc_21203_new_n3927_));
AND2X2 AND2X2_3942 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_12__1_), .Y(w_mem_inst__abc_21203_new_n3930_));
AND2X2 AND2X2_3943 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_13__1_), .Y(w_mem_inst__abc_21203_new_n3931_));
AND2X2 AND2X2_3944 ( .A(round_ctr_rst), .B(\block[97] ), .Y(w_mem_inst__abc_21203_new_n3932_));
AND2X2 AND2X2_3945 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3932_), .Y(w_mem_inst__abc_21203_new_n3933_));
AND2X2 AND2X2_3946 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_12__2_), .Y(w_mem_inst__abc_21203_new_n3936_));
AND2X2 AND2X2_3947 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_13__2_), .Y(w_mem_inst__abc_21203_new_n3937_));
AND2X2 AND2X2_3948 ( .A(round_ctr_rst), .B(\block[98] ), .Y(w_mem_inst__abc_21203_new_n3938_));
AND2X2 AND2X2_3949 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3938_), .Y(w_mem_inst__abc_21203_new_n3939_));
AND2X2 AND2X2_395 ( .A(_abc_15497_new_n1523_), .B(_abc_15497_new_n1521_), .Y(_abc_15497_new_n1524_));
AND2X2 AND2X2_3950 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_12__3_), .Y(w_mem_inst__abc_21203_new_n3942_));
AND2X2 AND2X2_3951 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_13__3_), .Y(w_mem_inst__abc_21203_new_n3943_));
AND2X2 AND2X2_3952 ( .A(round_ctr_rst), .B(\block[99] ), .Y(w_mem_inst__abc_21203_new_n3944_));
AND2X2 AND2X2_3953 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3944_), .Y(w_mem_inst__abc_21203_new_n3945_));
AND2X2 AND2X2_3954 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_12__4_), .Y(w_mem_inst__abc_21203_new_n3948_));
AND2X2 AND2X2_3955 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_13__4_), .Y(w_mem_inst__abc_21203_new_n3949_));
AND2X2 AND2X2_3956 ( .A(round_ctr_rst), .B(\block[100] ), .Y(w_mem_inst__abc_21203_new_n3950_));
AND2X2 AND2X2_3957 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3950_), .Y(w_mem_inst__abc_21203_new_n3951_));
AND2X2 AND2X2_3958 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_12__5_), .Y(w_mem_inst__abc_21203_new_n3954_));
AND2X2 AND2X2_3959 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_13__5_), .Y(w_mem_inst__abc_21203_new_n3955_));
AND2X2 AND2X2_396 ( .A(_abc_15497_new_n1524_), .B(digest_update), .Y(_abc_15497_new_n1525_));
AND2X2 AND2X2_3960 ( .A(round_ctr_rst), .B(\block[101] ), .Y(w_mem_inst__abc_21203_new_n3956_));
AND2X2 AND2X2_3961 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3956_), .Y(w_mem_inst__abc_21203_new_n3957_));
AND2X2 AND2X2_3962 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_12__6_), .Y(w_mem_inst__abc_21203_new_n3960_));
AND2X2 AND2X2_3963 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_13__6_), .Y(w_mem_inst__abc_21203_new_n3961_));
AND2X2 AND2X2_3964 ( .A(round_ctr_rst), .B(\block[102] ), .Y(w_mem_inst__abc_21203_new_n3962_));
AND2X2 AND2X2_3965 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3962_), .Y(w_mem_inst__abc_21203_new_n3963_));
AND2X2 AND2X2_3966 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_12__7_), .Y(w_mem_inst__abc_21203_new_n3966_));
AND2X2 AND2X2_3967 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_13__7_), .Y(w_mem_inst__abc_21203_new_n3967_));
AND2X2 AND2X2_3968 ( .A(round_ctr_rst), .B(\block[103] ), .Y(w_mem_inst__abc_21203_new_n3968_));
AND2X2 AND2X2_3969 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3968_), .Y(w_mem_inst__abc_21203_new_n3969_));
AND2X2 AND2X2_397 ( .A(_abc_15497_new_n1526_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n1527_));
AND2X2 AND2X2_3970 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_12__8_), .Y(w_mem_inst__abc_21203_new_n3972_));
AND2X2 AND2X2_3971 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_13__8_), .Y(w_mem_inst__abc_21203_new_n3973_));
AND2X2 AND2X2_3972 ( .A(round_ctr_rst), .B(\block[104] ), .Y(w_mem_inst__abc_21203_new_n3974_));
AND2X2 AND2X2_3973 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3974_), .Y(w_mem_inst__abc_21203_new_n3975_));
AND2X2 AND2X2_3974 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_12__9_), .Y(w_mem_inst__abc_21203_new_n3978_));
AND2X2 AND2X2_3975 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_13__9_), .Y(w_mem_inst__abc_21203_new_n3979_));
AND2X2 AND2X2_3976 ( .A(round_ctr_rst), .B(\block[105] ), .Y(w_mem_inst__abc_21203_new_n3980_));
AND2X2 AND2X2_3977 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3980_), .Y(w_mem_inst__abc_21203_new_n3981_));
AND2X2 AND2X2_3978 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_12__10_), .Y(w_mem_inst__abc_21203_new_n3984_));
AND2X2 AND2X2_3979 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_13__10_), .Y(w_mem_inst__abc_21203_new_n3985_));
AND2X2 AND2X2_398 ( .A(\digest[32] ), .B(d_reg_0_), .Y(_abc_15497_new_n1529_));
AND2X2 AND2X2_3980 ( .A(round_ctr_rst), .B(\block[106] ), .Y(w_mem_inst__abc_21203_new_n3986_));
AND2X2 AND2X2_3981 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3986_), .Y(w_mem_inst__abc_21203_new_n3987_));
AND2X2 AND2X2_3982 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_12__11_), .Y(w_mem_inst__abc_21203_new_n3990_));
AND2X2 AND2X2_3983 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_13__11_), .Y(w_mem_inst__abc_21203_new_n3991_));
AND2X2 AND2X2_3984 ( .A(round_ctr_rst), .B(\block[107] ), .Y(w_mem_inst__abc_21203_new_n3992_));
AND2X2 AND2X2_3985 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3992_), .Y(w_mem_inst__abc_21203_new_n3993_));
AND2X2 AND2X2_3986 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_12__12_), .Y(w_mem_inst__abc_21203_new_n3996_));
AND2X2 AND2X2_3987 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_13__12_), .Y(w_mem_inst__abc_21203_new_n3997_));
AND2X2 AND2X2_3988 ( .A(round_ctr_rst), .B(\block[108] ), .Y(w_mem_inst__abc_21203_new_n3998_));
AND2X2 AND2X2_3989 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n3998_), .Y(w_mem_inst__abc_21203_new_n3999_));
AND2X2 AND2X2_399 ( .A(_abc_15497_new_n1531_), .B(digest_update), .Y(_abc_15497_new_n1532_));
AND2X2 AND2X2_3990 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_12__13_), .Y(w_mem_inst__abc_21203_new_n4002_));
AND2X2 AND2X2_3991 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_13__13_), .Y(w_mem_inst__abc_21203_new_n4003_));
AND2X2 AND2X2_3992 ( .A(round_ctr_rst), .B(\block[109] ), .Y(w_mem_inst__abc_21203_new_n4004_));
AND2X2 AND2X2_3993 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4004_), .Y(w_mem_inst__abc_21203_new_n4005_));
AND2X2 AND2X2_3994 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_12__14_), .Y(w_mem_inst__abc_21203_new_n4008_));
AND2X2 AND2X2_3995 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_13__14_), .Y(w_mem_inst__abc_21203_new_n4009_));
AND2X2 AND2X2_3996 ( .A(round_ctr_rst), .B(\block[110] ), .Y(w_mem_inst__abc_21203_new_n4010_));
AND2X2 AND2X2_3997 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4010_), .Y(w_mem_inst__abc_21203_new_n4011_));
AND2X2 AND2X2_3998 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_12__15_), .Y(w_mem_inst__abc_21203_new_n4014_));
AND2X2 AND2X2_3999 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_13__15_), .Y(w_mem_inst__abc_21203_new_n4015_));
AND2X2 AND2X2_4 ( .A(c_reg_23_), .B(\digest[87] ), .Y(_abc_15497_new_n704_));
AND2X2 AND2X2_40 ( .A(_abc_15497_new_n776_), .B(_abc_15497_new_n766_), .Y(_abc_15497_new_n777_));
AND2X2 AND2X2_400 ( .A(_abc_15497_new_n1532_), .B(_abc_15497_new_n1530_), .Y(_abc_15497_new_n1533_));
AND2X2 AND2X2_4000 ( .A(round_ctr_rst), .B(\block[111] ), .Y(w_mem_inst__abc_21203_new_n4016_));
AND2X2 AND2X2_4001 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4016_), .Y(w_mem_inst__abc_21203_new_n4017_));
AND2X2 AND2X2_4002 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_12__16_), .Y(w_mem_inst__abc_21203_new_n4020_));
AND2X2 AND2X2_4003 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_13__16_), .Y(w_mem_inst__abc_21203_new_n4021_));
AND2X2 AND2X2_4004 ( .A(round_ctr_rst), .B(\block[112] ), .Y(w_mem_inst__abc_21203_new_n4022_));
AND2X2 AND2X2_4005 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4022_), .Y(w_mem_inst__abc_21203_new_n4023_));
AND2X2 AND2X2_4006 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_12__17_), .Y(w_mem_inst__abc_21203_new_n4026_));
AND2X2 AND2X2_4007 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_13__17_), .Y(w_mem_inst__abc_21203_new_n4027_));
AND2X2 AND2X2_4008 ( .A(round_ctr_rst), .B(\block[113] ), .Y(w_mem_inst__abc_21203_new_n4028_));
AND2X2 AND2X2_4009 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4028_), .Y(w_mem_inst__abc_21203_new_n4029_));
AND2X2 AND2X2_401 ( .A(_abc_15497_new_n701_), .B(\digest[32] ), .Y(_abc_15497_new_n1534_));
AND2X2 AND2X2_4010 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_12__18_), .Y(w_mem_inst__abc_21203_new_n4032_));
AND2X2 AND2X2_4011 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_13__18_), .Y(w_mem_inst__abc_21203_new_n4033_));
AND2X2 AND2X2_4012 ( .A(round_ctr_rst), .B(\block[114] ), .Y(w_mem_inst__abc_21203_new_n4034_));
AND2X2 AND2X2_4013 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4034_), .Y(w_mem_inst__abc_21203_new_n4035_));
AND2X2 AND2X2_4014 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_12__19_), .Y(w_mem_inst__abc_21203_new_n4038_));
AND2X2 AND2X2_4015 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_13__19_), .Y(w_mem_inst__abc_21203_new_n4039_));
AND2X2 AND2X2_4016 ( .A(round_ctr_rst), .B(\block[115] ), .Y(w_mem_inst__abc_21203_new_n4040_));
AND2X2 AND2X2_4017 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4040_), .Y(w_mem_inst__abc_21203_new_n4041_));
AND2X2 AND2X2_4018 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_12__20_), .Y(w_mem_inst__abc_21203_new_n4044_));
AND2X2 AND2X2_4019 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_13__20_), .Y(w_mem_inst__abc_21203_new_n4045_));
AND2X2 AND2X2_402 ( .A(\digest[33] ), .B(d_reg_1_), .Y(_abc_15497_new_n1537_));
AND2X2 AND2X2_4020 ( .A(round_ctr_rst), .B(\block[116] ), .Y(w_mem_inst__abc_21203_new_n4046_));
AND2X2 AND2X2_4021 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4046_), .Y(w_mem_inst__abc_21203_new_n4047_));
AND2X2 AND2X2_4022 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_12__21_), .Y(w_mem_inst__abc_21203_new_n4050_));
AND2X2 AND2X2_4023 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_13__21_), .Y(w_mem_inst__abc_21203_new_n4051_));
AND2X2 AND2X2_4024 ( .A(round_ctr_rst), .B(\block[117] ), .Y(w_mem_inst__abc_21203_new_n4052_));
AND2X2 AND2X2_4025 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4052_), .Y(w_mem_inst__abc_21203_new_n4053_));
AND2X2 AND2X2_4026 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_12__22_), .Y(w_mem_inst__abc_21203_new_n4056_));
AND2X2 AND2X2_4027 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_13__22_), .Y(w_mem_inst__abc_21203_new_n4057_));
AND2X2 AND2X2_4028 ( .A(round_ctr_rst), .B(\block[118] ), .Y(w_mem_inst__abc_21203_new_n4058_));
AND2X2 AND2X2_4029 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4058_), .Y(w_mem_inst__abc_21203_new_n4059_));
AND2X2 AND2X2_403 ( .A(_abc_15497_new_n1538_), .B(_abc_15497_new_n1536_), .Y(_abc_15497_new_n1539_));
AND2X2 AND2X2_4030 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_12__23_), .Y(w_mem_inst__abc_21203_new_n4062_));
AND2X2 AND2X2_4031 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_13__23_), .Y(w_mem_inst__abc_21203_new_n4063_));
AND2X2 AND2X2_4032 ( .A(round_ctr_rst), .B(\block[119] ), .Y(w_mem_inst__abc_21203_new_n4064_));
AND2X2 AND2X2_4033 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4064_), .Y(w_mem_inst__abc_21203_new_n4065_));
AND2X2 AND2X2_4034 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_12__24_), .Y(w_mem_inst__abc_21203_new_n4068_));
AND2X2 AND2X2_4035 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_13__24_), .Y(w_mem_inst__abc_21203_new_n4069_));
AND2X2 AND2X2_4036 ( .A(round_ctr_rst), .B(\block[120] ), .Y(w_mem_inst__abc_21203_new_n4070_));
AND2X2 AND2X2_4037 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4070_), .Y(w_mem_inst__abc_21203_new_n4071_));
AND2X2 AND2X2_4038 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_12__25_), .Y(w_mem_inst__abc_21203_new_n4074_));
AND2X2 AND2X2_4039 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_13__25_), .Y(w_mem_inst__abc_21203_new_n4075_));
AND2X2 AND2X2_404 ( .A(_abc_15497_new_n1539_), .B(_abc_15497_new_n1529_), .Y(_abc_15497_new_n1540_));
AND2X2 AND2X2_4040 ( .A(round_ctr_rst), .B(\block[121] ), .Y(w_mem_inst__abc_21203_new_n4076_));
AND2X2 AND2X2_4041 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4076_), .Y(w_mem_inst__abc_21203_new_n4077_));
AND2X2 AND2X2_4042 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_12__26_), .Y(w_mem_inst__abc_21203_new_n4080_));
AND2X2 AND2X2_4043 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_13__26_), .Y(w_mem_inst__abc_21203_new_n4081_));
AND2X2 AND2X2_4044 ( .A(round_ctr_rst), .B(\block[122] ), .Y(w_mem_inst__abc_21203_new_n4082_));
AND2X2 AND2X2_4045 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4082_), .Y(w_mem_inst__abc_21203_new_n4083_));
AND2X2 AND2X2_4046 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_12__27_), .Y(w_mem_inst__abc_21203_new_n4086_));
AND2X2 AND2X2_4047 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_13__27_), .Y(w_mem_inst__abc_21203_new_n4087_));
AND2X2 AND2X2_4048 ( .A(round_ctr_rst), .B(\block[123] ), .Y(w_mem_inst__abc_21203_new_n4088_));
AND2X2 AND2X2_4049 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4088_), .Y(w_mem_inst__abc_21203_new_n4089_));
AND2X2 AND2X2_405 ( .A(_abc_15497_new_n1541_), .B(_abc_15497_new_n1542_), .Y(_abc_15497_new_n1543_));
AND2X2 AND2X2_4050 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_12__28_), .Y(w_mem_inst__abc_21203_new_n4092_));
AND2X2 AND2X2_4051 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_13__28_), .Y(w_mem_inst__abc_21203_new_n4093_));
AND2X2 AND2X2_4052 ( .A(round_ctr_rst), .B(\block[124] ), .Y(w_mem_inst__abc_21203_new_n4094_));
AND2X2 AND2X2_4053 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4094_), .Y(w_mem_inst__abc_21203_new_n4095_));
AND2X2 AND2X2_4054 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_12__29_), .Y(w_mem_inst__abc_21203_new_n4098_));
AND2X2 AND2X2_4055 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_13__29_), .Y(w_mem_inst__abc_21203_new_n4099_));
AND2X2 AND2X2_4056 ( .A(round_ctr_rst), .B(\block[125] ), .Y(w_mem_inst__abc_21203_new_n4100_));
AND2X2 AND2X2_4057 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4100_), .Y(w_mem_inst__abc_21203_new_n4101_));
AND2X2 AND2X2_4058 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_12__30_), .Y(w_mem_inst__abc_21203_new_n4104_));
AND2X2 AND2X2_4059 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_13__30_), .Y(w_mem_inst__abc_21203_new_n4105_));
AND2X2 AND2X2_406 ( .A(_abc_15497_new_n1544_), .B(_abc_15497_new_n1546_), .Y(_0H3_reg_31_0__1_));
AND2X2 AND2X2_4060 ( .A(round_ctr_rst), .B(\block[126] ), .Y(w_mem_inst__abc_21203_new_n4106_));
AND2X2 AND2X2_4061 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4106_), .Y(w_mem_inst__abc_21203_new_n4107_));
AND2X2 AND2X2_4062 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_12__31_), .Y(w_mem_inst__abc_21203_new_n4110_));
AND2X2 AND2X2_4063 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_13__31_), .Y(w_mem_inst__abc_21203_new_n4111_));
AND2X2 AND2X2_4064 ( .A(round_ctr_rst), .B(\block[127] ), .Y(w_mem_inst__abc_21203_new_n4112_));
AND2X2 AND2X2_4065 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4112_), .Y(w_mem_inst__abc_21203_new_n4113_));
AND2X2 AND2X2_4066 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_11__0_), .Y(w_mem_inst__abc_21203_new_n4116_));
AND2X2 AND2X2_4067 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_12__0_), .Y(w_mem_inst__abc_21203_new_n4117_));
AND2X2 AND2X2_4068 ( .A(round_ctr_rst), .B(\block[128] ), .Y(w_mem_inst__abc_21203_new_n4118_));
AND2X2 AND2X2_4069 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4118_), .Y(w_mem_inst__abc_21203_new_n4119_));
AND2X2 AND2X2_407 ( .A(\digest[34] ), .B(d_reg_2_), .Y(_abc_15497_new_n1550_));
AND2X2 AND2X2_4070 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_11__1_), .Y(w_mem_inst__abc_21203_new_n4122_));
AND2X2 AND2X2_4071 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_12__1_), .Y(w_mem_inst__abc_21203_new_n4123_));
AND2X2 AND2X2_4072 ( .A(round_ctr_rst), .B(\block[129] ), .Y(w_mem_inst__abc_21203_new_n4124_));
AND2X2 AND2X2_4073 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4124_), .Y(w_mem_inst__abc_21203_new_n4125_));
AND2X2 AND2X2_4074 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_11__2_), .Y(w_mem_inst__abc_21203_new_n4128_));
AND2X2 AND2X2_4075 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_12__2_), .Y(w_mem_inst__abc_21203_new_n4129_));
AND2X2 AND2X2_4076 ( .A(round_ctr_rst), .B(\block[130] ), .Y(w_mem_inst__abc_21203_new_n4130_));
AND2X2 AND2X2_4077 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4130_), .Y(w_mem_inst__abc_21203_new_n4131_));
AND2X2 AND2X2_4078 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_11__3_), .Y(w_mem_inst__abc_21203_new_n4134_));
AND2X2 AND2X2_4079 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_12__3_), .Y(w_mem_inst__abc_21203_new_n4135_));
AND2X2 AND2X2_408 ( .A(_abc_15497_new_n1551_), .B(_abc_15497_new_n1549_), .Y(_abc_15497_new_n1552_));
AND2X2 AND2X2_4080 ( .A(round_ctr_rst), .B(\block[131] ), .Y(w_mem_inst__abc_21203_new_n4136_));
AND2X2 AND2X2_4081 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4136_), .Y(w_mem_inst__abc_21203_new_n4137_));
AND2X2 AND2X2_4082 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_11__4_), .Y(w_mem_inst__abc_21203_new_n4140_));
AND2X2 AND2X2_4083 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_12__4_), .Y(w_mem_inst__abc_21203_new_n4141_));
AND2X2 AND2X2_4084 ( .A(round_ctr_rst), .B(\block[132] ), .Y(w_mem_inst__abc_21203_new_n4142_));
AND2X2 AND2X2_4085 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4142_), .Y(w_mem_inst__abc_21203_new_n4143_));
AND2X2 AND2X2_4086 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_11__5_), .Y(w_mem_inst__abc_21203_new_n4146_));
AND2X2 AND2X2_4087 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_12__5_), .Y(w_mem_inst__abc_21203_new_n4147_));
AND2X2 AND2X2_4088 ( .A(round_ctr_rst), .B(\block[133] ), .Y(w_mem_inst__abc_21203_new_n4148_));
AND2X2 AND2X2_4089 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4148_), .Y(w_mem_inst__abc_21203_new_n4149_));
AND2X2 AND2X2_409 ( .A(_abc_15497_new_n1548_), .B(_abc_15497_new_n1552_), .Y(_abc_15497_new_n1553_));
AND2X2 AND2X2_4090 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_11__6_), .Y(w_mem_inst__abc_21203_new_n4152_));
AND2X2 AND2X2_4091 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_12__6_), .Y(w_mem_inst__abc_21203_new_n4153_));
AND2X2 AND2X2_4092 ( .A(round_ctr_rst), .B(\block[134] ), .Y(w_mem_inst__abc_21203_new_n4154_));
AND2X2 AND2X2_4093 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4154_), .Y(w_mem_inst__abc_21203_new_n4155_));
AND2X2 AND2X2_4094 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_11__7_), .Y(w_mem_inst__abc_21203_new_n4158_));
AND2X2 AND2X2_4095 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_12__7_), .Y(w_mem_inst__abc_21203_new_n4159_));
AND2X2 AND2X2_4096 ( .A(round_ctr_rst), .B(\block[135] ), .Y(w_mem_inst__abc_21203_new_n4160_));
AND2X2 AND2X2_4097 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4160_), .Y(w_mem_inst__abc_21203_new_n4161_));
AND2X2 AND2X2_4098 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_11__8_), .Y(w_mem_inst__abc_21203_new_n4164_));
AND2X2 AND2X2_4099 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_12__8_), .Y(w_mem_inst__abc_21203_new_n4165_));
AND2X2 AND2X2_41 ( .A(_abc_15497_new_n760_), .B(_abc_15497_new_n762_), .Y(_abc_15497_new_n778_));
AND2X2 AND2X2_410 ( .A(_abc_15497_new_n1554_), .B(_abc_15497_new_n1555_), .Y(_abc_15497_new_n1556_));
AND2X2 AND2X2_4100 ( .A(round_ctr_rst), .B(\block[136] ), .Y(w_mem_inst__abc_21203_new_n4166_));
AND2X2 AND2X2_4101 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4166_), .Y(w_mem_inst__abc_21203_new_n4167_));
AND2X2 AND2X2_4102 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_11__9_), .Y(w_mem_inst__abc_21203_new_n4170_));
AND2X2 AND2X2_4103 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_12__9_), .Y(w_mem_inst__abc_21203_new_n4171_));
AND2X2 AND2X2_4104 ( .A(round_ctr_rst), .B(\block[137] ), .Y(w_mem_inst__abc_21203_new_n4172_));
AND2X2 AND2X2_4105 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4172_), .Y(w_mem_inst__abc_21203_new_n4173_));
AND2X2 AND2X2_4106 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_11__10_), .Y(w_mem_inst__abc_21203_new_n4176_));
AND2X2 AND2X2_4107 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_12__10_), .Y(w_mem_inst__abc_21203_new_n4177_));
AND2X2 AND2X2_4108 ( .A(round_ctr_rst), .B(\block[138] ), .Y(w_mem_inst__abc_21203_new_n4178_));
AND2X2 AND2X2_4109 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4178_), .Y(w_mem_inst__abc_21203_new_n4179_));
AND2X2 AND2X2_411 ( .A(_abc_15497_new_n1557_), .B(_abc_15497_new_n1559_), .Y(_0H3_reg_31_0__2_));
AND2X2 AND2X2_4110 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_11__11_), .Y(w_mem_inst__abc_21203_new_n4182_));
AND2X2 AND2X2_4111 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_12__11_), .Y(w_mem_inst__abc_21203_new_n4183_));
AND2X2 AND2X2_4112 ( .A(round_ctr_rst), .B(\block[139] ), .Y(w_mem_inst__abc_21203_new_n4184_));
AND2X2 AND2X2_4113 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4184_), .Y(w_mem_inst__abc_21203_new_n4185_));
AND2X2 AND2X2_4114 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_11__12_), .Y(w_mem_inst__abc_21203_new_n4188_));
AND2X2 AND2X2_4115 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_12__12_), .Y(w_mem_inst__abc_21203_new_n4189_));
AND2X2 AND2X2_4116 ( .A(round_ctr_rst), .B(\block[140] ), .Y(w_mem_inst__abc_21203_new_n4190_));
AND2X2 AND2X2_4117 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4190_), .Y(w_mem_inst__abc_21203_new_n4191_));
AND2X2 AND2X2_4118 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_11__13_), .Y(w_mem_inst__abc_21203_new_n4194_));
AND2X2 AND2X2_4119 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_12__13_), .Y(w_mem_inst__abc_21203_new_n4195_));
AND2X2 AND2X2_412 ( .A(_abc_15497_new_n701_), .B(\digest[35] ), .Y(_abc_15497_new_n1561_));
AND2X2 AND2X2_4120 ( .A(round_ctr_rst), .B(\block[141] ), .Y(w_mem_inst__abc_21203_new_n4196_));
AND2X2 AND2X2_4121 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4196_), .Y(w_mem_inst__abc_21203_new_n4197_));
AND2X2 AND2X2_4122 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_11__14_), .Y(w_mem_inst__abc_21203_new_n4200_));
AND2X2 AND2X2_4123 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_12__14_), .Y(w_mem_inst__abc_21203_new_n4201_));
AND2X2 AND2X2_4124 ( .A(round_ctr_rst), .B(\block[142] ), .Y(w_mem_inst__abc_21203_new_n4202_));
AND2X2 AND2X2_4125 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4202_), .Y(w_mem_inst__abc_21203_new_n4203_));
AND2X2 AND2X2_4126 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_11__15_), .Y(w_mem_inst__abc_21203_new_n4206_));
AND2X2 AND2X2_4127 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_12__15_), .Y(w_mem_inst__abc_21203_new_n4207_));
AND2X2 AND2X2_4128 ( .A(round_ctr_rst), .B(\block[143] ), .Y(w_mem_inst__abc_21203_new_n4208_));
AND2X2 AND2X2_4129 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4208_), .Y(w_mem_inst__abc_21203_new_n4209_));
AND2X2 AND2X2_413 ( .A(\digest[35] ), .B(d_reg_3_), .Y(_abc_15497_new_n1564_));
AND2X2 AND2X2_4130 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_11__16_), .Y(w_mem_inst__abc_21203_new_n4212_));
AND2X2 AND2X2_4131 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_12__16_), .Y(w_mem_inst__abc_21203_new_n4213_));
AND2X2 AND2X2_4132 ( .A(round_ctr_rst), .B(\block[144] ), .Y(w_mem_inst__abc_21203_new_n4214_));
AND2X2 AND2X2_4133 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4214_), .Y(w_mem_inst__abc_21203_new_n4215_));
AND2X2 AND2X2_4134 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_11__17_), .Y(w_mem_inst__abc_21203_new_n4218_));
AND2X2 AND2X2_4135 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_12__17_), .Y(w_mem_inst__abc_21203_new_n4219_));
AND2X2 AND2X2_4136 ( .A(round_ctr_rst), .B(\block[145] ), .Y(w_mem_inst__abc_21203_new_n4220_));
AND2X2 AND2X2_4137 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4220_), .Y(w_mem_inst__abc_21203_new_n4221_));
AND2X2 AND2X2_4138 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_11__18_), .Y(w_mem_inst__abc_21203_new_n4224_));
AND2X2 AND2X2_4139 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_12__18_), .Y(w_mem_inst__abc_21203_new_n4225_));
AND2X2 AND2X2_414 ( .A(_abc_15497_new_n1565_), .B(_abc_15497_new_n1563_), .Y(_abc_15497_new_n1566_));
AND2X2 AND2X2_4140 ( .A(round_ctr_rst), .B(\block[146] ), .Y(w_mem_inst__abc_21203_new_n4226_));
AND2X2 AND2X2_4141 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4226_), .Y(w_mem_inst__abc_21203_new_n4227_));
AND2X2 AND2X2_4142 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_11__19_), .Y(w_mem_inst__abc_21203_new_n4230_));
AND2X2 AND2X2_4143 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_12__19_), .Y(w_mem_inst__abc_21203_new_n4231_));
AND2X2 AND2X2_4144 ( .A(round_ctr_rst), .B(\block[147] ), .Y(w_mem_inst__abc_21203_new_n4232_));
AND2X2 AND2X2_4145 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4232_), .Y(w_mem_inst__abc_21203_new_n4233_));
AND2X2 AND2X2_4146 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_11__20_), .Y(w_mem_inst__abc_21203_new_n4236_));
AND2X2 AND2X2_4147 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_12__20_), .Y(w_mem_inst__abc_21203_new_n4237_));
AND2X2 AND2X2_4148 ( .A(round_ctr_rst), .B(\block[148] ), .Y(w_mem_inst__abc_21203_new_n4238_));
AND2X2 AND2X2_4149 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4238_), .Y(w_mem_inst__abc_21203_new_n4239_));
AND2X2 AND2X2_415 ( .A(_abc_15497_new_n1570_), .B(_abc_15497_new_n1567_), .Y(_abc_15497_new_n1571_));
AND2X2 AND2X2_4150 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_11__21_), .Y(w_mem_inst__abc_21203_new_n4242_));
AND2X2 AND2X2_4151 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_12__21_), .Y(w_mem_inst__abc_21203_new_n4243_));
AND2X2 AND2X2_4152 ( .A(round_ctr_rst), .B(\block[149] ), .Y(w_mem_inst__abc_21203_new_n4244_));
AND2X2 AND2X2_4153 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4244_), .Y(w_mem_inst__abc_21203_new_n4245_));
AND2X2 AND2X2_4154 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_11__22_), .Y(w_mem_inst__abc_21203_new_n4248_));
AND2X2 AND2X2_4155 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_12__22_), .Y(w_mem_inst__abc_21203_new_n4249_));
AND2X2 AND2X2_4156 ( .A(round_ctr_rst), .B(\block[150] ), .Y(w_mem_inst__abc_21203_new_n4250_));
AND2X2 AND2X2_4157 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4250_), .Y(w_mem_inst__abc_21203_new_n4251_));
AND2X2 AND2X2_4158 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_11__23_), .Y(w_mem_inst__abc_21203_new_n4254_));
AND2X2 AND2X2_4159 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_12__23_), .Y(w_mem_inst__abc_21203_new_n4255_));
AND2X2 AND2X2_416 ( .A(_abc_15497_new_n1571_), .B(digest_update), .Y(_abc_15497_new_n1572_));
AND2X2 AND2X2_4160 ( .A(round_ctr_rst), .B(\block[151] ), .Y(w_mem_inst__abc_21203_new_n4256_));
AND2X2 AND2X2_4161 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4256_), .Y(w_mem_inst__abc_21203_new_n4257_));
AND2X2 AND2X2_4162 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_11__24_), .Y(w_mem_inst__abc_21203_new_n4260_));
AND2X2 AND2X2_4163 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_12__24_), .Y(w_mem_inst__abc_21203_new_n4261_));
AND2X2 AND2X2_4164 ( .A(round_ctr_rst), .B(\block[152] ), .Y(w_mem_inst__abc_21203_new_n4262_));
AND2X2 AND2X2_4165 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4262_), .Y(w_mem_inst__abc_21203_new_n4263_));
AND2X2 AND2X2_4166 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_11__25_), .Y(w_mem_inst__abc_21203_new_n4266_));
AND2X2 AND2X2_4167 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_12__25_), .Y(w_mem_inst__abc_21203_new_n4267_));
AND2X2 AND2X2_4168 ( .A(round_ctr_rst), .B(\block[153] ), .Y(w_mem_inst__abc_21203_new_n4268_));
AND2X2 AND2X2_4169 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4268_), .Y(w_mem_inst__abc_21203_new_n4269_));
AND2X2 AND2X2_417 ( .A(\digest[36] ), .B(d_reg_4_), .Y(_abc_15497_new_n1575_));
AND2X2 AND2X2_4170 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_11__26_), .Y(w_mem_inst__abc_21203_new_n4272_));
AND2X2 AND2X2_4171 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_12__26_), .Y(w_mem_inst__abc_21203_new_n4273_));
AND2X2 AND2X2_4172 ( .A(round_ctr_rst), .B(\block[154] ), .Y(w_mem_inst__abc_21203_new_n4274_));
AND2X2 AND2X2_4173 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4274_), .Y(w_mem_inst__abc_21203_new_n4275_));
AND2X2 AND2X2_4174 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_11__27_), .Y(w_mem_inst__abc_21203_new_n4278_));
AND2X2 AND2X2_4175 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_12__27_), .Y(w_mem_inst__abc_21203_new_n4279_));
AND2X2 AND2X2_4176 ( .A(round_ctr_rst), .B(\block[155] ), .Y(w_mem_inst__abc_21203_new_n4280_));
AND2X2 AND2X2_4177 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4280_), .Y(w_mem_inst__abc_21203_new_n4281_));
AND2X2 AND2X2_4178 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_11__28_), .Y(w_mem_inst__abc_21203_new_n4284_));
AND2X2 AND2X2_4179 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_12__28_), .Y(w_mem_inst__abc_21203_new_n4285_));
AND2X2 AND2X2_418 ( .A(_abc_15497_new_n1576_), .B(_abc_15497_new_n1574_), .Y(_abc_15497_new_n1577_));
AND2X2 AND2X2_4180 ( .A(round_ctr_rst), .B(\block[156] ), .Y(w_mem_inst__abc_21203_new_n4286_));
AND2X2 AND2X2_4181 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4286_), .Y(w_mem_inst__abc_21203_new_n4287_));
AND2X2 AND2X2_4182 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_11__29_), .Y(w_mem_inst__abc_21203_new_n4290_));
AND2X2 AND2X2_4183 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_12__29_), .Y(w_mem_inst__abc_21203_new_n4291_));
AND2X2 AND2X2_4184 ( .A(round_ctr_rst), .B(\block[157] ), .Y(w_mem_inst__abc_21203_new_n4292_));
AND2X2 AND2X2_4185 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4292_), .Y(w_mem_inst__abc_21203_new_n4293_));
AND2X2 AND2X2_4186 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_11__30_), .Y(w_mem_inst__abc_21203_new_n4296_));
AND2X2 AND2X2_4187 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_12__30_), .Y(w_mem_inst__abc_21203_new_n4297_));
AND2X2 AND2X2_4188 ( .A(round_ctr_rst), .B(\block[158] ), .Y(w_mem_inst__abc_21203_new_n4298_));
AND2X2 AND2X2_4189 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4298_), .Y(w_mem_inst__abc_21203_new_n4299_));
AND2X2 AND2X2_419 ( .A(_abc_15497_new_n1562_), .B(_abc_15497_new_n1563_), .Y(_abc_15497_new_n1578_));
AND2X2 AND2X2_4190 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_11__31_), .Y(w_mem_inst__abc_21203_new_n4302_));
AND2X2 AND2X2_4191 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_12__31_), .Y(w_mem_inst__abc_21203_new_n4303_));
AND2X2 AND2X2_4192 ( .A(round_ctr_rst), .B(\block[159] ), .Y(w_mem_inst__abc_21203_new_n4304_));
AND2X2 AND2X2_4193 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4304_), .Y(w_mem_inst__abc_21203_new_n4305_));
AND2X2 AND2X2_4194 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_7__0_), .Y(w_mem_inst__abc_21203_new_n4308_));
AND2X2 AND2X2_4195 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_8__0_), .Y(w_mem_inst__abc_21203_new_n4309_));
AND2X2 AND2X2_4196 ( .A(round_ctr_rst), .B(\block[256] ), .Y(w_mem_inst__abc_21203_new_n4310_));
AND2X2 AND2X2_4197 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4310_), .Y(w_mem_inst__abc_21203_new_n4311_));
AND2X2 AND2X2_4198 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_7__1_), .Y(w_mem_inst__abc_21203_new_n4314_));
AND2X2 AND2X2_4199 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_8__1_), .Y(w_mem_inst__abc_21203_new_n4315_));
AND2X2 AND2X2_42 ( .A(_abc_15497_new_n770_), .B(_abc_15497_new_n781_), .Y(_abc_15497_new_n782_));
AND2X2 AND2X2_420 ( .A(_abc_15497_new_n1579_), .B(_abc_15497_new_n1577_), .Y(_abc_15497_new_n1580_));
AND2X2 AND2X2_4200 ( .A(round_ctr_rst), .B(\block[257] ), .Y(w_mem_inst__abc_21203_new_n4316_));
AND2X2 AND2X2_4201 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4316_), .Y(w_mem_inst__abc_21203_new_n4317_));
AND2X2 AND2X2_4202 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_7__2_), .Y(w_mem_inst__abc_21203_new_n4320_));
AND2X2 AND2X2_4203 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_8__2_), .Y(w_mem_inst__abc_21203_new_n4321_));
AND2X2 AND2X2_4204 ( .A(round_ctr_rst), .B(\block[258] ), .Y(w_mem_inst__abc_21203_new_n4322_));
AND2X2 AND2X2_4205 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4322_), .Y(w_mem_inst__abc_21203_new_n4323_));
AND2X2 AND2X2_4206 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_7__3_), .Y(w_mem_inst__abc_21203_new_n4326_));
AND2X2 AND2X2_4207 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_8__3_), .Y(w_mem_inst__abc_21203_new_n4327_));
AND2X2 AND2X2_4208 ( .A(round_ctr_rst), .B(\block[259] ), .Y(w_mem_inst__abc_21203_new_n4328_));
AND2X2 AND2X2_4209 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4328_), .Y(w_mem_inst__abc_21203_new_n4329_));
AND2X2 AND2X2_421 ( .A(_abc_15497_new_n1581_), .B(_abc_15497_new_n1582_), .Y(_abc_15497_new_n1583_));
AND2X2 AND2X2_4210 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_7__4_), .Y(w_mem_inst__abc_21203_new_n4332_));
AND2X2 AND2X2_4211 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_8__4_), .Y(w_mem_inst__abc_21203_new_n4333_));
AND2X2 AND2X2_4212 ( .A(round_ctr_rst), .B(\block[260] ), .Y(w_mem_inst__abc_21203_new_n4334_));
AND2X2 AND2X2_4213 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4334_), .Y(w_mem_inst__abc_21203_new_n4335_));
AND2X2 AND2X2_4214 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_7__5_), .Y(w_mem_inst__abc_21203_new_n4338_));
AND2X2 AND2X2_4215 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_8__5_), .Y(w_mem_inst__abc_21203_new_n4339_));
AND2X2 AND2X2_4216 ( .A(round_ctr_rst), .B(\block[261] ), .Y(w_mem_inst__abc_21203_new_n4340_));
AND2X2 AND2X2_4217 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4340_), .Y(w_mem_inst__abc_21203_new_n4341_));
AND2X2 AND2X2_4218 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_7__6_), .Y(w_mem_inst__abc_21203_new_n4344_));
AND2X2 AND2X2_4219 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_8__6_), .Y(w_mem_inst__abc_21203_new_n4345_));
AND2X2 AND2X2_422 ( .A(_abc_15497_new_n1584_), .B(_abc_15497_new_n1586_), .Y(_0H3_reg_31_0__4_));
AND2X2 AND2X2_4220 ( .A(round_ctr_rst), .B(\block[262] ), .Y(w_mem_inst__abc_21203_new_n4346_));
AND2X2 AND2X2_4221 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4346_), .Y(w_mem_inst__abc_21203_new_n4347_));
AND2X2 AND2X2_4222 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_7__7_), .Y(w_mem_inst__abc_21203_new_n4350_));
AND2X2 AND2X2_4223 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_8__7_), .Y(w_mem_inst__abc_21203_new_n4351_));
AND2X2 AND2X2_4224 ( .A(round_ctr_rst), .B(\block[263] ), .Y(w_mem_inst__abc_21203_new_n4352_));
AND2X2 AND2X2_4225 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4352_), .Y(w_mem_inst__abc_21203_new_n4353_));
AND2X2 AND2X2_4226 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_7__8_), .Y(w_mem_inst__abc_21203_new_n4356_));
AND2X2 AND2X2_4227 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_8__8_), .Y(w_mem_inst__abc_21203_new_n4357_));
AND2X2 AND2X2_4228 ( .A(round_ctr_rst), .B(\block[264] ), .Y(w_mem_inst__abc_21203_new_n4358_));
AND2X2 AND2X2_4229 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4358_), .Y(w_mem_inst__abc_21203_new_n4359_));
AND2X2 AND2X2_423 ( .A(\digest[37] ), .B(d_reg_5_), .Y(_abc_15497_new_n1590_));
AND2X2 AND2X2_4230 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_7__9_), .Y(w_mem_inst__abc_21203_new_n4362_));
AND2X2 AND2X2_4231 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_8__9_), .Y(w_mem_inst__abc_21203_new_n4363_));
AND2X2 AND2X2_4232 ( .A(round_ctr_rst), .B(\block[265] ), .Y(w_mem_inst__abc_21203_new_n4364_));
AND2X2 AND2X2_4233 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4364_), .Y(w_mem_inst__abc_21203_new_n4365_));
AND2X2 AND2X2_4234 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_7__10_), .Y(w_mem_inst__abc_21203_new_n4368_));
AND2X2 AND2X2_4235 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_8__10_), .Y(w_mem_inst__abc_21203_new_n4369_));
AND2X2 AND2X2_4236 ( .A(round_ctr_rst), .B(\block[266] ), .Y(w_mem_inst__abc_21203_new_n4370_));
AND2X2 AND2X2_4237 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4370_), .Y(w_mem_inst__abc_21203_new_n4371_));
AND2X2 AND2X2_4238 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_7__11_), .Y(w_mem_inst__abc_21203_new_n4374_));
AND2X2 AND2X2_4239 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_8__11_), .Y(w_mem_inst__abc_21203_new_n4375_));
AND2X2 AND2X2_424 ( .A(_abc_15497_new_n1591_), .B(_abc_15497_new_n1589_), .Y(_abc_15497_new_n1592_));
AND2X2 AND2X2_4240 ( .A(round_ctr_rst), .B(\block[267] ), .Y(w_mem_inst__abc_21203_new_n4376_));
AND2X2 AND2X2_4241 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4376_), .Y(w_mem_inst__abc_21203_new_n4377_));
AND2X2 AND2X2_4242 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_7__12_), .Y(w_mem_inst__abc_21203_new_n4380_));
AND2X2 AND2X2_4243 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_8__12_), .Y(w_mem_inst__abc_21203_new_n4381_));
AND2X2 AND2X2_4244 ( .A(round_ctr_rst), .B(\block[268] ), .Y(w_mem_inst__abc_21203_new_n4382_));
AND2X2 AND2X2_4245 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4382_), .Y(w_mem_inst__abc_21203_new_n4383_));
AND2X2 AND2X2_4246 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_7__13_), .Y(w_mem_inst__abc_21203_new_n4386_));
AND2X2 AND2X2_4247 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_8__13_), .Y(w_mem_inst__abc_21203_new_n4387_));
AND2X2 AND2X2_4248 ( .A(round_ctr_rst), .B(\block[269] ), .Y(w_mem_inst__abc_21203_new_n4388_));
AND2X2 AND2X2_4249 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4388_), .Y(w_mem_inst__abc_21203_new_n4389_));
AND2X2 AND2X2_425 ( .A(_abc_15497_new_n1588_), .B(_abc_15497_new_n1592_), .Y(_abc_15497_new_n1594_));
AND2X2 AND2X2_4250 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_7__14_), .Y(w_mem_inst__abc_21203_new_n4392_));
AND2X2 AND2X2_4251 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_8__14_), .Y(w_mem_inst__abc_21203_new_n4393_));
AND2X2 AND2X2_4252 ( .A(round_ctr_rst), .B(\block[270] ), .Y(w_mem_inst__abc_21203_new_n4394_));
AND2X2 AND2X2_4253 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4394_), .Y(w_mem_inst__abc_21203_new_n4395_));
AND2X2 AND2X2_4254 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_7__15_), .Y(w_mem_inst__abc_21203_new_n4398_));
AND2X2 AND2X2_4255 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_8__15_), .Y(w_mem_inst__abc_21203_new_n4399_));
AND2X2 AND2X2_4256 ( .A(round_ctr_rst), .B(\block[271] ), .Y(w_mem_inst__abc_21203_new_n4400_));
AND2X2 AND2X2_4257 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4400_), .Y(w_mem_inst__abc_21203_new_n4401_));
AND2X2 AND2X2_4258 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_7__16_), .Y(w_mem_inst__abc_21203_new_n4404_));
AND2X2 AND2X2_4259 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_8__16_), .Y(w_mem_inst__abc_21203_new_n4405_));
AND2X2 AND2X2_426 ( .A(_abc_15497_new_n1595_), .B(_abc_15497_new_n1593_), .Y(_abc_15497_new_n1596_));
AND2X2 AND2X2_4260 ( .A(round_ctr_rst), .B(\block[272] ), .Y(w_mem_inst__abc_21203_new_n4406_));
AND2X2 AND2X2_4261 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4406_), .Y(w_mem_inst__abc_21203_new_n4407_));
AND2X2 AND2X2_4262 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_7__17_), .Y(w_mem_inst__abc_21203_new_n4410_));
AND2X2 AND2X2_4263 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_8__17_), .Y(w_mem_inst__abc_21203_new_n4411_));
AND2X2 AND2X2_4264 ( .A(round_ctr_rst), .B(\block[273] ), .Y(w_mem_inst__abc_21203_new_n4412_));
AND2X2 AND2X2_4265 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4412_), .Y(w_mem_inst__abc_21203_new_n4413_));
AND2X2 AND2X2_4266 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_7__18_), .Y(w_mem_inst__abc_21203_new_n4416_));
AND2X2 AND2X2_4267 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_8__18_), .Y(w_mem_inst__abc_21203_new_n4417_));
AND2X2 AND2X2_4268 ( .A(round_ctr_rst), .B(\block[274] ), .Y(w_mem_inst__abc_21203_new_n4418_));
AND2X2 AND2X2_4269 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4418_), .Y(w_mem_inst__abc_21203_new_n4419_));
AND2X2 AND2X2_427 ( .A(_abc_15497_new_n1596_), .B(digest_update), .Y(_abc_15497_new_n1597_));
AND2X2 AND2X2_4270 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_7__19_), .Y(w_mem_inst__abc_21203_new_n4422_));
AND2X2 AND2X2_4271 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_8__19_), .Y(w_mem_inst__abc_21203_new_n4423_));
AND2X2 AND2X2_4272 ( .A(round_ctr_rst), .B(\block[275] ), .Y(w_mem_inst__abc_21203_new_n4424_));
AND2X2 AND2X2_4273 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4424_), .Y(w_mem_inst__abc_21203_new_n4425_));
AND2X2 AND2X2_4274 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_7__20_), .Y(w_mem_inst__abc_21203_new_n4428_));
AND2X2 AND2X2_4275 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_8__20_), .Y(w_mem_inst__abc_21203_new_n4429_));
AND2X2 AND2X2_4276 ( .A(round_ctr_rst), .B(\block[276] ), .Y(w_mem_inst__abc_21203_new_n4430_));
AND2X2 AND2X2_4277 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4430_), .Y(w_mem_inst__abc_21203_new_n4431_));
AND2X2 AND2X2_4278 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_7__21_), .Y(w_mem_inst__abc_21203_new_n4434_));
AND2X2 AND2X2_4279 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_8__21_), .Y(w_mem_inst__abc_21203_new_n4435_));
AND2X2 AND2X2_428 ( .A(_abc_15497_new_n1598_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n1599_));
AND2X2 AND2X2_4280 ( .A(round_ctr_rst), .B(\block[277] ), .Y(w_mem_inst__abc_21203_new_n4436_));
AND2X2 AND2X2_4281 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4436_), .Y(w_mem_inst__abc_21203_new_n4437_));
AND2X2 AND2X2_4282 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_7__22_), .Y(w_mem_inst__abc_21203_new_n4440_));
AND2X2 AND2X2_4283 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_8__22_), .Y(w_mem_inst__abc_21203_new_n4441_));
AND2X2 AND2X2_4284 ( .A(round_ctr_rst), .B(\block[278] ), .Y(w_mem_inst__abc_21203_new_n4442_));
AND2X2 AND2X2_4285 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4442_), .Y(w_mem_inst__abc_21203_new_n4443_));
AND2X2 AND2X2_4286 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_7__23_), .Y(w_mem_inst__abc_21203_new_n4446_));
AND2X2 AND2X2_4287 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_8__23_), .Y(w_mem_inst__abc_21203_new_n4447_));
AND2X2 AND2X2_4288 ( .A(round_ctr_rst), .B(\block[279] ), .Y(w_mem_inst__abc_21203_new_n4448_));
AND2X2 AND2X2_4289 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4448_), .Y(w_mem_inst__abc_21203_new_n4449_));
AND2X2 AND2X2_429 ( .A(\digest[38] ), .B(d_reg_6_), .Y(_abc_15497_new_n1603_));
AND2X2 AND2X2_4290 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_7__24_), .Y(w_mem_inst__abc_21203_new_n4452_));
AND2X2 AND2X2_4291 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_8__24_), .Y(w_mem_inst__abc_21203_new_n4453_));
AND2X2 AND2X2_4292 ( .A(round_ctr_rst), .B(\block[280] ), .Y(w_mem_inst__abc_21203_new_n4454_));
AND2X2 AND2X2_4293 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4454_), .Y(w_mem_inst__abc_21203_new_n4455_));
AND2X2 AND2X2_4294 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_7__25_), .Y(w_mem_inst__abc_21203_new_n4458_));
AND2X2 AND2X2_4295 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_8__25_), .Y(w_mem_inst__abc_21203_new_n4459_));
AND2X2 AND2X2_4296 ( .A(round_ctr_rst), .B(\block[281] ), .Y(w_mem_inst__abc_21203_new_n4460_));
AND2X2 AND2X2_4297 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4460_), .Y(w_mem_inst__abc_21203_new_n4461_));
AND2X2 AND2X2_4298 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_7__26_), .Y(w_mem_inst__abc_21203_new_n4464_));
AND2X2 AND2X2_4299 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_8__26_), .Y(w_mem_inst__abc_21203_new_n4465_));
AND2X2 AND2X2_43 ( .A(_abc_15497_new_n772_), .B(_abc_15497_new_n782_), .Y(_abc_15497_new_n783_));
AND2X2 AND2X2_430 ( .A(_abc_15497_new_n1604_), .B(_abc_15497_new_n1602_), .Y(_abc_15497_new_n1605_));
AND2X2 AND2X2_4300 ( .A(round_ctr_rst), .B(\block[282] ), .Y(w_mem_inst__abc_21203_new_n4466_));
AND2X2 AND2X2_4301 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4466_), .Y(w_mem_inst__abc_21203_new_n4467_));
AND2X2 AND2X2_4302 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_7__27_), .Y(w_mem_inst__abc_21203_new_n4470_));
AND2X2 AND2X2_4303 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_8__27_), .Y(w_mem_inst__abc_21203_new_n4471_));
AND2X2 AND2X2_4304 ( .A(round_ctr_rst), .B(\block[283] ), .Y(w_mem_inst__abc_21203_new_n4472_));
AND2X2 AND2X2_4305 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4472_), .Y(w_mem_inst__abc_21203_new_n4473_));
AND2X2 AND2X2_4306 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_7__28_), .Y(w_mem_inst__abc_21203_new_n4476_));
AND2X2 AND2X2_4307 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_8__28_), .Y(w_mem_inst__abc_21203_new_n4477_));
AND2X2 AND2X2_4308 ( .A(round_ctr_rst), .B(\block[284] ), .Y(w_mem_inst__abc_21203_new_n4478_));
AND2X2 AND2X2_4309 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4478_), .Y(w_mem_inst__abc_21203_new_n4479_));
AND2X2 AND2X2_431 ( .A(_abc_15497_new_n1601_), .B(_abc_15497_new_n1605_), .Y(_abc_15497_new_n1607_));
AND2X2 AND2X2_4310 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_7__29_), .Y(w_mem_inst__abc_21203_new_n4482_));
AND2X2 AND2X2_4311 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_8__29_), .Y(w_mem_inst__abc_21203_new_n4483_));
AND2X2 AND2X2_4312 ( .A(round_ctr_rst), .B(\block[285] ), .Y(w_mem_inst__abc_21203_new_n4484_));
AND2X2 AND2X2_4313 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4484_), .Y(w_mem_inst__abc_21203_new_n4485_));
AND2X2 AND2X2_4314 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_7__30_), .Y(w_mem_inst__abc_21203_new_n4488_));
AND2X2 AND2X2_4315 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_8__30_), .Y(w_mem_inst__abc_21203_new_n4489_));
AND2X2 AND2X2_4316 ( .A(round_ctr_rst), .B(\block[286] ), .Y(w_mem_inst__abc_21203_new_n4490_));
AND2X2 AND2X2_4317 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4490_), .Y(w_mem_inst__abc_21203_new_n4491_));
AND2X2 AND2X2_4318 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_7__31_), .Y(w_mem_inst__abc_21203_new_n4494_));
AND2X2 AND2X2_4319 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_8__31_), .Y(w_mem_inst__abc_21203_new_n4495_));
AND2X2 AND2X2_432 ( .A(_abc_15497_new_n1608_), .B(_abc_15497_new_n1606_), .Y(_abc_15497_new_n1609_));
AND2X2 AND2X2_4320 ( .A(round_ctr_rst), .B(\block[287] ), .Y(w_mem_inst__abc_21203_new_n4496_));
AND2X2 AND2X2_4321 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4496_), .Y(w_mem_inst__abc_21203_new_n4497_));
AND2X2 AND2X2_4322 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_9__0_), .Y(w_mem_inst__abc_21203_new_n4500_));
AND2X2 AND2X2_4323 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_10__0_), .Y(w_mem_inst__abc_21203_new_n4501_));
AND2X2 AND2X2_4324 ( .A(round_ctr_rst), .B(\block[192] ), .Y(w_mem_inst__abc_21203_new_n4502_));
AND2X2 AND2X2_4325 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4502_), .Y(w_mem_inst__abc_21203_new_n4503_));
AND2X2 AND2X2_4326 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_9__1_), .Y(w_mem_inst__abc_21203_new_n4506_));
AND2X2 AND2X2_4327 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_10__1_), .Y(w_mem_inst__abc_21203_new_n4507_));
AND2X2 AND2X2_4328 ( .A(round_ctr_rst), .B(\block[193] ), .Y(w_mem_inst__abc_21203_new_n4508_));
AND2X2 AND2X2_4329 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4508_), .Y(w_mem_inst__abc_21203_new_n4509_));
AND2X2 AND2X2_433 ( .A(_abc_15497_new_n1609_), .B(digest_update), .Y(_abc_15497_new_n1610_));
AND2X2 AND2X2_4330 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_9__2_), .Y(w_mem_inst__abc_21203_new_n4512_));
AND2X2 AND2X2_4331 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_10__2_), .Y(w_mem_inst__abc_21203_new_n4513_));
AND2X2 AND2X2_4332 ( .A(round_ctr_rst), .B(\block[194] ), .Y(w_mem_inst__abc_21203_new_n4514_));
AND2X2 AND2X2_4333 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4514_), .Y(w_mem_inst__abc_21203_new_n4515_));
AND2X2 AND2X2_4334 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_9__3_), .Y(w_mem_inst__abc_21203_new_n4518_));
AND2X2 AND2X2_4335 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_10__3_), .Y(w_mem_inst__abc_21203_new_n4519_));
AND2X2 AND2X2_4336 ( .A(round_ctr_rst), .B(\block[195] ), .Y(w_mem_inst__abc_21203_new_n4520_));
AND2X2 AND2X2_4337 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4520_), .Y(w_mem_inst__abc_21203_new_n4521_));
AND2X2 AND2X2_4338 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_9__4_), .Y(w_mem_inst__abc_21203_new_n4524_));
AND2X2 AND2X2_4339 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_10__4_), .Y(w_mem_inst__abc_21203_new_n4525_));
AND2X2 AND2X2_434 ( .A(_abc_15497_new_n1611_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n1612_));
AND2X2 AND2X2_4340 ( .A(round_ctr_rst), .B(\block[196] ), .Y(w_mem_inst__abc_21203_new_n4526_));
AND2X2 AND2X2_4341 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4526_), .Y(w_mem_inst__abc_21203_new_n4527_));
AND2X2 AND2X2_4342 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_9__5_), .Y(w_mem_inst__abc_21203_new_n4530_));
AND2X2 AND2X2_4343 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_10__5_), .Y(w_mem_inst__abc_21203_new_n4531_));
AND2X2 AND2X2_4344 ( .A(round_ctr_rst), .B(\block[197] ), .Y(w_mem_inst__abc_21203_new_n4532_));
AND2X2 AND2X2_4345 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4532_), .Y(w_mem_inst__abc_21203_new_n4533_));
AND2X2 AND2X2_4346 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_9__6_), .Y(w_mem_inst__abc_21203_new_n4536_));
AND2X2 AND2X2_4347 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_10__6_), .Y(w_mem_inst__abc_21203_new_n4537_));
AND2X2 AND2X2_4348 ( .A(round_ctr_rst), .B(\block[198] ), .Y(w_mem_inst__abc_21203_new_n4538_));
AND2X2 AND2X2_4349 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4538_), .Y(w_mem_inst__abc_21203_new_n4539_));
AND2X2 AND2X2_435 ( .A(_abc_15497_new_n701_), .B(\digest[39] ), .Y(_abc_15497_new_n1614_));
AND2X2 AND2X2_4350 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_9__7_), .Y(w_mem_inst__abc_21203_new_n4542_));
AND2X2 AND2X2_4351 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_10__7_), .Y(w_mem_inst__abc_21203_new_n4543_));
AND2X2 AND2X2_4352 ( .A(round_ctr_rst), .B(\block[199] ), .Y(w_mem_inst__abc_21203_new_n4544_));
AND2X2 AND2X2_4353 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4544_), .Y(w_mem_inst__abc_21203_new_n4545_));
AND2X2 AND2X2_4354 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_9__8_), .Y(w_mem_inst__abc_21203_new_n4548_));
AND2X2 AND2X2_4355 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_10__8_), .Y(w_mem_inst__abc_21203_new_n4549_));
AND2X2 AND2X2_4356 ( .A(round_ctr_rst), .B(\block[200] ), .Y(w_mem_inst__abc_21203_new_n4550_));
AND2X2 AND2X2_4357 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4550_), .Y(w_mem_inst__abc_21203_new_n4551_));
AND2X2 AND2X2_4358 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_9__9_), .Y(w_mem_inst__abc_21203_new_n4554_));
AND2X2 AND2X2_4359 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_10__9_), .Y(w_mem_inst__abc_21203_new_n4555_));
AND2X2 AND2X2_436 ( .A(\digest[39] ), .B(d_reg_7_), .Y(_abc_15497_new_n1616_));
AND2X2 AND2X2_4360 ( .A(round_ctr_rst), .B(\block[201] ), .Y(w_mem_inst__abc_21203_new_n4556_));
AND2X2 AND2X2_4361 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4556_), .Y(w_mem_inst__abc_21203_new_n4557_));
AND2X2 AND2X2_4362 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_9__10_), .Y(w_mem_inst__abc_21203_new_n4560_));
AND2X2 AND2X2_4363 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_10__10_), .Y(w_mem_inst__abc_21203_new_n4561_));
AND2X2 AND2X2_4364 ( .A(round_ctr_rst), .B(\block[202] ), .Y(w_mem_inst__abc_21203_new_n4562_));
AND2X2 AND2X2_4365 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4562_), .Y(w_mem_inst__abc_21203_new_n4563_));
AND2X2 AND2X2_4366 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_9__11_), .Y(w_mem_inst__abc_21203_new_n4566_));
AND2X2 AND2X2_4367 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_10__11_), .Y(w_mem_inst__abc_21203_new_n4567_));
AND2X2 AND2X2_4368 ( .A(round_ctr_rst), .B(\block[203] ), .Y(w_mem_inst__abc_21203_new_n4568_));
AND2X2 AND2X2_4369 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4568_), .Y(w_mem_inst__abc_21203_new_n4569_));
AND2X2 AND2X2_437 ( .A(_abc_15497_new_n1617_), .B(_abc_15497_new_n1615_), .Y(_abc_15497_new_n1618_));
AND2X2 AND2X2_4370 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_9__12_), .Y(w_mem_inst__abc_21203_new_n4572_));
AND2X2 AND2X2_4371 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_10__12_), .Y(w_mem_inst__abc_21203_new_n4573_));
AND2X2 AND2X2_4372 ( .A(round_ctr_rst), .B(\block[204] ), .Y(w_mem_inst__abc_21203_new_n4574_));
AND2X2 AND2X2_4373 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4574_), .Y(w_mem_inst__abc_21203_new_n4575_));
AND2X2 AND2X2_4374 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_9__13_), .Y(w_mem_inst__abc_21203_new_n4578_));
AND2X2 AND2X2_4375 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_10__13_), .Y(w_mem_inst__abc_21203_new_n4579_));
AND2X2 AND2X2_4376 ( .A(round_ctr_rst), .B(\block[205] ), .Y(w_mem_inst__abc_21203_new_n4580_));
AND2X2 AND2X2_4377 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4580_), .Y(w_mem_inst__abc_21203_new_n4581_));
AND2X2 AND2X2_4378 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_9__14_), .Y(w_mem_inst__abc_21203_new_n4584_));
AND2X2 AND2X2_4379 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_10__14_), .Y(w_mem_inst__abc_21203_new_n4585_));
AND2X2 AND2X2_438 ( .A(_abc_15497_new_n1619_), .B(_abc_15497_new_n1618_), .Y(_abc_15497_new_n1621_));
AND2X2 AND2X2_4380 ( .A(round_ctr_rst), .B(\block[206] ), .Y(w_mem_inst__abc_21203_new_n4586_));
AND2X2 AND2X2_4381 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4586_), .Y(w_mem_inst__abc_21203_new_n4587_));
AND2X2 AND2X2_4382 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_9__15_), .Y(w_mem_inst__abc_21203_new_n4590_));
AND2X2 AND2X2_4383 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_10__15_), .Y(w_mem_inst__abc_21203_new_n4591_));
AND2X2 AND2X2_4384 ( .A(round_ctr_rst), .B(\block[207] ), .Y(w_mem_inst__abc_21203_new_n4592_));
AND2X2 AND2X2_4385 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4592_), .Y(w_mem_inst__abc_21203_new_n4593_));
AND2X2 AND2X2_4386 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_9__16_), .Y(w_mem_inst__abc_21203_new_n4596_));
AND2X2 AND2X2_4387 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_10__16_), .Y(w_mem_inst__abc_21203_new_n4597_));
AND2X2 AND2X2_4388 ( .A(round_ctr_rst), .B(\block[208] ), .Y(w_mem_inst__abc_21203_new_n4598_));
AND2X2 AND2X2_4389 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4598_), .Y(w_mem_inst__abc_21203_new_n4599_));
AND2X2 AND2X2_439 ( .A(_abc_15497_new_n1622_), .B(_abc_15497_new_n1620_), .Y(_abc_15497_new_n1623_));
AND2X2 AND2X2_4390 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_9__17_), .Y(w_mem_inst__abc_21203_new_n4602_));
AND2X2 AND2X2_4391 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_10__17_), .Y(w_mem_inst__abc_21203_new_n4603_));
AND2X2 AND2X2_4392 ( .A(round_ctr_rst), .B(\block[209] ), .Y(w_mem_inst__abc_21203_new_n4604_));
AND2X2 AND2X2_4393 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4604_), .Y(w_mem_inst__abc_21203_new_n4605_));
AND2X2 AND2X2_4394 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_9__18_), .Y(w_mem_inst__abc_21203_new_n4608_));
AND2X2 AND2X2_4395 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_10__18_), .Y(w_mem_inst__abc_21203_new_n4609_));
AND2X2 AND2X2_4396 ( .A(round_ctr_rst), .B(\block[210] ), .Y(w_mem_inst__abc_21203_new_n4610_));
AND2X2 AND2X2_4397 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4610_), .Y(w_mem_inst__abc_21203_new_n4611_));
AND2X2 AND2X2_4398 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_9__19_), .Y(w_mem_inst__abc_21203_new_n4614_));
AND2X2 AND2X2_4399 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_10__19_), .Y(w_mem_inst__abc_21203_new_n4615_));
AND2X2 AND2X2_44 ( .A(_abc_15497_new_n766_), .B(_abc_15497_new_n783_), .Y(_abc_15497_new_n784_));
AND2X2 AND2X2_440 ( .A(_abc_15497_new_n1623_), .B(digest_update), .Y(_abc_15497_new_n1624_));
AND2X2 AND2X2_4400 ( .A(round_ctr_rst), .B(\block[211] ), .Y(w_mem_inst__abc_21203_new_n4616_));
AND2X2 AND2X2_4401 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4616_), .Y(w_mem_inst__abc_21203_new_n4617_));
AND2X2 AND2X2_4402 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_9__20_), .Y(w_mem_inst__abc_21203_new_n4620_));
AND2X2 AND2X2_4403 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_10__20_), .Y(w_mem_inst__abc_21203_new_n4621_));
AND2X2 AND2X2_4404 ( .A(round_ctr_rst), .B(\block[212] ), .Y(w_mem_inst__abc_21203_new_n4622_));
AND2X2 AND2X2_4405 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4622_), .Y(w_mem_inst__abc_21203_new_n4623_));
AND2X2 AND2X2_4406 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_9__21_), .Y(w_mem_inst__abc_21203_new_n4626_));
AND2X2 AND2X2_4407 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_10__21_), .Y(w_mem_inst__abc_21203_new_n4627_));
AND2X2 AND2X2_4408 ( .A(round_ctr_rst), .B(\block[213] ), .Y(w_mem_inst__abc_21203_new_n4628_));
AND2X2 AND2X2_4409 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4628_), .Y(w_mem_inst__abc_21203_new_n4629_));
AND2X2 AND2X2_441 ( .A(_abc_15497_new_n701_), .B(\digest[40] ), .Y(_abc_15497_new_n1626_));
AND2X2 AND2X2_4410 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_9__22_), .Y(w_mem_inst__abc_21203_new_n4632_));
AND2X2 AND2X2_4411 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_10__22_), .Y(w_mem_inst__abc_21203_new_n4633_));
AND2X2 AND2X2_4412 ( .A(round_ctr_rst), .B(\block[214] ), .Y(w_mem_inst__abc_21203_new_n4634_));
AND2X2 AND2X2_4413 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4634_), .Y(w_mem_inst__abc_21203_new_n4635_));
AND2X2 AND2X2_4414 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_9__23_), .Y(w_mem_inst__abc_21203_new_n4638_));
AND2X2 AND2X2_4415 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_10__23_), .Y(w_mem_inst__abc_21203_new_n4639_));
AND2X2 AND2X2_4416 ( .A(round_ctr_rst), .B(\block[215] ), .Y(w_mem_inst__abc_21203_new_n4640_));
AND2X2 AND2X2_4417 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4640_), .Y(w_mem_inst__abc_21203_new_n4641_));
AND2X2 AND2X2_4418 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_9__24_), .Y(w_mem_inst__abc_21203_new_n4644_));
AND2X2 AND2X2_4419 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_10__24_), .Y(w_mem_inst__abc_21203_new_n4645_));
AND2X2 AND2X2_442 ( .A(\digest[40] ), .B(d_reg_8_), .Y(_abc_15497_new_n1629_));
AND2X2 AND2X2_4420 ( .A(round_ctr_rst), .B(\block[216] ), .Y(w_mem_inst__abc_21203_new_n4646_));
AND2X2 AND2X2_4421 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4646_), .Y(w_mem_inst__abc_21203_new_n4647_));
AND2X2 AND2X2_4422 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_9__25_), .Y(w_mem_inst__abc_21203_new_n4650_));
AND2X2 AND2X2_4423 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_10__25_), .Y(w_mem_inst__abc_21203_new_n4651_));
AND2X2 AND2X2_4424 ( .A(round_ctr_rst), .B(\block[217] ), .Y(w_mem_inst__abc_21203_new_n4652_));
AND2X2 AND2X2_4425 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4652_), .Y(w_mem_inst__abc_21203_new_n4653_));
AND2X2 AND2X2_4426 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_9__26_), .Y(w_mem_inst__abc_21203_new_n4656_));
AND2X2 AND2X2_4427 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_10__26_), .Y(w_mem_inst__abc_21203_new_n4657_));
AND2X2 AND2X2_4428 ( .A(round_ctr_rst), .B(\block[218] ), .Y(w_mem_inst__abc_21203_new_n4658_));
AND2X2 AND2X2_4429 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4658_), .Y(w_mem_inst__abc_21203_new_n4659_));
AND2X2 AND2X2_443 ( .A(_abc_15497_new_n1630_), .B(_abc_15497_new_n1628_), .Y(_abc_15497_new_n1631_));
AND2X2 AND2X2_4430 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_9__27_), .Y(w_mem_inst__abc_21203_new_n4662_));
AND2X2 AND2X2_4431 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_10__27_), .Y(w_mem_inst__abc_21203_new_n4663_));
AND2X2 AND2X2_4432 ( .A(round_ctr_rst), .B(\block[219] ), .Y(w_mem_inst__abc_21203_new_n4664_));
AND2X2 AND2X2_4433 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4664_), .Y(w_mem_inst__abc_21203_new_n4665_));
AND2X2 AND2X2_4434 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_9__28_), .Y(w_mem_inst__abc_21203_new_n4668_));
AND2X2 AND2X2_4435 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_10__28_), .Y(w_mem_inst__abc_21203_new_n4669_));
AND2X2 AND2X2_4436 ( .A(round_ctr_rst), .B(\block[220] ), .Y(w_mem_inst__abc_21203_new_n4670_));
AND2X2 AND2X2_4437 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4670_), .Y(w_mem_inst__abc_21203_new_n4671_));
AND2X2 AND2X2_4438 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_9__29_), .Y(w_mem_inst__abc_21203_new_n4674_));
AND2X2 AND2X2_4439 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_10__29_), .Y(w_mem_inst__abc_21203_new_n4675_));
AND2X2 AND2X2_444 ( .A(_abc_15497_new_n1627_), .B(_abc_15497_new_n1631_), .Y(_abc_15497_new_n1633_));
AND2X2 AND2X2_4440 ( .A(round_ctr_rst), .B(\block[221] ), .Y(w_mem_inst__abc_21203_new_n4676_));
AND2X2 AND2X2_4441 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4676_), .Y(w_mem_inst__abc_21203_new_n4677_));
AND2X2 AND2X2_4442 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_9__30_), .Y(w_mem_inst__abc_21203_new_n4680_));
AND2X2 AND2X2_4443 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_10__30_), .Y(w_mem_inst__abc_21203_new_n4681_));
AND2X2 AND2X2_4444 ( .A(round_ctr_rst), .B(\block[222] ), .Y(w_mem_inst__abc_21203_new_n4682_));
AND2X2 AND2X2_4445 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4682_), .Y(w_mem_inst__abc_21203_new_n4683_));
AND2X2 AND2X2_4446 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_9__31_), .Y(w_mem_inst__abc_21203_new_n4686_));
AND2X2 AND2X2_4447 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_10__31_), .Y(w_mem_inst__abc_21203_new_n4687_));
AND2X2 AND2X2_4448 ( .A(round_ctr_rst), .B(\block[223] ), .Y(w_mem_inst__abc_21203_new_n4688_));
AND2X2 AND2X2_4449 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4688_), .Y(w_mem_inst__abc_21203_new_n4689_));
AND2X2 AND2X2_445 ( .A(_abc_15497_new_n1634_), .B(_abc_15497_new_n1632_), .Y(_abc_15497_new_n1635_));
AND2X2 AND2X2_4450 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_8__0_), .Y(w_mem_inst__abc_21203_new_n4692_));
AND2X2 AND2X2_4451 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_9__0_), .Y(w_mem_inst__abc_21203_new_n4693_));
AND2X2 AND2X2_4452 ( .A(round_ctr_rst), .B(\block[224] ), .Y(w_mem_inst__abc_21203_new_n4694_));
AND2X2 AND2X2_4453 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4694_), .Y(w_mem_inst__abc_21203_new_n4695_));
AND2X2 AND2X2_4454 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_8__1_), .Y(w_mem_inst__abc_21203_new_n4698_));
AND2X2 AND2X2_4455 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_9__1_), .Y(w_mem_inst__abc_21203_new_n4699_));
AND2X2 AND2X2_4456 ( .A(round_ctr_rst), .B(\block[225] ), .Y(w_mem_inst__abc_21203_new_n4700_));
AND2X2 AND2X2_4457 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4700_), .Y(w_mem_inst__abc_21203_new_n4701_));
AND2X2 AND2X2_4458 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_8__2_), .Y(w_mem_inst__abc_21203_new_n4704_));
AND2X2 AND2X2_4459 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_9__2_), .Y(w_mem_inst__abc_21203_new_n4705_));
AND2X2 AND2X2_446 ( .A(_abc_15497_new_n1635_), .B(digest_update), .Y(_abc_15497_new_n1636_));
AND2X2 AND2X2_4460 ( .A(round_ctr_rst), .B(\block[226] ), .Y(w_mem_inst__abc_21203_new_n4706_));
AND2X2 AND2X2_4461 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4706_), .Y(w_mem_inst__abc_21203_new_n4707_));
AND2X2 AND2X2_4462 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_8__3_), .Y(w_mem_inst__abc_21203_new_n4710_));
AND2X2 AND2X2_4463 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_9__3_), .Y(w_mem_inst__abc_21203_new_n4711_));
AND2X2 AND2X2_4464 ( .A(round_ctr_rst), .B(\block[227] ), .Y(w_mem_inst__abc_21203_new_n4712_));
AND2X2 AND2X2_4465 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4712_), .Y(w_mem_inst__abc_21203_new_n4713_));
AND2X2 AND2X2_4466 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_8__4_), .Y(w_mem_inst__abc_21203_new_n4716_));
AND2X2 AND2X2_4467 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_9__4_), .Y(w_mem_inst__abc_21203_new_n4717_));
AND2X2 AND2X2_4468 ( .A(round_ctr_rst), .B(\block[228] ), .Y(w_mem_inst__abc_21203_new_n4718_));
AND2X2 AND2X2_4469 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4718_), .Y(w_mem_inst__abc_21203_new_n4719_));
AND2X2 AND2X2_447 ( .A(_abc_15497_new_n701_), .B(\digest[41] ), .Y(_abc_15497_new_n1638_));
AND2X2 AND2X2_4470 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_8__5_), .Y(w_mem_inst__abc_21203_new_n4722_));
AND2X2 AND2X2_4471 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_9__5_), .Y(w_mem_inst__abc_21203_new_n4723_));
AND2X2 AND2X2_4472 ( .A(round_ctr_rst), .B(\block[229] ), .Y(w_mem_inst__abc_21203_new_n4724_));
AND2X2 AND2X2_4473 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4724_), .Y(w_mem_inst__abc_21203_new_n4725_));
AND2X2 AND2X2_4474 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_8__6_), .Y(w_mem_inst__abc_21203_new_n4728_));
AND2X2 AND2X2_4475 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_9__6_), .Y(w_mem_inst__abc_21203_new_n4729_));
AND2X2 AND2X2_4476 ( .A(round_ctr_rst), .B(\block[230] ), .Y(w_mem_inst__abc_21203_new_n4730_));
AND2X2 AND2X2_4477 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4730_), .Y(w_mem_inst__abc_21203_new_n4731_));
AND2X2 AND2X2_4478 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_8__7_), .Y(w_mem_inst__abc_21203_new_n4734_));
AND2X2 AND2X2_4479 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_9__7_), .Y(w_mem_inst__abc_21203_new_n4735_));
AND2X2 AND2X2_448 ( .A(\digest[41] ), .B(d_reg_9_), .Y(_abc_15497_new_n1640_));
AND2X2 AND2X2_4480 ( .A(round_ctr_rst), .B(\block[231] ), .Y(w_mem_inst__abc_21203_new_n4736_));
AND2X2 AND2X2_4481 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4736_), .Y(w_mem_inst__abc_21203_new_n4737_));
AND2X2 AND2X2_4482 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_8__8_), .Y(w_mem_inst__abc_21203_new_n4740_));
AND2X2 AND2X2_4483 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_9__8_), .Y(w_mem_inst__abc_21203_new_n4741_));
AND2X2 AND2X2_4484 ( .A(round_ctr_rst), .B(\block[232] ), .Y(w_mem_inst__abc_21203_new_n4742_));
AND2X2 AND2X2_4485 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4742_), .Y(w_mem_inst__abc_21203_new_n4743_));
AND2X2 AND2X2_4486 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_8__9_), .Y(w_mem_inst__abc_21203_new_n4746_));
AND2X2 AND2X2_4487 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_9__9_), .Y(w_mem_inst__abc_21203_new_n4747_));
AND2X2 AND2X2_4488 ( .A(round_ctr_rst), .B(\block[233] ), .Y(w_mem_inst__abc_21203_new_n4748_));
AND2X2 AND2X2_4489 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4748_), .Y(w_mem_inst__abc_21203_new_n4749_));
AND2X2 AND2X2_449 ( .A(_abc_15497_new_n1641_), .B(_abc_15497_new_n1639_), .Y(_abc_15497_new_n1642_));
AND2X2 AND2X2_4490 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_8__10_), .Y(w_mem_inst__abc_21203_new_n4752_));
AND2X2 AND2X2_4491 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_9__10_), .Y(w_mem_inst__abc_21203_new_n4753_));
AND2X2 AND2X2_4492 ( .A(round_ctr_rst), .B(\block[234] ), .Y(w_mem_inst__abc_21203_new_n4754_));
AND2X2 AND2X2_4493 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4754_), .Y(w_mem_inst__abc_21203_new_n4755_));
AND2X2 AND2X2_4494 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_8__11_), .Y(w_mem_inst__abc_21203_new_n4758_));
AND2X2 AND2X2_4495 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_9__11_), .Y(w_mem_inst__abc_21203_new_n4759_));
AND2X2 AND2X2_4496 ( .A(round_ctr_rst), .B(\block[235] ), .Y(w_mem_inst__abc_21203_new_n4760_));
AND2X2 AND2X2_4497 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4760_), .Y(w_mem_inst__abc_21203_new_n4761_));
AND2X2 AND2X2_4498 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_8__12_), .Y(w_mem_inst__abc_21203_new_n4764_));
AND2X2 AND2X2_4499 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_9__12_), .Y(w_mem_inst__abc_21203_new_n4765_));
AND2X2 AND2X2_45 ( .A(c_reg_11_), .B(\digest[75] ), .Y(_abc_15497_new_n785_));
AND2X2 AND2X2_450 ( .A(_abc_15497_new_n1631_), .B(_abc_15497_new_n1642_), .Y(_abc_15497_new_n1645_));
AND2X2 AND2X2_4500 ( .A(round_ctr_rst), .B(\block[236] ), .Y(w_mem_inst__abc_21203_new_n4766_));
AND2X2 AND2X2_4501 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4766_), .Y(w_mem_inst__abc_21203_new_n4767_));
AND2X2 AND2X2_4502 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_8__13_), .Y(w_mem_inst__abc_21203_new_n4770_));
AND2X2 AND2X2_4503 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_9__13_), .Y(w_mem_inst__abc_21203_new_n4771_));
AND2X2 AND2X2_4504 ( .A(round_ctr_rst), .B(\block[237] ), .Y(w_mem_inst__abc_21203_new_n4772_));
AND2X2 AND2X2_4505 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4772_), .Y(w_mem_inst__abc_21203_new_n4773_));
AND2X2 AND2X2_4506 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_8__14_), .Y(w_mem_inst__abc_21203_new_n4776_));
AND2X2 AND2X2_4507 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_9__14_), .Y(w_mem_inst__abc_21203_new_n4777_));
AND2X2 AND2X2_4508 ( .A(round_ctr_rst), .B(\block[238] ), .Y(w_mem_inst__abc_21203_new_n4778_));
AND2X2 AND2X2_4509 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4778_), .Y(w_mem_inst__abc_21203_new_n4779_));
AND2X2 AND2X2_451 ( .A(_abc_15497_new_n1627_), .B(_abc_15497_new_n1645_), .Y(_abc_15497_new_n1646_));
AND2X2 AND2X2_4510 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_8__15_), .Y(w_mem_inst__abc_21203_new_n4782_));
AND2X2 AND2X2_4511 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_9__15_), .Y(w_mem_inst__abc_21203_new_n4783_));
AND2X2 AND2X2_4512 ( .A(round_ctr_rst), .B(\block[239] ), .Y(w_mem_inst__abc_21203_new_n4784_));
AND2X2 AND2X2_4513 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4784_), .Y(w_mem_inst__abc_21203_new_n4785_));
AND2X2 AND2X2_4514 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_8__16_), .Y(w_mem_inst__abc_21203_new_n4788_));
AND2X2 AND2X2_4515 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_9__16_), .Y(w_mem_inst__abc_21203_new_n4789_));
AND2X2 AND2X2_4516 ( .A(round_ctr_rst), .B(\block[240] ), .Y(w_mem_inst__abc_21203_new_n4790_));
AND2X2 AND2X2_4517 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4790_), .Y(w_mem_inst__abc_21203_new_n4791_));
AND2X2 AND2X2_4518 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_8__17_), .Y(w_mem_inst__abc_21203_new_n4794_));
AND2X2 AND2X2_4519 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_9__17_), .Y(w_mem_inst__abc_21203_new_n4795_));
AND2X2 AND2X2_452 ( .A(_abc_15497_new_n1642_), .B(_abc_15497_new_n1629_), .Y(_abc_15497_new_n1648_));
AND2X2 AND2X2_4520 ( .A(round_ctr_rst), .B(\block[241] ), .Y(w_mem_inst__abc_21203_new_n4796_));
AND2X2 AND2X2_4521 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4796_), .Y(w_mem_inst__abc_21203_new_n4797_));
AND2X2 AND2X2_4522 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_8__18_), .Y(w_mem_inst__abc_21203_new_n4800_));
AND2X2 AND2X2_4523 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_9__18_), .Y(w_mem_inst__abc_21203_new_n4801_));
AND2X2 AND2X2_4524 ( .A(round_ctr_rst), .B(\block[242] ), .Y(w_mem_inst__abc_21203_new_n4802_));
AND2X2 AND2X2_4525 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4802_), .Y(w_mem_inst__abc_21203_new_n4803_));
AND2X2 AND2X2_4526 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_8__19_), .Y(w_mem_inst__abc_21203_new_n4806_));
AND2X2 AND2X2_4527 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_9__19_), .Y(w_mem_inst__abc_21203_new_n4807_));
AND2X2 AND2X2_4528 ( .A(round_ctr_rst), .B(\block[243] ), .Y(w_mem_inst__abc_21203_new_n4808_));
AND2X2 AND2X2_4529 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4808_), .Y(w_mem_inst__abc_21203_new_n4809_));
AND2X2 AND2X2_453 ( .A(_abc_15497_new_n1649_), .B(digest_update), .Y(_abc_15497_new_n1650_));
AND2X2 AND2X2_4530 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_8__20_), .Y(w_mem_inst__abc_21203_new_n4812_));
AND2X2 AND2X2_4531 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_9__20_), .Y(w_mem_inst__abc_21203_new_n4813_));
AND2X2 AND2X2_4532 ( .A(round_ctr_rst), .B(\block[244] ), .Y(w_mem_inst__abc_21203_new_n4814_));
AND2X2 AND2X2_4533 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4814_), .Y(w_mem_inst__abc_21203_new_n4815_));
AND2X2 AND2X2_4534 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_8__21_), .Y(w_mem_inst__abc_21203_new_n4818_));
AND2X2 AND2X2_4535 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_9__21_), .Y(w_mem_inst__abc_21203_new_n4819_));
AND2X2 AND2X2_4536 ( .A(round_ctr_rst), .B(\block[245] ), .Y(w_mem_inst__abc_21203_new_n4820_));
AND2X2 AND2X2_4537 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4820_), .Y(w_mem_inst__abc_21203_new_n4821_));
AND2X2 AND2X2_4538 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_8__22_), .Y(w_mem_inst__abc_21203_new_n4824_));
AND2X2 AND2X2_4539 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_9__22_), .Y(w_mem_inst__abc_21203_new_n4825_));
AND2X2 AND2X2_454 ( .A(_abc_15497_new_n1647_), .B(_abc_15497_new_n1650_), .Y(_abc_15497_new_n1651_));
AND2X2 AND2X2_4540 ( .A(round_ctr_rst), .B(\block[246] ), .Y(w_mem_inst__abc_21203_new_n4826_));
AND2X2 AND2X2_4541 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4826_), .Y(w_mem_inst__abc_21203_new_n4827_));
AND2X2 AND2X2_4542 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_8__23_), .Y(w_mem_inst__abc_21203_new_n4830_));
AND2X2 AND2X2_4543 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_9__23_), .Y(w_mem_inst__abc_21203_new_n4831_));
AND2X2 AND2X2_4544 ( .A(round_ctr_rst), .B(\block[247] ), .Y(w_mem_inst__abc_21203_new_n4832_));
AND2X2 AND2X2_4545 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4832_), .Y(w_mem_inst__abc_21203_new_n4833_));
AND2X2 AND2X2_4546 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_8__24_), .Y(w_mem_inst__abc_21203_new_n4836_));
AND2X2 AND2X2_4547 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_9__24_), .Y(w_mem_inst__abc_21203_new_n4837_));
AND2X2 AND2X2_4548 ( .A(round_ctr_rst), .B(\block[248] ), .Y(w_mem_inst__abc_21203_new_n4838_));
AND2X2 AND2X2_4549 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4838_), .Y(w_mem_inst__abc_21203_new_n4839_));
AND2X2 AND2X2_455 ( .A(_abc_15497_new_n1651_), .B(_abc_15497_new_n1644_), .Y(_abc_15497_new_n1652_));
AND2X2 AND2X2_4550 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_8__25_), .Y(w_mem_inst__abc_21203_new_n4842_));
AND2X2 AND2X2_4551 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_9__25_), .Y(w_mem_inst__abc_21203_new_n4843_));
AND2X2 AND2X2_4552 ( .A(round_ctr_rst), .B(\block[249] ), .Y(w_mem_inst__abc_21203_new_n4844_));
AND2X2 AND2X2_4553 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4844_), .Y(w_mem_inst__abc_21203_new_n4845_));
AND2X2 AND2X2_4554 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_8__26_), .Y(w_mem_inst__abc_21203_new_n4848_));
AND2X2 AND2X2_4555 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_9__26_), .Y(w_mem_inst__abc_21203_new_n4849_));
AND2X2 AND2X2_4556 ( .A(round_ctr_rst), .B(\block[250] ), .Y(w_mem_inst__abc_21203_new_n4850_));
AND2X2 AND2X2_4557 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4850_), .Y(w_mem_inst__abc_21203_new_n4851_));
AND2X2 AND2X2_4558 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_8__27_), .Y(w_mem_inst__abc_21203_new_n4854_));
AND2X2 AND2X2_4559 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_9__27_), .Y(w_mem_inst__abc_21203_new_n4855_));
AND2X2 AND2X2_456 ( .A(_abc_15497_new_n1649_), .B(_abc_15497_new_n1641_), .Y(_abc_15497_new_n1654_));
AND2X2 AND2X2_4560 ( .A(round_ctr_rst), .B(\block[251] ), .Y(w_mem_inst__abc_21203_new_n4856_));
AND2X2 AND2X2_4561 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4856_), .Y(w_mem_inst__abc_21203_new_n4857_));
AND2X2 AND2X2_4562 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_8__28_), .Y(w_mem_inst__abc_21203_new_n4860_));
AND2X2 AND2X2_4563 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_9__28_), .Y(w_mem_inst__abc_21203_new_n4861_));
AND2X2 AND2X2_4564 ( .A(round_ctr_rst), .B(\block[252] ), .Y(w_mem_inst__abc_21203_new_n4862_));
AND2X2 AND2X2_4565 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4862_), .Y(w_mem_inst__abc_21203_new_n4863_));
AND2X2 AND2X2_4566 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_8__29_), .Y(w_mem_inst__abc_21203_new_n4866_));
AND2X2 AND2X2_4567 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_9__29_), .Y(w_mem_inst__abc_21203_new_n4867_));
AND2X2 AND2X2_4568 ( .A(round_ctr_rst), .B(\block[253] ), .Y(w_mem_inst__abc_21203_new_n4868_));
AND2X2 AND2X2_4569 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4868_), .Y(w_mem_inst__abc_21203_new_n4869_));
AND2X2 AND2X2_457 ( .A(_abc_15497_new_n1647_), .B(_abc_15497_new_n1654_), .Y(_abc_15497_new_n1655_));
AND2X2 AND2X2_4570 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_8__30_), .Y(w_mem_inst__abc_21203_new_n4872_));
AND2X2 AND2X2_4571 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_9__30_), .Y(w_mem_inst__abc_21203_new_n4873_));
AND2X2 AND2X2_4572 ( .A(round_ctr_rst), .B(\block[254] ), .Y(w_mem_inst__abc_21203_new_n4874_));
AND2X2 AND2X2_4573 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4874_), .Y(w_mem_inst__abc_21203_new_n4875_));
AND2X2 AND2X2_4574 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_8__31_), .Y(w_mem_inst__abc_21203_new_n4878_));
AND2X2 AND2X2_4575 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_9__31_), .Y(w_mem_inst__abc_21203_new_n4879_));
AND2X2 AND2X2_4576 ( .A(round_ctr_rst), .B(\block[255] ), .Y(w_mem_inst__abc_21203_new_n4880_));
AND2X2 AND2X2_4577 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4880_), .Y(w_mem_inst__abc_21203_new_n4881_));
AND2X2 AND2X2_4578 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_4__0_), .Y(w_mem_inst__abc_21203_new_n4884_));
AND2X2 AND2X2_4579 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_5__0_), .Y(w_mem_inst__abc_21203_new_n4885_));
AND2X2 AND2X2_458 ( .A(\digest[42] ), .B(d_reg_10_), .Y(_abc_15497_new_n1658_));
AND2X2 AND2X2_4580 ( .A(round_ctr_rst), .B(\block[352] ), .Y(w_mem_inst__abc_21203_new_n4886_));
AND2X2 AND2X2_4581 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4886_), .Y(w_mem_inst__abc_21203_new_n4887_));
AND2X2 AND2X2_4582 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_4__1_), .Y(w_mem_inst__abc_21203_new_n4890_));
AND2X2 AND2X2_4583 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_5__1_), .Y(w_mem_inst__abc_21203_new_n4891_));
AND2X2 AND2X2_4584 ( .A(round_ctr_rst), .B(\block[353] ), .Y(w_mem_inst__abc_21203_new_n4892_));
AND2X2 AND2X2_4585 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4892_), .Y(w_mem_inst__abc_21203_new_n4893_));
AND2X2 AND2X2_4586 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_4__2_), .Y(w_mem_inst__abc_21203_new_n4896_));
AND2X2 AND2X2_4587 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_5__2_), .Y(w_mem_inst__abc_21203_new_n4897_));
AND2X2 AND2X2_4588 ( .A(round_ctr_rst), .B(\block[354] ), .Y(w_mem_inst__abc_21203_new_n4898_));
AND2X2 AND2X2_4589 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4898_), .Y(w_mem_inst__abc_21203_new_n4899_));
AND2X2 AND2X2_459 ( .A(_abc_15497_new_n1659_), .B(_abc_15497_new_n1657_), .Y(_abc_15497_new_n1660_));
AND2X2 AND2X2_4590 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_4__3_), .Y(w_mem_inst__abc_21203_new_n4902_));
AND2X2 AND2X2_4591 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_5__3_), .Y(w_mem_inst__abc_21203_new_n4903_));
AND2X2 AND2X2_4592 ( .A(round_ctr_rst), .B(\block[355] ), .Y(w_mem_inst__abc_21203_new_n4904_));
AND2X2 AND2X2_4593 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4904_), .Y(w_mem_inst__abc_21203_new_n4905_));
AND2X2 AND2X2_4594 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_4__4_), .Y(w_mem_inst__abc_21203_new_n4908_));
AND2X2 AND2X2_4595 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_5__4_), .Y(w_mem_inst__abc_21203_new_n4909_));
AND2X2 AND2X2_4596 ( .A(round_ctr_rst), .B(\block[356] ), .Y(w_mem_inst__abc_21203_new_n4910_));
AND2X2 AND2X2_4597 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4910_), .Y(w_mem_inst__abc_21203_new_n4911_));
AND2X2 AND2X2_4598 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_4__5_), .Y(w_mem_inst__abc_21203_new_n4914_));
AND2X2 AND2X2_4599 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_5__5_), .Y(w_mem_inst__abc_21203_new_n4915_));
AND2X2 AND2X2_46 ( .A(c_reg_10_), .B(\digest[74] ), .Y(_abc_15497_new_n787_));
AND2X2 AND2X2_460 ( .A(_abc_15497_new_n1656_), .B(_abc_15497_new_n1660_), .Y(_abc_15497_new_n1662_));
AND2X2 AND2X2_4600 ( .A(round_ctr_rst), .B(\block[357] ), .Y(w_mem_inst__abc_21203_new_n4916_));
AND2X2 AND2X2_4601 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4916_), .Y(w_mem_inst__abc_21203_new_n4917_));
AND2X2 AND2X2_4602 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_4__6_), .Y(w_mem_inst__abc_21203_new_n4920_));
AND2X2 AND2X2_4603 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_5__6_), .Y(w_mem_inst__abc_21203_new_n4921_));
AND2X2 AND2X2_4604 ( .A(round_ctr_rst), .B(\block[358] ), .Y(w_mem_inst__abc_21203_new_n4922_));
AND2X2 AND2X2_4605 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4922_), .Y(w_mem_inst__abc_21203_new_n4923_));
AND2X2 AND2X2_4606 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_4__7_), .Y(w_mem_inst__abc_21203_new_n4926_));
AND2X2 AND2X2_4607 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_5__7_), .Y(w_mem_inst__abc_21203_new_n4927_));
AND2X2 AND2X2_4608 ( .A(round_ctr_rst), .B(\block[359] ), .Y(w_mem_inst__abc_21203_new_n4928_));
AND2X2 AND2X2_4609 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4928_), .Y(w_mem_inst__abc_21203_new_n4929_));
AND2X2 AND2X2_461 ( .A(_abc_15497_new_n1663_), .B(_abc_15497_new_n1661_), .Y(_abc_15497_new_n1664_));
AND2X2 AND2X2_4610 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_4__8_), .Y(w_mem_inst__abc_21203_new_n4932_));
AND2X2 AND2X2_4611 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_5__8_), .Y(w_mem_inst__abc_21203_new_n4933_));
AND2X2 AND2X2_4612 ( .A(round_ctr_rst), .B(\block[360] ), .Y(w_mem_inst__abc_21203_new_n4934_));
AND2X2 AND2X2_4613 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4934_), .Y(w_mem_inst__abc_21203_new_n4935_));
AND2X2 AND2X2_4614 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_4__9_), .Y(w_mem_inst__abc_21203_new_n4938_));
AND2X2 AND2X2_4615 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_5__9_), .Y(w_mem_inst__abc_21203_new_n4939_));
AND2X2 AND2X2_4616 ( .A(round_ctr_rst), .B(\block[361] ), .Y(w_mem_inst__abc_21203_new_n4940_));
AND2X2 AND2X2_4617 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4940_), .Y(w_mem_inst__abc_21203_new_n4941_));
AND2X2 AND2X2_4618 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_4__10_), .Y(w_mem_inst__abc_21203_new_n4944_));
AND2X2 AND2X2_4619 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_5__10_), .Y(w_mem_inst__abc_21203_new_n4945_));
AND2X2 AND2X2_462 ( .A(_abc_15497_new_n1664_), .B(digest_update), .Y(_abc_15497_new_n1665_));
AND2X2 AND2X2_4620 ( .A(round_ctr_rst), .B(\block[362] ), .Y(w_mem_inst__abc_21203_new_n4946_));
AND2X2 AND2X2_4621 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4946_), .Y(w_mem_inst__abc_21203_new_n4947_));
AND2X2 AND2X2_4622 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_4__11_), .Y(w_mem_inst__abc_21203_new_n4950_));
AND2X2 AND2X2_4623 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_5__11_), .Y(w_mem_inst__abc_21203_new_n4951_));
AND2X2 AND2X2_4624 ( .A(round_ctr_rst), .B(\block[363] ), .Y(w_mem_inst__abc_21203_new_n4952_));
AND2X2 AND2X2_4625 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4952_), .Y(w_mem_inst__abc_21203_new_n4953_));
AND2X2 AND2X2_4626 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_4__12_), .Y(w_mem_inst__abc_21203_new_n4956_));
AND2X2 AND2X2_4627 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_5__12_), .Y(w_mem_inst__abc_21203_new_n4957_));
AND2X2 AND2X2_4628 ( .A(round_ctr_rst), .B(\block[364] ), .Y(w_mem_inst__abc_21203_new_n4958_));
AND2X2 AND2X2_4629 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4958_), .Y(w_mem_inst__abc_21203_new_n4959_));
AND2X2 AND2X2_463 ( .A(_abc_15497_new_n1666_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n1667_));
AND2X2 AND2X2_4630 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_4__13_), .Y(w_mem_inst__abc_21203_new_n4962_));
AND2X2 AND2X2_4631 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_5__13_), .Y(w_mem_inst__abc_21203_new_n4963_));
AND2X2 AND2X2_4632 ( .A(round_ctr_rst), .B(\block[365] ), .Y(w_mem_inst__abc_21203_new_n4964_));
AND2X2 AND2X2_4633 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4964_), .Y(w_mem_inst__abc_21203_new_n4965_));
AND2X2 AND2X2_4634 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_4__14_), .Y(w_mem_inst__abc_21203_new_n4968_));
AND2X2 AND2X2_4635 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_5__14_), .Y(w_mem_inst__abc_21203_new_n4969_));
AND2X2 AND2X2_4636 ( .A(round_ctr_rst), .B(\block[366] ), .Y(w_mem_inst__abc_21203_new_n4970_));
AND2X2 AND2X2_4637 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4970_), .Y(w_mem_inst__abc_21203_new_n4971_));
AND2X2 AND2X2_4638 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_4__15_), .Y(w_mem_inst__abc_21203_new_n4974_));
AND2X2 AND2X2_4639 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_5__15_), .Y(w_mem_inst__abc_21203_new_n4975_));
AND2X2 AND2X2_464 ( .A(_abc_15497_new_n701_), .B(\digest[43] ), .Y(_abc_15497_new_n1669_));
AND2X2 AND2X2_4640 ( .A(round_ctr_rst), .B(\block[367] ), .Y(w_mem_inst__abc_21203_new_n4976_));
AND2X2 AND2X2_4641 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4976_), .Y(w_mem_inst__abc_21203_new_n4977_));
AND2X2 AND2X2_4642 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_4__16_), .Y(w_mem_inst__abc_21203_new_n4980_));
AND2X2 AND2X2_4643 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_5__16_), .Y(w_mem_inst__abc_21203_new_n4981_));
AND2X2 AND2X2_4644 ( .A(round_ctr_rst), .B(\block[368] ), .Y(w_mem_inst__abc_21203_new_n4982_));
AND2X2 AND2X2_4645 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4982_), .Y(w_mem_inst__abc_21203_new_n4983_));
AND2X2 AND2X2_4646 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_4__17_), .Y(w_mem_inst__abc_21203_new_n4986_));
AND2X2 AND2X2_4647 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_5__17_), .Y(w_mem_inst__abc_21203_new_n4987_));
AND2X2 AND2X2_4648 ( .A(round_ctr_rst), .B(\block[369] ), .Y(w_mem_inst__abc_21203_new_n4988_));
AND2X2 AND2X2_4649 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4988_), .Y(w_mem_inst__abc_21203_new_n4989_));
AND2X2 AND2X2_465 ( .A(_abc_15497_new_n1663_), .B(_abc_15497_new_n1659_), .Y(_abc_15497_new_n1670_));
AND2X2 AND2X2_4650 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_4__18_), .Y(w_mem_inst__abc_21203_new_n4992_));
AND2X2 AND2X2_4651 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_5__18_), .Y(w_mem_inst__abc_21203_new_n4993_));
AND2X2 AND2X2_4652 ( .A(round_ctr_rst), .B(\block[370] ), .Y(w_mem_inst__abc_21203_new_n4994_));
AND2X2 AND2X2_4653 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n4994_), .Y(w_mem_inst__abc_21203_new_n4995_));
AND2X2 AND2X2_4654 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_4__19_), .Y(w_mem_inst__abc_21203_new_n4998_));
AND2X2 AND2X2_4655 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_5__19_), .Y(w_mem_inst__abc_21203_new_n4999_));
AND2X2 AND2X2_4656 ( .A(round_ctr_rst), .B(\block[371] ), .Y(w_mem_inst__abc_21203_new_n5000_));
AND2X2 AND2X2_4657 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5000_), .Y(w_mem_inst__abc_21203_new_n5001_));
AND2X2 AND2X2_4658 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_4__20_), .Y(w_mem_inst__abc_21203_new_n5004_));
AND2X2 AND2X2_4659 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_5__20_), .Y(w_mem_inst__abc_21203_new_n5005_));
AND2X2 AND2X2_466 ( .A(\digest[43] ), .B(d_reg_11_), .Y(_abc_15497_new_n1673_));
AND2X2 AND2X2_4660 ( .A(round_ctr_rst), .B(\block[372] ), .Y(w_mem_inst__abc_21203_new_n5006_));
AND2X2 AND2X2_4661 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5006_), .Y(w_mem_inst__abc_21203_new_n5007_));
AND2X2 AND2X2_4662 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_4__21_), .Y(w_mem_inst__abc_21203_new_n5010_));
AND2X2 AND2X2_4663 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_5__21_), .Y(w_mem_inst__abc_21203_new_n5011_));
AND2X2 AND2X2_4664 ( .A(round_ctr_rst), .B(\block[373] ), .Y(w_mem_inst__abc_21203_new_n5012_));
AND2X2 AND2X2_4665 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5012_), .Y(w_mem_inst__abc_21203_new_n5013_));
AND2X2 AND2X2_4666 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_4__22_), .Y(w_mem_inst__abc_21203_new_n5016_));
AND2X2 AND2X2_4667 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_5__22_), .Y(w_mem_inst__abc_21203_new_n5017_));
AND2X2 AND2X2_4668 ( .A(round_ctr_rst), .B(\block[374] ), .Y(w_mem_inst__abc_21203_new_n5018_));
AND2X2 AND2X2_4669 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5018_), .Y(w_mem_inst__abc_21203_new_n5019_));
AND2X2 AND2X2_467 ( .A(_abc_15497_new_n1674_), .B(_abc_15497_new_n1672_), .Y(_abc_15497_new_n1675_));
AND2X2 AND2X2_4670 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_4__23_), .Y(w_mem_inst__abc_21203_new_n5022_));
AND2X2 AND2X2_4671 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_5__23_), .Y(w_mem_inst__abc_21203_new_n5023_));
AND2X2 AND2X2_4672 ( .A(round_ctr_rst), .B(\block[375] ), .Y(w_mem_inst__abc_21203_new_n5024_));
AND2X2 AND2X2_4673 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5024_), .Y(w_mem_inst__abc_21203_new_n5025_));
AND2X2 AND2X2_4674 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_4__24_), .Y(w_mem_inst__abc_21203_new_n5028_));
AND2X2 AND2X2_4675 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_5__24_), .Y(w_mem_inst__abc_21203_new_n5029_));
AND2X2 AND2X2_4676 ( .A(round_ctr_rst), .B(\block[376] ), .Y(w_mem_inst__abc_21203_new_n5030_));
AND2X2 AND2X2_4677 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5030_), .Y(w_mem_inst__abc_21203_new_n5031_));
AND2X2 AND2X2_4678 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_4__25_), .Y(w_mem_inst__abc_21203_new_n5034_));
AND2X2 AND2X2_4679 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_5__25_), .Y(w_mem_inst__abc_21203_new_n5035_));
AND2X2 AND2X2_468 ( .A(_abc_15497_new_n1678_), .B(digest_update), .Y(_abc_15497_new_n1679_));
AND2X2 AND2X2_4680 ( .A(round_ctr_rst), .B(\block[377] ), .Y(w_mem_inst__abc_21203_new_n5036_));
AND2X2 AND2X2_4681 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5036_), .Y(w_mem_inst__abc_21203_new_n5037_));
AND2X2 AND2X2_4682 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_4__26_), .Y(w_mem_inst__abc_21203_new_n5040_));
AND2X2 AND2X2_4683 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_5__26_), .Y(w_mem_inst__abc_21203_new_n5041_));
AND2X2 AND2X2_4684 ( .A(round_ctr_rst), .B(\block[378] ), .Y(w_mem_inst__abc_21203_new_n5042_));
AND2X2 AND2X2_4685 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5042_), .Y(w_mem_inst__abc_21203_new_n5043_));
AND2X2 AND2X2_4686 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_4__27_), .Y(w_mem_inst__abc_21203_new_n5046_));
AND2X2 AND2X2_4687 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_5__27_), .Y(w_mem_inst__abc_21203_new_n5047_));
AND2X2 AND2X2_4688 ( .A(round_ctr_rst), .B(\block[379] ), .Y(w_mem_inst__abc_21203_new_n5048_));
AND2X2 AND2X2_4689 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5048_), .Y(w_mem_inst__abc_21203_new_n5049_));
AND2X2 AND2X2_469 ( .A(_abc_15497_new_n1679_), .B(_abc_15497_new_n1676_), .Y(_abc_15497_new_n1680_));
AND2X2 AND2X2_4690 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_4__28_), .Y(w_mem_inst__abc_21203_new_n5052_));
AND2X2 AND2X2_4691 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_5__28_), .Y(w_mem_inst__abc_21203_new_n5053_));
AND2X2 AND2X2_4692 ( .A(round_ctr_rst), .B(\block[380] ), .Y(w_mem_inst__abc_21203_new_n5054_));
AND2X2 AND2X2_4693 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5054_), .Y(w_mem_inst__abc_21203_new_n5055_));
AND2X2 AND2X2_4694 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_4__29_), .Y(w_mem_inst__abc_21203_new_n5058_));
AND2X2 AND2X2_4695 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_5__29_), .Y(w_mem_inst__abc_21203_new_n5059_));
AND2X2 AND2X2_4696 ( .A(round_ctr_rst), .B(\block[381] ), .Y(w_mem_inst__abc_21203_new_n5060_));
AND2X2 AND2X2_4697 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5060_), .Y(w_mem_inst__abc_21203_new_n5061_));
AND2X2 AND2X2_4698 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_4__30_), .Y(w_mem_inst__abc_21203_new_n5064_));
AND2X2 AND2X2_4699 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_5__30_), .Y(w_mem_inst__abc_21203_new_n5065_));
AND2X2 AND2X2_47 ( .A(_abc_15497_new_n786_), .B(_abc_15497_new_n787_), .Y(_abc_15497_new_n788_));
AND2X2 AND2X2_470 ( .A(_abc_15497_new_n1660_), .B(_abc_15497_new_n1675_), .Y(_abc_15497_new_n1682_));
AND2X2 AND2X2_4700 ( .A(round_ctr_rst), .B(\block[382] ), .Y(w_mem_inst__abc_21203_new_n5066_));
AND2X2 AND2X2_4701 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5066_), .Y(w_mem_inst__abc_21203_new_n5067_));
AND2X2 AND2X2_4702 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_4__31_), .Y(w_mem_inst__abc_21203_new_n5070_));
AND2X2 AND2X2_4703 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_5__31_), .Y(w_mem_inst__abc_21203_new_n5071_));
AND2X2 AND2X2_4704 ( .A(round_ctr_rst), .B(\block[383] ), .Y(w_mem_inst__abc_21203_new_n5072_));
AND2X2 AND2X2_4705 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5072_), .Y(w_mem_inst__abc_21203_new_n5073_));
AND2X2 AND2X2_4706 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_6__0_), .Y(w_mem_inst__abc_21203_new_n5076_));
AND2X2 AND2X2_4707 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_7__0_), .Y(w_mem_inst__abc_21203_new_n5077_));
AND2X2 AND2X2_4708 ( .A(round_ctr_rst), .B(\block[288] ), .Y(w_mem_inst__abc_21203_new_n5078_));
AND2X2 AND2X2_4709 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5078_), .Y(w_mem_inst__abc_21203_new_n5079_));
AND2X2 AND2X2_471 ( .A(_abc_15497_new_n1645_), .B(_abc_15497_new_n1682_), .Y(_abc_15497_new_n1683_));
AND2X2 AND2X2_4710 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_6__1_), .Y(w_mem_inst__abc_21203_new_n5082_));
AND2X2 AND2X2_4711 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_7__1_), .Y(w_mem_inst__abc_21203_new_n5083_));
AND2X2 AND2X2_4712 ( .A(round_ctr_rst), .B(\block[289] ), .Y(w_mem_inst__abc_21203_new_n5084_));
AND2X2 AND2X2_4713 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5084_), .Y(w_mem_inst__abc_21203_new_n5085_));
AND2X2 AND2X2_4714 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_6__2_), .Y(w_mem_inst__abc_21203_new_n5088_));
AND2X2 AND2X2_4715 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_7__2_), .Y(w_mem_inst__abc_21203_new_n5089_));
AND2X2 AND2X2_4716 ( .A(round_ctr_rst), .B(\block[290] ), .Y(w_mem_inst__abc_21203_new_n5090_));
AND2X2 AND2X2_4717 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5090_), .Y(w_mem_inst__abc_21203_new_n5091_));
AND2X2 AND2X2_4718 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_6__3_), .Y(w_mem_inst__abc_21203_new_n5094_));
AND2X2 AND2X2_4719 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_7__3_), .Y(w_mem_inst__abc_21203_new_n5095_));
AND2X2 AND2X2_472 ( .A(_abc_15497_new_n1627_), .B(_abc_15497_new_n1683_), .Y(_abc_15497_new_n1684_));
AND2X2 AND2X2_4720 ( .A(round_ctr_rst), .B(\block[291] ), .Y(w_mem_inst__abc_21203_new_n5096_));
AND2X2 AND2X2_4721 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5096_), .Y(w_mem_inst__abc_21203_new_n5097_));
AND2X2 AND2X2_4722 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_6__4_), .Y(w_mem_inst__abc_21203_new_n5100_));
AND2X2 AND2X2_4723 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_7__4_), .Y(w_mem_inst__abc_21203_new_n5101_));
AND2X2 AND2X2_4724 ( .A(round_ctr_rst), .B(\block[292] ), .Y(w_mem_inst__abc_21203_new_n5102_));
AND2X2 AND2X2_4725 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5102_), .Y(w_mem_inst__abc_21203_new_n5103_));
AND2X2 AND2X2_4726 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_6__5_), .Y(w_mem_inst__abc_21203_new_n5106_));
AND2X2 AND2X2_4727 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_7__5_), .Y(w_mem_inst__abc_21203_new_n5107_));
AND2X2 AND2X2_4728 ( .A(round_ctr_rst), .B(\block[293] ), .Y(w_mem_inst__abc_21203_new_n5108_));
AND2X2 AND2X2_4729 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5108_), .Y(w_mem_inst__abc_21203_new_n5109_));
AND2X2 AND2X2_473 ( .A(_abc_15497_new_n1685_), .B(_abc_15497_new_n1682_), .Y(_abc_15497_new_n1686_));
AND2X2 AND2X2_4730 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_6__6_), .Y(w_mem_inst__abc_21203_new_n5112_));
AND2X2 AND2X2_4731 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_7__6_), .Y(w_mem_inst__abc_21203_new_n5113_));
AND2X2 AND2X2_4732 ( .A(round_ctr_rst), .B(\block[294] ), .Y(w_mem_inst__abc_21203_new_n5114_));
AND2X2 AND2X2_4733 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5114_), .Y(w_mem_inst__abc_21203_new_n5115_));
AND2X2 AND2X2_4734 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_6__7_), .Y(w_mem_inst__abc_21203_new_n5118_));
AND2X2 AND2X2_4735 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_7__7_), .Y(w_mem_inst__abc_21203_new_n5119_));
AND2X2 AND2X2_4736 ( .A(round_ctr_rst), .B(\block[295] ), .Y(w_mem_inst__abc_21203_new_n5120_));
AND2X2 AND2X2_4737 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5120_), .Y(w_mem_inst__abc_21203_new_n5121_));
AND2X2 AND2X2_4738 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_6__8_), .Y(w_mem_inst__abc_21203_new_n5124_));
AND2X2 AND2X2_4739 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_7__8_), .Y(w_mem_inst__abc_21203_new_n5125_));
AND2X2 AND2X2_474 ( .A(_abc_15497_new_n1672_), .B(_abc_15497_new_n1658_), .Y(_abc_15497_new_n1687_));
AND2X2 AND2X2_4740 ( .A(round_ctr_rst), .B(\block[296] ), .Y(w_mem_inst__abc_21203_new_n5126_));
AND2X2 AND2X2_4741 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5126_), .Y(w_mem_inst__abc_21203_new_n5127_));
AND2X2 AND2X2_4742 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_6__9_), .Y(w_mem_inst__abc_21203_new_n5130_));
AND2X2 AND2X2_4743 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_7__9_), .Y(w_mem_inst__abc_21203_new_n5131_));
AND2X2 AND2X2_4744 ( .A(round_ctr_rst), .B(\block[297] ), .Y(w_mem_inst__abc_21203_new_n5132_));
AND2X2 AND2X2_4745 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5132_), .Y(w_mem_inst__abc_21203_new_n5133_));
AND2X2 AND2X2_4746 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_6__10_), .Y(w_mem_inst__abc_21203_new_n5136_));
AND2X2 AND2X2_4747 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_7__10_), .Y(w_mem_inst__abc_21203_new_n5137_));
AND2X2 AND2X2_4748 ( .A(round_ctr_rst), .B(\block[298] ), .Y(w_mem_inst__abc_21203_new_n5138_));
AND2X2 AND2X2_4749 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5138_), .Y(w_mem_inst__abc_21203_new_n5139_));
AND2X2 AND2X2_475 ( .A(\digest[44] ), .B(d_reg_12_), .Y(_abc_15497_new_n1692_));
AND2X2 AND2X2_4750 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_6__11_), .Y(w_mem_inst__abc_21203_new_n5142_));
AND2X2 AND2X2_4751 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_7__11_), .Y(w_mem_inst__abc_21203_new_n5143_));
AND2X2 AND2X2_4752 ( .A(round_ctr_rst), .B(\block[299] ), .Y(w_mem_inst__abc_21203_new_n5144_));
AND2X2 AND2X2_4753 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5144_), .Y(w_mem_inst__abc_21203_new_n5145_));
AND2X2 AND2X2_4754 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_6__12_), .Y(w_mem_inst__abc_21203_new_n5148_));
AND2X2 AND2X2_4755 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_7__12_), .Y(w_mem_inst__abc_21203_new_n5149_));
AND2X2 AND2X2_4756 ( .A(round_ctr_rst), .B(\block[300] ), .Y(w_mem_inst__abc_21203_new_n5150_));
AND2X2 AND2X2_4757 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5150_), .Y(w_mem_inst__abc_21203_new_n5151_));
AND2X2 AND2X2_4758 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_6__13_), .Y(w_mem_inst__abc_21203_new_n5154_));
AND2X2 AND2X2_4759 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_7__13_), .Y(w_mem_inst__abc_21203_new_n5155_));
AND2X2 AND2X2_476 ( .A(_abc_15497_new_n1693_), .B(_abc_15497_new_n1691_), .Y(_abc_15497_new_n1694_));
AND2X2 AND2X2_4760 ( .A(round_ctr_rst), .B(\block[301] ), .Y(w_mem_inst__abc_21203_new_n5156_));
AND2X2 AND2X2_4761 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5156_), .Y(w_mem_inst__abc_21203_new_n5157_));
AND2X2 AND2X2_4762 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_6__14_), .Y(w_mem_inst__abc_21203_new_n5160_));
AND2X2 AND2X2_4763 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_7__14_), .Y(w_mem_inst__abc_21203_new_n5161_));
AND2X2 AND2X2_4764 ( .A(round_ctr_rst), .B(\block[302] ), .Y(w_mem_inst__abc_21203_new_n5162_));
AND2X2 AND2X2_4765 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5162_), .Y(w_mem_inst__abc_21203_new_n5163_));
AND2X2 AND2X2_4766 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_6__15_), .Y(w_mem_inst__abc_21203_new_n5166_));
AND2X2 AND2X2_4767 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_7__15_), .Y(w_mem_inst__abc_21203_new_n5167_));
AND2X2 AND2X2_4768 ( .A(round_ctr_rst), .B(\block[303] ), .Y(w_mem_inst__abc_21203_new_n5168_));
AND2X2 AND2X2_4769 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5168_), .Y(w_mem_inst__abc_21203_new_n5169_));
AND2X2 AND2X2_477 ( .A(_abc_15497_new_n1690_), .B(_abc_15497_new_n1694_), .Y(_abc_15497_new_n1696_));
AND2X2 AND2X2_4770 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_6__16_), .Y(w_mem_inst__abc_21203_new_n5172_));
AND2X2 AND2X2_4771 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_7__16_), .Y(w_mem_inst__abc_21203_new_n5173_));
AND2X2 AND2X2_4772 ( .A(round_ctr_rst), .B(\block[304] ), .Y(w_mem_inst__abc_21203_new_n5174_));
AND2X2 AND2X2_4773 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5174_), .Y(w_mem_inst__abc_21203_new_n5175_));
AND2X2 AND2X2_4774 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_6__17_), .Y(w_mem_inst__abc_21203_new_n5178_));
AND2X2 AND2X2_4775 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_7__17_), .Y(w_mem_inst__abc_21203_new_n5179_));
AND2X2 AND2X2_4776 ( .A(round_ctr_rst), .B(\block[305] ), .Y(w_mem_inst__abc_21203_new_n5180_));
AND2X2 AND2X2_4777 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5180_), .Y(w_mem_inst__abc_21203_new_n5181_));
AND2X2 AND2X2_4778 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_6__18_), .Y(w_mem_inst__abc_21203_new_n5184_));
AND2X2 AND2X2_4779 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_7__18_), .Y(w_mem_inst__abc_21203_new_n5185_));
AND2X2 AND2X2_478 ( .A(_abc_15497_new_n1697_), .B(_abc_15497_new_n1695_), .Y(_abc_15497_new_n1698_));
AND2X2 AND2X2_4780 ( .A(round_ctr_rst), .B(\block[306] ), .Y(w_mem_inst__abc_21203_new_n5186_));
AND2X2 AND2X2_4781 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5186_), .Y(w_mem_inst__abc_21203_new_n5187_));
AND2X2 AND2X2_4782 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_6__19_), .Y(w_mem_inst__abc_21203_new_n5190_));
AND2X2 AND2X2_4783 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_7__19_), .Y(w_mem_inst__abc_21203_new_n5191_));
AND2X2 AND2X2_4784 ( .A(round_ctr_rst), .B(\block[307] ), .Y(w_mem_inst__abc_21203_new_n5192_));
AND2X2 AND2X2_4785 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5192_), .Y(w_mem_inst__abc_21203_new_n5193_));
AND2X2 AND2X2_4786 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_6__20_), .Y(w_mem_inst__abc_21203_new_n5196_));
AND2X2 AND2X2_4787 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_7__20_), .Y(w_mem_inst__abc_21203_new_n5197_));
AND2X2 AND2X2_4788 ( .A(round_ctr_rst), .B(\block[308] ), .Y(w_mem_inst__abc_21203_new_n5198_));
AND2X2 AND2X2_4789 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5198_), .Y(w_mem_inst__abc_21203_new_n5199_));
AND2X2 AND2X2_479 ( .A(_abc_15497_new_n1698_), .B(digest_update), .Y(_abc_15497_new_n1699_));
AND2X2 AND2X2_4790 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_6__21_), .Y(w_mem_inst__abc_21203_new_n5202_));
AND2X2 AND2X2_4791 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_7__21_), .Y(w_mem_inst__abc_21203_new_n5203_));
AND2X2 AND2X2_4792 ( .A(round_ctr_rst), .B(\block[309] ), .Y(w_mem_inst__abc_21203_new_n5204_));
AND2X2 AND2X2_4793 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5204_), .Y(w_mem_inst__abc_21203_new_n5205_));
AND2X2 AND2X2_4794 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_6__22_), .Y(w_mem_inst__abc_21203_new_n5208_));
AND2X2 AND2X2_4795 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_7__22_), .Y(w_mem_inst__abc_21203_new_n5209_));
AND2X2 AND2X2_4796 ( .A(round_ctr_rst), .B(\block[310] ), .Y(w_mem_inst__abc_21203_new_n5210_));
AND2X2 AND2X2_4797 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5210_), .Y(w_mem_inst__abc_21203_new_n5211_));
AND2X2 AND2X2_4798 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_6__23_), .Y(w_mem_inst__abc_21203_new_n5214_));
AND2X2 AND2X2_4799 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_7__23_), .Y(w_mem_inst__abc_21203_new_n5215_));
AND2X2 AND2X2_48 ( .A(_abc_15497_new_n790_), .B(_abc_15497_new_n786_), .Y(_abc_15497_new_n791_));
AND2X2 AND2X2_480 ( .A(_abc_15497_new_n1700_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n1701_));
AND2X2 AND2X2_4800 ( .A(round_ctr_rst), .B(\block[311] ), .Y(w_mem_inst__abc_21203_new_n5216_));
AND2X2 AND2X2_4801 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5216_), .Y(w_mem_inst__abc_21203_new_n5217_));
AND2X2 AND2X2_4802 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_6__24_), .Y(w_mem_inst__abc_21203_new_n5220_));
AND2X2 AND2X2_4803 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_7__24_), .Y(w_mem_inst__abc_21203_new_n5221_));
AND2X2 AND2X2_4804 ( .A(round_ctr_rst), .B(\block[312] ), .Y(w_mem_inst__abc_21203_new_n5222_));
AND2X2 AND2X2_4805 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5222_), .Y(w_mem_inst__abc_21203_new_n5223_));
AND2X2 AND2X2_4806 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_6__25_), .Y(w_mem_inst__abc_21203_new_n5226_));
AND2X2 AND2X2_4807 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_7__25_), .Y(w_mem_inst__abc_21203_new_n5227_));
AND2X2 AND2X2_4808 ( .A(round_ctr_rst), .B(\block[313] ), .Y(w_mem_inst__abc_21203_new_n5228_));
AND2X2 AND2X2_4809 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5228_), .Y(w_mem_inst__abc_21203_new_n5229_));
AND2X2 AND2X2_481 ( .A(_abc_15497_new_n701_), .B(\digest[45] ), .Y(_abc_15497_new_n1703_));
AND2X2 AND2X2_4810 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_6__26_), .Y(w_mem_inst__abc_21203_new_n5232_));
AND2X2 AND2X2_4811 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_7__26_), .Y(w_mem_inst__abc_21203_new_n5233_));
AND2X2 AND2X2_4812 ( .A(round_ctr_rst), .B(\block[314] ), .Y(w_mem_inst__abc_21203_new_n5234_));
AND2X2 AND2X2_4813 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5234_), .Y(w_mem_inst__abc_21203_new_n5235_));
AND2X2 AND2X2_4814 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_6__27_), .Y(w_mem_inst__abc_21203_new_n5238_));
AND2X2 AND2X2_4815 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_7__27_), .Y(w_mem_inst__abc_21203_new_n5239_));
AND2X2 AND2X2_4816 ( .A(round_ctr_rst), .B(\block[315] ), .Y(w_mem_inst__abc_21203_new_n5240_));
AND2X2 AND2X2_4817 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5240_), .Y(w_mem_inst__abc_21203_new_n5241_));
AND2X2 AND2X2_4818 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_6__28_), .Y(w_mem_inst__abc_21203_new_n5244_));
AND2X2 AND2X2_4819 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_7__28_), .Y(w_mem_inst__abc_21203_new_n5245_));
AND2X2 AND2X2_482 ( .A(\digest[45] ), .B(d_reg_13_), .Y(_abc_15497_new_n1705_));
AND2X2 AND2X2_4820 ( .A(round_ctr_rst), .B(\block[316] ), .Y(w_mem_inst__abc_21203_new_n5246_));
AND2X2 AND2X2_4821 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5246_), .Y(w_mem_inst__abc_21203_new_n5247_));
AND2X2 AND2X2_4822 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_6__29_), .Y(w_mem_inst__abc_21203_new_n5250_));
AND2X2 AND2X2_4823 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_7__29_), .Y(w_mem_inst__abc_21203_new_n5251_));
AND2X2 AND2X2_4824 ( .A(round_ctr_rst), .B(\block[317] ), .Y(w_mem_inst__abc_21203_new_n5252_));
AND2X2 AND2X2_4825 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5252_), .Y(w_mem_inst__abc_21203_new_n5253_));
AND2X2 AND2X2_4826 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_6__30_), .Y(w_mem_inst__abc_21203_new_n5256_));
AND2X2 AND2X2_4827 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_7__30_), .Y(w_mem_inst__abc_21203_new_n5257_));
AND2X2 AND2X2_4828 ( .A(round_ctr_rst), .B(\block[318] ), .Y(w_mem_inst__abc_21203_new_n5258_));
AND2X2 AND2X2_4829 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5258_), .Y(w_mem_inst__abc_21203_new_n5259_));
AND2X2 AND2X2_483 ( .A(_abc_15497_new_n1706_), .B(_abc_15497_new_n1704_), .Y(_abc_15497_new_n1707_));
AND2X2 AND2X2_4830 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_6__31_), .Y(w_mem_inst__abc_21203_new_n5262_));
AND2X2 AND2X2_4831 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_7__31_), .Y(w_mem_inst__abc_21203_new_n5263_));
AND2X2 AND2X2_4832 ( .A(round_ctr_rst), .B(\block[319] ), .Y(w_mem_inst__abc_21203_new_n5264_));
AND2X2 AND2X2_4833 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5264_), .Y(w_mem_inst__abc_21203_new_n5265_));
AND2X2 AND2X2_4834 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_5__0_), .Y(w_mem_inst__abc_21203_new_n5268_));
AND2X2 AND2X2_4835 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_6__0_), .Y(w_mem_inst__abc_21203_new_n5269_));
AND2X2 AND2X2_4836 ( .A(round_ctr_rst), .B(\block[320] ), .Y(w_mem_inst__abc_21203_new_n5270_));
AND2X2 AND2X2_4837 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5270_), .Y(w_mem_inst__abc_21203_new_n5271_));
AND2X2 AND2X2_4838 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_5__1_), .Y(w_mem_inst__abc_21203_new_n5274_));
AND2X2 AND2X2_4839 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_6__1_), .Y(w_mem_inst__abc_21203_new_n5275_));
AND2X2 AND2X2_484 ( .A(_abc_15497_new_n1694_), .B(_abc_15497_new_n1707_), .Y(_abc_15497_new_n1710_));
AND2X2 AND2X2_4840 ( .A(round_ctr_rst), .B(\block[321] ), .Y(w_mem_inst__abc_21203_new_n5276_));
AND2X2 AND2X2_4841 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5276_), .Y(w_mem_inst__abc_21203_new_n5277_));
AND2X2 AND2X2_4842 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_5__2_), .Y(w_mem_inst__abc_21203_new_n5280_));
AND2X2 AND2X2_4843 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_6__2_), .Y(w_mem_inst__abc_21203_new_n5281_));
AND2X2 AND2X2_4844 ( .A(round_ctr_rst), .B(\block[322] ), .Y(w_mem_inst__abc_21203_new_n5282_));
AND2X2 AND2X2_4845 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5282_), .Y(w_mem_inst__abc_21203_new_n5283_));
AND2X2 AND2X2_4846 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_5__3_), .Y(w_mem_inst__abc_21203_new_n5286_));
AND2X2 AND2X2_4847 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_6__3_), .Y(w_mem_inst__abc_21203_new_n5287_));
AND2X2 AND2X2_4848 ( .A(round_ctr_rst), .B(\block[323] ), .Y(w_mem_inst__abc_21203_new_n5288_));
AND2X2 AND2X2_4849 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5288_), .Y(w_mem_inst__abc_21203_new_n5289_));
AND2X2 AND2X2_485 ( .A(_abc_15497_new_n1690_), .B(_abc_15497_new_n1710_), .Y(_abc_15497_new_n1711_));
AND2X2 AND2X2_4850 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_5__4_), .Y(w_mem_inst__abc_21203_new_n5292_));
AND2X2 AND2X2_4851 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_6__4_), .Y(w_mem_inst__abc_21203_new_n5293_));
AND2X2 AND2X2_4852 ( .A(round_ctr_rst), .B(\block[324] ), .Y(w_mem_inst__abc_21203_new_n5294_));
AND2X2 AND2X2_4853 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5294_), .Y(w_mem_inst__abc_21203_new_n5295_));
AND2X2 AND2X2_4854 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_5__5_), .Y(w_mem_inst__abc_21203_new_n5298_));
AND2X2 AND2X2_4855 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_6__5_), .Y(w_mem_inst__abc_21203_new_n5299_));
AND2X2 AND2X2_4856 ( .A(round_ctr_rst), .B(\block[325] ), .Y(w_mem_inst__abc_21203_new_n5300_));
AND2X2 AND2X2_4857 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5300_), .Y(w_mem_inst__abc_21203_new_n5301_));
AND2X2 AND2X2_4858 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_5__6_), .Y(w_mem_inst__abc_21203_new_n5304_));
AND2X2 AND2X2_4859 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_6__6_), .Y(w_mem_inst__abc_21203_new_n5305_));
AND2X2 AND2X2_486 ( .A(_abc_15497_new_n1707_), .B(_abc_15497_new_n1692_), .Y(_abc_15497_new_n1713_));
AND2X2 AND2X2_4860 ( .A(round_ctr_rst), .B(\block[326] ), .Y(w_mem_inst__abc_21203_new_n5306_));
AND2X2 AND2X2_4861 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5306_), .Y(w_mem_inst__abc_21203_new_n5307_));
AND2X2 AND2X2_4862 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_5__7_), .Y(w_mem_inst__abc_21203_new_n5310_));
AND2X2 AND2X2_4863 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_6__7_), .Y(w_mem_inst__abc_21203_new_n5311_));
AND2X2 AND2X2_4864 ( .A(round_ctr_rst), .B(\block[327] ), .Y(w_mem_inst__abc_21203_new_n5312_));
AND2X2 AND2X2_4865 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5312_), .Y(w_mem_inst__abc_21203_new_n5313_));
AND2X2 AND2X2_4866 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_5__8_), .Y(w_mem_inst__abc_21203_new_n5316_));
AND2X2 AND2X2_4867 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_6__8_), .Y(w_mem_inst__abc_21203_new_n5317_));
AND2X2 AND2X2_4868 ( .A(round_ctr_rst), .B(\block[328] ), .Y(w_mem_inst__abc_21203_new_n5318_));
AND2X2 AND2X2_4869 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5318_), .Y(w_mem_inst__abc_21203_new_n5319_));
AND2X2 AND2X2_487 ( .A(_abc_15497_new_n1714_), .B(digest_update), .Y(_abc_15497_new_n1715_));
AND2X2 AND2X2_4870 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_5__9_), .Y(w_mem_inst__abc_21203_new_n5322_));
AND2X2 AND2X2_4871 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_6__9_), .Y(w_mem_inst__abc_21203_new_n5323_));
AND2X2 AND2X2_4872 ( .A(round_ctr_rst), .B(\block[329] ), .Y(w_mem_inst__abc_21203_new_n5324_));
AND2X2 AND2X2_4873 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5324_), .Y(w_mem_inst__abc_21203_new_n5325_));
AND2X2 AND2X2_4874 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_5__10_), .Y(w_mem_inst__abc_21203_new_n5328_));
AND2X2 AND2X2_4875 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_6__10_), .Y(w_mem_inst__abc_21203_new_n5329_));
AND2X2 AND2X2_4876 ( .A(round_ctr_rst), .B(\block[330] ), .Y(w_mem_inst__abc_21203_new_n5330_));
AND2X2 AND2X2_4877 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5330_), .Y(w_mem_inst__abc_21203_new_n5331_));
AND2X2 AND2X2_4878 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_5__11_), .Y(w_mem_inst__abc_21203_new_n5334_));
AND2X2 AND2X2_4879 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_6__11_), .Y(w_mem_inst__abc_21203_new_n5335_));
AND2X2 AND2X2_488 ( .A(_abc_15497_new_n1712_), .B(_abc_15497_new_n1715_), .Y(_abc_15497_new_n1716_));
AND2X2 AND2X2_4880 ( .A(round_ctr_rst), .B(\block[331] ), .Y(w_mem_inst__abc_21203_new_n5336_));
AND2X2 AND2X2_4881 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5336_), .Y(w_mem_inst__abc_21203_new_n5337_));
AND2X2 AND2X2_4882 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_5__12_), .Y(w_mem_inst__abc_21203_new_n5340_));
AND2X2 AND2X2_4883 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_6__12_), .Y(w_mem_inst__abc_21203_new_n5341_));
AND2X2 AND2X2_4884 ( .A(round_ctr_rst), .B(\block[332] ), .Y(w_mem_inst__abc_21203_new_n5342_));
AND2X2 AND2X2_4885 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5342_), .Y(w_mem_inst__abc_21203_new_n5343_));
AND2X2 AND2X2_4886 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_5__13_), .Y(w_mem_inst__abc_21203_new_n5346_));
AND2X2 AND2X2_4887 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_6__13_), .Y(w_mem_inst__abc_21203_new_n5347_));
AND2X2 AND2X2_4888 ( .A(round_ctr_rst), .B(\block[333] ), .Y(w_mem_inst__abc_21203_new_n5348_));
AND2X2 AND2X2_4889 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5348_), .Y(w_mem_inst__abc_21203_new_n5349_));
AND2X2 AND2X2_489 ( .A(_abc_15497_new_n1716_), .B(_abc_15497_new_n1709_), .Y(_abc_15497_new_n1717_));
AND2X2 AND2X2_4890 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_5__14_), .Y(w_mem_inst__abc_21203_new_n5352_));
AND2X2 AND2X2_4891 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_6__14_), .Y(w_mem_inst__abc_21203_new_n5353_));
AND2X2 AND2X2_4892 ( .A(round_ctr_rst), .B(\block[334] ), .Y(w_mem_inst__abc_21203_new_n5354_));
AND2X2 AND2X2_4893 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5354_), .Y(w_mem_inst__abc_21203_new_n5355_));
AND2X2 AND2X2_4894 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_5__15_), .Y(w_mem_inst__abc_21203_new_n5358_));
AND2X2 AND2X2_4895 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_6__15_), .Y(w_mem_inst__abc_21203_new_n5359_));
AND2X2 AND2X2_4896 ( .A(round_ctr_rst), .B(\block[335] ), .Y(w_mem_inst__abc_21203_new_n5360_));
AND2X2 AND2X2_4897 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5360_), .Y(w_mem_inst__abc_21203_new_n5361_));
AND2X2 AND2X2_4898 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_5__16_), .Y(w_mem_inst__abc_21203_new_n5364_));
AND2X2 AND2X2_4899 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_6__16_), .Y(w_mem_inst__abc_21203_new_n5365_));
AND2X2 AND2X2_49 ( .A(_abc_15497_new_n792_), .B(_abc_15497_new_n793_), .Y(_abc_15497_new_n794_));
AND2X2 AND2X2_490 ( .A(_abc_15497_new_n1714_), .B(_abc_15497_new_n1706_), .Y(_abc_15497_new_n1719_));
AND2X2 AND2X2_4900 ( .A(round_ctr_rst), .B(\block[336] ), .Y(w_mem_inst__abc_21203_new_n5366_));
AND2X2 AND2X2_4901 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5366_), .Y(w_mem_inst__abc_21203_new_n5367_));
AND2X2 AND2X2_4902 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_5__17_), .Y(w_mem_inst__abc_21203_new_n5370_));
AND2X2 AND2X2_4903 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_6__17_), .Y(w_mem_inst__abc_21203_new_n5371_));
AND2X2 AND2X2_4904 ( .A(round_ctr_rst), .B(\block[337] ), .Y(w_mem_inst__abc_21203_new_n5372_));
AND2X2 AND2X2_4905 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5372_), .Y(w_mem_inst__abc_21203_new_n5373_));
AND2X2 AND2X2_4906 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_5__18_), .Y(w_mem_inst__abc_21203_new_n5376_));
AND2X2 AND2X2_4907 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_6__18_), .Y(w_mem_inst__abc_21203_new_n5377_));
AND2X2 AND2X2_4908 ( .A(round_ctr_rst), .B(\block[338] ), .Y(w_mem_inst__abc_21203_new_n5378_));
AND2X2 AND2X2_4909 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5378_), .Y(w_mem_inst__abc_21203_new_n5379_));
AND2X2 AND2X2_491 ( .A(_abc_15497_new_n1712_), .B(_abc_15497_new_n1719_), .Y(_abc_15497_new_n1720_));
AND2X2 AND2X2_4910 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_5__19_), .Y(w_mem_inst__abc_21203_new_n5382_));
AND2X2 AND2X2_4911 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_6__19_), .Y(w_mem_inst__abc_21203_new_n5383_));
AND2X2 AND2X2_4912 ( .A(round_ctr_rst), .B(\block[339] ), .Y(w_mem_inst__abc_21203_new_n5384_));
AND2X2 AND2X2_4913 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5384_), .Y(w_mem_inst__abc_21203_new_n5385_));
AND2X2 AND2X2_4914 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_5__20_), .Y(w_mem_inst__abc_21203_new_n5388_));
AND2X2 AND2X2_4915 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_6__20_), .Y(w_mem_inst__abc_21203_new_n5389_));
AND2X2 AND2X2_4916 ( .A(round_ctr_rst), .B(\block[340] ), .Y(w_mem_inst__abc_21203_new_n5390_));
AND2X2 AND2X2_4917 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5390_), .Y(w_mem_inst__abc_21203_new_n5391_));
AND2X2 AND2X2_4918 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_5__21_), .Y(w_mem_inst__abc_21203_new_n5394_));
AND2X2 AND2X2_4919 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_6__21_), .Y(w_mem_inst__abc_21203_new_n5395_));
AND2X2 AND2X2_492 ( .A(\digest[46] ), .B(d_reg_14_), .Y(_abc_15497_new_n1723_));
AND2X2 AND2X2_4920 ( .A(round_ctr_rst), .B(\block[341] ), .Y(w_mem_inst__abc_21203_new_n5396_));
AND2X2 AND2X2_4921 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5396_), .Y(w_mem_inst__abc_21203_new_n5397_));
AND2X2 AND2X2_4922 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_5__22_), .Y(w_mem_inst__abc_21203_new_n5400_));
AND2X2 AND2X2_4923 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_6__22_), .Y(w_mem_inst__abc_21203_new_n5401_));
AND2X2 AND2X2_4924 ( .A(round_ctr_rst), .B(\block[342] ), .Y(w_mem_inst__abc_21203_new_n5402_));
AND2X2 AND2X2_4925 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5402_), .Y(w_mem_inst__abc_21203_new_n5403_));
AND2X2 AND2X2_4926 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_5__23_), .Y(w_mem_inst__abc_21203_new_n5406_));
AND2X2 AND2X2_4927 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_6__23_), .Y(w_mem_inst__abc_21203_new_n5407_));
AND2X2 AND2X2_4928 ( .A(round_ctr_rst), .B(\block[343] ), .Y(w_mem_inst__abc_21203_new_n5408_));
AND2X2 AND2X2_4929 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5408_), .Y(w_mem_inst__abc_21203_new_n5409_));
AND2X2 AND2X2_493 ( .A(_abc_15497_new_n1724_), .B(_abc_15497_new_n1722_), .Y(_abc_15497_new_n1725_));
AND2X2 AND2X2_4930 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_5__24_), .Y(w_mem_inst__abc_21203_new_n5412_));
AND2X2 AND2X2_4931 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_6__24_), .Y(w_mem_inst__abc_21203_new_n5413_));
AND2X2 AND2X2_4932 ( .A(round_ctr_rst), .B(\block[344] ), .Y(w_mem_inst__abc_21203_new_n5414_));
AND2X2 AND2X2_4933 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5414_), .Y(w_mem_inst__abc_21203_new_n5415_));
AND2X2 AND2X2_4934 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_5__25_), .Y(w_mem_inst__abc_21203_new_n5418_));
AND2X2 AND2X2_4935 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_6__25_), .Y(w_mem_inst__abc_21203_new_n5419_));
AND2X2 AND2X2_4936 ( .A(round_ctr_rst), .B(\block[345] ), .Y(w_mem_inst__abc_21203_new_n5420_));
AND2X2 AND2X2_4937 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5420_), .Y(w_mem_inst__abc_21203_new_n5421_));
AND2X2 AND2X2_4938 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_5__26_), .Y(w_mem_inst__abc_21203_new_n5424_));
AND2X2 AND2X2_4939 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_6__26_), .Y(w_mem_inst__abc_21203_new_n5425_));
AND2X2 AND2X2_494 ( .A(_abc_15497_new_n1721_), .B(_abc_15497_new_n1725_), .Y(_abc_15497_new_n1727_));
AND2X2 AND2X2_4940 ( .A(round_ctr_rst), .B(\block[346] ), .Y(w_mem_inst__abc_21203_new_n5426_));
AND2X2 AND2X2_4941 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5426_), .Y(w_mem_inst__abc_21203_new_n5427_));
AND2X2 AND2X2_4942 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_5__27_), .Y(w_mem_inst__abc_21203_new_n5430_));
AND2X2 AND2X2_4943 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_6__27_), .Y(w_mem_inst__abc_21203_new_n5431_));
AND2X2 AND2X2_4944 ( .A(round_ctr_rst), .B(\block[347] ), .Y(w_mem_inst__abc_21203_new_n5432_));
AND2X2 AND2X2_4945 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5432_), .Y(w_mem_inst__abc_21203_new_n5433_));
AND2X2 AND2X2_4946 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_5__28_), .Y(w_mem_inst__abc_21203_new_n5436_));
AND2X2 AND2X2_4947 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_6__28_), .Y(w_mem_inst__abc_21203_new_n5437_));
AND2X2 AND2X2_4948 ( .A(round_ctr_rst), .B(\block[348] ), .Y(w_mem_inst__abc_21203_new_n5438_));
AND2X2 AND2X2_4949 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5438_), .Y(w_mem_inst__abc_21203_new_n5439_));
AND2X2 AND2X2_495 ( .A(_abc_15497_new_n1728_), .B(_abc_15497_new_n1726_), .Y(_abc_15497_new_n1729_));
AND2X2 AND2X2_4950 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_5__29_), .Y(w_mem_inst__abc_21203_new_n5442_));
AND2X2 AND2X2_4951 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_6__29_), .Y(w_mem_inst__abc_21203_new_n5443_));
AND2X2 AND2X2_4952 ( .A(round_ctr_rst), .B(\block[349] ), .Y(w_mem_inst__abc_21203_new_n5444_));
AND2X2 AND2X2_4953 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5444_), .Y(w_mem_inst__abc_21203_new_n5445_));
AND2X2 AND2X2_4954 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_5__30_), .Y(w_mem_inst__abc_21203_new_n5448_));
AND2X2 AND2X2_4955 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_6__30_), .Y(w_mem_inst__abc_21203_new_n5449_));
AND2X2 AND2X2_4956 ( .A(round_ctr_rst), .B(\block[350] ), .Y(w_mem_inst__abc_21203_new_n5450_));
AND2X2 AND2X2_4957 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5450_), .Y(w_mem_inst__abc_21203_new_n5451_));
AND2X2 AND2X2_4958 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_5__31_), .Y(w_mem_inst__abc_21203_new_n5454_));
AND2X2 AND2X2_4959 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_6__31_), .Y(w_mem_inst__abc_21203_new_n5455_));
AND2X2 AND2X2_496 ( .A(_abc_15497_new_n1729_), .B(digest_update), .Y(_abc_15497_new_n1730_));
AND2X2 AND2X2_4960 ( .A(round_ctr_rst), .B(\block[351] ), .Y(w_mem_inst__abc_21203_new_n5456_));
AND2X2 AND2X2_4961 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5456_), .Y(w_mem_inst__abc_21203_new_n5457_));
AND2X2 AND2X2_4962 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_1__0_), .Y(w_mem_inst__abc_21203_new_n5460_));
AND2X2 AND2X2_4963 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_2__0_), .Y(w_mem_inst__abc_21203_new_n5461_));
AND2X2 AND2X2_4964 ( .A(round_ctr_rst), .B(\block[448] ), .Y(w_mem_inst__abc_21203_new_n5462_));
AND2X2 AND2X2_4965 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5462_), .Y(w_mem_inst__abc_21203_new_n5463_));
AND2X2 AND2X2_4966 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_1__1_), .Y(w_mem_inst__abc_21203_new_n5466_));
AND2X2 AND2X2_4967 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_2__1_), .Y(w_mem_inst__abc_21203_new_n5467_));
AND2X2 AND2X2_4968 ( .A(round_ctr_rst), .B(\block[449] ), .Y(w_mem_inst__abc_21203_new_n5468_));
AND2X2 AND2X2_4969 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5468_), .Y(w_mem_inst__abc_21203_new_n5469_));
AND2X2 AND2X2_497 ( .A(_abc_15497_new_n1731_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n1732_));
AND2X2 AND2X2_4970 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_1__2_), .Y(w_mem_inst__abc_21203_new_n5472_));
AND2X2 AND2X2_4971 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_2__2_), .Y(w_mem_inst__abc_21203_new_n5473_));
AND2X2 AND2X2_4972 ( .A(round_ctr_rst), .B(\block[450] ), .Y(w_mem_inst__abc_21203_new_n5474_));
AND2X2 AND2X2_4973 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5474_), .Y(w_mem_inst__abc_21203_new_n5475_));
AND2X2 AND2X2_4974 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_1__3_), .Y(w_mem_inst__abc_21203_new_n5478_));
AND2X2 AND2X2_4975 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_2__3_), .Y(w_mem_inst__abc_21203_new_n5479_));
AND2X2 AND2X2_4976 ( .A(round_ctr_rst), .B(\block[451] ), .Y(w_mem_inst__abc_21203_new_n5480_));
AND2X2 AND2X2_4977 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5480_), .Y(w_mem_inst__abc_21203_new_n5481_));
AND2X2 AND2X2_4978 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_1__4_), .Y(w_mem_inst__abc_21203_new_n5484_));
AND2X2 AND2X2_4979 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_2__4_), .Y(w_mem_inst__abc_21203_new_n5485_));
AND2X2 AND2X2_498 ( .A(_abc_15497_new_n701_), .B(\digest[47] ), .Y(_abc_15497_new_n1734_));
AND2X2 AND2X2_4980 ( .A(round_ctr_rst), .B(\block[452] ), .Y(w_mem_inst__abc_21203_new_n5486_));
AND2X2 AND2X2_4981 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5486_), .Y(w_mem_inst__abc_21203_new_n5487_));
AND2X2 AND2X2_4982 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_1__5_), .Y(w_mem_inst__abc_21203_new_n5490_));
AND2X2 AND2X2_4983 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_2__5_), .Y(w_mem_inst__abc_21203_new_n5491_));
AND2X2 AND2X2_4984 ( .A(round_ctr_rst), .B(\block[453] ), .Y(w_mem_inst__abc_21203_new_n5492_));
AND2X2 AND2X2_4985 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5492_), .Y(w_mem_inst__abc_21203_new_n5493_));
AND2X2 AND2X2_4986 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_1__6_), .Y(w_mem_inst__abc_21203_new_n5496_));
AND2X2 AND2X2_4987 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_2__6_), .Y(w_mem_inst__abc_21203_new_n5497_));
AND2X2 AND2X2_4988 ( .A(round_ctr_rst), .B(\block[454] ), .Y(w_mem_inst__abc_21203_new_n5498_));
AND2X2 AND2X2_4989 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5498_), .Y(w_mem_inst__abc_21203_new_n5499_));
AND2X2 AND2X2_499 ( .A(_abc_15497_new_n1728_), .B(_abc_15497_new_n1724_), .Y(_abc_15497_new_n1735_));
AND2X2 AND2X2_4990 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_1__7_), .Y(w_mem_inst__abc_21203_new_n5502_));
AND2X2 AND2X2_4991 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_2__7_), .Y(w_mem_inst__abc_21203_new_n5503_));
AND2X2 AND2X2_4992 ( .A(round_ctr_rst), .B(\block[455] ), .Y(w_mem_inst__abc_21203_new_n5504_));
AND2X2 AND2X2_4993 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5504_), .Y(w_mem_inst__abc_21203_new_n5505_));
AND2X2 AND2X2_4994 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_1__8_), .Y(w_mem_inst__abc_21203_new_n5508_));
AND2X2 AND2X2_4995 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_2__8_), .Y(w_mem_inst__abc_21203_new_n5509_));
AND2X2 AND2X2_4996 ( .A(round_ctr_rst), .B(\block[456] ), .Y(w_mem_inst__abc_21203_new_n5510_));
AND2X2 AND2X2_4997 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5510_), .Y(w_mem_inst__abc_21203_new_n5511_));
AND2X2 AND2X2_4998 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_1__9_), .Y(w_mem_inst__abc_21203_new_n5514_));
AND2X2 AND2X2_4999 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_2__9_), .Y(w_mem_inst__abc_21203_new_n5515_));
AND2X2 AND2X2_5 ( .A(_abc_15497_new_n705_), .B(_abc_15497_new_n703_), .Y(_abc_15497_new_n706_));
AND2X2 AND2X2_50 ( .A(_abc_15497_new_n791_), .B(_abc_15497_new_n794_), .Y(_abc_15497_new_n795_));
AND2X2 AND2X2_500 ( .A(\digest[47] ), .B(d_reg_15_), .Y(_abc_15497_new_n1738_));
AND2X2 AND2X2_5000 ( .A(round_ctr_rst), .B(\block[457] ), .Y(w_mem_inst__abc_21203_new_n5516_));
AND2X2 AND2X2_5001 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5516_), .Y(w_mem_inst__abc_21203_new_n5517_));
AND2X2 AND2X2_5002 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_1__10_), .Y(w_mem_inst__abc_21203_new_n5520_));
AND2X2 AND2X2_5003 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_2__10_), .Y(w_mem_inst__abc_21203_new_n5521_));
AND2X2 AND2X2_5004 ( .A(round_ctr_rst), .B(\block[458] ), .Y(w_mem_inst__abc_21203_new_n5522_));
AND2X2 AND2X2_5005 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5522_), .Y(w_mem_inst__abc_21203_new_n5523_));
AND2X2 AND2X2_5006 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_1__11_), .Y(w_mem_inst__abc_21203_new_n5526_));
AND2X2 AND2X2_5007 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_2__11_), .Y(w_mem_inst__abc_21203_new_n5527_));
AND2X2 AND2X2_5008 ( .A(round_ctr_rst), .B(\block[459] ), .Y(w_mem_inst__abc_21203_new_n5528_));
AND2X2 AND2X2_5009 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5528_), .Y(w_mem_inst__abc_21203_new_n5529_));
AND2X2 AND2X2_501 ( .A(_abc_15497_new_n1739_), .B(_abc_15497_new_n1737_), .Y(_abc_15497_new_n1740_));
AND2X2 AND2X2_5010 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_1__12_), .Y(w_mem_inst__abc_21203_new_n5532_));
AND2X2 AND2X2_5011 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_2__12_), .Y(w_mem_inst__abc_21203_new_n5533_));
AND2X2 AND2X2_5012 ( .A(round_ctr_rst), .B(\block[460] ), .Y(w_mem_inst__abc_21203_new_n5534_));
AND2X2 AND2X2_5013 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5534_), .Y(w_mem_inst__abc_21203_new_n5535_));
AND2X2 AND2X2_5014 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_1__13_), .Y(w_mem_inst__abc_21203_new_n5538_));
AND2X2 AND2X2_5015 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_2__13_), .Y(w_mem_inst__abc_21203_new_n5539_));
AND2X2 AND2X2_5016 ( .A(round_ctr_rst), .B(\block[461] ), .Y(w_mem_inst__abc_21203_new_n5540_));
AND2X2 AND2X2_5017 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5540_), .Y(w_mem_inst__abc_21203_new_n5541_));
AND2X2 AND2X2_5018 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_1__14_), .Y(w_mem_inst__abc_21203_new_n5544_));
AND2X2 AND2X2_5019 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_2__14_), .Y(w_mem_inst__abc_21203_new_n5545_));
AND2X2 AND2X2_502 ( .A(_abc_15497_new_n1743_), .B(digest_update), .Y(_abc_15497_new_n1744_));
AND2X2 AND2X2_5020 ( .A(round_ctr_rst), .B(\block[462] ), .Y(w_mem_inst__abc_21203_new_n5546_));
AND2X2 AND2X2_5021 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5546_), .Y(w_mem_inst__abc_21203_new_n5547_));
AND2X2 AND2X2_5022 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_1__15_), .Y(w_mem_inst__abc_21203_new_n5550_));
AND2X2 AND2X2_5023 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_2__15_), .Y(w_mem_inst__abc_21203_new_n5551_));
AND2X2 AND2X2_5024 ( .A(round_ctr_rst), .B(\block[463] ), .Y(w_mem_inst__abc_21203_new_n5552_));
AND2X2 AND2X2_5025 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5552_), .Y(w_mem_inst__abc_21203_new_n5553_));
AND2X2 AND2X2_5026 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_1__16_), .Y(w_mem_inst__abc_21203_new_n5556_));
AND2X2 AND2X2_5027 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_2__16_), .Y(w_mem_inst__abc_21203_new_n5557_));
AND2X2 AND2X2_5028 ( .A(round_ctr_rst), .B(\block[464] ), .Y(w_mem_inst__abc_21203_new_n5558_));
AND2X2 AND2X2_5029 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5558_), .Y(w_mem_inst__abc_21203_new_n5559_));
AND2X2 AND2X2_503 ( .A(_abc_15497_new_n1744_), .B(_abc_15497_new_n1741_), .Y(_abc_15497_new_n1745_));
AND2X2 AND2X2_5030 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_1__17_), .Y(w_mem_inst__abc_21203_new_n5562_));
AND2X2 AND2X2_5031 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_2__17_), .Y(w_mem_inst__abc_21203_new_n5563_));
AND2X2 AND2X2_5032 ( .A(round_ctr_rst), .B(\block[465] ), .Y(w_mem_inst__abc_21203_new_n5564_));
AND2X2 AND2X2_5033 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5564_), .Y(w_mem_inst__abc_21203_new_n5565_));
AND2X2 AND2X2_5034 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_1__18_), .Y(w_mem_inst__abc_21203_new_n5568_));
AND2X2 AND2X2_5035 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_2__18_), .Y(w_mem_inst__abc_21203_new_n5569_));
AND2X2 AND2X2_5036 ( .A(round_ctr_rst), .B(\block[466] ), .Y(w_mem_inst__abc_21203_new_n5570_));
AND2X2 AND2X2_5037 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5570_), .Y(w_mem_inst__abc_21203_new_n5571_));
AND2X2 AND2X2_5038 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_1__19_), .Y(w_mem_inst__abc_21203_new_n5574_));
AND2X2 AND2X2_5039 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_2__19_), .Y(w_mem_inst__abc_21203_new_n5575_));
AND2X2 AND2X2_504 ( .A(_abc_15497_new_n701_), .B(\digest[48] ), .Y(_abc_15497_new_n1747_));
AND2X2 AND2X2_5040 ( .A(round_ctr_rst), .B(\block[467] ), .Y(w_mem_inst__abc_21203_new_n5576_));
AND2X2 AND2X2_5041 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5576_), .Y(w_mem_inst__abc_21203_new_n5577_));
AND2X2 AND2X2_5042 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_1__20_), .Y(w_mem_inst__abc_21203_new_n5580_));
AND2X2 AND2X2_5043 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_2__20_), .Y(w_mem_inst__abc_21203_new_n5581_));
AND2X2 AND2X2_5044 ( .A(round_ctr_rst), .B(\block[468] ), .Y(w_mem_inst__abc_21203_new_n5582_));
AND2X2 AND2X2_5045 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5582_), .Y(w_mem_inst__abc_21203_new_n5583_));
AND2X2 AND2X2_5046 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_1__21_), .Y(w_mem_inst__abc_21203_new_n5586_));
AND2X2 AND2X2_5047 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_2__21_), .Y(w_mem_inst__abc_21203_new_n5587_));
AND2X2 AND2X2_5048 ( .A(round_ctr_rst), .B(\block[469] ), .Y(w_mem_inst__abc_21203_new_n5588_));
AND2X2 AND2X2_5049 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5588_), .Y(w_mem_inst__abc_21203_new_n5589_));
AND2X2 AND2X2_505 ( .A(_abc_15497_new_n1725_), .B(_abc_15497_new_n1740_), .Y(_abc_15497_new_n1748_));
AND2X2 AND2X2_5050 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_1__22_), .Y(w_mem_inst__abc_21203_new_n5592_));
AND2X2 AND2X2_5051 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_2__22_), .Y(w_mem_inst__abc_21203_new_n5593_));
AND2X2 AND2X2_5052 ( .A(round_ctr_rst), .B(\block[470] ), .Y(w_mem_inst__abc_21203_new_n5594_));
AND2X2 AND2X2_5053 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5594_), .Y(w_mem_inst__abc_21203_new_n5595_));
AND2X2 AND2X2_5054 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_1__23_), .Y(w_mem_inst__abc_21203_new_n5598_));
AND2X2 AND2X2_5055 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_2__23_), .Y(w_mem_inst__abc_21203_new_n5599_));
AND2X2 AND2X2_5056 ( .A(round_ctr_rst), .B(\block[471] ), .Y(w_mem_inst__abc_21203_new_n5600_));
AND2X2 AND2X2_5057 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5600_), .Y(w_mem_inst__abc_21203_new_n5601_));
AND2X2 AND2X2_5058 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_1__24_), .Y(w_mem_inst__abc_21203_new_n5604_));
AND2X2 AND2X2_5059 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_2__24_), .Y(w_mem_inst__abc_21203_new_n5605_));
AND2X2 AND2X2_506 ( .A(_abc_15497_new_n1737_), .B(_abc_15497_new_n1723_), .Y(_abc_15497_new_n1751_));
AND2X2 AND2X2_5060 ( .A(round_ctr_rst), .B(\block[472] ), .Y(w_mem_inst__abc_21203_new_n5606_));
AND2X2 AND2X2_5061 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5606_), .Y(w_mem_inst__abc_21203_new_n5607_));
AND2X2 AND2X2_5062 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_1__25_), .Y(w_mem_inst__abc_21203_new_n5610_));
AND2X2 AND2X2_5063 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_2__25_), .Y(w_mem_inst__abc_21203_new_n5611_));
AND2X2 AND2X2_5064 ( .A(round_ctr_rst), .B(\block[473] ), .Y(w_mem_inst__abc_21203_new_n5612_));
AND2X2 AND2X2_5065 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5612_), .Y(w_mem_inst__abc_21203_new_n5613_));
AND2X2 AND2X2_5066 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_1__26_), .Y(w_mem_inst__abc_21203_new_n5616_));
AND2X2 AND2X2_5067 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_2__26_), .Y(w_mem_inst__abc_21203_new_n5617_));
AND2X2 AND2X2_5068 ( .A(round_ctr_rst), .B(\block[474] ), .Y(w_mem_inst__abc_21203_new_n5618_));
AND2X2 AND2X2_5069 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5618_), .Y(w_mem_inst__abc_21203_new_n5619_));
AND2X2 AND2X2_507 ( .A(_abc_15497_new_n1750_), .B(_abc_15497_new_n1753_), .Y(_abc_15497_new_n1754_));
AND2X2 AND2X2_5070 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_1__27_), .Y(w_mem_inst__abc_21203_new_n5622_));
AND2X2 AND2X2_5071 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_2__27_), .Y(w_mem_inst__abc_21203_new_n5623_));
AND2X2 AND2X2_5072 ( .A(round_ctr_rst), .B(\block[475] ), .Y(w_mem_inst__abc_21203_new_n5624_));
AND2X2 AND2X2_5073 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5624_), .Y(w_mem_inst__abc_21203_new_n5625_));
AND2X2 AND2X2_5074 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_1__28_), .Y(w_mem_inst__abc_21203_new_n5628_));
AND2X2 AND2X2_5075 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_2__28_), .Y(w_mem_inst__abc_21203_new_n5629_));
AND2X2 AND2X2_5076 ( .A(round_ctr_rst), .B(\block[476] ), .Y(w_mem_inst__abc_21203_new_n5630_));
AND2X2 AND2X2_5077 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5630_), .Y(w_mem_inst__abc_21203_new_n5631_));
AND2X2 AND2X2_5078 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_1__29_), .Y(w_mem_inst__abc_21203_new_n5634_));
AND2X2 AND2X2_5079 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_2__29_), .Y(w_mem_inst__abc_21203_new_n5635_));
AND2X2 AND2X2_508 ( .A(_abc_15497_new_n1710_), .B(_abc_15497_new_n1748_), .Y(_abc_15497_new_n1756_));
AND2X2 AND2X2_5080 ( .A(round_ctr_rst), .B(\block[477] ), .Y(w_mem_inst__abc_21203_new_n5636_));
AND2X2 AND2X2_5081 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5636_), .Y(w_mem_inst__abc_21203_new_n5637_));
AND2X2 AND2X2_5082 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_1__30_), .Y(w_mem_inst__abc_21203_new_n5640_));
AND2X2 AND2X2_5083 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_2__30_), .Y(w_mem_inst__abc_21203_new_n5641_));
AND2X2 AND2X2_5084 ( .A(round_ctr_rst), .B(\block[478] ), .Y(w_mem_inst__abc_21203_new_n5642_));
AND2X2 AND2X2_5085 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5642_), .Y(w_mem_inst__abc_21203_new_n5643_));
AND2X2 AND2X2_5086 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_1__31_), .Y(w_mem_inst__abc_21203_new_n5646_));
AND2X2 AND2X2_5087 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_2__31_), .Y(w_mem_inst__abc_21203_new_n5647_));
AND2X2 AND2X2_5088 ( .A(round_ctr_rst), .B(\block[479] ), .Y(w_mem_inst__abc_21203_new_n5648_));
AND2X2 AND2X2_5089 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5648_), .Y(w_mem_inst__abc_21203_new_n5649_));
AND2X2 AND2X2_509 ( .A(_abc_15497_new_n1690_), .B(_abc_15497_new_n1756_), .Y(_abc_15497_new_n1757_));
AND2X2 AND2X2_5090 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_3__0_), .Y(w_mem_inst__abc_21203_new_n5652_));
AND2X2 AND2X2_5091 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_4__0_), .Y(w_mem_inst__abc_21203_new_n5653_));
AND2X2 AND2X2_5092 ( .A(round_ctr_rst), .B(\block[384] ), .Y(w_mem_inst__abc_21203_new_n5654_));
AND2X2 AND2X2_5093 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5654_), .Y(w_mem_inst__abc_21203_new_n5655_));
AND2X2 AND2X2_5094 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_3__1_), .Y(w_mem_inst__abc_21203_new_n5658_));
AND2X2 AND2X2_5095 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_4__1_), .Y(w_mem_inst__abc_21203_new_n5659_));
AND2X2 AND2X2_5096 ( .A(round_ctr_rst), .B(\block[385] ), .Y(w_mem_inst__abc_21203_new_n5660_));
AND2X2 AND2X2_5097 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5660_), .Y(w_mem_inst__abc_21203_new_n5661_));
AND2X2 AND2X2_5098 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_3__2_), .Y(w_mem_inst__abc_21203_new_n5664_));
AND2X2 AND2X2_5099 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_4__2_), .Y(w_mem_inst__abc_21203_new_n5665_));
AND2X2 AND2X2_51 ( .A(c_reg_9_), .B(\digest[73] ), .Y(_abc_15497_new_n796_));
AND2X2 AND2X2_510 ( .A(\digest[48] ), .B(d_reg_16_), .Y(_abc_15497_new_n1760_));
AND2X2 AND2X2_5100 ( .A(round_ctr_rst), .B(\block[386] ), .Y(w_mem_inst__abc_21203_new_n5666_));
AND2X2 AND2X2_5101 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5666_), .Y(w_mem_inst__abc_21203_new_n5667_));
AND2X2 AND2X2_5102 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_3__3_), .Y(w_mem_inst__abc_21203_new_n5670_));
AND2X2 AND2X2_5103 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_4__3_), .Y(w_mem_inst__abc_21203_new_n5671_));
AND2X2 AND2X2_5104 ( .A(round_ctr_rst), .B(\block[387] ), .Y(w_mem_inst__abc_21203_new_n5672_));
AND2X2 AND2X2_5105 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5672_), .Y(w_mem_inst__abc_21203_new_n5673_));
AND2X2 AND2X2_5106 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_3__4_), .Y(w_mem_inst__abc_21203_new_n5676_));
AND2X2 AND2X2_5107 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_4__4_), .Y(w_mem_inst__abc_21203_new_n5677_));
AND2X2 AND2X2_5108 ( .A(round_ctr_rst), .B(\block[388] ), .Y(w_mem_inst__abc_21203_new_n5678_));
AND2X2 AND2X2_5109 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5678_), .Y(w_mem_inst__abc_21203_new_n5679_));
AND2X2 AND2X2_511 ( .A(_abc_15497_new_n1761_), .B(_abc_15497_new_n1759_), .Y(_abc_15497_new_n1762_));
AND2X2 AND2X2_5110 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_3__5_), .Y(w_mem_inst__abc_21203_new_n5682_));
AND2X2 AND2X2_5111 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_4__5_), .Y(w_mem_inst__abc_21203_new_n5683_));
AND2X2 AND2X2_5112 ( .A(round_ctr_rst), .B(\block[389] ), .Y(w_mem_inst__abc_21203_new_n5684_));
AND2X2 AND2X2_5113 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5684_), .Y(w_mem_inst__abc_21203_new_n5685_));
AND2X2 AND2X2_5114 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_3__6_), .Y(w_mem_inst__abc_21203_new_n5688_));
AND2X2 AND2X2_5115 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_4__6_), .Y(w_mem_inst__abc_21203_new_n5689_));
AND2X2 AND2X2_5116 ( .A(round_ctr_rst), .B(\block[390] ), .Y(w_mem_inst__abc_21203_new_n5690_));
AND2X2 AND2X2_5117 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5690_), .Y(w_mem_inst__abc_21203_new_n5691_));
AND2X2 AND2X2_5118 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_3__7_), .Y(w_mem_inst__abc_21203_new_n5694_));
AND2X2 AND2X2_5119 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_4__7_), .Y(w_mem_inst__abc_21203_new_n5695_));
AND2X2 AND2X2_512 ( .A(_abc_15497_new_n1758_), .B(_abc_15497_new_n1762_), .Y(_abc_15497_new_n1764_));
AND2X2 AND2X2_5120 ( .A(round_ctr_rst), .B(\block[391] ), .Y(w_mem_inst__abc_21203_new_n5696_));
AND2X2 AND2X2_5121 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5696_), .Y(w_mem_inst__abc_21203_new_n5697_));
AND2X2 AND2X2_5122 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_3__8_), .Y(w_mem_inst__abc_21203_new_n5700_));
AND2X2 AND2X2_5123 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_4__8_), .Y(w_mem_inst__abc_21203_new_n5701_));
AND2X2 AND2X2_5124 ( .A(round_ctr_rst), .B(\block[392] ), .Y(w_mem_inst__abc_21203_new_n5702_));
AND2X2 AND2X2_5125 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5702_), .Y(w_mem_inst__abc_21203_new_n5703_));
AND2X2 AND2X2_5126 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_3__9_), .Y(w_mem_inst__abc_21203_new_n5706_));
AND2X2 AND2X2_5127 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_4__9_), .Y(w_mem_inst__abc_21203_new_n5707_));
AND2X2 AND2X2_5128 ( .A(round_ctr_rst), .B(\block[393] ), .Y(w_mem_inst__abc_21203_new_n5708_));
AND2X2 AND2X2_5129 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5708_), .Y(w_mem_inst__abc_21203_new_n5709_));
AND2X2 AND2X2_513 ( .A(_abc_15497_new_n1765_), .B(_abc_15497_new_n1763_), .Y(_abc_15497_new_n1766_));
AND2X2 AND2X2_5130 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_3__10_), .Y(w_mem_inst__abc_21203_new_n5712_));
AND2X2 AND2X2_5131 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_4__10_), .Y(w_mem_inst__abc_21203_new_n5713_));
AND2X2 AND2X2_5132 ( .A(round_ctr_rst), .B(\block[394] ), .Y(w_mem_inst__abc_21203_new_n5714_));
AND2X2 AND2X2_5133 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5714_), .Y(w_mem_inst__abc_21203_new_n5715_));
AND2X2 AND2X2_5134 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_3__11_), .Y(w_mem_inst__abc_21203_new_n5718_));
AND2X2 AND2X2_5135 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_4__11_), .Y(w_mem_inst__abc_21203_new_n5719_));
AND2X2 AND2X2_5136 ( .A(round_ctr_rst), .B(\block[395] ), .Y(w_mem_inst__abc_21203_new_n5720_));
AND2X2 AND2X2_5137 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5720_), .Y(w_mem_inst__abc_21203_new_n5721_));
AND2X2 AND2X2_5138 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_3__12_), .Y(w_mem_inst__abc_21203_new_n5724_));
AND2X2 AND2X2_5139 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_4__12_), .Y(w_mem_inst__abc_21203_new_n5725_));
AND2X2 AND2X2_514 ( .A(_abc_15497_new_n1766_), .B(digest_update), .Y(_abc_15497_new_n1767_));
AND2X2 AND2X2_5140 ( .A(round_ctr_rst), .B(\block[396] ), .Y(w_mem_inst__abc_21203_new_n5726_));
AND2X2 AND2X2_5141 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5726_), .Y(w_mem_inst__abc_21203_new_n5727_));
AND2X2 AND2X2_5142 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_3__13_), .Y(w_mem_inst__abc_21203_new_n5730_));
AND2X2 AND2X2_5143 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_4__13_), .Y(w_mem_inst__abc_21203_new_n5731_));
AND2X2 AND2X2_5144 ( .A(round_ctr_rst), .B(\block[397] ), .Y(w_mem_inst__abc_21203_new_n5732_));
AND2X2 AND2X2_5145 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5732_), .Y(w_mem_inst__abc_21203_new_n5733_));
AND2X2 AND2X2_5146 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_3__14_), .Y(w_mem_inst__abc_21203_new_n5736_));
AND2X2 AND2X2_5147 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_4__14_), .Y(w_mem_inst__abc_21203_new_n5737_));
AND2X2 AND2X2_5148 ( .A(round_ctr_rst), .B(\block[398] ), .Y(w_mem_inst__abc_21203_new_n5738_));
AND2X2 AND2X2_5149 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5738_), .Y(w_mem_inst__abc_21203_new_n5739_));
AND2X2 AND2X2_515 ( .A(_abc_15497_new_n1765_), .B(_abc_15497_new_n1761_), .Y(_abc_15497_new_n1769_));
AND2X2 AND2X2_5150 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_3__15_), .Y(w_mem_inst__abc_21203_new_n5742_));
AND2X2 AND2X2_5151 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_4__15_), .Y(w_mem_inst__abc_21203_new_n5743_));
AND2X2 AND2X2_5152 ( .A(round_ctr_rst), .B(\block[399] ), .Y(w_mem_inst__abc_21203_new_n5744_));
AND2X2 AND2X2_5153 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5744_), .Y(w_mem_inst__abc_21203_new_n5745_));
AND2X2 AND2X2_5154 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_3__16_), .Y(w_mem_inst__abc_21203_new_n5748_));
AND2X2 AND2X2_5155 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_4__16_), .Y(w_mem_inst__abc_21203_new_n5749_));
AND2X2 AND2X2_5156 ( .A(round_ctr_rst), .B(\block[400] ), .Y(w_mem_inst__abc_21203_new_n5750_));
AND2X2 AND2X2_5157 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5750_), .Y(w_mem_inst__abc_21203_new_n5751_));
AND2X2 AND2X2_5158 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_3__17_), .Y(w_mem_inst__abc_21203_new_n5754_));
AND2X2 AND2X2_5159 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_4__17_), .Y(w_mem_inst__abc_21203_new_n5755_));
AND2X2 AND2X2_516 ( .A(\digest[49] ), .B(d_reg_17_), .Y(_abc_15497_new_n1771_));
AND2X2 AND2X2_5160 ( .A(round_ctr_rst), .B(\block[401] ), .Y(w_mem_inst__abc_21203_new_n5756_));
AND2X2 AND2X2_5161 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5756_), .Y(w_mem_inst__abc_21203_new_n5757_));
AND2X2 AND2X2_5162 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_3__18_), .Y(w_mem_inst__abc_21203_new_n5760_));
AND2X2 AND2X2_5163 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_4__18_), .Y(w_mem_inst__abc_21203_new_n5761_));
AND2X2 AND2X2_5164 ( .A(round_ctr_rst), .B(\block[402] ), .Y(w_mem_inst__abc_21203_new_n5762_));
AND2X2 AND2X2_5165 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5762_), .Y(w_mem_inst__abc_21203_new_n5763_));
AND2X2 AND2X2_5166 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_3__19_), .Y(w_mem_inst__abc_21203_new_n5766_));
AND2X2 AND2X2_5167 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_4__19_), .Y(w_mem_inst__abc_21203_new_n5767_));
AND2X2 AND2X2_5168 ( .A(round_ctr_rst), .B(\block[403] ), .Y(w_mem_inst__abc_21203_new_n5768_));
AND2X2 AND2X2_5169 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5768_), .Y(w_mem_inst__abc_21203_new_n5769_));
AND2X2 AND2X2_517 ( .A(_abc_15497_new_n1772_), .B(_abc_15497_new_n1770_), .Y(_abc_15497_new_n1773_));
AND2X2 AND2X2_5170 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_3__20_), .Y(w_mem_inst__abc_21203_new_n5772_));
AND2X2 AND2X2_5171 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_4__20_), .Y(w_mem_inst__abc_21203_new_n5773_));
AND2X2 AND2X2_5172 ( .A(round_ctr_rst), .B(\block[404] ), .Y(w_mem_inst__abc_21203_new_n5774_));
AND2X2 AND2X2_5173 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5774_), .Y(w_mem_inst__abc_21203_new_n5775_));
AND2X2 AND2X2_5174 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_3__21_), .Y(w_mem_inst__abc_21203_new_n5778_));
AND2X2 AND2X2_5175 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_4__21_), .Y(w_mem_inst__abc_21203_new_n5779_));
AND2X2 AND2X2_5176 ( .A(round_ctr_rst), .B(\block[405] ), .Y(w_mem_inst__abc_21203_new_n5780_));
AND2X2 AND2X2_5177 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5780_), .Y(w_mem_inst__abc_21203_new_n5781_));
AND2X2 AND2X2_5178 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_3__22_), .Y(w_mem_inst__abc_21203_new_n5784_));
AND2X2 AND2X2_5179 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_4__22_), .Y(w_mem_inst__abc_21203_new_n5785_));
AND2X2 AND2X2_518 ( .A(_abc_15497_new_n1769_), .B(_abc_15497_new_n1773_), .Y(_abc_15497_new_n1774_));
AND2X2 AND2X2_5180 ( .A(round_ctr_rst), .B(\block[406] ), .Y(w_mem_inst__abc_21203_new_n5786_));
AND2X2 AND2X2_5181 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5786_), .Y(w_mem_inst__abc_21203_new_n5787_));
AND2X2 AND2X2_5182 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_3__23_), .Y(w_mem_inst__abc_21203_new_n5790_));
AND2X2 AND2X2_5183 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_4__23_), .Y(w_mem_inst__abc_21203_new_n5791_));
AND2X2 AND2X2_5184 ( .A(round_ctr_rst), .B(\block[407] ), .Y(w_mem_inst__abc_21203_new_n5792_));
AND2X2 AND2X2_5185 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5792_), .Y(w_mem_inst__abc_21203_new_n5793_));
AND2X2 AND2X2_5186 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_3__24_), .Y(w_mem_inst__abc_21203_new_n5796_));
AND2X2 AND2X2_5187 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_4__24_), .Y(w_mem_inst__abc_21203_new_n5797_));
AND2X2 AND2X2_5188 ( .A(round_ctr_rst), .B(\block[408] ), .Y(w_mem_inst__abc_21203_new_n5798_));
AND2X2 AND2X2_5189 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5798_), .Y(w_mem_inst__abc_21203_new_n5799_));
AND2X2 AND2X2_519 ( .A(_abc_15497_new_n1775_), .B(_abc_15497_new_n1776_), .Y(_abc_15497_new_n1777_));
AND2X2 AND2X2_5190 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_3__25_), .Y(w_mem_inst__abc_21203_new_n5802_));
AND2X2 AND2X2_5191 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_4__25_), .Y(w_mem_inst__abc_21203_new_n5803_));
AND2X2 AND2X2_5192 ( .A(round_ctr_rst), .B(\block[409] ), .Y(w_mem_inst__abc_21203_new_n5804_));
AND2X2 AND2X2_5193 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5804_), .Y(w_mem_inst__abc_21203_new_n5805_));
AND2X2 AND2X2_5194 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_3__26_), .Y(w_mem_inst__abc_21203_new_n5808_));
AND2X2 AND2X2_5195 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_4__26_), .Y(w_mem_inst__abc_21203_new_n5809_));
AND2X2 AND2X2_5196 ( .A(round_ctr_rst), .B(\block[410] ), .Y(w_mem_inst__abc_21203_new_n5810_));
AND2X2 AND2X2_5197 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5810_), .Y(w_mem_inst__abc_21203_new_n5811_));
AND2X2 AND2X2_5198 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_3__27_), .Y(w_mem_inst__abc_21203_new_n5814_));
AND2X2 AND2X2_5199 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_4__27_), .Y(w_mem_inst__abc_21203_new_n5815_));
AND2X2 AND2X2_52 ( .A(c_reg_8_), .B(\digest[72] ), .Y(_abc_15497_new_n798_));
AND2X2 AND2X2_520 ( .A(_abc_15497_new_n1778_), .B(digest_update), .Y(_abc_15497_new_n1779_));
AND2X2 AND2X2_5200 ( .A(round_ctr_rst), .B(\block[411] ), .Y(w_mem_inst__abc_21203_new_n5816_));
AND2X2 AND2X2_5201 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5816_), .Y(w_mem_inst__abc_21203_new_n5817_));
AND2X2 AND2X2_5202 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_3__28_), .Y(w_mem_inst__abc_21203_new_n5820_));
AND2X2 AND2X2_5203 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_4__28_), .Y(w_mem_inst__abc_21203_new_n5821_));
AND2X2 AND2X2_5204 ( .A(round_ctr_rst), .B(\block[412] ), .Y(w_mem_inst__abc_21203_new_n5822_));
AND2X2 AND2X2_5205 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5822_), .Y(w_mem_inst__abc_21203_new_n5823_));
AND2X2 AND2X2_5206 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_3__29_), .Y(w_mem_inst__abc_21203_new_n5826_));
AND2X2 AND2X2_5207 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_4__29_), .Y(w_mem_inst__abc_21203_new_n5827_));
AND2X2 AND2X2_5208 ( .A(round_ctr_rst), .B(\block[413] ), .Y(w_mem_inst__abc_21203_new_n5828_));
AND2X2 AND2X2_5209 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5828_), .Y(w_mem_inst__abc_21203_new_n5829_));
AND2X2 AND2X2_521 ( .A(_abc_15497_new_n1780_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n1781_));
AND2X2 AND2X2_5210 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_3__30_), .Y(w_mem_inst__abc_21203_new_n5832_));
AND2X2 AND2X2_5211 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_4__30_), .Y(w_mem_inst__abc_21203_new_n5833_));
AND2X2 AND2X2_5212 ( .A(round_ctr_rst), .B(\block[414] ), .Y(w_mem_inst__abc_21203_new_n5834_));
AND2X2 AND2X2_5213 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5834_), .Y(w_mem_inst__abc_21203_new_n5835_));
AND2X2 AND2X2_5214 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_3__31_), .Y(w_mem_inst__abc_21203_new_n5838_));
AND2X2 AND2X2_5215 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_4__31_), .Y(w_mem_inst__abc_21203_new_n5839_));
AND2X2 AND2X2_5216 ( .A(round_ctr_rst), .B(\block[415] ), .Y(w_mem_inst__abc_21203_new_n5840_));
AND2X2 AND2X2_5217 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5840_), .Y(w_mem_inst__abc_21203_new_n5841_));
AND2X2 AND2X2_5218 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_2__0_), .Y(w_mem_inst__abc_21203_new_n5844_));
AND2X2 AND2X2_5219 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_3__0_), .Y(w_mem_inst__abc_21203_new_n5845_));
AND2X2 AND2X2_522 ( .A(_abc_15497_new_n701_), .B(\digest[50] ), .Y(_abc_15497_new_n1783_));
AND2X2 AND2X2_5220 ( .A(round_ctr_rst), .B(\block[416] ), .Y(w_mem_inst__abc_21203_new_n5846_));
AND2X2 AND2X2_5221 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5846_), .Y(w_mem_inst__abc_21203_new_n5847_));
AND2X2 AND2X2_5222 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_2__1_), .Y(w_mem_inst__abc_21203_new_n5850_));
AND2X2 AND2X2_5223 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_3__1_), .Y(w_mem_inst__abc_21203_new_n5851_));
AND2X2 AND2X2_5224 ( .A(round_ctr_rst), .B(\block[417] ), .Y(w_mem_inst__abc_21203_new_n5852_));
AND2X2 AND2X2_5225 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5852_), .Y(w_mem_inst__abc_21203_new_n5853_));
AND2X2 AND2X2_5226 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_2__2_), .Y(w_mem_inst__abc_21203_new_n5856_));
AND2X2 AND2X2_5227 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_3__2_), .Y(w_mem_inst__abc_21203_new_n5857_));
AND2X2 AND2X2_5228 ( .A(round_ctr_rst), .B(\block[418] ), .Y(w_mem_inst__abc_21203_new_n5858_));
AND2X2 AND2X2_5229 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5858_), .Y(w_mem_inst__abc_21203_new_n5859_));
AND2X2 AND2X2_523 ( .A(_abc_15497_new_n1773_), .B(_abc_15497_new_n1760_), .Y(_abc_15497_new_n1784_));
AND2X2 AND2X2_5230 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_2__3_), .Y(w_mem_inst__abc_21203_new_n5862_));
AND2X2 AND2X2_5231 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_3__3_), .Y(w_mem_inst__abc_21203_new_n5863_));
AND2X2 AND2X2_5232 ( .A(round_ctr_rst), .B(\block[419] ), .Y(w_mem_inst__abc_21203_new_n5864_));
AND2X2 AND2X2_5233 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5864_), .Y(w_mem_inst__abc_21203_new_n5865_));
AND2X2 AND2X2_5234 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_2__4_), .Y(w_mem_inst__abc_21203_new_n5868_));
AND2X2 AND2X2_5235 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_3__4_), .Y(w_mem_inst__abc_21203_new_n5869_));
AND2X2 AND2X2_5236 ( .A(round_ctr_rst), .B(\block[420] ), .Y(w_mem_inst__abc_21203_new_n5870_));
AND2X2 AND2X2_5237 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5870_), .Y(w_mem_inst__abc_21203_new_n5871_));
AND2X2 AND2X2_5238 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_2__5_), .Y(w_mem_inst__abc_21203_new_n5874_));
AND2X2 AND2X2_5239 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_3__5_), .Y(w_mem_inst__abc_21203_new_n5875_));
AND2X2 AND2X2_524 ( .A(_abc_15497_new_n1762_), .B(_abc_15497_new_n1773_), .Y(_abc_15497_new_n1786_));
AND2X2 AND2X2_5240 ( .A(round_ctr_rst), .B(\block[421] ), .Y(w_mem_inst__abc_21203_new_n5876_));
AND2X2 AND2X2_5241 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5876_), .Y(w_mem_inst__abc_21203_new_n5877_));
AND2X2 AND2X2_5242 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_2__6_), .Y(w_mem_inst__abc_21203_new_n5880_));
AND2X2 AND2X2_5243 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_3__6_), .Y(w_mem_inst__abc_21203_new_n5881_));
AND2X2 AND2X2_5244 ( .A(round_ctr_rst), .B(\block[422] ), .Y(w_mem_inst__abc_21203_new_n5882_));
AND2X2 AND2X2_5245 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5882_), .Y(w_mem_inst__abc_21203_new_n5883_));
AND2X2 AND2X2_5246 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_2__7_), .Y(w_mem_inst__abc_21203_new_n5886_));
AND2X2 AND2X2_5247 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_3__7_), .Y(w_mem_inst__abc_21203_new_n5887_));
AND2X2 AND2X2_5248 ( .A(round_ctr_rst), .B(\block[423] ), .Y(w_mem_inst__abc_21203_new_n5888_));
AND2X2 AND2X2_5249 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5888_), .Y(w_mem_inst__abc_21203_new_n5889_));
AND2X2 AND2X2_525 ( .A(_abc_15497_new_n1758_), .B(_abc_15497_new_n1786_), .Y(_abc_15497_new_n1787_));
AND2X2 AND2X2_5250 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_2__8_), .Y(w_mem_inst__abc_21203_new_n5892_));
AND2X2 AND2X2_5251 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_3__8_), .Y(w_mem_inst__abc_21203_new_n5893_));
AND2X2 AND2X2_5252 ( .A(round_ctr_rst), .B(\block[424] ), .Y(w_mem_inst__abc_21203_new_n5894_));
AND2X2 AND2X2_5253 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5894_), .Y(w_mem_inst__abc_21203_new_n5895_));
AND2X2 AND2X2_5254 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_2__9_), .Y(w_mem_inst__abc_21203_new_n5898_));
AND2X2 AND2X2_5255 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_3__9_), .Y(w_mem_inst__abc_21203_new_n5899_));
AND2X2 AND2X2_5256 ( .A(round_ctr_rst), .B(\block[425] ), .Y(w_mem_inst__abc_21203_new_n5900_));
AND2X2 AND2X2_5257 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5900_), .Y(w_mem_inst__abc_21203_new_n5901_));
AND2X2 AND2X2_5258 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_2__10_), .Y(w_mem_inst__abc_21203_new_n5904_));
AND2X2 AND2X2_5259 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_3__10_), .Y(w_mem_inst__abc_21203_new_n5905_));
AND2X2 AND2X2_526 ( .A(\digest[50] ), .B(d_reg_18_), .Y(_abc_15497_new_n1790_));
AND2X2 AND2X2_5260 ( .A(round_ctr_rst), .B(\block[426] ), .Y(w_mem_inst__abc_21203_new_n5906_));
AND2X2 AND2X2_5261 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5906_), .Y(w_mem_inst__abc_21203_new_n5907_));
AND2X2 AND2X2_5262 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_2__11_), .Y(w_mem_inst__abc_21203_new_n5910_));
AND2X2 AND2X2_5263 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_3__11_), .Y(w_mem_inst__abc_21203_new_n5911_));
AND2X2 AND2X2_5264 ( .A(round_ctr_rst), .B(\block[427] ), .Y(w_mem_inst__abc_21203_new_n5912_));
AND2X2 AND2X2_5265 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5912_), .Y(w_mem_inst__abc_21203_new_n5913_));
AND2X2 AND2X2_5266 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_2__12_), .Y(w_mem_inst__abc_21203_new_n5916_));
AND2X2 AND2X2_5267 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_3__12_), .Y(w_mem_inst__abc_21203_new_n5917_));
AND2X2 AND2X2_5268 ( .A(round_ctr_rst), .B(\block[428] ), .Y(w_mem_inst__abc_21203_new_n5918_));
AND2X2 AND2X2_5269 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5918_), .Y(w_mem_inst__abc_21203_new_n5919_));
AND2X2 AND2X2_527 ( .A(_abc_15497_new_n1791_), .B(_abc_15497_new_n1789_), .Y(_abc_15497_new_n1792_));
AND2X2 AND2X2_5270 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_2__13_), .Y(w_mem_inst__abc_21203_new_n5922_));
AND2X2 AND2X2_5271 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_3__13_), .Y(w_mem_inst__abc_21203_new_n5923_));
AND2X2 AND2X2_5272 ( .A(round_ctr_rst), .B(\block[429] ), .Y(w_mem_inst__abc_21203_new_n5924_));
AND2X2 AND2X2_5273 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5924_), .Y(w_mem_inst__abc_21203_new_n5925_));
AND2X2 AND2X2_5274 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_2__14_), .Y(w_mem_inst__abc_21203_new_n5928_));
AND2X2 AND2X2_5275 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_3__14_), .Y(w_mem_inst__abc_21203_new_n5929_));
AND2X2 AND2X2_5276 ( .A(round_ctr_rst), .B(\block[430] ), .Y(w_mem_inst__abc_21203_new_n5930_));
AND2X2 AND2X2_5277 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5930_), .Y(w_mem_inst__abc_21203_new_n5931_));
AND2X2 AND2X2_5278 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_2__15_), .Y(w_mem_inst__abc_21203_new_n5934_));
AND2X2 AND2X2_5279 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_3__15_), .Y(w_mem_inst__abc_21203_new_n5935_));
AND2X2 AND2X2_528 ( .A(_abc_15497_new_n1788_), .B(_abc_15497_new_n1792_), .Y(_abc_15497_new_n1794_));
AND2X2 AND2X2_5280 ( .A(round_ctr_rst), .B(\block[431] ), .Y(w_mem_inst__abc_21203_new_n5936_));
AND2X2 AND2X2_5281 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5936_), .Y(w_mem_inst__abc_21203_new_n5937_));
AND2X2 AND2X2_5282 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_2__16_), .Y(w_mem_inst__abc_21203_new_n5940_));
AND2X2 AND2X2_5283 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_3__16_), .Y(w_mem_inst__abc_21203_new_n5941_));
AND2X2 AND2X2_5284 ( .A(round_ctr_rst), .B(\block[432] ), .Y(w_mem_inst__abc_21203_new_n5942_));
AND2X2 AND2X2_5285 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5942_), .Y(w_mem_inst__abc_21203_new_n5943_));
AND2X2 AND2X2_5286 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_2__17_), .Y(w_mem_inst__abc_21203_new_n5946_));
AND2X2 AND2X2_5287 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_3__17_), .Y(w_mem_inst__abc_21203_new_n5947_));
AND2X2 AND2X2_5288 ( .A(round_ctr_rst), .B(\block[433] ), .Y(w_mem_inst__abc_21203_new_n5948_));
AND2X2 AND2X2_5289 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5948_), .Y(w_mem_inst__abc_21203_new_n5949_));
AND2X2 AND2X2_529 ( .A(_abc_15497_new_n1795_), .B(_abc_15497_new_n1793_), .Y(_abc_15497_new_n1796_));
AND2X2 AND2X2_5290 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_2__18_), .Y(w_mem_inst__abc_21203_new_n5952_));
AND2X2 AND2X2_5291 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_3__18_), .Y(w_mem_inst__abc_21203_new_n5953_));
AND2X2 AND2X2_5292 ( .A(round_ctr_rst), .B(\block[434] ), .Y(w_mem_inst__abc_21203_new_n5954_));
AND2X2 AND2X2_5293 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5954_), .Y(w_mem_inst__abc_21203_new_n5955_));
AND2X2 AND2X2_5294 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_2__19_), .Y(w_mem_inst__abc_21203_new_n5958_));
AND2X2 AND2X2_5295 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_3__19_), .Y(w_mem_inst__abc_21203_new_n5959_));
AND2X2 AND2X2_5296 ( .A(round_ctr_rst), .B(\block[435] ), .Y(w_mem_inst__abc_21203_new_n5960_));
AND2X2 AND2X2_5297 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5960_), .Y(w_mem_inst__abc_21203_new_n5961_));
AND2X2 AND2X2_5298 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_2__20_), .Y(w_mem_inst__abc_21203_new_n5964_));
AND2X2 AND2X2_5299 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_3__20_), .Y(w_mem_inst__abc_21203_new_n5965_));
AND2X2 AND2X2_53 ( .A(_abc_15497_new_n797_), .B(_abc_15497_new_n798_), .Y(_abc_15497_new_n799_));
AND2X2 AND2X2_530 ( .A(_abc_15497_new_n1796_), .B(digest_update), .Y(_abc_15497_new_n1797_));
AND2X2 AND2X2_5300 ( .A(round_ctr_rst), .B(\block[436] ), .Y(w_mem_inst__abc_21203_new_n5966_));
AND2X2 AND2X2_5301 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5966_), .Y(w_mem_inst__abc_21203_new_n5967_));
AND2X2 AND2X2_5302 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_2__21_), .Y(w_mem_inst__abc_21203_new_n5970_));
AND2X2 AND2X2_5303 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_3__21_), .Y(w_mem_inst__abc_21203_new_n5971_));
AND2X2 AND2X2_5304 ( .A(round_ctr_rst), .B(\block[437] ), .Y(w_mem_inst__abc_21203_new_n5972_));
AND2X2 AND2X2_5305 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5972_), .Y(w_mem_inst__abc_21203_new_n5973_));
AND2X2 AND2X2_5306 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_2__22_), .Y(w_mem_inst__abc_21203_new_n5976_));
AND2X2 AND2X2_5307 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_3__22_), .Y(w_mem_inst__abc_21203_new_n5977_));
AND2X2 AND2X2_5308 ( .A(round_ctr_rst), .B(\block[438] ), .Y(w_mem_inst__abc_21203_new_n5978_));
AND2X2 AND2X2_5309 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5978_), .Y(w_mem_inst__abc_21203_new_n5979_));
AND2X2 AND2X2_531 ( .A(_abc_15497_new_n701_), .B(\digest[51] ), .Y(_abc_15497_new_n1799_));
AND2X2 AND2X2_5310 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_2__23_), .Y(w_mem_inst__abc_21203_new_n5982_));
AND2X2 AND2X2_5311 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_3__23_), .Y(w_mem_inst__abc_21203_new_n5983_));
AND2X2 AND2X2_5312 ( .A(round_ctr_rst), .B(\block[439] ), .Y(w_mem_inst__abc_21203_new_n5984_));
AND2X2 AND2X2_5313 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5984_), .Y(w_mem_inst__abc_21203_new_n5985_));
AND2X2 AND2X2_5314 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_2__24_), .Y(w_mem_inst__abc_21203_new_n5988_));
AND2X2 AND2X2_5315 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_3__24_), .Y(w_mem_inst__abc_21203_new_n5989_));
AND2X2 AND2X2_5316 ( .A(round_ctr_rst), .B(\block[440] ), .Y(w_mem_inst__abc_21203_new_n5990_));
AND2X2 AND2X2_5317 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5990_), .Y(w_mem_inst__abc_21203_new_n5991_));
AND2X2 AND2X2_5318 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_2__25_), .Y(w_mem_inst__abc_21203_new_n5994_));
AND2X2 AND2X2_5319 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_3__25_), .Y(w_mem_inst__abc_21203_new_n5995_));
AND2X2 AND2X2_532 ( .A(_abc_15497_new_n1795_), .B(_abc_15497_new_n1791_), .Y(_abc_15497_new_n1800_));
AND2X2 AND2X2_5320 ( .A(round_ctr_rst), .B(\block[441] ), .Y(w_mem_inst__abc_21203_new_n5996_));
AND2X2 AND2X2_5321 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n5996_), .Y(w_mem_inst__abc_21203_new_n5997_));
AND2X2 AND2X2_5322 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_2__26_), .Y(w_mem_inst__abc_21203_new_n6000_));
AND2X2 AND2X2_5323 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_3__26_), .Y(w_mem_inst__abc_21203_new_n6001_));
AND2X2 AND2X2_5324 ( .A(round_ctr_rst), .B(\block[442] ), .Y(w_mem_inst__abc_21203_new_n6002_));
AND2X2 AND2X2_5325 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n6002_), .Y(w_mem_inst__abc_21203_new_n6003_));
AND2X2 AND2X2_5326 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_2__27_), .Y(w_mem_inst__abc_21203_new_n6006_));
AND2X2 AND2X2_5327 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_3__27_), .Y(w_mem_inst__abc_21203_new_n6007_));
AND2X2 AND2X2_5328 ( .A(round_ctr_rst), .B(\block[443] ), .Y(w_mem_inst__abc_21203_new_n6008_));
AND2X2 AND2X2_5329 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n6008_), .Y(w_mem_inst__abc_21203_new_n6009_));
AND2X2 AND2X2_533 ( .A(\digest[51] ), .B(d_reg_19_), .Y(_abc_15497_new_n1803_));
AND2X2 AND2X2_5330 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_2__28_), .Y(w_mem_inst__abc_21203_new_n6012_));
AND2X2 AND2X2_5331 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_3__28_), .Y(w_mem_inst__abc_21203_new_n6013_));
AND2X2 AND2X2_5332 ( .A(round_ctr_rst), .B(\block[444] ), .Y(w_mem_inst__abc_21203_new_n6014_));
AND2X2 AND2X2_5333 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n6014_), .Y(w_mem_inst__abc_21203_new_n6015_));
AND2X2 AND2X2_5334 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_2__29_), .Y(w_mem_inst__abc_21203_new_n6018_));
AND2X2 AND2X2_5335 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_3__29_), .Y(w_mem_inst__abc_21203_new_n6019_));
AND2X2 AND2X2_5336 ( .A(round_ctr_rst), .B(\block[445] ), .Y(w_mem_inst__abc_21203_new_n6020_));
AND2X2 AND2X2_5337 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n6020_), .Y(w_mem_inst__abc_21203_new_n6021_));
AND2X2 AND2X2_5338 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_2__30_), .Y(w_mem_inst__abc_21203_new_n6024_));
AND2X2 AND2X2_5339 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_3__30_), .Y(w_mem_inst__abc_21203_new_n6025_));
AND2X2 AND2X2_534 ( .A(_abc_15497_new_n1804_), .B(_abc_15497_new_n1802_), .Y(_abc_15497_new_n1805_));
AND2X2 AND2X2_5340 ( .A(round_ctr_rst), .B(\block[446] ), .Y(w_mem_inst__abc_21203_new_n6026_));
AND2X2 AND2X2_5341 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n6026_), .Y(w_mem_inst__abc_21203_new_n6027_));
AND2X2 AND2X2_5342 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_2__31_), .Y(w_mem_inst__abc_21203_new_n6030_));
AND2X2 AND2X2_5343 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_3__31_), .Y(w_mem_inst__abc_21203_new_n6031_));
AND2X2 AND2X2_5344 ( .A(round_ctr_rst), .B(\block[447] ), .Y(w_mem_inst__abc_21203_new_n6032_));
AND2X2 AND2X2_5345 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n6032_), .Y(w_mem_inst__abc_21203_new_n6033_));
AND2X2 AND2X2_5346 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_0__0_), .Y(w_mem_inst__abc_21203_new_n6036_));
AND2X2 AND2X2_5347 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_1__0_), .Y(w_mem_inst__abc_21203_new_n6037_));
AND2X2 AND2X2_5348 ( .A(round_ctr_rst), .B(\block[480] ), .Y(w_mem_inst__abc_21203_new_n6038_));
AND2X2 AND2X2_5349 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n6038_), .Y(w_mem_inst__abc_21203_new_n6039_));
AND2X2 AND2X2_535 ( .A(_abc_15497_new_n1808_), .B(digest_update), .Y(_abc_15497_new_n1809_));
AND2X2 AND2X2_5350 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_0__1_), .Y(w_mem_inst__abc_21203_new_n6042_));
AND2X2 AND2X2_5351 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_1__1_), .Y(w_mem_inst__abc_21203_new_n6043_));
AND2X2 AND2X2_5352 ( .A(round_ctr_rst), .B(\block[481] ), .Y(w_mem_inst__abc_21203_new_n6044_));
AND2X2 AND2X2_5353 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n6044_), .Y(w_mem_inst__abc_21203_new_n6045_));
AND2X2 AND2X2_5354 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_0__2_), .Y(w_mem_inst__abc_21203_new_n6048_));
AND2X2 AND2X2_5355 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_1__2_), .Y(w_mem_inst__abc_21203_new_n6049_));
AND2X2 AND2X2_5356 ( .A(round_ctr_rst), .B(\block[482] ), .Y(w_mem_inst__abc_21203_new_n6050_));
AND2X2 AND2X2_5357 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n6050_), .Y(w_mem_inst__abc_21203_new_n6051_));
AND2X2 AND2X2_5358 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_0__3_), .Y(w_mem_inst__abc_21203_new_n6054_));
AND2X2 AND2X2_5359 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_1__3_), .Y(w_mem_inst__abc_21203_new_n6055_));
AND2X2 AND2X2_536 ( .A(_abc_15497_new_n1809_), .B(_abc_15497_new_n1806_), .Y(_abc_15497_new_n1810_));
AND2X2 AND2X2_5360 ( .A(round_ctr_rst), .B(\block[483] ), .Y(w_mem_inst__abc_21203_new_n6056_));
AND2X2 AND2X2_5361 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n6056_), .Y(w_mem_inst__abc_21203_new_n6057_));
AND2X2 AND2X2_5362 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_0__4_), .Y(w_mem_inst__abc_21203_new_n6060_));
AND2X2 AND2X2_5363 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_1__4_), .Y(w_mem_inst__abc_21203_new_n6061_));
AND2X2 AND2X2_5364 ( .A(round_ctr_rst), .B(\block[484] ), .Y(w_mem_inst__abc_21203_new_n6062_));
AND2X2 AND2X2_5365 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n6062_), .Y(w_mem_inst__abc_21203_new_n6063_));
AND2X2 AND2X2_5366 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_0__5_), .Y(w_mem_inst__abc_21203_new_n6066_));
AND2X2 AND2X2_5367 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_1__5_), .Y(w_mem_inst__abc_21203_new_n6067_));
AND2X2 AND2X2_5368 ( .A(round_ctr_rst), .B(\block[485] ), .Y(w_mem_inst__abc_21203_new_n6068_));
AND2X2 AND2X2_5369 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n6068_), .Y(w_mem_inst__abc_21203_new_n6069_));
AND2X2 AND2X2_537 ( .A(_abc_15497_new_n1792_), .B(_abc_15497_new_n1805_), .Y(_abc_15497_new_n1812_));
AND2X2 AND2X2_5370 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_0__6_), .Y(w_mem_inst__abc_21203_new_n6072_));
AND2X2 AND2X2_5371 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_1__6_), .Y(w_mem_inst__abc_21203_new_n6073_));
AND2X2 AND2X2_5372 ( .A(round_ctr_rst), .B(\block[486] ), .Y(w_mem_inst__abc_21203_new_n6074_));
AND2X2 AND2X2_5373 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n6074_), .Y(w_mem_inst__abc_21203_new_n6075_));
AND2X2 AND2X2_5374 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_0__7_), .Y(w_mem_inst__abc_21203_new_n6078_));
AND2X2 AND2X2_5375 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_1__7_), .Y(w_mem_inst__abc_21203_new_n6079_));
AND2X2 AND2X2_5376 ( .A(round_ctr_rst), .B(\block[487] ), .Y(w_mem_inst__abc_21203_new_n6080_));
AND2X2 AND2X2_5377 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n6080_), .Y(w_mem_inst__abc_21203_new_n6081_));
AND2X2 AND2X2_5378 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_0__8_), .Y(w_mem_inst__abc_21203_new_n6084_));
AND2X2 AND2X2_5379 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_1__8_), .Y(w_mem_inst__abc_21203_new_n6085_));
AND2X2 AND2X2_538 ( .A(_abc_15497_new_n1786_), .B(_abc_15497_new_n1812_), .Y(_abc_15497_new_n1813_));
AND2X2 AND2X2_5380 ( .A(round_ctr_rst), .B(\block[488] ), .Y(w_mem_inst__abc_21203_new_n6086_));
AND2X2 AND2X2_5381 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n6086_), .Y(w_mem_inst__abc_21203_new_n6087_));
AND2X2 AND2X2_5382 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_0__9_), .Y(w_mem_inst__abc_21203_new_n6090_));
AND2X2 AND2X2_5383 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_1__9_), .Y(w_mem_inst__abc_21203_new_n6091_));
AND2X2 AND2X2_5384 ( .A(round_ctr_rst), .B(\block[489] ), .Y(w_mem_inst__abc_21203_new_n6092_));
AND2X2 AND2X2_5385 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n6092_), .Y(w_mem_inst__abc_21203_new_n6093_));
AND2X2 AND2X2_5386 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_0__10_), .Y(w_mem_inst__abc_21203_new_n6096_));
AND2X2 AND2X2_5387 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_1__10_), .Y(w_mem_inst__abc_21203_new_n6097_));
AND2X2 AND2X2_5388 ( .A(round_ctr_rst), .B(\block[490] ), .Y(w_mem_inst__abc_21203_new_n6098_));
AND2X2 AND2X2_5389 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n6098_), .Y(w_mem_inst__abc_21203_new_n6099_));
AND2X2 AND2X2_539 ( .A(_abc_15497_new_n1758_), .B(_abc_15497_new_n1813_), .Y(_abc_15497_new_n1814_));
AND2X2 AND2X2_5390 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_0__11_), .Y(w_mem_inst__abc_21203_new_n6102_));
AND2X2 AND2X2_5391 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_1__11_), .Y(w_mem_inst__abc_21203_new_n6103_));
AND2X2 AND2X2_5392 ( .A(round_ctr_rst), .B(\block[491] ), .Y(w_mem_inst__abc_21203_new_n6104_));
AND2X2 AND2X2_5393 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n6104_), .Y(w_mem_inst__abc_21203_new_n6105_));
AND2X2 AND2X2_5394 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_0__12_), .Y(w_mem_inst__abc_21203_new_n6108_));
AND2X2 AND2X2_5395 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_1__12_), .Y(w_mem_inst__abc_21203_new_n6109_));
AND2X2 AND2X2_5396 ( .A(round_ctr_rst), .B(\block[492] ), .Y(w_mem_inst__abc_21203_new_n6110_));
AND2X2 AND2X2_5397 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n6110_), .Y(w_mem_inst__abc_21203_new_n6111_));
AND2X2 AND2X2_5398 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_0__13_), .Y(w_mem_inst__abc_21203_new_n6114_));
AND2X2 AND2X2_5399 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_1__13_), .Y(w_mem_inst__abc_21203_new_n6115_));
AND2X2 AND2X2_54 ( .A(c_reg_7_), .B(\digest[71] ), .Y(_abc_15497_new_n801_));
AND2X2 AND2X2_540 ( .A(_abc_15497_new_n1785_), .B(_abc_15497_new_n1812_), .Y(_abc_15497_new_n1815_));
AND2X2 AND2X2_5400 ( .A(round_ctr_rst), .B(\block[493] ), .Y(w_mem_inst__abc_21203_new_n6116_));
AND2X2 AND2X2_5401 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n6116_), .Y(w_mem_inst__abc_21203_new_n6117_));
AND2X2 AND2X2_5402 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_0__14_), .Y(w_mem_inst__abc_21203_new_n6120_));
AND2X2 AND2X2_5403 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_1__14_), .Y(w_mem_inst__abc_21203_new_n6121_));
AND2X2 AND2X2_5404 ( .A(round_ctr_rst), .B(\block[494] ), .Y(w_mem_inst__abc_21203_new_n6122_));
AND2X2 AND2X2_5405 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n6122_), .Y(w_mem_inst__abc_21203_new_n6123_));
AND2X2 AND2X2_5406 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_0__15_), .Y(w_mem_inst__abc_21203_new_n6126_));
AND2X2 AND2X2_5407 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_1__15_), .Y(w_mem_inst__abc_21203_new_n6127_));
AND2X2 AND2X2_5408 ( .A(round_ctr_rst), .B(\block[495] ), .Y(w_mem_inst__abc_21203_new_n6128_));
AND2X2 AND2X2_5409 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n6128_), .Y(w_mem_inst__abc_21203_new_n6129_));
AND2X2 AND2X2_541 ( .A(_abc_15497_new_n1802_), .B(_abc_15497_new_n1790_), .Y(_abc_15497_new_n1816_));
AND2X2 AND2X2_5410 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_0__16_), .Y(w_mem_inst__abc_21203_new_n6132_));
AND2X2 AND2X2_5411 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_1__16_), .Y(w_mem_inst__abc_21203_new_n6133_));
AND2X2 AND2X2_5412 ( .A(round_ctr_rst), .B(\block[496] ), .Y(w_mem_inst__abc_21203_new_n6134_));
AND2X2 AND2X2_5413 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n6134_), .Y(w_mem_inst__abc_21203_new_n6135_));
AND2X2 AND2X2_5414 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_0__17_), .Y(w_mem_inst__abc_21203_new_n6138_));
AND2X2 AND2X2_5415 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_1__17_), .Y(w_mem_inst__abc_21203_new_n6139_));
AND2X2 AND2X2_5416 ( .A(round_ctr_rst), .B(\block[497] ), .Y(w_mem_inst__abc_21203_new_n6140_));
AND2X2 AND2X2_5417 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n6140_), .Y(w_mem_inst__abc_21203_new_n6141_));
AND2X2 AND2X2_5418 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_0__18_), .Y(w_mem_inst__abc_21203_new_n6144_));
AND2X2 AND2X2_5419 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_1__18_), .Y(w_mem_inst__abc_21203_new_n6145_));
AND2X2 AND2X2_542 ( .A(\digest[52] ), .B(d_reg_20_), .Y(_abc_15497_new_n1821_));
AND2X2 AND2X2_5420 ( .A(round_ctr_rst), .B(\block[498] ), .Y(w_mem_inst__abc_21203_new_n6146_));
AND2X2 AND2X2_5421 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n6146_), .Y(w_mem_inst__abc_21203_new_n6147_));
AND2X2 AND2X2_5422 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_0__19_), .Y(w_mem_inst__abc_21203_new_n6150_));
AND2X2 AND2X2_5423 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_1__19_), .Y(w_mem_inst__abc_21203_new_n6151_));
AND2X2 AND2X2_5424 ( .A(round_ctr_rst), .B(\block[499] ), .Y(w_mem_inst__abc_21203_new_n6152_));
AND2X2 AND2X2_5425 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n6152_), .Y(w_mem_inst__abc_21203_new_n6153_));
AND2X2 AND2X2_5426 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_0__20_), .Y(w_mem_inst__abc_21203_new_n6156_));
AND2X2 AND2X2_5427 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_1__20_), .Y(w_mem_inst__abc_21203_new_n6157_));
AND2X2 AND2X2_5428 ( .A(round_ctr_rst), .B(\block[500] ), .Y(w_mem_inst__abc_21203_new_n6158_));
AND2X2 AND2X2_5429 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n6158_), .Y(w_mem_inst__abc_21203_new_n6159_));
AND2X2 AND2X2_543 ( .A(_abc_15497_new_n1822_), .B(_abc_15497_new_n1820_), .Y(_abc_15497_new_n1823_));
AND2X2 AND2X2_5430 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_0__21_), .Y(w_mem_inst__abc_21203_new_n6162_));
AND2X2 AND2X2_5431 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_1__21_), .Y(w_mem_inst__abc_21203_new_n6163_));
AND2X2 AND2X2_5432 ( .A(round_ctr_rst), .B(\block[501] ), .Y(w_mem_inst__abc_21203_new_n6164_));
AND2X2 AND2X2_5433 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n6164_), .Y(w_mem_inst__abc_21203_new_n6165_));
AND2X2 AND2X2_5434 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_0__22_), .Y(w_mem_inst__abc_21203_new_n6168_));
AND2X2 AND2X2_5435 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_1__22_), .Y(w_mem_inst__abc_21203_new_n6169_));
AND2X2 AND2X2_5436 ( .A(round_ctr_rst), .B(\block[502] ), .Y(w_mem_inst__abc_21203_new_n6170_));
AND2X2 AND2X2_5437 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n6170_), .Y(w_mem_inst__abc_21203_new_n6171_));
AND2X2 AND2X2_5438 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_0__23_), .Y(w_mem_inst__abc_21203_new_n6174_));
AND2X2 AND2X2_5439 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_1__23_), .Y(w_mem_inst__abc_21203_new_n6175_));
AND2X2 AND2X2_544 ( .A(_abc_15497_new_n1819_), .B(_abc_15497_new_n1823_), .Y(_abc_15497_new_n1825_));
AND2X2 AND2X2_5440 ( .A(round_ctr_rst), .B(\block[503] ), .Y(w_mem_inst__abc_21203_new_n6176_));
AND2X2 AND2X2_5441 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n6176_), .Y(w_mem_inst__abc_21203_new_n6177_));
AND2X2 AND2X2_5442 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_0__24_), .Y(w_mem_inst__abc_21203_new_n6180_));
AND2X2 AND2X2_5443 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_1__24_), .Y(w_mem_inst__abc_21203_new_n6181_));
AND2X2 AND2X2_5444 ( .A(round_ctr_rst), .B(\block[504] ), .Y(w_mem_inst__abc_21203_new_n6182_));
AND2X2 AND2X2_5445 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n6182_), .Y(w_mem_inst__abc_21203_new_n6183_));
AND2X2 AND2X2_5446 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_0__25_), .Y(w_mem_inst__abc_21203_new_n6186_));
AND2X2 AND2X2_5447 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_1__25_), .Y(w_mem_inst__abc_21203_new_n6187_));
AND2X2 AND2X2_5448 ( .A(round_ctr_rst), .B(\block[505] ), .Y(w_mem_inst__abc_21203_new_n6188_));
AND2X2 AND2X2_5449 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n6188_), .Y(w_mem_inst__abc_21203_new_n6189_));
AND2X2 AND2X2_545 ( .A(_abc_15497_new_n1826_), .B(_abc_15497_new_n1824_), .Y(_abc_15497_new_n1827_));
AND2X2 AND2X2_5450 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_0__26_), .Y(w_mem_inst__abc_21203_new_n6192_));
AND2X2 AND2X2_5451 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_1__26_), .Y(w_mem_inst__abc_21203_new_n6193_));
AND2X2 AND2X2_5452 ( .A(round_ctr_rst), .B(\block[506] ), .Y(w_mem_inst__abc_21203_new_n6194_));
AND2X2 AND2X2_5453 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n6194_), .Y(w_mem_inst__abc_21203_new_n6195_));
AND2X2 AND2X2_5454 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_0__27_), .Y(w_mem_inst__abc_21203_new_n6198_));
AND2X2 AND2X2_5455 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_1__27_), .Y(w_mem_inst__abc_21203_new_n6199_));
AND2X2 AND2X2_5456 ( .A(round_ctr_rst), .B(\block[507] ), .Y(w_mem_inst__abc_21203_new_n6200_));
AND2X2 AND2X2_5457 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n6200_), .Y(w_mem_inst__abc_21203_new_n6201_));
AND2X2 AND2X2_5458 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_0__28_), .Y(w_mem_inst__abc_21203_new_n6204_));
AND2X2 AND2X2_5459 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_1__28_), .Y(w_mem_inst__abc_21203_new_n6205_));
AND2X2 AND2X2_546 ( .A(_abc_15497_new_n1827_), .B(digest_update), .Y(_abc_15497_new_n1828_));
AND2X2 AND2X2_5460 ( .A(round_ctr_rst), .B(\block[508] ), .Y(w_mem_inst__abc_21203_new_n6206_));
AND2X2 AND2X2_5461 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n6206_), .Y(w_mem_inst__abc_21203_new_n6207_));
AND2X2 AND2X2_5462 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_0__29_), .Y(w_mem_inst__abc_21203_new_n6210_));
AND2X2 AND2X2_5463 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_1__29_), .Y(w_mem_inst__abc_21203_new_n6211_));
AND2X2 AND2X2_5464 ( .A(round_ctr_rst), .B(\block[509] ), .Y(w_mem_inst__abc_21203_new_n6212_));
AND2X2 AND2X2_5465 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n6212_), .Y(w_mem_inst__abc_21203_new_n6213_));
AND2X2 AND2X2_5466 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_0__30_), .Y(w_mem_inst__abc_21203_new_n6216_));
AND2X2 AND2X2_5467 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_1__30_), .Y(w_mem_inst__abc_21203_new_n6217_));
AND2X2 AND2X2_5468 ( .A(round_ctr_rst), .B(\block[510] ), .Y(w_mem_inst__abc_21203_new_n6218_));
AND2X2 AND2X2_5469 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n6218_), .Y(w_mem_inst__abc_21203_new_n6219_));
AND2X2 AND2X2_547 ( .A(_abc_15497_new_n1829_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n1830_));
AND2X2 AND2X2_5470 ( .A(w_mem_inst__abc_21203_new_n3155_), .B(w_mem_inst_w_mem_0__31_), .Y(w_mem_inst__abc_21203_new_n6222_));
AND2X2 AND2X2_5471 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst_w_mem_1__31_), .Y(w_mem_inst__abc_21203_new_n6223_));
AND2X2 AND2X2_5472 ( .A(round_ctr_rst), .B(\block[511] ), .Y(w_mem_inst__abc_21203_new_n6224_));
AND2X2 AND2X2_5473 ( .A(w_mem_inst__abc_21203_new_n3154_), .B(w_mem_inst__abc_21203_new_n6224_), .Y(w_mem_inst__abc_21203_new_n6225_));
AND2X2 AND2X2_5474 ( .A(w_mem_inst__abc_21203_new_n6229_), .B(w_mem_inst__abc_21203_new_n3152_), .Y(w_mem_inst__abc_21203_new_n6230_));
AND2X2 AND2X2_5475 ( .A(w_mem_inst__abc_21203_new_n6231_), .B(w_mem_inst__abc_21203_new_n6228_), .Y(w_mem_inst__0w_ctr_reg_6_0__0_));
AND2X2 AND2X2_5476 ( .A(w_mem_inst__abc_21203_new_n6230_), .B(w_mem_inst_w_ctr_reg_1_), .Y(w_mem_inst__abc_21203_new_n6233_));
AND2X2 AND2X2_5477 ( .A(w_mem_inst__abc_21203_new_n6234_), .B(round_ctr_inc), .Y(w_mem_inst__abc_21203_new_n6235_));
AND2X2 AND2X2_5478 ( .A(w_mem_inst__abc_21203_new_n6237_), .B(w_mem_inst_w_ctr_reg_2_), .Y(w_mem_inst__abc_21203_new_n6238_));
AND2X2 AND2X2_5479 ( .A(w_mem_inst__abc_21203_new_n1616_), .B(round_ctr_inc), .Y(w_mem_inst__abc_21203_new_n6239_));
AND2X2 AND2X2_548 ( .A(_abc_15497_new_n1826_), .B(_abc_15497_new_n1822_), .Y(_abc_15497_new_n1832_));
AND2X2 AND2X2_5480 ( .A(w_mem_inst__abc_21203_new_n1616_), .B(w_mem_inst_w_ctr_reg_2_), .Y(w_mem_inst__abc_21203_new_n6241_));
AND2X2 AND2X2_5481 ( .A(w_mem_inst__abc_21203_new_n6241_), .B(round_ctr_inc), .Y(w_mem_inst__abc_21203_new_n6242_));
AND2X2 AND2X2_5482 ( .A(w_mem_inst__abc_21203_new_n6240_), .B(w_mem_inst__abc_21203_new_n6243_), .Y(w_mem_inst__0w_ctr_reg_6_0__2_));
AND2X2 AND2X2_5483 ( .A(w_mem_inst__abc_21203_new_n6237_), .B(w_mem_inst_w_ctr_reg_3_), .Y(w_mem_inst__abc_21203_new_n6245_));
AND2X2 AND2X2_5484 ( .A(w_mem_inst__abc_21203_new_n1624_), .B(round_ctr_inc), .Y(w_mem_inst__abc_21203_new_n6247_));
AND2X2 AND2X2_5485 ( .A(w_mem_inst__abc_21203_new_n6246_), .B(w_mem_inst__abc_21203_new_n6248_), .Y(w_mem_inst__0w_ctr_reg_6_0__3_));
AND2X2 AND2X2_5486 ( .A(w_mem_inst__abc_21203_new_n6237_), .B(w_mem_inst_w_ctr_reg_4_), .Y(w_mem_inst__abc_21203_new_n6250_));
AND2X2 AND2X2_5487 ( .A(w_mem_inst__abc_21203_new_n6247_), .B(w_mem_inst_w_ctr_reg_4_), .Y(w_mem_inst__abc_21203_new_n6252_));
AND2X2 AND2X2_5488 ( .A(w_mem_inst__abc_21203_new_n6253_), .B(w_mem_inst__abc_21203_new_n6251_), .Y(w_mem_inst__0w_ctr_reg_6_0__4_));
AND2X2 AND2X2_5489 ( .A(w_mem_inst__abc_21203_new_n6237_), .B(w_mem_inst_w_ctr_reg_5_), .Y(w_mem_inst__abc_21203_new_n6255_));
AND2X2 AND2X2_549 ( .A(\digest[53] ), .B(d_reg_21_), .Y(_abc_15497_new_n1835_));
AND2X2 AND2X2_5490 ( .A(w_mem_inst__abc_21203_new_n6252_), .B(w_mem_inst_w_ctr_reg_5_), .Y(w_mem_inst__abc_21203_new_n6257_));
AND2X2 AND2X2_5491 ( .A(w_mem_inst__abc_21203_new_n6258_), .B(w_mem_inst__abc_21203_new_n6256_), .Y(w_mem_inst__0w_ctr_reg_6_0__5_));
AND2X2 AND2X2_5492 ( .A(w_mem_inst__abc_21203_new_n6237_), .B(w_mem_inst_w_ctr_reg_6_), .Y(w_mem_inst__abc_21203_new_n6260_));
AND2X2 AND2X2_5493 ( .A(w_mem_inst__abc_21203_new_n6257_), .B(w_mem_inst_w_ctr_reg_6_), .Y(w_mem_inst__abc_21203_new_n6262_));
AND2X2 AND2X2_5494 ( .A(w_mem_inst__abc_21203_new_n6263_), .B(w_mem_inst__abc_21203_new_n6261_), .Y(w_mem_inst__0w_ctr_reg_6_0__6_));
AND2X2 AND2X2_55 ( .A(c_reg_6_), .B(\digest[70] ), .Y(_abc_15497_new_n803_));
AND2X2 AND2X2_550 ( .A(_abc_15497_new_n1836_), .B(_abc_15497_new_n1834_), .Y(_abc_15497_new_n1837_));
AND2X2 AND2X2_551 ( .A(_abc_15497_new_n1838_), .B(_abc_15497_new_n1840_), .Y(_abc_15497_new_n1841_));
AND2X2 AND2X2_552 ( .A(_abc_15497_new_n1841_), .B(digest_update), .Y(_abc_15497_new_n1842_));
AND2X2 AND2X2_553 ( .A(_abc_15497_new_n1843_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n1844_));
AND2X2 AND2X2_554 ( .A(_abc_15497_new_n701_), .B(\digest[54] ), .Y(_abc_15497_new_n1846_));
AND2X2 AND2X2_555 ( .A(\digest[54] ), .B(d_reg_22_), .Y(_abc_15497_new_n1848_));
AND2X2 AND2X2_556 ( .A(_abc_15497_new_n1849_), .B(_abc_15497_new_n1847_), .Y(_abc_15497_new_n1850_));
AND2X2 AND2X2_557 ( .A(_abc_15497_new_n1822_), .B(_abc_15497_new_n1836_), .Y(_abc_15497_new_n1852_));
AND2X2 AND2X2_558 ( .A(_abc_15497_new_n1826_), .B(_abc_15497_new_n1852_), .Y(_abc_15497_new_n1853_));
AND2X2 AND2X2_559 ( .A(_abc_15497_new_n1855_), .B(_abc_15497_new_n1850_), .Y(_abc_15497_new_n1857_));
AND2X2 AND2X2_56 ( .A(_abc_15497_new_n802_), .B(_abc_15497_new_n803_), .Y(_abc_15497_new_n804_));
AND2X2 AND2X2_560 ( .A(_abc_15497_new_n1858_), .B(_abc_15497_new_n1856_), .Y(_abc_15497_new_n1859_));
AND2X2 AND2X2_561 ( .A(_abc_15497_new_n1859_), .B(digest_update), .Y(_abc_15497_new_n1860_));
AND2X2 AND2X2_562 ( .A(_abc_15497_new_n701_), .B(\digest[55] ), .Y(_abc_15497_new_n1862_));
AND2X2 AND2X2_563 ( .A(\digest[55] ), .B(d_reg_23_), .Y(_abc_15497_new_n1865_));
AND2X2 AND2X2_564 ( .A(_abc_15497_new_n1866_), .B(_abc_15497_new_n1864_), .Y(_abc_15497_new_n1867_));
AND2X2 AND2X2_565 ( .A(_abc_15497_new_n1871_), .B(_abc_15497_new_n1868_), .Y(_abc_15497_new_n1872_));
AND2X2 AND2X2_566 ( .A(_abc_15497_new_n1872_), .B(digest_update), .Y(_abc_15497_new_n1873_));
AND2X2 AND2X2_567 ( .A(_abc_15497_new_n701_), .B(\digest[56] ), .Y(_abc_15497_new_n1875_));
AND2X2 AND2X2_568 ( .A(_abc_15497_new_n1864_), .B(_abc_15497_new_n1848_), .Y(_abc_15497_new_n1876_));
AND2X2 AND2X2_569 ( .A(_abc_15497_new_n1850_), .B(_abc_15497_new_n1867_), .Y(_abc_15497_new_n1880_));
AND2X2 AND2X2_57 ( .A(_abc_15497_new_n806_), .B(_abc_15497_new_n802_), .Y(_abc_15497_new_n807_));
AND2X2 AND2X2_570 ( .A(_abc_15497_new_n1882_), .B(_abc_15497_new_n1878_), .Y(_abc_15497_new_n1883_));
AND2X2 AND2X2_571 ( .A(_abc_15497_new_n1823_), .B(_abc_15497_new_n1837_), .Y(_abc_15497_new_n1885_));
AND2X2 AND2X2_572 ( .A(_abc_15497_new_n1885_), .B(_abc_15497_new_n1880_), .Y(_abc_15497_new_n1886_));
AND2X2 AND2X2_573 ( .A(_abc_15497_new_n1819_), .B(_abc_15497_new_n1886_), .Y(_abc_15497_new_n1887_));
AND2X2 AND2X2_574 ( .A(\digest[56] ), .B(d_reg_24_), .Y(_abc_15497_new_n1890_));
AND2X2 AND2X2_575 ( .A(_abc_15497_new_n1891_), .B(_abc_15497_new_n1889_), .Y(_abc_15497_new_n1892_));
AND2X2 AND2X2_576 ( .A(_abc_15497_new_n1888_), .B(_abc_15497_new_n1892_), .Y(_abc_15497_new_n1894_));
AND2X2 AND2X2_577 ( .A(_abc_15497_new_n1895_), .B(_abc_15497_new_n1893_), .Y(_abc_15497_new_n1896_));
AND2X2 AND2X2_578 ( .A(_abc_15497_new_n1896_), .B(digest_update), .Y(_abc_15497_new_n1897_));
AND2X2 AND2X2_579 ( .A(_abc_15497_new_n701_), .B(\digest[57] ), .Y(_abc_15497_new_n1899_));
AND2X2 AND2X2_58 ( .A(_abc_15497_new_n808_), .B(_abc_15497_new_n809_), .Y(_abc_15497_new_n810_));
AND2X2 AND2X2_580 ( .A(\digest[57] ), .B(d_reg_25_), .Y(_abc_15497_new_n1901_));
AND2X2 AND2X2_581 ( .A(_abc_15497_new_n1902_), .B(_abc_15497_new_n1900_), .Y(_abc_15497_new_n1903_));
AND2X2 AND2X2_582 ( .A(_abc_15497_new_n1892_), .B(_abc_15497_new_n1903_), .Y(_abc_15497_new_n1906_));
AND2X2 AND2X2_583 ( .A(_abc_15497_new_n1888_), .B(_abc_15497_new_n1906_), .Y(_abc_15497_new_n1907_));
AND2X2 AND2X2_584 ( .A(_abc_15497_new_n1903_), .B(_abc_15497_new_n1890_), .Y(_abc_15497_new_n1909_));
AND2X2 AND2X2_585 ( .A(_abc_15497_new_n1910_), .B(digest_update), .Y(_abc_15497_new_n1911_));
AND2X2 AND2X2_586 ( .A(_abc_15497_new_n1908_), .B(_abc_15497_new_n1911_), .Y(_abc_15497_new_n1912_));
AND2X2 AND2X2_587 ( .A(_abc_15497_new_n1912_), .B(_abc_15497_new_n1905_), .Y(_abc_15497_new_n1913_));
AND2X2 AND2X2_588 ( .A(_abc_15497_new_n701_), .B(\digest[58] ), .Y(_abc_15497_new_n1915_));
AND2X2 AND2X2_589 ( .A(_abc_15497_new_n1910_), .B(_abc_15497_new_n1902_), .Y(_abc_15497_new_n1916_));
AND2X2 AND2X2_59 ( .A(_abc_15497_new_n807_), .B(_abc_15497_new_n810_), .Y(_abc_15497_new_n811_));
AND2X2 AND2X2_590 ( .A(_abc_15497_new_n1908_), .B(_abc_15497_new_n1916_), .Y(_abc_15497_new_n1917_));
AND2X2 AND2X2_591 ( .A(\digest[58] ), .B(d_reg_26_), .Y(_abc_15497_new_n1920_));
AND2X2 AND2X2_592 ( .A(_abc_15497_new_n1921_), .B(_abc_15497_new_n1919_), .Y(_abc_15497_new_n1922_));
AND2X2 AND2X2_593 ( .A(_abc_15497_new_n1918_), .B(_abc_15497_new_n1922_), .Y(_abc_15497_new_n1924_));
AND2X2 AND2X2_594 ( .A(_abc_15497_new_n1925_), .B(_abc_15497_new_n1923_), .Y(_abc_15497_new_n1926_));
AND2X2 AND2X2_595 ( .A(_abc_15497_new_n1926_), .B(digest_update), .Y(_abc_15497_new_n1927_));
AND2X2 AND2X2_596 ( .A(_abc_15497_new_n701_), .B(\digest[59] ), .Y(_abc_15497_new_n1929_));
AND2X2 AND2X2_597 ( .A(\digest[59] ), .B(d_reg_27_), .Y(_abc_15497_new_n1931_));
AND2X2 AND2X2_598 ( .A(_abc_15497_new_n1932_), .B(_abc_15497_new_n1930_), .Y(_abc_15497_new_n1933_));
AND2X2 AND2X2_599 ( .A(_abc_15497_new_n1922_), .B(_abc_15497_new_n1933_), .Y(_abc_15497_new_n1936_));
AND2X2 AND2X2_6 ( .A(c_reg_22_), .B(\digest[86] ), .Y(_abc_15497_new_n707_));
AND2X2 AND2X2_60 ( .A(c_reg_5_), .B(\digest[69] ), .Y(_abc_15497_new_n812_));
AND2X2 AND2X2_600 ( .A(_abc_15497_new_n1933_), .B(_abc_15497_new_n1920_), .Y(_abc_15497_new_n1939_));
AND2X2 AND2X2_601 ( .A(_abc_15497_new_n1940_), .B(digest_update), .Y(_abc_15497_new_n1941_));
AND2X2 AND2X2_602 ( .A(_abc_15497_new_n1938_), .B(_abc_15497_new_n1941_), .Y(_abc_15497_new_n1942_));
AND2X2 AND2X2_603 ( .A(_abc_15497_new_n1935_), .B(_abc_15497_new_n1942_), .Y(_abc_15497_new_n1943_));
AND2X2 AND2X2_604 ( .A(_abc_15497_new_n1906_), .B(_abc_15497_new_n1936_), .Y(_abc_15497_new_n1945_));
AND2X2 AND2X2_605 ( .A(_abc_15497_new_n1888_), .B(_abc_15497_new_n1945_), .Y(_abc_15497_new_n1946_));
AND2X2 AND2X2_606 ( .A(_abc_15497_new_n1940_), .B(_abc_15497_new_n1932_), .Y(_abc_15497_new_n1947_));
AND2X2 AND2X2_607 ( .A(_abc_15497_new_n1948_), .B(_abc_15497_new_n1947_), .Y(_abc_15497_new_n1949_));
AND2X2 AND2X2_608 ( .A(\digest[60] ), .B(d_reg_28_), .Y(_abc_15497_new_n1953_));
AND2X2 AND2X2_609 ( .A(_abc_15497_new_n1954_), .B(_abc_15497_new_n1952_), .Y(_abc_15497_new_n1955_));
AND2X2 AND2X2_61 ( .A(c_reg_4_), .B(\digest[68] ), .Y(_abc_15497_new_n814_));
AND2X2 AND2X2_610 ( .A(_abc_15497_new_n1951_), .B(_abc_15497_new_n1955_), .Y(_abc_15497_new_n1957_));
AND2X2 AND2X2_611 ( .A(_abc_15497_new_n1958_), .B(_abc_15497_new_n1956_), .Y(_abc_15497_new_n1959_));
AND2X2 AND2X2_612 ( .A(_abc_15497_new_n1959_), .B(digest_update), .Y(_abc_15497_new_n1960_));
AND2X2 AND2X2_613 ( .A(_abc_15497_new_n1961_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n1962_));
AND2X2 AND2X2_614 ( .A(_abc_15497_new_n701_), .B(\digest[61] ), .Y(_abc_15497_new_n1964_));
AND2X2 AND2X2_615 ( .A(_abc_15497_new_n1958_), .B(_abc_15497_new_n1954_), .Y(_abc_15497_new_n1965_));
AND2X2 AND2X2_616 ( .A(\digest[61] ), .B(d_reg_29_), .Y(_abc_15497_new_n1968_));
AND2X2 AND2X2_617 ( .A(_abc_15497_new_n1969_), .B(_abc_15497_new_n1967_), .Y(_abc_15497_new_n1970_));
AND2X2 AND2X2_618 ( .A(_abc_15497_new_n1973_), .B(digest_update), .Y(_abc_15497_new_n1974_));
AND2X2 AND2X2_619 ( .A(_abc_15497_new_n1974_), .B(_abc_15497_new_n1971_), .Y(_abc_15497_new_n1975_));
AND2X2 AND2X2_62 ( .A(c_reg_3_), .B(\digest[67] ), .Y(_abc_15497_new_n815_));
AND2X2 AND2X2_620 ( .A(_abc_15497_new_n701_), .B(\digest[62] ), .Y(_abc_15497_new_n1977_));
AND2X2 AND2X2_621 ( .A(\digest[62] ), .B(d_reg_30_), .Y(_abc_15497_new_n1978_));
AND2X2 AND2X2_622 ( .A(_abc_15497_new_n1979_), .B(_abc_15497_new_n1980_), .Y(_abc_15497_new_n1981_));
AND2X2 AND2X2_623 ( .A(_abc_15497_new_n1970_), .B(_abc_15497_new_n1953_), .Y(_abc_15497_new_n1982_));
AND2X2 AND2X2_624 ( .A(_abc_15497_new_n1955_), .B(_abc_15497_new_n1970_), .Y(_abc_15497_new_n1984_));
AND2X2 AND2X2_625 ( .A(_abc_15497_new_n1951_), .B(_abc_15497_new_n1984_), .Y(_abc_15497_new_n1985_));
AND2X2 AND2X2_626 ( .A(_abc_15497_new_n1986_), .B(_abc_15497_new_n1981_), .Y(_abc_15497_new_n1987_));
AND2X2 AND2X2_627 ( .A(_abc_15497_new_n1989_), .B(digest_update), .Y(_abc_15497_new_n1990_));
AND2X2 AND2X2_628 ( .A(_abc_15497_new_n1990_), .B(_abc_15497_new_n1988_), .Y(_abc_15497_new_n1991_));
AND2X2 AND2X2_629 ( .A(_abc_15497_new_n701_), .B(\digest[63] ), .Y(_abc_15497_new_n1993_));
AND2X2 AND2X2_63 ( .A(c_reg_2_), .B(\digest[66] ), .Y(_abc_15497_new_n817_));
AND2X2 AND2X2_630 ( .A(\digest[63] ), .B(d_reg_31_), .Y(_abc_15497_new_n1997_));
AND2X2 AND2X2_631 ( .A(_abc_15497_new_n1998_), .B(_abc_15497_new_n1996_), .Y(_abc_15497_new_n1999_));
AND2X2 AND2X2_632 ( .A(_abc_15497_new_n2002_), .B(digest_update), .Y(_abc_15497_new_n2003_));
AND2X2 AND2X2_633 ( .A(_abc_15497_new_n2003_), .B(_abc_15497_new_n2001_), .Y(_abc_15497_new_n2004_));
AND2X2 AND2X2_634 ( .A(_abc_15497_new_n2006_), .B(ready), .Y(round_ctr_rst));
AND2X2 AND2X2_635 ( .A(_abc_15497_new_n2009_), .B(_abc_15497_new_n2008_), .Y(_abc_15497_new_n2010_));
AND2X2 AND2X2_636 ( .A(_abc_15497_new_n2010_), .B(e_reg_0_), .Y(_abc_15497_new_n2011_));
AND2X2 AND2X2_637 ( .A(_abc_15497_new_n700_), .B(\digest[0] ), .Y(_abc_15497_new_n2012_));
AND2X2 AND2X2_638 ( .A(round_ctr_rst), .B(_abc_15497_new_n2008_), .Y(_abc_15497_new_n2013_));
AND2X2 AND2X2_639 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n2012_), .Y(_abc_15497_new_n2014_));
AND2X2 AND2X2_64 ( .A(c_reg_1_), .B(\digest[65] ), .Y(_abc_15497_new_n818_));
AND2X2 AND2X2_640 ( .A(d_reg_0_), .B(round_ctr_inc), .Y(_abc_15497_new_n2015_));
AND2X2 AND2X2_641 ( .A(_abc_15497_new_n2010_), .B(e_reg_1_), .Y(_abc_15497_new_n2018_));
AND2X2 AND2X2_642 ( .A(_abc_15497_new_n700_), .B(\digest[1] ), .Y(_abc_15497_new_n2019_));
AND2X2 AND2X2_643 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n2019_), .Y(_abc_15497_new_n2020_));
AND2X2 AND2X2_644 ( .A(d_reg_1_), .B(round_ctr_inc), .Y(_abc_15497_new_n2021_));
AND2X2 AND2X2_645 ( .A(_abc_15497_new_n2010_), .B(e_reg_2_), .Y(_abc_15497_new_n2024_));
AND2X2 AND2X2_646 ( .A(_abc_15497_new_n700_), .B(\digest[2] ), .Y(_abc_15497_new_n2025_));
AND2X2 AND2X2_647 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n2025_), .Y(_abc_15497_new_n2026_));
AND2X2 AND2X2_648 ( .A(d_reg_2_), .B(round_ctr_inc), .Y(_abc_15497_new_n2027_));
AND2X2 AND2X2_649 ( .A(_abc_15497_new_n2010_), .B(e_reg_3_), .Y(_abc_15497_new_n2030_));
AND2X2 AND2X2_65 ( .A(c_reg_0_), .B(\digest[64] ), .Y(_abc_15497_new_n819_));
AND2X2 AND2X2_650 ( .A(_abc_15497_new_n700_), .B(\digest[3] ), .Y(_abc_15497_new_n2031_));
AND2X2 AND2X2_651 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n2031_), .Y(_abc_15497_new_n2032_));
AND2X2 AND2X2_652 ( .A(d_reg_3_), .B(round_ctr_inc), .Y(_abc_15497_new_n2033_));
AND2X2 AND2X2_653 ( .A(_abc_15497_new_n2010_), .B(e_reg_4_), .Y(_abc_15497_new_n2036_));
AND2X2 AND2X2_654 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n1070_), .Y(_abc_15497_new_n2037_));
AND2X2 AND2X2_655 ( .A(d_reg_4_), .B(round_ctr_inc), .Y(_abc_15497_new_n2038_));
AND2X2 AND2X2_656 ( .A(_abc_15497_new_n2010_), .B(e_reg_5_), .Y(_abc_15497_new_n2041_));
AND2X2 AND2X2_657 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n1085_), .Y(_abc_15497_new_n2042_));
AND2X2 AND2X2_658 ( .A(d_reg_5_), .B(round_ctr_inc), .Y(_abc_15497_new_n2043_));
AND2X2 AND2X2_659 ( .A(_abc_15497_new_n2010_), .B(e_reg_6_), .Y(_abc_15497_new_n2046_));
AND2X2 AND2X2_66 ( .A(_abc_15497_new_n820_), .B(_abc_15497_new_n821_), .Y(_abc_15497_new_n822_));
AND2X2 AND2X2_660 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n1100_), .Y(_abc_15497_new_n2047_));
AND2X2 AND2X2_661 ( .A(d_reg_6_), .B(round_ctr_inc), .Y(_abc_15497_new_n2048_));
AND2X2 AND2X2_662 ( .A(_abc_15497_new_n2010_), .B(e_reg_7_), .Y(_abc_15497_new_n2051_));
AND2X2 AND2X2_663 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n1103_), .Y(_abc_15497_new_n2052_));
AND2X2 AND2X2_664 ( .A(d_reg_7_), .B(round_ctr_inc), .Y(_abc_15497_new_n2053_));
AND2X2 AND2X2_665 ( .A(_abc_15497_new_n2010_), .B(e_reg_8_), .Y(_abc_15497_new_n2056_));
AND2X2 AND2X2_666 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n1129_), .Y(_abc_15497_new_n2057_));
AND2X2 AND2X2_667 ( .A(d_reg_8_), .B(round_ctr_inc), .Y(_abc_15497_new_n2058_));
AND2X2 AND2X2_668 ( .A(_abc_15497_new_n2010_), .B(e_reg_9_), .Y(_abc_15497_new_n2061_));
AND2X2 AND2X2_669 ( .A(_abc_15497_new_n700_), .B(\digest[9] ), .Y(_abc_15497_new_n2062_));
AND2X2 AND2X2_67 ( .A(_abc_15497_new_n822_), .B(_abc_15497_new_n819_), .Y(_abc_15497_new_n823_));
AND2X2 AND2X2_670 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n2062_), .Y(_abc_15497_new_n2063_));
AND2X2 AND2X2_671 ( .A(d_reg_9_), .B(round_ctr_inc), .Y(_abc_15497_new_n2064_));
AND2X2 AND2X2_672 ( .A(_abc_15497_new_n2010_), .B(e_reg_10_), .Y(_abc_15497_new_n2067_));
AND2X2 AND2X2_673 ( .A(_abc_15497_new_n700_), .B(\digest[10] ), .Y(_abc_15497_new_n2068_));
AND2X2 AND2X2_674 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n2068_), .Y(_abc_15497_new_n2069_));
AND2X2 AND2X2_675 ( .A(d_reg_10_), .B(round_ctr_inc), .Y(_abc_15497_new_n2070_));
AND2X2 AND2X2_676 ( .A(_abc_15497_new_n2010_), .B(e_reg_11_), .Y(_abc_15497_new_n2073_));
AND2X2 AND2X2_677 ( .A(_abc_15497_new_n700_), .B(\digest[11] ), .Y(_abc_15497_new_n2074_));
AND2X2 AND2X2_678 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n2074_), .Y(_abc_15497_new_n2075_));
AND2X2 AND2X2_679 ( .A(d_reg_11_), .B(round_ctr_inc), .Y(_abc_15497_new_n2076_));
AND2X2 AND2X2_68 ( .A(_abc_15497_new_n825_), .B(_abc_15497_new_n826_), .Y(_abc_15497_new_n827_));
AND2X2 AND2X2_680 ( .A(_abc_15497_new_n2010_), .B(e_reg_12_), .Y(_abc_15497_new_n2079_));
AND2X2 AND2X2_681 ( .A(_abc_15497_new_n700_), .B(\digest[12] ), .Y(_abc_15497_new_n2080_));
AND2X2 AND2X2_682 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n2080_), .Y(_abc_15497_new_n2081_));
AND2X2 AND2X2_683 ( .A(d_reg_12_), .B(round_ctr_inc), .Y(_abc_15497_new_n2082_));
AND2X2 AND2X2_684 ( .A(_abc_15497_new_n2010_), .B(e_reg_13_), .Y(_abc_15497_new_n2085_));
AND2X2 AND2X2_685 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n1208_), .Y(_abc_15497_new_n2086_));
AND2X2 AND2X2_686 ( .A(d_reg_13_), .B(round_ctr_inc), .Y(_abc_15497_new_n2087_));
AND2X2 AND2X2_687 ( .A(_abc_15497_new_n2010_), .B(e_reg_14_), .Y(_abc_15497_new_n2090_));
AND2X2 AND2X2_688 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n1225_), .Y(_abc_15497_new_n2091_));
AND2X2 AND2X2_689 ( .A(d_reg_14_), .B(round_ctr_inc), .Y(_abc_15497_new_n2092_));
AND2X2 AND2X2_69 ( .A(_abc_15497_new_n824_), .B(_abc_15497_new_n827_), .Y(_abc_15497_new_n828_));
AND2X2 AND2X2_690 ( .A(_abc_15497_new_n2010_), .B(e_reg_15_), .Y(_abc_15497_new_n2095_));
AND2X2 AND2X2_691 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n1239_), .Y(_abc_15497_new_n2096_));
AND2X2 AND2X2_692 ( .A(d_reg_15_), .B(round_ctr_inc), .Y(_abc_15497_new_n2097_));
AND2X2 AND2X2_693 ( .A(_abc_15497_new_n2010_), .B(e_reg_16_), .Y(_abc_15497_new_n2100_));
AND2X2 AND2X2_694 ( .A(_abc_15497_new_n700_), .B(\digest[16] ), .Y(_abc_15497_new_n2101_));
AND2X2 AND2X2_695 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n2101_), .Y(_abc_15497_new_n2102_));
AND2X2 AND2X2_696 ( .A(d_reg_16_), .B(round_ctr_inc), .Y(_abc_15497_new_n2103_));
AND2X2 AND2X2_697 ( .A(_abc_15497_new_n2010_), .B(e_reg_17_), .Y(_abc_15497_new_n2106_));
AND2X2 AND2X2_698 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n1278_), .Y(_abc_15497_new_n2107_));
AND2X2 AND2X2_699 ( .A(d_reg_17_), .B(round_ctr_inc), .Y(_abc_15497_new_n2108_));
AND2X2 AND2X2_7 ( .A(_abc_15497_new_n708_), .B(_abc_15497_new_n709_), .Y(_abc_15497_new_n710_));
AND2X2 AND2X2_70 ( .A(_abc_15497_new_n829_), .B(_abc_15497_new_n816_), .Y(_abc_15497_new_n830_));
AND2X2 AND2X2_700 ( .A(_abc_15497_new_n2010_), .B(e_reg_18_), .Y(_abc_15497_new_n2111_));
AND2X2 AND2X2_701 ( .A(_abc_15497_new_n700_), .B(\digest[18] ), .Y(_abc_15497_new_n2112_));
AND2X2 AND2X2_702 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n2112_), .Y(_abc_15497_new_n2113_));
AND2X2 AND2X2_703 ( .A(d_reg_18_), .B(round_ctr_inc), .Y(_abc_15497_new_n2114_));
AND2X2 AND2X2_704 ( .A(_abc_15497_new_n2010_), .B(e_reg_19_), .Y(_abc_15497_new_n2117_));
AND2X2 AND2X2_705 ( .A(_abc_15497_new_n700_), .B(\digest[19] ), .Y(_abc_15497_new_n2118_));
AND2X2 AND2X2_706 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n2118_), .Y(_abc_15497_new_n2119_));
AND2X2 AND2X2_707 ( .A(d_reg_19_), .B(round_ctr_inc), .Y(_abc_15497_new_n2120_));
AND2X2 AND2X2_708 ( .A(_abc_15497_new_n2010_), .B(e_reg_20_), .Y(_abc_15497_new_n2123_));
AND2X2 AND2X2_709 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n1332_), .Y(_abc_15497_new_n2124_));
AND2X2 AND2X2_71 ( .A(_abc_15497_new_n832_), .B(_abc_15497_new_n833_), .Y(_abc_15497_new_n834_));
AND2X2 AND2X2_710 ( .A(d_reg_20_), .B(round_ctr_inc), .Y(_abc_15497_new_n2125_));
AND2X2 AND2X2_711 ( .A(_abc_15497_new_n2010_), .B(e_reg_21_), .Y(_abc_15497_new_n2128_));
AND2X2 AND2X2_712 ( .A(_abc_15497_new_n700_), .B(\digest[21] ), .Y(_abc_15497_new_n2129_));
AND2X2 AND2X2_713 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n2129_), .Y(_abc_15497_new_n2130_));
AND2X2 AND2X2_714 ( .A(d_reg_21_), .B(round_ctr_inc), .Y(_abc_15497_new_n2131_));
AND2X2 AND2X2_715 ( .A(_abc_15497_new_n2010_), .B(e_reg_22_), .Y(_abc_15497_new_n2134_));
AND2X2 AND2X2_716 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n1363_), .Y(_abc_15497_new_n2135_));
AND2X2 AND2X2_717 ( .A(d_reg_22_), .B(round_ctr_inc), .Y(_abc_15497_new_n2136_));
AND2X2 AND2X2_718 ( .A(_abc_15497_new_n2010_), .B(e_reg_23_), .Y(_abc_15497_new_n2139_));
AND2X2 AND2X2_719 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n1377_), .Y(_abc_15497_new_n2140_));
AND2X2 AND2X2_72 ( .A(_abc_15497_new_n831_), .B(_abc_15497_new_n834_), .Y(_abc_15497_new_n835_));
AND2X2 AND2X2_720 ( .A(d_reg_23_), .B(round_ctr_inc), .Y(_abc_15497_new_n2141_));
AND2X2 AND2X2_721 ( .A(_abc_15497_new_n2010_), .B(e_reg_24_), .Y(_abc_15497_new_n2144_));
AND2X2 AND2X2_722 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n1401_), .Y(_abc_15497_new_n2145_));
AND2X2 AND2X2_723 ( .A(d_reg_24_), .B(round_ctr_inc), .Y(_abc_15497_new_n2146_));
AND2X2 AND2X2_724 ( .A(_abc_15497_new_n2010_), .B(e_reg_25_), .Y(_abc_15497_new_n2149_));
AND2X2 AND2X2_725 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n1415_), .Y(_abc_15497_new_n2150_));
AND2X2 AND2X2_726 ( .A(d_reg_25_), .B(round_ctr_inc), .Y(_abc_15497_new_n2151_));
AND2X2 AND2X2_727 ( .A(_abc_15497_new_n2010_), .B(e_reg_26_), .Y(_abc_15497_new_n2154_));
AND2X2 AND2X2_728 ( .A(_abc_15497_new_n700_), .B(\digest[26] ), .Y(_abc_15497_new_n2155_));
AND2X2 AND2X2_729 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n2155_), .Y(_abc_15497_new_n2156_));
AND2X2 AND2X2_73 ( .A(_abc_15497_new_n836_), .B(_abc_15497_new_n813_), .Y(_abc_15497_new_n837_));
AND2X2 AND2X2_730 ( .A(d_reg_26_), .B(round_ctr_inc), .Y(_abc_15497_new_n2157_));
AND2X2 AND2X2_731 ( .A(_abc_15497_new_n2010_), .B(e_reg_27_), .Y(_abc_15497_new_n2160_));
AND2X2 AND2X2_732 ( .A(_abc_15497_new_n700_), .B(\digest[27] ), .Y(_abc_15497_new_n2161_));
AND2X2 AND2X2_733 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n2161_), .Y(_abc_15497_new_n2162_));
AND2X2 AND2X2_734 ( .A(d_reg_27_), .B(round_ctr_inc), .Y(_abc_15497_new_n2163_));
AND2X2 AND2X2_735 ( .A(_abc_15497_new_n2010_), .B(e_reg_28_), .Y(_abc_15497_new_n2166_));
AND2X2 AND2X2_736 ( .A(_abc_15497_new_n700_), .B(\digest[28] ), .Y(_abc_15497_new_n2167_));
AND2X2 AND2X2_737 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n2167_), .Y(_abc_15497_new_n2168_));
AND2X2 AND2X2_738 ( .A(d_reg_28_), .B(round_ctr_inc), .Y(_abc_15497_new_n2169_));
AND2X2 AND2X2_739 ( .A(_abc_15497_new_n2010_), .B(e_reg_29_), .Y(_abc_15497_new_n2172_));
AND2X2 AND2X2_74 ( .A(_abc_15497_new_n838_), .B(_abc_15497_new_n811_), .Y(_abc_15497_new_n839_));
AND2X2 AND2X2_740 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n1481_), .Y(_abc_15497_new_n2173_));
AND2X2 AND2X2_741 ( .A(d_reg_29_), .B(round_ctr_inc), .Y(_abc_15497_new_n2174_));
AND2X2 AND2X2_742 ( .A(_abc_15497_new_n2010_), .B(e_reg_30_), .Y(_abc_15497_new_n2177_));
AND2X2 AND2X2_743 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n1510_), .Y(_abc_15497_new_n2178_));
AND2X2 AND2X2_744 ( .A(d_reg_30_), .B(round_ctr_inc), .Y(_abc_15497_new_n2179_));
AND2X2 AND2X2_745 ( .A(_abc_15497_new_n2010_), .B(e_reg_31_), .Y(_abc_15497_new_n2182_));
AND2X2 AND2X2_746 ( .A(_abc_15497_new_n2013_), .B(_abc_15497_new_n1526_), .Y(_abc_15497_new_n2183_));
AND2X2 AND2X2_747 ( .A(d_reg_31_), .B(round_ctr_inc), .Y(_abc_15497_new_n2184_));
AND2X2 AND2X2_748 ( .A(\digest[96] ), .B(b_reg_0_), .Y(_abc_15497_new_n2188_));
AND2X2 AND2X2_749 ( .A(_abc_15497_new_n2189_), .B(digest_update), .Y(_abc_15497_new_n2190_));
AND2X2 AND2X2_75 ( .A(_abc_15497_new_n841_), .B(_abc_15497_new_n797_), .Y(_abc_15497_new_n842_));
AND2X2 AND2X2_750 ( .A(_abc_15497_new_n2190_), .B(_abc_15497_new_n2187_), .Y(_abc_15497_new_n2191_));
AND2X2 AND2X2_751 ( .A(_abc_15497_new_n2192_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n2193_));
AND2X2 AND2X2_752 ( .A(\digest[97] ), .B(b_reg_1_), .Y(_abc_15497_new_n2197_));
AND2X2 AND2X2_753 ( .A(_abc_15497_new_n2200_), .B(_abc_15497_new_n2195_), .Y(_abc_15497_new_n2201_));
AND2X2 AND2X2_754 ( .A(_abc_15497_new_n2202_), .B(digest_update), .Y(_abc_15497_new_n2203_));
AND2X2 AND2X2_755 ( .A(_abc_15497_new_n2203_), .B(_abc_15497_new_n2199_), .Y(_abc_15497_new_n2204_));
AND2X2 AND2X2_756 ( .A(_abc_15497_new_n701_), .B(\digest[97] ), .Y(_abc_15497_new_n2205_));
AND2X2 AND2X2_757 ( .A(_abc_15497_new_n2199_), .B(_abc_15497_new_n2200_), .Y(_abc_15497_new_n2207_));
AND2X2 AND2X2_758 ( .A(\digest[98] ), .B(b_reg_2_), .Y(_abc_15497_new_n2209_));
AND2X2 AND2X2_759 ( .A(_abc_15497_new_n2210_), .B(_abc_15497_new_n2208_), .Y(_abc_15497_new_n2211_));
AND2X2 AND2X2_76 ( .A(_abc_15497_new_n843_), .B(_abc_15497_new_n844_), .Y(_abc_15497_new_n845_));
AND2X2 AND2X2_760 ( .A(_abc_15497_new_n2201_), .B(_abc_15497_new_n2188_), .Y(_abc_15497_new_n2214_));
AND2X2 AND2X2_761 ( .A(_abc_15497_new_n2216_), .B(digest_update), .Y(_abc_15497_new_n2217_));
AND2X2 AND2X2_762 ( .A(_abc_15497_new_n2217_), .B(_abc_15497_new_n2213_), .Y(_abc_15497_new_n2218_));
AND2X2 AND2X2_763 ( .A(_abc_15497_new_n701_), .B(\digest[98] ), .Y(_abc_15497_new_n2219_));
AND2X2 AND2X2_764 ( .A(_abc_15497_new_n2215_), .B(_abc_15497_new_n2211_), .Y(_abc_15497_new_n2221_));
AND2X2 AND2X2_765 ( .A(\digest[99] ), .B(b_reg_3_), .Y(_abc_15497_new_n2224_));
AND2X2 AND2X2_766 ( .A(_abc_15497_new_n2225_), .B(_abc_15497_new_n2223_), .Y(_abc_15497_new_n2226_));
AND2X2 AND2X2_767 ( .A(_abc_15497_new_n2213_), .B(_abc_15497_new_n2210_), .Y(_abc_15497_new_n2228_));
AND2X2 AND2X2_768 ( .A(_abc_15497_new_n2230_), .B(_abc_15497_new_n2227_), .Y(_abc_15497_new_n2231_));
AND2X2 AND2X2_769 ( .A(_abc_15497_new_n2231_), .B(digest_update), .Y(_abc_15497_new_n2232_));
AND2X2 AND2X2_77 ( .A(_abc_15497_new_n842_), .B(_abc_15497_new_n845_), .Y(_abc_15497_new_n846_));
AND2X2 AND2X2_770 ( .A(_abc_15497_new_n2233_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n2234_));
AND2X2 AND2X2_771 ( .A(\digest[100] ), .B(b_reg_4_), .Y(_abc_15497_new_n2237_));
AND2X2 AND2X2_772 ( .A(_abc_15497_new_n2238_), .B(_abc_15497_new_n2236_), .Y(_abc_15497_new_n2239_));
AND2X2 AND2X2_773 ( .A(_abc_15497_new_n2242_), .B(_abc_15497_new_n2225_), .Y(_abc_15497_new_n2243_));
AND2X2 AND2X2_774 ( .A(_abc_15497_new_n2222_), .B(_abc_15497_new_n2223_), .Y(_abc_15497_new_n2245_));
AND2X2 AND2X2_775 ( .A(_abc_15497_new_n2247_), .B(digest_update), .Y(_abc_15497_new_n2248_));
AND2X2 AND2X2_776 ( .A(_abc_15497_new_n2248_), .B(_abc_15497_new_n2244_), .Y(_abc_15497_new_n2249_));
AND2X2 AND2X2_777 ( .A(_abc_15497_new_n701_), .B(\digest[100] ), .Y(_abc_15497_new_n2250_));
AND2X2 AND2X2_778 ( .A(_abc_15497_new_n701_), .B(\digest[101] ), .Y(_abc_15497_new_n2252_));
AND2X2 AND2X2_779 ( .A(_abc_15497_new_n2246_), .B(_abc_15497_new_n2239_), .Y(_abc_15497_new_n2253_));
AND2X2 AND2X2_78 ( .A(_abc_15497_new_n840_), .B(_abc_15497_new_n846_), .Y(_abc_15497_new_n847_));
AND2X2 AND2X2_780 ( .A(\digest[101] ), .B(b_reg_5_), .Y(_abc_15497_new_n2256_));
AND2X2 AND2X2_781 ( .A(_abc_15497_new_n2257_), .B(_abc_15497_new_n2255_), .Y(_abc_15497_new_n2258_));
AND2X2 AND2X2_782 ( .A(_abc_15497_new_n2244_), .B(_abc_15497_new_n2238_), .Y(_abc_15497_new_n2260_));
AND2X2 AND2X2_783 ( .A(_abc_15497_new_n2262_), .B(_abc_15497_new_n2259_), .Y(_abc_15497_new_n2263_));
AND2X2 AND2X2_784 ( .A(_abc_15497_new_n2263_), .B(digest_update), .Y(_abc_15497_new_n2264_));
AND2X2 AND2X2_785 ( .A(_abc_15497_new_n701_), .B(\digest[102] ), .Y(_abc_15497_new_n2266_));
AND2X2 AND2X2_786 ( .A(_abc_15497_new_n2254_), .B(_abc_15497_new_n2258_), .Y(_abc_15497_new_n2267_));
AND2X2 AND2X2_787 ( .A(\digest[102] ), .B(b_reg_6_), .Y(_abc_15497_new_n2270_));
AND2X2 AND2X2_788 ( .A(_abc_15497_new_n2271_), .B(_abc_15497_new_n2269_), .Y(_abc_15497_new_n2272_));
AND2X2 AND2X2_789 ( .A(_abc_15497_new_n2262_), .B(_abc_15497_new_n2257_), .Y(_abc_15497_new_n2274_));
AND2X2 AND2X2_79 ( .A(_abc_15497_new_n848_), .B(_abc_15497_new_n795_), .Y(_abc_15497_new_n849_));
AND2X2 AND2X2_790 ( .A(_abc_15497_new_n2276_), .B(_abc_15497_new_n2273_), .Y(_abc_15497_new_n2277_));
AND2X2 AND2X2_791 ( .A(_abc_15497_new_n2277_), .B(digest_update), .Y(_abc_15497_new_n2278_));
AND2X2 AND2X2_792 ( .A(_abc_15497_new_n2276_), .B(_abc_15497_new_n2271_), .Y(_abc_15497_new_n2282_));
AND2X2 AND2X2_793 ( .A(\digest[103] ), .B(b_reg_7_), .Y(_abc_15497_new_n2284_));
AND2X2 AND2X2_794 ( .A(_abc_15497_new_n2285_), .B(_abc_15497_new_n2283_), .Y(_abc_15497_new_n2286_));
AND2X2 AND2X2_795 ( .A(_abc_15497_new_n2282_), .B(_abc_15497_new_n2286_), .Y(_abc_15497_new_n2287_));
AND2X2 AND2X2_796 ( .A(_abc_15497_new_n2268_), .B(_abc_15497_new_n2272_), .Y(_abc_15497_new_n2288_));
AND2X2 AND2X2_797 ( .A(_abc_15497_new_n2289_), .B(_abc_15497_new_n2290_), .Y(_abc_15497_new_n2291_));
AND2X2 AND2X2_798 ( .A(_abc_15497_new_n2293_), .B(_abc_15497_new_n2281_), .Y(_0H1_reg_31_0__7_));
AND2X2 AND2X2_799 ( .A(\digest[104] ), .B(b_reg_8_), .Y(_abc_15497_new_n2296_));
AND2X2 AND2X2_8 ( .A(_abc_15497_new_n706_), .B(_abc_15497_new_n710_), .Y(_abc_15497_new_n711_));
AND2X2 AND2X2_80 ( .A(_abc_15497_new_n850_), .B(_abc_15497_new_n784_), .Y(_abc_15497_new_n851_));
AND2X2 AND2X2_800 ( .A(_abc_15497_new_n2297_), .B(_abc_15497_new_n2295_), .Y(_abc_15497_new_n2298_));
AND2X2 AND2X2_801 ( .A(_abc_15497_new_n2289_), .B(_abc_15497_new_n2283_), .Y(_abc_15497_new_n2299_));
AND2X2 AND2X2_802 ( .A(_abc_15497_new_n2300_), .B(_abc_15497_new_n2298_), .Y(_abc_15497_new_n2302_));
AND2X2 AND2X2_803 ( .A(_abc_15497_new_n2303_), .B(_abc_15497_new_n2301_), .Y(_abc_15497_new_n2304_));
AND2X2 AND2X2_804 ( .A(_abc_15497_new_n2304_), .B(digest_update), .Y(_abc_15497_new_n2305_));
AND2X2 AND2X2_805 ( .A(_abc_15497_new_n2306_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n2307_));
AND2X2 AND2X2_806 ( .A(_abc_15497_new_n2303_), .B(_abc_15497_new_n2297_), .Y(_abc_15497_new_n2309_));
AND2X2 AND2X2_807 ( .A(\digest[105] ), .B(b_reg_9_), .Y(_abc_15497_new_n2312_));
AND2X2 AND2X2_808 ( .A(_abc_15497_new_n2313_), .B(_abc_15497_new_n2311_), .Y(_abc_15497_new_n2314_));
AND2X2 AND2X2_809 ( .A(_abc_15497_new_n2315_), .B(_abc_15497_new_n2317_), .Y(_abc_15497_new_n2318_));
AND2X2 AND2X2_81 ( .A(_abc_15497_new_n746_), .B(_abc_15497_new_n853_), .Y(_abc_15497_new_n854_));
AND2X2 AND2X2_810 ( .A(_abc_15497_new_n2318_), .B(digest_update), .Y(_abc_15497_new_n2319_));
AND2X2 AND2X2_811 ( .A(_abc_15497_new_n2320_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n2321_));
AND2X2 AND2X2_812 ( .A(_abc_15497_new_n701_), .B(\digest[106] ), .Y(_abc_15497_new_n2323_));
AND2X2 AND2X2_813 ( .A(_abc_15497_new_n2298_), .B(_abc_15497_new_n2314_), .Y(_abc_15497_new_n2324_));
AND2X2 AND2X2_814 ( .A(_abc_15497_new_n2300_), .B(_abc_15497_new_n2324_), .Y(_abc_15497_new_n2325_));
AND2X2 AND2X2_815 ( .A(_abc_15497_new_n2326_), .B(_abc_15497_new_n2313_), .Y(_abc_15497_new_n2327_));
AND2X2 AND2X2_816 ( .A(\digest[106] ), .B(b_reg_10_), .Y(_abc_15497_new_n2331_));
AND2X2 AND2X2_817 ( .A(_abc_15497_new_n2332_), .B(_abc_15497_new_n2330_), .Y(_abc_15497_new_n2333_));
AND2X2 AND2X2_818 ( .A(_abc_15497_new_n2329_), .B(_abc_15497_new_n2333_), .Y(_abc_15497_new_n2335_));
AND2X2 AND2X2_819 ( .A(_abc_15497_new_n2336_), .B(_abc_15497_new_n2334_), .Y(_abc_15497_new_n2337_));
AND2X2 AND2X2_82 ( .A(_abc_15497_new_n743_), .B(_abc_15497_new_n854_), .Y(_abc_15497_new_n855_));
AND2X2 AND2X2_820 ( .A(_abc_15497_new_n2337_), .B(digest_update), .Y(_abc_15497_new_n2338_));
AND2X2 AND2X2_821 ( .A(_abc_15497_new_n2336_), .B(_abc_15497_new_n2332_), .Y(_abc_15497_new_n2340_));
AND2X2 AND2X2_822 ( .A(\digest[107] ), .B(b_reg_11_), .Y(_abc_15497_new_n2342_));
AND2X2 AND2X2_823 ( .A(_abc_15497_new_n2343_), .B(_abc_15497_new_n2341_), .Y(_abc_15497_new_n2344_));
AND2X2 AND2X2_824 ( .A(_abc_15497_new_n2340_), .B(_abc_15497_new_n2344_), .Y(_abc_15497_new_n2345_));
AND2X2 AND2X2_825 ( .A(_abc_15497_new_n2346_), .B(_abc_15497_new_n2347_), .Y(_abc_15497_new_n2348_));
AND2X2 AND2X2_826 ( .A(_abc_15497_new_n2349_), .B(digest_update), .Y(_abc_15497_new_n2350_));
AND2X2 AND2X2_827 ( .A(_abc_15497_new_n2351_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n2352_));
AND2X2 AND2X2_828 ( .A(_abc_15497_new_n701_), .B(\digest[108] ), .Y(_abc_15497_new_n2354_));
AND2X2 AND2X2_829 ( .A(\digest[108] ), .B(b_reg_12_), .Y(_abc_15497_new_n2356_));
AND2X2 AND2X2_83 ( .A(_abc_15497_new_n739_), .B(_abc_15497_new_n855_), .Y(_abc_15497_new_n856_));
AND2X2 AND2X2_830 ( .A(_abc_15497_new_n2357_), .B(_abc_15497_new_n2355_), .Y(_abc_15497_new_n2358_));
AND2X2 AND2X2_831 ( .A(_abc_15497_new_n2341_), .B(_abc_15497_new_n2331_), .Y(_abc_15497_new_n2359_));
AND2X2 AND2X2_832 ( .A(_abc_15497_new_n2333_), .B(_abc_15497_new_n2344_), .Y(_abc_15497_new_n2361_));
AND2X2 AND2X2_833 ( .A(_abc_15497_new_n2328_), .B(_abc_15497_new_n2361_), .Y(_abc_15497_new_n2362_));
AND2X2 AND2X2_834 ( .A(_abc_15497_new_n2324_), .B(_abc_15497_new_n2361_), .Y(_abc_15497_new_n2364_));
AND2X2 AND2X2_835 ( .A(_abc_15497_new_n2300_), .B(_abc_15497_new_n2364_), .Y(_abc_15497_new_n2365_));
AND2X2 AND2X2_836 ( .A(_abc_15497_new_n2366_), .B(_abc_15497_new_n2358_), .Y(_abc_15497_new_n2368_));
AND2X2 AND2X2_837 ( .A(_abc_15497_new_n2369_), .B(_abc_15497_new_n2367_), .Y(_abc_15497_new_n2370_));
AND2X2 AND2X2_838 ( .A(_abc_15497_new_n2370_), .B(digest_update), .Y(_abc_15497_new_n2371_));
AND2X2 AND2X2_839 ( .A(_abc_15497_new_n2369_), .B(_abc_15497_new_n2357_), .Y(_abc_15497_new_n2373_));
AND2X2 AND2X2_84 ( .A(_abc_15497_new_n730_), .B(_abc_15497_new_n856_), .Y(_abc_15497_new_n857_));
AND2X2 AND2X2_840 ( .A(\digest[109] ), .B(b_reg_13_), .Y(_abc_15497_new_n2376_));
AND2X2 AND2X2_841 ( .A(_abc_15497_new_n2377_), .B(_abc_15497_new_n2375_), .Y(_abc_15497_new_n2378_));
AND2X2 AND2X2_842 ( .A(_abc_15497_new_n2379_), .B(_abc_15497_new_n2381_), .Y(_abc_15497_new_n2382_));
AND2X2 AND2X2_843 ( .A(_abc_15497_new_n2382_), .B(digest_update), .Y(_abc_15497_new_n2383_));
AND2X2 AND2X2_844 ( .A(_abc_15497_new_n2384_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n2385_));
AND2X2 AND2X2_845 ( .A(_abc_15497_new_n701_), .B(\digest[110] ), .Y(_abc_15497_new_n2387_));
AND2X2 AND2X2_846 ( .A(\digest[110] ), .B(b_reg_14_), .Y(_abc_15497_new_n2389_));
AND2X2 AND2X2_847 ( .A(_abc_15497_new_n2390_), .B(_abc_15497_new_n2388_), .Y(_abc_15497_new_n2391_));
AND2X2 AND2X2_848 ( .A(_abc_15497_new_n2357_), .B(_abc_15497_new_n2377_), .Y(_abc_15497_new_n2393_));
AND2X2 AND2X2_849 ( .A(_abc_15497_new_n2369_), .B(_abc_15497_new_n2393_), .Y(_abc_15497_new_n2394_));
AND2X2 AND2X2_85 ( .A(_abc_15497_new_n852_), .B(_abc_15497_new_n857_), .Y(_abc_15497_new_n858_));
AND2X2 AND2X2_850 ( .A(_abc_15497_new_n2396_), .B(_abc_15497_new_n2391_), .Y(_abc_15497_new_n2398_));
AND2X2 AND2X2_851 ( .A(_abc_15497_new_n2399_), .B(_abc_15497_new_n2397_), .Y(_abc_15497_new_n2400_));
AND2X2 AND2X2_852 ( .A(_abc_15497_new_n2400_), .B(digest_update), .Y(_abc_15497_new_n2401_));
AND2X2 AND2X2_853 ( .A(_abc_15497_new_n2399_), .B(_abc_15497_new_n2390_), .Y(_abc_15497_new_n2403_));
AND2X2 AND2X2_854 ( .A(\digest[111] ), .B(b_reg_15_), .Y(_abc_15497_new_n2406_));
AND2X2 AND2X2_855 ( .A(_abc_15497_new_n2407_), .B(_abc_15497_new_n2405_), .Y(_abc_15497_new_n2408_));
AND2X2 AND2X2_856 ( .A(_abc_15497_new_n2409_), .B(_abc_15497_new_n2411_), .Y(_abc_15497_new_n2412_));
AND2X2 AND2X2_857 ( .A(_abc_15497_new_n2412_), .B(digest_update), .Y(_abc_15497_new_n2413_));
AND2X2 AND2X2_858 ( .A(_abc_15497_new_n2414_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n2415_));
AND2X2 AND2X2_859 ( .A(_abc_15497_new_n2408_), .B(_abc_15497_new_n2389_), .Y(_abc_15497_new_n2417_));
AND2X2 AND2X2_86 ( .A(c_reg_25_), .B(\digest[89] ), .Y(_abc_15497_new_n860_));
AND2X2 AND2X2_860 ( .A(_abc_15497_new_n2391_), .B(_abc_15497_new_n2408_), .Y(_abc_15497_new_n2421_));
AND2X2 AND2X2_861 ( .A(_abc_15497_new_n2423_), .B(_abc_15497_new_n2419_), .Y(_abc_15497_new_n2424_));
AND2X2 AND2X2_862 ( .A(_abc_15497_new_n2358_), .B(_abc_15497_new_n2378_), .Y(_abc_15497_new_n2426_));
AND2X2 AND2X2_863 ( .A(_abc_15497_new_n2426_), .B(_abc_15497_new_n2421_), .Y(_abc_15497_new_n2427_));
AND2X2 AND2X2_864 ( .A(_abc_15497_new_n2366_), .B(_abc_15497_new_n2427_), .Y(_abc_15497_new_n2428_));
AND2X2 AND2X2_865 ( .A(\digest[112] ), .B(b_reg_16_), .Y(_abc_15497_new_n2431_));
AND2X2 AND2X2_866 ( .A(_abc_15497_new_n2432_), .B(_abc_15497_new_n2430_), .Y(_abc_15497_new_n2433_));
AND2X2 AND2X2_867 ( .A(_abc_15497_new_n2429_), .B(_abc_15497_new_n2433_), .Y(_abc_15497_new_n2435_));
AND2X2 AND2X2_868 ( .A(_abc_15497_new_n2436_), .B(_abc_15497_new_n2434_), .Y(_abc_15497_new_n2437_));
AND2X2 AND2X2_869 ( .A(_abc_15497_new_n2437_), .B(digest_update), .Y(_abc_15497_new_n2438_));
AND2X2 AND2X2_87 ( .A(_abc_15497_new_n861_), .B(_abc_15497_new_n862_), .Y(_abc_15497_new_n863_));
AND2X2 AND2X2_870 ( .A(_abc_15497_new_n2439_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n2440_));
AND2X2 AND2X2_871 ( .A(_abc_15497_new_n701_), .B(\digest[113] ), .Y(_abc_15497_new_n2442_));
AND2X2 AND2X2_872 ( .A(\digest[113] ), .B(b_reg_17_), .Y(_abc_15497_new_n2444_));
AND2X2 AND2X2_873 ( .A(_abc_15497_new_n2445_), .B(_abc_15497_new_n2443_), .Y(_abc_15497_new_n2446_));
AND2X2 AND2X2_874 ( .A(_abc_15497_new_n2433_), .B(_abc_15497_new_n2446_), .Y(_abc_15497_new_n2449_));
AND2X2 AND2X2_875 ( .A(_abc_15497_new_n2429_), .B(_abc_15497_new_n2449_), .Y(_abc_15497_new_n2450_));
AND2X2 AND2X2_876 ( .A(_abc_15497_new_n2446_), .B(_abc_15497_new_n2431_), .Y(_abc_15497_new_n2452_));
AND2X2 AND2X2_877 ( .A(_abc_15497_new_n2453_), .B(digest_update), .Y(_abc_15497_new_n2454_));
AND2X2 AND2X2_878 ( .A(_abc_15497_new_n2451_), .B(_abc_15497_new_n2454_), .Y(_abc_15497_new_n2455_));
AND2X2 AND2X2_879 ( .A(_abc_15497_new_n2455_), .B(_abc_15497_new_n2448_), .Y(_abc_15497_new_n2456_));
AND2X2 AND2X2_88 ( .A(c_reg_24_), .B(\digest[88] ), .Y(_abc_15497_new_n864_));
AND2X2 AND2X2_880 ( .A(_abc_15497_new_n2453_), .B(_abc_15497_new_n2445_), .Y(_abc_15497_new_n2458_));
AND2X2 AND2X2_881 ( .A(_abc_15497_new_n2451_), .B(_abc_15497_new_n2458_), .Y(_abc_15497_new_n2459_));
AND2X2 AND2X2_882 ( .A(\digest[114] ), .B(b_reg_18_), .Y(_abc_15497_new_n2462_));
AND2X2 AND2X2_883 ( .A(_abc_15497_new_n2463_), .B(_abc_15497_new_n2461_), .Y(_abc_15497_new_n2464_));
AND2X2 AND2X2_884 ( .A(_abc_15497_new_n2460_), .B(_abc_15497_new_n2464_), .Y(_abc_15497_new_n2466_));
AND2X2 AND2X2_885 ( .A(_abc_15497_new_n2467_), .B(_abc_15497_new_n2465_), .Y(_abc_15497_new_n2468_));
AND2X2 AND2X2_886 ( .A(_abc_15497_new_n2468_), .B(digest_update), .Y(_abc_15497_new_n2469_));
AND2X2 AND2X2_887 ( .A(_abc_15497_new_n2470_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n2471_));
AND2X2 AND2X2_888 ( .A(_abc_15497_new_n2467_), .B(_abc_15497_new_n2463_), .Y(_abc_15497_new_n2473_));
AND2X2 AND2X2_889 ( .A(\digest[115] ), .B(b_reg_19_), .Y(_abc_15497_new_n2475_));
AND2X2 AND2X2_89 ( .A(_abc_15497_new_n865_), .B(_abc_15497_new_n866_), .Y(_abc_15497_new_n867_));
AND2X2 AND2X2_890 ( .A(_abc_15497_new_n2476_), .B(_abc_15497_new_n2474_), .Y(_abc_15497_new_n2477_));
AND2X2 AND2X2_891 ( .A(_abc_15497_new_n2473_), .B(_abc_15497_new_n2477_), .Y(_abc_15497_new_n2478_));
AND2X2 AND2X2_892 ( .A(_abc_15497_new_n2479_), .B(_abc_15497_new_n2480_), .Y(_abc_15497_new_n2481_));
AND2X2 AND2X2_893 ( .A(_abc_15497_new_n2482_), .B(digest_update), .Y(_abc_15497_new_n2483_));
AND2X2 AND2X2_894 ( .A(_abc_15497_new_n2484_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n2485_));
AND2X2 AND2X2_895 ( .A(_abc_15497_new_n701_), .B(\digest[116] ), .Y(_abc_15497_new_n2487_));
AND2X2 AND2X2_896 ( .A(_abc_15497_new_n2464_), .B(_abc_15497_new_n2477_), .Y(_abc_15497_new_n2488_));
AND2X2 AND2X2_897 ( .A(_abc_15497_new_n2474_), .B(_abc_15497_new_n2462_), .Y(_abc_15497_new_n2491_));
AND2X2 AND2X2_898 ( .A(_abc_15497_new_n2490_), .B(_abc_15497_new_n2493_), .Y(_abc_15497_new_n2494_));
AND2X2 AND2X2_899 ( .A(_abc_15497_new_n2449_), .B(_abc_15497_new_n2488_), .Y(_abc_15497_new_n2496_));
AND2X2 AND2X2_9 ( .A(c_reg_21_), .B(\digest[85] ), .Y(_abc_15497_new_n713_));
AND2X2 AND2X2_90 ( .A(_abc_15497_new_n863_), .B(_abc_15497_new_n867_), .Y(_abc_15497_new_n868_));
AND2X2 AND2X2_900 ( .A(_abc_15497_new_n2429_), .B(_abc_15497_new_n2496_), .Y(_abc_15497_new_n2497_));
AND2X2 AND2X2_901 ( .A(\digest[116] ), .B(b_reg_20_), .Y(_abc_15497_new_n2500_));
AND2X2 AND2X2_902 ( .A(_abc_15497_new_n2501_), .B(_abc_15497_new_n2499_), .Y(_abc_15497_new_n2502_));
AND2X2 AND2X2_903 ( .A(_abc_15497_new_n2498_), .B(_abc_15497_new_n2502_), .Y(_abc_15497_new_n2504_));
AND2X2 AND2X2_904 ( .A(_abc_15497_new_n2505_), .B(_abc_15497_new_n2503_), .Y(_abc_15497_new_n2506_));
AND2X2 AND2X2_905 ( .A(_abc_15497_new_n2506_), .B(digest_update), .Y(_abc_15497_new_n2507_));
AND2X2 AND2X2_906 ( .A(_abc_15497_new_n701_), .B(\digest[117] ), .Y(_abc_15497_new_n2509_));
AND2X2 AND2X2_907 ( .A(\digest[117] ), .B(b_reg_21_), .Y(_abc_15497_new_n2511_));
AND2X2 AND2X2_908 ( .A(_abc_15497_new_n2512_), .B(_abc_15497_new_n2510_), .Y(_abc_15497_new_n2513_));
AND2X2 AND2X2_909 ( .A(_abc_15497_new_n2502_), .B(_abc_15497_new_n2513_), .Y(_abc_15497_new_n2516_));
AND2X2 AND2X2_91 ( .A(_abc_15497_new_n859_), .B(_abc_15497_new_n868_), .Y(_abc_15497_new_n869_));
AND2X2 AND2X2_910 ( .A(_abc_15497_new_n2498_), .B(_abc_15497_new_n2516_), .Y(_abc_15497_new_n2517_));
AND2X2 AND2X2_911 ( .A(_abc_15497_new_n2513_), .B(_abc_15497_new_n2500_), .Y(_abc_15497_new_n2518_));
AND2X2 AND2X2_912 ( .A(_abc_15497_new_n2520_), .B(digest_update), .Y(_abc_15497_new_n2521_));
AND2X2 AND2X2_913 ( .A(_abc_15497_new_n2521_), .B(_abc_15497_new_n2515_), .Y(_abc_15497_new_n2522_));
AND2X2 AND2X2_914 ( .A(_abc_15497_new_n2520_), .B(_abc_15497_new_n2512_), .Y(_abc_15497_new_n2524_));
AND2X2 AND2X2_915 ( .A(\digest[118] ), .B(b_reg_22_), .Y(_abc_15497_new_n2527_));
AND2X2 AND2X2_916 ( .A(_abc_15497_new_n2528_), .B(_abc_15497_new_n2526_), .Y(_abc_15497_new_n2529_));
AND2X2 AND2X2_917 ( .A(_abc_15497_new_n2525_), .B(_abc_15497_new_n2529_), .Y(_abc_15497_new_n2531_));
AND2X2 AND2X2_918 ( .A(_abc_15497_new_n2532_), .B(_abc_15497_new_n2530_), .Y(_abc_15497_new_n2533_));
AND2X2 AND2X2_919 ( .A(_abc_15497_new_n2533_), .B(digest_update), .Y(_abc_15497_new_n2534_));
AND2X2 AND2X2_92 ( .A(_abc_15497_new_n862_), .B(_abc_15497_new_n864_), .Y(_abc_15497_new_n870_));
AND2X2 AND2X2_920 ( .A(_abc_15497_new_n2535_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n2536_));
AND2X2 AND2X2_921 ( .A(\digest[119] ), .B(b_reg_23_), .Y(_abc_15497_new_n2541_));
AND2X2 AND2X2_922 ( .A(_abc_15497_new_n2542_), .B(_abc_15497_new_n2540_), .Y(_abc_15497_new_n2543_));
AND2X2 AND2X2_923 ( .A(_abc_15497_new_n2539_), .B(_abc_15497_new_n2543_), .Y(_abc_15497_new_n2544_));
AND2X2 AND2X2_924 ( .A(_abc_15497_new_n2538_), .B(_abc_15497_new_n2545_), .Y(_abc_15497_new_n2546_));
AND2X2 AND2X2_925 ( .A(_abc_15497_new_n2547_), .B(digest_update), .Y(_abc_15497_new_n2548_));
AND2X2 AND2X2_926 ( .A(_abc_15497_new_n2549_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n2550_));
AND2X2 AND2X2_927 ( .A(_abc_15497_new_n2529_), .B(_abc_15497_new_n2543_), .Y(_abc_15497_new_n2552_));
AND2X2 AND2X2_928 ( .A(_abc_15497_new_n2516_), .B(_abc_15497_new_n2552_), .Y(_abc_15497_new_n2553_));
AND2X2 AND2X2_929 ( .A(_abc_15497_new_n2495_), .B(_abc_15497_new_n2553_), .Y(_abc_15497_new_n2554_));
AND2X2 AND2X2_93 ( .A(\digest[90] ), .B(c_reg_26_), .Y(_abc_15497_new_n874_));
AND2X2 AND2X2_930 ( .A(_abc_15497_new_n2540_), .B(_abc_15497_new_n2527_), .Y(_abc_15497_new_n2555_));
AND2X2 AND2X2_931 ( .A(_abc_15497_new_n2557_), .B(_abc_15497_new_n2552_), .Y(_abc_15497_new_n2558_));
AND2X2 AND2X2_932 ( .A(_abc_15497_new_n2496_), .B(_abc_15497_new_n2553_), .Y(_abc_15497_new_n2561_));
AND2X2 AND2X2_933 ( .A(_abc_15497_new_n2429_), .B(_abc_15497_new_n2561_), .Y(_abc_15497_new_n2562_));
AND2X2 AND2X2_934 ( .A(\digest[120] ), .B(b_reg_24_), .Y(_abc_15497_new_n2565_));
AND2X2 AND2X2_935 ( .A(_abc_15497_new_n2566_), .B(_abc_15497_new_n2564_), .Y(_abc_15497_new_n2567_));
AND2X2 AND2X2_936 ( .A(_abc_15497_new_n2563_), .B(_abc_15497_new_n2567_), .Y(_abc_15497_new_n2569_));
AND2X2 AND2X2_937 ( .A(_abc_15497_new_n2570_), .B(_abc_15497_new_n2568_), .Y(_abc_15497_new_n2571_));
AND2X2 AND2X2_938 ( .A(_abc_15497_new_n2571_), .B(digest_update), .Y(_abc_15497_new_n2572_));
AND2X2 AND2X2_939 ( .A(_abc_15497_new_n2573_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n2574_));
AND2X2 AND2X2_94 ( .A(_abc_15497_new_n875_), .B(_abc_15497_new_n873_), .Y(_abc_15497_new_n876_));
AND2X2 AND2X2_940 ( .A(_abc_15497_new_n2570_), .B(_abc_15497_new_n2566_), .Y(_abc_15497_new_n2576_));
AND2X2 AND2X2_941 ( .A(\digest[121] ), .B(b_reg_25_), .Y(_abc_15497_new_n2579_));
AND2X2 AND2X2_942 ( .A(_abc_15497_new_n2580_), .B(_abc_15497_new_n2578_), .Y(_abc_15497_new_n2581_));
AND2X2 AND2X2_943 ( .A(_abc_15497_new_n2582_), .B(_abc_15497_new_n2584_), .Y(_abc_15497_new_n2585_));
AND2X2 AND2X2_944 ( .A(_abc_15497_new_n2585_), .B(digest_update), .Y(_abc_15497_new_n2586_));
AND2X2 AND2X2_945 ( .A(_abc_15497_new_n2587_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n2588_));
AND2X2 AND2X2_946 ( .A(_abc_15497_new_n2567_), .B(_abc_15497_new_n2581_), .Y(_abc_15497_new_n2590_));
AND2X2 AND2X2_947 ( .A(_abc_15497_new_n2563_), .B(_abc_15497_new_n2590_), .Y(_abc_15497_new_n2591_));
AND2X2 AND2X2_948 ( .A(_abc_15497_new_n2578_), .B(_abc_15497_new_n2565_), .Y(_abc_15497_new_n2592_));
AND2X2 AND2X2_949 ( .A(\digest[122] ), .B(b_reg_26_), .Y(_abc_15497_new_n2596_));
AND2X2 AND2X2_95 ( .A(_abc_15497_new_n872_), .B(_abc_15497_new_n876_), .Y(_abc_15497_new_n878_));
AND2X2 AND2X2_950 ( .A(_abc_15497_new_n2597_), .B(_abc_15497_new_n2595_), .Y(_abc_15497_new_n2598_));
AND2X2 AND2X2_951 ( .A(_abc_15497_new_n2594_), .B(_abc_15497_new_n2598_), .Y(_abc_15497_new_n2600_));
AND2X2 AND2X2_952 ( .A(_abc_15497_new_n2601_), .B(_abc_15497_new_n2599_), .Y(_abc_15497_new_n2602_));
AND2X2 AND2X2_953 ( .A(_abc_15497_new_n2602_), .B(digest_update), .Y(_abc_15497_new_n2603_));
AND2X2 AND2X2_954 ( .A(_abc_15497_new_n2604_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n2605_));
AND2X2 AND2X2_955 ( .A(_abc_15497_new_n2601_), .B(_abc_15497_new_n2597_), .Y(_abc_15497_new_n2607_));
AND2X2 AND2X2_956 ( .A(\digest[123] ), .B(b_reg_27_), .Y(_abc_15497_new_n2610_));
AND2X2 AND2X2_957 ( .A(_abc_15497_new_n2611_), .B(_abc_15497_new_n2609_), .Y(_abc_15497_new_n2612_));
AND2X2 AND2X2_958 ( .A(_abc_15497_new_n2613_), .B(_abc_15497_new_n2615_), .Y(_abc_15497_new_n2616_));
AND2X2 AND2X2_959 ( .A(_abc_15497_new_n2616_), .B(digest_update), .Y(_abc_15497_new_n2617_));
AND2X2 AND2X2_96 ( .A(_abc_15497_new_n879_), .B(_abc_15497_new_n877_), .Y(_abc_15497_new_n880_));
AND2X2 AND2X2_960 ( .A(_abc_15497_new_n2618_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n2619_));
AND2X2 AND2X2_961 ( .A(_abc_15497_new_n701_), .B(\digest[124] ), .Y(_abc_15497_new_n2621_));
AND2X2 AND2X2_962 ( .A(_abc_15497_new_n2609_), .B(_abc_15497_new_n2596_), .Y(_abc_15497_new_n2622_));
AND2X2 AND2X2_963 ( .A(_abc_15497_new_n2598_), .B(_abc_15497_new_n2612_), .Y(_abc_15497_new_n2624_));
AND2X2 AND2X2_964 ( .A(_abc_15497_new_n2594_), .B(_abc_15497_new_n2624_), .Y(_abc_15497_new_n2625_));
AND2X2 AND2X2_965 ( .A(\digest[124] ), .B(b_reg_28_), .Y(_abc_15497_new_n2628_));
AND2X2 AND2X2_966 ( .A(_abc_15497_new_n2629_), .B(_abc_15497_new_n2627_), .Y(_abc_15497_new_n2630_));
AND2X2 AND2X2_967 ( .A(_abc_15497_new_n2626_), .B(_abc_15497_new_n2630_), .Y(_abc_15497_new_n2632_));
AND2X2 AND2X2_968 ( .A(_abc_15497_new_n2633_), .B(_abc_15497_new_n2631_), .Y(_abc_15497_new_n2634_));
AND2X2 AND2X2_969 ( .A(_abc_15497_new_n2634_), .B(digest_update), .Y(_abc_15497_new_n2635_));
AND2X2 AND2X2_97 ( .A(_abc_15497_new_n880_), .B(digest_update), .Y(_abc_15497_new_n881_));
AND2X2 AND2X2_970 ( .A(\digest[125] ), .B(b_reg_29_), .Y(_abc_15497_new_n2642_));
AND2X2 AND2X2_971 ( .A(_abc_15497_new_n2643_), .B(_abc_15497_new_n2641_), .Y(_abc_15497_new_n2644_));
AND2X2 AND2X2_972 ( .A(_abc_15497_new_n2640_), .B(_abc_15497_new_n2644_), .Y(_abc_15497_new_n2645_));
AND2X2 AND2X2_973 ( .A(_abc_15497_new_n2639_), .B(_abc_15497_new_n2646_), .Y(_abc_15497_new_n2647_));
AND2X2 AND2X2_974 ( .A(_abc_15497_new_n2649_), .B(_abc_15497_new_n2638_), .Y(_0H1_reg_31_0__29_));
AND2X2 AND2X2_975 ( .A(\digest[126] ), .B(b_reg_30_), .Y(_abc_15497_new_n2652_));
AND2X2 AND2X2_976 ( .A(_abc_15497_new_n2653_), .B(_abc_15497_new_n2651_), .Y(_abc_15497_new_n2654_));
AND2X2 AND2X2_977 ( .A(_abc_15497_new_n2644_), .B(_abc_15497_new_n2628_), .Y(_abc_15497_new_n2655_));
AND2X2 AND2X2_978 ( .A(_abc_15497_new_n2630_), .B(_abc_15497_new_n2644_), .Y(_abc_15497_new_n2657_));
AND2X2 AND2X2_979 ( .A(_abc_15497_new_n2626_), .B(_abc_15497_new_n2657_), .Y(_abc_15497_new_n2658_));
AND2X2 AND2X2_98 ( .A(_abc_15497_new_n879_), .B(_abc_15497_new_n875_), .Y(_abc_15497_new_n883_));
AND2X2 AND2X2_980 ( .A(_abc_15497_new_n2667_), .B(_abc_15497_new_n2285_), .Y(_abc_15497_new_n2668_));
AND2X2 AND2X2_981 ( .A(_abc_15497_new_n2670_), .B(_abc_15497_new_n2665_), .Y(_abc_15497_new_n2671_));
AND2X2 AND2X2_982 ( .A(_abc_15497_new_n2673_), .B(_abc_15497_new_n2424_), .Y(_abc_15497_new_n2674_));
AND2X2 AND2X2_983 ( .A(_abc_15497_new_n2676_), .B(_abc_15497_new_n2664_), .Y(_abc_15497_new_n2677_));
AND2X2 AND2X2_984 ( .A(_abc_15497_new_n2679_), .B(_abc_15497_new_n2680_), .Y(_abc_15497_new_n2681_));
AND2X2 AND2X2_985 ( .A(_abc_15497_new_n2683_), .B(_abc_15497_new_n2663_), .Y(_abc_15497_new_n2684_));
AND2X2 AND2X2_986 ( .A(_abc_15497_new_n2686_), .B(_abc_15497_new_n2662_), .Y(_abc_15497_new_n2687_));
AND2X2 AND2X2_987 ( .A(_abc_15497_new_n2688_), .B(_abc_15497_new_n2660_), .Y(_abc_15497_new_n2689_));
AND2X2 AND2X2_988 ( .A(_abc_15497_new_n2689_), .B(digest_update), .Y(_abc_15497_new_n2690_));
AND2X2 AND2X2_989 ( .A(_abc_15497_new_n2691_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n2692_));
AND2X2 AND2X2_99 ( .A(\digest[91] ), .B(c_reg_27_), .Y(_abc_15497_new_n886_));
AND2X2 AND2X2_990 ( .A(_abc_15497_new_n2659_), .B(_abc_15497_new_n2654_), .Y(_abc_15497_new_n2694_));
AND2X2 AND2X2_991 ( .A(_abc_15497_new_n2697_), .B(_abc_15497_new_n2699_), .Y(_abc_15497_new_n2700_));
AND2X2 AND2X2_992 ( .A(_abc_15497_new_n2688_), .B(_abc_15497_new_n2653_), .Y(_abc_15497_new_n2703_));
AND2X2 AND2X2_993 ( .A(_abc_15497_new_n2704_), .B(_abc_15497_new_n2702_), .Y(_abc_15497_new_n2705_));
AND2X2 AND2X2_994 ( .A(_abc_15497_new_n2705_), .B(digest_update), .Y(_abc_15497_new_n2706_));
AND2X2 AND2X2_995 ( .A(_abc_15497_new_n2707_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n2708_));
AND2X2 AND2X2_996 ( .A(\digest[128] ), .B(a_reg_0_), .Y(_abc_15497_new_n2711_));
AND2X2 AND2X2_997 ( .A(_abc_15497_new_n2712_), .B(digest_update), .Y(_abc_15497_new_n2713_));
AND2X2 AND2X2_998 ( .A(_abc_15497_new_n2713_), .B(_abc_15497_new_n2710_), .Y(_abc_15497_new_n2714_));
AND2X2 AND2X2_999 ( .A(_abc_15497_new_n2715_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n2716_));
DFFSR DFFSR_1 ( .CLK(clk), .D(_0a_reg_31_0__0_), .Q(a_reg_0_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_10 ( .CLK(clk), .D(_0a_reg_31_0__9_), .Q(a_reg_9_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_100 ( .CLK(clk), .D(_0d_reg_31_0__3_), .Q(d_reg_3_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_101 ( .CLK(clk), .D(_0d_reg_31_0__4_), .Q(d_reg_4_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_102 ( .CLK(clk), .D(_0d_reg_31_0__5_), .Q(d_reg_5_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_103 ( .CLK(clk), .D(_0d_reg_31_0__6_), .Q(d_reg_6_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_104 ( .CLK(clk), .D(_0d_reg_31_0__7_), .Q(d_reg_7_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_105 ( .CLK(clk), .D(_0d_reg_31_0__8_), .Q(d_reg_8_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_106 ( .CLK(clk), .D(_0d_reg_31_0__9_), .Q(d_reg_9_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_107 ( .CLK(clk), .D(_0d_reg_31_0__10_), .Q(d_reg_10_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_108 ( .CLK(clk), .D(_0d_reg_31_0__11_), .Q(d_reg_11_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_109 ( .CLK(clk), .D(_0d_reg_31_0__12_), .Q(d_reg_12_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_11 ( .CLK(clk), .D(_0a_reg_31_0__10_), .Q(a_reg_10_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_110 ( .CLK(clk), .D(_0d_reg_31_0__13_), .Q(d_reg_13_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_111 ( .CLK(clk), .D(_0d_reg_31_0__14_), .Q(d_reg_14_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_112 ( .CLK(clk), .D(_0d_reg_31_0__15_), .Q(d_reg_15_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_113 ( .CLK(clk), .D(_0d_reg_31_0__16_), .Q(d_reg_16_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_114 ( .CLK(clk), .D(_0d_reg_31_0__17_), .Q(d_reg_17_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_115 ( .CLK(clk), .D(_0d_reg_31_0__18_), .Q(d_reg_18_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_116 ( .CLK(clk), .D(_0d_reg_31_0__19_), .Q(d_reg_19_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_117 ( .CLK(clk), .D(_0d_reg_31_0__20_), .Q(d_reg_20_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_118 ( .CLK(clk), .D(_0d_reg_31_0__21_), .Q(d_reg_21_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_119 ( .CLK(clk), .D(_0d_reg_31_0__22_), .Q(d_reg_22_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_12 ( .CLK(clk), .D(_0a_reg_31_0__11_), .Q(a_reg_11_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_120 ( .CLK(clk), .D(_0d_reg_31_0__23_), .Q(d_reg_23_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_121 ( .CLK(clk), .D(_0d_reg_31_0__24_), .Q(d_reg_24_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_122 ( .CLK(clk), .D(_0d_reg_31_0__25_), .Q(d_reg_25_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_123 ( .CLK(clk), .D(_0d_reg_31_0__26_), .Q(d_reg_26_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_124 ( .CLK(clk), .D(_0d_reg_31_0__27_), .Q(d_reg_27_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_125 ( .CLK(clk), .D(_0d_reg_31_0__28_), .Q(d_reg_28_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_126 ( .CLK(clk), .D(_0d_reg_31_0__29_), .Q(d_reg_29_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_127 ( .CLK(clk), .D(_0d_reg_31_0__30_), .Q(d_reg_30_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_128 ( .CLK(clk), .D(_0d_reg_31_0__31_), .Q(d_reg_31_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_129 ( .CLK(clk), .D(_0e_reg_31_0__0_), .Q(e_reg_0_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_13 ( .CLK(clk), .D(_0a_reg_31_0__12_), .Q(a_reg_12_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_130 ( .CLK(clk), .D(_0e_reg_31_0__1_), .Q(e_reg_1_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_131 ( .CLK(clk), .D(_0e_reg_31_0__2_), .Q(e_reg_2_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_132 ( .CLK(clk), .D(_0e_reg_31_0__3_), .Q(e_reg_3_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_133 ( .CLK(clk), .D(_0e_reg_31_0__4_), .Q(e_reg_4_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_134 ( .CLK(clk), .D(_0e_reg_31_0__5_), .Q(e_reg_5_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_135 ( .CLK(clk), .D(_0e_reg_31_0__6_), .Q(e_reg_6_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_136 ( .CLK(clk), .D(_0e_reg_31_0__7_), .Q(e_reg_7_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_137 ( .CLK(clk), .D(_0e_reg_31_0__8_), .Q(e_reg_8_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_138 ( .CLK(clk), .D(_0e_reg_31_0__9_), .Q(e_reg_9_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_139 ( .CLK(clk), .D(_0e_reg_31_0__10_), .Q(e_reg_10_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_14 ( .CLK(clk), .D(_0a_reg_31_0__13_), .Q(a_reg_13_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_140 ( .CLK(clk), .D(_0e_reg_31_0__11_), .Q(e_reg_11_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_141 ( .CLK(clk), .D(_0e_reg_31_0__12_), .Q(e_reg_12_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_142 ( .CLK(clk), .D(_0e_reg_31_0__13_), .Q(e_reg_13_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_143 ( .CLK(clk), .D(_0e_reg_31_0__14_), .Q(e_reg_14_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_144 ( .CLK(clk), .D(_0e_reg_31_0__15_), .Q(e_reg_15_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_145 ( .CLK(clk), .D(_0e_reg_31_0__16_), .Q(e_reg_16_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_146 ( .CLK(clk), .D(_0e_reg_31_0__17_), .Q(e_reg_17_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_147 ( .CLK(clk), .D(_0e_reg_31_0__18_), .Q(e_reg_18_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_148 ( .CLK(clk), .D(_0e_reg_31_0__19_), .Q(e_reg_19_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_149 ( .CLK(clk), .D(_0e_reg_31_0__20_), .Q(e_reg_20_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_15 ( .CLK(clk), .D(_0a_reg_31_0__14_), .Q(a_reg_14_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_150 ( .CLK(clk), .D(_0e_reg_31_0__21_), .Q(e_reg_21_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_151 ( .CLK(clk), .D(_0e_reg_31_0__22_), .Q(e_reg_22_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_152 ( .CLK(clk), .D(_0e_reg_31_0__23_), .Q(e_reg_23_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_153 ( .CLK(clk), .D(_0e_reg_31_0__24_), .Q(e_reg_24_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_154 ( .CLK(clk), .D(_0e_reg_31_0__25_), .Q(e_reg_25_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_155 ( .CLK(clk), .D(_0e_reg_31_0__26_), .Q(e_reg_26_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_156 ( .CLK(clk), .D(_0e_reg_31_0__27_), .Q(e_reg_27_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_157 ( .CLK(clk), .D(_0e_reg_31_0__28_), .Q(e_reg_28_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_158 ( .CLK(clk), .D(_0e_reg_31_0__29_), .Q(e_reg_29_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_159 ( .CLK(clk), .D(_0e_reg_31_0__30_), .Q(e_reg_30_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_16 ( .CLK(clk), .D(_0a_reg_31_0__15_), .Q(a_reg_15_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_160 ( .CLK(clk), .D(_0e_reg_31_0__31_), .Q(e_reg_31_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_161 ( .CLK(clk), .D(_0H0_reg_31_0__0_), .Q(\digest[128] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_162 ( .CLK(clk), .D(_0H0_reg_31_0__1_), .Q(\digest[129] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_163 ( .CLK(clk), .D(_0H0_reg_31_0__2_), .Q(\digest[130] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_164 ( .CLK(clk), .D(_0H0_reg_31_0__3_), .Q(\digest[131] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_165 ( .CLK(clk), .D(_0H0_reg_31_0__4_), .Q(\digest[132] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_166 ( .CLK(clk), .D(_0H0_reg_31_0__5_), .Q(\digest[133] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_167 ( .CLK(clk), .D(_0H0_reg_31_0__6_), .Q(\digest[134] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_168 ( .CLK(clk), .D(_0H0_reg_31_0__7_), .Q(\digest[135] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_169 ( .CLK(clk), .D(_0H0_reg_31_0__8_), .Q(\digest[136] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_17 ( .CLK(clk), .D(_0a_reg_31_0__16_), .Q(a_reg_16_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_170 ( .CLK(clk), .D(_0H0_reg_31_0__9_), .Q(\digest[137] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_171 ( .CLK(clk), .D(_0H0_reg_31_0__10_), .Q(\digest[138] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_172 ( .CLK(clk), .D(_0H0_reg_31_0__11_), .Q(\digest[139] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_173 ( .CLK(clk), .D(_0H0_reg_31_0__12_), .Q(\digest[140] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_174 ( .CLK(clk), .D(_0H0_reg_31_0__13_), .Q(\digest[141] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_175 ( .CLK(clk), .D(_0H0_reg_31_0__14_), .Q(\digest[142] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_176 ( .CLK(clk), .D(_0H0_reg_31_0__15_), .Q(\digest[143] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_177 ( .CLK(clk), .D(_0H0_reg_31_0__16_), .Q(\digest[144] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_178 ( .CLK(clk), .D(_0H0_reg_31_0__17_), .Q(\digest[145] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_179 ( .CLK(clk), .D(_0H0_reg_31_0__18_), .Q(\digest[146] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_18 ( .CLK(clk), .D(_0a_reg_31_0__17_), .Q(a_reg_17_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_180 ( .CLK(clk), .D(_0H0_reg_31_0__19_), .Q(\digest[147] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_181 ( .CLK(clk), .D(_0H0_reg_31_0__20_), .Q(\digest[148] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_182 ( .CLK(clk), .D(_0H0_reg_31_0__21_), .Q(\digest[149] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_183 ( .CLK(clk), .D(_0H0_reg_31_0__22_), .Q(\digest[150] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_184 ( .CLK(clk), .D(_0H0_reg_31_0__23_), .Q(\digest[151] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_185 ( .CLK(clk), .D(_0H0_reg_31_0__24_), .Q(\digest[152] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_186 ( .CLK(clk), .D(_0H0_reg_31_0__25_), .Q(\digest[153] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_187 ( .CLK(clk), .D(_0H0_reg_31_0__26_), .Q(\digest[154] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_188 ( .CLK(clk), .D(_0H0_reg_31_0__27_), .Q(\digest[155] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_189 ( .CLK(clk), .D(_0H0_reg_31_0__28_), .Q(\digest[156] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_19 ( .CLK(clk), .D(_0a_reg_31_0__18_), .Q(a_reg_18_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_190 ( .CLK(clk), .D(_0H0_reg_31_0__29_), .Q(\digest[157] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_191 ( .CLK(clk), .D(_0H0_reg_31_0__30_), .Q(\digest[158] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_192 ( .CLK(clk), .D(_0H0_reg_31_0__31_), .Q(\digest[159] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_193 ( .CLK(clk), .D(_0H1_reg_31_0__0_), .Q(\digest[96] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_194 ( .CLK(clk), .D(_0H1_reg_31_0__1_), .Q(\digest[97] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_195 ( .CLK(clk), .D(_0H1_reg_31_0__2_), .Q(\digest[98] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_196 ( .CLK(clk), .D(_0H1_reg_31_0__3_), .Q(\digest[99] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_197 ( .CLK(clk), .D(_0H1_reg_31_0__4_), .Q(\digest[100] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_198 ( .CLK(clk), .D(_0H1_reg_31_0__5_), .Q(\digest[101] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_199 ( .CLK(clk), .D(_0H1_reg_31_0__6_), .Q(\digest[102] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_2 ( .CLK(clk), .D(_0a_reg_31_0__1_), .Q(a_reg_1_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_20 ( .CLK(clk), .D(_0a_reg_31_0__19_), .Q(a_reg_19_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_200 ( .CLK(clk), .D(_0H1_reg_31_0__7_), .Q(\digest[103] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_201 ( .CLK(clk), .D(_0H1_reg_31_0__8_), .Q(\digest[104] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_202 ( .CLK(clk), .D(_0H1_reg_31_0__9_), .Q(\digest[105] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_203 ( .CLK(clk), .D(_0H1_reg_31_0__10_), .Q(\digest[106] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_204 ( .CLK(clk), .D(_0H1_reg_31_0__11_), .Q(\digest[107] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_205 ( .CLK(clk), .D(_0H1_reg_31_0__12_), .Q(\digest[108] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_206 ( .CLK(clk), .D(_0H1_reg_31_0__13_), .Q(\digest[109] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_207 ( .CLK(clk), .D(_0H1_reg_31_0__14_), .Q(\digest[110] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_208 ( .CLK(clk), .D(_0H1_reg_31_0__15_), .Q(\digest[111] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_209 ( .CLK(clk), .D(_0H1_reg_31_0__16_), .Q(\digest[112] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_21 ( .CLK(clk), .D(_0a_reg_31_0__20_), .Q(a_reg_20_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_210 ( .CLK(clk), .D(_0H1_reg_31_0__17_), .Q(\digest[113] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_211 ( .CLK(clk), .D(_0H1_reg_31_0__18_), .Q(\digest[114] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_212 ( .CLK(clk), .D(_0H1_reg_31_0__19_), .Q(\digest[115] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_213 ( .CLK(clk), .D(_0H1_reg_31_0__20_), .Q(\digest[116] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_214 ( .CLK(clk), .D(_0H1_reg_31_0__21_), .Q(\digest[117] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_215 ( .CLK(clk), .D(_0H1_reg_31_0__22_), .Q(\digest[118] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_216 ( .CLK(clk), .D(_0H1_reg_31_0__23_), .Q(\digest[119] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_217 ( .CLK(clk), .D(_0H1_reg_31_0__24_), .Q(\digest[120] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_218 ( .CLK(clk), .D(_0H1_reg_31_0__25_), .Q(\digest[121] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_219 ( .CLK(clk), .D(_0H1_reg_31_0__26_), .Q(\digest[122] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_22 ( .CLK(clk), .D(_0a_reg_31_0__21_), .Q(a_reg_21_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_220 ( .CLK(clk), .D(_0H1_reg_31_0__27_), .Q(\digest[123] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_221 ( .CLK(clk), .D(_0H1_reg_31_0__28_), .Q(\digest[124] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_222 ( .CLK(clk), .D(_0H1_reg_31_0__29_), .Q(\digest[125] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_223 ( .CLK(clk), .D(_0H1_reg_31_0__30_), .Q(\digest[126] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_224 ( .CLK(clk), .D(_0H1_reg_31_0__31_), .Q(\digest[127] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_225 ( .CLK(clk), .D(_0H2_reg_31_0__0_), .Q(\digest[64] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_226 ( .CLK(clk), .D(_0H2_reg_31_0__1_), .Q(\digest[65] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_227 ( .CLK(clk), .D(_0H2_reg_31_0__2_), .Q(\digest[66] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_228 ( .CLK(clk), .D(_0H2_reg_31_0__3_), .Q(\digest[67] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_229 ( .CLK(clk), .D(_0H2_reg_31_0__4_), .Q(\digest[68] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_23 ( .CLK(clk), .D(_0a_reg_31_0__22_), .Q(a_reg_22_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_230 ( .CLK(clk), .D(_0H2_reg_31_0__5_), .Q(\digest[69] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_231 ( .CLK(clk), .D(_0H2_reg_31_0__6_), .Q(\digest[70] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_232 ( .CLK(clk), .D(_0H2_reg_31_0__7_), .Q(\digest[71] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_233 ( .CLK(clk), .D(_0H2_reg_31_0__8_), .Q(\digest[72] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_234 ( .CLK(clk), .D(_0H2_reg_31_0__9_), .Q(\digest[73] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_235 ( .CLK(clk), .D(_0H2_reg_31_0__10_), .Q(\digest[74] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_236 ( .CLK(clk), .D(_0H2_reg_31_0__11_), .Q(\digest[75] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_237 ( .CLK(clk), .D(_0H2_reg_31_0__12_), .Q(\digest[76] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_238 ( .CLK(clk), .D(_0H2_reg_31_0__13_), .Q(\digest[77] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_239 ( .CLK(clk), .D(_0H2_reg_31_0__14_), .Q(\digest[78] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_24 ( .CLK(clk), .D(_0a_reg_31_0__23_), .Q(a_reg_23_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_240 ( .CLK(clk), .D(_0H2_reg_31_0__15_), .Q(\digest[79] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_241 ( .CLK(clk), .D(_0H2_reg_31_0__16_), .Q(\digest[80] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_242 ( .CLK(clk), .D(_0H2_reg_31_0__17_), .Q(\digest[81] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_243 ( .CLK(clk), .D(_0H2_reg_31_0__18_), .Q(\digest[82] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_244 ( .CLK(clk), .D(_0H2_reg_31_0__19_), .Q(\digest[83] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_245 ( .CLK(clk), .D(_0H2_reg_31_0__20_), .Q(\digest[84] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_246 ( .CLK(clk), .D(_0H2_reg_31_0__21_), .Q(\digest[85] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_247 ( .CLK(clk), .D(_0H2_reg_31_0__22_), .Q(\digest[86] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_248 ( .CLK(clk), .D(_0H2_reg_31_0__23_), .Q(\digest[87] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_249 ( .CLK(clk), .D(_0H2_reg_31_0__24_), .Q(\digest[88] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_25 ( .CLK(clk), .D(_0a_reg_31_0__24_), .Q(a_reg_24_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_250 ( .CLK(clk), .D(_0H2_reg_31_0__25_), .Q(\digest[89] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_251 ( .CLK(clk), .D(_0H2_reg_31_0__26_), .Q(\digest[90] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_252 ( .CLK(clk), .D(_0H2_reg_31_0__27_), .Q(\digest[91] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_253 ( .CLK(clk), .D(_0H2_reg_31_0__28_), .Q(\digest[92] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_254 ( .CLK(clk), .D(_0H2_reg_31_0__29_), .Q(\digest[93] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_255 ( .CLK(clk), .D(_0H2_reg_31_0__30_), .Q(\digest[94] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_256 ( .CLK(clk), .D(_0H2_reg_31_0__31_), .Q(\digest[95] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_257 ( .CLK(clk), .D(_0H3_reg_31_0__0_), .Q(\digest[32] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_258 ( .CLK(clk), .D(_0H3_reg_31_0__1_), .Q(\digest[33] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_259 ( .CLK(clk), .D(_0H3_reg_31_0__2_), .Q(\digest[34] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_26 ( .CLK(clk), .D(_0a_reg_31_0__25_), .Q(a_reg_25_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_260 ( .CLK(clk), .D(_0H3_reg_31_0__3_), .Q(\digest[35] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_261 ( .CLK(clk), .D(_0H3_reg_31_0__4_), .Q(\digest[36] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_262 ( .CLK(clk), .D(_0H3_reg_31_0__5_), .Q(\digest[37] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_263 ( .CLK(clk), .D(_0H3_reg_31_0__6_), .Q(\digest[38] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_264 ( .CLK(clk), .D(_0H3_reg_31_0__7_), .Q(\digest[39] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_265 ( .CLK(clk), .D(_0H3_reg_31_0__8_), .Q(\digest[40] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_266 ( .CLK(clk), .D(_0H3_reg_31_0__9_), .Q(\digest[41] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_267 ( .CLK(clk), .D(_0H3_reg_31_0__10_), .Q(\digest[42] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_268 ( .CLK(clk), .D(_0H3_reg_31_0__11_), .Q(\digest[43] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_269 ( .CLK(clk), .D(_0H3_reg_31_0__12_), .Q(\digest[44] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_27 ( .CLK(clk), .D(_0a_reg_31_0__26_), .Q(a_reg_26_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_270 ( .CLK(clk), .D(_0H3_reg_31_0__13_), .Q(\digest[45] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_271 ( .CLK(clk), .D(_0H3_reg_31_0__14_), .Q(\digest[46] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_272 ( .CLK(clk), .D(_0H3_reg_31_0__15_), .Q(\digest[47] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_273 ( .CLK(clk), .D(_0H3_reg_31_0__16_), .Q(\digest[48] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_274 ( .CLK(clk), .D(_0H3_reg_31_0__17_), .Q(\digest[49] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_275 ( .CLK(clk), .D(_0H3_reg_31_0__18_), .Q(\digest[50] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_276 ( .CLK(clk), .D(_0H3_reg_31_0__19_), .Q(\digest[51] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_277 ( .CLK(clk), .D(_0H3_reg_31_0__20_), .Q(\digest[52] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_278 ( .CLK(clk), .D(_0H3_reg_31_0__21_), .Q(\digest[53] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_279 ( .CLK(clk), .D(_0H3_reg_31_0__22_), .Q(\digest[54] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_28 ( .CLK(clk), .D(_0a_reg_31_0__27_), .Q(a_reg_27_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_280 ( .CLK(clk), .D(_0H3_reg_31_0__23_), .Q(\digest[55] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_281 ( .CLK(clk), .D(_0H3_reg_31_0__24_), .Q(\digest[56] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_282 ( .CLK(clk), .D(_0H3_reg_31_0__25_), .Q(\digest[57] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_283 ( .CLK(clk), .D(_0H3_reg_31_0__26_), .Q(\digest[58] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_284 ( .CLK(clk), .D(_0H3_reg_31_0__27_), .Q(\digest[59] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_285 ( .CLK(clk), .D(_0H3_reg_31_0__28_), .Q(\digest[60] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_286 ( .CLK(clk), .D(_0H3_reg_31_0__29_), .Q(\digest[61] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_287 ( .CLK(clk), .D(_0H3_reg_31_0__30_), .Q(\digest[62] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_288 ( .CLK(clk), .D(_0H3_reg_31_0__31_), .Q(\digest[63] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_289 ( .CLK(clk), .D(_0H4_reg_31_0__0_), .Q(\digest[0] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_29 ( .CLK(clk), .D(_0a_reg_31_0__28_), .Q(a_reg_28_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_290 ( .CLK(clk), .D(_0H4_reg_31_0__1_), .Q(\digest[1] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_291 ( .CLK(clk), .D(_0H4_reg_31_0__2_), .Q(\digest[2] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_292 ( .CLK(clk), .D(_0H4_reg_31_0__3_), .Q(\digest[3] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_293 ( .CLK(clk), .D(_0H4_reg_31_0__4_), .Q(\digest[4] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_294 ( .CLK(clk), .D(_0H4_reg_31_0__5_), .Q(\digest[5] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_295 ( .CLK(clk), .D(_0H4_reg_31_0__6_), .Q(\digest[6] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_296 ( .CLK(clk), .D(_0H4_reg_31_0__7_), .Q(\digest[7] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_297 ( .CLK(clk), .D(_0H4_reg_31_0__8_), .Q(\digest[8] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_298 ( .CLK(clk), .D(_0H4_reg_31_0__9_), .Q(\digest[9] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_299 ( .CLK(clk), .D(_0H4_reg_31_0__10_), .Q(\digest[10] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_3 ( .CLK(clk), .D(_0a_reg_31_0__2_), .Q(a_reg_2_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_30 ( .CLK(clk), .D(_0a_reg_31_0__29_), .Q(a_reg_29_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_300 ( .CLK(clk), .D(_0H4_reg_31_0__11_), .Q(\digest[11] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_301 ( .CLK(clk), .D(_0H4_reg_31_0__12_), .Q(\digest[12] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_302 ( .CLK(clk), .D(_0H4_reg_31_0__13_), .Q(\digest[13] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_303 ( .CLK(clk), .D(_0H4_reg_31_0__14_), .Q(\digest[14] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_304 ( .CLK(clk), .D(_0H4_reg_31_0__15_), .Q(\digest[15] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_305 ( .CLK(clk), .D(_0H4_reg_31_0__16_), .Q(\digest[16] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_306 ( .CLK(clk), .D(_0H4_reg_31_0__17_), .Q(\digest[17] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_307 ( .CLK(clk), .D(_0H4_reg_31_0__18_), .Q(\digest[18] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_308 ( .CLK(clk), .D(_0H4_reg_31_0__19_), .Q(\digest[19] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_309 ( .CLK(clk), .D(_0H4_reg_31_0__20_), .Q(\digest[20] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_31 ( .CLK(clk), .D(_0a_reg_31_0__30_), .Q(a_reg_30_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_310 ( .CLK(clk), .D(_0H4_reg_31_0__21_), .Q(\digest[21] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_311 ( .CLK(clk), .D(_0H4_reg_31_0__22_), .Q(\digest[22] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_312 ( .CLK(clk), .D(_0H4_reg_31_0__23_), .Q(\digest[23] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_313 ( .CLK(clk), .D(_0H4_reg_31_0__24_), .Q(\digest[24] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_314 ( .CLK(clk), .D(_0H4_reg_31_0__25_), .Q(\digest[25] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_315 ( .CLK(clk), .D(_0H4_reg_31_0__26_), .Q(\digest[26] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_316 ( .CLK(clk), .D(_0H4_reg_31_0__27_), .Q(\digest[27] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_317 ( .CLK(clk), .D(_0H4_reg_31_0__28_), .Q(\digest[28] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_318 ( .CLK(clk), .D(_0H4_reg_31_0__29_), .Q(\digest[29] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_319 ( .CLK(clk), .D(_0H4_reg_31_0__30_), .Q(\digest[30] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_32 ( .CLK(clk), .D(_0a_reg_31_0__31_), .Q(a_reg_31_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_320 ( .CLK(clk), .D(_0H4_reg_31_0__31_), .Q(\digest[31] ), .R(reset_n), .S(1'h1));
DFFSR DFFSR_321 ( .CLK(clk), .D(_0round_ctr_reg_6_0__0_), .Q(round_ctr_reg_0_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_322 ( .CLK(clk), .D(_0round_ctr_reg_6_0__1_), .Q(round_ctr_reg_1_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_323 ( .CLK(clk), .D(_0round_ctr_reg_6_0__2_), .Q(round_ctr_reg_2_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_324 ( .CLK(clk), .D(_0round_ctr_reg_6_0__3_), .Q(round_ctr_reg_3_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_325 ( .CLK(clk), .D(_0round_ctr_reg_6_0__4_), .Q(round_ctr_reg_4_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_326 ( .CLK(clk), .D(_0round_ctr_reg_6_0__5_), .Q(round_ctr_reg_5_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_327 ( .CLK(clk), .D(_0round_ctr_reg_6_0__6_), .Q(round_ctr_reg_6_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_328 ( .CLK(clk), .D(_0digest_valid_reg_0_0_), .Q(digest_valid), .R(reset_n), .S(1'h1));
DFFSR DFFSR_329 ( .CLK(clk), .D(_abc_15497_abc_9717_auto_fsm_map_cc_170_map_fsm_844_0_), .Q(ready), .R(1'h1), .S(reset_n));
DFFSR DFFSR_33 ( .CLK(clk), .D(_0b_reg_31_0__0_), .Q(b_reg_0_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_330 ( .CLK(clk), .D(_abc_15497_abc_9717_auto_fsm_map_cc_118_implement_pattern_cache_863), .Q(digest_update), .R(reset_n), .S(1'h1));
DFFSR DFFSR_331 ( .CLK(clk), .D(_abc_15497_abc_9717_auto_fsm_map_cc_170_map_fsm_844_2_), .Q(round_ctr_inc), .R(reset_n), .S(1'h1));
DFFSR DFFSR_332 ( .CLK(clk), .D(w_mem_inst__0w_ctr_reg_6_0__0_), .Q(w_mem_inst_w_ctr_reg_0_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_333 ( .CLK(clk), .D(w_mem_inst__0w_ctr_reg_6_0__1_), .Q(w_mem_inst_w_ctr_reg_1_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_334 ( .CLK(clk), .D(w_mem_inst__0w_ctr_reg_6_0__2_), .Q(w_mem_inst_w_ctr_reg_2_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_335 ( .CLK(clk), .D(w_mem_inst__0w_ctr_reg_6_0__3_), .Q(w_mem_inst_w_ctr_reg_3_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_336 ( .CLK(clk), .D(w_mem_inst__0w_ctr_reg_6_0__4_), .Q(w_mem_inst_w_ctr_reg_4_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_337 ( .CLK(clk), .D(w_mem_inst__0w_ctr_reg_6_0__5_), .Q(w_mem_inst_w_ctr_reg_5_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_338 ( .CLK(clk), .D(w_mem_inst__0w_ctr_reg_6_0__6_), .Q(w_mem_inst_w_ctr_reg_6_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_339 ( .CLK(clk), .D(w_mem_inst__0w_mem_0__31_0__0_), .Q(w_mem_inst_w_mem_0__0_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_34 ( .CLK(clk), .D(_0b_reg_31_0__1_), .Q(b_reg_1_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_340 ( .CLK(clk), .D(w_mem_inst__0w_mem_0__31_0__1_), .Q(w_mem_inst_w_mem_0__1_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_341 ( .CLK(clk), .D(w_mem_inst__0w_mem_0__31_0__2_), .Q(w_mem_inst_w_mem_0__2_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_342 ( .CLK(clk), .D(w_mem_inst__0w_mem_0__31_0__3_), .Q(w_mem_inst_w_mem_0__3_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_343 ( .CLK(clk), .D(w_mem_inst__0w_mem_0__31_0__4_), .Q(w_mem_inst_w_mem_0__4_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_344 ( .CLK(clk), .D(w_mem_inst__0w_mem_0__31_0__5_), .Q(w_mem_inst_w_mem_0__5_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_345 ( .CLK(clk), .D(w_mem_inst__0w_mem_0__31_0__6_), .Q(w_mem_inst_w_mem_0__6_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_346 ( .CLK(clk), .D(w_mem_inst__0w_mem_0__31_0__7_), .Q(w_mem_inst_w_mem_0__7_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_347 ( .CLK(clk), .D(w_mem_inst__0w_mem_0__31_0__8_), .Q(w_mem_inst_w_mem_0__8_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_348 ( .CLK(clk), .D(w_mem_inst__0w_mem_0__31_0__9_), .Q(w_mem_inst_w_mem_0__9_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_349 ( .CLK(clk), .D(w_mem_inst__0w_mem_0__31_0__10_), .Q(w_mem_inst_w_mem_0__10_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_35 ( .CLK(clk), .D(_0b_reg_31_0__2_), .Q(b_reg_2_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_350 ( .CLK(clk), .D(w_mem_inst__0w_mem_0__31_0__11_), .Q(w_mem_inst_w_mem_0__11_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_351 ( .CLK(clk), .D(w_mem_inst__0w_mem_0__31_0__12_), .Q(w_mem_inst_w_mem_0__12_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_352 ( .CLK(clk), .D(w_mem_inst__0w_mem_0__31_0__13_), .Q(w_mem_inst_w_mem_0__13_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_353 ( .CLK(clk), .D(w_mem_inst__0w_mem_0__31_0__14_), .Q(w_mem_inst_w_mem_0__14_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_354 ( .CLK(clk), .D(w_mem_inst__0w_mem_0__31_0__15_), .Q(w_mem_inst_w_mem_0__15_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_355 ( .CLK(clk), .D(w_mem_inst__0w_mem_0__31_0__16_), .Q(w_mem_inst_w_mem_0__16_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_356 ( .CLK(clk), .D(w_mem_inst__0w_mem_0__31_0__17_), .Q(w_mem_inst_w_mem_0__17_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_357 ( .CLK(clk), .D(w_mem_inst__0w_mem_0__31_0__18_), .Q(w_mem_inst_w_mem_0__18_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_358 ( .CLK(clk), .D(w_mem_inst__0w_mem_0__31_0__19_), .Q(w_mem_inst_w_mem_0__19_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_359 ( .CLK(clk), .D(w_mem_inst__0w_mem_0__31_0__20_), .Q(w_mem_inst_w_mem_0__20_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_36 ( .CLK(clk), .D(_0b_reg_31_0__3_), .Q(b_reg_3_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_360 ( .CLK(clk), .D(w_mem_inst__0w_mem_0__31_0__21_), .Q(w_mem_inst_w_mem_0__21_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_361 ( .CLK(clk), .D(w_mem_inst__0w_mem_0__31_0__22_), .Q(w_mem_inst_w_mem_0__22_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_362 ( .CLK(clk), .D(w_mem_inst__0w_mem_0__31_0__23_), .Q(w_mem_inst_w_mem_0__23_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_363 ( .CLK(clk), .D(w_mem_inst__0w_mem_0__31_0__24_), .Q(w_mem_inst_w_mem_0__24_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_364 ( .CLK(clk), .D(w_mem_inst__0w_mem_0__31_0__25_), .Q(w_mem_inst_w_mem_0__25_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_365 ( .CLK(clk), .D(w_mem_inst__0w_mem_0__31_0__26_), .Q(w_mem_inst_w_mem_0__26_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_366 ( .CLK(clk), .D(w_mem_inst__0w_mem_0__31_0__27_), .Q(w_mem_inst_w_mem_0__27_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_367 ( .CLK(clk), .D(w_mem_inst__0w_mem_0__31_0__28_), .Q(w_mem_inst_w_mem_0__28_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_368 ( .CLK(clk), .D(w_mem_inst__0w_mem_0__31_0__29_), .Q(w_mem_inst_w_mem_0__29_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_369 ( .CLK(clk), .D(w_mem_inst__0w_mem_0__31_0__30_), .Q(w_mem_inst_w_mem_0__30_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_37 ( .CLK(clk), .D(_0b_reg_31_0__4_), .Q(b_reg_4_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_370 ( .CLK(clk), .D(w_mem_inst__0w_mem_0__31_0__31_), .Q(w_mem_inst_w_mem_0__31_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_371 ( .CLK(clk), .D(w_mem_inst__0w_mem_1__31_0__0_), .Q(w_mem_inst_w_mem_1__0_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_372 ( .CLK(clk), .D(w_mem_inst__0w_mem_1__31_0__1_), .Q(w_mem_inst_w_mem_1__1_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_373 ( .CLK(clk), .D(w_mem_inst__0w_mem_1__31_0__2_), .Q(w_mem_inst_w_mem_1__2_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_374 ( .CLK(clk), .D(w_mem_inst__0w_mem_1__31_0__3_), .Q(w_mem_inst_w_mem_1__3_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_375 ( .CLK(clk), .D(w_mem_inst__0w_mem_1__31_0__4_), .Q(w_mem_inst_w_mem_1__4_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_376 ( .CLK(clk), .D(w_mem_inst__0w_mem_1__31_0__5_), .Q(w_mem_inst_w_mem_1__5_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_377 ( .CLK(clk), .D(w_mem_inst__0w_mem_1__31_0__6_), .Q(w_mem_inst_w_mem_1__6_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_378 ( .CLK(clk), .D(w_mem_inst__0w_mem_1__31_0__7_), .Q(w_mem_inst_w_mem_1__7_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_379 ( .CLK(clk), .D(w_mem_inst__0w_mem_1__31_0__8_), .Q(w_mem_inst_w_mem_1__8_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_38 ( .CLK(clk), .D(_0b_reg_31_0__5_), .Q(b_reg_5_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_380 ( .CLK(clk), .D(w_mem_inst__0w_mem_1__31_0__9_), .Q(w_mem_inst_w_mem_1__9_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_381 ( .CLK(clk), .D(w_mem_inst__0w_mem_1__31_0__10_), .Q(w_mem_inst_w_mem_1__10_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_382 ( .CLK(clk), .D(w_mem_inst__0w_mem_1__31_0__11_), .Q(w_mem_inst_w_mem_1__11_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_383 ( .CLK(clk), .D(w_mem_inst__0w_mem_1__31_0__12_), .Q(w_mem_inst_w_mem_1__12_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_384 ( .CLK(clk), .D(w_mem_inst__0w_mem_1__31_0__13_), .Q(w_mem_inst_w_mem_1__13_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_385 ( .CLK(clk), .D(w_mem_inst__0w_mem_1__31_0__14_), .Q(w_mem_inst_w_mem_1__14_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_386 ( .CLK(clk), .D(w_mem_inst__0w_mem_1__31_0__15_), .Q(w_mem_inst_w_mem_1__15_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_387 ( .CLK(clk), .D(w_mem_inst__0w_mem_1__31_0__16_), .Q(w_mem_inst_w_mem_1__16_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_388 ( .CLK(clk), .D(w_mem_inst__0w_mem_1__31_0__17_), .Q(w_mem_inst_w_mem_1__17_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_389 ( .CLK(clk), .D(w_mem_inst__0w_mem_1__31_0__18_), .Q(w_mem_inst_w_mem_1__18_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_39 ( .CLK(clk), .D(_0b_reg_31_0__6_), .Q(b_reg_6_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_390 ( .CLK(clk), .D(w_mem_inst__0w_mem_1__31_0__19_), .Q(w_mem_inst_w_mem_1__19_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_391 ( .CLK(clk), .D(w_mem_inst__0w_mem_1__31_0__20_), .Q(w_mem_inst_w_mem_1__20_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_392 ( .CLK(clk), .D(w_mem_inst__0w_mem_1__31_0__21_), .Q(w_mem_inst_w_mem_1__21_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_393 ( .CLK(clk), .D(w_mem_inst__0w_mem_1__31_0__22_), .Q(w_mem_inst_w_mem_1__22_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_394 ( .CLK(clk), .D(w_mem_inst__0w_mem_1__31_0__23_), .Q(w_mem_inst_w_mem_1__23_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_395 ( .CLK(clk), .D(w_mem_inst__0w_mem_1__31_0__24_), .Q(w_mem_inst_w_mem_1__24_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_396 ( .CLK(clk), .D(w_mem_inst__0w_mem_1__31_0__25_), .Q(w_mem_inst_w_mem_1__25_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_397 ( .CLK(clk), .D(w_mem_inst__0w_mem_1__31_0__26_), .Q(w_mem_inst_w_mem_1__26_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_398 ( .CLK(clk), .D(w_mem_inst__0w_mem_1__31_0__27_), .Q(w_mem_inst_w_mem_1__27_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_399 ( .CLK(clk), .D(w_mem_inst__0w_mem_1__31_0__28_), .Q(w_mem_inst_w_mem_1__28_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_4 ( .CLK(clk), .D(_0a_reg_31_0__3_), .Q(a_reg_3_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_40 ( .CLK(clk), .D(_0b_reg_31_0__7_), .Q(b_reg_7_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_400 ( .CLK(clk), .D(w_mem_inst__0w_mem_1__31_0__29_), .Q(w_mem_inst_w_mem_1__29_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_401 ( .CLK(clk), .D(w_mem_inst__0w_mem_1__31_0__30_), .Q(w_mem_inst_w_mem_1__30_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_402 ( .CLK(clk), .D(w_mem_inst__0w_mem_1__31_0__31_), .Q(w_mem_inst_w_mem_1__31_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_403 ( .CLK(clk), .D(w_mem_inst__0w_mem_2__31_0__0_), .Q(w_mem_inst_w_mem_2__0_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_404 ( .CLK(clk), .D(w_mem_inst__0w_mem_2__31_0__1_), .Q(w_mem_inst_w_mem_2__1_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_405 ( .CLK(clk), .D(w_mem_inst__0w_mem_2__31_0__2_), .Q(w_mem_inst_w_mem_2__2_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_406 ( .CLK(clk), .D(w_mem_inst__0w_mem_2__31_0__3_), .Q(w_mem_inst_w_mem_2__3_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_407 ( .CLK(clk), .D(w_mem_inst__0w_mem_2__31_0__4_), .Q(w_mem_inst_w_mem_2__4_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_408 ( .CLK(clk), .D(w_mem_inst__0w_mem_2__31_0__5_), .Q(w_mem_inst_w_mem_2__5_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_409 ( .CLK(clk), .D(w_mem_inst__0w_mem_2__31_0__6_), .Q(w_mem_inst_w_mem_2__6_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_41 ( .CLK(clk), .D(_0b_reg_31_0__8_), .Q(b_reg_8_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_410 ( .CLK(clk), .D(w_mem_inst__0w_mem_2__31_0__7_), .Q(w_mem_inst_w_mem_2__7_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_411 ( .CLK(clk), .D(w_mem_inst__0w_mem_2__31_0__8_), .Q(w_mem_inst_w_mem_2__8_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_412 ( .CLK(clk), .D(w_mem_inst__0w_mem_2__31_0__9_), .Q(w_mem_inst_w_mem_2__9_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_413 ( .CLK(clk), .D(w_mem_inst__0w_mem_2__31_0__10_), .Q(w_mem_inst_w_mem_2__10_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_414 ( .CLK(clk), .D(w_mem_inst__0w_mem_2__31_0__11_), .Q(w_mem_inst_w_mem_2__11_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_415 ( .CLK(clk), .D(w_mem_inst__0w_mem_2__31_0__12_), .Q(w_mem_inst_w_mem_2__12_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_416 ( .CLK(clk), .D(w_mem_inst__0w_mem_2__31_0__13_), .Q(w_mem_inst_w_mem_2__13_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_417 ( .CLK(clk), .D(w_mem_inst__0w_mem_2__31_0__14_), .Q(w_mem_inst_w_mem_2__14_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_418 ( .CLK(clk), .D(w_mem_inst__0w_mem_2__31_0__15_), .Q(w_mem_inst_w_mem_2__15_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_419 ( .CLK(clk), .D(w_mem_inst__0w_mem_2__31_0__16_), .Q(w_mem_inst_w_mem_2__16_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_42 ( .CLK(clk), .D(_0b_reg_31_0__9_), .Q(b_reg_9_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_420 ( .CLK(clk), .D(w_mem_inst__0w_mem_2__31_0__17_), .Q(w_mem_inst_w_mem_2__17_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_421 ( .CLK(clk), .D(w_mem_inst__0w_mem_2__31_0__18_), .Q(w_mem_inst_w_mem_2__18_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_422 ( .CLK(clk), .D(w_mem_inst__0w_mem_2__31_0__19_), .Q(w_mem_inst_w_mem_2__19_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_423 ( .CLK(clk), .D(w_mem_inst__0w_mem_2__31_0__20_), .Q(w_mem_inst_w_mem_2__20_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_424 ( .CLK(clk), .D(w_mem_inst__0w_mem_2__31_0__21_), .Q(w_mem_inst_w_mem_2__21_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_425 ( .CLK(clk), .D(w_mem_inst__0w_mem_2__31_0__22_), .Q(w_mem_inst_w_mem_2__22_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_426 ( .CLK(clk), .D(w_mem_inst__0w_mem_2__31_0__23_), .Q(w_mem_inst_w_mem_2__23_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_427 ( .CLK(clk), .D(w_mem_inst__0w_mem_2__31_0__24_), .Q(w_mem_inst_w_mem_2__24_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_428 ( .CLK(clk), .D(w_mem_inst__0w_mem_2__31_0__25_), .Q(w_mem_inst_w_mem_2__25_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_429 ( .CLK(clk), .D(w_mem_inst__0w_mem_2__31_0__26_), .Q(w_mem_inst_w_mem_2__26_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_43 ( .CLK(clk), .D(_0b_reg_31_0__10_), .Q(b_reg_10_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_430 ( .CLK(clk), .D(w_mem_inst__0w_mem_2__31_0__27_), .Q(w_mem_inst_w_mem_2__27_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_431 ( .CLK(clk), .D(w_mem_inst__0w_mem_2__31_0__28_), .Q(w_mem_inst_w_mem_2__28_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_432 ( .CLK(clk), .D(w_mem_inst__0w_mem_2__31_0__29_), .Q(w_mem_inst_w_mem_2__29_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_433 ( .CLK(clk), .D(w_mem_inst__0w_mem_2__31_0__30_), .Q(w_mem_inst_w_mem_2__30_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_434 ( .CLK(clk), .D(w_mem_inst__0w_mem_2__31_0__31_), .Q(w_mem_inst_w_mem_2__31_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_435 ( .CLK(clk), .D(w_mem_inst__0w_mem_3__31_0__0_), .Q(w_mem_inst_w_mem_3__0_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_436 ( .CLK(clk), .D(w_mem_inst__0w_mem_3__31_0__1_), .Q(w_mem_inst_w_mem_3__1_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_437 ( .CLK(clk), .D(w_mem_inst__0w_mem_3__31_0__2_), .Q(w_mem_inst_w_mem_3__2_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_438 ( .CLK(clk), .D(w_mem_inst__0w_mem_3__31_0__3_), .Q(w_mem_inst_w_mem_3__3_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_439 ( .CLK(clk), .D(w_mem_inst__0w_mem_3__31_0__4_), .Q(w_mem_inst_w_mem_3__4_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_44 ( .CLK(clk), .D(_0b_reg_31_0__11_), .Q(b_reg_11_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_440 ( .CLK(clk), .D(w_mem_inst__0w_mem_3__31_0__5_), .Q(w_mem_inst_w_mem_3__5_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_441 ( .CLK(clk), .D(w_mem_inst__0w_mem_3__31_0__6_), .Q(w_mem_inst_w_mem_3__6_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_442 ( .CLK(clk), .D(w_mem_inst__0w_mem_3__31_0__7_), .Q(w_mem_inst_w_mem_3__7_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_443 ( .CLK(clk), .D(w_mem_inst__0w_mem_3__31_0__8_), .Q(w_mem_inst_w_mem_3__8_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_444 ( .CLK(clk), .D(w_mem_inst__0w_mem_3__31_0__9_), .Q(w_mem_inst_w_mem_3__9_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_445 ( .CLK(clk), .D(w_mem_inst__0w_mem_3__31_0__10_), .Q(w_mem_inst_w_mem_3__10_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_446 ( .CLK(clk), .D(w_mem_inst__0w_mem_3__31_0__11_), .Q(w_mem_inst_w_mem_3__11_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_447 ( .CLK(clk), .D(w_mem_inst__0w_mem_3__31_0__12_), .Q(w_mem_inst_w_mem_3__12_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_448 ( .CLK(clk), .D(w_mem_inst__0w_mem_3__31_0__13_), .Q(w_mem_inst_w_mem_3__13_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_449 ( .CLK(clk), .D(w_mem_inst__0w_mem_3__31_0__14_), .Q(w_mem_inst_w_mem_3__14_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_45 ( .CLK(clk), .D(_0b_reg_31_0__12_), .Q(b_reg_12_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_450 ( .CLK(clk), .D(w_mem_inst__0w_mem_3__31_0__15_), .Q(w_mem_inst_w_mem_3__15_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_451 ( .CLK(clk), .D(w_mem_inst__0w_mem_3__31_0__16_), .Q(w_mem_inst_w_mem_3__16_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_452 ( .CLK(clk), .D(w_mem_inst__0w_mem_3__31_0__17_), .Q(w_mem_inst_w_mem_3__17_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_453 ( .CLK(clk), .D(w_mem_inst__0w_mem_3__31_0__18_), .Q(w_mem_inst_w_mem_3__18_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_454 ( .CLK(clk), .D(w_mem_inst__0w_mem_3__31_0__19_), .Q(w_mem_inst_w_mem_3__19_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_455 ( .CLK(clk), .D(w_mem_inst__0w_mem_3__31_0__20_), .Q(w_mem_inst_w_mem_3__20_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_456 ( .CLK(clk), .D(w_mem_inst__0w_mem_3__31_0__21_), .Q(w_mem_inst_w_mem_3__21_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_457 ( .CLK(clk), .D(w_mem_inst__0w_mem_3__31_0__22_), .Q(w_mem_inst_w_mem_3__22_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_458 ( .CLK(clk), .D(w_mem_inst__0w_mem_3__31_0__23_), .Q(w_mem_inst_w_mem_3__23_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_459 ( .CLK(clk), .D(w_mem_inst__0w_mem_3__31_0__24_), .Q(w_mem_inst_w_mem_3__24_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_46 ( .CLK(clk), .D(_0b_reg_31_0__13_), .Q(b_reg_13_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_460 ( .CLK(clk), .D(w_mem_inst__0w_mem_3__31_0__25_), .Q(w_mem_inst_w_mem_3__25_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_461 ( .CLK(clk), .D(w_mem_inst__0w_mem_3__31_0__26_), .Q(w_mem_inst_w_mem_3__26_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_462 ( .CLK(clk), .D(w_mem_inst__0w_mem_3__31_0__27_), .Q(w_mem_inst_w_mem_3__27_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_463 ( .CLK(clk), .D(w_mem_inst__0w_mem_3__31_0__28_), .Q(w_mem_inst_w_mem_3__28_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_464 ( .CLK(clk), .D(w_mem_inst__0w_mem_3__31_0__29_), .Q(w_mem_inst_w_mem_3__29_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_465 ( .CLK(clk), .D(w_mem_inst__0w_mem_3__31_0__30_), .Q(w_mem_inst_w_mem_3__30_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_466 ( .CLK(clk), .D(w_mem_inst__0w_mem_3__31_0__31_), .Q(w_mem_inst_w_mem_3__31_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_467 ( .CLK(clk), .D(w_mem_inst__0w_mem_4__31_0__0_), .Q(w_mem_inst_w_mem_4__0_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_468 ( .CLK(clk), .D(w_mem_inst__0w_mem_4__31_0__1_), .Q(w_mem_inst_w_mem_4__1_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_469 ( .CLK(clk), .D(w_mem_inst__0w_mem_4__31_0__2_), .Q(w_mem_inst_w_mem_4__2_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_47 ( .CLK(clk), .D(_0b_reg_31_0__14_), .Q(b_reg_14_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_470 ( .CLK(clk), .D(w_mem_inst__0w_mem_4__31_0__3_), .Q(w_mem_inst_w_mem_4__3_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_471 ( .CLK(clk), .D(w_mem_inst__0w_mem_4__31_0__4_), .Q(w_mem_inst_w_mem_4__4_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_472 ( .CLK(clk), .D(w_mem_inst__0w_mem_4__31_0__5_), .Q(w_mem_inst_w_mem_4__5_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_473 ( .CLK(clk), .D(w_mem_inst__0w_mem_4__31_0__6_), .Q(w_mem_inst_w_mem_4__6_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_474 ( .CLK(clk), .D(w_mem_inst__0w_mem_4__31_0__7_), .Q(w_mem_inst_w_mem_4__7_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_475 ( .CLK(clk), .D(w_mem_inst__0w_mem_4__31_0__8_), .Q(w_mem_inst_w_mem_4__8_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_476 ( .CLK(clk), .D(w_mem_inst__0w_mem_4__31_0__9_), .Q(w_mem_inst_w_mem_4__9_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_477 ( .CLK(clk), .D(w_mem_inst__0w_mem_4__31_0__10_), .Q(w_mem_inst_w_mem_4__10_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_478 ( .CLK(clk), .D(w_mem_inst__0w_mem_4__31_0__11_), .Q(w_mem_inst_w_mem_4__11_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_479 ( .CLK(clk), .D(w_mem_inst__0w_mem_4__31_0__12_), .Q(w_mem_inst_w_mem_4__12_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_48 ( .CLK(clk), .D(_0b_reg_31_0__15_), .Q(b_reg_15_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_480 ( .CLK(clk), .D(w_mem_inst__0w_mem_4__31_0__13_), .Q(w_mem_inst_w_mem_4__13_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_481 ( .CLK(clk), .D(w_mem_inst__0w_mem_4__31_0__14_), .Q(w_mem_inst_w_mem_4__14_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_482 ( .CLK(clk), .D(w_mem_inst__0w_mem_4__31_0__15_), .Q(w_mem_inst_w_mem_4__15_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_483 ( .CLK(clk), .D(w_mem_inst__0w_mem_4__31_0__16_), .Q(w_mem_inst_w_mem_4__16_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_484 ( .CLK(clk), .D(w_mem_inst__0w_mem_4__31_0__17_), .Q(w_mem_inst_w_mem_4__17_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_485 ( .CLK(clk), .D(w_mem_inst__0w_mem_4__31_0__18_), .Q(w_mem_inst_w_mem_4__18_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_486 ( .CLK(clk), .D(w_mem_inst__0w_mem_4__31_0__19_), .Q(w_mem_inst_w_mem_4__19_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_487 ( .CLK(clk), .D(w_mem_inst__0w_mem_4__31_0__20_), .Q(w_mem_inst_w_mem_4__20_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_488 ( .CLK(clk), .D(w_mem_inst__0w_mem_4__31_0__21_), .Q(w_mem_inst_w_mem_4__21_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_489 ( .CLK(clk), .D(w_mem_inst__0w_mem_4__31_0__22_), .Q(w_mem_inst_w_mem_4__22_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_49 ( .CLK(clk), .D(_0b_reg_31_0__16_), .Q(b_reg_16_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_490 ( .CLK(clk), .D(w_mem_inst__0w_mem_4__31_0__23_), .Q(w_mem_inst_w_mem_4__23_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_491 ( .CLK(clk), .D(w_mem_inst__0w_mem_4__31_0__24_), .Q(w_mem_inst_w_mem_4__24_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_492 ( .CLK(clk), .D(w_mem_inst__0w_mem_4__31_0__25_), .Q(w_mem_inst_w_mem_4__25_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_493 ( .CLK(clk), .D(w_mem_inst__0w_mem_4__31_0__26_), .Q(w_mem_inst_w_mem_4__26_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_494 ( .CLK(clk), .D(w_mem_inst__0w_mem_4__31_0__27_), .Q(w_mem_inst_w_mem_4__27_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_495 ( .CLK(clk), .D(w_mem_inst__0w_mem_4__31_0__28_), .Q(w_mem_inst_w_mem_4__28_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_496 ( .CLK(clk), .D(w_mem_inst__0w_mem_4__31_0__29_), .Q(w_mem_inst_w_mem_4__29_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_497 ( .CLK(clk), .D(w_mem_inst__0w_mem_4__31_0__30_), .Q(w_mem_inst_w_mem_4__30_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_498 ( .CLK(clk), .D(w_mem_inst__0w_mem_4__31_0__31_), .Q(w_mem_inst_w_mem_4__31_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_499 ( .CLK(clk), .D(w_mem_inst__0w_mem_5__31_0__0_), .Q(w_mem_inst_w_mem_5__0_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_5 ( .CLK(clk), .D(_0a_reg_31_0__4_), .Q(a_reg_4_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_50 ( .CLK(clk), .D(_0b_reg_31_0__17_), .Q(b_reg_17_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_500 ( .CLK(clk), .D(w_mem_inst__0w_mem_5__31_0__1_), .Q(w_mem_inst_w_mem_5__1_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_501 ( .CLK(clk), .D(w_mem_inst__0w_mem_5__31_0__2_), .Q(w_mem_inst_w_mem_5__2_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_502 ( .CLK(clk), .D(w_mem_inst__0w_mem_5__31_0__3_), .Q(w_mem_inst_w_mem_5__3_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_503 ( .CLK(clk), .D(w_mem_inst__0w_mem_5__31_0__4_), .Q(w_mem_inst_w_mem_5__4_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_504 ( .CLK(clk), .D(w_mem_inst__0w_mem_5__31_0__5_), .Q(w_mem_inst_w_mem_5__5_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_505 ( .CLK(clk), .D(w_mem_inst__0w_mem_5__31_0__6_), .Q(w_mem_inst_w_mem_5__6_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_506 ( .CLK(clk), .D(w_mem_inst__0w_mem_5__31_0__7_), .Q(w_mem_inst_w_mem_5__7_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_507 ( .CLK(clk), .D(w_mem_inst__0w_mem_5__31_0__8_), .Q(w_mem_inst_w_mem_5__8_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_508 ( .CLK(clk), .D(w_mem_inst__0w_mem_5__31_0__9_), .Q(w_mem_inst_w_mem_5__9_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_509 ( .CLK(clk), .D(w_mem_inst__0w_mem_5__31_0__10_), .Q(w_mem_inst_w_mem_5__10_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_51 ( .CLK(clk), .D(_0b_reg_31_0__18_), .Q(b_reg_18_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_510 ( .CLK(clk), .D(w_mem_inst__0w_mem_5__31_0__11_), .Q(w_mem_inst_w_mem_5__11_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_511 ( .CLK(clk), .D(w_mem_inst__0w_mem_5__31_0__12_), .Q(w_mem_inst_w_mem_5__12_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_512 ( .CLK(clk), .D(w_mem_inst__0w_mem_5__31_0__13_), .Q(w_mem_inst_w_mem_5__13_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_513 ( .CLK(clk), .D(w_mem_inst__0w_mem_5__31_0__14_), .Q(w_mem_inst_w_mem_5__14_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_514 ( .CLK(clk), .D(w_mem_inst__0w_mem_5__31_0__15_), .Q(w_mem_inst_w_mem_5__15_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_515 ( .CLK(clk), .D(w_mem_inst__0w_mem_5__31_0__16_), .Q(w_mem_inst_w_mem_5__16_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_516 ( .CLK(clk), .D(w_mem_inst__0w_mem_5__31_0__17_), .Q(w_mem_inst_w_mem_5__17_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_517 ( .CLK(clk), .D(w_mem_inst__0w_mem_5__31_0__18_), .Q(w_mem_inst_w_mem_5__18_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_518 ( .CLK(clk), .D(w_mem_inst__0w_mem_5__31_0__19_), .Q(w_mem_inst_w_mem_5__19_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_519 ( .CLK(clk), .D(w_mem_inst__0w_mem_5__31_0__20_), .Q(w_mem_inst_w_mem_5__20_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_52 ( .CLK(clk), .D(_0b_reg_31_0__19_), .Q(b_reg_19_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_520 ( .CLK(clk), .D(w_mem_inst__0w_mem_5__31_0__21_), .Q(w_mem_inst_w_mem_5__21_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_521 ( .CLK(clk), .D(w_mem_inst__0w_mem_5__31_0__22_), .Q(w_mem_inst_w_mem_5__22_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_522 ( .CLK(clk), .D(w_mem_inst__0w_mem_5__31_0__23_), .Q(w_mem_inst_w_mem_5__23_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_523 ( .CLK(clk), .D(w_mem_inst__0w_mem_5__31_0__24_), .Q(w_mem_inst_w_mem_5__24_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_524 ( .CLK(clk), .D(w_mem_inst__0w_mem_5__31_0__25_), .Q(w_mem_inst_w_mem_5__25_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_525 ( .CLK(clk), .D(w_mem_inst__0w_mem_5__31_0__26_), .Q(w_mem_inst_w_mem_5__26_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_526 ( .CLK(clk), .D(w_mem_inst__0w_mem_5__31_0__27_), .Q(w_mem_inst_w_mem_5__27_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_527 ( .CLK(clk), .D(w_mem_inst__0w_mem_5__31_0__28_), .Q(w_mem_inst_w_mem_5__28_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_528 ( .CLK(clk), .D(w_mem_inst__0w_mem_5__31_0__29_), .Q(w_mem_inst_w_mem_5__29_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_529 ( .CLK(clk), .D(w_mem_inst__0w_mem_5__31_0__30_), .Q(w_mem_inst_w_mem_5__30_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_53 ( .CLK(clk), .D(_0b_reg_31_0__20_), .Q(b_reg_20_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_530 ( .CLK(clk), .D(w_mem_inst__0w_mem_5__31_0__31_), .Q(w_mem_inst_w_mem_5__31_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_531 ( .CLK(clk), .D(w_mem_inst__0w_mem_6__31_0__0_), .Q(w_mem_inst_w_mem_6__0_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_532 ( .CLK(clk), .D(w_mem_inst__0w_mem_6__31_0__1_), .Q(w_mem_inst_w_mem_6__1_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_533 ( .CLK(clk), .D(w_mem_inst__0w_mem_6__31_0__2_), .Q(w_mem_inst_w_mem_6__2_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_534 ( .CLK(clk), .D(w_mem_inst__0w_mem_6__31_0__3_), .Q(w_mem_inst_w_mem_6__3_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_535 ( .CLK(clk), .D(w_mem_inst__0w_mem_6__31_0__4_), .Q(w_mem_inst_w_mem_6__4_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_536 ( .CLK(clk), .D(w_mem_inst__0w_mem_6__31_0__5_), .Q(w_mem_inst_w_mem_6__5_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_537 ( .CLK(clk), .D(w_mem_inst__0w_mem_6__31_0__6_), .Q(w_mem_inst_w_mem_6__6_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_538 ( .CLK(clk), .D(w_mem_inst__0w_mem_6__31_0__7_), .Q(w_mem_inst_w_mem_6__7_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_539 ( .CLK(clk), .D(w_mem_inst__0w_mem_6__31_0__8_), .Q(w_mem_inst_w_mem_6__8_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_54 ( .CLK(clk), .D(_0b_reg_31_0__21_), .Q(b_reg_21_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_540 ( .CLK(clk), .D(w_mem_inst__0w_mem_6__31_0__9_), .Q(w_mem_inst_w_mem_6__9_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_541 ( .CLK(clk), .D(w_mem_inst__0w_mem_6__31_0__10_), .Q(w_mem_inst_w_mem_6__10_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_542 ( .CLK(clk), .D(w_mem_inst__0w_mem_6__31_0__11_), .Q(w_mem_inst_w_mem_6__11_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_543 ( .CLK(clk), .D(w_mem_inst__0w_mem_6__31_0__12_), .Q(w_mem_inst_w_mem_6__12_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_544 ( .CLK(clk), .D(w_mem_inst__0w_mem_6__31_0__13_), .Q(w_mem_inst_w_mem_6__13_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_545 ( .CLK(clk), .D(w_mem_inst__0w_mem_6__31_0__14_), .Q(w_mem_inst_w_mem_6__14_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_546 ( .CLK(clk), .D(w_mem_inst__0w_mem_6__31_0__15_), .Q(w_mem_inst_w_mem_6__15_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_547 ( .CLK(clk), .D(w_mem_inst__0w_mem_6__31_0__16_), .Q(w_mem_inst_w_mem_6__16_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_548 ( .CLK(clk), .D(w_mem_inst__0w_mem_6__31_0__17_), .Q(w_mem_inst_w_mem_6__17_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_549 ( .CLK(clk), .D(w_mem_inst__0w_mem_6__31_0__18_), .Q(w_mem_inst_w_mem_6__18_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_55 ( .CLK(clk), .D(_0b_reg_31_0__22_), .Q(b_reg_22_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_550 ( .CLK(clk), .D(w_mem_inst__0w_mem_6__31_0__19_), .Q(w_mem_inst_w_mem_6__19_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_551 ( .CLK(clk), .D(w_mem_inst__0w_mem_6__31_0__20_), .Q(w_mem_inst_w_mem_6__20_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_552 ( .CLK(clk), .D(w_mem_inst__0w_mem_6__31_0__21_), .Q(w_mem_inst_w_mem_6__21_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_553 ( .CLK(clk), .D(w_mem_inst__0w_mem_6__31_0__22_), .Q(w_mem_inst_w_mem_6__22_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_554 ( .CLK(clk), .D(w_mem_inst__0w_mem_6__31_0__23_), .Q(w_mem_inst_w_mem_6__23_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_555 ( .CLK(clk), .D(w_mem_inst__0w_mem_6__31_0__24_), .Q(w_mem_inst_w_mem_6__24_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_556 ( .CLK(clk), .D(w_mem_inst__0w_mem_6__31_0__25_), .Q(w_mem_inst_w_mem_6__25_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_557 ( .CLK(clk), .D(w_mem_inst__0w_mem_6__31_0__26_), .Q(w_mem_inst_w_mem_6__26_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_558 ( .CLK(clk), .D(w_mem_inst__0w_mem_6__31_0__27_), .Q(w_mem_inst_w_mem_6__27_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_559 ( .CLK(clk), .D(w_mem_inst__0w_mem_6__31_0__28_), .Q(w_mem_inst_w_mem_6__28_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_56 ( .CLK(clk), .D(_0b_reg_31_0__23_), .Q(b_reg_23_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_560 ( .CLK(clk), .D(w_mem_inst__0w_mem_6__31_0__29_), .Q(w_mem_inst_w_mem_6__29_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_561 ( .CLK(clk), .D(w_mem_inst__0w_mem_6__31_0__30_), .Q(w_mem_inst_w_mem_6__30_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_562 ( .CLK(clk), .D(w_mem_inst__0w_mem_6__31_0__31_), .Q(w_mem_inst_w_mem_6__31_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_563 ( .CLK(clk), .D(w_mem_inst__0w_mem_7__31_0__0_), .Q(w_mem_inst_w_mem_7__0_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_564 ( .CLK(clk), .D(w_mem_inst__0w_mem_7__31_0__1_), .Q(w_mem_inst_w_mem_7__1_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_565 ( .CLK(clk), .D(w_mem_inst__0w_mem_7__31_0__2_), .Q(w_mem_inst_w_mem_7__2_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_566 ( .CLK(clk), .D(w_mem_inst__0w_mem_7__31_0__3_), .Q(w_mem_inst_w_mem_7__3_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_567 ( .CLK(clk), .D(w_mem_inst__0w_mem_7__31_0__4_), .Q(w_mem_inst_w_mem_7__4_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_568 ( .CLK(clk), .D(w_mem_inst__0w_mem_7__31_0__5_), .Q(w_mem_inst_w_mem_7__5_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_569 ( .CLK(clk), .D(w_mem_inst__0w_mem_7__31_0__6_), .Q(w_mem_inst_w_mem_7__6_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_57 ( .CLK(clk), .D(_0b_reg_31_0__24_), .Q(b_reg_24_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_570 ( .CLK(clk), .D(w_mem_inst__0w_mem_7__31_0__7_), .Q(w_mem_inst_w_mem_7__7_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_571 ( .CLK(clk), .D(w_mem_inst__0w_mem_7__31_0__8_), .Q(w_mem_inst_w_mem_7__8_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_572 ( .CLK(clk), .D(w_mem_inst__0w_mem_7__31_0__9_), .Q(w_mem_inst_w_mem_7__9_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_573 ( .CLK(clk), .D(w_mem_inst__0w_mem_7__31_0__10_), .Q(w_mem_inst_w_mem_7__10_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_574 ( .CLK(clk), .D(w_mem_inst__0w_mem_7__31_0__11_), .Q(w_mem_inst_w_mem_7__11_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_575 ( .CLK(clk), .D(w_mem_inst__0w_mem_7__31_0__12_), .Q(w_mem_inst_w_mem_7__12_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_576 ( .CLK(clk), .D(w_mem_inst__0w_mem_7__31_0__13_), .Q(w_mem_inst_w_mem_7__13_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_577 ( .CLK(clk), .D(w_mem_inst__0w_mem_7__31_0__14_), .Q(w_mem_inst_w_mem_7__14_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_578 ( .CLK(clk), .D(w_mem_inst__0w_mem_7__31_0__15_), .Q(w_mem_inst_w_mem_7__15_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_579 ( .CLK(clk), .D(w_mem_inst__0w_mem_7__31_0__16_), .Q(w_mem_inst_w_mem_7__16_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_58 ( .CLK(clk), .D(_0b_reg_31_0__25_), .Q(b_reg_25_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_580 ( .CLK(clk), .D(w_mem_inst__0w_mem_7__31_0__17_), .Q(w_mem_inst_w_mem_7__17_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_581 ( .CLK(clk), .D(w_mem_inst__0w_mem_7__31_0__18_), .Q(w_mem_inst_w_mem_7__18_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_582 ( .CLK(clk), .D(w_mem_inst__0w_mem_7__31_0__19_), .Q(w_mem_inst_w_mem_7__19_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_583 ( .CLK(clk), .D(w_mem_inst__0w_mem_7__31_0__20_), .Q(w_mem_inst_w_mem_7__20_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_584 ( .CLK(clk), .D(w_mem_inst__0w_mem_7__31_0__21_), .Q(w_mem_inst_w_mem_7__21_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_585 ( .CLK(clk), .D(w_mem_inst__0w_mem_7__31_0__22_), .Q(w_mem_inst_w_mem_7__22_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_586 ( .CLK(clk), .D(w_mem_inst__0w_mem_7__31_0__23_), .Q(w_mem_inst_w_mem_7__23_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_587 ( .CLK(clk), .D(w_mem_inst__0w_mem_7__31_0__24_), .Q(w_mem_inst_w_mem_7__24_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_588 ( .CLK(clk), .D(w_mem_inst__0w_mem_7__31_0__25_), .Q(w_mem_inst_w_mem_7__25_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_589 ( .CLK(clk), .D(w_mem_inst__0w_mem_7__31_0__26_), .Q(w_mem_inst_w_mem_7__26_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_59 ( .CLK(clk), .D(_0b_reg_31_0__26_), .Q(b_reg_26_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_590 ( .CLK(clk), .D(w_mem_inst__0w_mem_7__31_0__27_), .Q(w_mem_inst_w_mem_7__27_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_591 ( .CLK(clk), .D(w_mem_inst__0w_mem_7__31_0__28_), .Q(w_mem_inst_w_mem_7__28_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_592 ( .CLK(clk), .D(w_mem_inst__0w_mem_7__31_0__29_), .Q(w_mem_inst_w_mem_7__29_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_593 ( .CLK(clk), .D(w_mem_inst__0w_mem_7__31_0__30_), .Q(w_mem_inst_w_mem_7__30_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_594 ( .CLK(clk), .D(w_mem_inst__0w_mem_7__31_0__31_), .Q(w_mem_inst_w_mem_7__31_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_595 ( .CLK(clk), .D(w_mem_inst__0w_mem_8__31_0__0_), .Q(w_mem_inst_w_mem_8__0_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_596 ( .CLK(clk), .D(w_mem_inst__0w_mem_8__31_0__1_), .Q(w_mem_inst_w_mem_8__1_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_597 ( .CLK(clk), .D(w_mem_inst__0w_mem_8__31_0__2_), .Q(w_mem_inst_w_mem_8__2_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_598 ( .CLK(clk), .D(w_mem_inst__0w_mem_8__31_0__3_), .Q(w_mem_inst_w_mem_8__3_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_599 ( .CLK(clk), .D(w_mem_inst__0w_mem_8__31_0__4_), .Q(w_mem_inst_w_mem_8__4_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_6 ( .CLK(clk), .D(_0a_reg_31_0__5_), .Q(a_reg_5_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_60 ( .CLK(clk), .D(_0b_reg_31_0__27_), .Q(b_reg_27_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_600 ( .CLK(clk), .D(w_mem_inst__0w_mem_8__31_0__5_), .Q(w_mem_inst_w_mem_8__5_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_601 ( .CLK(clk), .D(w_mem_inst__0w_mem_8__31_0__6_), .Q(w_mem_inst_w_mem_8__6_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_602 ( .CLK(clk), .D(w_mem_inst__0w_mem_8__31_0__7_), .Q(w_mem_inst_w_mem_8__7_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_603 ( .CLK(clk), .D(w_mem_inst__0w_mem_8__31_0__8_), .Q(w_mem_inst_w_mem_8__8_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_604 ( .CLK(clk), .D(w_mem_inst__0w_mem_8__31_0__9_), .Q(w_mem_inst_w_mem_8__9_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_605 ( .CLK(clk), .D(w_mem_inst__0w_mem_8__31_0__10_), .Q(w_mem_inst_w_mem_8__10_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_606 ( .CLK(clk), .D(w_mem_inst__0w_mem_8__31_0__11_), .Q(w_mem_inst_w_mem_8__11_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_607 ( .CLK(clk), .D(w_mem_inst__0w_mem_8__31_0__12_), .Q(w_mem_inst_w_mem_8__12_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_608 ( .CLK(clk), .D(w_mem_inst__0w_mem_8__31_0__13_), .Q(w_mem_inst_w_mem_8__13_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_609 ( .CLK(clk), .D(w_mem_inst__0w_mem_8__31_0__14_), .Q(w_mem_inst_w_mem_8__14_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_61 ( .CLK(clk), .D(_0b_reg_31_0__28_), .Q(b_reg_28_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_610 ( .CLK(clk), .D(w_mem_inst__0w_mem_8__31_0__15_), .Q(w_mem_inst_w_mem_8__15_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_611 ( .CLK(clk), .D(w_mem_inst__0w_mem_8__31_0__16_), .Q(w_mem_inst_w_mem_8__16_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_612 ( .CLK(clk), .D(w_mem_inst__0w_mem_8__31_0__17_), .Q(w_mem_inst_w_mem_8__17_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_613 ( .CLK(clk), .D(w_mem_inst__0w_mem_8__31_0__18_), .Q(w_mem_inst_w_mem_8__18_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_614 ( .CLK(clk), .D(w_mem_inst__0w_mem_8__31_0__19_), .Q(w_mem_inst_w_mem_8__19_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_615 ( .CLK(clk), .D(w_mem_inst__0w_mem_8__31_0__20_), .Q(w_mem_inst_w_mem_8__20_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_616 ( .CLK(clk), .D(w_mem_inst__0w_mem_8__31_0__21_), .Q(w_mem_inst_w_mem_8__21_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_617 ( .CLK(clk), .D(w_mem_inst__0w_mem_8__31_0__22_), .Q(w_mem_inst_w_mem_8__22_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_618 ( .CLK(clk), .D(w_mem_inst__0w_mem_8__31_0__23_), .Q(w_mem_inst_w_mem_8__23_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_619 ( .CLK(clk), .D(w_mem_inst__0w_mem_8__31_0__24_), .Q(w_mem_inst_w_mem_8__24_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_62 ( .CLK(clk), .D(_0b_reg_31_0__29_), .Q(b_reg_29_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_620 ( .CLK(clk), .D(w_mem_inst__0w_mem_8__31_0__25_), .Q(w_mem_inst_w_mem_8__25_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_621 ( .CLK(clk), .D(w_mem_inst__0w_mem_8__31_0__26_), .Q(w_mem_inst_w_mem_8__26_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_622 ( .CLK(clk), .D(w_mem_inst__0w_mem_8__31_0__27_), .Q(w_mem_inst_w_mem_8__27_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_623 ( .CLK(clk), .D(w_mem_inst__0w_mem_8__31_0__28_), .Q(w_mem_inst_w_mem_8__28_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_624 ( .CLK(clk), .D(w_mem_inst__0w_mem_8__31_0__29_), .Q(w_mem_inst_w_mem_8__29_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_625 ( .CLK(clk), .D(w_mem_inst__0w_mem_8__31_0__30_), .Q(w_mem_inst_w_mem_8__30_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_626 ( .CLK(clk), .D(w_mem_inst__0w_mem_8__31_0__31_), .Q(w_mem_inst_w_mem_8__31_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_627 ( .CLK(clk), .D(w_mem_inst__0w_mem_9__31_0__0_), .Q(w_mem_inst_w_mem_9__0_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_628 ( .CLK(clk), .D(w_mem_inst__0w_mem_9__31_0__1_), .Q(w_mem_inst_w_mem_9__1_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_629 ( .CLK(clk), .D(w_mem_inst__0w_mem_9__31_0__2_), .Q(w_mem_inst_w_mem_9__2_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_63 ( .CLK(clk), .D(_0b_reg_31_0__30_), .Q(b_reg_30_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_630 ( .CLK(clk), .D(w_mem_inst__0w_mem_9__31_0__3_), .Q(w_mem_inst_w_mem_9__3_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_631 ( .CLK(clk), .D(w_mem_inst__0w_mem_9__31_0__4_), .Q(w_mem_inst_w_mem_9__4_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_632 ( .CLK(clk), .D(w_mem_inst__0w_mem_9__31_0__5_), .Q(w_mem_inst_w_mem_9__5_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_633 ( .CLK(clk), .D(w_mem_inst__0w_mem_9__31_0__6_), .Q(w_mem_inst_w_mem_9__6_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_634 ( .CLK(clk), .D(w_mem_inst__0w_mem_9__31_0__7_), .Q(w_mem_inst_w_mem_9__7_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_635 ( .CLK(clk), .D(w_mem_inst__0w_mem_9__31_0__8_), .Q(w_mem_inst_w_mem_9__8_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_636 ( .CLK(clk), .D(w_mem_inst__0w_mem_9__31_0__9_), .Q(w_mem_inst_w_mem_9__9_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_637 ( .CLK(clk), .D(w_mem_inst__0w_mem_9__31_0__10_), .Q(w_mem_inst_w_mem_9__10_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_638 ( .CLK(clk), .D(w_mem_inst__0w_mem_9__31_0__11_), .Q(w_mem_inst_w_mem_9__11_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_639 ( .CLK(clk), .D(w_mem_inst__0w_mem_9__31_0__12_), .Q(w_mem_inst_w_mem_9__12_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_64 ( .CLK(clk), .D(_0b_reg_31_0__31_), .Q(b_reg_31_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_640 ( .CLK(clk), .D(w_mem_inst__0w_mem_9__31_0__13_), .Q(w_mem_inst_w_mem_9__13_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_641 ( .CLK(clk), .D(w_mem_inst__0w_mem_9__31_0__14_), .Q(w_mem_inst_w_mem_9__14_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_642 ( .CLK(clk), .D(w_mem_inst__0w_mem_9__31_0__15_), .Q(w_mem_inst_w_mem_9__15_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_643 ( .CLK(clk), .D(w_mem_inst__0w_mem_9__31_0__16_), .Q(w_mem_inst_w_mem_9__16_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_644 ( .CLK(clk), .D(w_mem_inst__0w_mem_9__31_0__17_), .Q(w_mem_inst_w_mem_9__17_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_645 ( .CLK(clk), .D(w_mem_inst__0w_mem_9__31_0__18_), .Q(w_mem_inst_w_mem_9__18_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_646 ( .CLK(clk), .D(w_mem_inst__0w_mem_9__31_0__19_), .Q(w_mem_inst_w_mem_9__19_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_647 ( .CLK(clk), .D(w_mem_inst__0w_mem_9__31_0__20_), .Q(w_mem_inst_w_mem_9__20_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_648 ( .CLK(clk), .D(w_mem_inst__0w_mem_9__31_0__21_), .Q(w_mem_inst_w_mem_9__21_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_649 ( .CLK(clk), .D(w_mem_inst__0w_mem_9__31_0__22_), .Q(w_mem_inst_w_mem_9__22_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_65 ( .CLK(clk), .D(_0c_reg_31_0__0_), .Q(c_reg_0_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_650 ( .CLK(clk), .D(w_mem_inst__0w_mem_9__31_0__23_), .Q(w_mem_inst_w_mem_9__23_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_651 ( .CLK(clk), .D(w_mem_inst__0w_mem_9__31_0__24_), .Q(w_mem_inst_w_mem_9__24_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_652 ( .CLK(clk), .D(w_mem_inst__0w_mem_9__31_0__25_), .Q(w_mem_inst_w_mem_9__25_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_653 ( .CLK(clk), .D(w_mem_inst__0w_mem_9__31_0__26_), .Q(w_mem_inst_w_mem_9__26_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_654 ( .CLK(clk), .D(w_mem_inst__0w_mem_9__31_0__27_), .Q(w_mem_inst_w_mem_9__27_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_655 ( .CLK(clk), .D(w_mem_inst__0w_mem_9__31_0__28_), .Q(w_mem_inst_w_mem_9__28_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_656 ( .CLK(clk), .D(w_mem_inst__0w_mem_9__31_0__29_), .Q(w_mem_inst_w_mem_9__29_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_657 ( .CLK(clk), .D(w_mem_inst__0w_mem_9__31_0__30_), .Q(w_mem_inst_w_mem_9__30_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_658 ( .CLK(clk), .D(w_mem_inst__0w_mem_9__31_0__31_), .Q(w_mem_inst_w_mem_9__31_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_659 ( .CLK(clk), .D(w_mem_inst__0w_mem_10__31_0__0_), .Q(w_mem_inst_w_mem_10__0_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_66 ( .CLK(clk), .D(_0c_reg_31_0__1_), .Q(c_reg_1_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_660 ( .CLK(clk), .D(w_mem_inst__0w_mem_10__31_0__1_), .Q(w_mem_inst_w_mem_10__1_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_661 ( .CLK(clk), .D(w_mem_inst__0w_mem_10__31_0__2_), .Q(w_mem_inst_w_mem_10__2_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_662 ( .CLK(clk), .D(w_mem_inst__0w_mem_10__31_0__3_), .Q(w_mem_inst_w_mem_10__3_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_663 ( .CLK(clk), .D(w_mem_inst__0w_mem_10__31_0__4_), .Q(w_mem_inst_w_mem_10__4_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_664 ( .CLK(clk), .D(w_mem_inst__0w_mem_10__31_0__5_), .Q(w_mem_inst_w_mem_10__5_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_665 ( .CLK(clk), .D(w_mem_inst__0w_mem_10__31_0__6_), .Q(w_mem_inst_w_mem_10__6_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_666 ( .CLK(clk), .D(w_mem_inst__0w_mem_10__31_0__7_), .Q(w_mem_inst_w_mem_10__7_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_667 ( .CLK(clk), .D(w_mem_inst__0w_mem_10__31_0__8_), .Q(w_mem_inst_w_mem_10__8_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_668 ( .CLK(clk), .D(w_mem_inst__0w_mem_10__31_0__9_), .Q(w_mem_inst_w_mem_10__9_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_669 ( .CLK(clk), .D(w_mem_inst__0w_mem_10__31_0__10_), .Q(w_mem_inst_w_mem_10__10_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_67 ( .CLK(clk), .D(_0c_reg_31_0__2_), .Q(c_reg_2_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_670 ( .CLK(clk), .D(w_mem_inst__0w_mem_10__31_0__11_), .Q(w_mem_inst_w_mem_10__11_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_671 ( .CLK(clk), .D(w_mem_inst__0w_mem_10__31_0__12_), .Q(w_mem_inst_w_mem_10__12_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_672 ( .CLK(clk), .D(w_mem_inst__0w_mem_10__31_0__13_), .Q(w_mem_inst_w_mem_10__13_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_673 ( .CLK(clk), .D(w_mem_inst__0w_mem_10__31_0__14_), .Q(w_mem_inst_w_mem_10__14_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_674 ( .CLK(clk), .D(w_mem_inst__0w_mem_10__31_0__15_), .Q(w_mem_inst_w_mem_10__15_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_675 ( .CLK(clk), .D(w_mem_inst__0w_mem_10__31_0__16_), .Q(w_mem_inst_w_mem_10__16_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_676 ( .CLK(clk), .D(w_mem_inst__0w_mem_10__31_0__17_), .Q(w_mem_inst_w_mem_10__17_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_677 ( .CLK(clk), .D(w_mem_inst__0w_mem_10__31_0__18_), .Q(w_mem_inst_w_mem_10__18_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_678 ( .CLK(clk), .D(w_mem_inst__0w_mem_10__31_0__19_), .Q(w_mem_inst_w_mem_10__19_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_679 ( .CLK(clk), .D(w_mem_inst__0w_mem_10__31_0__20_), .Q(w_mem_inst_w_mem_10__20_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_68 ( .CLK(clk), .D(_0c_reg_31_0__3_), .Q(c_reg_3_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_680 ( .CLK(clk), .D(w_mem_inst__0w_mem_10__31_0__21_), .Q(w_mem_inst_w_mem_10__21_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_681 ( .CLK(clk), .D(w_mem_inst__0w_mem_10__31_0__22_), .Q(w_mem_inst_w_mem_10__22_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_682 ( .CLK(clk), .D(w_mem_inst__0w_mem_10__31_0__23_), .Q(w_mem_inst_w_mem_10__23_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_683 ( .CLK(clk), .D(w_mem_inst__0w_mem_10__31_0__24_), .Q(w_mem_inst_w_mem_10__24_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_684 ( .CLK(clk), .D(w_mem_inst__0w_mem_10__31_0__25_), .Q(w_mem_inst_w_mem_10__25_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_685 ( .CLK(clk), .D(w_mem_inst__0w_mem_10__31_0__26_), .Q(w_mem_inst_w_mem_10__26_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_686 ( .CLK(clk), .D(w_mem_inst__0w_mem_10__31_0__27_), .Q(w_mem_inst_w_mem_10__27_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_687 ( .CLK(clk), .D(w_mem_inst__0w_mem_10__31_0__28_), .Q(w_mem_inst_w_mem_10__28_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_688 ( .CLK(clk), .D(w_mem_inst__0w_mem_10__31_0__29_), .Q(w_mem_inst_w_mem_10__29_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_689 ( .CLK(clk), .D(w_mem_inst__0w_mem_10__31_0__30_), .Q(w_mem_inst_w_mem_10__30_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_69 ( .CLK(clk), .D(_0c_reg_31_0__4_), .Q(c_reg_4_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_690 ( .CLK(clk), .D(w_mem_inst__0w_mem_10__31_0__31_), .Q(w_mem_inst_w_mem_10__31_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_691 ( .CLK(clk), .D(w_mem_inst__0w_mem_11__31_0__0_), .Q(w_mem_inst_w_mem_11__0_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_692 ( .CLK(clk), .D(w_mem_inst__0w_mem_11__31_0__1_), .Q(w_mem_inst_w_mem_11__1_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_693 ( .CLK(clk), .D(w_mem_inst__0w_mem_11__31_0__2_), .Q(w_mem_inst_w_mem_11__2_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_694 ( .CLK(clk), .D(w_mem_inst__0w_mem_11__31_0__3_), .Q(w_mem_inst_w_mem_11__3_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_695 ( .CLK(clk), .D(w_mem_inst__0w_mem_11__31_0__4_), .Q(w_mem_inst_w_mem_11__4_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_696 ( .CLK(clk), .D(w_mem_inst__0w_mem_11__31_0__5_), .Q(w_mem_inst_w_mem_11__5_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_697 ( .CLK(clk), .D(w_mem_inst__0w_mem_11__31_0__6_), .Q(w_mem_inst_w_mem_11__6_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_698 ( .CLK(clk), .D(w_mem_inst__0w_mem_11__31_0__7_), .Q(w_mem_inst_w_mem_11__7_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_699 ( .CLK(clk), .D(w_mem_inst__0w_mem_11__31_0__8_), .Q(w_mem_inst_w_mem_11__8_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_7 ( .CLK(clk), .D(_0a_reg_31_0__6_), .Q(a_reg_6_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_70 ( .CLK(clk), .D(_0c_reg_31_0__5_), .Q(c_reg_5_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_700 ( .CLK(clk), .D(w_mem_inst__0w_mem_11__31_0__9_), .Q(w_mem_inst_w_mem_11__9_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_701 ( .CLK(clk), .D(w_mem_inst__0w_mem_11__31_0__10_), .Q(w_mem_inst_w_mem_11__10_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_702 ( .CLK(clk), .D(w_mem_inst__0w_mem_11__31_0__11_), .Q(w_mem_inst_w_mem_11__11_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_703 ( .CLK(clk), .D(w_mem_inst__0w_mem_11__31_0__12_), .Q(w_mem_inst_w_mem_11__12_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_704 ( .CLK(clk), .D(w_mem_inst__0w_mem_11__31_0__13_), .Q(w_mem_inst_w_mem_11__13_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_705 ( .CLK(clk), .D(w_mem_inst__0w_mem_11__31_0__14_), .Q(w_mem_inst_w_mem_11__14_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_706 ( .CLK(clk), .D(w_mem_inst__0w_mem_11__31_0__15_), .Q(w_mem_inst_w_mem_11__15_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_707 ( .CLK(clk), .D(w_mem_inst__0w_mem_11__31_0__16_), .Q(w_mem_inst_w_mem_11__16_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_708 ( .CLK(clk), .D(w_mem_inst__0w_mem_11__31_0__17_), .Q(w_mem_inst_w_mem_11__17_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_709 ( .CLK(clk), .D(w_mem_inst__0w_mem_11__31_0__18_), .Q(w_mem_inst_w_mem_11__18_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_71 ( .CLK(clk), .D(_0c_reg_31_0__6_), .Q(c_reg_6_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_710 ( .CLK(clk), .D(w_mem_inst__0w_mem_11__31_0__19_), .Q(w_mem_inst_w_mem_11__19_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_711 ( .CLK(clk), .D(w_mem_inst__0w_mem_11__31_0__20_), .Q(w_mem_inst_w_mem_11__20_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_712 ( .CLK(clk), .D(w_mem_inst__0w_mem_11__31_0__21_), .Q(w_mem_inst_w_mem_11__21_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_713 ( .CLK(clk), .D(w_mem_inst__0w_mem_11__31_0__22_), .Q(w_mem_inst_w_mem_11__22_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_714 ( .CLK(clk), .D(w_mem_inst__0w_mem_11__31_0__23_), .Q(w_mem_inst_w_mem_11__23_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_715 ( .CLK(clk), .D(w_mem_inst__0w_mem_11__31_0__24_), .Q(w_mem_inst_w_mem_11__24_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_716 ( .CLK(clk), .D(w_mem_inst__0w_mem_11__31_0__25_), .Q(w_mem_inst_w_mem_11__25_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_717 ( .CLK(clk), .D(w_mem_inst__0w_mem_11__31_0__26_), .Q(w_mem_inst_w_mem_11__26_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_718 ( .CLK(clk), .D(w_mem_inst__0w_mem_11__31_0__27_), .Q(w_mem_inst_w_mem_11__27_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_719 ( .CLK(clk), .D(w_mem_inst__0w_mem_11__31_0__28_), .Q(w_mem_inst_w_mem_11__28_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_72 ( .CLK(clk), .D(_0c_reg_31_0__7_), .Q(c_reg_7_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_720 ( .CLK(clk), .D(w_mem_inst__0w_mem_11__31_0__29_), .Q(w_mem_inst_w_mem_11__29_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_721 ( .CLK(clk), .D(w_mem_inst__0w_mem_11__31_0__30_), .Q(w_mem_inst_w_mem_11__30_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_722 ( .CLK(clk), .D(w_mem_inst__0w_mem_11__31_0__31_), .Q(w_mem_inst_w_mem_11__31_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_723 ( .CLK(clk), .D(w_mem_inst__0w_mem_12__31_0__0_), .Q(w_mem_inst_w_mem_12__0_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_724 ( .CLK(clk), .D(w_mem_inst__0w_mem_12__31_0__1_), .Q(w_mem_inst_w_mem_12__1_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_725 ( .CLK(clk), .D(w_mem_inst__0w_mem_12__31_0__2_), .Q(w_mem_inst_w_mem_12__2_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_726 ( .CLK(clk), .D(w_mem_inst__0w_mem_12__31_0__3_), .Q(w_mem_inst_w_mem_12__3_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_727 ( .CLK(clk), .D(w_mem_inst__0w_mem_12__31_0__4_), .Q(w_mem_inst_w_mem_12__4_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_728 ( .CLK(clk), .D(w_mem_inst__0w_mem_12__31_0__5_), .Q(w_mem_inst_w_mem_12__5_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_729 ( .CLK(clk), .D(w_mem_inst__0w_mem_12__31_0__6_), .Q(w_mem_inst_w_mem_12__6_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_73 ( .CLK(clk), .D(_0c_reg_31_0__8_), .Q(c_reg_8_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_730 ( .CLK(clk), .D(w_mem_inst__0w_mem_12__31_0__7_), .Q(w_mem_inst_w_mem_12__7_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_731 ( .CLK(clk), .D(w_mem_inst__0w_mem_12__31_0__8_), .Q(w_mem_inst_w_mem_12__8_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_732 ( .CLK(clk), .D(w_mem_inst__0w_mem_12__31_0__9_), .Q(w_mem_inst_w_mem_12__9_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_733 ( .CLK(clk), .D(w_mem_inst__0w_mem_12__31_0__10_), .Q(w_mem_inst_w_mem_12__10_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_734 ( .CLK(clk), .D(w_mem_inst__0w_mem_12__31_0__11_), .Q(w_mem_inst_w_mem_12__11_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_735 ( .CLK(clk), .D(w_mem_inst__0w_mem_12__31_0__12_), .Q(w_mem_inst_w_mem_12__12_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_736 ( .CLK(clk), .D(w_mem_inst__0w_mem_12__31_0__13_), .Q(w_mem_inst_w_mem_12__13_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_737 ( .CLK(clk), .D(w_mem_inst__0w_mem_12__31_0__14_), .Q(w_mem_inst_w_mem_12__14_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_738 ( .CLK(clk), .D(w_mem_inst__0w_mem_12__31_0__15_), .Q(w_mem_inst_w_mem_12__15_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_739 ( .CLK(clk), .D(w_mem_inst__0w_mem_12__31_0__16_), .Q(w_mem_inst_w_mem_12__16_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_74 ( .CLK(clk), .D(_0c_reg_31_0__9_), .Q(c_reg_9_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_740 ( .CLK(clk), .D(w_mem_inst__0w_mem_12__31_0__17_), .Q(w_mem_inst_w_mem_12__17_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_741 ( .CLK(clk), .D(w_mem_inst__0w_mem_12__31_0__18_), .Q(w_mem_inst_w_mem_12__18_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_742 ( .CLK(clk), .D(w_mem_inst__0w_mem_12__31_0__19_), .Q(w_mem_inst_w_mem_12__19_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_743 ( .CLK(clk), .D(w_mem_inst__0w_mem_12__31_0__20_), .Q(w_mem_inst_w_mem_12__20_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_744 ( .CLK(clk), .D(w_mem_inst__0w_mem_12__31_0__21_), .Q(w_mem_inst_w_mem_12__21_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_745 ( .CLK(clk), .D(w_mem_inst__0w_mem_12__31_0__22_), .Q(w_mem_inst_w_mem_12__22_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_746 ( .CLK(clk), .D(w_mem_inst__0w_mem_12__31_0__23_), .Q(w_mem_inst_w_mem_12__23_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_747 ( .CLK(clk), .D(w_mem_inst__0w_mem_12__31_0__24_), .Q(w_mem_inst_w_mem_12__24_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_748 ( .CLK(clk), .D(w_mem_inst__0w_mem_12__31_0__25_), .Q(w_mem_inst_w_mem_12__25_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_749 ( .CLK(clk), .D(w_mem_inst__0w_mem_12__31_0__26_), .Q(w_mem_inst_w_mem_12__26_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_75 ( .CLK(clk), .D(_0c_reg_31_0__10_), .Q(c_reg_10_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_750 ( .CLK(clk), .D(w_mem_inst__0w_mem_12__31_0__27_), .Q(w_mem_inst_w_mem_12__27_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_751 ( .CLK(clk), .D(w_mem_inst__0w_mem_12__31_0__28_), .Q(w_mem_inst_w_mem_12__28_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_752 ( .CLK(clk), .D(w_mem_inst__0w_mem_12__31_0__29_), .Q(w_mem_inst_w_mem_12__29_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_753 ( .CLK(clk), .D(w_mem_inst__0w_mem_12__31_0__30_), .Q(w_mem_inst_w_mem_12__30_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_754 ( .CLK(clk), .D(w_mem_inst__0w_mem_12__31_0__31_), .Q(w_mem_inst_w_mem_12__31_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_755 ( .CLK(clk), .D(w_mem_inst__0w_mem_13__31_0__0_), .Q(w_mem_inst_w_mem_13__0_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_756 ( .CLK(clk), .D(w_mem_inst__0w_mem_13__31_0__1_), .Q(w_mem_inst_w_mem_13__1_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_757 ( .CLK(clk), .D(w_mem_inst__0w_mem_13__31_0__2_), .Q(w_mem_inst_w_mem_13__2_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_758 ( .CLK(clk), .D(w_mem_inst__0w_mem_13__31_0__3_), .Q(w_mem_inst_w_mem_13__3_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_759 ( .CLK(clk), .D(w_mem_inst__0w_mem_13__31_0__4_), .Q(w_mem_inst_w_mem_13__4_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_76 ( .CLK(clk), .D(_0c_reg_31_0__11_), .Q(c_reg_11_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_760 ( .CLK(clk), .D(w_mem_inst__0w_mem_13__31_0__5_), .Q(w_mem_inst_w_mem_13__5_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_761 ( .CLK(clk), .D(w_mem_inst__0w_mem_13__31_0__6_), .Q(w_mem_inst_w_mem_13__6_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_762 ( .CLK(clk), .D(w_mem_inst__0w_mem_13__31_0__7_), .Q(w_mem_inst_w_mem_13__7_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_763 ( .CLK(clk), .D(w_mem_inst__0w_mem_13__31_0__8_), .Q(w_mem_inst_w_mem_13__8_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_764 ( .CLK(clk), .D(w_mem_inst__0w_mem_13__31_0__9_), .Q(w_mem_inst_w_mem_13__9_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_765 ( .CLK(clk), .D(w_mem_inst__0w_mem_13__31_0__10_), .Q(w_mem_inst_w_mem_13__10_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_766 ( .CLK(clk), .D(w_mem_inst__0w_mem_13__31_0__11_), .Q(w_mem_inst_w_mem_13__11_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_767 ( .CLK(clk), .D(w_mem_inst__0w_mem_13__31_0__12_), .Q(w_mem_inst_w_mem_13__12_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_768 ( .CLK(clk), .D(w_mem_inst__0w_mem_13__31_0__13_), .Q(w_mem_inst_w_mem_13__13_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_769 ( .CLK(clk), .D(w_mem_inst__0w_mem_13__31_0__14_), .Q(w_mem_inst_w_mem_13__14_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_77 ( .CLK(clk), .D(_0c_reg_31_0__12_), .Q(c_reg_12_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_770 ( .CLK(clk), .D(w_mem_inst__0w_mem_13__31_0__15_), .Q(w_mem_inst_w_mem_13__15_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_771 ( .CLK(clk), .D(w_mem_inst__0w_mem_13__31_0__16_), .Q(w_mem_inst_w_mem_13__16_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_772 ( .CLK(clk), .D(w_mem_inst__0w_mem_13__31_0__17_), .Q(w_mem_inst_w_mem_13__17_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_773 ( .CLK(clk), .D(w_mem_inst__0w_mem_13__31_0__18_), .Q(w_mem_inst_w_mem_13__18_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_774 ( .CLK(clk), .D(w_mem_inst__0w_mem_13__31_0__19_), .Q(w_mem_inst_w_mem_13__19_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_775 ( .CLK(clk), .D(w_mem_inst__0w_mem_13__31_0__20_), .Q(w_mem_inst_w_mem_13__20_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_776 ( .CLK(clk), .D(w_mem_inst__0w_mem_13__31_0__21_), .Q(w_mem_inst_w_mem_13__21_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_777 ( .CLK(clk), .D(w_mem_inst__0w_mem_13__31_0__22_), .Q(w_mem_inst_w_mem_13__22_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_778 ( .CLK(clk), .D(w_mem_inst__0w_mem_13__31_0__23_), .Q(w_mem_inst_w_mem_13__23_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_779 ( .CLK(clk), .D(w_mem_inst__0w_mem_13__31_0__24_), .Q(w_mem_inst_w_mem_13__24_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_78 ( .CLK(clk), .D(_0c_reg_31_0__13_), .Q(c_reg_13_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_780 ( .CLK(clk), .D(w_mem_inst__0w_mem_13__31_0__25_), .Q(w_mem_inst_w_mem_13__25_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_781 ( .CLK(clk), .D(w_mem_inst__0w_mem_13__31_0__26_), .Q(w_mem_inst_w_mem_13__26_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_782 ( .CLK(clk), .D(w_mem_inst__0w_mem_13__31_0__27_), .Q(w_mem_inst_w_mem_13__27_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_783 ( .CLK(clk), .D(w_mem_inst__0w_mem_13__31_0__28_), .Q(w_mem_inst_w_mem_13__28_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_784 ( .CLK(clk), .D(w_mem_inst__0w_mem_13__31_0__29_), .Q(w_mem_inst_w_mem_13__29_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_785 ( .CLK(clk), .D(w_mem_inst__0w_mem_13__31_0__30_), .Q(w_mem_inst_w_mem_13__30_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_786 ( .CLK(clk), .D(w_mem_inst__0w_mem_13__31_0__31_), .Q(w_mem_inst_w_mem_13__31_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_787 ( .CLK(clk), .D(w_mem_inst__0w_mem_14__31_0__0_), .Q(w_mem_inst_w_mem_14__0_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_788 ( .CLK(clk), .D(w_mem_inst__0w_mem_14__31_0__1_), .Q(w_mem_inst_w_mem_14__1_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_789 ( .CLK(clk), .D(w_mem_inst__0w_mem_14__31_0__2_), .Q(w_mem_inst_w_mem_14__2_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_79 ( .CLK(clk), .D(_0c_reg_31_0__14_), .Q(c_reg_14_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_790 ( .CLK(clk), .D(w_mem_inst__0w_mem_14__31_0__3_), .Q(w_mem_inst_w_mem_14__3_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_791 ( .CLK(clk), .D(w_mem_inst__0w_mem_14__31_0__4_), .Q(w_mem_inst_w_mem_14__4_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_792 ( .CLK(clk), .D(w_mem_inst__0w_mem_14__31_0__5_), .Q(w_mem_inst_w_mem_14__5_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_793 ( .CLK(clk), .D(w_mem_inst__0w_mem_14__31_0__6_), .Q(w_mem_inst_w_mem_14__6_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_794 ( .CLK(clk), .D(w_mem_inst__0w_mem_14__31_0__7_), .Q(w_mem_inst_w_mem_14__7_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_795 ( .CLK(clk), .D(w_mem_inst__0w_mem_14__31_0__8_), .Q(w_mem_inst_w_mem_14__8_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_796 ( .CLK(clk), .D(w_mem_inst__0w_mem_14__31_0__9_), .Q(w_mem_inst_w_mem_14__9_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_797 ( .CLK(clk), .D(w_mem_inst__0w_mem_14__31_0__10_), .Q(w_mem_inst_w_mem_14__10_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_798 ( .CLK(clk), .D(w_mem_inst__0w_mem_14__31_0__11_), .Q(w_mem_inst_w_mem_14__11_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_799 ( .CLK(clk), .D(w_mem_inst__0w_mem_14__31_0__12_), .Q(w_mem_inst_w_mem_14__12_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_8 ( .CLK(clk), .D(_0a_reg_31_0__7_), .Q(a_reg_7_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_80 ( .CLK(clk), .D(_0c_reg_31_0__15_), .Q(c_reg_15_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_800 ( .CLK(clk), .D(w_mem_inst__0w_mem_14__31_0__13_), .Q(w_mem_inst_w_mem_14__13_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_801 ( .CLK(clk), .D(w_mem_inst__0w_mem_14__31_0__14_), .Q(w_mem_inst_w_mem_14__14_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_802 ( .CLK(clk), .D(w_mem_inst__0w_mem_14__31_0__15_), .Q(w_mem_inst_w_mem_14__15_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_803 ( .CLK(clk), .D(w_mem_inst__0w_mem_14__31_0__16_), .Q(w_mem_inst_w_mem_14__16_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_804 ( .CLK(clk), .D(w_mem_inst__0w_mem_14__31_0__17_), .Q(w_mem_inst_w_mem_14__17_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_805 ( .CLK(clk), .D(w_mem_inst__0w_mem_14__31_0__18_), .Q(w_mem_inst_w_mem_14__18_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_806 ( .CLK(clk), .D(w_mem_inst__0w_mem_14__31_0__19_), .Q(w_mem_inst_w_mem_14__19_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_807 ( .CLK(clk), .D(w_mem_inst__0w_mem_14__31_0__20_), .Q(w_mem_inst_w_mem_14__20_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_808 ( .CLK(clk), .D(w_mem_inst__0w_mem_14__31_0__21_), .Q(w_mem_inst_w_mem_14__21_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_809 ( .CLK(clk), .D(w_mem_inst__0w_mem_14__31_0__22_), .Q(w_mem_inst_w_mem_14__22_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_81 ( .CLK(clk), .D(_0c_reg_31_0__16_), .Q(c_reg_16_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_810 ( .CLK(clk), .D(w_mem_inst__0w_mem_14__31_0__23_), .Q(w_mem_inst_w_mem_14__23_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_811 ( .CLK(clk), .D(w_mem_inst__0w_mem_14__31_0__24_), .Q(w_mem_inst_w_mem_14__24_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_812 ( .CLK(clk), .D(w_mem_inst__0w_mem_14__31_0__25_), .Q(w_mem_inst_w_mem_14__25_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_813 ( .CLK(clk), .D(w_mem_inst__0w_mem_14__31_0__26_), .Q(w_mem_inst_w_mem_14__26_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_814 ( .CLK(clk), .D(w_mem_inst__0w_mem_14__31_0__27_), .Q(w_mem_inst_w_mem_14__27_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_815 ( .CLK(clk), .D(w_mem_inst__0w_mem_14__31_0__28_), .Q(w_mem_inst_w_mem_14__28_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_816 ( .CLK(clk), .D(w_mem_inst__0w_mem_14__31_0__29_), .Q(w_mem_inst_w_mem_14__29_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_817 ( .CLK(clk), .D(w_mem_inst__0w_mem_14__31_0__30_), .Q(w_mem_inst_w_mem_14__30_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_818 ( .CLK(clk), .D(w_mem_inst__0w_mem_14__31_0__31_), .Q(w_mem_inst_w_mem_14__31_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_819 ( .CLK(clk), .D(w_mem_inst__0w_mem_15__31_0__0_), .Q(w_mem_inst_w_mem_15__0_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_82 ( .CLK(clk), .D(_0c_reg_31_0__17_), .Q(c_reg_17_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_820 ( .CLK(clk), .D(w_mem_inst__0w_mem_15__31_0__1_), .Q(w_mem_inst_w_mem_15__1_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_821 ( .CLK(clk), .D(w_mem_inst__0w_mem_15__31_0__2_), .Q(w_mem_inst_w_mem_15__2_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_822 ( .CLK(clk), .D(w_mem_inst__0w_mem_15__31_0__3_), .Q(w_mem_inst_w_mem_15__3_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_823 ( .CLK(clk), .D(w_mem_inst__0w_mem_15__31_0__4_), .Q(w_mem_inst_w_mem_15__4_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_824 ( .CLK(clk), .D(w_mem_inst__0w_mem_15__31_0__5_), .Q(w_mem_inst_w_mem_15__5_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_825 ( .CLK(clk), .D(w_mem_inst__0w_mem_15__31_0__6_), .Q(w_mem_inst_w_mem_15__6_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_826 ( .CLK(clk), .D(w_mem_inst__0w_mem_15__31_0__7_), .Q(w_mem_inst_w_mem_15__7_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_827 ( .CLK(clk), .D(w_mem_inst__0w_mem_15__31_0__8_), .Q(w_mem_inst_w_mem_15__8_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_828 ( .CLK(clk), .D(w_mem_inst__0w_mem_15__31_0__9_), .Q(w_mem_inst_w_mem_15__9_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_829 ( .CLK(clk), .D(w_mem_inst__0w_mem_15__31_0__10_), .Q(w_mem_inst_w_mem_15__10_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_83 ( .CLK(clk), .D(_0c_reg_31_0__18_), .Q(c_reg_18_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_830 ( .CLK(clk), .D(w_mem_inst__0w_mem_15__31_0__11_), .Q(w_mem_inst_w_mem_15__11_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_831 ( .CLK(clk), .D(w_mem_inst__0w_mem_15__31_0__12_), .Q(w_mem_inst_w_mem_15__12_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_832 ( .CLK(clk), .D(w_mem_inst__0w_mem_15__31_0__13_), .Q(w_mem_inst_w_mem_15__13_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_833 ( .CLK(clk), .D(w_mem_inst__0w_mem_15__31_0__14_), .Q(w_mem_inst_w_mem_15__14_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_834 ( .CLK(clk), .D(w_mem_inst__0w_mem_15__31_0__15_), .Q(w_mem_inst_w_mem_15__15_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_835 ( .CLK(clk), .D(w_mem_inst__0w_mem_15__31_0__16_), .Q(w_mem_inst_w_mem_15__16_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_836 ( .CLK(clk), .D(w_mem_inst__0w_mem_15__31_0__17_), .Q(w_mem_inst_w_mem_15__17_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_837 ( .CLK(clk), .D(w_mem_inst__0w_mem_15__31_0__18_), .Q(w_mem_inst_w_mem_15__18_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_838 ( .CLK(clk), .D(w_mem_inst__0w_mem_15__31_0__19_), .Q(w_mem_inst_w_mem_15__19_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_839 ( .CLK(clk), .D(w_mem_inst__0w_mem_15__31_0__20_), .Q(w_mem_inst_w_mem_15__20_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_84 ( .CLK(clk), .D(_0c_reg_31_0__19_), .Q(c_reg_19_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_840 ( .CLK(clk), .D(w_mem_inst__0w_mem_15__31_0__21_), .Q(w_mem_inst_w_mem_15__21_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_841 ( .CLK(clk), .D(w_mem_inst__0w_mem_15__31_0__22_), .Q(w_mem_inst_w_mem_15__22_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_842 ( .CLK(clk), .D(w_mem_inst__0w_mem_15__31_0__23_), .Q(w_mem_inst_w_mem_15__23_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_843 ( .CLK(clk), .D(w_mem_inst__0w_mem_15__31_0__24_), .Q(w_mem_inst_w_mem_15__24_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_844 ( .CLK(clk), .D(w_mem_inst__0w_mem_15__31_0__25_), .Q(w_mem_inst_w_mem_15__25_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_845 ( .CLK(clk), .D(w_mem_inst__0w_mem_15__31_0__26_), .Q(w_mem_inst_w_mem_15__26_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_846 ( .CLK(clk), .D(w_mem_inst__0w_mem_15__31_0__27_), .Q(w_mem_inst_w_mem_15__27_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_847 ( .CLK(clk), .D(w_mem_inst__0w_mem_15__31_0__28_), .Q(w_mem_inst_w_mem_15__28_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_848 ( .CLK(clk), .D(w_mem_inst__0w_mem_15__31_0__29_), .Q(w_mem_inst_w_mem_15__29_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_849 ( .CLK(clk), .D(w_mem_inst__0w_mem_15__31_0__30_), .Q(w_mem_inst_w_mem_15__30_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_85 ( .CLK(clk), .D(_0c_reg_31_0__20_), .Q(c_reg_20_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_850 ( .CLK(clk), .D(w_mem_inst__0w_mem_15__31_0__31_), .Q(w_mem_inst_w_mem_15__31_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_86 ( .CLK(clk), .D(_0c_reg_31_0__21_), .Q(c_reg_21_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_87 ( .CLK(clk), .D(_0c_reg_31_0__22_), .Q(c_reg_22_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_88 ( .CLK(clk), .D(_0c_reg_31_0__23_), .Q(c_reg_23_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_89 ( .CLK(clk), .D(_0c_reg_31_0__24_), .Q(c_reg_24_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_9 ( .CLK(clk), .D(_0a_reg_31_0__8_), .Q(a_reg_8_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_90 ( .CLK(clk), .D(_0c_reg_31_0__25_), .Q(c_reg_25_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_91 ( .CLK(clk), .D(_0c_reg_31_0__26_), .Q(c_reg_26_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_92 ( .CLK(clk), .D(_0c_reg_31_0__27_), .Q(c_reg_27_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_93 ( .CLK(clk), .D(_0c_reg_31_0__28_), .Q(c_reg_28_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_94 ( .CLK(clk), .D(_0c_reg_31_0__29_), .Q(c_reg_29_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_95 ( .CLK(clk), .D(_0c_reg_31_0__30_), .Q(c_reg_30_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_96 ( .CLK(clk), .D(_0c_reg_31_0__31_), .Q(c_reg_31_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_97 ( .CLK(clk), .D(_0d_reg_31_0__0_), .Q(d_reg_0_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_98 ( .CLK(clk), .D(_0d_reg_31_0__1_), .Q(d_reg_1_), .R(reset_n), .S(1'h1));
DFFSR DFFSR_99 ( .CLK(clk), .D(_0d_reg_31_0__2_), .Q(d_reg_2_), .R(reset_n), .S(1'h1));
INVX1 INVX1_1 ( .A(digest_update), .Y(_abc_15497_new_n698_));
INVX1 INVX1_10 ( .A(_abc_15497_new_n731_), .Y(_abc_15497_new_n732_));
INVX1 INVX1_100 ( .A(_abc_15497_new_n1176_), .Y(_abc_15497_new_n1177_));
INVX1 INVX1_1000 ( .A(_abc_15497_new_n5887_), .Y(_abc_15497_new_n5888_));
INVX1 INVX1_1001 ( .A(_abc_15497_new_n5890_), .Y(_abc_15497_new_n5891_));
INVX1 INVX1_1002 ( .A(_abc_15497_new_n5893_), .Y(_abc_15497_new_n5894_));
INVX1 INVX1_1003 ( .A(w_28_), .Y(_abc_15497_new_n5896_));
INVX1 INVX1_1004 ( .A(_abc_15497_new_n5898_), .Y(_abc_15497_new_n5899_));
INVX1 INVX1_1005 ( .A(_abc_15497_new_n5900_), .Y(_abc_15497_new_n5901_));
INVX1 INVX1_1006 ( .A(_abc_15497_new_n5904_), .Y(_abc_15497_new_n5905_));
INVX1 INVX1_1007 ( .A(_abc_15497_new_n5906_), .Y(_abc_15497_new_n5907_));
INVX1 INVX1_1008 ( .A(_abc_15497_new_n5910_), .Y(_abc_15497_new_n5911_));
INVX1 INVX1_1009 ( .A(_abc_15497_new_n5913_), .Y(_abc_15497_new_n5914_));
INVX1 INVX1_101 ( .A(_abc_15497_new_n1180_), .Y(_abc_15497_new_n1181_));
INVX1 INVX1_1010 ( .A(_abc_15497_new_n5916_), .Y(_abc_15497_new_n5917_));
INVX1 INVX1_1011 ( .A(_abc_15497_new_n5918_), .Y(_abc_15497_new_n5919_));
INVX1 INVX1_1012 ( .A(_abc_15497_new_n5924_), .Y(_abc_15497_new_n5925_));
INVX1 INVX1_1013 ( .A(_abc_15497_new_n5926_), .Y(_abc_15497_new_n5927_));
INVX1 INVX1_1014 ( .A(_abc_15497_new_n5929_), .Y(_abc_15497_new_n5930_));
INVX1 INVX1_1015 ( .A(_abc_15497_new_n5939_), .Y(_abc_15497_new_n5940_));
INVX1 INVX1_1016 ( .A(b_reg_29_), .Y(_abc_15497_new_n5943_));
INVX1 INVX1_1017 ( .A(d_reg_29_), .Y(_abc_15497_new_n5947_));
INVX1 INVX1_1018 ( .A(_abc_15497_new_n5942_), .Y(_abc_15497_new_n5948_));
INVX1 INVX1_1019 ( .A(_abc_15497_new_n5951_), .Y(_abc_15497_new_n5952_));
INVX1 INVX1_102 ( .A(_abc_15497_new_n1182_), .Y(_abc_15497_new_n1183_));
INVX1 INVX1_1020 ( .A(_abc_15497_new_n5956_), .Y(_abc_15497_new_n5957_));
INVX1 INVX1_1021 ( .A(_abc_15497_new_n5960_), .Y(_abc_15497_new_n5961_));
INVX1 INVX1_1022 ( .A(_abc_15497_new_n5962_), .Y(_abc_15497_new_n5963_));
INVX1 INVX1_1023 ( .A(w_29_), .Y(_abc_15497_new_n5966_));
INVX1 INVX1_1024 ( .A(_abc_15497_new_n5968_), .Y(_abc_15497_new_n5969_));
INVX1 INVX1_1025 ( .A(_abc_15497_new_n5970_), .Y(_abc_15497_new_n5971_));
INVX1 INVX1_1026 ( .A(_abc_15497_new_n5974_), .Y(_abc_15497_new_n5975_));
INVX1 INVX1_1027 ( .A(_abc_15497_new_n5976_), .Y(_abc_15497_new_n5977_));
INVX1 INVX1_1028 ( .A(_abc_15497_new_n5980_), .Y(_abc_15497_new_n5981_));
INVX1 INVX1_1029 ( .A(_abc_15497_new_n5983_), .Y(_abc_15497_new_n5984_));
INVX1 INVX1_103 ( .A(_abc_15497_new_n1188_), .Y(_abc_15497_new_n1189_));
INVX1 INVX1_1030 ( .A(_abc_15497_new_n5986_), .Y(_abc_15497_new_n5987_));
INVX1 INVX1_1031 ( .A(_abc_15497_new_n5990_), .Y(_abc_15497_new_n5991_));
INVX1 INVX1_1032 ( .A(_abc_15497_new_n5994_), .Y(_abc_15497_new_n5995_));
INVX1 INVX1_1033 ( .A(_abc_15497_new_n5938_), .Y(_abc_15497_new_n5998_));
INVX1 INVX1_1034 ( .A(_abc_15497_new_n5996_), .Y(_abc_15497_new_n5999_));
INVX1 INVX1_1035 ( .A(_abc_15497_new_n6007_), .Y(_abc_15497_new_n6008_));
INVX1 INVX1_1036 ( .A(_abc_15497_new_n6011_), .Y(_abc_15497_new_n6012_));
INVX1 INVX1_1037 ( .A(_abc_15497_new_n6013_), .Y(_abc_15497_new_n6014_));
INVX1 INVX1_1038 ( .A(b_reg_30_), .Y(_abc_15497_new_n6018_));
INVX1 INVX1_1039 ( .A(d_reg_30_), .Y(_abc_15497_new_n6022_));
INVX1 INVX1_104 ( .A(_abc_15497_new_n1192_), .Y(_abc_15497_new_n1193_));
INVX1 INVX1_1040 ( .A(_abc_15497_new_n6017_), .Y(_abc_15497_new_n6023_));
INVX1 INVX1_1041 ( .A(_abc_15497_new_n6026_), .Y(_abc_15497_new_n6027_));
INVX1 INVX1_1042 ( .A(_abc_15497_new_n6031_), .Y(_abc_15497_new_n6032_));
INVX1 INVX1_1043 ( .A(_abc_15497_new_n6035_), .Y(_abc_15497_new_n6036_));
INVX1 INVX1_1044 ( .A(_abc_15497_new_n6037_), .Y(_abc_15497_new_n6038_));
INVX1 INVX1_1045 ( .A(w_30_), .Y(_abc_15497_new_n6041_));
INVX1 INVX1_1046 ( .A(_abc_15497_new_n6043_), .Y(_abc_15497_new_n6044_));
INVX1 INVX1_1047 ( .A(_abc_15497_new_n6045_), .Y(_abc_15497_new_n6046_));
INVX1 INVX1_1048 ( .A(_abc_15497_new_n6049_), .Y(_abc_15497_new_n6050_));
INVX1 INVX1_1049 ( .A(_abc_15497_new_n6051_), .Y(_abc_15497_new_n6052_));
INVX1 INVX1_105 ( .A(_abc_15497_new_n1199_), .Y(_abc_15497_new_n1200_));
INVX1 INVX1_1050 ( .A(_abc_15497_new_n6055_), .Y(_abc_15497_new_n6056_));
INVX1 INVX1_1051 ( .A(_abc_15497_new_n6058_), .Y(_abc_15497_new_n6059_));
INVX1 INVX1_1052 ( .A(_abc_15497_new_n6061_), .Y(_abc_15497_new_n6062_));
INVX1 INVX1_1053 ( .A(_abc_15497_new_n6063_), .Y(_abc_15497_new_n6064_));
INVX1 INVX1_1054 ( .A(_abc_15497_new_n6069_), .Y(_abc_15497_new_n6070_));
INVX1 INVX1_1055 ( .A(_abc_15497_new_n6071_), .Y(_abc_15497_new_n6072_));
INVX1 INVX1_1056 ( .A(_abc_15497_new_n6081_), .Y(_abc_15497_new_n6082_));
INVX1 INVX1_1057 ( .A(_abc_15497_new_n6083_), .Y(_abc_15497_new_n6084_));
INVX1 INVX1_1058 ( .A(_abc_15497_new_n6085_), .Y(_abc_15497_new_n6086_));
INVX1 INVX1_1059 ( .A(_abc_15497_new_n6087_), .Y(_abc_15497_new_n6088_));
INVX1 INVX1_106 ( .A(_abc_15497_new_n1197_), .Y(_abc_15497_new_n1203_));
INVX1 INVX1_1060 ( .A(d_reg_31_), .Y(_abc_15497_new_n6089_));
INVX1 INVX1_1061 ( .A(_abc_15497_new_n6093_), .Y(_abc_15497_new_n6094_));
INVX1 INVX1_1062 ( .A(_abc_15497_new_n6096_), .Y(_abc_15497_new_n6097_));
INVX1 INVX1_1063 ( .A(_abc_15497_new_n6106_), .Y(_abc_15497_new_n6107_));
INVX1 INVX1_1064 ( .A(_abc_15497_new_n6108_), .Y(_abc_15497_new_n6109_));
INVX1 INVX1_1065 ( .A(_abc_15497_new_n6111_), .Y(_abc_15497_new_n6112_));
INVX1 INVX1_1066 ( .A(_abc_15497_new_n6114_), .Y(_abc_15497_new_n6115_));
INVX1 INVX1_1067 ( .A(_abc_15497_new_n6117_), .Y(_abc_15497_new_n6118_));
INVX1 INVX1_1068 ( .A(_abc_15497_new_n6121_), .Y(_abc_15497_new_n6122_));
INVX1 INVX1_1069 ( .A(_abc_15497_new_n6126_), .Y(_abc_15497_new_n6127_));
INVX1 INVX1_107 ( .A(_abc_15497_new_n1201_), .Y(_abc_15497_new_n1204_));
INVX1 INVX1_1070 ( .A(_abc_15497_new_n6129_), .Y(_abc_15497_new_n6131_));
INVX1 INVX1_1071 ( .A(_abc_15497_new_n6134_), .Y(_abc_15497_new_n6135_));
INVX1 INVX1_1072 ( .A(_abc_15497_new_n6137_), .Y(_abc_15497_new_n6139_));
INVX1 INVX1_1073 ( .A(_abc_15497_new_n2006_), .Y(_abc_15497_new_n6153_));
INVX1 INVX1_1074 ( .A(_abc_15497_new_n6151_), .Y(_abc_15497_new_n6154_));
INVX1 INVX1_1075 ( .A(round_ctr_reg_0_), .Y(_abc_15497_new_n6161_));
INVX1 INVX1_1076 ( .A(_abc_15497_new_n6148_), .Y(_abc_15497_new_n6166_));
INVX1 INVX1_1077 ( .A(_abc_15497_new_n6172_), .Y(_abc_15497_new_n6173_));
INVX1 INVX1_1078 ( .A(_abc_15497_new_n2013_), .Y(_abc_15497_new_n6178_));
INVX1 INVX1_1079 ( .A(_abc_15497_new_n6182_), .Y(_abc_15497_new_n6183_));
INVX1 INVX1_108 ( .A(_abc_15497_new_n1212_), .Y(_abc_15497_new_n1213_));
INVX1 INVX1_1080 ( .A(_abc_15497_new_n6187_), .Y(_abc_15497_new_n6188_));
INVX1 INVX1_1081 ( .A(_abc_15497_new_n6193_), .Y(_abc_15497_new_n6194_));
INVX1 INVX1_1082 ( .A(_abc_15497_new_n6217_), .Y(_abc_15497_new_n6219_));
INVX1 INVX1_1083 ( .A(_abc_15497_new_n6231_), .Y(_abc_15497_new_n6233_));
INVX1 INVX1_1084 ( .A(_abc_15497_new_n6239_), .Y(_abc_15497_new_n6240_));
INVX1 INVX1_1085 ( .A(_abc_15497_new_n6245_), .Y(_abc_15497_new_n6246_));
INVX1 INVX1_1086 ( .A(_abc_15497_new_n807_), .Y(_abc_15497_new_n6248_));
INVX1 INVX1_1087 ( .A(_abc_15497_new_n6256_), .Y(_abc_15497_new_n6257_));
INVX1 INVX1_1088 ( .A(_abc_15497_new_n6262_), .Y(_abc_15497_new_n6263_));
INVX1 INVX1_1089 ( .A(_abc_15497_new_n842_), .Y(_abc_15497_new_n6265_));
INVX1 INVX1_109 ( .A(_abc_15497_new_n1198_), .Y(_abc_15497_new_n1215_));
INVX1 INVX1_1090 ( .A(_abc_15497_new_n6271_), .Y(_abc_15497_new_n6272_));
INVX1 INVX1_1091 ( .A(_abc_15497_new_n6277_), .Y(_abc_15497_new_n6278_));
INVX1 INVX1_1092 ( .A(_abc_15497_new_n791_), .Y(_abc_15497_new_n6280_));
INVX1 INVX1_1093 ( .A(_abc_15497_new_n6287_), .Y(_abc_15497_new_n6288_));
INVX1 INVX1_1094 ( .A(_abc_15497_new_n6294_), .Y(_abc_15497_new_n6295_));
INVX1 INVX1_1095 ( .A(_abc_15497_new_n6304_), .Y(_abc_15497_new_n6305_));
INVX1 INVX1_1096 ( .A(_abc_15497_new_n6310_), .Y(_abc_15497_new_n6311_));
INVX1 INVX1_1097 ( .A(_abc_15497_new_n761_), .Y(_abc_15497_new_n6313_));
INVX1 INVX1_1098 ( .A(_abc_15497_new_n6321_), .Y(_abc_15497_new_n6322_));
INVX1 INVX1_1099 ( .A(_abc_15497_new_n6326_), .Y(_abc_15497_new_n6327_));
INVX1 INVX1_11 ( .A(_abc_15497_new_n735_), .Y(_abc_15497_new_n736_));
INVX1 INVX1_110 ( .A(_abc_15497_new_n1218_), .Y(_abc_15497_new_n1219_));
INVX1 INVX1_1100 ( .A(_abc_15497_new_n6338_), .Y(_abc_15497_new_n6339_));
INVX1 INVX1_1101 ( .A(_abc_15497_new_n734_), .Y(_abc_15497_new_n6345_));
INVX1 INVX1_1102 ( .A(_abc_15497_new_n6343_), .Y(_abc_15497_new_n6346_));
INVX1 INVX1_1103 ( .A(_abc_15497_new_n6355_), .Y(_abc_15497_new_n6356_));
INVX1 INVX1_1104 ( .A(_abc_15497_new_n6362_), .Y(_abc_15497_new_n6363_));
INVX1 INVX1_1105 ( .A(_abc_15497_new_n6373_), .Y(_abc_15497_new_n6374_));
INVX1 INVX1_1106 ( .A(_abc_15497_new_n6378_), .Y(_abc_15497_new_n6379_));
INVX1 INVX1_1107 ( .A(_abc_15497_new_n706_), .Y(_abc_15497_new_n6381_));
INVX1 INVX1_1108 ( .A(_abc_15497_new_n6389_), .Y(_abc_15497_new_n6390_));
INVX1 INVX1_1109 ( .A(_abc_15497_new_n6395_), .Y(_abc_15497_new_n6396_));
INVX1 INVX1_111 ( .A(_abc_15497_new_n1221_), .Y(_abc_15497_new_n1222_));
INVX1 INVX1_1110 ( .A(_abc_15497_new_n863_), .Y(_abc_15497_new_n6398_));
INVX1 INVX1_1111 ( .A(w_mem_inst__abc_21203_new_n1586_), .Y(w_mem_inst__abc_21203_new_n1587_));
INVX1 INVX1_1112 ( .A(w_mem_inst_w_mem_8__31_), .Y(w_mem_inst__abc_21203_new_n1588_));
INVX1 INVX1_1113 ( .A(w_mem_inst_w_mem_13__31_), .Y(w_mem_inst__abc_21203_new_n1590_));
INVX1 INVX1_1114 ( .A(w_mem_inst__abc_21203_new_n1592_), .Y(w_mem_inst__abc_21203_new_n1593_));
INVX1 INVX1_1115 ( .A(w_mem_inst__abc_21203_new_n1595_), .Y(w_mem_inst__abc_21203_new_n1596_));
INVX1 INVX1_1116 ( .A(w_mem_inst__abc_21203_new_n1597_), .Y(w_mem_inst__abc_21203_new_n1599_));
INVX1 INVX1_1117 ( .A(w_mem_inst_w_ctr_reg_1_), .Y(w_mem_inst__abc_21203_new_n1603_));
INVX1 INVX1_1118 ( .A(w_mem_inst_w_ctr_reg_3_), .Y(w_mem_inst__abc_21203_new_n1605_));
INVX1 INVX1_1119 ( .A(w_mem_inst_w_ctr_reg_0_), .Y(w_mem_inst__abc_21203_new_n1610_));
INVX1 INVX1_112 ( .A(_abc_15497_new_n1230_), .Y(_abc_15497_new_n1231_));
INVX1 INVX1_1120 ( .A(w_mem_inst_w_ctr_reg_2_), .Y(w_mem_inst__abc_21203_new_n1612_));
INVX1 INVX1_1121 ( .A(w_mem_inst_w_mem_13__0_), .Y(w_mem_inst__abc_21203_new_n1664_));
INVX1 INVX1_1122 ( .A(w_mem_inst_w_mem_8__0_), .Y(w_mem_inst__abc_21203_new_n1666_));
INVX1 INVX1_1123 ( .A(w_mem_inst__abc_21203_new_n1668_), .Y(w_mem_inst__abc_21203_new_n1669_));
INVX1 INVX1_1124 ( .A(w_mem_inst__abc_21203_new_n1671_), .Y(w_mem_inst__abc_21203_new_n1672_));
INVX1 INVX1_1125 ( .A(w_mem_inst__abc_21203_new_n1673_), .Y(w_mem_inst__abc_21203_new_n1675_));
INVX1 INVX1_1126 ( .A(w_mem_inst_w_mem_13__1_), .Y(w_mem_inst__abc_21203_new_n1712_));
INVX1 INVX1_1127 ( .A(w_mem_inst_w_mem_8__1_), .Y(w_mem_inst__abc_21203_new_n1714_));
INVX1 INVX1_1128 ( .A(w_mem_inst__abc_21203_new_n1716_), .Y(w_mem_inst__abc_21203_new_n1717_));
INVX1 INVX1_1129 ( .A(w_mem_inst__abc_21203_new_n1719_), .Y(w_mem_inst__abc_21203_new_n1720_));
INVX1 INVX1_113 ( .A(_abc_15497_new_n1228_), .Y(_abc_15497_new_n1234_));
INVX1 INVX1_1130 ( .A(w_mem_inst__abc_21203_new_n1721_), .Y(w_mem_inst__abc_21203_new_n1723_));
INVX1 INVX1_1131 ( .A(w_mem_inst_w_mem_13__2_), .Y(w_mem_inst__abc_21203_new_n1760_));
INVX1 INVX1_1132 ( .A(w_mem_inst_w_mem_8__2_), .Y(w_mem_inst__abc_21203_new_n1762_));
INVX1 INVX1_1133 ( .A(w_mem_inst__abc_21203_new_n1764_), .Y(w_mem_inst__abc_21203_new_n1765_));
INVX1 INVX1_1134 ( .A(w_mem_inst__abc_21203_new_n1767_), .Y(w_mem_inst__abc_21203_new_n1768_));
INVX1 INVX1_1135 ( .A(w_mem_inst__abc_21203_new_n1769_), .Y(w_mem_inst__abc_21203_new_n1771_));
INVX1 INVX1_1136 ( .A(w_mem_inst_w_mem_13__3_), .Y(w_mem_inst__abc_21203_new_n1808_));
INVX1 INVX1_1137 ( .A(w_mem_inst_w_mem_8__3_), .Y(w_mem_inst__abc_21203_new_n1810_));
INVX1 INVX1_1138 ( .A(w_mem_inst__abc_21203_new_n1812_), .Y(w_mem_inst__abc_21203_new_n1813_));
INVX1 INVX1_1139 ( .A(w_mem_inst__abc_21203_new_n1815_), .Y(w_mem_inst__abc_21203_new_n1816_));
INVX1 INVX1_114 ( .A(_abc_15497_new_n1232_), .Y(_abc_15497_new_n1235_));
INVX1 INVX1_1140 ( .A(w_mem_inst__abc_21203_new_n1817_), .Y(w_mem_inst__abc_21203_new_n1819_));
INVX1 INVX1_1141 ( .A(w_mem_inst_w_mem_13__4_), .Y(w_mem_inst__abc_21203_new_n1856_));
INVX1 INVX1_1142 ( .A(w_mem_inst_w_mem_8__4_), .Y(w_mem_inst__abc_21203_new_n1858_));
INVX1 INVX1_1143 ( .A(w_mem_inst__abc_21203_new_n1860_), .Y(w_mem_inst__abc_21203_new_n1861_));
INVX1 INVX1_1144 ( .A(w_mem_inst__abc_21203_new_n1863_), .Y(w_mem_inst__abc_21203_new_n1864_));
INVX1 INVX1_1145 ( .A(w_mem_inst__abc_21203_new_n1865_), .Y(w_mem_inst__abc_21203_new_n1867_));
INVX1 INVX1_1146 ( .A(w_mem_inst_w_mem_13__5_), .Y(w_mem_inst__abc_21203_new_n1904_));
INVX1 INVX1_1147 ( .A(w_mem_inst_w_mem_8__5_), .Y(w_mem_inst__abc_21203_new_n1906_));
INVX1 INVX1_1148 ( .A(w_mem_inst__abc_21203_new_n1908_), .Y(w_mem_inst__abc_21203_new_n1909_));
INVX1 INVX1_1149 ( .A(w_mem_inst__abc_21203_new_n1911_), .Y(w_mem_inst__abc_21203_new_n1912_));
INVX1 INVX1_115 ( .A(_abc_15497_new_n1249_), .Y(_abc_15497_new_n1250_));
INVX1 INVX1_1150 ( .A(w_mem_inst__abc_21203_new_n1913_), .Y(w_mem_inst__abc_21203_new_n1915_));
INVX1 INVX1_1151 ( .A(w_mem_inst_w_mem_13__6_), .Y(w_mem_inst__abc_21203_new_n1952_));
INVX1 INVX1_1152 ( .A(w_mem_inst_w_mem_8__6_), .Y(w_mem_inst__abc_21203_new_n1954_));
INVX1 INVX1_1153 ( .A(w_mem_inst__abc_21203_new_n1956_), .Y(w_mem_inst__abc_21203_new_n1957_));
INVX1 INVX1_1154 ( .A(w_mem_inst__abc_21203_new_n1959_), .Y(w_mem_inst__abc_21203_new_n1960_));
INVX1 INVX1_1155 ( .A(w_mem_inst__abc_21203_new_n1961_), .Y(w_mem_inst__abc_21203_new_n1963_));
INVX1 INVX1_1156 ( .A(w_mem_inst_w_mem_13__7_), .Y(w_mem_inst__abc_21203_new_n2000_));
INVX1 INVX1_1157 ( .A(w_mem_inst_w_mem_8__7_), .Y(w_mem_inst__abc_21203_new_n2002_));
INVX1 INVX1_1158 ( .A(w_mem_inst__abc_21203_new_n2004_), .Y(w_mem_inst__abc_21203_new_n2005_));
INVX1 INVX1_1159 ( .A(w_mem_inst__abc_21203_new_n2007_), .Y(w_mem_inst__abc_21203_new_n2008_));
INVX1 INVX1_116 ( .A(_abc_15497_new_n1258_), .Y(_abc_15497_new_n1259_));
INVX1 INVX1_1160 ( .A(w_mem_inst__abc_21203_new_n2009_), .Y(w_mem_inst__abc_21203_new_n2011_));
INVX1 INVX1_1161 ( .A(w_mem_inst_w_mem_13__8_), .Y(w_mem_inst__abc_21203_new_n2048_));
INVX1 INVX1_1162 ( .A(w_mem_inst_w_mem_8__8_), .Y(w_mem_inst__abc_21203_new_n2050_));
INVX1 INVX1_1163 ( .A(w_mem_inst__abc_21203_new_n2052_), .Y(w_mem_inst__abc_21203_new_n2053_));
INVX1 INVX1_1164 ( .A(w_mem_inst__abc_21203_new_n2055_), .Y(w_mem_inst__abc_21203_new_n2056_));
INVX1 INVX1_1165 ( .A(w_mem_inst__abc_21203_new_n2057_), .Y(w_mem_inst__abc_21203_new_n2059_));
INVX1 INVX1_1166 ( .A(w_mem_inst_w_mem_13__9_), .Y(w_mem_inst__abc_21203_new_n2096_));
INVX1 INVX1_1167 ( .A(w_mem_inst_w_mem_8__9_), .Y(w_mem_inst__abc_21203_new_n2098_));
INVX1 INVX1_1168 ( .A(w_mem_inst__abc_21203_new_n2100_), .Y(w_mem_inst__abc_21203_new_n2101_));
INVX1 INVX1_1169 ( .A(w_mem_inst__abc_21203_new_n2103_), .Y(w_mem_inst__abc_21203_new_n2104_));
INVX1 INVX1_117 ( .A(_abc_15497_new_n1262_), .Y(_abc_15497_new_n1263_));
INVX1 INVX1_1170 ( .A(w_mem_inst__abc_21203_new_n2105_), .Y(w_mem_inst__abc_21203_new_n2107_));
INVX1 INVX1_1171 ( .A(w_mem_inst_w_mem_13__10_), .Y(w_mem_inst__abc_21203_new_n2144_));
INVX1 INVX1_1172 ( .A(w_mem_inst_w_mem_8__10_), .Y(w_mem_inst__abc_21203_new_n2146_));
INVX1 INVX1_1173 ( .A(w_mem_inst__abc_21203_new_n2148_), .Y(w_mem_inst__abc_21203_new_n2149_));
INVX1 INVX1_1174 ( .A(w_mem_inst__abc_21203_new_n2151_), .Y(w_mem_inst__abc_21203_new_n2152_));
INVX1 INVX1_1175 ( .A(w_mem_inst__abc_21203_new_n2153_), .Y(w_mem_inst__abc_21203_new_n2155_));
INVX1 INVX1_1176 ( .A(w_mem_inst_w_mem_13__11_), .Y(w_mem_inst__abc_21203_new_n2192_));
INVX1 INVX1_1177 ( .A(w_mem_inst_w_mem_8__11_), .Y(w_mem_inst__abc_21203_new_n2194_));
INVX1 INVX1_1178 ( .A(w_mem_inst__abc_21203_new_n2196_), .Y(w_mem_inst__abc_21203_new_n2197_));
INVX1 INVX1_1179 ( .A(w_mem_inst__abc_21203_new_n2199_), .Y(w_mem_inst__abc_21203_new_n2200_));
INVX1 INVX1_118 ( .A(_abc_15497_new_n1267_), .Y(_abc_15497_new_n1268_));
INVX1 INVX1_1180 ( .A(w_mem_inst__abc_21203_new_n2201_), .Y(w_mem_inst__abc_21203_new_n2203_));
INVX1 INVX1_1181 ( .A(w_mem_inst_w_mem_13__12_), .Y(w_mem_inst__abc_21203_new_n2240_));
INVX1 INVX1_1182 ( .A(w_mem_inst_w_mem_8__12_), .Y(w_mem_inst__abc_21203_new_n2242_));
INVX1 INVX1_1183 ( .A(w_mem_inst__abc_21203_new_n2244_), .Y(w_mem_inst__abc_21203_new_n2245_));
INVX1 INVX1_1184 ( .A(w_mem_inst__abc_21203_new_n2247_), .Y(w_mem_inst__abc_21203_new_n2248_));
INVX1 INVX1_1185 ( .A(w_mem_inst__abc_21203_new_n2249_), .Y(w_mem_inst__abc_21203_new_n2251_));
INVX1 INVX1_1186 ( .A(w_mem_inst_w_mem_13__13_), .Y(w_mem_inst__abc_21203_new_n2288_));
INVX1 INVX1_1187 ( .A(w_mem_inst_w_mem_8__13_), .Y(w_mem_inst__abc_21203_new_n2290_));
INVX1 INVX1_1188 ( .A(w_mem_inst__abc_21203_new_n2292_), .Y(w_mem_inst__abc_21203_new_n2293_));
INVX1 INVX1_1189 ( .A(w_mem_inst__abc_21203_new_n2295_), .Y(w_mem_inst__abc_21203_new_n2296_));
INVX1 INVX1_119 ( .A(_abc_15497_new_n1270_), .Y(_abc_15497_new_n1271_));
INVX1 INVX1_1190 ( .A(w_mem_inst__abc_21203_new_n2297_), .Y(w_mem_inst__abc_21203_new_n2299_));
INVX1 INVX1_1191 ( .A(w_mem_inst_w_mem_13__14_), .Y(w_mem_inst__abc_21203_new_n2336_));
INVX1 INVX1_1192 ( .A(w_mem_inst_w_mem_8__14_), .Y(w_mem_inst__abc_21203_new_n2338_));
INVX1 INVX1_1193 ( .A(w_mem_inst__abc_21203_new_n2340_), .Y(w_mem_inst__abc_21203_new_n2341_));
INVX1 INVX1_1194 ( .A(w_mem_inst__abc_21203_new_n2343_), .Y(w_mem_inst__abc_21203_new_n2344_));
INVX1 INVX1_1195 ( .A(w_mem_inst__abc_21203_new_n2345_), .Y(w_mem_inst__abc_21203_new_n2347_));
INVX1 INVX1_1196 ( .A(w_mem_inst_w_mem_13__15_), .Y(w_mem_inst__abc_21203_new_n2384_));
INVX1 INVX1_1197 ( .A(w_mem_inst_w_mem_8__15_), .Y(w_mem_inst__abc_21203_new_n2386_));
INVX1 INVX1_1198 ( .A(w_mem_inst__abc_21203_new_n2388_), .Y(w_mem_inst__abc_21203_new_n2389_));
INVX1 INVX1_1199 ( .A(w_mem_inst__abc_21203_new_n2391_), .Y(w_mem_inst__abc_21203_new_n2392_));
INVX1 INVX1_12 ( .A(_abc_15497_new_n740_), .Y(_abc_15497_new_n741_));
INVX1 INVX1_120 ( .A(_abc_15497_new_n1272_), .Y(_abc_15497_new_n1274_));
INVX1 INVX1_1200 ( .A(w_mem_inst__abc_21203_new_n2393_), .Y(w_mem_inst__abc_21203_new_n2395_));
INVX1 INVX1_1201 ( .A(w_mem_inst_w_mem_13__16_), .Y(w_mem_inst__abc_21203_new_n2432_));
INVX1 INVX1_1202 ( .A(w_mem_inst_w_mem_8__16_), .Y(w_mem_inst__abc_21203_new_n2434_));
INVX1 INVX1_1203 ( .A(w_mem_inst__abc_21203_new_n2436_), .Y(w_mem_inst__abc_21203_new_n2437_));
INVX1 INVX1_1204 ( .A(w_mem_inst__abc_21203_new_n2439_), .Y(w_mem_inst__abc_21203_new_n2440_));
INVX1 INVX1_1205 ( .A(w_mem_inst__abc_21203_new_n2441_), .Y(w_mem_inst__abc_21203_new_n2443_));
INVX1 INVX1_1206 ( .A(w_mem_inst_w_mem_13__17_), .Y(w_mem_inst__abc_21203_new_n2480_));
INVX1 INVX1_1207 ( .A(w_mem_inst_w_mem_8__17_), .Y(w_mem_inst__abc_21203_new_n2482_));
INVX1 INVX1_1208 ( .A(w_mem_inst__abc_21203_new_n2484_), .Y(w_mem_inst__abc_21203_new_n2485_));
INVX1 INVX1_1209 ( .A(w_mem_inst__abc_21203_new_n2487_), .Y(w_mem_inst__abc_21203_new_n2488_));
INVX1 INVX1_121 ( .A(_abc_15497_new_n1283_), .Y(_abc_15497_new_n1284_));
INVX1 INVX1_1210 ( .A(w_mem_inst__abc_21203_new_n2489_), .Y(w_mem_inst__abc_21203_new_n2491_));
INVX1 INVX1_1211 ( .A(w_mem_inst_w_mem_13__18_), .Y(w_mem_inst__abc_21203_new_n2528_));
INVX1 INVX1_1212 ( .A(w_mem_inst_w_mem_8__18_), .Y(w_mem_inst__abc_21203_new_n2530_));
INVX1 INVX1_1213 ( .A(w_mem_inst__abc_21203_new_n2532_), .Y(w_mem_inst__abc_21203_new_n2533_));
INVX1 INVX1_1214 ( .A(w_mem_inst__abc_21203_new_n2535_), .Y(w_mem_inst__abc_21203_new_n2536_));
INVX1 INVX1_1215 ( .A(w_mem_inst__abc_21203_new_n2537_), .Y(w_mem_inst__abc_21203_new_n2539_));
INVX1 INVX1_1216 ( .A(w_mem_inst_w_mem_13__19_), .Y(w_mem_inst__abc_21203_new_n2576_));
INVX1 INVX1_1217 ( .A(w_mem_inst_w_mem_8__19_), .Y(w_mem_inst__abc_21203_new_n2578_));
INVX1 INVX1_1218 ( .A(w_mem_inst__abc_21203_new_n2580_), .Y(w_mem_inst__abc_21203_new_n2581_));
INVX1 INVX1_1219 ( .A(w_mem_inst__abc_21203_new_n2583_), .Y(w_mem_inst__abc_21203_new_n2584_));
INVX1 INVX1_122 ( .A(_abc_15497_new_n1269_), .Y(_abc_15497_new_n1286_));
INVX1 INVX1_1220 ( .A(w_mem_inst__abc_21203_new_n2585_), .Y(w_mem_inst__abc_21203_new_n2587_));
INVX1 INVX1_1221 ( .A(w_mem_inst_w_mem_13__20_), .Y(w_mem_inst__abc_21203_new_n2624_));
INVX1 INVX1_1222 ( .A(w_mem_inst_w_mem_8__20_), .Y(w_mem_inst__abc_21203_new_n2626_));
INVX1 INVX1_1223 ( .A(w_mem_inst__abc_21203_new_n2628_), .Y(w_mem_inst__abc_21203_new_n2629_));
INVX1 INVX1_1224 ( .A(w_mem_inst__abc_21203_new_n2631_), .Y(w_mem_inst__abc_21203_new_n2632_));
INVX1 INVX1_1225 ( .A(w_mem_inst__abc_21203_new_n2633_), .Y(w_mem_inst__abc_21203_new_n2635_));
INVX1 INVX1_1226 ( .A(w_mem_inst_w_mem_13__21_), .Y(w_mem_inst__abc_21203_new_n2672_));
INVX1 INVX1_1227 ( .A(w_mem_inst_w_mem_8__21_), .Y(w_mem_inst__abc_21203_new_n2674_));
INVX1 INVX1_1228 ( .A(w_mem_inst__abc_21203_new_n2676_), .Y(w_mem_inst__abc_21203_new_n2677_));
INVX1 INVX1_1229 ( .A(w_mem_inst__abc_21203_new_n2679_), .Y(w_mem_inst__abc_21203_new_n2680_));
INVX1 INVX1_123 ( .A(_abc_15497_new_n1289_), .Y(_abc_15497_new_n1290_));
INVX1 INVX1_1230 ( .A(w_mem_inst__abc_21203_new_n2681_), .Y(w_mem_inst__abc_21203_new_n2683_));
INVX1 INVX1_1231 ( .A(w_mem_inst_w_mem_13__22_), .Y(w_mem_inst__abc_21203_new_n2720_));
INVX1 INVX1_1232 ( .A(w_mem_inst_w_mem_8__22_), .Y(w_mem_inst__abc_21203_new_n2722_));
INVX1 INVX1_1233 ( .A(w_mem_inst__abc_21203_new_n2724_), .Y(w_mem_inst__abc_21203_new_n2725_));
INVX1 INVX1_1234 ( .A(w_mem_inst__abc_21203_new_n2727_), .Y(w_mem_inst__abc_21203_new_n2728_));
INVX1 INVX1_1235 ( .A(w_mem_inst__abc_21203_new_n2729_), .Y(w_mem_inst__abc_21203_new_n2731_));
INVX1 INVX1_1236 ( .A(w_mem_inst_w_mem_13__23_), .Y(w_mem_inst__abc_21203_new_n2768_));
INVX1 INVX1_1237 ( .A(w_mem_inst_w_mem_8__23_), .Y(w_mem_inst__abc_21203_new_n2770_));
INVX1 INVX1_1238 ( .A(w_mem_inst__abc_21203_new_n2772_), .Y(w_mem_inst__abc_21203_new_n2773_));
INVX1 INVX1_1239 ( .A(w_mem_inst__abc_21203_new_n2775_), .Y(w_mem_inst__abc_21203_new_n2776_));
INVX1 INVX1_124 ( .A(_abc_15497_new_n1292_), .Y(_abc_15497_new_n1293_));
INVX1 INVX1_1240 ( .A(w_mem_inst__abc_21203_new_n2777_), .Y(w_mem_inst__abc_21203_new_n2779_));
INVX1 INVX1_1241 ( .A(w_mem_inst_w_mem_13__24_), .Y(w_mem_inst__abc_21203_new_n2816_));
INVX1 INVX1_1242 ( .A(w_mem_inst_w_mem_8__24_), .Y(w_mem_inst__abc_21203_new_n2818_));
INVX1 INVX1_1243 ( .A(w_mem_inst__abc_21203_new_n2820_), .Y(w_mem_inst__abc_21203_new_n2821_));
INVX1 INVX1_1244 ( .A(w_mem_inst__abc_21203_new_n2823_), .Y(w_mem_inst__abc_21203_new_n2824_));
INVX1 INVX1_1245 ( .A(w_mem_inst__abc_21203_new_n2825_), .Y(w_mem_inst__abc_21203_new_n2827_));
INVX1 INVX1_1246 ( .A(w_mem_inst_w_mem_13__25_), .Y(w_mem_inst__abc_21203_new_n2864_));
INVX1 INVX1_1247 ( .A(w_mem_inst_w_mem_8__25_), .Y(w_mem_inst__abc_21203_new_n2866_));
INVX1 INVX1_1248 ( .A(w_mem_inst__abc_21203_new_n2868_), .Y(w_mem_inst__abc_21203_new_n2869_));
INVX1 INVX1_1249 ( .A(w_mem_inst__abc_21203_new_n2871_), .Y(w_mem_inst__abc_21203_new_n2872_));
INVX1 INVX1_125 ( .A(_abc_15497_new_n1298_), .Y(_abc_15497_new_n1299_));
INVX1 INVX1_1250 ( .A(w_mem_inst__abc_21203_new_n2873_), .Y(w_mem_inst__abc_21203_new_n2875_));
INVX1 INVX1_1251 ( .A(w_mem_inst_w_mem_13__26_), .Y(w_mem_inst__abc_21203_new_n2912_));
INVX1 INVX1_1252 ( .A(w_mem_inst_w_mem_8__26_), .Y(w_mem_inst__abc_21203_new_n2914_));
INVX1 INVX1_1253 ( .A(w_mem_inst__abc_21203_new_n2916_), .Y(w_mem_inst__abc_21203_new_n2917_));
INVX1 INVX1_1254 ( .A(w_mem_inst__abc_21203_new_n2919_), .Y(w_mem_inst__abc_21203_new_n2920_));
INVX1 INVX1_1255 ( .A(w_mem_inst__abc_21203_new_n2921_), .Y(w_mem_inst__abc_21203_new_n2923_));
INVX1 INVX1_1256 ( .A(w_mem_inst_w_mem_13__27_), .Y(w_mem_inst__abc_21203_new_n2960_));
INVX1 INVX1_1257 ( .A(w_mem_inst_w_mem_8__27_), .Y(w_mem_inst__abc_21203_new_n2962_));
INVX1 INVX1_1258 ( .A(w_mem_inst__abc_21203_new_n2964_), .Y(w_mem_inst__abc_21203_new_n2965_));
INVX1 INVX1_1259 ( .A(w_mem_inst__abc_21203_new_n2967_), .Y(w_mem_inst__abc_21203_new_n2968_));
INVX1 INVX1_126 ( .A(_abc_15497_new_n1301_), .Y(_abc_15497_new_n1302_));
INVX1 INVX1_1260 ( .A(w_mem_inst__abc_21203_new_n2969_), .Y(w_mem_inst__abc_21203_new_n2971_));
INVX1 INVX1_1261 ( .A(w_mem_inst_w_mem_13__28_), .Y(w_mem_inst__abc_21203_new_n3008_));
INVX1 INVX1_1262 ( .A(w_mem_inst_w_mem_8__28_), .Y(w_mem_inst__abc_21203_new_n3010_));
INVX1 INVX1_1263 ( .A(w_mem_inst__abc_21203_new_n3012_), .Y(w_mem_inst__abc_21203_new_n3013_));
INVX1 INVX1_1264 ( .A(w_mem_inst__abc_21203_new_n3015_), .Y(w_mem_inst__abc_21203_new_n3016_));
INVX1 INVX1_1265 ( .A(w_mem_inst__abc_21203_new_n3017_), .Y(w_mem_inst__abc_21203_new_n3019_));
INVX1 INVX1_1266 ( .A(w_mem_inst_w_mem_13__29_), .Y(w_mem_inst__abc_21203_new_n3056_));
INVX1 INVX1_1267 ( .A(w_mem_inst_w_mem_8__29_), .Y(w_mem_inst__abc_21203_new_n3058_));
INVX1 INVX1_1268 ( .A(w_mem_inst__abc_21203_new_n3060_), .Y(w_mem_inst__abc_21203_new_n3061_));
INVX1 INVX1_1269 ( .A(w_mem_inst__abc_21203_new_n3063_), .Y(w_mem_inst__abc_21203_new_n3064_));
INVX1 INVX1_127 ( .A(_abc_15497_new_n1303_), .Y(_abc_15497_new_n1305_));
INVX1 INVX1_1270 ( .A(w_mem_inst__abc_21203_new_n3065_), .Y(w_mem_inst__abc_21203_new_n3067_));
INVX1 INVX1_1271 ( .A(w_mem_inst_w_mem_13__30_), .Y(w_mem_inst__abc_21203_new_n3104_));
INVX1 INVX1_1272 ( .A(w_mem_inst_w_mem_8__30_), .Y(w_mem_inst__abc_21203_new_n3106_));
INVX1 INVX1_1273 ( .A(w_mem_inst__abc_21203_new_n3108_), .Y(w_mem_inst__abc_21203_new_n3109_));
INVX1 INVX1_1274 ( .A(w_mem_inst__abc_21203_new_n3111_), .Y(w_mem_inst__abc_21203_new_n3112_));
INVX1 INVX1_1275 ( .A(w_mem_inst__abc_21203_new_n3113_), .Y(w_mem_inst__abc_21203_new_n3115_));
INVX1 INVX1_1276 ( .A(round_ctr_rst), .Y(w_mem_inst__abc_21203_new_n3152_));
INVX1 INVX1_1277 ( .A(w_mem_inst__abc_21203_new_n3153_), .Y(w_mem_inst__abc_21203_new_n3154_));
INVX1 INVX1_1278 ( .A(round_ctr_inc), .Y(w_mem_inst__abc_21203_new_n6229_));
INVX1 INVX1_1279 ( .A(w_mem_inst__abc_21203_new_n6242_), .Y(w_mem_inst__abc_21203_new_n6243_));
INVX1 INVX1_128 ( .A(_abc_15497_new_n1311_), .Y(_abc_15497_new_n1312_));
INVX1 INVX1_1280 ( .A(w_mem_inst__abc_21203_new_n6247_), .Y(w_mem_inst__abc_21203_new_n6248_));
INVX1 INVX1_1281 ( .A(w_mem_inst__abc_21203_new_n6252_), .Y(w_mem_inst__abc_21203_new_n6253_));
INVX1 INVX1_1282 ( .A(w_mem_inst__abc_21203_new_n6257_), .Y(w_mem_inst__abc_21203_new_n6258_));
INVX1 INVX1_1283 ( .A(w_mem_inst__abc_21203_new_n6262_), .Y(w_mem_inst__abc_21203_new_n6263_));
INVX1 INVX1_129 ( .A(_abc_15497_new_n1314_), .Y(_abc_15497_new_n1315_));
INVX1 INVX1_13 ( .A(_abc_15497_new_n743_), .Y(_abc_15497_new_n744_));
INVX1 INVX1_130 ( .A(_abc_15497_new_n1317_), .Y(_abc_15497_new_n1318_));
INVX1 INVX1_131 ( .A(_abc_15497_new_n1324_), .Y(_abc_15497_new_n1325_));
INVX1 INVX1_132 ( .A(_abc_15497_new_n1328_), .Y(_abc_15497_new_n1329_));
INVX1 INVX1_133 ( .A(_abc_15497_new_n1337_), .Y(_abc_15497_new_n1338_));
INVX1 INVX1_134 ( .A(_abc_15497_new_n1343_), .Y(_abc_15497_new_n1344_));
INVX1 INVX1_135 ( .A(_abc_15497_new_n1345_), .Y(_abc_15497_new_n1346_));
INVX1 INVX1_136 ( .A(_abc_15497_new_n1352_), .Y(_abc_15497_new_n1353_));
INVX1 INVX1_137 ( .A(_abc_15497_new_n1355_), .Y(_abc_15497_new_n1356_));
INVX1 INVX1_138 ( .A(_abc_15497_new_n1359_), .Y(_abc_15497_new_n1360_));
INVX1 INVX1_139 ( .A(_abc_15497_new_n1368_), .Y(_abc_15497_new_n1369_));
INVX1 INVX1_14 ( .A(_abc_15497_new_n745_), .Y(_abc_15497_new_n746_));
INVX1 INVX1_140 ( .A(_abc_15497_new_n1366_), .Y(_abc_15497_new_n1372_));
INVX1 INVX1_141 ( .A(_abc_15497_new_n1370_), .Y(_abc_15497_new_n1373_));
INVX1 INVX1_142 ( .A(_abc_15497_new_n1351_), .Y(_abc_15497_new_n1385_));
INVX1 INVX1_143 ( .A(_abc_15497_new_n1393_), .Y(_abc_15497_new_n1394_));
INVX1 INVX1_144 ( .A(_abc_15497_new_n1397_), .Y(_abc_15497_new_n1398_));
INVX1 INVX1_145 ( .A(_abc_15497_new_n1404_), .Y(_abc_15497_new_n1405_));
INVX1 INVX1_146 ( .A(_abc_15497_new_n1407_), .Y(_abc_15497_new_n1408_));
INVX1 INVX1_147 ( .A(_abc_15497_new_n1409_), .Y(_abc_15497_new_n1411_));
INVX1 INVX1_148 ( .A(_abc_15497_new_n1425_), .Y(_abc_15497_new_n1426_));
INVX1 INVX1_149 ( .A(_abc_15497_new_n1429_), .Y(_abc_15497_new_n1430_));
INVX1 INVX1_15 ( .A(_abc_15497_new_n748_), .Y(_abc_15497_new_n749_));
INVX1 INVX1_150 ( .A(_abc_15497_new_n1436_), .Y(_abc_15497_new_n1437_));
INVX1 INVX1_151 ( .A(_abc_15497_new_n1388_), .Y(_abc_15497_new_n1441_));
INVX1 INVX1_152 ( .A(_abc_15497_new_n1253_), .Y(_abc_15497_new_n1442_));
INVX1 INVX1_153 ( .A(_abc_15497_new_n1106_), .Y(_abc_15497_new_n1443_));
INVX1 INVX1_154 ( .A(_abc_15497_new_n1254_), .Y(_abc_15497_new_n1446_));
INVX1 INVX1_155 ( .A(_abc_15497_new_n1389_), .Y(_abc_15497_new_n1449_));
INVX1 INVX1_156 ( .A(_abc_15497_new_n1419_), .Y(_abc_15497_new_n1452_));
INVX1 INVX1_157 ( .A(_abc_15497_new_n1422_), .Y(_abc_15497_new_n1454_));
INVX1 INVX1_158 ( .A(_abc_15497_new_n1456_), .Y(_abc_15497_new_n1457_));
INVX1 INVX1_159 ( .A(_abc_15497_new_n1459_), .Y(_abc_15497_new_n1460_));
INVX1 INVX1_16 ( .A(_abc_15497_new_n754_), .Y(_abc_15497_new_n755_));
INVX1 INVX1_160 ( .A(_abc_15497_new_n1467_), .Y(_abc_15497_new_n1468_));
INVX1 INVX1_161 ( .A(_abc_15497_new_n1471_), .Y(_abc_15497_new_n1472_));
INVX1 INVX1_162 ( .A(_abc_15497_new_n1473_), .Y(_abc_15497_new_n1476_));
INVX1 INVX1_163 ( .A(_abc_15497_new_n1485_), .Y(_abc_15497_new_n1486_));
INVX1 INVX1_164 ( .A(_abc_15497_new_n1487_), .Y(_abc_15497_new_n1491_));
INVX1 INVX1_165 ( .A(_abc_15497_new_n1497_), .Y(_abc_15497_new_n1498_));
INVX1 INVX1_166 ( .A(_abc_15497_new_n1499_), .Y(_abc_15497_new_n1503_));
INVX1 INVX1_167 ( .A(_abc_15497_new_n1484_), .Y(_abc_15497_new_n1504_));
INVX1 INVX1_168 ( .A(e_reg_31_), .Y(_abc_15497_new_n1515_));
INVX1 INVX1_169 ( .A(\digest[31] ), .Y(_abc_15497_new_n1517_));
INVX1 INVX1_17 ( .A(_abc_15497_new_n756_), .Y(_abc_15497_new_n757_));
INVX1 INVX1_170 ( .A(_abc_15497_new_n1519_), .Y(_abc_15497_new_n1520_));
INVX1 INVX1_171 ( .A(_abc_15497_new_n1529_), .Y(_abc_15497_new_n1530_));
INVX1 INVX1_172 ( .A(_abc_15497_new_n1537_), .Y(_abc_15497_new_n1538_));
INVX1 INVX1_173 ( .A(_abc_15497_new_n1540_), .Y(_abc_15497_new_n1541_));
INVX1 INVX1_174 ( .A(_abc_15497_new_n1550_), .Y(_abc_15497_new_n1551_));
INVX1 INVX1_175 ( .A(_abc_15497_new_n1553_), .Y(_abc_15497_new_n1554_));
INVX1 INVX1_176 ( .A(_abc_15497_new_n1564_), .Y(_abc_15497_new_n1565_));
INVX1 INVX1_177 ( .A(_abc_15497_new_n1562_), .Y(_abc_15497_new_n1568_));
INVX1 INVX1_178 ( .A(_abc_15497_new_n1566_), .Y(_abc_15497_new_n1569_));
INVX1 INVX1_179 ( .A(_abc_15497_new_n1575_), .Y(_abc_15497_new_n1576_));
INVX1 INVX1_18 ( .A(_abc_15497_new_n758_), .Y(_abc_15497_new_n759_));
INVX1 INVX1_180 ( .A(_abc_15497_new_n1580_), .Y(_abc_15497_new_n1581_));
INVX1 INVX1_181 ( .A(_abc_15497_new_n1590_), .Y(_abc_15497_new_n1591_));
INVX1 INVX1_182 ( .A(_abc_15497_new_n1594_), .Y(_abc_15497_new_n1595_));
INVX1 INVX1_183 ( .A(_abc_15497_new_n1603_), .Y(_abc_15497_new_n1604_));
INVX1 INVX1_184 ( .A(_abc_15497_new_n1607_), .Y(_abc_15497_new_n1608_));
INVX1 INVX1_185 ( .A(_abc_15497_new_n1616_), .Y(_abc_15497_new_n1617_));
INVX1 INVX1_186 ( .A(_abc_15497_new_n1621_), .Y(_abc_15497_new_n1622_));
INVX1 INVX1_187 ( .A(_abc_15497_new_n1629_), .Y(_abc_15497_new_n1630_));
INVX1 INVX1_188 ( .A(_abc_15497_new_n1633_), .Y(_abc_15497_new_n1634_));
INVX1 INVX1_189 ( .A(_abc_15497_new_n1640_), .Y(_abc_15497_new_n1641_));
INVX1 INVX1_19 ( .A(_abc_15497_new_n762_), .Y(_abc_15497_new_n763_));
INVX1 INVX1_190 ( .A(_abc_15497_new_n1646_), .Y(_abc_15497_new_n1647_));
INVX1 INVX1_191 ( .A(_abc_15497_new_n1648_), .Y(_abc_15497_new_n1649_));
INVX1 INVX1_192 ( .A(_abc_15497_new_n1655_), .Y(_abc_15497_new_n1656_));
INVX1 INVX1_193 ( .A(_abc_15497_new_n1658_), .Y(_abc_15497_new_n1659_));
INVX1 INVX1_194 ( .A(_abc_15497_new_n1662_), .Y(_abc_15497_new_n1663_));
INVX1 INVX1_195 ( .A(_abc_15497_new_n1670_), .Y(_abc_15497_new_n1671_));
INVX1 INVX1_196 ( .A(_abc_15497_new_n1673_), .Y(_abc_15497_new_n1674_));
INVX1 INVX1_197 ( .A(_abc_15497_new_n1675_), .Y(_abc_15497_new_n1677_));
INVX1 INVX1_198 ( .A(_abc_15497_new_n1654_), .Y(_abc_15497_new_n1685_));
INVX1 INVX1_199 ( .A(_abc_15497_new_n1692_), .Y(_abc_15497_new_n1693_));
INVX1 INVX1_2 ( .A(_abc_15497_new_n699_), .Y(_abc_15497_new_n700_));
INVX1 INVX1_20 ( .A(_abc_15497_new_n767_), .Y(_abc_15497_new_n768_));
INVX1 INVX1_200 ( .A(_abc_15497_new_n1696_), .Y(_abc_15497_new_n1697_));
INVX1 INVX1_201 ( .A(_abc_15497_new_n1705_), .Y(_abc_15497_new_n1706_));
INVX1 INVX1_202 ( .A(_abc_15497_new_n1711_), .Y(_abc_15497_new_n1712_));
INVX1 INVX1_203 ( .A(_abc_15497_new_n1713_), .Y(_abc_15497_new_n1714_));
INVX1 INVX1_204 ( .A(_abc_15497_new_n1720_), .Y(_abc_15497_new_n1721_));
INVX1 INVX1_205 ( .A(_abc_15497_new_n1723_), .Y(_abc_15497_new_n1724_));
INVX1 INVX1_206 ( .A(_abc_15497_new_n1727_), .Y(_abc_15497_new_n1728_));
INVX1 INVX1_207 ( .A(_abc_15497_new_n1735_), .Y(_abc_15497_new_n1736_));
INVX1 INVX1_208 ( .A(_abc_15497_new_n1738_), .Y(_abc_15497_new_n1739_));
INVX1 INVX1_209 ( .A(_abc_15497_new_n1740_), .Y(_abc_15497_new_n1742_));
INVX1 INVX1_21 ( .A(_abc_15497_new_n769_), .Y(_abc_15497_new_n770_));
INVX1 INVX1_210 ( .A(_abc_15497_new_n1748_), .Y(_abc_15497_new_n1749_));
INVX1 INVX1_211 ( .A(_abc_15497_new_n1752_), .Y(_abc_15497_new_n1753_));
INVX1 INVX1_212 ( .A(_abc_15497_new_n1754_), .Y(_abc_15497_new_n1755_));
INVX1 INVX1_213 ( .A(_abc_15497_new_n1760_), .Y(_abc_15497_new_n1761_));
INVX1 INVX1_214 ( .A(_abc_15497_new_n1764_), .Y(_abc_15497_new_n1765_));
INVX1 INVX1_215 ( .A(_abc_15497_new_n1771_), .Y(_abc_15497_new_n1772_));
INVX1 INVX1_216 ( .A(_abc_15497_new_n1769_), .Y(_abc_15497_new_n1775_));
INVX1 INVX1_217 ( .A(_abc_15497_new_n1773_), .Y(_abc_15497_new_n1776_));
INVX1 INVX1_218 ( .A(_abc_15497_new_n1790_), .Y(_abc_15497_new_n1791_));
INVX1 INVX1_219 ( .A(_abc_15497_new_n1794_), .Y(_abc_15497_new_n1795_));
INVX1 INVX1_22 ( .A(_abc_15497_new_n772_), .Y(_abc_15497_new_n773_));
INVX1 INVX1_220 ( .A(_abc_15497_new_n1800_), .Y(_abc_15497_new_n1801_));
INVX1 INVX1_221 ( .A(_abc_15497_new_n1803_), .Y(_abc_15497_new_n1804_));
INVX1 INVX1_222 ( .A(_abc_15497_new_n1805_), .Y(_abc_15497_new_n1807_));
INVX1 INVX1_223 ( .A(_abc_15497_new_n1821_), .Y(_abc_15497_new_n1822_));
INVX1 INVX1_224 ( .A(_abc_15497_new_n1825_), .Y(_abc_15497_new_n1826_));
INVX1 INVX1_225 ( .A(_abc_15497_new_n1832_), .Y(_abc_15497_new_n1833_));
INVX1 INVX1_226 ( .A(_abc_15497_new_n1835_), .Y(_abc_15497_new_n1836_));
INVX1 INVX1_227 ( .A(_abc_15497_new_n1837_), .Y(_abc_15497_new_n1839_));
INVX1 INVX1_228 ( .A(_abc_15497_new_n1848_), .Y(_abc_15497_new_n1849_));
INVX1 INVX1_229 ( .A(_abc_15497_new_n1834_), .Y(_abc_15497_new_n1851_));
INVX1 INVX1_23 ( .A(_abc_15497_new_n775_), .Y(_abc_15497_new_n776_));
INVX1 INVX1_230 ( .A(_abc_15497_new_n1854_), .Y(_abc_15497_new_n1855_));
INVX1 INVX1_231 ( .A(_abc_15497_new_n1857_), .Y(_abc_15497_new_n1858_));
INVX1 INVX1_232 ( .A(_abc_15497_new_n1865_), .Y(_abc_15497_new_n1866_));
INVX1 INVX1_233 ( .A(_abc_15497_new_n1863_), .Y(_abc_15497_new_n1869_));
INVX1 INVX1_234 ( .A(_abc_15497_new_n1867_), .Y(_abc_15497_new_n1870_));
INVX1 INVX1_235 ( .A(_abc_15497_new_n1877_), .Y(_abc_15497_new_n1878_));
INVX1 INVX1_236 ( .A(_abc_15497_new_n1880_), .Y(_abc_15497_new_n1881_));
INVX1 INVX1_237 ( .A(_abc_15497_new_n1883_), .Y(_abc_15497_new_n1884_));
INVX1 INVX1_238 ( .A(_abc_15497_new_n1890_), .Y(_abc_15497_new_n1891_));
INVX1 INVX1_239 ( .A(_abc_15497_new_n1894_), .Y(_abc_15497_new_n1895_));
INVX1 INVX1_24 ( .A(_abc_15497_new_n785_), .Y(_abc_15497_new_n790_));
INVX1 INVX1_240 ( .A(_abc_15497_new_n1901_), .Y(_abc_15497_new_n1902_));
INVX1 INVX1_241 ( .A(_abc_15497_new_n1907_), .Y(_abc_15497_new_n1908_));
INVX1 INVX1_242 ( .A(_abc_15497_new_n1909_), .Y(_abc_15497_new_n1910_));
INVX1 INVX1_243 ( .A(_abc_15497_new_n1917_), .Y(_abc_15497_new_n1918_));
INVX1 INVX1_244 ( .A(_abc_15497_new_n1920_), .Y(_abc_15497_new_n1921_));
INVX1 INVX1_245 ( .A(_abc_15497_new_n1924_), .Y(_abc_15497_new_n1925_));
INVX1 INVX1_246 ( .A(_abc_15497_new_n1931_), .Y(_abc_15497_new_n1932_));
INVX1 INVX1_247 ( .A(_abc_15497_new_n1936_), .Y(_abc_15497_new_n1937_));
INVX1 INVX1_248 ( .A(_abc_15497_new_n1939_), .Y(_abc_15497_new_n1940_));
INVX1 INVX1_249 ( .A(_abc_15497_new_n1949_), .Y(_abc_15497_new_n1950_));
INVX1 INVX1_25 ( .A(_abc_15497_new_n787_), .Y(_abc_15497_new_n792_));
INVX1 INVX1_250 ( .A(_abc_15497_new_n1953_), .Y(_abc_15497_new_n1954_));
INVX1 INVX1_251 ( .A(_abc_15497_new_n1957_), .Y(_abc_15497_new_n1958_));
INVX1 INVX1_252 ( .A(_abc_15497_new_n1965_), .Y(_abc_15497_new_n1966_));
INVX1 INVX1_253 ( .A(_abc_15497_new_n1968_), .Y(_abc_15497_new_n1969_));
INVX1 INVX1_254 ( .A(_abc_15497_new_n1970_), .Y(_abc_15497_new_n1972_));
INVX1 INVX1_255 ( .A(_abc_15497_new_n1978_), .Y(_abc_15497_new_n1979_));
INVX1 INVX1_256 ( .A(_abc_15497_new_n1987_), .Y(_abc_15497_new_n1988_));
INVX1 INVX1_257 ( .A(_abc_15497_new_n1994_), .Y(_abc_15497_new_n1995_));
INVX1 INVX1_258 ( .A(_abc_15497_new_n1997_), .Y(_abc_15497_new_n1998_));
INVX1 INVX1_259 ( .A(_abc_15497_new_n1999_), .Y(_abc_15497_new_n2000_));
INVX1 INVX1_26 ( .A(_abc_15497_new_n801_), .Y(_abc_15497_new_n806_));
INVX1 INVX1_260 ( .A(round_ctr_inc), .Y(_abc_15497_new_n2008_));
INVX1 INVX1_261 ( .A(round_ctr_rst), .Y(_abc_15497_new_n2009_));
INVX1 INVX1_262 ( .A(_abc_15497_new_n2188_), .Y(_abc_15497_new_n2189_));
INVX1 INVX1_263 ( .A(_abc_15497_new_n2195_), .Y(_abc_15497_new_n2196_));
INVX1 INVX1_264 ( .A(_abc_15497_new_n2197_), .Y(_abc_15497_new_n2200_));
INVX1 INVX1_265 ( .A(_abc_15497_new_n2209_), .Y(_abc_15497_new_n2210_));
INVX1 INVX1_266 ( .A(_abc_15497_new_n2211_), .Y(_abc_15497_new_n2212_));
INVX1 INVX1_267 ( .A(_abc_15497_new_n2224_), .Y(_abc_15497_new_n2225_));
INVX1 INVX1_268 ( .A(_abc_15497_new_n2226_), .Y(_abc_15497_new_n2229_));
INVX1 INVX1_269 ( .A(_abc_15497_new_n2237_), .Y(_abc_15497_new_n2238_));
INVX1 INVX1_27 ( .A(_abc_15497_new_n803_), .Y(_abc_15497_new_n808_));
INVX1 INVX1_270 ( .A(_abc_15497_new_n2239_), .Y(_abc_15497_new_n2240_));
INVX1 INVX1_271 ( .A(_abc_15497_new_n2223_), .Y(_abc_15497_new_n2241_));
INVX1 INVX1_272 ( .A(_abc_15497_new_n2256_), .Y(_abc_15497_new_n2257_));
INVX1 INVX1_273 ( .A(_abc_15497_new_n2258_), .Y(_abc_15497_new_n2261_));
INVX1 INVX1_274 ( .A(_abc_15497_new_n2270_), .Y(_abc_15497_new_n2271_));
INVX1 INVX1_275 ( .A(_abc_15497_new_n2272_), .Y(_abc_15497_new_n2275_));
INVX1 INVX1_276 ( .A(_abc_15497_new_n2284_), .Y(_abc_15497_new_n2285_));
INVX1 INVX1_277 ( .A(_abc_15497_new_n2286_), .Y(_abc_15497_new_n2290_));
INVX1 INVX1_278 ( .A(_abc_15497_new_n2296_), .Y(_abc_15497_new_n2297_));
INVX1 INVX1_279 ( .A(_abc_15497_new_n2302_), .Y(_abc_15497_new_n2303_));
INVX1 INVX1_28 ( .A(_abc_15497_new_n818_), .Y(_abc_15497_new_n820_));
INVX1 INVX1_280 ( .A(_abc_15497_new_n2309_), .Y(_abc_15497_new_n2310_));
INVX1 INVX1_281 ( .A(_abc_15497_new_n2312_), .Y(_abc_15497_new_n2313_));
INVX1 INVX1_282 ( .A(_abc_15497_new_n2314_), .Y(_abc_15497_new_n2316_));
INVX1 INVX1_283 ( .A(_abc_15497_new_n2327_), .Y(_abc_15497_new_n2328_));
INVX1 INVX1_284 ( .A(_abc_15497_new_n2331_), .Y(_abc_15497_new_n2332_));
INVX1 INVX1_285 ( .A(_abc_15497_new_n2335_), .Y(_abc_15497_new_n2336_));
INVX1 INVX1_286 ( .A(_abc_15497_new_n2342_), .Y(_abc_15497_new_n2343_));
INVX1 INVX1_287 ( .A(_abc_15497_new_n2340_), .Y(_abc_15497_new_n2346_));
INVX1 INVX1_288 ( .A(_abc_15497_new_n2344_), .Y(_abc_15497_new_n2347_));
INVX1 INVX1_289 ( .A(_abc_15497_new_n2356_), .Y(_abc_15497_new_n2357_));
INVX1 INVX1_29 ( .A(_abc_15497_new_n817_), .Y(_abc_15497_new_n825_));
INVX1 INVX1_290 ( .A(_abc_15497_new_n2368_), .Y(_abc_15497_new_n2369_));
INVX1 INVX1_291 ( .A(_abc_15497_new_n2373_), .Y(_abc_15497_new_n2374_));
INVX1 INVX1_292 ( .A(_abc_15497_new_n2376_), .Y(_abc_15497_new_n2377_));
INVX1 INVX1_293 ( .A(_abc_15497_new_n2378_), .Y(_abc_15497_new_n2380_));
INVX1 INVX1_294 ( .A(_abc_15497_new_n2389_), .Y(_abc_15497_new_n2390_));
INVX1 INVX1_295 ( .A(_abc_15497_new_n2375_), .Y(_abc_15497_new_n2392_));
INVX1 INVX1_296 ( .A(_abc_15497_new_n2395_), .Y(_abc_15497_new_n2396_));
INVX1 INVX1_297 ( .A(_abc_15497_new_n2398_), .Y(_abc_15497_new_n2399_));
INVX1 INVX1_298 ( .A(_abc_15497_new_n2403_), .Y(_abc_15497_new_n2404_));
INVX1 INVX1_299 ( .A(_abc_15497_new_n2406_), .Y(_abc_15497_new_n2407_));
INVX1 INVX1_3 ( .A(_abc_15497_new_n704_), .Y(_abc_15497_new_n705_));
INVX1 INVX1_30 ( .A(_abc_15497_new_n814_), .Y(_abc_15497_new_n832_));
INVX1 INVX1_300 ( .A(_abc_15497_new_n2408_), .Y(_abc_15497_new_n2410_));
INVX1 INVX1_301 ( .A(_abc_15497_new_n2418_), .Y(_abc_15497_new_n2419_));
INVX1 INVX1_302 ( .A(_abc_15497_new_n2421_), .Y(_abc_15497_new_n2422_));
INVX1 INVX1_303 ( .A(_abc_15497_new_n2424_), .Y(_abc_15497_new_n2425_));
INVX1 INVX1_304 ( .A(_abc_15497_new_n2431_), .Y(_abc_15497_new_n2432_));
INVX1 INVX1_305 ( .A(_abc_15497_new_n2435_), .Y(_abc_15497_new_n2436_));
INVX1 INVX1_306 ( .A(_abc_15497_new_n2444_), .Y(_abc_15497_new_n2445_));
INVX1 INVX1_307 ( .A(_abc_15497_new_n2450_), .Y(_abc_15497_new_n2451_));
INVX1 INVX1_308 ( .A(_abc_15497_new_n2452_), .Y(_abc_15497_new_n2453_));
INVX1 INVX1_309 ( .A(_abc_15497_new_n2459_), .Y(_abc_15497_new_n2460_));
INVX1 INVX1_31 ( .A(_abc_15497_new_n796_), .Y(_abc_15497_new_n841_));
INVX1 INVX1_310 ( .A(_abc_15497_new_n2462_), .Y(_abc_15497_new_n2463_));
INVX1 INVX1_311 ( .A(_abc_15497_new_n2466_), .Y(_abc_15497_new_n2467_));
INVX1 INVX1_312 ( .A(_abc_15497_new_n2475_), .Y(_abc_15497_new_n2476_));
INVX1 INVX1_313 ( .A(_abc_15497_new_n2473_), .Y(_abc_15497_new_n2479_));
INVX1 INVX1_314 ( .A(_abc_15497_new_n2477_), .Y(_abc_15497_new_n2480_));
INVX1 INVX1_315 ( .A(_abc_15497_new_n2488_), .Y(_abc_15497_new_n2489_));
INVX1 INVX1_316 ( .A(_abc_15497_new_n2492_), .Y(_abc_15497_new_n2493_));
INVX1 INVX1_317 ( .A(_abc_15497_new_n2494_), .Y(_abc_15497_new_n2495_));
INVX1 INVX1_318 ( .A(_abc_15497_new_n2500_), .Y(_abc_15497_new_n2501_));
INVX1 INVX1_319 ( .A(_abc_15497_new_n2504_), .Y(_abc_15497_new_n2505_));
INVX1 INVX1_32 ( .A(_abc_15497_new_n798_), .Y(_abc_15497_new_n843_));
INVX1 INVX1_320 ( .A(_abc_15497_new_n2511_), .Y(_abc_15497_new_n2512_));
INVX1 INVX1_321 ( .A(_abc_15497_new_n2519_), .Y(_abc_15497_new_n2520_));
INVX1 INVX1_322 ( .A(_abc_15497_new_n2524_), .Y(_abc_15497_new_n2525_));
INVX1 INVX1_323 ( .A(_abc_15497_new_n2527_), .Y(_abc_15497_new_n2528_));
INVX1 INVX1_324 ( .A(_abc_15497_new_n2531_), .Y(_abc_15497_new_n2532_));
INVX1 INVX1_325 ( .A(_abc_15497_new_n2538_), .Y(_abc_15497_new_n2539_));
INVX1 INVX1_326 ( .A(_abc_15497_new_n2541_), .Y(_abc_15497_new_n2542_));
INVX1 INVX1_327 ( .A(_abc_15497_new_n2543_), .Y(_abc_15497_new_n2545_));
INVX1 INVX1_328 ( .A(_abc_15497_new_n2565_), .Y(_abc_15497_new_n2566_));
INVX1 INVX1_329 ( .A(_abc_15497_new_n2569_), .Y(_abc_15497_new_n2570_));
INVX1 INVX1_33 ( .A(_abc_15497_new_n860_), .Y(_abc_15497_new_n861_));
INVX1 INVX1_330 ( .A(_abc_15497_new_n2576_), .Y(_abc_15497_new_n2577_));
INVX1 INVX1_331 ( .A(_abc_15497_new_n2579_), .Y(_abc_15497_new_n2580_));
INVX1 INVX1_332 ( .A(_abc_15497_new_n2581_), .Y(_abc_15497_new_n2583_));
INVX1 INVX1_333 ( .A(_abc_15497_new_n2596_), .Y(_abc_15497_new_n2597_));
INVX1 INVX1_334 ( .A(_abc_15497_new_n2600_), .Y(_abc_15497_new_n2601_));
INVX1 INVX1_335 ( .A(_abc_15497_new_n2607_), .Y(_abc_15497_new_n2608_));
INVX1 INVX1_336 ( .A(_abc_15497_new_n2610_), .Y(_abc_15497_new_n2611_));
INVX1 INVX1_337 ( .A(_abc_15497_new_n2612_), .Y(_abc_15497_new_n2614_));
INVX1 INVX1_338 ( .A(_abc_15497_new_n2628_), .Y(_abc_15497_new_n2629_));
INVX1 INVX1_339 ( .A(_abc_15497_new_n2632_), .Y(_abc_15497_new_n2633_));
INVX1 INVX1_34 ( .A(_abc_15497_new_n864_), .Y(_abc_15497_new_n865_));
INVX1 INVX1_340 ( .A(_abc_15497_new_n2639_), .Y(_abc_15497_new_n2640_));
INVX1 INVX1_341 ( .A(_abc_15497_new_n2642_), .Y(_abc_15497_new_n2643_));
INVX1 INVX1_342 ( .A(_abc_15497_new_n2644_), .Y(_abc_15497_new_n2646_));
INVX1 INVX1_343 ( .A(_abc_15497_new_n2652_), .Y(_abc_15497_new_n2653_));
INVX1 INVX1_344 ( .A(_abc_15497_new_n2654_), .Y(_abc_15497_new_n2661_));
INVX1 INVX1_345 ( .A(_abc_15497_new_n2656_), .Y(_abc_15497_new_n2662_));
INVX1 INVX1_346 ( .A(_abc_15497_new_n2623_), .Y(_abc_15497_new_n2663_));
INVX1 INVX1_347 ( .A(_abc_15497_new_n2560_), .Y(_abc_15497_new_n2664_));
INVX1 INVX1_348 ( .A(_abc_15497_new_n2363_), .Y(_abc_15497_new_n2665_));
INVX1 INVX1_349 ( .A(_abc_15497_new_n2283_), .Y(_abc_15497_new_n2666_));
INVX1 INVX1_35 ( .A(_abc_15497_new_n874_), .Y(_abc_15497_new_n875_));
INVX1 INVX1_350 ( .A(_abc_15497_new_n2364_), .Y(_abc_15497_new_n2669_));
INVX1 INVX1_351 ( .A(_abc_15497_new_n2427_), .Y(_abc_15497_new_n2672_));
INVX1 INVX1_352 ( .A(_abc_15497_new_n2561_), .Y(_abc_15497_new_n2675_));
INVX1 INVX1_353 ( .A(_abc_15497_new_n2590_), .Y(_abc_15497_new_n2678_));
INVX1 INVX1_354 ( .A(_abc_15497_new_n2593_), .Y(_abc_15497_new_n2680_));
INVX1 INVX1_355 ( .A(_abc_15497_new_n2624_), .Y(_abc_15497_new_n2682_));
INVX1 INVX1_356 ( .A(_abc_15497_new_n2657_), .Y(_abc_15497_new_n2685_));
INVX1 INVX1_357 ( .A(\digest[127] ), .Y(_abc_15497_new_n2696_));
INVX1 INVX1_358 ( .A(b_reg_31_), .Y(_abc_15497_new_n2698_));
INVX1 INVX1_359 ( .A(_abc_15497_new_n2700_), .Y(_abc_15497_new_n2701_));
INVX1 INVX1_36 ( .A(_abc_15497_new_n878_), .Y(_abc_15497_new_n879_));
INVX1 INVX1_360 ( .A(_abc_15497_new_n2711_), .Y(_abc_15497_new_n2712_));
INVX1 INVX1_361 ( .A(_abc_15497_new_n2719_), .Y(_abc_15497_new_n2720_));
INVX1 INVX1_362 ( .A(_abc_15497_new_n2722_), .Y(_abc_15497_new_n2723_));
INVX1 INVX1_363 ( .A(_abc_15497_new_n2729_), .Y(_abc_15497_new_n2730_));
INVX1 INVX1_364 ( .A(_abc_15497_new_n2732_), .Y(_abc_15497_new_n2733_));
INVX1 INVX1_365 ( .A(_abc_15497_new_n2734_), .Y(_abc_15497_new_n2736_));
INVX1 INVX1_366 ( .A(_abc_15497_new_n2743_), .Y(_abc_15497_new_n2744_));
INVX1 INVX1_367 ( .A(_abc_15497_new_n2746_), .Y(_abc_15497_new_n2747_));
INVX1 INVX1_368 ( .A(_abc_15497_new_n2748_), .Y(_abc_15497_new_n2750_));
INVX1 INVX1_369 ( .A(_abc_15497_new_n2756_), .Y(_abc_15497_new_n2757_));
INVX1 INVX1_37 ( .A(_abc_15497_new_n883_), .Y(_abc_15497_new_n884_));
INVX1 INVX1_370 ( .A(_abc_15497_new_n2745_), .Y(_abc_15497_new_n2759_));
INVX1 INVX1_371 ( .A(_abc_15497_new_n2761_), .Y(_abc_15497_new_n2762_));
INVX1 INVX1_372 ( .A(_abc_15497_new_n2758_), .Y(_abc_15497_new_n2764_));
INVX1 INVX1_373 ( .A(_abc_15497_new_n2771_), .Y(_abc_15497_new_n2772_));
INVX1 INVX1_374 ( .A(_abc_15497_new_n2774_), .Y(_abc_15497_new_n2775_));
INVX1 INVX1_375 ( .A(_abc_15497_new_n2776_), .Y(_abc_15497_new_n2778_));
INVX1 INVX1_376 ( .A(_abc_15497_new_n2784_), .Y(_abc_15497_new_n2785_));
INVX1 INVX1_377 ( .A(_abc_15497_new_n2787_), .Y(_abc_15497_new_n2788_));
INVX1 INVX1_378 ( .A(_abc_15497_new_n2789_), .Y(_abc_15497_new_n2791_));
INVX1 INVX1_379 ( .A(_abc_15497_new_n2792_), .Y(_abc_15497_new_n2797_));
INVX1 INVX1_38 ( .A(_abc_15497_new_n886_), .Y(_abc_15497_new_n887_));
INVX1 INVX1_380 ( .A(_abc_15497_new_n2799_), .Y(_abc_15497_new_n2800_));
INVX1 INVX1_381 ( .A(_abc_15497_new_n2801_), .Y(_abc_15497_new_n2804_));
INVX1 INVX1_382 ( .A(_abc_15497_new_n2806_), .Y(_abc_15497_new_n2807_));
INVX1 INVX1_383 ( .A(_abc_15497_new_n2805_), .Y(_abc_15497_new_n2812_));
INVX1 INVX1_384 ( .A(_abc_15497_new_n2816_), .Y(_abc_15497_new_n2817_));
INVX1 INVX1_385 ( .A(_abc_15497_new_n2820_), .Y(_abc_15497_new_n2821_));
INVX1 INVX1_386 ( .A(_abc_15497_new_n2827_), .Y(_abc_15497_new_n2828_));
INVX1 INVX1_387 ( .A(_abc_15497_new_n2830_), .Y(_abc_15497_new_n2831_));
INVX1 INVX1_388 ( .A(_abc_15497_new_n2832_), .Y(_abc_15497_new_n2834_));
INVX1 INVX1_389 ( .A(_abc_15497_new_n2843_), .Y(_abc_15497_new_n2844_));
INVX1 INVX1_39 ( .A(_abc_15497_new_n888_), .Y(_abc_15497_new_n890_));
INVX1 INVX1_390 ( .A(_abc_15497_new_n2847_), .Y(_abc_15497_new_n2848_));
INVX1 INVX1_391 ( .A(_abc_15497_new_n2853_), .Y(_abc_15497_new_n2854_));
INVX1 INVX1_392 ( .A(_abc_15497_new_n2859_), .Y(_abc_15497_new_n2860_));
INVX1 INVX1_393 ( .A(_abc_15497_new_n2862_), .Y(_abc_15497_new_n2863_));
INVX1 INVX1_394 ( .A(_abc_15497_new_n2864_), .Y(_abc_15497_new_n2866_));
INVX1 INVX1_395 ( .A(_abc_15497_new_n2875_), .Y(_abc_15497_new_n2876_));
INVX1 INVX1_396 ( .A(_abc_15497_new_n2879_), .Y(_abc_15497_new_n2880_));
INVX1 INVX1_397 ( .A(_abc_15497_new_n2883_), .Y(_abc_15497_new_n2884_));
INVX1 INVX1_398 ( .A(_abc_15497_new_n2887_), .Y(_abc_15497_new_n2888_));
INVX1 INVX1_399 ( .A(_abc_15497_new_n2892_), .Y(_abc_15497_new_n2893_));
INVX1 INVX1_4 ( .A(_abc_15497_new_n707_), .Y(_abc_15497_new_n708_));
INVX1 INVX1_40 ( .A(_abc_15497_new_n903_), .Y(_abc_15497_new_n904_));
INVX1 INVX1_400 ( .A(_abc_15497_new_n2895_), .Y(_abc_15497_new_n2896_));
INVX1 INVX1_401 ( .A(_abc_15497_new_n2897_), .Y(_abc_15497_new_n2899_));
INVX1 INVX1_402 ( .A(_abc_15497_new_n2908_), .Y(_abc_15497_new_n2909_));
INVX1 INVX1_403 ( .A(_abc_15497_new_n2894_), .Y(_abc_15497_new_n2911_));
INVX1 INVX1_404 ( .A(_abc_15497_new_n2914_), .Y(_abc_15497_new_n2915_));
INVX1 INVX1_405 ( .A(_abc_15497_new_n2917_), .Y(_abc_15497_new_n2918_));
INVX1 INVX1_406 ( .A(_abc_15497_new_n2923_), .Y(_abc_15497_new_n2924_));
INVX1 INVX1_407 ( .A(_abc_15497_new_n2926_), .Y(_abc_15497_new_n2927_));
INVX1 INVX1_408 ( .A(_abc_15497_new_n2928_), .Y(_abc_15497_new_n2930_));
INVX1 INVX1_409 ( .A(_abc_15497_new_n2936_), .Y(_abc_15497_new_n2937_));
INVX1 INVX1_41 ( .A(_abc_15497_new_n907_), .Y(_abc_15497_new_n908_));
INVX1 INVX1_410 ( .A(_abc_15497_new_n2939_), .Y(_abc_15497_new_n2940_));
INVX1 INVX1_411 ( .A(_abc_15497_new_n2942_), .Y(_abc_15497_new_n2943_));
INVX1 INVX1_412 ( .A(_abc_15497_new_n2949_), .Y(_abc_15497_new_n2950_));
INVX1 INVX1_413 ( .A(_abc_15497_new_n2953_), .Y(_abc_15497_new_n2954_));
INVX1 INVX1_414 ( .A(_abc_15497_new_n2962_), .Y(_abc_15497_new_n2963_));
INVX1 INVX1_415 ( .A(_abc_15497_new_n2968_), .Y(_abc_15497_new_n2969_));
INVX1 INVX1_416 ( .A(_abc_15497_new_n2970_), .Y(_abc_15497_new_n2971_));
INVX1 INVX1_417 ( .A(_abc_15497_new_n2977_), .Y(_abc_15497_new_n2978_));
INVX1 INVX1_418 ( .A(_abc_15497_new_n2980_), .Y(_abc_15497_new_n2981_));
INVX1 INVX1_419 ( .A(_abc_15497_new_n2984_), .Y(_abc_15497_new_n2985_));
INVX1 INVX1_42 ( .A(_abc_15497_new_n915_), .Y(_abc_15497_new_n916_));
INVX1 INVX1_420 ( .A(_abc_15497_new_n2992_), .Y(_abc_15497_new_n2993_));
INVX1 INVX1_421 ( .A(_abc_15497_new_n2995_), .Y(_abc_15497_new_n2996_));
INVX1 INVX1_422 ( .A(_abc_15497_new_n2997_), .Y(_abc_15497_new_n2999_));
INVX1 INVX1_423 ( .A(_abc_15497_new_n2976_), .Y(_abc_15497_new_n3008_));
INVX1 INVX1_424 ( .A(_abc_15497_new_n3015_), .Y(_abc_15497_new_n3016_));
INVX1 INVX1_425 ( .A(_abc_15497_new_n3019_), .Y(_abc_15497_new_n3020_));
INVX1 INVX1_426 ( .A(_abc_15497_new_n3026_), .Y(_abc_15497_new_n3027_));
INVX1 INVX1_427 ( .A(_abc_15497_new_n3034_), .Y(_abc_15497_new_n3035_));
INVX1 INVX1_428 ( .A(_abc_15497_new_n3039_), .Y(_abc_15497_new_n3040_));
INVX1 INVX1_429 ( .A(_abc_15497_new_n3042_), .Y(_abc_15497_new_n3043_));
INVX1 INVX1_43 ( .A(_abc_15497_new_n918_), .Y(_abc_15497_new_n919_));
INVX1 INVX1_430 ( .A(_abc_15497_new_n3046_), .Y(_abc_15497_new_n3047_));
INVX1 INVX1_431 ( .A(_abc_15497_new_n3054_), .Y(_abc_15497_new_n3055_));
INVX1 INVX1_432 ( .A(_abc_15497_new_n3057_), .Y(_abc_15497_new_n3058_));
INVX1 INVX1_433 ( .A(_abc_15497_new_n3059_), .Y(_abc_15497_new_n3061_));
INVX1 INVX1_434 ( .A(_abc_15497_new_n3076_), .Y(_abc_15497_new_n3077_));
INVX1 INVX1_435 ( .A(_abc_15497_new_n3080_), .Y(_abc_15497_new_n3081_));
INVX1 INVX1_436 ( .A(_abc_15497_new_n3087_), .Y(_abc_15497_new_n3088_));
INVX1 INVX1_437 ( .A(_abc_15497_new_n3090_), .Y(_abc_15497_new_n3091_));
INVX1 INVX1_438 ( .A(_abc_15497_new_n3092_), .Y(_abc_15497_new_n3094_));
INVX1 INVX1_439 ( .A(_abc_15497_new_n3107_), .Y(_abc_15497_new_n3108_));
INVX1 INVX1_44 ( .A(_abc_15497_new_n920_), .Y(_abc_15497_new_n922_));
INVX1 INVX1_440 ( .A(_abc_15497_new_n3111_), .Y(_abc_15497_new_n3112_));
INVX1 INVX1_441 ( .A(_abc_15497_new_n3120_), .Y(_abc_15497_new_n3121_));
INVX1 INVX1_442 ( .A(_abc_15497_new_n3122_), .Y(_abc_15497_new_n3125_));
INVX1 INVX1_443 ( .A(_abc_15497_new_n3135_), .Y(_abc_15497_new_n3136_));
INVX1 INVX1_444 ( .A(_abc_15497_new_n3138_), .Y(_abc_15497_new_n3139_));
INVX1 INVX1_445 ( .A(_abc_15497_new_n3140_), .Y(_abc_15497_new_n3141_));
INVX1 INVX1_446 ( .A(_abc_15497_new_n3144_), .Y(_abc_15497_new_n3145_));
INVX1 INVX1_447 ( .A(_abc_15497_new_n3148_), .Y(_abc_15497_new_n3149_));
INVX1 INVX1_448 ( .A(_abc_15497_new_n3155_), .Y(_abc_15497_new_n3156_));
INVX1 INVX1_449 ( .A(_abc_15497_new_n3157_), .Y(_abc_15497_new_n3158_));
INVX1 INVX1_45 ( .A(_abc_15497_new_n928_), .Y(_abc_15497_new_n929_));
INVX1 INVX1_450 ( .A(_abc_15497_new_n3153_), .Y(_abc_15497_new_n3160_));
INVX1 INVX1_451 ( .A(_abc_15497_new_n3168_), .Y(_abc_15497_new_n3169_));
INVX1 INVX1_452 ( .A(_abc_15497_new_n3177_), .Y(_abc_15497_new_n3178_));
INVX1 INVX1_453 ( .A(_abc_15497_new_n3185_), .Y(_abc_15497_new_n3186_));
INVX1 INVX1_454 ( .A(_abc_15497_new_n3188_), .Y(_abc_15497_new_n3189_));
INVX1 INVX1_455 ( .A(_abc_15497_new_n3190_), .Y(_abc_15497_new_n3191_));
INVX1 INVX1_456 ( .A(_abc_15497_new_n3738_), .Y(_abc_15497_new_n3739_));
INVX1 INVX1_457 ( .A(round_ctr_reg_6_), .Y(_abc_15497_new_n3740_));
INVX1 INVX1_458 ( .A(_abc_15497_new_n3741_), .Y(_abc_15497_new_n3742_));
INVX1 INVX1_459 ( .A(round_ctr_reg_5_), .Y(_abc_15497_new_n3745_));
INVX1 INVX1_46 ( .A(_abc_15497_new_n931_), .Y(_abc_15497_new_n932_));
INVX1 INVX1_460 ( .A(round_ctr_reg_4_), .Y(_abc_15497_new_n3746_));
INVX1 INVX1_461 ( .A(round_ctr_reg_2_), .Y(_abc_15497_new_n3748_));
INVX1 INVX1_462 ( .A(round_ctr_reg_3_), .Y(_abc_15497_new_n3749_));
INVX1 INVX1_463 ( .A(c_reg_0_), .Y(_abc_15497_new_n3754_));
INVX1 INVX1_464 ( .A(d_reg_0_), .Y(_abc_15497_new_n3756_));
INVX1 INVX1_465 ( .A(_abc_15497_new_n3757_), .Y(_abc_15497_new_n3758_));
INVX1 INVX1_466 ( .A(_abc_15497_new_n3763_), .Y(_abc_15497_new_n3764_));
INVX1 INVX1_467 ( .A(_abc_15497_new_n3771_), .Y(_abc_15497_new_n3772_));
INVX1 INVX1_468 ( .A(_abc_15497_new_n3762_), .Y(_abc_15497_new_n3781_));
INVX1 INVX1_469 ( .A(_abc_15497_new_n3790_), .Y(_abc_15497_new_n3791_));
INVX1 INVX1_47 ( .A(_abc_15497_new_n934_), .Y(_abc_15497_new_n935_));
INVX1 INVX1_470 ( .A(w_0_), .Y(_abc_15497_new_n3794_));
INVX1 INVX1_471 ( .A(_abc_15497_new_n3792_), .Y(_abc_15497_new_n3795_));
INVX1 INVX1_472 ( .A(_abc_15497_new_n3761_), .Y(_abc_15497_new_n3799_));
INVX1 INVX1_473 ( .A(_abc_15497_new_n3765_), .Y(_abc_15497_new_n3800_));
INVX1 INVX1_474 ( .A(_abc_15497_new_n3766_), .Y(_abc_15497_new_n3801_));
INVX1 INVX1_475 ( .A(_abc_15497_new_n3782_), .Y(_abc_15497_new_n3805_));
INVX1 INVX1_476 ( .A(_abc_15497_new_n3797_), .Y(_abc_15497_new_n3810_));
INVX1 INVX1_477 ( .A(_abc_15497_new_n3812_), .Y(_abc_15497_new_n3813_));
INVX1 INVX1_478 ( .A(_abc_15497_new_n3815_), .Y(_abc_15497_new_n3816_));
INVX1 INVX1_479 ( .A(_abc_15497_new_n3825_), .Y(_abc_15497_new_n3826_));
INVX1 INVX1_48 ( .A(_abc_15497_new_n898_), .Y(_abc_15497_new_n936_));
INVX1 INVX1_480 ( .A(_abc_15497_new_n3828_), .Y(_abc_15497_new_n3829_));
INVX1 INVX1_481 ( .A(d_reg_1_), .Y(_abc_15497_new_n3833_));
INVX1 INVX1_482 ( .A(_abc_15497_new_n3824_), .Y(_abc_15497_new_n3837_));
INVX1 INVX1_483 ( .A(_abc_15497_new_n3845_), .Y(_abc_15497_new_n3846_));
INVX1 INVX1_484 ( .A(_abc_15497_new_n3849_), .Y(_abc_15497_new_n3850_));
INVX1 INVX1_485 ( .A(_abc_15497_new_n3852_), .Y(_abc_15497_new_n3853_));
INVX1 INVX1_486 ( .A(_abc_15497_new_n3830_), .Y(_abc_15497_new_n3857_));
INVX1 INVX1_487 ( .A(_abc_15497_new_n3835_), .Y(_abc_15497_new_n3860_));
INVX1 INVX1_488 ( .A(_abc_15497_new_n3839_), .Y(_abc_15497_new_n3862_));
INVX1 INVX1_489 ( .A(_abc_15497_new_n3843_), .Y(_abc_15497_new_n3866_));
INVX1 INVX1_49 ( .A(_abc_15497_new_n780_), .Y(_abc_15497_new_n937_));
INVX1 INVX1_490 ( .A(_abc_15497_new_n3848_), .Y(_abc_15497_new_n3867_));
INVX1 INVX1_491 ( .A(_abc_15497_new_n3884_), .Y(_abc_15497_new_n3885_));
INVX1 INVX1_492 ( .A(_abc_15497_new_n3887_), .Y(_abc_15497_new_n3895_));
INVX1 INVX1_493 ( .A(_abc_15497_new_n3901_), .Y(_abc_15497_new_n3902_));
INVX1 INVX1_494 ( .A(_abc_15497_new_n3905_), .Y(_abc_15497_new_n3906_));
INVX1 INVX1_495 ( .A(_abc_15497_new_n3907_), .Y(_abc_15497_new_n3908_));
INVX1 INVX1_496 ( .A(d_reg_2_), .Y(_abc_15497_new_n3910_));
INVX1 INVX1_497 ( .A(_abc_15497_new_n3900_), .Y(_abc_15497_new_n3914_));
INVX1 INVX1_498 ( .A(_abc_15497_new_n3922_), .Y(_abc_15497_new_n3923_));
INVX1 INVX1_499 ( .A(_abc_15497_new_n3926_), .Y(_abc_15497_new_n3927_));
INVX1 INVX1_5 ( .A(_abc_15497_new_n711_), .Y(_abc_15497_new_n712_));
INVX1 INVX1_50 ( .A(_abc_15497_new_n784_), .Y(_abc_15497_new_n938_));
INVX1 INVX1_500 ( .A(_abc_15497_new_n3920_), .Y(_abc_15497_new_n3930_));
INVX1 INVX1_501 ( .A(_abc_15497_new_n3925_), .Y(_abc_15497_new_n3931_));
INVX1 INVX1_502 ( .A(_abc_15497_new_n3912_), .Y(_abc_15497_new_n3937_));
INVX1 INVX1_503 ( .A(_abc_15497_new_n3916_), .Y(_abc_15497_new_n3939_));
INVX1 INVX1_504 ( .A(_abc_15497_new_n3929_), .Y(_abc_15497_new_n3943_));
INVX1 INVX1_505 ( .A(_abc_15497_new_n3981_), .Y(_abc_15497_new_n3982_));
INVX1 INVX1_506 ( .A(d_reg_3_), .Y(_abc_15497_new_n3984_));
INVX1 INVX1_507 ( .A(_abc_15497_new_n3986_), .Y(_abc_15497_new_n3987_));
INVX1 INVX1_508 ( .A(_abc_15497_new_n3988_), .Y(_abc_15497_new_n3989_));
INVX1 INVX1_509 ( .A(_abc_15497_new_n3985_), .Y(_abc_15497_new_n3997_));
INVX1 INVX1_51 ( .A(_abc_15497_new_n789_), .Y(_abc_15497_new_n939_));
INVX1 INVX1_510 ( .A(_abc_15497_new_n4003_), .Y(_abc_15497_new_n4004_));
INVX1 INVX1_511 ( .A(w_3_), .Y(_abc_15497_new_n4005_));
INVX1 INVX1_512 ( .A(_abc_15497_new_n4007_), .Y(_abc_15497_new_n4008_));
INVX1 INVX1_513 ( .A(_abc_15497_new_n4009_), .Y(_abc_15497_new_n4010_));
INVX1 INVX1_514 ( .A(_abc_15497_new_n4013_), .Y(_abc_15497_new_n4014_));
INVX1 INVX1_515 ( .A(_abc_15497_new_n4018_), .Y(_abc_15497_new_n4019_));
INVX1 INVX1_516 ( .A(_abc_15497_new_n3983_), .Y(_abc_15497_new_n4023_));
INVX1 INVX1_517 ( .A(_abc_15497_new_n4020_), .Y(_abc_15497_new_n4024_));
INVX1 INVX1_518 ( .A(_abc_15497_new_n3980_), .Y(_abc_15497_new_n4041_));
INVX1 INVX1_519 ( .A(_abc_15497_new_n4059_), .Y(_abc_15497_new_n4060_));
INVX1 INVX1_52 ( .A(_abc_15497_new_n795_), .Y(_abc_15497_new_n940_));
INVX1 INVX1_520 ( .A(_abc_15497_new_n4015_), .Y(_abc_15497_new_n4061_));
INVX1 INVX1_521 ( .A(d_reg_4_), .Y(_abc_15497_new_n4063_));
INVX1 INVX1_522 ( .A(_abc_15497_new_n4065_), .Y(_abc_15497_new_n4066_));
INVX1 INVX1_523 ( .A(_abc_15497_new_n4067_), .Y(_abc_15497_new_n4068_));
INVX1 INVX1_524 ( .A(_abc_15497_new_n4071_), .Y(_abc_15497_new_n4072_));
INVX1 INVX1_525 ( .A(b_reg_4_), .Y(_abc_15497_new_n4074_));
INVX1 INVX1_526 ( .A(_abc_15497_new_n4064_), .Y(_abc_15497_new_n4078_));
INVX1 INVX1_527 ( .A(_abc_15497_new_n4080_), .Y(_abc_15497_new_n4081_));
INVX1 INVX1_528 ( .A(w_4_), .Y(_abc_15497_new_n4086_));
INVX1 INVX1_529 ( .A(_abc_15497_new_n4088_), .Y(_abc_15497_new_n4089_));
INVX1 INVX1_53 ( .A(_abc_15497_new_n800_), .Y(_abc_15497_new_n941_));
INVX1 INVX1_530 ( .A(_abc_15497_new_n4090_), .Y(_abc_15497_new_n4091_));
INVX1 INVX1_531 ( .A(_abc_15497_new_n4094_), .Y(_abc_15497_new_n4095_));
INVX1 INVX1_532 ( .A(_abc_15497_new_n4085_), .Y(_abc_15497_new_n4097_));
INVX1 INVX1_533 ( .A(_abc_15497_new_n4099_), .Y(_abc_15497_new_n4100_));
INVX1 INVX1_534 ( .A(_abc_15497_new_n4084_), .Y(_abc_15497_new_n4102_));
INVX1 INVX1_535 ( .A(_abc_15497_new_n4062_), .Y(_abc_15497_new_n4106_));
INVX1 INVX1_536 ( .A(_abc_15497_new_n4124_), .Y(_abc_15497_new_n4125_));
INVX1 INVX1_537 ( .A(_abc_15497_new_n4127_), .Y(_abc_15497_new_n4128_));
INVX1 INVX1_538 ( .A(_abc_15497_new_n4137_), .Y(_abc_15497_new_n4138_));
INVX1 INVX1_539 ( .A(d_reg_5_), .Y(_abc_15497_new_n4141_));
INVX1 INVX1_54 ( .A(_abc_15497_new_n805_), .Y(_abc_15497_new_n942_));
INVX1 INVX1_540 ( .A(_abc_15497_new_n4143_), .Y(_abc_15497_new_n4144_));
INVX1 INVX1_541 ( .A(_abc_15497_new_n4145_), .Y(_abc_15497_new_n4146_));
INVX1 INVX1_542 ( .A(_abc_15497_new_n4149_), .Y(_abc_15497_new_n4150_));
INVX1 INVX1_543 ( .A(b_reg_5_), .Y(_abc_15497_new_n4152_));
INVX1 INVX1_544 ( .A(_abc_15497_new_n4142_), .Y(_abc_15497_new_n4156_));
INVX1 INVX1_545 ( .A(_abc_15497_new_n4158_), .Y(_abc_15497_new_n4159_));
INVX1 INVX1_546 ( .A(_abc_15497_new_n4162_), .Y(_abc_15497_new_n4163_));
INVX1 INVX1_547 ( .A(w_5_), .Y(_abc_15497_new_n4165_));
INVX1 INVX1_548 ( .A(_abc_15497_new_n4167_), .Y(_abc_15497_new_n4168_));
INVX1 INVX1_549 ( .A(_abc_15497_new_n4169_), .Y(_abc_15497_new_n4170_));
INVX1 INVX1_55 ( .A(_abc_15497_new_n811_), .Y(_abc_15497_new_n943_));
INVX1 INVX1_550 ( .A(_abc_15497_new_n4173_), .Y(_abc_15497_new_n4174_));
INVX1 INVX1_551 ( .A(_abc_15497_new_n4164_), .Y(_abc_15497_new_n4176_));
INVX1 INVX1_552 ( .A(_abc_15497_new_n4178_), .Y(_abc_15497_new_n4180_));
INVX1 INVX1_553 ( .A(_abc_15497_new_n4096_), .Y(_abc_15497_new_n4184_));
INVX1 INVX1_554 ( .A(_abc_15497_new_n4203_), .Y(_abc_15497_new_n4204_));
INVX1 INVX1_555 ( .A(_abc_15497_new_n4214_), .Y(_abc_15497_new_n4215_));
INVX1 INVX1_556 ( .A(_abc_15497_new_n4197_), .Y(_abc_15497_new_n4217_));
INVX1 INVX1_557 ( .A(_abc_15497_new_n4219_), .Y(_abc_15497_new_n4220_));
INVX1 INVX1_558 ( .A(d_reg_6_), .Y(_abc_15497_new_n4224_));
INVX1 INVX1_559 ( .A(_abc_15497_new_n4226_), .Y(_abc_15497_new_n4227_));
INVX1 INVX1_56 ( .A(_abc_15497_new_n812_), .Y(_abc_15497_new_n944_));
INVX1 INVX1_560 ( .A(_abc_15497_new_n4228_), .Y(_abc_15497_new_n4229_));
INVX1 INVX1_561 ( .A(_abc_15497_new_n4232_), .Y(_abc_15497_new_n4233_));
INVX1 INVX1_562 ( .A(b_reg_6_), .Y(_abc_15497_new_n4235_));
INVX1 INVX1_563 ( .A(_abc_15497_new_n4225_), .Y(_abc_15497_new_n4239_));
INVX1 INVX1_564 ( .A(_abc_15497_new_n4241_), .Y(_abc_15497_new_n4242_));
INVX1 INVX1_565 ( .A(_abc_15497_new_n4245_), .Y(_abc_15497_new_n4246_));
INVX1 INVX1_566 ( .A(w_6_), .Y(_abc_15497_new_n4248_));
INVX1 INVX1_567 ( .A(_abc_15497_new_n4250_), .Y(_abc_15497_new_n4251_));
INVX1 INVX1_568 ( .A(_abc_15497_new_n4252_), .Y(_abc_15497_new_n4253_));
INVX1 INVX1_569 ( .A(_abc_15497_new_n4256_), .Y(_abc_15497_new_n4257_));
INVX1 INVX1_57 ( .A(_abc_15497_new_n813_), .Y(_abc_15497_new_n945_));
INVX1 INVX1_570 ( .A(_abc_15497_new_n4247_), .Y(_abc_15497_new_n4259_));
INVX1 INVX1_571 ( .A(_abc_15497_new_n4261_), .Y(_abc_15497_new_n4263_));
INVX1 INVX1_572 ( .A(_abc_15497_new_n4175_), .Y(_abc_15497_new_n4267_));
INVX1 INVX1_573 ( .A(_abc_15497_new_n4286_), .Y(_abc_15497_new_n4287_));
INVX1 INVX1_574 ( .A(_abc_15497_new_n4289_), .Y(_abc_15497_new_n4290_));
INVX1 INVX1_575 ( .A(_abc_15497_new_n4280_), .Y(_abc_15497_new_n4298_));
INVX1 INVX1_576 ( .A(_abc_15497_new_n4258_), .Y(_abc_15497_new_n4301_));
INVX1 INVX1_577 ( .A(_abc_15497_new_n4302_), .Y(_abc_15497_new_n4303_));
INVX1 INVX1_578 ( .A(d_reg_7_), .Y(_abc_15497_new_n4304_));
INVX1 INVX1_579 ( .A(_abc_15497_new_n4306_), .Y(_abc_15497_new_n4307_));
INVX1 INVX1_58 ( .A(_abc_15497_new_n815_), .Y(_abc_15497_new_n946_));
INVX1 INVX1_580 ( .A(_abc_15497_new_n4308_), .Y(_abc_15497_new_n4309_));
INVX1 INVX1_581 ( .A(b_reg_7_), .Y(_abc_15497_new_n4314_));
INVX1 INVX1_582 ( .A(_abc_15497_new_n4317_), .Y(_abc_15497_new_n4318_));
INVX1 INVX1_583 ( .A(_abc_15497_new_n4305_), .Y(_abc_15497_new_n4319_));
INVX1 INVX1_584 ( .A(_abc_15497_new_n4324_), .Y(_abc_15497_new_n4325_));
INVX1 INVX1_585 ( .A(w_7_), .Y(_abc_15497_new_n4327_));
INVX1 INVX1_586 ( .A(_abc_15497_new_n4329_), .Y(_abc_15497_new_n4330_));
INVX1 INVX1_587 ( .A(_abc_15497_new_n4331_), .Y(_abc_15497_new_n4332_));
INVX1 INVX1_588 ( .A(_abc_15497_new_n4335_), .Y(_abc_15497_new_n4336_));
INVX1 INVX1_589 ( .A(_abc_15497_new_n4337_), .Y(_abc_15497_new_n4338_));
INVX1 INVX1_59 ( .A(_abc_15497_new_n816_), .Y(_abc_15497_new_n947_));
INVX1 INVX1_590 ( .A(_abc_15497_new_n4339_), .Y(_abc_15497_new_n4342_));
INVX1 INVX1_591 ( .A(_abc_15497_new_n4345_), .Y(_abc_15497_new_n4346_));
INVX1 INVX1_592 ( .A(_abc_15497_new_n4349_), .Y(_abc_15497_new_n4352_));
INVX1 INVX1_593 ( .A(_abc_15497_new_n4299_), .Y(_abc_15497_new_n4356_));
INVX1 INVX1_594 ( .A(_abc_15497_new_n4354_), .Y(_abc_15497_new_n4357_));
INVX1 INVX1_595 ( .A(_abc_15497_new_n4348_), .Y(_abc_15497_new_n4366_));
INVX1 INVX1_596 ( .A(d_reg_8_), .Y(_abc_15497_new_n4368_));
INVX1 INVX1_597 ( .A(_abc_15497_new_n4370_), .Y(_abc_15497_new_n4371_));
INVX1 INVX1_598 ( .A(_abc_15497_new_n4372_), .Y(_abc_15497_new_n4373_));
INVX1 INVX1_599 ( .A(b_reg_8_), .Y(_abc_15497_new_n4378_));
INVX1 INVX1_6 ( .A(_abc_15497_new_n713_), .Y(_abc_15497_new_n714_));
INVX1 INVX1_60 ( .A(_abc_15497_new_n819_), .Y(_abc_15497_new_n948_));
INVX1 INVX1_600 ( .A(_abc_15497_new_n4381_), .Y(_abc_15497_new_n4382_));
INVX1 INVX1_601 ( .A(_abc_15497_new_n4369_), .Y(_abc_15497_new_n4383_));
INVX1 INVX1_602 ( .A(w_8_), .Y(_abc_15497_new_n4390_));
INVX1 INVX1_603 ( .A(_abc_15497_new_n4392_), .Y(_abc_15497_new_n4393_));
INVX1 INVX1_604 ( .A(_abc_15497_new_n4394_), .Y(_abc_15497_new_n4395_));
INVX1 INVX1_605 ( .A(_abc_15497_new_n4398_), .Y(_abc_15497_new_n4399_));
INVX1 INVX1_606 ( .A(_abc_15497_new_n4401_), .Y(_abc_15497_new_n4402_));
INVX1 INVX1_607 ( .A(_abc_15497_new_n4388_), .Y(_abc_15497_new_n4405_));
INVX1 INVX1_608 ( .A(_abc_15497_new_n4400_), .Y(_abc_15497_new_n4406_));
INVX1 INVX1_609 ( .A(_abc_15497_new_n4423_), .Y(_abc_15497_new_n4424_));
INVX1 INVX1_61 ( .A(_abc_15497_new_n821_), .Y(_abc_15497_new_n949_));
INVX1 INVX1_610 ( .A(_abc_15497_new_n4427_), .Y(_abc_15497_new_n4428_));
INVX1 INVX1_611 ( .A(_abc_15497_new_n4055_), .Y(_abc_15497_new_n4430_));
INVX1 INVX1_612 ( .A(_abc_15497_new_n4350_), .Y(_abc_15497_new_n4436_));
INVX1 INVX1_613 ( .A(_abc_15497_new_n4441_), .Y(_abc_15497_new_n4442_));
INVX1 INVX1_614 ( .A(_abc_15497_new_n4444_), .Y(_abc_15497_new_n4445_));
INVX1 INVX1_615 ( .A(_abc_15497_new_n4455_), .Y(_abc_15497_new_n4456_));
INVX1 INVX1_616 ( .A(d_reg_9_), .Y(_abc_15497_new_n4458_));
INVX1 INVX1_617 ( .A(_abc_15497_new_n4460_), .Y(_abc_15497_new_n4461_));
INVX1 INVX1_618 ( .A(_abc_15497_new_n4462_), .Y(_abc_15497_new_n4463_));
INVX1 INVX1_619 ( .A(b_reg_9_), .Y(_abc_15497_new_n4468_));
INVX1 INVX1_62 ( .A(_abc_15497_new_n827_), .Y(_abc_15497_new_n953_));
INVX1 INVX1_620 ( .A(_abc_15497_new_n4471_), .Y(_abc_15497_new_n4472_));
INVX1 INVX1_621 ( .A(_abc_15497_new_n4459_), .Y(_abc_15497_new_n4473_));
INVX1 INVX1_622 ( .A(_abc_15497_new_n4478_), .Y(_abc_15497_new_n4479_));
INVX1 INVX1_623 ( .A(w_9_), .Y(_abc_15497_new_n4481_));
INVX1 INVX1_624 ( .A(_abc_15497_new_n4483_), .Y(_abc_15497_new_n4484_));
INVX1 INVX1_625 ( .A(_abc_15497_new_n4485_), .Y(_abc_15497_new_n4486_));
INVX1 INVX1_626 ( .A(_abc_15497_new_n4489_), .Y(_abc_15497_new_n4490_));
INVX1 INVX1_627 ( .A(_abc_15497_new_n4491_), .Y(_abc_15497_new_n4492_));
INVX1 INVX1_628 ( .A(_abc_15497_new_n4493_), .Y(_abc_15497_new_n4496_));
INVX1 INVX1_629 ( .A(_abc_15497_new_n4512_), .Y(_abc_15497_new_n4513_));
INVX1 INVX1_63 ( .A(_abc_15497_new_n834_), .Y(_abc_15497_new_n958_));
INVX1 INVX1_630 ( .A(_abc_15497_new_n4453_), .Y(_abc_15497_new_n4518_));
INVX1 INVX1_631 ( .A(_abc_15497_new_n4516_), .Y(_abc_15497_new_n4519_));
INVX1 INVX1_632 ( .A(_abc_15497_new_n4514_), .Y(_abc_15497_new_n4527_));
INVX1 INVX1_633 ( .A(_abc_15497_new_n4529_), .Y(_abc_15497_new_n4530_));
INVX1 INVX1_634 ( .A(_abc_15497_new_n4531_), .Y(_abc_15497_new_n4532_));
INVX1 INVX1_635 ( .A(d_reg_10_), .Y(_abc_15497_new_n4537_));
INVX1 INVX1_636 ( .A(_abc_15497_new_n4539_), .Y(_abc_15497_new_n4540_));
INVX1 INVX1_637 ( .A(_abc_15497_new_n4541_), .Y(_abc_15497_new_n4542_));
INVX1 INVX1_638 ( .A(b_reg_10_), .Y(_abc_15497_new_n4547_));
INVX1 INVX1_639 ( .A(_abc_15497_new_n4550_), .Y(_abc_15497_new_n4551_));
INVX1 INVX1_64 ( .A(_abc_15497_new_n846_), .Y(_abc_15497_new_n965_));
INVX1 INVX1_640 ( .A(_abc_15497_new_n4538_), .Y(_abc_15497_new_n4552_));
INVX1 INVX1_641 ( .A(w_10_), .Y(_abc_15497_new_n4559_));
INVX1 INVX1_642 ( .A(_abc_15497_new_n4561_), .Y(_abc_15497_new_n4562_));
INVX1 INVX1_643 ( .A(_abc_15497_new_n4563_), .Y(_abc_15497_new_n4564_));
INVX1 INVX1_644 ( .A(_abc_15497_new_n4567_), .Y(_abc_15497_new_n4568_));
INVX1 INVX1_645 ( .A(_abc_15497_new_n4570_), .Y(_abc_15497_new_n4571_));
INVX1 INVX1_646 ( .A(_abc_15497_new_n4557_), .Y(_abc_15497_new_n4574_));
INVX1 INVX1_647 ( .A(_abc_15497_new_n4569_), .Y(_abc_15497_new_n4575_));
INVX1 INVX1_648 ( .A(_abc_15497_new_n4599_), .Y(_abc_15497_new_n4600_));
INVX1 INVX1_649 ( .A(_abc_15497_new_n4602_), .Y(_abc_15497_new_n4603_));
INVX1 INVX1_65 ( .A(_abc_15497_new_n857_), .Y(_abc_15497_new_n972_));
INVX1 INVX1_650 ( .A(_abc_15497_new_n4592_), .Y(_abc_15497_new_n4611_));
INVX1 INVX1_651 ( .A(d_reg_11_), .Y(_abc_15497_new_n4615_));
INVX1 INVX1_652 ( .A(_abc_15497_new_n4617_), .Y(_abc_15497_new_n4618_));
INVX1 INVX1_653 ( .A(_abc_15497_new_n4619_), .Y(_abc_15497_new_n4620_));
INVX1 INVX1_654 ( .A(b_reg_11_), .Y(_abc_15497_new_n4625_));
INVX1 INVX1_655 ( .A(_abc_15497_new_n4628_), .Y(_abc_15497_new_n4629_));
INVX1 INVX1_656 ( .A(_abc_15497_new_n4616_), .Y(_abc_15497_new_n4630_));
INVX1 INVX1_657 ( .A(_abc_15497_new_n4635_), .Y(_abc_15497_new_n4636_));
INVX1 INVX1_658 ( .A(w_11_), .Y(_abc_15497_new_n4638_));
INVX1 INVX1_659 ( .A(_abc_15497_new_n4640_), .Y(_abc_15497_new_n4641_));
INVX1 INVX1_66 ( .A(_abc_15497_new_n868_), .Y(_abc_15497_new_n975_));
INVX1 INVX1_660 ( .A(_abc_15497_new_n4642_), .Y(_abc_15497_new_n4643_));
INVX1 INVX1_661 ( .A(_abc_15497_new_n4646_), .Y(_abc_15497_new_n4647_));
INVX1 INVX1_662 ( .A(_abc_15497_new_n4648_), .Y(_abc_15497_new_n4649_));
INVX1 INVX1_663 ( .A(_abc_15497_new_n4650_), .Y(_abc_15497_new_n4653_));
INVX1 INVX1_664 ( .A(_abc_15497_new_n4612_), .Y(_abc_15497_new_n4678_));
INVX1 INVX1_665 ( .A(_abc_15497_new_n4676_), .Y(_abc_15497_new_n4679_));
INVX1 INVX1_666 ( .A(_abc_15497_new_n4670_), .Y(_abc_15497_new_n4690_));
INVX1 INVX1_667 ( .A(_abc_15497_new_n4693_), .Y(_abc_15497_new_n4694_));
INVX1 INVX1_668 ( .A(_abc_15497_new_n4695_), .Y(_abc_15497_new_n4696_));
INVX1 INVX1_669 ( .A(_abc_15497_new_n4700_), .Y(_abc_15497_new_n4701_));
INVX1 INVX1_67 ( .A(_abc_15497_new_n871_), .Y(_abc_15497_new_n977_));
INVX1 INVX1_670 ( .A(_abc_15497_new_n4703_), .Y(_abc_15497_new_n4704_));
INVX1 INVX1_671 ( .A(_abc_15497_new_n4707_), .Y(_abc_15497_new_n4708_));
INVX1 INVX1_672 ( .A(_abc_15497_new_n4710_), .Y(_abc_15497_new_n4711_));
INVX1 INVX1_673 ( .A(d_reg_12_), .Y(_abc_15497_new_n4712_));
INVX1 INVX1_674 ( .A(_abc_15497_new_n4702_), .Y(_abc_15497_new_n4716_));
INVX1 INVX1_675 ( .A(_abc_15497_new_n4721_), .Y(_abc_15497_new_n4722_));
INVX1 INVX1_676 ( .A(w_12_), .Y(_abc_15497_new_n4724_));
INVX1 INVX1_677 ( .A(_abc_15497_new_n4726_), .Y(_abc_15497_new_n4727_));
INVX1 INVX1_678 ( .A(_abc_15497_new_n4728_), .Y(_abc_15497_new_n4729_));
INVX1 INVX1_679 ( .A(_abc_15497_new_n4732_), .Y(_abc_15497_new_n4733_));
INVX1 INVX1_68 ( .A(_abc_15497_new_n899_), .Y(_abc_15497_new_n979_));
INVX1 INVX1_680 ( .A(_abc_15497_new_n4734_), .Y(_abc_15497_new_n4735_));
INVX1 INVX1_681 ( .A(_abc_15497_new_n4738_), .Y(_abc_15497_new_n4739_));
INVX1 INVX1_682 ( .A(_abc_15497_new_n4743_), .Y(_abc_15497_new_n4744_));
INVX1 INVX1_683 ( .A(_abc_15497_new_n4740_), .Y(_abc_15497_new_n4747_));
INVX1 INVX1_684 ( .A(_abc_15497_new_n4699_), .Y(_abc_15497_new_n4754_));
INVX1 INVX1_685 ( .A(_abc_15497_new_n4759_), .Y(_abc_15497_new_n4760_));
INVX1 INVX1_686 ( .A(_abc_15497_new_n4762_), .Y(_abc_15497_new_n4763_));
INVX1 INVX1_687 ( .A(_abc_15497_new_n4776_), .Y(_abc_15497_new_n4777_));
INVX1 INVX1_688 ( .A(_abc_15497_new_n4780_), .Y(_abc_15497_new_n4781_));
INVX1 INVX1_689 ( .A(_abc_15497_new_n4783_), .Y(_abc_15497_new_n4784_));
INVX1 INVX1_69 ( .A(_abc_15497_new_n982_), .Y(_abc_15497_new_n983_));
INVX1 INVX1_690 ( .A(d_reg_13_), .Y(_abc_15497_new_n4785_));
INVX1 INVX1_691 ( .A(_abc_15497_new_n4775_), .Y(_abc_15497_new_n4789_));
INVX1 INVX1_692 ( .A(_abc_15497_new_n4794_), .Y(_abc_15497_new_n4795_));
INVX1 INVX1_693 ( .A(w_13_), .Y(_abc_15497_new_n4797_));
INVX1 INVX1_694 ( .A(_abc_15497_new_n4799_), .Y(_abc_15497_new_n4800_));
INVX1 INVX1_695 ( .A(_abc_15497_new_n4801_), .Y(_abc_15497_new_n4802_));
INVX1 INVX1_696 ( .A(_abc_15497_new_n4805_), .Y(_abc_15497_new_n4806_));
INVX1 INVX1_697 ( .A(_abc_15497_new_n4807_), .Y(_abc_15497_new_n4808_));
INVX1 INVX1_698 ( .A(_abc_15497_new_n4811_), .Y(_abc_15497_new_n4812_));
INVX1 INVX1_699 ( .A(_abc_15497_new_n4816_), .Y(_abc_15497_new_n4817_));
INVX1 INVX1_7 ( .A(_abc_15497_new_n715_), .Y(_abc_15497_new_n716_));
INVX1 INVX1_70 ( .A(\digest[95] ), .Y(_abc_15497_new_n995_));
INVX1 INVX1_700 ( .A(_abc_15497_new_n4774_), .Y(_abc_15497_new_n4820_));
INVX1 INVX1_701 ( .A(_abc_15497_new_n4813_), .Y(_abc_15497_new_n4821_));
INVX1 INVX1_702 ( .A(_abc_15497_new_n4772_), .Y(_abc_15497_new_n4835_));
INVX1 INVX1_703 ( .A(_abc_15497_new_n4833_), .Y(_abc_15497_new_n4836_));
INVX1 INVX1_704 ( .A(_abc_15497_new_n4827_), .Y(_abc_15497_new_n4844_));
INVX1 INVX1_705 ( .A(_abc_15497_new_n4846_), .Y(_abc_15497_new_n4847_));
INVX1 INVX1_706 ( .A(_abc_15497_new_n4848_), .Y(_abc_15497_new_n4849_));
INVX1 INVX1_707 ( .A(_abc_15497_new_n4855_), .Y(_abc_15497_new_n4856_));
INVX1 INVX1_708 ( .A(_abc_15497_new_n4859_), .Y(_abc_15497_new_n4860_));
INVX1 INVX1_709 ( .A(_abc_15497_new_n4862_), .Y(_abc_15497_new_n4863_));
INVX1 INVX1_71 ( .A(c_reg_31_), .Y(_abc_15497_new_n997_));
INVX1 INVX1_710 ( .A(d_reg_14_), .Y(_abc_15497_new_n4864_));
INVX1 INVX1_711 ( .A(_abc_15497_new_n4868_), .Y(_abc_15497_new_n4869_));
INVX1 INVX1_712 ( .A(_abc_15497_new_n4871_), .Y(_abc_15497_new_n4872_));
INVX1 INVX1_713 ( .A(_abc_15497_new_n4874_), .Y(_abc_15497_new_n4875_));
INVX1 INVX1_714 ( .A(_abc_15497_new_n4878_), .Y(_abc_15497_new_n4879_));
INVX1 INVX1_715 ( .A(_abc_15497_new_n4882_), .Y(_abc_15497_new_n4883_));
INVX1 INVX1_716 ( .A(_abc_15497_new_n4885_), .Y(_abc_15497_new_n4886_));
INVX1 INVX1_717 ( .A(_abc_15497_new_n4889_), .Y(_abc_15497_new_n4890_));
INVX1 INVX1_718 ( .A(_abc_15497_new_n4853_), .Y(_abc_15497_new_n4894_));
INVX1 INVX1_719 ( .A(_abc_15497_new_n4891_), .Y(_abc_15497_new_n4895_));
INVX1 INVX1_72 ( .A(_abc_15497_new_n999_), .Y(_abc_15497_new_n1000_));
INVX1 INVX1_720 ( .A(_abc_15497_new_n4911_), .Y(_abc_15497_new_n4912_));
INVX1 INVX1_721 ( .A(_abc_15497_new_n4914_), .Y(_abc_15497_new_n4915_));
INVX1 INVX1_722 ( .A(_abc_15497_new_n4905_), .Y(_abc_15497_new_n4923_));
INVX1 INVX1_723 ( .A(_abc_15497_new_n4928_), .Y(_abc_15497_new_n4929_));
INVX1 INVX1_724 ( .A(_abc_15497_new_n4932_), .Y(_abc_15497_new_n4933_));
INVX1 INVX1_725 ( .A(_abc_15497_new_n4935_), .Y(_abc_15497_new_n4936_));
INVX1 INVX1_726 ( .A(d_reg_15_), .Y(_abc_15497_new_n4937_));
INVX1 INVX1_727 ( .A(_abc_15497_new_n4941_), .Y(_abc_15497_new_n4942_));
INVX1 INVX1_728 ( .A(_abc_15497_new_n4944_), .Y(_abc_15497_new_n4945_));
INVX1 INVX1_729 ( .A(_abc_15497_new_n4947_), .Y(_abc_15497_new_n4948_));
INVX1 INVX1_73 ( .A(_abc_15497_new_n1009_), .Y(_abc_15497_new_n1010_));
INVX1 INVX1_730 ( .A(_abc_15497_new_n4951_), .Y(_abc_15497_new_n4952_));
INVX1 INVX1_731 ( .A(_abc_15497_new_n4955_), .Y(_abc_15497_new_n4956_));
INVX1 INVX1_732 ( .A(_abc_15497_new_n4958_), .Y(_abc_15497_new_n4959_));
INVX1 INVX1_733 ( .A(_abc_15497_new_n4962_), .Y(_abc_15497_new_n4963_));
INVX1 INVX1_734 ( .A(_abc_15497_new_n4967_), .Y(_abc_15497_new_n4968_));
INVX1 INVX1_735 ( .A(_abc_15497_new_n4926_), .Y(_abc_15497_new_n4971_));
INVX1 INVX1_736 ( .A(_abc_15497_new_n4964_), .Y(_abc_15497_new_n4972_));
INVX1 INVX1_737 ( .A(_abc_15497_new_n4924_), .Y(_abc_15497_new_n4986_));
INVX1 INVX1_738 ( .A(_abc_15497_new_n4984_), .Y(_abc_15497_new_n4987_));
INVX1 INVX1_739 ( .A(_abc_15497_new_n4978_), .Y(_abc_15497_new_n5000_));
INVX1 INVX1_74 ( .A(_abc_15497_new_n1016_), .Y(_abc_15497_new_n1017_));
INVX1 INVX1_740 ( .A(_abc_15497_new_n5007_), .Y(_abc_15497_new_n5008_));
INVX1 INVX1_741 ( .A(_abc_15497_new_n5010_), .Y(_abc_15497_new_n5011_));
INVX1 INVX1_742 ( .A(_abc_15497_new_n5012_), .Y(_abc_15497_new_n5013_));
INVX1 INVX1_743 ( .A(_abc_15497_new_n5015_), .Y(_abc_15497_new_n5016_));
INVX1 INVX1_744 ( .A(_abc_15497_new_n5018_), .Y(_abc_15497_new_n5019_));
INVX1 INVX1_745 ( .A(_abc_15497_new_n5022_), .Y(_abc_15497_new_n5023_));
INVX1 INVX1_746 ( .A(_abc_15497_new_n5014_), .Y(_abc_15497_new_n5024_));
INVX1 INVX1_747 ( .A(c_reg_16_), .Y(_abc_15497_new_n5025_));
INVX1 INVX1_748 ( .A(_abc_15497_new_n5031_), .Y(_abc_15497_new_n5032_));
INVX1 INVX1_749 ( .A(_abc_15497_new_n5035_), .Y(_abc_15497_new_n5036_));
INVX1 INVX1_75 ( .A(_abc_15497_new_n1018_), .Y(_abc_15497_new_n1021_));
INVX1 INVX1_750 ( .A(w_16_), .Y(_abc_15497_new_n5037_));
INVX1 INVX1_751 ( .A(_abc_15497_new_n5039_), .Y(_abc_15497_new_n5040_));
INVX1 INVX1_752 ( .A(_abc_15497_new_n5041_), .Y(_abc_15497_new_n5042_));
INVX1 INVX1_753 ( .A(_abc_15497_new_n5045_), .Y(_abc_15497_new_n5046_));
INVX1 INVX1_754 ( .A(_abc_15497_new_n5051_), .Y(_abc_15497_new_n5052_));
INVX1 INVX1_755 ( .A(_abc_15497_new_n5055_), .Y(_abc_15497_new_n5056_));
INVX1 INVX1_756 ( .A(_abc_15497_new_n5057_), .Y(_abc_15497_new_n5059_));
INVX1 INVX1_757 ( .A(_abc_15497_new_n5063_), .Y(_abc_15497_new_n5064_));
INVX1 INVX1_758 ( .A(_abc_15497_new_n5065_), .Y(_abc_15497_new_n5066_));
INVX1 INVX1_759 ( .A(_abc_15497_new_n5068_), .Y(_abc_15497_new_n5069_));
INVX1 INVX1_76 ( .A(_abc_15497_new_n1030_), .Y(_abc_15497_new_n1031_));
INVX1 INVX1_760 ( .A(_abc_15497_new_n5076_), .Y(_abc_15497_new_n5077_));
INVX1 INVX1_761 ( .A(_abc_15497_new_n5058_), .Y(_abc_15497_new_n5078_));
INVX1 INVX1_762 ( .A(_abc_15497_new_n5079_), .Y(_abc_15497_new_n5080_));
INVX1 INVX1_763 ( .A(_abc_15497_new_n5047_), .Y(_abc_15497_new_n5081_));
INVX1 INVX1_764 ( .A(_abc_15497_new_n5084_), .Y(_abc_15497_new_n5085_));
INVX1 INVX1_765 ( .A(_abc_15497_new_n5088_), .Y(_abc_15497_new_n5089_));
INVX1 INVX1_766 ( .A(_abc_15497_new_n5091_), .Y(_abc_15497_new_n5092_));
INVX1 INVX1_767 ( .A(d_reg_17_), .Y(_abc_15497_new_n5093_));
INVX1 INVX1_768 ( .A(_abc_15497_new_n5083_), .Y(_abc_15497_new_n5097_));
INVX1 INVX1_769 ( .A(_abc_15497_new_n5102_), .Y(_abc_15497_new_n5103_));
INVX1 INVX1_77 ( .A(_abc_15497_new_n1032_), .Y(_abc_15497_new_n1033_));
INVX1 INVX1_770 ( .A(w_17_), .Y(_abc_15497_new_n5105_));
INVX1 INVX1_771 ( .A(_abc_15497_new_n5107_), .Y(_abc_15497_new_n5108_));
INVX1 INVX1_772 ( .A(_abc_15497_new_n5109_), .Y(_abc_15497_new_n5110_));
INVX1 INVX1_773 ( .A(_abc_15497_new_n5113_), .Y(_abc_15497_new_n5114_));
INVX1 INVX1_774 ( .A(_abc_15497_new_n5115_), .Y(_abc_15497_new_n5116_));
INVX1 INVX1_775 ( .A(_abc_15497_new_n5119_), .Y(_abc_15497_new_n5120_));
INVX1 INVX1_776 ( .A(_abc_15497_new_n5122_), .Y(_abc_15497_new_n5123_));
INVX1 INVX1_777 ( .A(_abc_15497_new_n5125_), .Y(_abc_15497_new_n5126_));
INVX1 INVX1_778 ( .A(_abc_15497_new_n5128_), .Y(_abc_15497_new_n5129_));
INVX1 INVX1_779 ( .A(_abc_15497_new_n5131_), .Y(_abc_15497_new_n5132_));
INVX1 INVX1_78 ( .A(_abc_15497_new_n1046_), .Y(_abc_15497_new_n1047_));
INVX1 INVX1_780 ( .A(_abc_15497_new_n5135_), .Y(_abc_15497_new_n5136_));
INVX1 INVX1_781 ( .A(_abc_15497_new_n5133_), .Y(_abc_15497_new_n5147_));
INVX1 INVX1_782 ( .A(_abc_15497_new_n5149_), .Y(_abc_15497_new_n5150_));
INVX1 INVX1_783 ( .A(_abc_15497_new_n5152_), .Y(_abc_15497_new_n5153_));
INVX1 INVX1_784 ( .A(_abc_15497_new_n5154_), .Y(_abc_15497_new_n5155_));
INVX1 INVX1_785 ( .A(_abc_15497_new_n5157_), .Y(_abc_15497_new_n5158_));
INVX1 INVX1_786 ( .A(_abc_15497_new_n5160_), .Y(_abc_15497_new_n5161_));
INVX1 INVX1_787 ( .A(_abc_15497_new_n5164_), .Y(_abc_15497_new_n5165_));
INVX1 INVX1_788 ( .A(_abc_15497_new_n5156_), .Y(_abc_15497_new_n5166_));
INVX1 INVX1_789 ( .A(c_reg_18_), .Y(_abc_15497_new_n5167_));
INVX1 INVX1_79 ( .A(_abc_15497_new_n1048_), .Y(_abc_15497_new_n1051_));
INVX1 INVX1_790 ( .A(_abc_15497_new_n5173_), .Y(_abc_15497_new_n5174_));
INVX1 INVX1_791 ( .A(w_18_), .Y(_abc_15497_new_n5178_));
INVX1 INVX1_792 ( .A(_abc_15497_new_n5180_), .Y(_abc_15497_new_n5181_));
INVX1 INVX1_793 ( .A(_abc_15497_new_n5182_), .Y(_abc_15497_new_n5183_));
INVX1 INVX1_794 ( .A(_abc_15497_new_n5186_), .Y(_abc_15497_new_n5187_));
INVX1 INVX1_795 ( .A(_abc_15497_new_n5188_), .Y(_abc_15497_new_n5189_));
INVX1 INVX1_796 ( .A(_abc_15497_new_n5191_), .Y(_abc_15497_new_n5192_));
INVX1 INVX1_797 ( .A(_abc_15497_new_n5176_), .Y(_abc_15497_new_n5194_));
INVX1 INVX1_798 ( .A(_abc_15497_new_n5196_), .Y(_abc_15497_new_n5197_));
INVX1 INVX1_799 ( .A(_abc_15497_new_n5200_), .Y(_abc_15497_new_n5201_));
INVX1 INVX1_8 ( .A(_abc_15497_new_n718_), .Y(_abc_15497_new_n719_));
INVX1 INVX1_80 ( .A(_abc_15497_new_n1057_), .Y(_abc_15497_new_n1058_));
INVX1 INVX1_800 ( .A(_abc_15497_new_n5204_), .Y(_abc_15497_new_n5205_));
INVX1 INVX1_801 ( .A(_abc_15497_new_n5207_), .Y(_abc_15497_new_n5208_));
INVX1 INVX1_802 ( .A(_abc_15497_new_n5202_), .Y(_abc_15497_new_n5215_));
INVX1 INVX1_803 ( .A(_abc_15497_new_n5217_), .Y(_abc_15497_new_n5218_));
INVX1 INVX1_804 ( .A(_abc_15497_new_n5220_), .Y(_abc_15497_new_n5221_));
INVX1 INVX1_805 ( .A(_abc_15497_new_n5223_), .Y(_abc_15497_new_n5224_));
INVX1 INVX1_806 ( .A(_abc_15497_new_n5227_), .Y(_abc_15497_new_n5228_));
INVX1 INVX1_807 ( .A(_abc_15497_new_n5219_), .Y(_abc_15497_new_n5229_));
INVX1 INVX1_808 ( .A(c_reg_19_), .Y(_abc_15497_new_n5230_));
INVX1 INVX1_809 ( .A(_abc_15497_new_n5236_), .Y(_abc_15497_new_n5237_));
INVX1 INVX1_81 ( .A(_abc_15497_new_n1059_), .Y(_abc_15497_new_n1060_));
INVX1 INVX1_810 ( .A(_abc_15497_new_n5239_), .Y(_abc_15497_new_n5240_));
INVX1 INVX1_811 ( .A(w_19_), .Y(_abc_15497_new_n5242_));
INVX1 INVX1_812 ( .A(_abc_15497_new_n5244_), .Y(_abc_15497_new_n5245_));
INVX1 INVX1_813 ( .A(_abc_15497_new_n5246_), .Y(_abc_15497_new_n5247_));
INVX1 INVX1_814 ( .A(_abc_15497_new_n5250_), .Y(_abc_15497_new_n5251_));
INVX1 INVX1_815 ( .A(_abc_15497_new_n5252_), .Y(_abc_15497_new_n5253_));
INVX1 INVX1_816 ( .A(_abc_15497_new_n5256_), .Y(_abc_15497_new_n5257_));
INVX1 INVX1_817 ( .A(_abc_15497_new_n5259_), .Y(_abc_15497_new_n5260_));
INVX1 INVX1_818 ( .A(_abc_15497_new_n5263_), .Y(_abc_15497_new_n5264_));
INVX1 INVX1_819 ( .A(_abc_15497_new_n5267_), .Y(_abc_15497_new_n5268_));
INVX1 INVX1_82 ( .A(_abc_15497_new_n1045_), .Y(_abc_15497_new_n1061_));
INVX1 INVX1_820 ( .A(_abc_15497_new_n5198_), .Y(_abc_15497_new_n5270_));
INVX1 INVX1_821 ( .A(_abc_15497_new_n5216_), .Y(_abc_15497_new_n5274_));
INVX1 INVX1_822 ( .A(_abc_15497_new_n5272_), .Y(_abc_15497_new_n5275_));
INVX1 INVX1_823 ( .A(_abc_15497_new_n5271_), .Y(_abc_15497_new_n5286_));
INVX1 INVX1_824 ( .A(_abc_15497_new_n5288_), .Y(_abc_15497_new_n5289_));
INVX1 INVX1_825 ( .A(_abc_15497_new_n5294_), .Y(_abc_15497_new_n5295_));
INVX1 INVX1_826 ( .A(_abc_15497_new_n5262_), .Y(_abc_15497_new_n5296_));
INVX1 INVX1_827 ( .A(_abc_15497_new_n5265_), .Y(_abc_15497_new_n5297_));
INVX1 INVX1_828 ( .A(_abc_15497_new_n5298_), .Y(_abc_15497_new_n5299_));
INVX1 INVX1_829 ( .A(_abc_15497_new_n5300_), .Y(_abc_15497_new_n5301_));
INVX1 INVX1_83 ( .A(_abc_15497_new_n1076_), .Y(_abc_15497_new_n1077_));
INVX1 INVX1_830 ( .A(_abc_15497_new_n5303_), .Y(_abc_15497_new_n5304_));
INVX1 INVX1_831 ( .A(_abc_15497_new_n5306_), .Y(_abc_15497_new_n5307_));
INVX1 INVX1_832 ( .A(_abc_15497_new_n5310_), .Y(_abc_15497_new_n5311_));
INVX1 INVX1_833 ( .A(_abc_15497_new_n5302_), .Y(_abc_15497_new_n5312_));
INVX1 INVX1_834 ( .A(c_reg_20_), .Y(_abc_15497_new_n5313_));
INVX1 INVX1_835 ( .A(_abc_15497_new_n5319_), .Y(_abc_15497_new_n5320_));
INVX1 INVX1_836 ( .A(_abc_15497_new_n5322_), .Y(_abc_15497_new_n5323_));
INVX1 INVX1_837 ( .A(w_20_), .Y(_abc_15497_new_n5325_));
INVX1 INVX1_838 ( .A(_abc_15497_new_n5327_), .Y(_abc_15497_new_n5328_));
INVX1 INVX1_839 ( .A(_abc_15497_new_n5329_), .Y(_abc_15497_new_n5330_));
INVX1 INVX1_84 ( .A(_abc_15497_new_n1078_), .Y(_abc_15497_new_n1081_));
INVX1 INVX1_840 ( .A(_abc_15497_new_n5333_), .Y(_abc_15497_new_n5334_));
INVX1 INVX1_841 ( .A(_abc_15497_new_n5335_), .Y(_abc_15497_new_n5336_));
INVX1 INVX1_842 ( .A(_abc_15497_new_n5339_), .Y(_abc_15497_new_n5340_));
INVX1 INVX1_843 ( .A(_abc_15497_new_n5342_), .Y(_abc_15497_new_n5343_));
INVX1 INVX1_844 ( .A(_abc_15497_new_n5347_), .Y(_abc_15497_new_n5348_));
INVX1 INVX1_845 ( .A(_abc_15497_new_n5350_), .Y(_abc_15497_new_n5351_));
INVX1 INVX1_846 ( .A(_abc_15497_new_n5354_), .Y(_abc_15497_new_n5355_));
INVX1 INVX1_847 ( .A(_abc_15497_new_n5352_), .Y(_abc_15497_new_n5365_));
INVX1 INVX1_848 ( .A(_abc_15497_new_n5366_), .Y(_abc_15497_new_n5367_));
INVX1 INVX1_849 ( .A(_abc_15497_new_n5369_), .Y(_abc_15497_new_n5370_));
INVX1 INVX1_85 ( .A(_abc_15497_new_n1091_), .Y(_abc_15497_new_n1092_));
INVX1 INVX1_850 ( .A(_abc_15497_new_n5372_), .Y(_abc_15497_new_n5373_));
INVX1 INVX1_851 ( .A(_abc_15497_new_n5375_), .Y(_abc_15497_new_n5376_));
INVX1 INVX1_852 ( .A(_abc_15497_new_n5379_), .Y(_abc_15497_new_n5380_));
INVX1 INVX1_853 ( .A(_abc_15497_new_n5371_), .Y(_abc_15497_new_n5381_));
INVX1 INVX1_854 ( .A(c_reg_21_), .Y(_abc_15497_new_n5382_));
INVX1 INVX1_855 ( .A(_abc_15497_new_n5388_), .Y(_abc_15497_new_n5389_));
INVX1 INVX1_856 ( .A(_abc_15497_new_n5391_), .Y(_abc_15497_new_n5392_));
INVX1 INVX1_857 ( .A(w_21_), .Y(_abc_15497_new_n5394_));
INVX1 INVX1_858 ( .A(_abc_15497_new_n5396_), .Y(_abc_15497_new_n5397_));
INVX1 INVX1_859 ( .A(_abc_15497_new_n5398_), .Y(_abc_15497_new_n5399_));
INVX1 INVX1_86 ( .A(_abc_15497_new_n1093_), .Y(_abc_15497_new_n1096_));
INVX1 INVX1_860 ( .A(_abc_15497_new_n5402_), .Y(_abc_15497_new_n5403_));
INVX1 INVX1_861 ( .A(_abc_15497_new_n5404_), .Y(_abc_15497_new_n5405_));
INVX1 INVX1_862 ( .A(_abc_15497_new_n5408_), .Y(_abc_15497_new_n5409_));
INVX1 INVX1_863 ( .A(_abc_15497_new_n5411_), .Y(_abc_15497_new_n5412_));
INVX1 INVX1_864 ( .A(_abc_15497_new_n5415_), .Y(_abc_15497_new_n5416_));
INVX1 INVX1_865 ( .A(_abc_15497_new_n5419_), .Y(_abc_15497_new_n5420_));
INVX1 INVX1_866 ( .A(_abc_15497_new_n5368_), .Y(_abc_15497_new_n5422_));
INVX1 INVX1_867 ( .A(_abc_15497_new_n5424_), .Y(_abc_15497_new_n5425_));
INVX1 INVX1_868 ( .A(_abc_15497_new_n5421_), .Y(_abc_15497_new_n5437_));
INVX1 INVX1_869 ( .A(_abc_15497_new_n5440_), .Y(_abc_15497_new_n5441_));
INVX1 INVX1_87 ( .A(_abc_15497_new_n1107_), .Y(_abc_15497_new_n1108_));
INVX1 INVX1_870 ( .A(_abc_15497_new_n5414_), .Y(_abc_15497_new_n5442_));
INVX1 INVX1_871 ( .A(_abc_15497_new_n5417_), .Y(_abc_15497_new_n5443_));
INVX1 INVX1_872 ( .A(_abc_15497_new_n5444_), .Y(_abc_15497_new_n5445_));
INVX1 INVX1_873 ( .A(_abc_15497_new_n5448_), .Y(_abc_15497_new_n5449_));
INVX1 INVX1_874 ( .A(_abc_15497_new_n5451_), .Y(_abc_15497_new_n5452_));
INVX1 INVX1_875 ( .A(_abc_15497_new_n5455_), .Y(_abc_15497_new_n5456_));
INVX1 INVX1_876 ( .A(_abc_15497_new_n5447_), .Y(_abc_15497_new_n5457_));
INVX1 INVX1_877 ( .A(c_reg_22_), .Y(_abc_15497_new_n5458_));
INVX1 INVX1_878 ( .A(_abc_15497_new_n5464_), .Y(_abc_15497_new_n5465_));
INVX1 INVX1_879 ( .A(_abc_15497_new_n5467_), .Y(_abc_15497_new_n5468_));
INVX1 INVX1_88 ( .A(_abc_15497_new_n1109_), .Y(_abc_15497_new_n1113_));
INVX1 INVX1_880 ( .A(w_22_), .Y(_abc_15497_new_n5470_));
INVX1 INVX1_881 ( .A(_abc_15497_new_n5472_), .Y(_abc_15497_new_n5473_));
INVX1 INVX1_882 ( .A(_abc_15497_new_n5474_), .Y(_abc_15497_new_n5475_));
INVX1 INVX1_883 ( .A(_abc_15497_new_n5478_), .Y(_abc_15497_new_n5479_));
INVX1 INVX1_884 ( .A(_abc_15497_new_n5480_), .Y(_abc_15497_new_n5481_));
INVX1 INVX1_885 ( .A(_abc_15497_new_n5484_), .Y(_abc_15497_new_n5485_));
INVX1 INVX1_886 ( .A(_abc_15497_new_n5487_), .Y(_abc_15497_new_n5488_));
INVX1 INVX1_887 ( .A(_abc_15497_new_n5490_), .Y(_abc_15497_new_n5491_));
INVX1 INVX1_888 ( .A(_abc_15497_new_n5492_), .Y(_abc_15497_new_n5493_));
INVX1 INVX1_889 ( .A(_abc_15497_new_n5496_), .Y(_abc_15497_new_n5497_));
INVX1 INVX1_89 ( .A(_abc_15497_new_n1119_), .Y(_abc_15497_new_n1120_));
INVX1 INVX1_890 ( .A(_abc_15497_new_n5500_), .Y(_abc_15497_new_n5501_));
INVX1 INVX1_891 ( .A(_abc_15497_new_n5498_), .Y(_abc_15497_new_n5510_));
INVX1 INVX1_892 ( .A(_abc_15497_new_n5511_), .Y(_abc_15497_new_n5512_));
INVX1 INVX1_893 ( .A(_abc_15497_new_n5516_), .Y(_abc_15497_new_n5517_));
INVX1 INVX1_894 ( .A(_abc_15497_new_n5520_), .Y(_abc_15497_new_n5521_));
INVX1 INVX1_895 ( .A(_abc_15497_new_n5523_), .Y(_abc_15497_new_n5524_));
INVX1 INVX1_896 ( .A(d_reg_23_), .Y(_abc_15497_new_n5525_));
INVX1 INVX1_897 ( .A(_abc_15497_new_n5515_), .Y(_abc_15497_new_n5529_));
INVX1 INVX1_898 ( .A(_abc_15497_new_n5534_), .Y(_abc_15497_new_n5535_));
INVX1 INVX1_899 ( .A(w_23_), .Y(_abc_15497_new_n5537_));
INVX1 INVX1_9 ( .A(_abc_15497_new_n724_), .Y(_abc_15497_new_n725_));
INVX1 INVX1_90 ( .A(_abc_15497_new_n1125_), .Y(_abc_15497_new_n1126_));
INVX1 INVX1_900 ( .A(_abc_15497_new_n5539_), .Y(_abc_15497_new_n5540_));
INVX1 INVX1_901 ( .A(_abc_15497_new_n5541_), .Y(_abc_15497_new_n5542_));
INVX1 INVX1_902 ( .A(_abc_15497_new_n5545_), .Y(_abc_15497_new_n5546_));
INVX1 INVX1_903 ( .A(_abc_15497_new_n5547_), .Y(_abc_15497_new_n5548_));
INVX1 INVX1_904 ( .A(_abc_15497_new_n5551_), .Y(_abc_15497_new_n5552_));
INVX1 INVX1_905 ( .A(_abc_15497_new_n5554_), .Y(_abc_15497_new_n5555_));
INVX1 INVX1_906 ( .A(_abc_15497_new_n5556_), .Y(_abc_15497_new_n5557_));
INVX1 INVX1_907 ( .A(_abc_15497_new_n5560_), .Y(_abc_15497_new_n5561_));
INVX1 INVX1_908 ( .A(_abc_15497_new_n5513_), .Y(_abc_15497_new_n5565_));
INVX1 INVX1_909 ( .A(_abc_15497_new_n5563_), .Y(_abc_15497_new_n5566_));
INVX1 INVX1_91 ( .A(_abc_15497_new_n1134_), .Y(_abc_15497_new_n1135_));
INVX1 INVX1_910 ( .A(_abc_15497_new_n5568_), .Y(_abc_15497_new_n5569_));
INVX1 INVX1_911 ( .A(_abc_15497_new_n5564_), .Y(_abc_15497_new_n5583_));
INVX1 INVX1_912 ( .A(_abc_15497_new_n5590_), .Y(_abc_15497_new_n5591_));
INVX1 INVX1_913 ( .A(_abc_15497_new_n5592_), .Y(_abc_15497_new_n5593_));
INVX1 INVX1_914 ( .A(_abc_15497_new_n5596_), .Y(_abc_15497_new_n5597_));
INVX1 INVX1_915 ( .A(_abc_15497_new_n5600_), .Y(_abc_15497_new_n5601_));
INVX1 INVX1_916 ( .A(_abc_15497_new_n5603_), .Y(_abc_15497_new_n5604_));
INVX1 INVX1_917 ( .A(d_reg_24_), .Y(_abc_15497_new_n5605_));
INVX1 INVX1_918 ( .A(_abc_15497_new_n5595_), .Y(_abc_15497_new_n5609_));
INVX1 INVX1_919 ( .A(_abc_15497_new_n5614_), .Y(_abc_15497_new_n5615_));
INVX1 INVX1_92 ( .A(_abc_15497_new_n1138_), .Y(_abc_15497_new_n1139_));
INVX1 INVX1_920 ( .A(w_24_), .Y(_abc_15497_new_n5617_));
INVX1 INVX1_921 ( .A(_abc_15497_new_n5619_), .Y(_abc_15497_new_n5620_));
INVX1 INVX1_922 ( .A(_abc_15497_new_n5621_), .Y(_abc_15497_new_n5622_));
INVX1 INVX1_923 ( .A(_abc_15497_new_n5625_), .Y(_abc_15497_new_n5626_));
INVX1 INVX1_924 ( .A(_abc_15497_new_n5627_), .Y(_abc_15497_new_n5628_));
INVX1 INVX1_925 ( .A(_abc_15497_new_n5631_), .Y(_abc_15497_new_n5632_));
INVX1 INVX1_926 ( .A(_abc_15497_new_n5634_), .Y(_abc_15497_new_n5635_));
INVX1 INVX1_927 ( .A(_abc_15497_new_n5637_), .Y(_abc_15497_new_n5638_));
INVX1 INVX1_928 ( .A(_abc_15497_new_n5639_), .Y(_abc_15497_new_n5640_));
INVX1 INVX1_929 ( .A(_abc_15497_new_n5643_), .Y(_abc_15497_new_n5644_));
INVX1 INVX1_93 ( .A(_abc_15497_new_n1142_), .Y(_abc_15497_new_n1143_));
INVX1 INVX1_930 ( .A(_abc_15497_new_n5647_), .Y(_abc_15497_new_n5648_));
INVX1 INVX1_931 ( .A(_abc_15497_new_n5650_), .Y(_abc_15497_new_n5651_));
INVX1 INVX1_932 ( .A(_abc_15497_new_n5645_), .Y(_abc_15497_new_n5658_));
INVX1 INVX1_933 ( .A(_abc_15497_new_n5660_), .Y(_abc_15497_new_n5661_));
INVX1 INVX1_934 ( .A(_abc_15497_new_n5664_), .Y(_abc_15497_new_n5665_));
INVX1 INVX1_935 ( .A(_abc_15497_new_n5668_), .Y(_abc_15497_new_n5669_));
INVX1 INVX1_936 ( .A(_abc_15497_new_n5671_), .Y(_abc_15497_new_n5672_));
INVX1 INVX1_937 ( .A(d_reg_25_), .Y(_abc_15497_new_n5673_));
INVX1 INVX1_938 ( .A(_abc_15497_new_n5663_), .Y(_abc_15497_new_n5677_));
INVX1 INVX1_939 ( .A(_abc_15497_new_n5682_), .Y(_abc_15497_new_n5683_));
INVX1 INVX1_94 ( .A(_abc_15497_new_n1150_), .Y(_abc_15497_new_n1151_));
INVX1 INVX1_940 ( .A(w_25_), .Y(_abc_15497_new_n5685_));
INVX1 INVX1_941 ( .A(_abc_15497_new_n5687_), .Y(_abc_15497_new_n5688_));
INVX1 INVX1_942 ( .A(_abc_15497_new_n5689_), .Y(_abc_15497_new_n5690_));
INVX1 INVX1_943 ( .A(_abc_15497_new_n5693_), .Y(_abc_15497_new_n5694_));
INVX1 INVX1_944 ( .A(_abc_15497_new_n5695_), .Y(_abc_15497_new_n5696_));
INVX1 INVX1_945 ( .A(_abc_15497_new_n5699_), .Y(_abc_15497_new_n5700_));
INVX1 INVX1_946 ( .A(_abc_15497_new_n5702_), .Y(_abc_15497_new_n5703_));
INVX1 INVX1_947 ( .A(_abc_15497_new_n5704_), .Y(_abc_15497_new_n5705_));
INVX1 INVX1_948 ( .A(_abc_15497_new_n5709_), .Y(_abc_15497_new_n5710_));
INVX1 INVX1_949 ( .A(_abc_15497_new_n5659_), .Y(_abc_15497_new_n5713_));
INVX1 INVX1_95 ( .A(_abc_15497_new_n1153_), .Y(_abc_15497_new_n1154_));
INVX1 INVX1_950 ( .A(_abc_15497_new_n5711_), .Y(_abc_15497_new_n5714_));
INVX1 INVX1_951 ( .A(_abc_15497_new_n5724_), .Y(_abc_15497_new_n5725_));
INVX1 INVX1_952 ( .A(_abc_15497_new_n5726_), .Y(_abc_15497_new_n5727_));
INVX1 INVX1_953 ( .A(_abc_15497_new_n5728_), .Y(_abc_15497_new_n5729_));
INVX1 INVX1_954 ( .A(_abc_15497_new_n5731_), .Y(_abc_15497_new_n5732_));
INVX1 INVX1_955 ( .A(_abc_15497_new_n5735_), .Y(_abc_15497_new_n5736_));
INVX1 INVX1_956 ( .A(_abc_15497_new_n5739_), .Y(_abc_15497_new_n5740_));
INVX1 INVX1_957 ( .A(d_reg_26_), .Y(_abc_15497_new_n5741_));
INVX1 INVX1_958 ( .A(_abc_15497_new_n5745_), .Y(_abc_15497_new_n5746_));
INVX1 INVX1_959 ( .A(_abc_15497_new_n5748_), .Y(_abc_15497_new_n5749_));
INVX1 INVX1_96 ( .A(_abc_15497_new_n1157_), .Y(_abc_15497_new_n1158_));
INVX1 INVX1_960 ( .A(_abc_15497_new_n5751_), .Y(_abc_15497_new_n5752_));
INVX1 INVX1_961 ( .A(w_26_), .Y(_abc_15497_new_n5754_));
INVX1 INVX1_962 ( .A(_abc_15497_new_n5756_), .Y(_abc_15497_new_n5757_));
INVX1 INVX1_963 ( .A(_abc_15497_new_n5758_), .Y(_abc_15497_new_n5759_));
INVX1 INVX1_964 ( .A(_abc_15497_new_n5762_), .Y(_abc_15497_new_n5763_));
INVX1 INVX1_965 ( .A(_abc_15497_new_n5764_), .Y(_abc_15497_new_n5765_));
INVX1 INVX1_966 ( .A(_abc_15497_new_n5768_), .Y(_abc_15497_new_n5769_));
INVX1 INVX1_967 ( .A(_abc_15497_new_n5771_), .Y(_abc_15497_new_n5772_));
INVX1 INVX1_968 ( .A(_abc_15497_new_n5774_), .Y(_abc_15497_new_n5775_));
INVX1 INVX1_969 ( .A(_abc_15497_new_n5776_), .Y(_abc_15497_new_n5777_));
INVX1 INVX1_97 ( .A(_abc_15497_new_n1163_), .Y(_abc_15497_new_n1164_));
INVX1 INVX1_970 ( .A(_abc_15497_new_n5780_), .Y(_abc_15497_new_n5781_));
INVX1 INVX1_971 ( .A(_abc_15497_new_n5784_), .Y(_abc_15497_new_n5785_));
INVX1 INVX1_972 ( .A(_abc_15497_new_n5787_), .Y(_abc_15497_new_n5788_));
INVX1 INVX1_973 ( .A(_abc_15497_new_n5795_), .Y(_abc_15497_new_n5796_));
INVX1 INVX1_974 ( .A(_abc_15497_new_n5797_), .Y(_abc_15497_new_n5798_));
INVX1 INVX1_975 ( .A(_abc_15497_new_n5800_), .Y(_abc_15497_new_n5801_));
INVX1 INVX1_976 ( .A(_abc_15497_new_n5804_), .Y(_abc_15497_new_n5805_));
INVX1 INVX1_977 ( .A(_abc_15497_new_n5808_), .Y(_abc_15497_new_n5809_));
INVX1 INVX1_978 ( .A(d_reg_27_), .Y(_abc_15497_new_n5810_));
INVX1 INVX1_979 ( .A(_abc_15497_new_n5814_), .Y(_abc_15497_new_n5815_));
INVX1 INVX1_98 ( .A(_abc_15497_new_n1166_), .Y(_abc_15497_new_n1167_));
INVX1 INVX1_980 ( .A(_abc_15497_new_n5817_), .Y(_abc_15497_new_n5818_));
INVX1 INVX1_981 ( .A(_abc_15497_new_n5820_), .Y(_abc_15497_new_n5821_));
INVX1 INVX1_982 ( .A(w_27_), .Y(_abc_15497_new_n5823_));
INVX1 INVX1_983 ( .A(_abc_15497_new_n5825_), .Y(_abc_15497_new_n5826_));
INVX1 INVX1_984 ( .A(_abc_15497_new_n5827_), .Y(_abc_15497_new_n5828_));
INVX1 INVX1_985 ( .A(_abc_15497_new_n5831_), .Y(_abc_15497_new_n5832_));
INVX1 INVX1_986 ( .A(_abc_15497_new_n5833_), .Y(_abc_15497_new_n5834_));
INVX1 INVX1_987 ( .A(_abc_15497_new_n5837_), .Y(_abc_15497_new_n5838_));
INVX1 INVX1_988 ( .A(_abc_15497_new_n5840_), .Y(_abc_15497_new_n5841_));
INVX1 INVX1_989 ( .A(_abc_15497_new_n5842_), .Y(_abc_15497_new_n5843_));
INVX1 INVX1_99 ( .A(_abc_15497_new_n1168_), .Y(_abc_15497_new_n1170_));
INVX1 INVX1_990 ( .A(_abc_15497_new_n5847_), .Y(_abc_15497_new_n5848_));
INVX1 INVX1_991 ( .A(_abc_15497_new_n5849_), .Y(_abc_15497_new_n5851_));
INVX1 INVX1_992 ( .A(_abc_15497_new_n5861_), .Y(_abc_15497_new_n5862_));
INVX1 INVX1_993 ( .A(_abc_15497_new_n5860_), .Y(_abc_15497_new_n5864_));
INVX1 INVX1_994 ( .A(_abc_15497_new_n5867_), .Y(_abc_15497_new_n5868_));
INVX1 INVX1_995 ( .A(_abc_15497_new_n5870_), .Y(_abc_15497_new_n5871_));
INVX1 INVX1_996 ( .A(_abc_15497_new_n5873_), .Y(_abc_15497_new_n5874_));
INVX1 INVX1_997 ( .A(_abc_15497_new_n5877_), .Y(_abc_15497_new_n5878_));
INVX1 INVX1_998 ( .A(_abc_15497_new_n5881_), .Y(_abc_15497_new_n5882_));
INVX1 INVX1_999 ( .A(d_reg_28_), .Y(_abc_15497_new_n5883_));
OR2X2 OR2X2_1 ( .A(c_reg_23_), .B(\digest[87] ), .Y(_abc_15497_new_n703_));
OR2X2 OR2X2_10 ( .A(c_reg_17_), .B(\digest[81] ), .Y(_abc_15497_new_n742_));
OR2X2 OR2X2_100 ( .A(_abc_15497_new_n1022_), .B(_abc_15497_new_n1009_), .Y(_abc_15497_new_n1023_));
OR2X2 OR2X2_1000 ( .A(_abc_15497_new_n3683_), .B(_abc_15497_new_n3684_), .Y(_abc_15497_new_n3685_));
OR2X2 OR2X2_1001 ( .A(_abc_15497_new_n3685_), .B(_abc_15497_new_n3681_), .Y(_0c_reg_31_0__22_));
OR2X2 OR2X2_1002 ( .A(_abc_15497_new_n699_), .B(\digest[87] ), .Y(_abc_15497_new_n3688_));
OR2X2 OR2X2_1003 ( .A(_abc_15497_new_n3689_), .B(_abc_15497_new_n3690_), .Y(_abc_15497_new_n3691_));
OR2X2 OR2X2_1004 ( .A(_abc_15497_new_n3691_), .B(_abc_15497_new_n3687_), .Y(_0c_reg_31_0__23_));
OR2X2 OR2X2_1005 ( .A(_abc_15497_new_n3695_), .B(_abc_15497_new_n3696_), .Y(_abc_15497_new_n3697_));
OR2X2 OR2X2_1006 ( .A(_abc_15497_new_n3697_), .B(_abc_15497_new_n3693_), .Y(_0c_reg_31_0__24_));
OR2X2 OR2X2_1007 ( .A(_abc_15497_new_n3701_), .B(_abc_15497_new_n3702_), .Y(_abc_15497_new_n3703_));
OR2X2 OR2X2_1008 ( .A(_abc_15497_new_n3703_), .B(_abc_15497_new_n3699_), .Y(_0c_reg_31_0__25_));
OR2X2 OR2X2_1009 ( .A(_abc_15497_new_n3707_), .B(_abc_15497_new_n3708_), .Y(_abc_15497_new_n3709_));
OR2X2 OR2X2_101 ( .A(_abc_15497_new_n1025_), .B(_abc_15497_new_n1026_), .Y(_0H4_reg_31_0__1_));
OR2X2 OR2X2_1010 ( .A(_abc_15497_new_n3709_), .B(_abc_15497_new_n3705_), .Y(_0c_reg_31_0__26_));
OR2X2 OR2X2_1011 ( .A(_abc_15497_new_n3712_), .B(_abc_15497_new_n3713_), .Y(_abc_15497_new_n3714_));
OR2X2 OR2X2_1012 ( .A(_abc_15497_new_n3714_), .B(_abc_15497_new_n3711_), .Y(_0c_reg_31_0__27_));
OR2X2 OR2X2_1013 ( .A(_abc_15497_new_n3717_), .B(_abc_15497_new_n3718_), .Y(_abc_15497_new_n3719_));
OR2X2 OR2X2_1014 ( .A(_abc_15497_new_n3719_), .B(_abc_15497_new_n3716_), .Y(_0c_reg_31_0__28_));
OR2X2 OR2X2_1015 ( .A(_abc_15497_new_n3723_), .B(_abc_15497_new_n3724_), .Y(_abc_15497_new_n3725_));
OR2X2 OR2X2_1016 ( .A(_abc_15497_new_n3725_), .B(_abc_15497_new_n3721_), .Y(_0c_reg_31_0__29_));
OR2X2 OR2X2_1017 ( .A(_abc_15497_new_n3729_), .B(_abc_15497_new_n3730_), .Y(_abc_15497_new_n3731_));
OR2X2 OR2X2_1018 ( .A(_abc_15497_new_n3731_), .B(_abc_15497_new_n3727_), .Y(_0c_reg_31_0__30_));
OR2X2 OR2X2_1019 ( .A(_abc_15497_new_n3734_), .B(_abc_15497_new_n3735_), .Y(_abc_15497_new_n3736_));
OR2X2 OR2X2_102 ( .A(e_reg_2_), .B(\digest[2] ), .Y(_abc_15497_new_n1029_));
OR2X2 OR2X2_1020 ( .A(_abc_15497_new_n3736_), .B(_abc_15497_new_n3733_), .Y(_0c_reg_31_0__31_));
OR2X2 OR2X2_1021 ( .A(_abc_15497_new_n3751_), .B(_abc_15497_new_n3747_), .Y(_abc_15497_new_n3752_));
OR2X2 OR2X2_1022 ( .A(_abc_15497_new_n3759_), .B(_abc_15497_new_n3755_), .Y(_abc_15497_new_n3760_));
OR2X2 OR2X2_1023 ( .A(b_reg_0_), .B(c_reg_0_), .Y(_abc_15497_new_n3762_));
OR2X2 OR2X2_1024 ( .A(_abc_15497_new_n3765_), .B(_abc_15497_new_n3766_), .Y(_abc_15497_new_n3767_));
OR2X2 OR2X2_1025 ( .A(_abc_15497_new_n3741_), .B(round_ctr_reg_6_), .Y(_abc_15497_new_n3768_));
OR2X2 OR2X2_1026 ( .A(_abc_15497_new_n3768_), .B(_abc_15497_new_n3738_), .Y(_abc_15497_new_n3769_));
OR2X2 OR2X2_1027 ( .A(_abc_15497_new_n3753_), .B(_abc_15497_new_n3774_), .Y(_abc_15497_new_n3775_));
OR2X2 OR2X2_1028 ( .A(_abc_15497_new_n3775_), .B(_abc_15497_new_n3767_), .Y(_abc_15497_new_n3776_));
OR2X2 OR2X2_1029 ( .A(round_ctr_reg_3_), .B(round_ctr_reg_2_), .Y(_abc_15497_new_n3777_));
OR2X2 OR2X2_103 ( .A(_abc_15497_new_n1028_), .B(_abc_15497_new_n1033_), .Y(_abc_15497_new_n1034_));
OR2X2 OR2X2_1030 ( .A(_abc_15497_new_n3778_), .B(round_ctr_reg_5_), .Y(_abc_15497_new_n3779_));
OR2X2 OR2X2_1031 ( .A(_abc_15497_new_n3779_), .B(round_ctr_reg_6_), .Y(_abc_15497_new_n3780_));
OR2X2 OR2X2_1032 ( .A(_abc_15497_new_n3759_), .B(_abc_15497_new_n3781_), .Y(_abc_15497_new_n3782_));
OR2X2 OR2X2_1033 ( .A(_abc_15497_new_n3771_), .B(round_ctr_reg_6_), .Y(_abc_15497_new_n3783_));
OR2X2 OR2X2_1034 ( .A(_abc_15497_new_n3744_), .B(_abc_15497_new_n3783_), .Y(_abc_15497_new_n3784_));
OR2X2 OR2X2_1035 ( .A(_abc_15497_new_n3784_), .B(_abc_15497_new_n3782_), .Y(_abc_15497_new_n3785_));
OR2X2 OR2X2_1036 ( .A(_abc_15497_new_n3787_), .B(_abc_15497_new_n3761_), .Y(_abc_15497_new_n3788_));
OR2X2 OR2X2_1037 ( .A(e_reg_0_), .B(a_reg_27_), .Y(_abc_15497_new_n3789_));
OR2X2 OR2X2_1038 ( .A(_abc_15497_new_n3796_), .B(_abc_15497_new_n3793_), .Y(_abc_15497_new_n3797_));
OR2X2 OR2X2_1039 ( .A(_abc_15497_new_n3806_), .B(_abc_15497_new_n3753_), .Y(_abc_15497_new_n3807_));
OR2X2 OR2X2_104 ( .A(_abc_15497_new_n1035_), .B(_abc_15497_new_n1018_), .Y(_abc_15497_new_n1036_));
OR2X2 OR2X2_1040 ( .A(_abc_15497_new_n3804_), .B(_abc_15497_new_n3807_), .Y(_abc_15497_new_n3808_));
OR2X2 OR2X2_1041 ( .A(_abc_15497_new_n3798_), .B(_abc_15497_new_n3811_), .Y(_abc_15497_new_n3812_));
OR2X2 OR2X2_1042 ( .A(_abc_15497_new_n3813_), .B(_abc_15497_new_n3744_), .Y(_abc_15497_new_n3814_));
OR2X2 OR2X2_1043 ( .A(_abc_15497_new_n3819_), .B(_abc_15497_new_n3820_), .Y(_abc_15497_new_n3821_));
OR2X2 OR2X2_1044 ( .A(_abc_15497_new_n3818_), .B(_abc_15497_new_n3821_), .Y(_0a_reg_31_0__0_));
OR2X2 OR2X2_1045 ( .A(_abc_15497_new_n3788_), .B(_abc_15497_new_n3797_), .Y(_abc_15497_new_n3823_));
OR2X2 OR2X2_1046 ( .A(b_reg_1_), .B(c_reg_1_), .Y(_abc_15497_new_n3824_));
OR2X2 OR2X2_1047 ( .A(_abc_15497_new_n3827_), .B(d_reg_1_), .Y(_abc_15497_new_n3828_));
OR2X2 OR2X2_1048 ( .A(_abc_15497_new_n3829_), .B(_abc_15497_new_n3830_), .Y(_abc_15497_new_n3831_));
OR2X2 OR2X2_1049 ( .A(_abc_15497_new_n3775_), .B(_abc_15497_new_n3831_), .Y(_abc_15497_new_n3832_));
OR2X2 OR2X2_105 ( .A(_abc_15497_new_n1036_), .B(_abc_15497_new_n1032_), .Y(_abc_15497_new_n1037_));
OR2X2 OR2X2_1050 ( .A(_abc_15497_new_n3833_), .B(b_reg_1_), .Y(_abc_15497_new_n3834_));
OR2X2 OR2X2_1051 ( .A(_abc_15497_new_n3780_), .B(_abc_15497_new_n3835_), .Y(_abc_15497_new_n3836_));
OR2X2 OR2X2_1052 ( .A(_abc_15497_new_n3838_), .B(_abc_15497_new_n3837_), .Y(_abc_15497_new_n3839_));
OR2X2 OR2X2_1053 ( .A(_abc_15497_new_n3784_), .B(_abc_15497_new_n3839_), .Y(_abc_15497_new_n3840_));
OR2X2 OR2X2_1054 ( .A(_abc_15497_new_n3793_), .B(_abc_15497_new_n3790_), .Y(_abc_15497_new_n3843_));
OR2X2 OR2X2_1055 ( .A(e_reg_1_), .B(a_reg_28_), .Y(_abc_15497_new_n3844_));
OR2X2 OR2X2_1056 ( .A(_abc_15497_new_n3847_), .B(w_1_), .Y(_abc_15497_new_n3848_));
OR2X2 OR2X2_1057 ( .A(_abc_15497_new_n3851_), .B(_abc_15497_new_n3843_), .Y(_abc_15497_new_n3854_));
OR2X2 OR2X2_1058 ( .A(_abc_15497_new_n3842_), .B(_abc_15497_new_n3855_), .Y(_abc_15497_new_n3856_));
OR2X2 OR2X2_1059 ( .A(_abc_15497_new_n3861_), .B(_abc_15497_new_n3863_), .Y(_abc_15497_new_n3864_));
OR2X2 OR2X2_106 ( .A(_abc_15497_new_n1039_), .B(_abc_15497_new_n1040_), .Y(_0H4_reg_31_0__2_));
OR2X2 OR2X2_1060 ( .A(_abc_15497_new_n3864_), .B(_abc_15497_new_n3859_), .Y(_abc_15497_new_n3865_));
OR2X2 OR2X2_1061 ( .A(_abc_15497_new_n3867_), .B(_abc_15497_new_n3849_), .Y(_abc_15497_new_n3868_));
OR2X2 OR2X2_1062 ( .A(_abc_15497_new_n3869_), .B(_abc_15497_new_n3852_), .Y(_abc_15497_new_n3870_));
OR2X2 OR2X2_1063 ( .A(_abc_15497_new_n3865_), .B(_abc_15497_new_n3870_), .Y(_abc_15497_new_n3871_));
OR2X2 OR2X2_1064 ( .A(_abc_15497_new_n3823_), .B(_abc_15497_new_n3872_), .Y(_abc_15497_new_n3873_));
OR2X2 OR2X2_1065 ( .A(_abc_15497_new_n3842_), .B(_abc_15497_new_n3870_), .Y(_abc_15497_new_n3874_));
OR2X2 OR2X2_1066 ( .A(_abc_15497_new_n3865_), .B(_abc_15497_new_n3855_), .Y(_abc_15497_new_n3875_));
OR2X2 OR2X2_1067 ( .A(_abc_15497_new_n3876_), .B(_abc_15497_new_n3811_), .Y(_abc_15497_new_n3877_));
OR2X2 OR2X2_1068 ( .A(_abc_15497_new_n3881_), .B(_abc_15497_new_n3880_), .Y(_abc_15497_new_n3882_));
OR2X2 OR2X2_1069 ( .A(_abc_15497_new_n3879_), .B(_abc_15497_new_n3883_), .Y(_abc_15497_new_n3884_));
OR2X2 OR2X2_107 ( .A(_abc_15497_new_n1043_), .B(_abc_15497_new_n1030_), .Y(_abc_15497_new_n1044_));
OR2X2 OR2X2_1070 ( .A(_abc_15497_new_n3885_), .B(_abc_15497_new_n3815_), .Y(_abc_15497_new_n3886_));
OR2X2 OR2X2_1071 ( .A(_abc_15497_new_n3884_), .B(_abc_15497_new_n3816_), .Y(_abc_15497_new_n3887_));
OR2X2 OR2X2_1072 ( .A(_abc_15497_new_n3890_), .B(_abc_15497_new_n3892_), .Y(_abc_15497_new_n3893_));
OR2X2 OR2X2_1073 ( .A(_abc_15497_new_n3889_), .B(_abc_15497_new_n3893_), .Y(_0a_reg_31_0__1_));
OR2X2 OR2X2_1074 ( .A(_abc_15497_new_n3882_), .B(_abc_15497_new_n3773_), .Y(_abc_15497_new_n3896_));
OR2X2 OR2X2_1075 ( .A(_abc_15497_new_n3898_), .B(_abc_15497_new_n3852_), .Y(_abc_15497_new_n3899_));
OR2X2 OR2X2_1076 ( .A(b_reg_2_), .B(c_reg_2_), .Y(_abc_15497_new_n3900_));
OR2X2 OR2X2_1077 ( .A(_abc_15497_new_n3903_), .B(d_reg_2_), .Y(_abc_15497_new_n3904_));
OR2X2 OR2X2_1078 ( .A(_abc_15497_new_n3775_), .B(_abc_15497_new_n3908_), .Y(_abc_15497_new_n3909_));
OR2X2 OR2X2_1079 ( .A(_abc_15497_new_n3910_), .B(b_reg_2_), .Y(_abc_15497_new_n3911_));
OR2X2 OR2X2_108 ( .A(e_reg_3_), .B(\digest[3] ), .Y(_abc_15497_new_n1045_));
OR2X2 OR2X2_1080 ( .A(_abc_15497_new_n3780_), .B(_abc_15497_new_n3912_), .Y(_abc_15497_new_n3913_));
OR2X2 OR2X2_1081 ( .A(_abc_15497_new_n3915_), .B(_abc_15497_new_n3914_), .Y(_abc_15497_new_n3916_));
OR2X2 OR2X2_1082 ( .A(_abc_15497_new_n3784_), .B(_abc_15497_new_n3916_), .Y(_abc_15497_new_n3917_));
OR2X2 OR2X2_1083 ( .A(_abc_15497_new_n3849_), .B(_abc_15497_new_n3845_), .Y(_abc_15497_new_n3920_));
OR2X2 OR2X2_1084 ( .A(e_reg_2_), .B(a_reg_29_), .Y(_abc_15497_new_n3921_));
OR2X2 OR2X2_1085 ( .A(_abc_15497_new_n3924_), .B(w_2_), .Y(_abc_15497_new_n3925_));
OR2X2 OR2X2_1086 ( .A(_abc_15497_new_n3931_), .B(_abc_15497_new_n3926_), .Y(_abc_15497_new_n3932_));
OR2X2 OR2X2_1087 ( .A(_abc_15497_new_n3933_), .B(_abc_15497_new_n3929_), .Y(_abc_15497_new_n3934_));
OR2X2 OR2X2_1088 ( .A(_abc_15497_new_n3919_), .B(_abc_15497_new_n3934_), .Y(_abc_15497_new_n3935_));
OR2X2 OR2X2_1089 ( .A(_abc_15497_new_n3938_), .B(_abc_15497_new_n3940_), .Y(_abc_15497_new_n3941_));
OR2X2 OR2X2_109 ( .A(_abc_15497_new_n1044_), .B(_abc_15497_new_n1048_), .Y(_abc_15497_new_n1049_));
OR2X2 OR2X2_1090 ( .A(_abc_15497_new_n3941_), .B(_abc_15497_new_n3936_), .Y(_abc_15497_new_n3942_));
OR2X2 OR2X2_1091 ( .A(_abc_15497_new_n3928_), .B(_abc_15497_new_n3920_), .Y(_abc_15497_new_n3944_));
OR2X2 OR2X2_1092 ( .A(_abc_15497_new_n3942_), .B(_abc_15497_new_n3945_), .Y(_abc_15497_new_n3946_));
OR2X2 OR2X2_1093 ( .A(_abc_15497_new_n3919_), .B(_abc_15497_new_n3945_), .Y(_abc_15497_new_n3950_));
OR2X2 OR2X2_1094 ( .A(_abc_15497_new_n3942_), .B(_abc_15497_new_n3934_), .Y(_abc_15497_new_n3951_));
OR2X2 OR2X2_1095 ( .A(_abc_15497_new_n3948_), .B(_abc_15497_new_n3953_), .Y(_abc_15497_new_n3954_));
OR2X2 OR2X2_1096 ( .A(_abc_15497_new_n3952_), .B(_abc_15497_new_n3949_), .Y(_abc_15497_new_n3956_));
OR2X2 OR2X2_1097 ( .A(_abc_15497_new_n3947_), .B(_abc_15497_new_n3899_), .Y(_abc_15497_new_n3957_));
OR2X2 OR2X2_1098 ( .A(_abc_15497_new_n3955_), .B(_abc_15497_new_n3959_), .Y(_abc_15497_new_n3960_));
OR2X2 OR2X2_1099 ( .A(_abc_15497_new_n3960_), .B(_abc_15497_new_n3897_), .Y(_abc_15497_new_n3961_));
OR2X2 OR2X2_11 ( .A(_abc_15497_new_n744_), .B(_abc_15497_new_n746_), .Y(_abc_15497_new_n747_));
OR2X2 OR2X2_110 ( .A(_abc_15497_new_n1050_), .B(_abc_15497_new_n1051_), .Y(_abc_15497_new_n1052_));
OR2X2 OR2X2_1100 ( .A(_abc_15497_new_n3879_), .B(_abc_15497_new_n3880_), .Y(_abc_15497_new_n3962_));
OR2X2 OR2X2_1101 ( .A(_abc_15497_new_n3958_), .B(_abc_15497_new_n3769_), .Y(_abc_15497_new_n3963_));
OR2X2 OR2X2_1102 ( .A(_abc_15497_new_n3954_), .B(_abc_15497_new_n3744_), .Y(_abc_15497_new_n3964_));
OR2X2 OR2X2_1103 ( .A(_abc_15497_new_n3965_), .B(_abc_15497_new_n3962_), .Y(_abc_15497_new_n3966_));
OR2X2 OR2X2_1104 ( .A(_abc_15497_new_n3967_), .B(_abc_15497_new_n3895_), .Y(_abc_15497_new_n3968_));
OR2X2 OR2X2_1105 ( .A(_abc_15497_new_n3970_), .B(_abc_15497_new_n3969_), .Y(_abc_15497_new_n3971_));
OR2X2 OR2X2_1106 ( .A(_abc_15497_new_n3971_), .B(_abc_15497_new_n3887_), .Y(_abc_15497_new_n3972_));
OR2X2 OR2X2_1107 ( .A(_abc_15497_new_n3975_), .B(_abc_15497_new_n3977_), .Y(_abc_15497_new_n3978_));
OR2X2 OR2X2_1108 ( .A(_abc_15497_new_n3974_), .B(_abc_15497_new_n3978_), .Y(_0a_reg_31_0__2_));
OR2X2 OR2X2_1109 ( .A(b_reg_3_), .B(c_reg_3_), .Y(_abc_15497_new_n3985_));
OR2X2 OR2X2_111 ( .A(_abc_15497_new_n1054_), .B(_abc_15497_new_n1042_), .Y(_0H4_reg_31_0__3_));
OR2X2 OR2X2_1110 ( .A(_abc_15497_new_n3990_), .B(_abc_15497_new_n3991_), .Y(_abc_15497_new_n3992_));
OR2X2 OR2X2_1111 ( .A(_abc_15497_new_n3775_), .B(_abc_15497_new_n3992_), .Y(_abc_15497_new_n3993_));
OR2X2 OR2X2_1112 ( .A(_abc_15497_new_n3984_), .B(b_reg_3_), .Y(_abc_15497_new_n3994_));
OR2X2 OR2X2_1113 ( .A(_abc_15497_new_n3780_), .B(_abc_15497_new_n3995_), .Y(_abc_15497_new_n3996_));
OR2X2 OR2X2_1114 ( .A(_abc_15497_new_n3998_), .B(_abc_15497_new_n3997_), .Y(_abc_15497_new_n3999_));
OR2X2 OR2X2_1115 ( .A(_abc_15497_new_n3784_), .B(_abc_15497_new_n3999_), .Y(_abc_15497_new_n4000_));
OR2X2 OR2X2_1116 ( .A(e_reg_3_), .B(a_reg_30_), .Y(_abc_15497_new_n4006_));
OR2X2 OR2X2_1117 ( .A(_abc_15497_new_n4011_), .B(_abc_15497_new_n4012_), .Y(_abc_15497_new_n4013_));
OR2X2 OR2X2_1118 ( .A(_abc_15497_new_n4015_), .B(_abc_15497_new_n4016_), .Y(_abc_15497_new_n4017_));
OR2X2 OR2X2_1119 ( .A(_abc_15497_new_n4017_), .B(_abc_15497_new_n4002_), .Y(_abc_15497_new_n4018_));
OR2X2 OR2X2_112 ( .A(e_reg_4_), .B(\digest[4] ), .Y(_abc_15497_new_n1056_));
OR2X2 OR2X2_1120 ( .A(_abc_15497_new_n4019_), .B(_abc_15497_new_n4020_), .Y(_abc_15497_new_n4021_));
OR2X2 OR2X2_1121 ( .A(_abc_15497_new_n4021_), .B(_abc_15497_new_n3983_), .Y(_abc_15497_new_n4022_));
OR2X2 OR2X2_1122 ( .A(_abc_15497_new_n4023_), .B(_abc_15497_new_n4025_), .Y(_abc_15497_new_n4026_));
OR2X2 OR2X2_1123 ( .A(_abc_15497_new_n4027_), .B(_abc_15497_new_n3775_), .Y(_abc_15497_new_n4028_));
OR2X2 OR2X2_1124 ( .A(_abc_15497_new_n4030_), .B(_abc_15497_new_n4029_), .Y(_abc_15497_new_n4031_));
OR2X2 OR2X2_1125 ( .A(_abc_15497_new_n4031_), .B(_abc_15497_new_n3803_), .Y(_abc_15497_new_n4032_));
OR2X2 OR2X2_1126 ( .A(_abc_15497_new_n4035_), .B(_abc_15497_new_n4036_), .Y(_abc_15497_new_n4037_));
OR2X2 OR2X2_1127 ( .A(_abc_15497_new_n4038_), .B(_abc_15497_new_n4034_), .Y(_abc_15497_new_n4039_));
OR2X2 OR2X2_1128 ( .A(_abc_15497_new_n3980_), .B(_abc_15497_new_n4039_), .Y(_abc_15497_new_n4040_));
OR2X2 OR2X2_1129 ( .A(_abc_15497_new_n4037_), .B(_abc_15497_new_n3981_), .Y(_abc_15497_new_n4042_));
OR2X2 OR2X2_113 ( .A(_abc_15497_new_n1050_), .B(_abc_15497_new_n1061_), .Y(_abc_15497_new_n1062_));
OR2X2 OR2X2_1130 ( .A(_abc_15497_new_n4033_), .B(_abc_15497_new_n3982_), .Y(_abc_15497_new_n4043_));
OR2X2 OR2X2_1131 ( .A(_abc_15497_new_n4041_), .B(_abc_15497_new_n4044_), .Y(_abc_15497_new_n4045_));
OR2X2 OR2X2_1132 ( .A(_abc_15497_new_n4048_), .B(_abc_15497_new_n4050_), .Y(_abc_15497_new_n4051_));
OR2X2 OR2X2_1133 ( .A(_abc_15497_new_n4047_), .B(_abc_15497_new_n4051_), .Y(_0a_reg_31_0__3_));
OR2X2 OR2X2_1134 ( .A(_abc_15497_new_n4055_), .B(_abc_15497_new_n4034_), .Y(_abc_15497_new_n4056_));
OR2X2 OR2X2_1135 ( .A(_abc_15497_new_n4054_), .B(_abc_15497_new_n4056_), .Y(_abc_15497_new_n4057_));
OR2X2 OR2X2_1136 ( .A(b_reg_4_), .B(c_reg_4_), .Y(_abc_15497_new_n4064_));
OR2X2 OR2X2_1137 ( .A(_abc_15497_new_n4069_), .B(_abc_15497_new_n4070_), .Y(_abc_15497_new_n4071_));
OR2X2 OR2X2_1138 ( .A(_abc_15497_new_n4075_), .B(_abc_15497_new_n4065_), .Y(_abc_15497_new_n4076_));
OR2X2 OR2X2_1139 ( .A(_abc_15497_new_n4079_), .B(_abc_15497_new_n4078_), .Y(_abc_15497_new_n4080_));
OR2X2 OR2X2_114 ( .A(_abc_15497_new_n1063_), .B(_abc_15497_new_n1060_), .Y(_abc_15497_new_n1064_));
OR2X2 OR2X2_1140 ( .A(_abc_15497_new_n4077_), .B(_abc_15497_new_n4082_), .Y(_abc_15497_new_n4083_));
OR2X2 OR2X2_1141 ( .A(_abc_15497_new_n4073_), .B(_abc_15497_new_n4083_), .Y(_abc_15497_new_n4084_));
OR2X2 OR2X2_1142 ( .A(_abc_15497_new_n4012_), .B(_abc_15497_new_n4007_), .Y(_abc_15497_new_n4085_));
OR2X2 OR2X2_1143 ( .A(e_reg_4_), .B(a_reg_31_), .Y(_abc_15497_new_n4087_));
OR2X2 OR2X2_1144 ( .A(_abc_15497_new_n4092_), .B(_abc_15497_new_n4093_), .Y(_abc_15497_new_n4094_));
OR2X2 OR2X2_1145 ( .A(_abc_15497_new_n4096_), .B(_abc_15497_new_n4098_), .Y(_abc_15497_new_n4099_));
OR2X2 OR2X2_1146 ( .A(_abc_15497_new_n4103_), .B(_abc_15497_new_n4101_), .Y(_abc_15497_new_n4104_));
OR2X2 OR2X2_1147 ( .A(_abc_15497_new_n4104_), .B(_abc_15497_new_n4062_), .Y(_abc_15497_new_n4105_));
OR2X2 OR2X2_1148 ( .A(_abc_15497_new_n4102_), .B(_abc_15497_new_n4099_), .Y(_abc_15497_new_n4107_));
OR2X2 OR2X2_1149 ( .A(_abc_15497_new_n4100_), .B(_abc_15497_new_n4084_), .Y(_abc_15497_new_n4108_));
OR2X2 OR2X2_115 ( .A(_abc_15497_new_n1065_), .B(_abc_15497_new_n1046_), .Y(_abc_15497_new_n1066_));
OR2X2 OR2X2_1150 ( .A(_abc_15497_new_n4109_), .B(_abc_15497_new_n4106_), .Y(_abc_15497_new_n4110_));
OR2X2 OR2X2_1151 ( .A(_abc_15497_new_n4114_), .B(_abc_15497_new_n4113_), .Y(_abc_15497_new_n4115_));
OR2X2 OR2X2_1152 ( .A(_abc_15497_new_n4116_), .B(_abc_15497_new_n4112_), .Y(_abc_15497_new_n4117_));
OR2X2 OR2X2_1153 ( .A(_abc_15497_new_n4036_), .B(_abc_15497_new_n4029_), .Y(_abc_15497_new_n4119_));
OR2X2 OR2X2_1154 ( .A(_abc_15497_new_n4115_), .B(_abc_15497_new_n4059_), .Y(_abc_15497_new_n4120_));
OR2X2 OR2X2_1155 ( .A(_abc_15497_new_n4111_), .B(_abc_15497_new_n4060_), .Y(_abc_15497_new_n4121_));
OR2X2 OR2X2_1156 ( .A(_abc_15497_new_n4118_), .B(_abc_15497_new_n4123_), .Y(_abc_15497_new_n4124_));
OR2X2 OR2X2_1157 ( .A(_abc_15497_new_n4057_), .B(_abc_15497_new_n4125_), .Y(_abc_15497_new_n4126_));
OR2X2 OR2X2_1158 ( .A(_abc_15497_new_n4131_), .B(_abc_15497_new_n4133_), .Y(_abc_15497_new_n4134_));
OR2X2 OR2X2_1159 ( .A(_abc_15497_new_n4130_), .B(_abc_15497_new_n4134_), .Y(_0a_reg_31_0__4_));
OR2X2 OR2X2_116 ( .A(_abc_15497_new_n1066_), .B(_abc_15497_new_n1059_), .Y(_abc_15497_new_n1067_));
OR2X2 OR2X2_1160 ( .A(_abc_15497_new_n4117_), .B(_abc_15497_new_n4058_), .Y(_abc_15497_new_n4136_));
OR2X2 OR2X2_1161 ( .A(_abc_15497_new_n4112_), .B(_abc_15497_new_n4113_), .Y(_abc_15497_new_n4139_));
OR2X2 OR2X2_1162 ( .A(_abc_15497_new_n4101_), .B(_abc_15497_new_n4096_), .Y(_abc_15497_new_n4140_));
OR2X2 OR2X2_1163 ( .A(b_reg_5_), .B(c_reg_5_), .Y(_abc_15497_new_n4142_));
OR2X2 OR2X2_1164 ( .A(_abc_15497_new_n4147_), .B(_abc_15497_new_n4148_), .Y(_abc_15497_new_n4149_));
OR2X2 OR2X2_1165 ( .A(_abc_15497_new_n4153_), .B(_abc_15497_new_n4143_), .Y(_abc_15497_new_n4154_));
OR2X2 OR2X2_1166 ( .A(_abc_15497_new_n4157_), .B(_abc_15497_new_n4156_), .Y(_abc_15497_new_n4158_));
OR2X2 OR2X2_1167 ( .A(_abc_15497_new_n4155_), .B(_abc_15497_new_n4160_), .Y(_abc_15497_new_n4161_));
OR2X2 OR2X2_1168 ( .A(_abc_15497_new_n4151_), .B(_abc_15497_new_n4161_), .Y(_abc_15497_new_n4162_));
OR2X2 OR2X2_1169 ( .A(_abc_15497_new_n4093_), .B(_abc_15497_new_n4088_), .Y(_abc_15497_new_n4164_));
OR2X2 OR2X2_117 ( .A(_abc_15497_new_n1068_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n1069_));
OR2X2 OR2X2_1170 ( .A(e_reg_5_), .B(a_reg_0_), .Y(_abc_15497_new_n4166_));
OR2X2 OR2X2_1171 ( .A(_abc_15497_new_n4171_), .B(_abc_15497_new_n4172_), .Y(_abc_15497_new_n4173_));
OR2X2 OR2X2_1172 ( .A(_abc_15497_new_n4175_), .B(_abc_15497_new_n4177_), .Y(_abc_15497_new_n4178_));
OR2X2 OR2X2_1173 ( .A(_abc_15497_new_n4163_), .B(_abc_15497_new_n4178_), .Y(_abc_15497_new_n4179_));
OR2X2 OR2X2_1174 ( .A(_abc_15497_new_n4180_), .B(_abc_15497_new_n4162_), .Y(_abc_15497_new_n4181_));
OR2X2 OR2X2_1175 ( .A(_abc_15497_new_n4182_), .B(_abc_15497_new_n4140_), .Y(_abc_15497_new_n4183_));
OR2X2 OR2X2_1176 ( .A(_abc_15497_new_n4187_), .B(_abc_15497_new_n4186_), .Y(_abc_15497_new_n4188_));
OR2X2 OR2X2_1177 ( .A(_abc_15497_new_n4188_), .B(_abc_15497_new_n4185_), .Y(_abc_15497_new_n4189_));
OR2X2 OR2X2_1178 ( .A(_abc_15497_new_n4190_), .B(_abc_15497_new_n4059_), .Y(_abc_15497_new_n4191_));
OR2X2 OR2X2_1179 ( .A(_abc_15497_new_n4192_), .B(_abc_15497_new_n4193_), .Y(_abc_15497_new_n4194_));
OR2X2 OR2X2_118 ( .A(_abc_15497_new_n699_), .B(\digest[4] ), .Y(_abc_15497_new_n1070_));
OR2X2 OR2X2_1180 ( .A(_abc_15497_new_n4194_), .B(_abc_15497_new_n4060_), .Y(_abc_15497_new_n4195_));
OR2X2 OR2X2_1181 ( .A(_abc_15497_new_n4199_), .B(_abc_15497_new_n4200_), .Y(_abc_15497_new_n4201_));
OR2X2 OR2X2_1182 ( .A(_abc_15497_new_n4202_), .B(_abc_15497_new_n4197_), .Y(_abc_15497_new_n4203_));
OR2X2 OR2X2_1183 ( .A(_abc_15497_new_n4138_), .B(_abc_15497_new_n4204_), .Y(_abc_15497_new_n4205_));
OR2X2 OR2X2_1184 ( .A(_abc_15497_new_n4137_), .B(_abc_15497_new_n4203_), .Y(_abc_15497_new_n4206_));
OR2X2 OR2X2_1185 ( .A(_abc_15497_new_n4209_), .B(_abc_15497_new_n4211_), .Y(_abc_15497_new_n4212_));
OR2X2 OR2X2_1186 ( .A(_abc_15497_new_n4208_), .B(_abc_15497_new_n4212_), .Y(_0a_reg_31_0__5_));
OR2X2 OR2X2_1187 ( .A(_abc_15497_new_n4124_), .B(_abc_15497_new_n4203_), .Y(_abc_15497_new_n4214_));
OR2X2 OR2X2_1188 ( .A(_abc_15497_new_n4136_), .B(_abc_15497_new_n4202_), .Y(_abc_15497_new_n4218_));
OR2X2 OR2X2_1189 ( .A(_abc_15497_new_n4216_), .B(_abc_15497_new_n4220_), .Y(_abc_15497_new_n4221_));
OR2X2 OR2X2_119 ( .A(_abc_15497_new_n1070_), .B(digest_update), .Y(_abc_15497_new_n1071_));
OR2X2 OR2X2_1190 ( .A(_abc_15497_new_n4200_), .B(_abc_15497_new_n4193_), .Y(_abc_15497_new_n4222_));
OR2X2 OR2X2_1191 ( .A(_abc_15497_new_n4186_), .B(_abc_15497_new_n4175_), .Y(_abc_15497_new_n4223_));
OR2X2 OR2X2_1192 ( .A(b_reg_6_), .B(c_reg_6_), .Y(_abc_15497_new_n4225_));
OR2X2 OR2X2_1193 ( .A(_abc_15497_new_n4230_), .B(_abc_15497_new_n4231_), .Y(_abc_15497_new_n4232_));
OR2X2 OR2X2_1194 ( .A(_abc_15497_new_n4236_), .B(_abc_15497_new_n4226_), .Y(_abc_15497_new_n4237_));
OR2X2 OR2X2_1195 ( .A(_abc_15497_new_n4240_), .B(_abc_15497_new_n4239_), .Y(_abc_15497_new_n4241_));
OR2X2 OR2X2_1196 ( .A(_abc_15497_new_n4238_), .B(_abc_15497_new_n4243_), .Y(_abc_15497_new_n4244_));
OR2X2 OR2X2_1197 ( .A(_abc_15497_new_n4234_), .B(_abc_15497_new_n4244_), .Y(_abc_15497_new_n4245_));
OR2X2 OR2X2_1198 ( .A(_abc_15497_new_n4172_), .B(_abc_15497_new_n4167_), .Y(_abc_15497_new_n4247_));
OR2X2 OR2X2_1199 ( .A(e_reg_6_), .B(a_reg_1_), .Y(_abc_15497_new_n4249_));
OR2X2 OR2X2_12 ( .A(_abc_15497_new_n751_), .B(_abc_15497_new_n731_), .Y(_abc_15497_new_n752_));
OR2X2 OR2X2_120 ( .A(_abc_15497_new_n1073_), .B(_abc_15497_new_n1057_), .Y(_abc_15497_new_n1074_));
OR2X2 OR2X2_1200 ( .A(_abc_15497_new_n4254_), .B(_abc_15497_new_n4255_), .Y(_abc_15497_new_n4256_));
OR2X2 OR2X2_1201 ( .A(_abc_15497_new_n4258_), .B(_abc_15497_new_n4260_), .Y(_abc_15497_new_n4261_));
OR2X2 OR2X2_1202 ( .A(_abc_15497_new_n4246_), .B(_abc_15497_new_n4261_), .Y(_abc_15497_new_n4262_));
OR2X2 OR2X2_1203 ( .A(_abc_15497_new_n4263_), .B(_abc_15497_new_n4245_), .Y(_abc_15497_new_n4264_));
OR2X2 OR2X2_1204 ( .A(_abc_15497_new_n4265_), .B(_abc_15497_new_n4223_), .Y(_abc_15497_new_n4266_));
OR2X2 OR2X2_1205 ( .A(_abc_15497_new_n4270_), .B(_abc_15497_new_n4269_), .Y(_abc_15497_new_n4271_));
OR2X2 OR2X2_1206 ( .A(_abc_15497_new_n4271_), .B(_abc_15497_new_n4268_), .Y(_abc_15497_new_n4272_));
OR2X2 OR2X2_1207 ( .A(_abc_15497_new_n4273_), .B(_abc_15497_new_n3769_), .Y(_abc_15497_new_n4274_));
OR2X2 OR2X2_1208 ( .A(_abc_15497_new_n4275_), .B(_abc_15497_new_n4276_), .Y(_abc_15497_new_n4277_));
OR2X2 OR2X2_1209 ( .A(_abc_15497_new_n4277_), .B(_abc_15497_new_n3744_), .Y(_abc_15497_new_n4278_));
OR2X2 OR2X2_121 ( .A(e_reg_5_), .B(\digest[5] ), .Y(_abc_15497_new_n1075_));
OR2X2 OR2X2_1210 ( .A(_abc_15497_new_n4282_), .B(_abc_15497_new_n4283_), .Y(_abc_15497_new_n4284_));
OR2X2 OR2X2_1211 ( .A(_abc_15497_new_n4285_), .B(_abc_15497_new_n4280_), .Y(_abc_15497_new_n4286_));
OR2X2 OR2X2_1212 ( .A(_abc_15497_new_n4221_), .B(_abc_15497_new_n4287_), .Y(_abc_15497_new_n4288_));
OR2X2 OR2X2_1213 ( .A(_abc_15497_new_n4293_), .B(_abc_15497_new_n4295_), .Y(_abc_15497_new_n4296_));
OR2X2 OR2X2_1214 ( .A(_abc_15497_new_n4292_), .B(_abc_15497_new_n4296_), .Y(_0a_reg_31_0__6_));
OR2X2 OR2X2_1215 ( .A(_abc_15497_new_n4283_), .B(_abc_15497_new_n4276_), .Y(_abc_15497_new_n4300_));
OR2X2 OR2X2_1216 ( .A(b_reg_7_), .B(c_reg_7_), .Y(_abc_15497_new_n4305_));
OR2X2 OR2X2_1217 ( .A(_abc_15497_new_n4310_), .B(_abc_15497_new_n4311_), .Y(_abc_15497_new_n4312_));
OR2X2 OR2X2_1218 ( .A(_abc_15497_new_n3775_), .B(_abc_15497_new_n4312_), .Y(_abc_15497_new_n4313_));
OR2X2 OR2X2_1219 ( .A(_abc_15497_new_n4315_), .B(_abc_15497_new_n4306_), .Y(_abc_15497_new_n4316_));
OR2X2 OR2X2_122 ( .A(_abc_15497_new_n1074_), .B(_abc_15497_new_n1078_), .Y(_abc_15497_new_n1079_));
OR2X2 OR2X2_1220 ( .A(_abc_15497_new_n4320_), .B(_abc_15497_new_n4319_), .Y(_abc_15497_new_n4321_));
OR2X2 OR2X2_1221 ( .A(_abc_15497_new_n3784_), .B(_abc_15497_new_n4321_), .Y(_abc_15497_new_n4322_));
OR2X2 OR2X2_1222 ( .A(_abc_15497_new_n4255_), .B(_abc_15497_new_n4250_), .Y(_abc_15497_new_n4326_));
OR2X2 OR2X2_1223 ( .A(e_reg_7_), .B(a_reg_2_), .Y(_abc_15497_new_n4328_));
OR2X2 OR2X2_1224 ( .A(_abc_15497_new_n4333_), .B(_abc_15497_new_n4334_), .Y(_abc_15497_new_n4335_));
OR2X2 OR2X2_1225 ( .A(_abc_15497_new_n4336_), .B(_abc_15497_new_n4326_), .Y(_abc_15497_new_n4339_));
OR2X2 OR2X2_1226 ( .A(_abc_15497_new_n4342_), .B(_abc_15497_new_n4337_), .Y(_abc_15497_new_n4343_));
OR2X2 OR2X2_1227 ( .A(_abc_15497_new_n4341_), .B(_abc_15497_new_n4344_), .Y(_abc_15497_new_n4345_));
OR2X2 OR2X2_1228 ( .A(_abc_15497_new_n4347_), .B(_abc_15497_new_n4348_), .Y(_abc_15497_new_n4349_));
OR2X2 OR2X2_1229 ( .A(_abc_15497_new_n4350_), .B(_abc_15497_new_n4353_), .Y(_abc_15497_new_n4354_));
OR2X2 OR2X2_123 ( .A(_abc_15497_new_n1080_), .B(_abc_15497_new_n1081_), .Y(_abc_15497_new_n1082_));
OR2X2 OR2X2_1230 ( .A(_abc_15497_new_n4299_), .B(_abc_15497_new_n4354_), .Y(_abc_15497_new_n4355_));
OR2X2 OR2X2_1231 ( .A(_abc_15497_new_n4356_), .B(_abc_15497_new_n4357_), .Y(_abc_15497_new_n4358_));
OR2X2 OR2X2_1232 ( .A(_abc_15497_new_n4361_), .B(_abc_15497_new_n4363_), .Y(_abc_15497_new_n4364_));
OR2X2 OR2X2_1233 ( .A(_abc_15497_new_n4360_), .B(_abc_15497_new_n4364_), .Y(_0a_reg_31_0__7_));
OR2X2 OR2X2_1234 ( .A(_abc_15497_new_n4341_), .B(_abc_15497_new_n4337_), .Y(_abc_15497_new_n4367_));
OR2X2 OR2X2_1235 ( .A(b_reg_8_), .B(c_reg_8_), .Y(_abc_15497_new_n4369_));
OR2X2 OR2X2_1236 ( .A(_abc_15497_new_n4374_), .B(_abc_15497_new_n4375_), .Y(_abc_15497_new_n4376_));
OR2X2 OR2X2_1237 ( .A(_abc_15497_new_n3775_), .B(_abc_15497_new_n4376_), .Y(_abc_15497_new_n4377_));
OR2X2 OR2X2_1238 ( .A(_abc_15497_new_n4379_), .B(_abc_15497_new_n4370_), .Y(_abc_15497_new_n4380_));
OR2X2 OR2X2_1239 ( .A(_abc_15497_new_n4384_), .B(_abc_15497_new_n4383_), .Y(_abc_15497_new_n4385_));
OR2X2 OR2X2_124 ( .A(_abc_15497_new_n699_), .B(\digest[5] ), .Y(_abc_15497_new_n1085_));
OR2X2 OR2X2_1240 ( .A(_abc_15497_new_n3784_), .B(_abc_15497_new_n4385_), .Y(_abc_15497_new_n4386_));
OR2X2 OR2X2_1241 ( .A(_abc_15497_new_n4334_), .B(_abc_15497_new_n4329_), .Y(_abc_15497_new_n4389_));
OR2X2 OR2X2_1242 ( .A(e_reg_8_), .B(a_reg_3_), .Y(_abc_15497_new_n4391_));
OR2X2 OR2X2_1243 ( .A(_abc_15497_new_n4396_), .B(_abc_15497_new_n4397_), .Y(_abc_15497_new_n4398_));
OR2X2 OR2X2_1244 ( .A(_abc_15497_new_n4399_), .B(_abc_15497_new_n4389_), .Y(_abc_15497_new_n4401_));
OR2X2 OR2X2_1245 ( .A(_abc_15497_new_n4402_), .B(_abc_15497_new_n4400_), .Y(_abc_15497_new_n4403_));
OR2X2 OR2X2_1246 ( .A(_abc_15497_new_n4403_), .B(_abc_15497_new_n4388_), .Y(_abc_15497_new_n4404_));
OR2X2 OR2X2_1247 ( .A(_abc_15497_new_n4405_), .B(_abc_15497_new_n4407_), .Y(_abc_15497_new_n4408_));
OR2X2 OR2X2_1248 ( .A(_abc_15497_new_n4343_), .B(_abc_15497_new_n4324_), .Y(_abc_15497_new_n4411_));
OR2X2 OR2X2_1249 ( .A(_abc_15497_new_n4413_), .B(_abc_15497_new_n4414_), .Y(_abc_15497_new_n4415_));
OR2X2 OR2X2_125 ( .A(_abc_15497_new_n1084_), .B(_abc_15497_new_n1086_), .Y(_0H4_reg_31_0__5_));
OR2X2 OR2X2_1250 ( .A(_abc_15497_new_n4410_), .B(_abc_15497_new_n4416_), .Y(_abc_15497_new_n4417_));
OR2X2 OR2X2_1251 ( .A(_abc_15497_new_n4415_), .B(_abc_15497_new_n4412_), .Y(_abc_15497_new_n4419_));
OR2X2 OR2X2_1252 ( .A(_abc_15497_new_n4409_), .B(_abc_15497_new_n4367_), .Y(_abc_15497_new_n4420_));
OR2X2 OR2X2_1253 ( .A(_abc_15497_new_n4418_), .B(_abc_15497_new_n4422_), .Y(_abc_15497_new_n4423_));
OR2X2 OR2X2_1254 ( .A(_abc_15497_new_n4425_), .B(_abc_15497_new_n4426_), .Y(_abc_15497_new_n4427_));
OR2X2 OR2X2_1255 ( .A(_abc_15497_new_n3972_), .B(_abc_15497_new_n4039_), .Y(_abc_15497_new_n4429_));
OR2X2 OR2X2_1256 ( .A(_abc_15497_new_n4286_), .B(_abc_15497_new_n4354_), .Y(_abc_15497_new_n4433_));
OR2X2 OR2X2_1257 ( .A(_abc_15497_new_n4214_), .B(_abc_15497_new_n4433_), .Y(_abc_15497_new_n4434_));
OR2X2 OR2X2_1258 ( .A(_abc_15497_new_n4432_), .B(_abc_15497_new_n4434_), .Y(_abc_15497_new_n4435_));
OR2X2 OR2X2_1259 ( .A(_abc_15497_new_n4437_), .B(_abc_15497_new_n4353_), .Y(_abc_15497_new_n4438_));
OR2X2 OR2X2_126 ( .A(_abc_15497_new_n1088_), .B(_abc_15497_new_n1076_), .Y(_abc_15497_new_n1089_));
OR2X2 OR2X2_1260 ( .A(_abc_15497_new_n4433_), .B(_abc_15497_new_n4219_), .Y(_abc_15497_new_n4439_));
OR2X2 OR2X2_1261 ( .A(_abc_15497_new_n4442_), .B(_abc_15497_new_n4428_), .Y(_abc_15497_new_n4443_));
OR2X2 OR2X2_1262 ( .A(_abc_15497_new_n4448_), .B(_abc_15497_new_n4449_), .Y(_abc_15497_new_n4450_));
OR2X2 OR2X2_1263 ( .A(_abc_15497_new_n4447_), .B(_abc_15497_new_n4450_), .Y(_0a_reg_31_0__8_));
OR2X2 OR2X2_1264 ( .A(_abc_15497_new_n4423_), .B(_abc_15497_new_n4348_), .Y(_abc_15497_new_n4452_));
OR2X2 OR2X2_1265 ( .A(_abc_15497_new_n4417_), .B(_abc_15497_new_n3774_), .Y(_abc_15497_new_n4454_));
OR2X2 OR2X2_1266 ( .A(b_reg_9_), .B(c_reg_9_), .Y(_abc_15497_new_n4459_));
OR2X2 OR2X2_1267 ( .A(_abc_15497_new_n4464_), .B(_abc_15497_new_n4465_), .Y(_abc_15497_new_n4466_));
OR2X2 OR2X2_1268 ( .A(_abc_15497_new_n3775_), .B(_abc_15497_new_n4466_), .Y(_abc_15497_new_n4467_));
OR2X2 OR2X2_1269 ( .A(_abc_15497_new_n4469_), .B(_abc_15497_new_n4460_), .Y(_abc_15497_new_n4470_));
OR2X2 OR2X2_127 ( .A(e_reg_6_), .B(\digest[6] ), .Y(_abc_15497_new_n1090_));
OR2X2 OR2X2_1270 ( .A(_abc_15497_new_n4474_), .B(_abc_15497_new_n4473_), .Y(_abc_15497_new_n4475_));
OR2X2 OR2X2_1271 ( .A(_abc_15497_new_n3784_), .B(_abc_15497_new_n4475_), .Y(_abc_15497_new_n4476_));
OR2X2 OR2X2_1272 ( .A(_abc_15497_new_n4397_), .B(_abc_15497_new_n4392_), .Y(_abc_15497_new_n4480_));
OR2X2 OR2X2_1273 ( .A(e_reg_9_), .B(a_reg_4_), .Y(_abc_15497_new_n4482_));
OR2X2 OR2X2_1274 ( .A(_abc_15497_new_n4487_), .B(_abc_15497_new_n4488_), .Y(_abc_15497_new_n4489_));
OR2X2 OR2X2_1275 ( .A(_abc_15497_new_n4490_), .B(_abc_15497_new_n4480_), .Y(_abc_15497_new_n4493_));
OR2X2 OR2X2_1276 ( .A(_abc_15497_new_n4496_), .B(_abc_15497_new_n4491_), .Y(_abc_15497_new_n4497_));
OR2X2 OR2X2_1277 ( .A(_abc_15497_new_n4495_), .B(_abc_15497_new_n4498_), .Y(_abc_15497_new_n4499_));
OR2X2 OR2X2_1278 ( .A(_abc_15497_new_n4413_), .B(_abc_15497_new_n4400_), .Y(_abc_15497_new_n4501_));
OR2X2 OR2X2_1279 ( .A(_abc_15497_new_n4497_), .B(_abc_15497_new_n4478_), .Y(_abc_15497_new_n4502_));
OR2X2 OR2X2_128 ( .A(_abc_15497_new_n1089_), .B(_abc_15497_new_n1093_), .Y(_abc_15497_new_n1094_));
OR2X2 OR2X2_1280 ( .A(_abc_15497_new_n4479_), .B(_abc_15497_new_n4494_), .Y(_abc_15497_new_n4503_));
OR2X2 OR2X2_1281 ( .A(_abc_15497_new_n4505_), .B(_abc_15497_new_n4500_), .Y(_abc_15497_new_n4506_));
OR2X2 OR2X2_1282 ( .A(_abc_15497_new_n4504_), .B(_abc_15497_new_n4501_), .Y(_abc_15497_new_n4508_));
OR2X2 OR2X2_1283 ( .A(_abc_15497_new_n4499_), .B(_abc_15497_new_n4457_), .Y(_abc_15497_new_n4509_));
OR2X2 OR2X2_1284 ( .A(_abc_15497_new_n4507_), .B(_abc_15497_new_n4511_), .Y(_abc_15497_new_n4512_));
OR2X2 OR2X2_1285 ( .A(_abc_15497_new_n4514_), .B(_abc_15497_new_n4515_), .Y(_abc_15497_new_n4516_));
OR2X2 OR2X2_1286 ( .A(_abc_15497_new_n4453_), .B(_abc_15497_new_n4516_), .Y(_abc_15497_new_n4517_));
OR2X2 OR2X2_1287 ( .A(_abc_15497_new_n4518_), .B(_abc_15497_new_n4519_), .Y(_abc_15497_new_n4520_));
OR2X2 OR2X2_1288 ( .A(_abc_15497_new_n4523_), .B(_abc_15497_new_n4524_), .Y(_abc_15497_new_n4525_));
OR2X2 OR2X2_1289 ( .A(_abc_15497_new_n4522_), .B(_abc_15497_new_n4525_), .Y(_0a_reg_31_0__9_));
OR2X2 OR2X2_129 ( .A(_abc_15497_new_n1095_), .B(_abc_15497_new_n1096_), .Y(_abc_15497_new_n1097_));
OR2X2 OR2X2_1290 ( .A(_abc_15497_new_n4452_), .B(_abc_15497_new_n4515_), .Y(_abc_15497_new_n4528_));
OR2X2 OR2X2_1291 ( .A(_abc_15497_new_n4516_), .B(_abc_15497_new_n4427_), .Y(_abc_15497_new_n4531_));
OR2X2 OR2X2_1292 ( .A(_abc_15497_new_n4533_), .B(_abc_15497_new_n4530_), .Y(_abc_15497_new_n4534_));
OR2X2 OR2X2_1293 ( .A(_abc_15497_new_n4511_), .B(_abc_15497_new_n4505_), .Y(_abc_15497_new_n4535_));
OR2X2 OR2X2_1294 ( .A(_abc_15497_new_n4495_), .B(_abc_15497_new_n4491_), .Y(_abc_15497_new_n4536_));
OR2X2 OR2X2_1295 ( .A(b_reg_10_), .B(c_reg_10_), .Y(_abc_15497_new_n4538_));
OR2X2 OR2X2_1296 ( .A(_abc_15497_new_n4543_), .B(_abc_15497_new_n4544_), .Y(_abc_15497_new_n4545_));
OR2X2 OR2X2_1297 ( .A(_abc_15497_new_n3775_), .B(_abc_15497_new_n4545_), .Y(_abc_15497_new_n4546_));
OR2X2 OR2X2_1298 ( .A(_abc_15497_new_n4548_), .B(_abc_15497_new_n4539_), .Y(_abc_15497_new_n4549_));
OR2X2 OR2X2_1299 ( .A(_abc_15497_new_n4553_), .B(_abc_15497_new_n4552_), .Y(_abc_15497_new_n4554_));
OR2X2 OR2X2_13 ( .A(_abc_15497_new_n750_), .B(_abc_15497_new_n752_), .Y(_abc_15497_new_n753_));
OR2X2 OR2X2_130 ( .A(_abc_15497_new_n699_), .B(\digest[6] ), .Y(_abc_15497_new_n1100_));
OR2X2 OR2X2_1300 ( .A(_abc_15497_new_n3784_), .B(_abc_15497_new_n4554_), .Y(_abc_15497_new_n4555_));
OR2X2 OR2X2_1301 ( .A(_abc_15497_new_n4488_), .B(_abc_15497_new_n4483_), .Y(_abc_15497_new_n4558_));
OR2X2 OR2X2_1302 ( .A(e_reg_10_), .B(a_reg_5_), .Y(_abc_15497_new_n4560_));
OR2X2 OR2X2_1303 ( .A(_abc_15497_new_n4565_), .B(_abc_15497_new_n4566_), .Y(_abc_15497_new_n4567_));
OR2X2 OR2X2_1304 ( .A(_abc_15497_new_n4568_), .B(_abc_15497_new_n4558_), .Y(_abc_15497_new_n4570_));
OR2X2 OR2X2_1305 ( .A(_abc_15497_new_n4571_), .B(_abc_15497_new_n4569_), .Y(_abc_15497_new_n4572_));
OR2X2 OR2X2_1306 ( .A(_abc_15497_new_n4572_), .B(_abc_15497_new_n4557_), .Y(_abc_15497_new_n4573_));
OR2X2 OR2X2_1307 ( .A(_abc_15497_new_n4574_), .B(_abc_15497_new_n4576_), .Y(_abc_15497_new_n4577_));
OR2X2 OR2X2_1308 ( .A(_abc_15497_new_n4578_), .B(_abc_15497_new_n4536_), .Y(_abc_15497_new_n4579_));
OR2X2 OR2X2_1309 ( .A(_abc_15497_new_n4581_), .B(_abc_15497_new_n4582_), .Y(_abc_15497_new_n4583_));
OR2X2 OR2X2_131 ( .A(_abc_15497_new_n1099_), .B(_abc_15497_new_n1101_), .Y(_0H4_reg_31_0__6_));
OR2X2 OR2X2_1310 ( .A(_abc_15497_new_n4583_), .B(_abc_15497_new_n4580_), .Y(_abc_15497_new_n4584_));
OR2X2 OR2X2_1311 ( .A(_abc_15497_new_n4585_), .B(_abc_15497_new_n3774_), .Y(_abc_15497_new_n4586_));
OR2X2 OR2X2_1312 ( .A(_abc_15497_new_n4588_), .B(_abc_15497_new_n4587_), .Y(_abc_15497_new_n4589_));
OR2X2 OR2X2_1313 ( .A(_abc_15497_new_n4589_), .B(_abc_15497_new_n3784_), .Y(_abc_15497_new_n4590_));
OR2X2 OR2X2_1314 ( .A(_abc_15497_new_n4506_), .B(_abc_15497_new_n4060_), .Y(_abc_15497_new_n4593_));
OR2X2 OR2X2_1315 ( .A(_abc_15497_new_n4595_), .B(_abc_15497_new_n4596_), .Y(_abc_15497_new_n4597_));
OR2X2 OR2X2_1316 ( .A(_abc_15497_new_n4598_), .B(_abc_15497_new_n4592_), .Y(_abc_15497_new_n4599_));
OR2X2 OR2X2_1317 ( .A(_abc_15497_new_n4534_), .B(_abc_15497_new_n4600_), .Y(_abc_15497_new_n4601_));
OR2X2 OR2X2_1318 ( .A(_abc_15497_new_n4606_), .B(_abc_15497_new_n4608_), .Y(_abc_15497_new_n4609_));
OR2X2 OR2X2_1319 ( .A(_abc_15497_new_n4605_), .B(_abc_15497_new_n4609_), .Y(_0a_reg_31_0__10_));
OR2X2 OR2X2_132 ( .A(_abc_15497_new_n699_), .B(\digest[7] ), .Y(_abc_15497_new_n1103_));
OR2X2 OR2X2_1320 ( .A(_abc_15497_new_n4596_), .B(_abc_15497_new_n4588_), .Y(_abc_15497_new_n4613_));
OR2X2 OR2X2_1321 ( .A(b_reg_11_), .B(c_reg_11_), .Y(_abc_15497_new_n4616_));
OR2X2 OR2X2_1322 ( .A(_abc_15497_new_n4621_), .B(_abc_15497_new_n4622_), .Y(_abc_15497_new_n4623_));
OR2X2 OR2X2_1323 ( .A(_abc_15497_new_n3775_), .B(_abc_15497_new_n4623_), .Y(_abc_15497_new_n4624_));
OR2X2 OR2X2_1324 ( .A(_abc_15497_new_n4626_), .B(_abc_15497_new_n4617_), .Y(_abc_15497_new_n4627_));
OR2X2 OR2X2_1325 ( .A(_abc_15497_new_n4631_), .B(_abc_15497_new_n4630_), .Y(_abc_15497_new_n4632_));
OR2X2 OR2X2_1326 ( .A(_abc_15497_new_n3784_), .B(_abc_15497_new_n4632_), .Y(_abc_15497_new_n4633_));
OR2X2 OR2X2_1327 ( .A(_abc_15497_new_n4566_), .B(_abc_15497_new_n4561_), .Y(_abc_15497_new_n4637_));
OR2X2 OR2X2_1328 ( .A(e_reg_11_), .B(a_reg_6_), .Y(_abc_15497_new_n4639_));
OR2X2 OR2X2_1329 ( .A(_abc_15497_new_n4644_), .B(_abc_15497_new_n4645_), .Y(_abc_15497_new_n4646_));
OR2X2 OR2X2_133 ( .A(_abc_15497_new_n1103_), .B(digest_update), .Y(_abc_15497_new_n1104_));
OR2X2 OR2X2_1330 ( .A(_abc_15497_new_n4647_), .B(_abc_15497_new_n4637_), .Y(_abc_15497_new_n4650_));
OR2X2 OR2X2_1331 ( .A(_abc_15497_new_n4653_), .B(_abc_15497_new_n4648_), .Y(_abc_15497_new_n4654_));
OR2X2 OR2X2_1332 ( .A(_abc_15497_new_n4652_), .B(_abc_15497_new_n4655_), .Y(_abc_15497_new_n4656_));
OR2X2 OR2X2_1333 ( .A(_abc_15497_new_n4656_), .B(_abc_15497_new_n4614_), .Y(_abc_15497_new_n4657_));
OR2X2 OR2X2_1334 ( .A(_abc_15497_new_n4581_), .B(_abc_15497_new_n4569_), .Y(_abc_15497_new_n4658_));
OR2X2 OR2X2_1335 ( .A(_abc_15497_new_n4654_), .B(_abc_15497_new_n4635_), .Y(_abc_15497_new_n4659_));
OR2X2 OR2X2_1336 ( .A(_abc_15497_new_n4636_), .B(_abc_15497_new_n4651_), .Y(_abc_15497_new_n4660_));
OR2X2 OR2X2_1337 ( .A(_abc_15497_new_n4661_), .B(_abc_15497_new_n4658_), .Y(_abc_15497_new_n4662_));
OR2X2 OR2X2_1338 ( .A(_abc_15497_new_n4663_), .B(_abc_15497_new_n3773_), .Y(_abc_15497_new_n4664_));
OR2X2 OR2X2_1339 ( .A(_abc_15497_new_n4665_), .B(_abc_15497_new_n4666_), .Y(_abc_15497_new_n4667_));
OR2X2 OR2X2_134 ( .A(e_reg_7_), .B(\digest[7] ), .Y(_abc_15497_new_n1106_));
OR2X2 OR2X2_1340 ( .A(_abc_15497_new_n4667_), .B(_abc_15497_new_n3783_), .Y(_abc_15497_new_n4668_));
OR2X2 OR2X2_1341 ( .A(_abc_15497_new_n4672_), .B(_abc_15497_new_n4673_), .Y(_abc_15497_new_n4674_));
OR2X2 OR2X2_1342 ( .A(_abc_15497_new_n4675_), .B(_abc_15497_new_n4670_), .Y(_abc_15497_new_n4676_));
OR2X2 OR2X2_1343 ( .A(_abc_15497_new_n4612_), .B(_abc_15497_new_n4676_), .Y(_abc_15497_new_n4677_));
OR2X2 OR2X2_1344 ( .A(_abc_15497_new_n4678_), .B(_abc_15497_new_n4679_), .Y(_abc_15497_new_n4680_));
OR2X2 OR2X2_1345 ( .A(_abc_15497_new_n4683_), .B(_abc_15497_new_n4685_), .Y(_abc_15497_new_n4686_));
OR2X2 OR2X2_1346 ( .A(_abc_15497_new_n4682_), .B(_abc_15497_new_n4686_), .Y(_0a_reg_31_0__11_));
OR2X2 OR2X2_1347 ( .A(_abc_15497_new_n4599_), .B(_abc_15497_new_n4676_), .Y(_abc_15497_new_n4688_));
OR2X2 OR2X2_1348 ( .A(_abc_15497_new_n4688_), .B(_abc_15497_new_n4529_), .Y(_abc_15497_new_n4689_));
OR2X2 OR2X2_1349 ( .A(_abc_15497_new_n4611_), .B(_abc_15497_new_n4675_), .Y(_abc_15497_new_n4691_));
OR2X2 OR2X2_135 ( .A(_abc_15497_new_n1111_), .B(_abc_15497_new_n1091_), .Y(_abc_15497_new_n1112_));
OR2X2 OR2X2_1350 ( .A(_abc_15497_new_n4531_), .B(_abc_15497_new_n4688_), .Y(_abc_15497_new_n4695_));
OR2X2 OR2X2_1351 ( .A(_abc_15497_new_n4697_), .B(_abc_15497_new_n4694_), .Y(_abc_15497_new_n4698_));
OR2X2 OR2X2_1352 ( .A(b_reg_12_), .B(c_reg_12_), .Y(_abc_15497_new_n4702_));
OR2X2 OR2X2_1353 ( .A(_abc_15497_new_n4705_), .B(d_reg_12_), .Y(_abc_15497_new_n4706_));
OR2X2 OR2X2_1354 ( .A(_abc_15497_new_n4712_), .B(b_reg_12_), .Y(_abc_15497_new_n4713_));
OR2X2 OR2X2_1355 ( .A(_abc_15497_new_n3780_), .B(_abc_15497_new_n4714_), .Y(_abc_15497_new_n4715_));
OR2X2 OR2X2_1356 ( .A(_abc_15497_new_n4717_), .B(_abc_15497_new_n4716_), .Y(_abc_15497_new_n4718_));
OR2X2 OR2X2_1357 ( .A(_abc_15497_new_n3784_), .B(_abc_15497_new_n4718_), .Y(_abc_15497_new_n4719_));
OR2X2 OR2X2_1358 ( .A(_abc_15497_new_n4645_), .B(_abc_15497_new_n4640_), .Y(_abc_15497_new_n4723_));
OR2X2 OR2X2_1359 ( .A(e_reg_12_), .B(a_reg_7_), .Y(_abc_15497_new_n4725_));
OR2X2 OR2X2_136 ( .A(_abc_15497_new_n1114_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n1115_));
OR2X2 OR2X2_1360 ( .A(_abc_15497_new_n4730_), .B(_abc_15497_new_n4731_), .Y(_abc_15497_new_n4732_));
OR2X2 OR2X2_1361 ( .A(_abc_15497_new_n4733_), .B(_abc_15497_new_n4723_), .Y(_abc_15497_new_n4736_));
OR2X2 OR2X2_1362 ( .A(_abc_15497_new_n4722_), .B(_abc_15497_new_n4737_), .Y(_abc_15497_new_n4740_));
OR2X2 OR2X2_1363 ( .A(_abc_15497_new_n4701_), .B(_abc_15497_new_n4741_), .Y(_abc_15497_new_n4742_));
OR2X2 OR2X2_1364 ( .A(_abc_15497_new_n4747_), .B(_abc_15497_new_n4738_), .Y(_abc_15497_new_n4748_));
OR2X2 OR2X2_1365 ( .A(_abc_15497_new_n4749_), .B(_abc_15497_new_n4743_), .Y(_abc_15497_new_n4750_));
OR2X2 OR2X2_1366 ( .A(_abc_15497_new_n4746_), .B(_abc_15497_new_n4751_), .Y(_abc_15497_new_n4752_));
OR2X2 OR2X2_1367 ( .A(_abc_15497_new_n4750_), .B(_abc_15497_new_n3803_), .Y(_abc_15497_new_n4755_));
OR2X2 OR2X2_1368 ( .A(_abc_15497_new_n4745_), .B(_abc_15497_new_n3775_), .Y(_abc_15497_new_n4756_));
OR2X2 OR2X2_1369 ( .A(_abc_15497_new_n4753_), .B(_abc_15497_new_n4758_), .Y(_abc_15497_new_n4759_));
OR2X2 OR2X2_137 ( .A(_abc_15497_new_n1115_), .B(_abc_15497_new_n1110_), .Y(_abc_15497_new_n1116_));
OR2X2 OR2X2_1370 ( .A(_abc_15497_new_n4698_), .B(_abc_15497_new_n4760_), .Y(_abc_15497_new_n4761_));
OR2X2 OR2X2_1371 ( .A(_abc_15497_new_n4766_), .B(_abc_15497_new_n4768_), .Y(_abc_15497_new_n4769_));
OR2X2 OR2X2_1372 ( .A(_abc_15497_new_n4765_), .B(_abc_15497_new_n4769_), .Y(_0a_reg_31_0__12_));
OR2X2 OR2X2_1373 ( .A(_abc_15497_new_n4752_), .B(_abc_15497_new_n4699_), .Y(_abc_15497_new_n4771_));
OR2X2 OR2X2_1374 ( .A(_abc_15497_new_n4746_), .B(_abc_15497_new_n4743_), .Y(_abc_15497_new_n4773_));
OR2X2 OR2X2_1375 ( .A(_abc_15497_new_n4738_), .B(_abc_15497_new_n4734_), .Y(_abc_15497_new_n4774_));
OR2X2 OR2X2_1376 ( .A(b_reg_13_), .B(c_reg_13_), .Y(_abc_15497_new_n4775_));
OR2X2 OR2X2_1377 ( .A(_abc_15497_new_n4778_), .B(d_reg_13_), .Y(_abc_15497_new_n4779_));
OR2X2 OR2X2_1378 ( .A(_abc_15497_new_n4785_), .B(b_reg_13_), .Y(_abc_15497_new_n4786_));
OR2X2 OR2X2_1379 ( .A(_abc_15497_new_n3780_), .B(_abc_15497_new_n4787_), .Y(_abc_15497_new_n4788_));
OR2X2 OR2X2_138 ( .A(e_reg_8_), .B(\digest[8] ), .Y(_abc_15497_new_n1118_));
OR2X2 OR2X2_1380 ( .A(_abc_15497_new_n4790_), .B(_abc_15497_new_n4789_), .Y(_abc_15497_new_n4791_));
OR2X2 OR2X2_1381 ( .A(_abc_15497_new_n3784_), .B(_abc_15497_new_n4791_), .Y(_abc_15497_new_n4792_));
OR2X2 OR2X2_1382 ( .A(_abc_15497_new_n4731_), .B(_abc_15497_new_n4726_), .Y(_abc_15497_new_n4796_));
OR2X2 OR2X2_1383 ( .A(e_reg_13_), .B(a_reg_8_), .Y(_abc_15497_new_n4798_));
OR2X2 OR2X2_1384 ( .A(_abc_15497_new_n4803_), .B(_abc_15497_new_n4804_), .Y(_abc_15497_new_n4805_));
OR2X2 OR2X2_1385 ( .A(_abc_15497_new_n4806_), .B(_abc_15497_new_n4796_), .Y(_abc_15497_new_n4809_));
OR2X2 OR2X2_1386 ( .A(_abc_15497_new_n4795_), .B(_abc_15497_new_n4810_), .Y(_abc_15497_new_n4813_));
OR2X2 OR2X2_1387 ( .A(_abc_15497_new_n4814_), .B(_abc_15497_new_n4774_), .Y(_abc_15497_new_n4815_));
OR2X2 OR2X2_1388 ( .A(_abc_15497_new_n4818_), .B(_abc_15497_new_n3773_), .Y(_abc_15497_new_n4819_));
OR2X2 OR2X2_1389 ( .A(_abc_15497_new_n4821_), .B(_abc_15497_new_n4811_), .Y(_abc_15497_new_n4822_));
OR2X2 OR2X2_139 ( .A(_abc_15497_new_n1122_), .B(_abc_15497_new_n1107_), .Y(_abc_15497_new_n1123_));
OR2X2 OR2X2_1390 ( .A(_abc_15497_new_n4823_), .B(_abc_15497_new_n4816_), .Y(_abc_15497_new_n4824_));
OR2X2 OR2X2_1391 ( .A(_abc_15497_new_n4824_), .B(_abc_15497_new_n3783_), .Y(_abc_15497_new_n4825_));
OR2X2 OR2X2_1392 ( .A(_abc_15497_new_n4830_), .B(_abc_15497_new_n4829_), .Y(_abc_15497_new_n4831_));
OR2X2 OR2X2_1393 ( .A(_abc_15497_new_n4827_), .B(_abc_15497_new_n4832_), .Y(_abc_15497_new_n4833_));
OR2X2 OR2X2_1394 ( .A(_abc_15497_new_n4772_), .B(_abc_15497_new_n4833_), .Y(_abc_15497_new_n4834_));
OR2X2 OR2X2_1395 ( .A(_abc_15497_new_n4835_), .B(_abc_15497_new_n4836_), .Y(_abc_15497_new_n4837_));
OR2X2 OR2X2_1396 ( .A(_abc_15497_new_n4840_), .B(_abc_15497_new_n4841_), .Y(_abc_15497_new_n4842_));
OR2X2 OR2X2_1397 ( .A(_abc_15497_new_n4839_), .B(_abc_15497_new_n4842_), .Y(_0a_reg_31_0__13_));
OR2X2 OR2X2_1398 ( .A(_abc_15497_new_n4771_), .B(_abc_15497_new_n4832_), .Y(_abc_15497_new_n4845_));
OR2X2 OR2X2_1399 ( .A(_abc_15497_new_n4759_), .B(_abc_15497_new_n4833_), .Y(_abc_15497_new_n4848_));
OR2X2 OR2X2_14 ( .A(c_reg_15_), .B(\digest[79] ), .Y(_abc_15497_new_n760_));
OR2X2 OR2X2_140 ( .A(_abc_15497_new_n1123_), .B(_abc_15497_new_n1121_), .Y(_abc_15497_new_n1124_));
OR2X2 OR2X2_1400 ( .A(_abc_15497_new_n4850_), .B(_abc_15497_new_n4847_), .Y(_abc_15497_new_n4851_));
OR2X2 OR2X2_1401 ( .A(_abc_15497_new_n4830_), .B(_abc_15497_new_n4816_), .Y(_abc_15497_new_n4852_));
OR2X2 OR2X2_1402 ( .A(_abc_15497_new_n4811_), .B(_abc_15497_new_n4807_), .Y(_abc_15497_new_n4853_));
OR2X2 OR2X2_1403 ( .A(b_reg_14_), .B(c_reg_14_), .Y(_abc_15497_new_n4854_));
OR2X2 OR2X2_1404 ( .A(_abc_15497_new_n4857_), .B(d_reg_14_), .Y(_abc_15497_new_n4858_));
OR2X2 OR2X2_1405 ( .A(_abc_15497_new_n4864_), .B(b_reg_14_), .Y(_abc_15497_new_n4865_));
OR2X2 OR2X2_1406 ( .A(_abc_15497_new_n3780_), .B(_abc_15497_new_n4866_), .Y(_abc_15497_new_n4867_));
OR2X2 OR2X2_1407 ( .A(_abc_15497_new_n4804_), .B(_abc_15497_new_n4799_), .Y(_abc_15497_new_n4876_));
OR2X2 OR2X2_1408 ( .A(e_reg_14_), .B(a_reg_9_), .Y(_abc_15497_new_n4877_));
OR2X2 OR2X2_1409 ( .A(_abc_15497_new_n4880_), .B(w_14_), .Y(_abc_15497_new_n4881_));
OR2X2 OR2X2_141 ( .A(_abc_15497_new_n699_), .B(\digest[8] ), .Y(_abc_15497_new_n1129_));
OR2X2 OR2X2_1410 ( .A(_abc_15497_new_n4884_), .B(_abc_15497_new_n4876_), .Y(_abc_15497_new_n4887_));
OR2X2 OR2X2_1411 ( .A(_abc_15497_new_n4875_), .B(_abc_15497_new_n4888_), .Y(_abc_15497_new_n4891_));
OR2X2 OR2X2_1412 ( .A(_abc_15497_new_n4892_), .B(_abc_15497_new_n4853_), .Y(_abc_15497_new_n4893_));
OR2X2 OR2X2_1413 ( .A(_abc_15497_new_n4895_), .B(_abc_15497_new_n4889_), .Y(_abc_15497_new_n4896_));
OR2X2 OR2X2_1414 ( .A(_abc_15497_new_n4896_), .B(_abc_15497_new_n4894_), .Y(_abc_15497_new_n4897_));
OR2X2 OR2X2_1415 ( .A(_abc_15497_new_n4898_), .B(_abc_15497_new_n3784_), .Y(_abc_15497_new_n4899_));
OR2X2 OR2X2_1416 ( .A(_abc_15497_new_n4900_), .B(_abc_15497_new_n4901_), .Y(_abc_15497_new_n4902_));
OR2X2 OR2X2_1417 ( .A(_abc_15497_new_n4902_), .B(_abc_15497_new_n3774_), .Y(_abc_15497_new_n4903_));
OR2X2 OR2X2_1418 ( .A(_abc_15497_new_n4907_), .B(_abc_15497_new_n4908_), .Y(_abc_15497_new_n4909_));
OR2X2 OR2X2_1419 ( .A(_abc_15497_new_n4905_), .B(_abc_15497_new_n4910_), .Y(_abc_15497_new_n4911_));
OR2X2 OR2X2_142 ( .A(_abc_15497_new_n1128_), .B(_abc_15497_new_n1130_), .Y(_0H4_reg_31_0__8_));
OR2X2 OR2X2_1420 ( .A(_abc_15497_new_n4851_), .B(_abc_15497_new_n4912_), .Y(_abc_15497_new_n4913_));
OR2X2 OR2X2_1421 ( .A(_abc_15497_new_n4918_), .B(_abc_15497_new_n4920_), .Y(_abc_15497_new_n4921_));
OR2X2 OR2X2_1422 ( .A(_abc_15497_new_n4917_), .B(_abc_15497_new_n4921_), .Y(_0a_reg_31_0__14_));
OR2X2 OR2X2_1423 ( .A(_abc_15497_new_n4908_), .B(_abc_15497_new_n4901_), .Y(_abc_15497_new_n4925_));
OR2X2 OR2X2_1424 ( .A(_abc_15497_new_n4889_), .B(_abc_15497_new_n4885_), .Y(_abc_15497_new_n4926_));
OR2X2 OR2X2_1425 ( .A(b_reg_15_), .B(c_reg_15_), .Y(_abc_15497_new_n4927_));
OR2X2 OR2X2_1426 ( .A(_abc_15497_new_n4930_), .B(d_reg_15_), .Y(_abc_15497_new_n4931_));
OR2X2 OR2X2_1427 ( .A(_abc_15497_new_n4937_), .B(b_reg_15_), .Y(_abc_15497_new_n4938_));
OR2X2 OR2X2_1428 ( .A(_abc_15497_new_n3780_), .B(_abc_15497_new_n4939_), .Y(_abc_15497_new_n4940_));
OR2X2 OR2X2_1429 ( .A(_abc_15497_new_n4882_), .B(_abc_15497_new_n4878_), .Y(_abc_15497_new_n4949_));
OR2X2 OR2X2_143 ( .A(e_reg_9_), .B(\digest[9] ), .Y(_abc_15497_new_n1133_));
OR2X2 OR2X2_1430 ( .A(e_reg_15_), .B(a_reg_10_), .Y(_abc_15497_new_n4950_));
OR2X2 OR2X2_1431 ( .A(_abc_15497_new_n4953_), .B(w_15_), .Y(_abc_15497_new_n4954_));
OR2X2 OR2X2_1432 ( .A(_abc_15497_new_n4957_), .B(_abc_15497_new_n4949_), .Y(_abc_15497_new_n4960_));
OR2X2 OR2X2_1433 ( .A(_abc_15497_new_n4948_), .B(_abc_15497_new_n4961_), .Y(_abc_15497_new_n4964_));
OR2X2 OR2X2_1434 ( .A(_abc_15497_new_n4965_), .B(_abc_15497_new_n4926_), .Y(_abc_15497_new_n4966_));
OR2X2 OR2X2_1435 ( .A(_abc_15497_new_n4969_), .B(_abc_15497_new_n3780_), .Y(_abc_15497_new_n4970_));
OR2X2 OR2X2_1436 ( .A(_abc_15497_new_n4972_), .B(_abc_15497_new_n4962_), .Y(_abc_15497_new_n4973_));
OR2X2 OR2X2_1437 ( .A(_abc_15497_new_n4974_), .B(_abc_15497_new_n4967_), .Y(_abc_15497_new_n4975_));
OR2X2 OR2X2_1438 ( .A(_abc_15497_new_n4975_), .B(_abc_15497_new_n3753_), .Y(_abc_15497_new_n4976_));
OR2X2 OR2X2_1439 ( .A(_abc_15497_new_n4981_), .B(_abc_15497_new_n4980_), .Y(_abc_15497_new_n4982_));
OR2X2 OR2X2_144 ( .A(_abc_15497_new_n1136_), .B(_abc_15497_new_n1119_), .Y(_abc_15497_new_n1140_));
OR2X2 OR2X2_1440 ( .A(_abc_15497_new_n4983_), .B(_abc_15497_new_n4978_), .Y(_abc_15497_new_n4984_));
OR2X2 OR2X2_1441 ( .A(_abc_15497_new_n4924_), .B(_abc_15497_new_n4984_), .Y(_abc_15497_new_n4985_));
OR2X2 OR2X2_1442 ( .A(_abc_15497_new_n4986_), .B(_abc_15497_new_n4987_), .Y(_abc_15497_new_n4988_));
OR2X2 OR2X2_1443 ( .A(_abc_15497_new_n4991_), .B(_abc_15497_new_n4993_), .Y(_abc_15497_new_n4994_));
OR2X2 OR2X2_1444 ( .A(_abc_15497_new_n4990_), .B(_abc_15497_new_n4994_), .Y(_0a_reg_31_0__15_));
OR2X2 OR2X2_1445 ( .A(_abc_15497_new_n4984_), .B(_abc_15497_new_n4911_), .Y(_abc_15497_new_n4996_));
OR2X2 OR2X2_1446 ( .A(_abc_15497_new_n4848_), .B(_abc_15497_new_n4996_), .Y(_abc_15497_new_n4997_));
OR2X2 OR2X2_1447 ( .A(_abc_15497_new_n4693_), .B(_abc_15497_new_n4997_), .Y(_abc_15497_new_n4998_));
OR2X2 OR2X2_1448 ( .A(_abc_15497_new_n4996_), .B(_abc_15497_new_n4846_), .Y(_abc_15497_new_n4999_));
OR2X2 OR2X2_1449 ( .A(_abc_15497_new_n4923_), .B(_abc_15497_new_n4983_), .Y(_abc_15497_new_n5001_));
OR2X2 OR2X2_145 ( .A(_abc_15497_new_n1125_), .B(_abc_15497_new_n1140_), .Y(_abc_15497_new_n1141_));
OR2X2 OR2X2_1450 ( .A(_abc_15497_new_n4997_), .B(_abc_15497_new_n4695_), .Y(_abc_15497_new_n5005_));
OR2X2 OR2X2_1451 ( .A(_abc_15497_new_n4441_), .B(_abc_15497_new_n5005_), .Y(_abc_15497_new_n5006_));
OR2X2 OR2X2_1452 ( .A(d_reg_16_), .B(b_reg_16_), .Y(_abc_15497_new_n5014_));
OR2X2 OR2X2_1453 ( .A(_abc_15497_new_n5017_), .B(c_reg_16_), .Y(_abc_15497_new_n5020_));
OR2X2 OR2X2_1454 ( .A(_abc_15497_new_n5024_), .B(_abc_15497_new_n5026_), .Y(_abc_15497_new_n5027_));
OR2X2 OR2X2_1455 ( .A(_abc_15497_new_n3780_), .B(_abc_15497_new_n5027_), .Y(_abc_15497_new_n5028_));
OR2X2 OR2X2_1456 ( .A(_abc_15497_new_n5029_), .B(_abc_15497_new_n5015_), .Y(_abc_15497_new_n5030_));
OR2X2 OR2X2_1457 ( .A(e_reg_16_), .B(a_reg_11_), .Y(_abc_15497_new_n5038_));
OR2X2 OR2X2_1458 ( .A(_abc_15497_new_n5043_), .B(_abc_15497_new_n5044_), .Y(_abc_15497_new_n5045_));
OR2X2 OR2X2_1459 ( .A(_abc_15497_new_n5047_), .B(_abc_15497_new_n5048_), .Y(_abc_15497_new_n5049_));
OR2X2 OR2X2_146 ( .A(_abc_15497_new_n1146_), .B(_abc_15497_new_n1132_), .Y(_0H4_reg_31_0__9_));
OR2X2 OR2X2_1460 ( .A(_abc_15497_new_n5034_), .B(_abc_15497_new_n5049_), .Y(_abc_15497_new_n5050_));
OR2X2 OR2X2_1461 ( .A(_abc_15497_new_n5013_), .B(_abc_15497_new_n5053_), .Y(_abc_15497_new_n5054_));
OR2X2 OR2X2_1462 ( .A(_abc_15497_new_n5060_), .B(_abc_15497_new_n5058_), .Y(_abc_15497_new_n5061_));
OR2X2 OR2X2_1463 ( .A(_abc_15497_new_n5061_), .B(_abc_15497_new_n5009_), .Y(_abc_15497_new_n5063_));
OR2X2 OR2X2_1464 ( .A(_abc_15497_new_n5064_), .B(_abc_15497_new_n5062_), .Y(_abc_15497_new_n5065_));
OR2X2 OR2X2_1465 ( .A(_abc_15497_new_n5008_), .B(_abc_15497_new_n5066_), .Y(_abc_15497_new_n5067_));
OR2X2 OR2X2_1466 ( .A(_abc_15497_new_n5072_), .B(_abc_15497_new_n5073_), .Y(_abc_15497_new_n5074_));
OR2X2 OR2X2_1467 ( .A(_abc_15497_new_n5071_), .B(_abc_15497_new_n5074_), .Y(_0a_reg_31_0__16_));
OR2X2 OR2X2_1468 ( .A(b_reg_17_), .B(c_reg_17_), .Y(_abc_15497_new_n5083_));
OR2X2 OR2X2_1469 ( .A(_abc_15497_new_n5086_), .B(d_reg_17_), .Y(_abc_15497_new_n5087_));
OR2X2 OR2X2_147 ( .A(e_reg_10_), .B(\digest[10] ), .Y(_abc_15497_new_n1152_));
OR2X2 OR2X2_1470 ( .A(_abc_15497_new_n5093_), .B(b_reg_17_), .Y(_abc_15497_new_n5094_));
OR2X2 OR2X2_1471 ( .A(_abc_15497_new_n3780_), .B(_abc_15497_new_n5095_), .Y(_abc_15497_new_n5096_));
OR2X2 OR2X2_1472 ( .A(_abc_15497_new_n5098_), .B(_abc_15497_new_n5097_), .Y(_abc_15497_new_n5099_));
OR2X2 OR2X2_1473 ( .A(_abc_15497_new_n3784_), .B(_abc_15497_new_n5099_), .Y(_abc_15497_new_n5100_));
OR2X2 OR2X2_1474 ( .A(_abc_15497_new_n5044_), .B(_abc_15497_new_n5039_), .Y(_abc_15497_new_n5104_));
OR2X2 OR2X2_1475 ( .A(e_reg_17_), .B(a_reg_12_), .Y(_abc_15497_new_n5106_));
OR2X2 OR2X2_1476 ( .A(_abc_15497_new_n5111_), .B(_abc_15497_new_n5112_), .Y(_abc_15497_new_n5113_));
OR2X2 OR2X2_1477 ( .A(_abc_15497_new_n5114_), .B(_abc_15497_new_n5104_), .Y(_abc_15497_new_n5117_));
OR2X2 OR2X2_1478 ( .A(_abc_15497_new_n5103_), .B(_abc_15497_new_n5118_), .Y(_abc_15497_new_n5121_));
OR2X2 OR2X2_1479 ( .A(_abc_15497_new_n5123_), .B(_abc_15497_new_n5082_), .Y(_abc_15497_new_n5125_));
OR2X2 OR2X2_148 ( .A(_abc_15497_new_n1151_), .B(_abc_15497_new_n1155_), .Y(_abc_15497_new_n1156_));
OR2X2 OR2X2_1480 ( .A(_abc_15497_new_n5126_), .B(_abc_15497_new_n5124_), .Y(_abc_15497_new_n5127_));
OR2X2 OR2X2_1481 ( .A(_abc_15497_new_n5127_), .B(_abc_15497_new_n4059_), .Y(_abc_15497_new_n5128_));
OR2X2 OR2X2_1482 ( .A(_abc_15497_new_n5129_), .B(_abc_15497_new_n5130_), .Y(_abc_15497_new_n5131_));
OR2X2 OR2X2_1483 ( .A(_abc_15497_new_n5133_), .B(_abc_15497_new_n5134_), .Y(_abc_15497_new_n5135_));
OR2X2 OR2X2_1484 ( .A(_abc_15497_new_n5077_), .B(_abc_15497_new_n5136_), .Y(_abc_15497_new_n5137_));
OR2X2 OR2X2_1485 ( .A(_abc_15497_new_n5076_), .B(_abc_15497_new_n5135_), .Y(_abc_15497_new_n5138_));
OR2X2 OR2X2_1486 ( .A(_abc_15497_new_n5141_), .B(_abc_15497_new_n5143_), .Y(_abc_15497_new_n5144_));
OR2X2 OR2X2_1487 ( .A(_abc_15497_new_n5140_), .B(_abc_15497_new_n5144_), .Y(_0a_reg_31_0__17_));
OR2X2 OR2X2_1488 ( .A(_abc_15497_new_n5134_), .B(_abc_15497_new_n5063_), .Y(_abc_15497_new_n5148_));
OR2X2 OR2X2_1489 ( .A(_abc_15497_new_n5146_), .B(_abc_15497_new_n5150_), .Y(_abc_15497_new_n5151_));
OR2X2 OR2X2_149 ( .A(_abc_15497_new_n1160_), .B(_abc_15497_new_n1148_), .Y(_0H4_reg_31_0__10_));
OR2X2 OR2X2_1490 ( .A(d_reg_18_), .B(b_reg_18_), .Y(_abc_15497_new_n5156_));
OR2X2 OR2X2_1491 ( .A(_abc_15497_new_n5159_), .B(c_reg_18_), .Y(_abc_15497_new_n5162_));
OR2X2 OR2X2_1492 ( .A(_abc_15497_new_n5166_), .B(_abc_15497_new_n5168_), .Y(_abc_15497_new_n5169_));
OR2X2 OR2X2_1493 ( .A(_abc_15497_new_n3780_), .B(_abc_15497_new_n5169_), .Y(_abc_15497_new_n5170_));
OR2X2 OR2X2_1494 ( .A(_abc_15497_new_n5171_), .B(_abc_15497_new_n5157_), .Y(_abc_15497_new_n5172_));
OR2X2 OR2X2_1495 ( .A(_abc_15497_new_n5112_), .B(_abc_15497_new_n5107_), .Y(_abc_15497_new_n5177_));
OR2X2 OR2X2_1496 ( .A(e_reg_18_), .B(a_reg_13_), .Y(_abc_15497_new_n5179_));
OR2X2 OR2X2_1497 ( .A(_abc_15497_new_n5184_), .B(_abc_15497_new_n5185_), .Y(_abc_15497_new_n5186_));
OR2X2 OR2X2_1498 ( .A(_abc_15497_new_n5187_), .B(_abc_15497_new_n5177_), .Y(_abc_15497_new_n5190_));
OR2X2 OR2X2_1499 ( .A(_abc_15497_new_n5193_), .B(_abc_15497_new_n5195_), .Y(_abc_15497_new_n5196_));
OR2X2 OR2X2_15 ( .A(c_reg_14_), .B(\digest[78] ), .Y(_abc_15497_new_n764_));
OR2X2 OR2X2_150 ( .A(e_reg_11_), .B(\digest[11] ), .Y(_abc_15497_new_n1165_));
OR2X2 OR2X2_1500 ( .A(_abc_15497_new_n5198_), .B(_abc_15497_new_n5199_), .Y(_abc_15497_new_n5200_));
OR2X2 OR2X2_1501 ( .A(_abc_15497_new_n5202_), .B(_abc_15497_new_n5203_), .Y(_abc_15497_new_n5204_));
OR2X2 OR2X2_1502 ( .A(_abc_15497_new_n5151_), .B(_abc_15497_new_n5205_), .Y(_abc_15497_new_n5206_));
OR2X2 OR2X2_1503 ( .A(_abc_15497_new_n5211_), .B(_abc_15497_new_n5212_), .Y(_abc_15497_new_n5213_));
OR2X2 OR2X2_1504 ( .A(_abc_15497_new_n5210_), .B(_abc_15497_new_n5213_), .Y(_0a_reg_31_0__18_));
OR2X2 OR2X2_1505 ( .A(_abc_15497_new_n5195_), .B(_abc_15497_new_n5188_), .Y(_abc_15497_new_n5217_));
OR2X2 OR2X2_1506 ( .A(d_reg_19_), .B(b_reg_19_), .Y(_abc_15497_new_n5219_));
OR2X2 OR2X2_1507 ( .A(_abc_15497_new_n5222_), .B(c_reg_19_), .Y(_abc_15497_new_n5225_));
OR2X2 OR2X2_1508 ( .A(_abc_15497_new_n5229_), .B(_abc_15497_new_n5231_), .Y(_abc_15497_new_n5232_));
OR2X2 OR2X2_1509 ( .A(_abc_15497_new_n3780_), .B(_abc_15497_new_n5232_), .Y(_abc_15497_new_n5233_));
OR2X2 OR2X2_151 ( .A(_abc_15497_new_n1164_), .B(_abc_15497_new_n1168_), .Y(_abc_15497_new_n1169_));
OR2X2 OR2X2_1510 ( .A(_abc_15497_new_n5234_), .B(_abc_15497_new_n5220_), .Y(_abc_15497_new_n5235_));
OR2X2 OR2X2_1511 ( .A(_abc_15497_new_n5185_), .B(_abc_15497_new_n5180_), .Y(_abc_15497_new_n5241_));
OR2X2 OR2X2_1512 ( .A(e_reg_19_), .B(a_reg_14_), .Y(_abc_15497_new_n5243_));
OR2X2 OR2X2_1513 ( .A(_abc_15497_new_n5248_), .B(_abc_15497_new_n5249_), .Y(_abc_15497_new_n5250_));
OR2X2 OR2X2_1514 ( .A(_abc_15497_new_n5251_), .B(_abc_15497_new_n5241_), .Y(_abc_15497_new_n5254_));
OR2X2 OR2X2_1515 ( .A(_abc_15497_new_n5240_), .B(_abc_15497_new_n5255_), .Y(_abc_15497_new_n5258_));
OR2X2 OR2X2_1516 ( .A(_abc_15497_new_n5261_), .B(_abc_15497_new_n5262_), .Y(_abc_15497_new_n5263_));
OR2X2 OR2X2_1517 ( .A(_abc_15497_new_n5265_), .B(_abc_15497_new_n5266_), .Y(_abc_15497_new_n5267_));
OR2X2 OR2X2_1518 ( .A(_abc_15497_new_n5269_), .B(_abc_15497_new_n5271_), .Y(_abc_15497_new_n5272_));
OR2X2 OR2X2_1519 ( .A(_abc_15497_new_n5216_), .B(_abc_15497_new_n5272_), .Y(_abc_15497_new_n5273_));
OR2X2 OR2X2_152 ( .A(_abc_15497_new_n1163_), .B(_abc_15497_new_n1170_), .Y(_abc_15497_new_n1171_));
OR2X2 OR2X2_1520 ( .A(_abc_15497_new_n5274_), .B(_abc_15497_new_n5275_), .Y(_abc_15497_new_n5276_));
OR2X2 OR2X2_1521 ( .A(_abc_15497_new_n5279_), .B(_abc_15497_new_n5281_), .Y(_abc_15497_new_n5282_));
OR2X2 OR2X2_1522 ( .A(_abc_15497_new_n5278_), .B(_abc_15497_new_n5282_), .Y(_0a_reg_31_0__19_));
OR2X2 OR2X2_1523 ( .A(_abc_15497_new_n5204_), .B(_abc_15497_new_n5272_), .Y(_abc_15497_new_n5284_));
OR2X2 OR2X2_1524 ( .A(_abc_15497_new_n5149_), .B(_abc_15497_new_n5284_), .Y(_abc_15497_new_n5285_));
OR2X2 OR2X2_1525 ( .A(_abc_15497_new_n5202_), .B(_abc_15497_new_n5269_), .Y(_abc_15497_new_n5287_));
OR2X2 OR2X2_1526 ( .A(_abc_15497_new_n5135_), .B(_abc_15497_new_n5065_), .Y(_abc_15497_new_n5291_));
OR2X2 OR2X2_1527 ( .A(_abc_15497_new_n5291_), .B(_abc_15497_new_n5284_), .Y(_abc_15497_new_n5292_));
OR2X2 OR2X2_1528 ( .A(_abc_15497_new_n5007_), .B(_abc_15497_new_n5292_), .Y(_abc_15497_new_n5293_));
OR2X2 OR2X2_1529 ( .A(_abc_15497_new_n5256_), .B(_abc_15497_new_n5252_), .Y(_abc_15497_new_n5300_));
OR2X2 OR2X2_153 ( .A(_abc_15497_new_n1173_), .B(_abc_15497_new_n1162_), .Y(_0H4_reg_31_0__11_));
OR2X2 OR2X2_1530 ( .A(d_reg_20_), .B(b_reg_20_), .Y(_abc_15497_new_n5302_));
OR2X2 OR2X2_1531 ( .A(_abc_15497_new_n5305_), .B(c_reg_20_), .Y(_abc_15497_new_n5308_));
OR2X2 OR2X2_1532 ( .A(_abc_15497_new_n5312_), .B(_abc_15497_new_n5314_), .Y(_abc_15497_new_n5315_));
OR2X2 OR2X2_1533 ( .A(_abc_15497_new_n3780_), .B(_abc_15497_new_n5315_), .Y(_abc_15497_new_n5316_));
OR2X2 OR2X2_1534 ( .A(_abc_15497_new_n5317_), .B(_abc_15497_new_n5303_), .Y(_abc_15497_new_n5318_));
OR2X2 OR2X2_1535 ( .A(_abc_15497_new_n5249_), .B(_abc_15497_new_n5244_), .Y(_abc_15497_new_n5324_));
OR2X2 OR2X2_1536 ( .A(e_reg_20_), .B(a_reg_15_), .Y(_abc_15497_new_n5326_));
OR2X2 OR2X2_1537 ( .A(_abc_15497_new_n5331_), .B(_abc_15497_new_n5332_), .Y(_abc_15497_new_n5333_));
OR2X2 OR2X2_1538 ( .A(_abc_15497_new_n5334_), .B(_abc_15497_new_n5324_), .Y(_abc_15497_new_n5337_));
OR2X2 OR2X2_1539 ( .A(_abc_15497_new_n5323_), .B(_abc_15497_new_n5338_), .Y(_abc_15497_new_n5341_));
OR2X2 OR2X2_154 ( .A(_abc_15497_new_n1149_), .B(_abc_15497_new_n1177_), .Y(_abc_15497_new_n1178_));
OR2X2 OR2X2_1540 ( .A(_abc_15497_new_n5344_), .B(_abc_15497_new_n5345_), .Y(_abc_15497_new_n5346_));
OR2X2 OR2X2_1541 ( .A(_abc_15497_new_n5346_), .B(_abc_15497_new_n5010_), .Y(_abc_15497_new_n5347_));
OR2X2 OR2X2_1542 ( .A(_abc_15497_new_n5348_), .B(_abc_15497_new_n5349_), .Y(_abc_15497_new_n5350_));
OR2X2 OR2X2_1543 ( .A(_abc_15497_new_n5352_), .B(_abc_15497_new_n5353_), .Y(_abc_15497_new_n5354_));
OR2X2 OR2X2_1544 ( .A(_abc_15497_new_n5295_), .B(_abc_15497_new_n5355_), .Y(_abc_15497_new_n5356_));
OR2X2 OR2X2_1545 ( .A(_abc_15497_new_n5294_), .B(_abc_15497_new_n5354_), .Y(_abc_15497_new_n5357_));
OR2X2 OR2X2_1546 ( .A(_abc_15497_new_n5360_), .B(_abc_15497_new_n5362_), .Y(_abc_15497_new_n5363_));
OR2X2 OR2X2_1547 ( .A(_abc_15497_new_n5359_), .B(_abc_15497_new_n5363_), .Y(_0a_reg_31_0__20_));
OR2X2 OR2X2_1548 ( .A(_abc_15497_new_n5348_), .B(_abc_15497_new_n5345_), .Y(_abc_15497_new_n5368_));
OR2X2 OR2X2_1549 ( .A(_abc_15497_new_n5339_), .B(_abc_15497_new_n5335_), .Y(_abc_15497_new_n5369_));
OR2X2 OR2X2_155 ( .A(_abc_15497_new_n1179_), .B(_abc_15497_new_n1166_), .Y(_abc_15497_new_n1180_));
OR2X2 OR2X2_1550 ( .A(d_reg_21_), .B(b_reg_21_), .Y(_abc_15497_new_n5371_));
OR2X2 OR2X2_1551 ( .A(_abc_15497_new_n5374_), .B(c_reg_21_), .Y(_abc_15497_new_n5377_));
OR2X2 OR2X2_1552 ( .A(_abc_15497_new_n5381_), .B(_abc_15497_new_n5383_), .Y(_abc_15497_new_n5384_));
OR2X2 OR2X2_1553 ( .A(_abc_15497_new_n3780_), .B(_abc_15497_new_n5384_), .Y(_abc_15497_new_n5385_));
OR2X2 OR2X2_1554 ( .A(_abc_15497_new_n5386_), .B(_abc_15497_new_n5372_), .Y(_abc_15497_new_n5387_));
OR2X2 OR2X2_1555 ( .A(_abc_15497_new_n5332_), .B(_abc_15497_new_n5327_), .Y(_abc_15497_new_n5393_));
OR2X2 OR2X2_1556 ( .A(e_reg_21_), .B(a_reg_16_), .Y(_abc_15497_new_n5395_));
OR2X2 OR2X2_1557 ( .A(_abc_15497_new_n5400_), .B(_abc_15497_new_n5401_), .Y(_abc_15497_new_n5402_));
OR2X2 OR2X2_1558 ( .A(_abc_15497_new_n5403_), .B(_abc_15497_new_n5393_), .Y(_abc_15497_new_n5406_));
OR2X2 OR2X2_1559 ( .A(_abc_15497_new_n5392_), .B(_abc_15497_new_n5407_), .Y(_abc_15497_new_n5410_));
OR2X2 OR2X2_156 ( .A(_abc_15497_new_n1185_), .B(_abc_15497_new_n1183_), .Y(_abc_15497_new_n1186_));
OR2X2 OR2X2_1560 ( .A(_abc_15497_new_n5413_), .B(_abc_15497_new_n5414_), .Y(_abc_15497_new_n5415_));
OR2X2 OR2X2_1561 ( .A(_abc_15497_new_n5417_), .B(_abc_15497_new_n5418_), .Y(_abc_15497_new_n5419_));
OR2X2 OR2X2_1562 ( .A(_abc_15497_new_n5423_), .B(_abc_15497_new_n5421_), .Y(_abc_15497_new_n5424_));
OR2X2 OR2X2_1563 ( .A(_abc_15497_new_n5367_), .B(_abc_15497_new_n5425_), .Y(_abc_15497_new_n5426_));
OR2X2 OR2X2_1564 ( .A(_abc_15497_new_n5366_), .B(_abc_15497_new_n5424_), .Y(_abc_15497_new_n5427_));
OR2X2 OR2X2_1565 ( .A(_abc_15497_new_n5430_), .B(_abc_15497_new_n5432_), .Y(_abc_15497_new_n5433_));
OR2X2 OR2X2_1566 ( .A(_abc_15497_new_n5429_), .B(_abc_15497_new_n5433_), .Y(_0a_reg_31_0__21_));
OR2X2 OR2X2_1567 ( .A(_abc_15497_new_n5354_), .B(_abc_15497_new_n5424_), .Y(_abc_15497_new_n5435_));
OR2X2 OR2X2_1568 ( .A(_abc_15497_new_n5294_), .B(_abc_15497_new_n5435_), .Y(_abc_15497_new_n5436_));
OR2X2 OR2X2_1569 ( .A(_abc_15497_new_n5365_), .B(_abc_15497_new_n5423_), .Y(_abc_15497_new_n5438_));
OR2X2 OR2X2_157 ( .A(e_reg_12_), .B(\digest[12] ), .Y(_abc_15497_new_n1187_));
OR2X2 OR2X2_1570 ( .A(d_reg_22_), .B(b_reg_22_), .Y(_abc_15497_new_n5447_));
OR2X2 OR2X2_1571 ( .A(_abc_15497_new_n5450_), .B(c_reg_22_), .Y(_abc_15497_new_n5453_));
OR2X2 OR2X2_1572 ( .A(_abc_15497_new_n5457_), .B(_abc_15497_new_n5459_), .Y(_abc_15497_new_n5460_));
OR2X2 OR2X2_1573 ( .A(_abc_15497_new_n3780_), .B(_abc_15497_new_n5460_), .Y(_abc_15497_new_n5461_));
OR2X2 OR2X2_1574 ( .A(_abc_15497_new_n5462_), .B(_abc_15497_new_n5448_), .Y(_abc_15497_new_n5463_));
OR2X2 OR2X2_1575 ( .A(_abc_15497_new_n5401_), .B(_abc_15497_new_n5396_), .Y(_abc_15497_new_n5469_));
OR2X2 OR2X2_1576 ( .A(e_reg_22_), .B(a_reg_17_), .Y(_abc_15497_new_n5471_));
OR2X2 OR2X2_1577 ( .A(_abc_15497_new_n5476_), .B(_abc_15497_new_n5477_), .Y(_abc_15497_new_n5478_));
OR2X2 OR2X2_1578 ( .A(_abc_15497_new_n5479_), .B(_abc_15497_new_n5469_), .Y(_abc_15497_new_n5482_));
OR2X2 OR2X2_1579 ( .A(_abc_15497_new_n5468_), .B(_abc_15497_new_n5483_), .Y(_abc_15497_new_n5486_));
OR2X2 OR2X2_158 ( .A(_abc_15497_new_n1186_), .B(_abc_15497_new_n1190_), .Y(_abc_15497_new_n1191_));
OR2X2 OR2X2_1580 ( .A(_abc_15497_new_n5488_), .B(_abc_15497_new_n5446_), .Y(_abc_15497_new_n5490_));
OR2X2 OR2X2_1581 ( .A(_abc_15497_new_n5491_), .B(_abc_15497_new_n5489_), .Y(_abc_15497_new_n5492_));
OR2X2 OR2X2_1582 ( .A(_abc_15497_new_n5494_), .B(_abc_15497_new_n5495_), .Y(_abc_15497_new_n5496_));
OR2X2 OR2X2_1583 ( .A(_abc_15497_new_n5498_), .B(_abc_15497_new_n5499_), .Y(_abc_15497_new_n5500_));
OR2X2 OR2X2_1584 ( .A(_abc_15497_new_n5441_), .B(_abc_15497_new_n5501_), .Y(_abc_15497_new_n5502_));
OR2X2 OR2X2_1585 ( .A(_abc_15497_new_n5440_), .B(_abc_15497_new_n5500_), .Y(_abc_15497_new_n5503_));
OR2X2 OR2X2_1586 ( .A(_abc_15497_new_n5506_), .B(_abc_15497_new_n5507_), .Y(_abc_15497_new_n5508_));
OR2X2 OR2X2_1587 ( .A(_abc_15497_new_n5505_), .B(_abc_15497_new_n5508_), .Y(_0a_reg_31_0__22_));
OR2X2 OR2X2_1588 ( .A(_abc_15497_new_n5494_), .B(_abc_15497_new_n5491_), .Y(_abc_15497_new_n5513_));
OR2X2 OR2X2_1589 ( .A(b_reg_23_), .B(c_reg_23_), .Y(_abc_15497_new_n5515_));
OR2X2 OR2X2_159 ( .A(_abc_15497_new_n1195_), .B(_abc_15497_new_n1175_), .Y(_0H4_reg_31_0__12_));
OR2X2 OR2X2_1590 ( .A(_abc_15497_new_n5518_), .B(d_reg_23_), .Y(_abc_15497_new_n5519_));
OR2X2 OR2X2_1591 ( .A(_abc_15497_new_n5525_), .B(b_reg_23_), .Y(_abc_15497_new_n5526_));
OR2X2 OR2X2_1592 ( .A(_abc_15497_new_n3780_), .B(_abc_15497_new_n5527_), .Y(_abc_15497_new_n5528_));
OR2X2 OR2X2_1593 ( .A(_abc_15497_new_n5530_), .B(_abc_15497_new_n5529_), .Y(_abc_15497_new_n5531_));
OR2X2 OR2X2_1594 ( .A(_abc_15497_new_n3784_), .B(_abc_15497_new_n5531_), .Y(_abc_15497_new_n5532_));
OR2X2 OR2X2_1595 ( .A(_abc_15497_new_n5477_), .B(_abc_15497_new_n5472_), .Y(_abc_15497_new_n5536_));
OR2X2 OR2X2_1596 ( .A(e_reg_23_), .B(a_reg_18_), .Y(_abc_15497_new_n5538_));
OR2X2 OR2X2_1597 ( .A(_abc_15497_new_n5543_), .B(_abc_15497_new_n5544_), .Y(_abc_15497_new_n5545_));
OR2X2 OR2X2_1598 ( .A(_abc_15497_new_n5546_), .B(_abc_15497_new_n5536_), .Y(_abc_15497_new_n5549_));
OR2X2 OR2X2_1599 ( .A(_abc_15497_new_n5535_), .B(_abc_15497_new_n5550_), .Y(_abc_15497_new_n5553_));
OR2X2 OR2X2_16 ( .A(c_reg_13_), .B(\digest[77] ), .Y(_abc_15497_new_n771_));
OR2X2 OR2X2_160 ( .A(e_reg_13_), .B(\digest[13] ), .Y(_abc_15497_new_n1198_));
OR2X2 OR2X2_1600 ( .A(_abc_15497_new_n5555_), .B(_abc_15497_new_n5514_), .Y(_abc_15497_new_n5558_));
OR2X2 OR2X2_1601 ( .A(_abc_15497_new_n5559_), .B(_abc_15497_new_n3744_), .Y(_abc_15497_new_n5562_));
OR2X2 OR2X2_1602 ( .A(_abc_15497_new_n5567_), .B(_abc_15497_new_n5564_), .Y(_abc_15497_new_n5568_));
OR2X2 OR2X2_1603 ( .A(_abc_15497_new_n5512_), .B(_abc_15497_new_n5569_), .Y(_abc_15497_new_n5570_));
OR2X2 OR2X2_1604 ( .A(_abc_15497_new_n5511_), .B(_abc_15497_new_n5568_), .Y(_abc_15497_new_n5571_));
OR2X2 OR2X2_1605 ( .A(_abc_15497_new_n5574_), .B(_abc_15497_new_n5576_), .Y(_abc_15497_new_n5577_));
OR2X2 OR2X2_1606 ( .A(_abc_15497_new_n5573_), .B(_abc_15497_new_n5577_), .Y(_0a_reg_31_0__23_));
OR2X2 OR2X2_1607 ( .A(_abc_15497_new_n5500_), .B(_abc_15497_new_n5568_), .Y(_abc_15497_new_n5579_));
OR2X2 OR2X2_1608 ( .A(_abc_15497_new_n5579_), .B(_abc_15497_new_n5435_), .Y(_abc_15497_new_n5580_));
OR2X2 OR2X2_1609 ( .A(_abc_15497_new_n5290_), .B(_abc_15497_new_n5580_), .Y(_abc_15497_new_n5581_));
OR2X2 OR2X2_161 ( .A(_abc_15497_new_n1205_), .B(_abc_15497_new_n1202_), .Y(_abc_15497_new_n1206_));
OR2X2 OR2X2_1610 ( .A(_abc_15497_new_n5439_), .B(_abc_15497_new_n5579_), .Y(_abc_15497_new_n5582_));
OR2X2 OR2X2_1611 ( .A(_abc_15497_new_n5510_), .B(_abc_15497_new_n5567_), .Y(_abc_15497_new_n5584_));
OR2X2 OR2X2_1612 ( .A(_abc_15497_new_n5292_), .B(_abc_15497_new_n5580_), .Y(_abc_15497_new_n5588_));
OR2X2 OR2X2_1613 ( .A(_abc_15497_new_n5007_), .B(_abc_15497_new_n5588_), .Y(_abc_15497_new_n5589_));
OR2X2 OR2X2_1614 ( .A(b_reg_24_), .B(c_reg_24_), .Y(_abc_15497_new_n5595_));
OR2X2 OR2X2_1615 ( .A(_abc_15497_new_n5598_), .B(d_reg_24_), .Y(_abc_15497_new_n5599_));
OR2X2 OR2X2_1616 ( .A(_abc_15497_new_n5605_), .B(b_reg_24_), .Y(_abc_15497_new_n5606_));
OR2X2 OR2X2_1617 ( .A(_abc_15497_new_n3780_), .B(_abc_15497_new_n5607_), .Y(_abc_15497_new_n5608_));
OR2X2 OR2X2_1618 ( .A(_abc_15497_new_n5610_), .B(_abc_15497_new_n5609_), .Y(_abc_15497_new_n5611_));
OR2X2 OR2X2_1619 ( .A(_abc_15497_new_n3784_), .B(_abc_15497_new_n5611_), .Y(_abc_15497_new_n5612_));
OR2X2 OR2X2_162 ( .A(_abc_15497_new_n699_), .B(\digest[13] ), .Y(_abc_15497_new_n1208_));
OR2X2 OR2X2_1620 ( .A(_abc_15497_new_n5544_), .B(_abc_15497_new_n5539_), .Y(_abc_15497_new_n5616_));
OR2X2 OR2X2_1621 ( .A(e_reg_24_), .B(a_reg_19_), .Y(_abc_15497_new_n5618_));
OR2X2 OR2X2_1622 ( .A(_abc_15497_new_n5623_), .B(_abc_15497_new_n5624_), .Y(_abc_15497_new_n5625_));
OR2X2 OR2X2_1623 ( .A(_abc_15497_new_n5626_), .B(_abc_15497_new_n5616_), .Y(_abc_15497_new_n5629_));
OR2X2 OR2X2_1624 ( .A(_abc_15497_new_n5615_), .B(_abc_15497_new_n5630_), .Y(_abc_15497_new_n5633_));
OR2X2 OR2X2_1625 ( .A(_abc_15497_new_n5635_), .B(_abc_15497_new_n5594_), .Y(_abc_15497_new_n5637_));
OR2X2 OR2X2_1626 ( .A(_abc_15497_new_n5638_), .B(_abc_15497_new_n5636_), .Y(_abc_15497_new_n5639_));
OR2X2 OR2X2_1627 ( .A(_abc_15497_new_n5641_), .B(_abc_15497_new_n5642_), .Y(_abc_15497_new_n5643_));
OR2X2 OR2X2_1628 ( .A(_abc_15497_new_n5645_), .B(_abc_15497_new_n5646_), .Y(_abc_15497_new_n5647_));
OR2X2 OR2X2_1629 ( .A(_abc_15497_new_n5591_), .B(_abc_15497_new_n5648_), .Y(_abc_15497_new_n5649_));
OR2X2 OR2X2_163 ( .A(_abc_15497_new_n1207_), .B(_abc_15497_new_n1209_), .Y(_0H4_reg_31_0__13_));
OR2X2 OR2X2_1630 ( .A(_abc_15497_new_n5654_), .B(_abc_15497_new_n5655_), .Y(_abc_15497_new_n5656_));
OR2X2 OR2X2_1631 ( .A(_abc_15497_new_n5653_), .B(_abc_15497_new_n5656_), .Y(_0a_reg_31_0__24_));
OR2X2 OR2X2_1632 ( .A(_abc_15497_new_n5641_), .B(_abc_15497_new_n5638_), .Y(_abc_15497_new_n5660_));
OR2X2 OR2X2_1633 ( .A(b_reg_25_), .B(c_reg_25_), .Y(_abc_15497_new_n5663_));
OR2X2 OR2X2_1634 ( .A(_abc_15497_new_n5666_), .B(d_reg_25_), .Y(_abc_15497_new_n5667_));
OR2X2 OR2X2_1635 ( .A(_abc_15497_new_n5673_), .B(b_reg_25_), .Y(_abc_15497_new_n5674_));
OR2X2 OR2X2_1636 ( .A(_abc_15497_new_n3780_), .B(_abc_15497_new_n5675_), .Y(_abc_15497_new_n5676_));
OR2X2 OR2X2_1637 ( .A(_abc_15497_new_n5678_), .B(_abc_15497_new_n5677_), .Y(_abc_15497_new_n5679_));
OR2X2 OR2X2_1638 ( .A(_abc_15497_new_n3784_), .B(_abc_15497_new_n5679_), .Y(_abc_15497_new_n5680_));
OR2X2 OR2X2_1639 ( .A(_abc_15497_new_n5624_), .B(_abc_15497_new_n5619_), .Y(_abc_15497_new_n5684_));
OR2X2 OR2X2_164 ( .A(e_reg_14_), .B(\digest[14] ), .Y(_abc_15497_new_n1211_));
OR2X2 OR2X2_1640 ( .A(e_reg_25_), .B(a_reg_20_), .Y(_abc_15497_new_n5686_));
OR2X2 OR2X2_1641 ( .A(_abc_15497_new_n5691_), .B(_abc_15497_new_n5692_), .Y(_abc_15497_new_n5693_));
OR2X2 OR2X2_1642 ( .A(_abc_15497_new_n5694_), .B(_abc_15497_new_n5684_), .Y(_abc_15497_new_n5697_));
OR2X2 OR2X2_1643 ( .A(_abc_15497_new_n5683_), .B(_abc_15497_new_n5698_), .Y(_abc_15497_new_n5701_));
OR2X2 OR2X2_1644 ( .A(_abc_15497_new_n5703_), .B(_abc_15497_new_n5662_), .Y(_abc_15497_new_n5706_));
OR2X2 OR2X2_1645 ( .A(_abc_15497_new_n5661_), .B(_abc_15497_new_n5707_), .Y(_abc_15497_new_n5709_));
OR2X2 OR2X2_1646 ( .A(_abc_15497_new_n5710_), .B(_abc_15497_new_n5708_), .Y(_abc_15497_new_n5711_));
OR2X2 OR2X2_1647 ( .A(_abc_15497_new_n5659_), .B(_abc_15497_new_n5711_), .Y(_abc_15497_new_n5712_));
OR2X2 OR2X2_1648 ( .A(_abc_15497_new_n5713_), .B(_abc_15497_new_n5714_), .Y(_abc_15497_new_n5715_));
OR2X2 OR2X2_1649 ( .A(_abc_15497_new_n5718_), .B(_abc_15497_new_n5719_), .Y(_abc_15497_new_n5720_));
OR2X2 OR2X2_165 ( .A(_abc_15497_new_n1217_), .B(_abc_15497_new_n1215_), .Y(_abc_15497_new_n1218_));
OR2X2 OR2X2_1650 ( .A(_abc_15497_new_n5717_), .B(_abc_15497_new_n5720_), .Y(_0a_reg_31_0__25_));
OR2X2 OR2X2_1651 ( .A(_abc_15497_new_n5711_), .B(_abc_15497_new_n5658_), .Y(_abc_15497_new_n5722_));
OR2X2 OR2X2_1652 ( .A(_abc_15497_new_n5711_), .B(_abc_15497_new_n5647_), .Y(_abc_15497_new_n5724_));
OR2X2 OR2X2_1653 ( .A(c_reg_26_), .B(b_reg_26_), .Y(_abc_15497_new_n5733_));
OR2X2 OR2X2_1654 ( .A(_abc_15497_new_n5734_), .B(d_reg_26_), .Y(_abc_15497_new_n5737_));
OR2X2 OR2X2_1655 ( .A(_abc_15497_new_n5741_), .B(b_reg_26_), .Y(_abc_15497_new_n5742_));
OR2X2 OR2X2_1656 ( .A(_abc_15497_new_n3780_), .B(_abc_15497_new_n5743_), .Y(_abc_15497_new_n5744_));
OR2X2 OR2X2_1657 ( .A(_abc_15497_new_n5692_), .B(_abc_15497_new_n5687_), .Y(_abc_15497_new_n5753_));
OR2X2 OR2X2_1658 ( .A(e_reg_26_), .B(a_reg_21_), .Y(_abc_15497_new_n5755_));
OR2X2 OR2X2_1659 ( .A(_abc_15497_new_n5760_), .B(_abc_15497_new_n5761_), .Y(_abc_15497_new_n5762_));
OR2X2 OR2X2_166 ( .A(_abc_15497_new_n1219_), .B(_abc_15497_new_n1214_), .Y(_abc_15497_new_n1220_));
OR2X2 OR2X2_1660 ( .A(_abc_15497_new_n5763_), .B(_abc_15497_new_n5753_), .Y(_abc_15497_new_n5766_));
OR2X2 OR2X2_1661 ( .A(_abc_15497_new_n5752_), .B(_abc_15497_new_n5767_), .Y(_abc_15497_new_n5770_));
OR2X2 OR2X2_1662 ( .A(_abc_15497_new_n5772_), .B(_abc_15497_new_n5730_), .Y(_abc_15497_new_n5774_));
OR2X2 OR2X2_1663 ( .A(_abc_15497_new_n5775_), .B(_abc_15497_new_n5773_), .Y(_abc_15497_new_n5776_));
OR2X2 OR2X2_1664 ( .A(_abc_15497_new_n5778_), .B(_abc_15497_new_n5779_), .Y(_abc_15497_new_n5780_));
OR2X2 OR2X2_1665 ( .A(_abc_15497_new_n5782_), .B(_abc_15497_new_n5783_), .Y(_abc_15497_new_n5784_));
OR2X2 OR2X2_1666 ( .A(_abc_15497_new_n5729_), .B(_abc_15497_new_n5785_), .Y(_abc_15497_new_n5786_));
OR2X2 OR2X2_1667 ( .A(_abc_15497_new_n5791_), .B(_abc_15497_new_n5792_), .Y(_abc_15497_new_n5793_));
OR2X2 OR2X2_1668 ( .A(_abc_15497_new_n5790_), .B(_abc_15497_new_n5793_), .Y(_0a_reg_31_0__26_));
OR2X2 OR2X2_1669 ( .A(_abc_15497_new_n5787_), .B(_abc_15497_new_n5782_), .Y(_abc_15497_new_n5795_));
OR2X2 OR2X2_167 ( .A(_abc_15497_new_n699_), .B(\digest[14] ), .Y(_abc_15497_new_n1225_));
OR2X2 OR2X2_1670 ( .A(_abc_15497_new_n5778_), .B(_abc_15497_new_n5775_), .Y(_abc_15497_new_n5797_));
OR2X2 OR2X2_1671 ( .A(c_reg_27_), .B(b_reg_27_), .Y(_abc_15497_new_n5802_));
OR2X2 OR2X2_1672 ( .A(_abc_15497_new_n5803_), .B(d_reg_27_), .Y(_abc_15497_new_n5806_));
OR2X2 OR2X2_1673 ( .A(_abc_15497_new_n5810_), .B(b_reg_27_), .Y(_abc_15497_new_n5811_));
OR2X2 OR2X2_1674 ( .A(_abc_15497_new_n3780_), .B(_abc_15497_new_n5812_), .Y(_abc_15497_new_n5813_));
OR2X2 OR2X2_1675 ( .A(_abc_15497_new_n5761_), .B(_abc_15497_new_n5756_), .Y(_abc_15497_new_n5822_));
OR2X2 OR2X2_1676 ( .A(e_reg_27_), .B(a_reg_22_), .Y(_abc_15497_new_n5824_));
OR2X2 OR2X2_1677 ( .A(_abc_15497_new_n5829_), .B(_abc_15497_new_n5830_), .Y(_abc_15497_new_n5831_));
OR2X2 OR2X2_1678 ( .A(_abc_15497_new_n5832_), .B(_abc_15497_new_n5822_), .Y(_abc_15497_new_n5835_));
OR2X2 OR2X2_1679 ( .A(_abc_15497_new_n5821_), .B(_abc_15497_new_n5836_), .Y(_abc_15497_new_n5839_));
OR2X2 OR2X2_168 ( .A(_abc_15497_new_n1224_), .B(_abc_15497_new_n1226_), .Y(_0H4_reg_31_0__14_));
OR2X2 OR2X2_1680 ( .A(_abc_15497_new_n5841_), .B(_abc_15497_new_n5799_), .Y(_abc_15497_new_n5844_));
OR2X2 OR2X2_1681 ( .A(_abc_15497_new_n5798_), .B(_abc_15497_new_n5845_), .Y(_abc_15497_new_n5847_));
OR2X2 OR2X2_1682 ( .A(_abc_15497_new_n5848_), .B(_abc_15497_new_n5846_), .Y(_abc_15497_new_n5849_));
OR2X2 OR2X2_1683 ( .A(_abc_15497_new_n5796_), .B(_abc_15497_new_n5849_), .Y(_abc_15497_new_n5850_));
OR2X2 OR2X2_1684 ( .A(_abc_15497_new_n5795_), .B(_abc_15497_new_n5851_), .Y(_abc_15497_new_n5852_));
OR2X2 OR2X2_1685 ( .A(_abc_15497_new_n5855_), .B(_abc_15497_new_n5857_), .Y(_abc_15497_new_n5858_));
OR2X2 OR2X2_1686 ( .A(_abc_15497_new_n5854_), .B(_abc_15497_new_n5858_), .Y(_0a_reg_31_0__27_));
OR2X2 OR2X2_1687 ( .A(_abc_15497_new_n5590_), .B(_abc_15497_new_n5862_), .Y(_abc_15497_new_n5863_));
OR2X2 OR2X2_1688 ( .A(_abc_15497_new_n5864_), .B(_abc_15497_new_n5723_), .Y(_abc_15497_new_n5865_));
OR2X2 OR2X2_1689 ( .A(_abc_15497_new_n5866_), .B(_abc_15497_new_n5848_), .Y(_abc_15497_new_n5867_));
OR2X2 OR2X2_169 ( .A(e_reg_15_), .B(\digest[15] ), .Y(_abc_15497_new_n1229_));
OR2X2 OR2X2_1690 ( .A(c_reg_28_), .B(b_reg_28_), .Y(_abc_15497_new_n5875_));
OR2X2 OR2X2_1691 ( .A(_abc_15497_new_n5876_), .B(d_reg_28_), .Y(_abc_15497_new_n5879_));
OR2X2 OR2X2_1692 ( .A(_abc_15497_new_n5883_), .B(b_reg_28_), .Y(_abc_15497_new_n5884_));
OR2X2 OR2X2_1693 ( .A(_abc_15497_new_n3780_), .B(_abc_15497_new_n5885_), .Y(_abc_15497_new_n5886_));
OR2X2 OR2X2_1694 ( .A(_abc_15497_new_n5830_), .B(_abc_15497_new_n5825_), .Y(_abc_15497_new_n5895_));
OR2X2 OR2X2_1695 ( .A(e_reg_28_), .B(a_reg_23_), .Y(_abc_15497_new_n5897_));
OR2X2 OR2X2_1696 ( .A(_abc_15497_new_n5902_), .B(_abc_15497_new_n5903_), .Y(_abc_15497_new_n5904_));
OR2X2 OR2X2_1697 ( .A(_abc_15497_new_n5905_), .B(_abc_15497_new_n5895_), .Y(_abc_15497_new_n5908_));
OR2X2 OR2X2_1698 ( .A(_abc_15497_new_n5894_), .B(_abc_15497_new_n5909_), .Y(_abc_15497_new_n5912_));
OR2X2 OR2X2_1699 ( .A(_abc_15497_new_n5914_), .B(_abc_15497_new_n5872_), .Y(_abc_15497_new_n5916_));
OR2X2 OR2X2_17 ( .A(_abc_15497_new_n773_), .B(_abc_15497_new_n770_), .Y(_abc_15497_new_n774_));
OR2X2 OR2X2_170 ( .A(_abc_15497_new_n1236_), .B(_abc_15497_new_n1233_), .Y(_abc_15497_new_n1237_));
OR2X2 OR2X2_1700 ( .A(_abc_15497_new_n5917_), .B(_abc_15497_new_n5915_), .Y(_abc_15497_new_n5918_));
OR2X2 OR2X2_1701 ( .A(_abc_15497_new_n5920_), .B(_abc_15497_new_n5921_), .Y(_abc_15497_new_n5922_));
OR2X2 OR2X2_1702 ( .A(_abc_15497_new_n5922_), .B(_abc_15497_new_n5842_), .Y(_abc_15497_new_n5924_));
OR2X2 OR2X2_1703 ( .A(_abc_15497_new_n5925_), .B(_abc_15497_new_n5923_), .Y(_abc_15497_new_n5926_));
OR2X2 OR2X2_1704 ( .A(_abc_15497_new_n5871_), .B(_abc_15497_new_n5927_), .Y(_abc_15497_new_n5928_));
OR2X2 OR2X2_1705 ( .A(_abc_15497_new_n5933_), .B(_abc_15497_new_n5935_), .Y(_abc_15497_new_n5936_));
OR2X2 OR2X2_1706 ( .A(_abc_15497_new_n5932_), .B(_abc_15497_new_n5936_), .Y(_0a_reg_31_0__28_));
OR2X2 OR2X2_1707 ( .A(_abc_15497_new_n5920_), .B(_abc_15497_new_n5917_), .Y(_abc_15497_new_n5939_));
OR2X2 OR2X2_1708 ( .A(_abc_15497_new_n5944_), .B(_abc_15497_new_n5942_), .Y(_abc_15497_new_n5945_));
OR2X2 OR2X2_1709 ( .A(_abc_15497_new_n3780_), .B(_abc_15497_new_n5945_), .Y(_abc_15497_new_n5946_));
OR2X2 OR2X2_171 ( .A(_abc_15497_new_n699_), .B(\digest[15] ), .Y(_abc_15497_new_n1239_));
OR2X2 OR2X2_1710 ( .A(c_reg_29_), .B(b_reg_29_), .Y(_abc_15497_new_n5949_));
OR2X2 OR2X2_1711 ( .A(_abc_15497_new_n5950_), .B(_abc_15497_new_n5947_), .Y(_abc_15497_new_n5953_));
OR2X2 OR2X2_1712 ( .A(_abc_15497_new_n3775_), .B(_abc_15497_new_n5954_), .Y(_abc_15497_new_n5955_));
OR2X2 OR2X2_1713 ( .A(_abc_15497_new_n5959_), .B(_abc_15497_new_n3753_), .Y(_abc_15497_new_n5960_));
OR2X2 OR2X2_1714 ( .A(_abc_15497_new_n5903_), .B(_abc_15497_new_n5898_), .Y(_abc_15497_new_n5965_));
OR2X2 OR2X2_1715 ( .A(e_reg_29_), .B(a_reg_24_), .Y(_abc_15497_new_n5967_));
OR2X2 OR2X2_1716 ( .A(_abc_15497_new_n5972_), .B(_abc_15497_new_n5973_), .Y(_abc_15497_new_n5974_));
OR2X2 OR2X2_1717 ( .A(_abc_15497_new_n5975_), .B(_abc_15497_new_n5965_), .Y(_abc_15497_new_n5978_));
OR2X2 OR2X2_1718 ( .A(_abc_15497_new_n5964_), .B(_abc_15497_new_n5979_), .Y(_abc_15497_new_n5982_));
OR2X2 OR2X2_1719 ( .A(_abc_15497_new_n5984_), .B(_abc_15497_new_n5941_), .Y(_abc_15497_new_n5986_));
OR2X2 OR2X2_172 ( .A(_abc_15497_new_n1238_), .B(_abc_15497_new_n1240_), .Y(_0H4_reg_31_0__15_));
OR2X2 OR2X2_1720 ( .A(_abc_15497_new_n5987_), .B(_abc_15497_new_n5985_), .Y(_abc_15497_new_n5988_));
OR2X2 OR2X2_1721 ( .A(_abc_15497_new_n5988_), .B(_abc_15497_new_n4060_), .Y(_abc_15497_new_n5990_));
OR2X2 OR2X2_1722 ( .A(_abc_15497_new_n5991_), .B(_abc_15497_new_n5989_), .Y(_abc_15497_new_n5992_));
OR2X2 OR2X2_1723 ( .A(_abc_15497_new_n5992_), .B(_abc_15497_new_n5940_), .Y(_abc_15497_new_n5994_));
OR2X2 OR2X2_1724 ( .A(_abc_15497_new_n5995_), .B(_abc_15497_new_n5993_), .Y(_abc_15497_new_n5996_));
OR2X2 OR2X2_1725 ( .A(_abc_15497_new_n5938_), .B(_abc_15497_new_n5996_), .Y(_abc_15497_new_n5997_));
OR2X2 OR2X2_1726 ( .A(_abc_15497_new_n5998_), .B(_abc_15497_new_n5999_), .Y(_abc_15497_new_n6000_));
OR2X2 OR2X2_1727 ( .A(_abc_15497_new_n6003_), .B(_abc_15497_new_n6004_), .Y(_abc_15497_new_n6005_));
OR2X2 OR2X2_1728 ( .A(_abc_15497_new_n6002_), .B(_abc_15497_new_n6005_), .Y(_0a_reg_31_0__29_));
OR2X2 OR2X2_1729 ( .A(_abc_15497_new_n5870_), .B(_abc_15497_new_n6008_), .Y(_abc_15497_new_n6009_));
OR2X2 OR2X2_173 ( .A(_abc_15497_new_n1247_), .B(_abc_15497_new_n1230_), .Y(_abc_15497_new_n1248_));
OR2X2 OR2X2_1730 ( .A(_abc_15497_new_n6010_), .B(_abc_15497_new_n5995_), .Y(_abc_15497_new_n6011_));
OR2X2 OR2X2_1731 ( .A(_abc_15497_new_n6019_), .B(_abc_15497_new_n6017_), .Y(_abc_15497_new_n6020_));
OR2X2 OR2X2_1732 ( .A(_abc_15497_new_n3780_), .B(_abc_15497_new_n6020_), .Y(_abc_15497_new_n6021_));
OR2X2 OR2X2_1733 ( .A(c_reg_30_), .B(b_reg_30_), .Y(_abc_15497_new_n6024_));
OR2X2 OR2X2_1734 ( .A(_abc_15497_new_n6025_), .B(_abc_15497_new_n6022_), .Y(_abc_15497_new_n6028_));
OR2X2 OR2X2_1735 ( .A(_abc_15497_new_n3775_), .B(_abc_15497_new_n6029_), .Y(_abc_15497_new_n6030_));
OR2X2 OR2X2_1736 ( .A(_abc_15497_new_n6034_), .B(_abc_15497_new_n3753_), .Y(_abc_15497_new_n6035_));
OR2X2 OR2X2_1737 ( .A(_abc_15497_new_n5973_), .B(_abc_15497_new_n5968_), .Y(_abc_15497_new_n6040_));
OR2X2 OR2X2_1738 ( .A(e_reg_30_), .B(a_reg_25_), .Y(_abc_15497_new_n6042_));
OR2X2 OR2X2_1739 ( .A(_abc_15497_new_n6047_), .B(_abc_15497_new_n6048_), .Y(_abc_15497_new_n6049_));
OR2X2 OR2X2_174 ( .A(_abc_15497_new_n1216_), .B(_abc_15497_new_n1215_), .Y(_abc_15497_new_n1249_));
OR2X2 OR2X2_1740 ( .A(_abc_15497_new_n6050_), .B(_abc_15497_new_n6040_), .Y(_abc_15497_new_n6053_));
OR2X2 OR2X2_1741 ( .A(_abc_15497_new_n6039_), .B(_abc_15497_new_n6054_), .Y(_abc_15497_new_n6057_));
OR2X2 OR2X2_1742 ( .A(_abc_15497_new_n6059_), .B(_abc_15497_new_n6016_), .Y(_abc_15497_new_n6061_));
OR2X2 OR2X2_1743 ( .A(_abc_15497_new_n6062_), .B(_abc_15497_new_n6060_), .Y(_abc_15497_new_n6063_));
OR2X2 OR2X2_1744 ( .A(_abc_15497_new_n6065_), .B(_abc_15497_new_n6066_), .Y(_abc_15497_new_n6067_));
OR2X2 OR2X2_1745 ( .A(_abc_15497_new_n6067_), .B(_abc_15497_new_n6015_), .Y(_abc_15497_new_n6069_));
OR2X2 OR2X2_1746 ( .A(_abc_15497_new_n6070_), .B(_abc_15497_new_n6068_), .Y(_abc_15497_new_n6071_));
OR2X2 OR2X2_1747 ( .A(_abc_15497_new_n6014_), .B(_abc_15497_new_n6072_), .Y(_abc_15497_new_n6073_));
OR2X2 OR2X2_1748 ( .A(_abc_15497_new_n6013_), .B(_abc_15497_new_n6071_), .Y(_abc_15497_new_n6074_));
OR2X2 OR2X2_1749 ( .A(_abc_15497_new_n6077_), .B(_abc_15497_new_n6078_), .Y(_abc_15497_new_n6079_));
OR2X2 OR2X2_175 ( .A(_abc_15497_new_n1251_), .B(_abc_15497_new_n1248_), .Y(_abc_15497_new_n1252_));
OR2X2 OR2X2_1750 ( .A(_abc_15497_new_n6076_), .B(_abc_15497_new_n6079_), .Y(_0a_reg_31_0__30_));
OR2X2 OR2X2_1751 ( .A(_abc_15497_new_n6065_), .B(_abc_15497_new_n6062_), .Y(_abc_15497_new_n6083_));
OR2X2 OR2X2_1752 ( .A(_abc_15497_new_n6089_), .B(b_reg_31_), .Y(_abc_15497_new_n6090_));
OR2X2 OR2X2_1753 ( .A(_abc_15497_new_n6095_), .B(_abc_15497_new_n6089_), .Y(_abc_15497_new_n6098_));
OR2X2 OR2X2_1754 ( .A(_abc_15497_new_n3775_), .B(_abc_15497_new_n6099_), .Y(_abc_15497_new_n6100_));
OR2X2 OR2X2_1755 ( .A(_abc_15497_new_n6101_), .B(_abc_15497_new_n6093_), .Y(_abc_15497_new_n6102_));
OR2X2 OR2X2_1756 ( .A(_abc_15497_new_n3784_), .B(_abc_15497_new_n6102_), .Y(_abc_15497_new_n6103_));
OR2X2 OR2X2_1757 ( .A(_abc_15497_new_n6105_), .B(_abc_15497_new_n6092_), .Y(_abc_15497_new_n6106_));
OR2X2 OR2X2_1758 ( .A(_abc_15497_new_n6048_), .B(_abc_15497_new_n6043_), .Y(_abc_15497_new_n6108_));
OR2X2 OR2X2_1759 ( .A(e_reg_31_), .B(w_31_), .Y(_abc_15497_new_n6110_));
OR2X2 OR2X2_176 ( .A(_abc_15497_new_n1246_), .B(_abc_15497_new_n1252_), .Y(_abc_15497_new_n1253_));
OR2X2 OR2X2_1760 ( .A(_abc_15497_new_n6113_), .B(a_reg_26_), .Y(_abc_15497_new_n6116_));
OR2X2 OR2X2_1761 ( .A(_abc_15497_new_n6119_), .B(_abc_15497_new_n6120_), .Y(_abc_15497_new_n6121_));
OR2X2 OR2X2_1762 ( .A(_abc_15497_new_n6123_), .B(_abc_15497_new_n6124_), .Y(_abc_15497_new_n6125_));
OR2X2 OR2X2_1763 ( .A(_abc_15497_new_n6086_), .B(_abc_15497_new_n6125_), .Y(_abc_15497_new_n6128_));
OR2X2 OR2X2_1764 ( .A(_abc_15497_new_n6129_), .B(_abc_15497_new_n3769_), .Y(_abc_15497_new_n6130_));
OR2X2 OR2X2_1765 ( .A(_abc_15497_new_n6131_), .B(_abc_15497_new_n3744_), .Y(_abc_15497_new_n6132_));
OR2X2 OR2X2_1766 ( .A(_abc_15497_new_n6084_), .B(_abc_15497_new_n6133_), .Y(_abc_15497_new_n6136_));
OR2X2 OR2X2_1767 ( .A(_abc_15497_new_n6082_), .B(_abc_15497_new_n6137_), .Y(_abc_15497_new_n6138_));
OR2X2 OR2X2_1768 ( .A(_abc_15497_new_n6081_), .B(_abc_15497_new_n6139_), .Y(_abc_15497_new_n6140_));
OR2X2 OR2X2_1769 ( .A(_abc_15497_new_n6143_), .B(_abc_15497_new_n6145_), .Y(_abc_15497_new_n6146_));
OR2X2 OR2X2_177 ( .A(_abc_15497_new_n1255_), .B(_abc_15497_new_n1253_), .Y(_abc_15497_new_n1256_));
OR2X2 OR2X2_1770 ( .A(_abc_15497_new_n6142_), .B(_abc_15497_new_n6146_), .Y(_0a_reg_31_0__31_));
OR2X2 OR2X2_1771 ( .A(_abc_15497_new_n6155_), .B(_abc_15497_new_n6153_), .Y(_abc_15497_new_n6156_));
OR2X2 OR2X2_1772 ( .A(_abc_15497_new_n6157_), .B(digest_update), .Y(_abc_15497_abc_9717_auto_fsm_map_cc_170_map_fsm_844_0_));
OR2X2 OR2X2_1773 ( .A(_abc_15497_new_n6159_), .B(round_ctr_rst), .Y(_abc_15497_abc_9717_auto_fsm_map_cc_170_map_fsm_844_2_));
OR2X2 OR2X2_1774 ( .A(_abc_15497_new_n2010_), .B(_abc_15497_new_n6161_), .Y(_abc_15497_new_n6162_));
OR2X2 OR2X2_1775 ( .A(round_ctr_inc), .B(round_ctr_reg_0_), .Y(_abc_15497_new_n6163_));
OR2X2 OR2X2_1776 ( .A(round_ctr_reg_1_), .B(round_ctr_reg_0_), .Y(_abc_15497_new_n6167_));
OR2X2 OR2X2_1777 ( .A(_abc_15497_new_n6165_), .B(_abc_15497_new_n6169_), .Y(_0round_ctr_reg_6_0__1_));
OR2X2 OR2X2_1778 ( .A(_abc_15497_new_n6148_), .B(round_ctr_reg_2_), .Y(_abc_15497_new_n6174_));
OR2X2 OR2X2_1779 ( .A(_abc_15497_new_n6171_), .B(_abc_15497_new_n6176_), .Y(_0round_ctr_reg_6_0__2_));
OR2X2 OR2X2_178 ( .A(e_reg_16_), .B(\digest[16] ), .Y(_abc_15497_new_n1257_));
OR2X2 OR2X2_1780 ( .A(_abc_15497_new_n6179_), .B(_abc_15497_new_n6180_), .Y(_abc_15497_new_n6181_));
OR2X2 OR2X2_1781 ( .A(_abc_15497_new_n6185_), .B(_abc_15497_new_n6182_), .Y(_abc_15497_new_n6186_));
OR2X2 OR2X2_1782 ( .A(_abc_15497_new_n6190_), .B(_abc_15497_new_n6187_), .Y(_abc_15497_new_n6191_));
OR2X2 OR2X2_1783 ( .A(_abc_15497_new_n6196_), .B(_abc_15497_new_n3740_), .Y(_abc_15497_new_n6197_));
OR2X2 OR2X2_1784 ( .A(_abc_15497_new_n6193_), .B(round_ctr_reg_6_), .Y(_abc_15497_new_n6198_));
OR2X2 OR2X2_1785 ( .A(_abc_15497_new_n6200_), .B(digest_update), .Y(_0digest_valid_reg_0_0_));
OR2X2 OR2X2_1786 ( .A(c_reg_0_), .B(\digest[64] ), .Y(_abc_15497_new_n6202_));
OR2X2 OR2X2_1787 ( .A(_abc_15497_new_n6204_), .B(_abc_15497_new_n6205_), .Y(_0H2_reg_31_0__0_));
OR2X2 OR2X2_1788 ( .A(_abc_15497_new_n822_), .B(_abc_15497_new_n819_), .Y(_abc_15497_new_n6207_));
OR2X2 OR2X2_1789 ( .A(_abc_15497_new_n6208_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n6209_));
OR2X2 OR2X2_179 ( .A(_abc_15497_new_n1256_), .B(_abc_15497_new_n1260_), .Y(_abc_15497_new_n1261_));
OR2X2 OR2X2_1790 ( .A(_abc_15497_new_n3556_), .B(digest_update), .Y(_abc_15497_new_n6210_));
OR2X2 OR2X2_1791 ( .A(_abc_15497_new_n824_), .B(_abc_15497_new_n827_), .Y(_abc_15497_new_n6212_));
OR2X2 OR2X2_1792 ( .A(_abc_15497_new_n6213_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n6214_));
OR2X2 OR2X2_1793 ( .A(_abc_15497_new_n3562_), .B(digest_update), .Y(_abc_15497_new_n6215_));
OR2X2 OR2X2_1794 ( .A(_abc_15497_new_n829_), .B(_abc_15497_new_n6217_), .Y(_abc_15497_new_n6218_));
OR2X2 OR2X2_1795 ( .A(_abc_15497_new_n955_), .B(_abc_15497_new_n6219_), .Y(_abc_15497_new_n6220_));
OR2X2 OR2X2_1796 ( .A(_abc_15497_new_n6222_), .B(_abc_15497_new_n6223_), .Y(_0H2_reg_31_0__3_));
OR2X2 OR2X2_1797 ( .A(_abc_15497_new_n831_), .B(_abc_15497_new_n834_), .Y(_abc_15497_new_n6225_));
OR2X2 OR2X2_1798 ( .A(_abc_15497_new_n6226_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n6227_));
OR2X2 OR2X2_1799 ( .A(_abc_15497_new_n3574_), .B(digest_update), .Y(_abc_15497_new_n6228_));
OR2X2 OR2X2_18 ( .A(_abc_15497_new_n778_), .B(_abc_15497_new_n758_), .Y(_abc_15497_new_n779_));
OR2X2 OR2X2_180 ( .A(_abc_15497_new_n1265_), .B(_abc_15497_new_n1242_), .Y(_0H4_reg_31_0__16_));
OR2X2 OR2X2_1800 ( .A(_abc_15497_new_n3580_), .B(digest_update), .Y(_abc_15497_new_n6230_));
OR2X2 OR2X2_1801 ( .A(_abc_15497_new_n6234_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n6235_));
OR2X2 OR2X2_1802 ( .A(_abc_15497_new_n6235_), .B(_abc_15497_new_n6232_), .Y(_abc_15497_new_n6236_));
OR2X2 OR2X2_1803 ( .A(_abc_15497_new_n838_), .B(_abc_15497_new_n810_), .Y(_abc_15497_new_n6238_));
OR2X2 OR2X2_1804 ( .A(_abc_15497_new_n6242_), .B(_abc_15497_new_n6243_), .Y(_0H2_reg_31_0__6_));
OR2X2 OR2X2_1805 ( .A(_abc_15497_new_n6246_), .B(_abc_15497_new_n807_), .Y(_abc_15497_new_n6247_));
OR2X2 OR2X2_1806 ( .A(_abc_15497_new_n6245_), .B(_abc_15497_new_n6248_), .Y(_abc_15497_new_n6249_));
OR2X2 OR2X2_1807 ( .A(_abc_15497_new_n6251_), .B(_abc_15497_new_n6252_), .Y(_0H2_reg_31_0__7_));
OR2X2 OR2X2_1808 ( .A(_abc_15497_new_n840_), .B(_abc_15497_new_n845_), .Y(_abc_15497_new_n6255_));
OR2X2 OR2X2_1809 ( .A(_abc_15497_new_n6259_), .B(_abc_15497_new_n6254_), .Y(_0H2_reg_31_0__8_));
OR2X2 OR2X2_181 ( .A(e_reg_17_), .B(\digest[17] ), .Y(_abc_15497_new_n1269_));
OR2X2 OR2X2_1810 ( .A(_abc_15497_new_n6263_), .B(_abc_15497_new_n842_), .Y(_abc_15497_new_n6264_));
OR2X2 OR2X2_1811 ( .A(_abc_15497_new_n6262_), .B(_abc_15497_new_n6265_), .Y(_abc_15497_new_n6266_));
OR2X2 OR2X2_1812 ( .A(_abc_15497_new_n6268_), .B(_abc_15497_new_n6261_), .Y(_0H2_reg_31_0__9_));
OR2X2 OR2X2_1813 ( .A(_abc_15497_new_n848_), .B(_abc_15497_new_n794_), .Y(_abc_15497_new_n6270_));
OR2X2 OR2X2_1814 ( .A(_abc_15497_new_n6274_), .B(_abc_15497_new_n6275_), .Y(_0H2_reg_31_0__10_));
OR2X2 OR2X2_1815 ( .A(_abc_15497_new_n6278_), .B(_abc_15497_new_n791_), .Y(_abc_15497_new_n6279_));
OR2X2 OR2X2_1816 ( .A(_abc_15497_new_n6277_), .B(_abc_15497_new_n6280_), .Y(_abc_15497_new_n6281_));
OR2X2 OR2X2_1817 ( .A(_abc_15497_new_n6283_), .B(_abc_15497_new_n6284_), .Y(_0H2_reg_31_0__11_));
OR2X2 OR2X2_1818 ( .A(_abc_15497_new_n850_), .B(_abc_15497_new_n782_), .Y(_abc_15497_new_n6286_));
OR2X2 OR2X2_1819 ( .A(_abc_15497_new_n6290_), .B(_abc_15497_new_n6291_), .Y(_0H2_reg_31_0__12_));
OR2X2 OR2X2_182 ( .A(_abc_15497_new_n1268_), .B(_abc_15497_new_n1272_), .Y(_abc_15497_new_n1273_));
OR2X2 OR2X2_1820 ( .A(_abc_15497_new_n6295_), .B(_abc_15497_new_n772_), .Y(_abc_15497_new_n6296_));
OR2X2 OR2X2_1821 ( .A(_abc_15497_new_n6294_), .B(_abc_15497_new_n773_), .Y(_abc_15497_new_n6297_));
OR2X2 OR2X2_1822 ( .A(_abc_15497_new_n6299_), .B(_abc_15497_new_n6293_), .Y(_0H2_reg_31_0__13_));
OR2X2 OR2X2_1823 ( .A(_abc_15497_new_n6301_), .B(_abc_15497_new_n776_), .Y(_abc_15497_new_n6302_));
OR2X2 OR2X2_1824 ( .A(_abc_15497_new_n6302_), .B(_abc_15497_new_n765_), .Y(_abc_15497_new_n6303_));
OR2X2 OR2X2_1825 ( .A(_abc_15497_new_n6307_), .B(_abc_15497_new_n6308_), .Y(_0H2_reg_31_0__14_));
OR2X2 OR2X2_1826 ( .A(_abc_15497_new_n6311_), .B(_abc_15497_new_n761_), .Y(_abc_15497_new_n6312_));
OR2X2 OR2X2_1827 ( .A(_abc_15497_new_n6310_), .B(_abc_15497_new_n6313_), .Y(_abc_15497_new_n6314_));
OR2X2 OR2X2_1828 ( .A(_abc_15497_new_n6316_), .B(_abc_15497_new_n6317_), .Y(_0H2_reg_31_0__15_));
OR2X2 OR2X2_1829 ( .A(_abc_15497_new_n852_), .B(_abc_15497_new_n854_), .Y(_abc_15497_new_n6320_));
OR2X2 OR2X2_183 ( .A(_abc_15497_new_n1267_), .B(_abc_15497_new_n1274_), .Y(_abc_15497_new_n1275_));
OR2X2 OR2X2_1830 ( .A(_abc_15497_new_n6324_), .B(_abc_15497_new_n6319_), .Y(_0H2_reg_31_0__16_));
OR2X2 OR2X2_1831 ( .A(_abc_15497_new_n6327_), .B(_abc_15497_new_n743_), .Y(_abc_15497_new_n6328_));
OR2X2 OR2X2_1832 ( .A(_abc_15497_new_n6326_), .B(_abc_15497_new_n744_), .Y(_abc_15497_new_n6329_));
OR2X2 OR2X2_1833 ( .A(_abc_15497_new_n6331_), .B(_abc_15497_new_n6332_), .Y(_0H2_reg_31_0__17_));
OR2X2 OR2X2_1834 ( .A(_abc_15497_new_n6335_), .B(_abc_15497_new_n749_), .Y(_abc_15497_new_n6336_));
OR2X2 OR2X2_1835 ( .A(_abc_15497_new_n6336_), .B(_abc_15497_new_n738_), .Y(_abc_15497_new_n6337_));
OR2X2 OR2X2_1836 ( .A(_abc_15497_new_n6341_), .B(_abc_15497_new_n6334_), .Y(_0H2_reg_31_0__18_));
OR2X2 OR2X2_1837 ( .A(_abc_15497_new_n6347_), .B(_abc_15497_new_n6344_), .Y(_abc_15497_new_n6348_));
OR2X2 OR2X2_1838 ( .A(_abc_15497_new_n6349_), .B(_abc_15497_new_n6350_), .Y(_0H2_reg_31_0__19_));
OR2X2 OR2X2_1839 ( .A(_abc_15497_new_n6352_), .B(_abc_15497_new_n753_), .Y(_abc_15497_new_n6353_));
OR2X2 OR2X2_184 ( .A(_abc_15497_new_n699_), .B(\digest[17] ), .Y(_abc_15497_new_n1278_));
OR2X2 OR2X2_1840 ( .A(_abc_15497_new_n6353_), .B(_abc_15497_new_n728_), .Y(_abc_15497_new_n6354_));
OR2X2 OR2X2_1841 ( .A(_abc_15497_new_n6358_), .B(_abc_15497_new_n6359_), .Y(_0H2_reg_31_0__20_));
OR2X2 OR2X2_1842 ( .A(_abc_15497_new_n3676_), .B(digest_update), .Y(_abc_15497_new_n6361_));
OR2X2 OR2X2_1843 ( .A(_abc_15497_new_n6355_), .B(_abc_15497_new_n715_), .Y(_abc_15497_new_n6362_));
OR2X2 OR2X2_1844 ( .A(_abc_15497_new_n6365_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n6366_));
OR2X2 OR2X2_1845 ( .A(_abc_15497_new_n6366_), .B(_abc_15497_new_n6364_), .Y(_abc_15497_new_n6367_));
OR2X2 OR2X2_1846 ( .A(_abc_15497_new_n6370_), .B(_abc_15497_new_n713_), .Y(_abc_15497_new_n6371_));
OR2X2 OR2X2_1847 ( .A(_abc_15497_new_n6371_), .B(_abc_15497_new_n710_), .Y(_abc_15497_new_n6372_));
OR2X2 OR2X2_1848 ( .A(_abc_15497_new_n6376_), .B(_abc_15497_new_n6369_), .Y(_0H2_reg_31_0__22_));
OR2X2 OR2X2_1849 ( .A(_abc_15497_new_n6373_), .B(_abc_15497_new_n707_), .Y(_abc_15497_new_n6378_));
OR2X2 OR2X2_185 ( .A(_abc_15497_new_n1277_), .B(_abc_15497_new_n1279_), .Y(_0H4_reg_31_0__17_));
OR2X2 OR2X2_1850 ( .A(_abc_15497_new_n6382_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n6383_));
OR2X2 OR2X2_1851 ( .A(_abc_15497_new_n6383_), .B(_abc_15497_new_n6380_), .Y(_abc_15497_new_n6384_));
OR2X2 OR2X2_1852 ( .A(_abc_15497_new_n3688_), .B(digest_update), .Y(_abc_15497_new_n6385_));
OR2X2 OR2X2_1853 ( .A(_abc_15497_new_n859_), .B(_abc_15497_new_n867_), .Y(_abc_15497_new_n6388_));
OR2X2 OR2X2_1854 ( .A(_abc_15497_new_n6392_), .B(_abc_15497_new_n6387_), .Y(_0H2_reg_31_0__24_));
OR2X2 OR2X2_1855 ( .A(_abc_15497_new_n6396_), .B(_abc_15497_new_n863_), .Y(_abc_15497_new_n6397_));
OR2X2 OR2X2_1856 ( .A(_abc_15497_new_n6395_), .B(_abc_15497_new_n6398_), .Y(_abc_15497_new_n6399_));
OR2X2 OR2X2_1857 ( .A(_abc_15497_new_n6401_), .B(_abc_15497_new_n6394_), .Y(_0H2_reg_31_0__25_));
OR2X2 OR2X2_1858 ( .A(w_mem_inst_w_ctr_reg_4_), .B(w_mem_inst_w_ctr_reg_5_), .Y(w_mem_inst__abc_21203_new_n1585_));
OR2X2 OR2X2_1859 ( .A(w_mem_inst__abc_21203_new_n1585_), .B(w_mem_inst_w_ctr_reg_6_), .Y(w_mem_inst__abc_21203_new_n1586_));
OR2X2 OR2X2_186 ( .A(e_reg_18_), .B(\digest[18] ), .Y(_abc_15497_new_n1282_));
OR2X2 OR2X2_1860 ( .A(w_mem_inst__abc_21203_new_n1588_), .B(w_mem_inst_w_mem_13__31_), .Y(w_mem_inst__abc_21203_new_n1589_));
OR2X2 OR2X2_1861 ( .A(w_mem_inst__abc_21203_new_n1590_), .B(w_mem_inst_w_mem_8__31_), .Y(w_mem_inst__abc_21203_new_n1591_));
OR2X2 OR2X2_1862 ( .A(w_mem_inst_w_mem_2__31_), .B(w_mem_inst_w_mem_0__31_), .Y(w_mem_inst__abc_21203_new_n1594_));
OR2X2 OR2X2_1863 ( .A(w_mem_inst__abc_21203_new_n1593_), .B(w_mem_inst__abc_21203_new_n1597_), .Y(w_mem_inst__abc_21203_new_n1598_));
OR2X2 OR2X2_1864 ( .A(w_mem_inst__abc_21203_new_n1599_), .B(w_mem_inst__abc_21203_new_n1592_), .Y(w_mem_inst__abc_21203_new_n1600_));
OR2X2 OR2X2_1865 ( .A(w_mem_inst__abc_21203_new_n1601_), .B(w_mem_inst__abc_21203_new_n1587_), .Y(w_mem_inst__abc_21203_new_n1602_));
OR2X2 OR2X2_1866 ( .A(w_mem_inst__abc_21203_new_n1608_), .B(w_mem_inst__abc_21203_new_n1586_), .Y(w_mem_inst__abc_21203_new_n1609_));
OR2X2 OR2X2_1867 ( .A(w_mem_inst__abc_21203_new_n1615_), .B(w_mem_inst__abc_21203_new_n1618_), .Y(w_mem_inst__abc_21203_new_n1619_));
OR2X2 OR2X2_1868 ( .A(w_mem_inst__abc_21203_new_n1619_), .B(w_mem_inst__abc_21203_new_n1609_), .Y(w_mem_inst__abc_21203_new_n1620_));
OR2X2 OR2X2_1869 ( .A(w_mem_inst__abc_21203_new_n1622_), .B(w_mem_inst__abc_21203_new_n1625_), .Y(w_mem_inst__abc_21203_new_n1626_));
OR2X2 OR2X2_187 ( .A(_abc_15497_new_n1288_), .B(_abc_15497_new_n1286_), .Y(_abc_15497_new_n1289_));
OR2X2 OR2X2_1870 ( .A(w_mem_inst__abc_21203_new_n1620_), .B(w_mem_inst__abc_21203_new_n1626_), .Y(w_mem_inst__abc_21203_new_n1627_));
OR2X2 OR2X2_1871 ( .A(w_mem_inst__abc_21203_new_n1632_), .B(w_mem_inst__abc_21203_new_n1634_), .Y(w_mem_inst__abc_21203_new_n1635_));
OR2X2 OR2X2_1872 ( .A(w_mem_inst__abc_21203_new_n1635_), .B(w_mem_inst__abc_21203_new_n1629_), .Y(w_mem_inst__abc_21203_new_n1636_));
OR2X2 OR2X2_1873 ( .A(w_mem_inst__abc_21203_new_n1638_), .B(w_mem_inst__abc_21203_new_n1641_), .Y(w_mem_inst__abc_21203_new_n1642_));
OR2X2 OR2X2_1874 ( .A(w_mem_inst__abc_21203_new_n1644_), .B(w_mem_inst__abc_21203_new_n1646_), .Y(w_mem_inst__abc_21203_new_n1647_));
OR2X2 OR2X2_1875 ( .A(w_mem_inst__abc_21203_new_n1642_), .B(w_mem_inst__abc_21203_new_n1647_), .Y(w_mem_inst__abc_21203_new_n1648_));
OR2X2 OR2X2_1876 ( .A(w_mem_inst__abc_21203_new_n1650_), .B(w_mem_inst__abc_21203_new_n1652_), .Y(w_mem_inst__abc_21203_new_n1653_));
OR2X2 OR2X2_1877 ( .A(w_mem_inst__abc_21203_new_n1655_), .B(w_mem_inst__abc_21203_new_n1657_), .Y(w_mem_inst__abc_21203_new_n1658_));
OR2X2 OR2X2_1878 ( .A(w_mem_inst__abc_21203_new_n1653_), .B(w_mem_inst__abc_21203_new_n1658_), .Y(w_mem_inst__abc_21203_new_n1659_));
OR2X2 OR2X2_1879 ( .A(w_mem_inst__abc_21203_new_n1648_), .B(w_mem_inst__abc_21203_new_n1659_), .Y(w_mem_inst__abc_21203_new_n1660_));
OR2X2 OR2X2_188 ( .A(_abc_15497_new_n1290_), .B(_abc_15497_new_n1285_), .Y(_abc_15497_new_n1291_));
OR2X2 OR2X2_1880 ( .A(w_mem_inst__abc_21203_new_n1660_), .B(w_mem_inst__abc_21203_new_n1636_), .Y(w_mem_inst__abc_21203_new_n1661_));
OR2X2 OR2X2_1881 ( .A(w_mem_inst__abc_21203_new_n1661_), .B(w_mem_inst__abc_21203_new_n1627_), .Y(w_mem_inst__abc_21203_new_n1662_));
OR2X2 OR2X2_1882 ( .A(w_mem_inst__abc_21203_new_n1664_), .B(w_mem_inst_w_mem_8__0_), .Y(w_mem_inst__abc_21203_new_n1665_));
OR2X2 OR2X2_1883 ( .A(w_mem_inst__abc_21203_new_n1666_), .B(w_mem_inst_w_mem_13__0_), .Y(w_mem_inst__abc_21203_new_n1667_));
OR2X2 OR2X2_1884 ( .A(w_mem_inst_w_mem_2__0_), .B(w_mem_inst_w_mem_0__0_), .Y(w_mem_inst__abc_21203_new_n1670_));
OR2X2 OR2X2_1885 ( .A(w_mem_inst__abc_21203_new_n1669_), .B(w_mem_inst__abc_21203_new_n1673_), .Y(w_mem_inst__abc_21203_new_n1674_));
OR2X2 OR2X2_1886 ( .A(w_mem_inst__abc_21203_new_n1675_), .B(w_mem_inst__abc_21203_new_n1668_), .Y(w_mem_inst__abc_21203_new_n1676_));
OR2X2 OR2X2_1887 ( .A(w_mem_inst__abc_21203_new_n1677_), .B(w_mem_inst__abc_21203_new_n1587_), .Y(w_mem_inst__abc_21203_new_n1678_));
OR2X2 OR2X2_1888 ( .A(w_mem_inst__abc_21203_new_n1679_), .B(w_mem_inst__abc_21203_new_n1586_), .Y(w_mem_inst__abc_21203_new_n1680_));
OR2X2 OR2X2_1889 ( .A(w_mem_inst__abc_21203_new_n1681_), .B(w_mem_inst__abc_21203_new_n1682_), .Y(w_mem_inst__abc_21203_new_n1683_));
OR2X2 OR2X2_189 ( .A(_abc_15497_new_n1295_), .B(_abc_15497_new_n1281_), .Y(_0H4_reg_31_0__18_));
OR2X2 OR2X2_1890 ( .A(w_mem_inst__abc_21203_new_n1683_), .B(w_mem_inst__abc_21203_new_n1680_), .Y(w_mem_inst__abc_21203_new_n1684_));
OR2X2 OR2X2_1891 ( .A(w_mem_inst__abc_21203_new_n1685_), .B(w_mem_inst__abc_21203_new_n1686_), .Y(w_mem_inst__abc_21203_new_n1687_));
OR2X2 OR2X2_1892 ( .A(w_mem_inst__abc_21203_new_n1684_), .B(w_mem_inst__abc_21203_new_n1687_), .Y(w_mem_inst__abc_21203_new_n1688_));
OR2X2 OR2X2_1893 ( .A(w_mem_inst__abc_21203_new_n1690_), .B(w_mem_inst__abc_21203_new_n1691_), .Y(w_mem_inst__abc_21203_new_n1692_));
OR2X2 OR2X2_1894 ( .A(w_mem_inst__abc_21203_new_n1692_), .B(w_mem_inst__abc_21203_new_n1689_), .Y(w_mem_inst__abc_21203_new_n1693_));
OR2X2 OR2X2_1895 ( .A(w_mem_inst__abc_21203_new_n1694_), .B(w_mem_inst__abc_21203_new_n1695_), .Y(w_mem_inst__abc_21203_new_n1696_));
OR2X2 OR2X2_1896 ( .A(w_mem_inst__abc_21203_new_n1697_), .B(w_mem_inst__abc_21203_new_n1698_), .Y(w_mem_inst__abc_21203_new_n1699_));
OR2X2 OR2X2_1897 ( .A(w_mem_inst__abc_21203_new_n1696_), .B(w_mem_inst__abc_21203_new_n1699_), .Y(w_mem_inst__abc_21203_new_n1700_));
OR2X2 OR2X2_1898 ( .A(w_mem_inst__abc_21203_new_n1701_), .B(w_mem_inst__abc_21203_new_n1702_), .Y(w_mem_inst__abc_21203_new_n1703_));
OR2X2 OR2X2_1899 ( .A(w_mem_inst__abc_21203_new_n1704_), .B(w_mem_inst__abc_21203_new_n1705_), .Y(w_mem_inst__abc_21203_new_n1706_));
OR2X2 OR2X2_19 ( .A(_abc_15497_new_n777_), .B(_abc_15497_new_n779_), .Y(_abc_15497_new_n780_));
OR2X2 OR2X2_190 ( .A(e_reg_19_), .B(\digest[19] ), .Y(_abc_15497_new_n1300_));
OR2X2 OR2X2_1900 ( .A(w_mem_inst__abc_21203_new_n1703_), .B(w_mem_inst__abc_21203_new_n1706_), .Y(w_mem_inst__abc_21203_new_n1707_));
OR2X2 OR2X2_1901 ( .A(w_mem_inst__abc_21203_new_n1700_), .B(w_mem_inst__abc_21203_new_n1707_), .Y(w_mem_inst__abc_21203_new_n1708_));
OR2X2 OR2X2_1902 ( .A(w_mem_inst__abc_21203_new_n1708_), .B(w_mem_inst__abc_21203_new_n1693_), .Y(w_mem_inst__abc_21203_new_n1709_));
OR2X2 OR2X2_1903 ( .A(w_mem_inst__abc_21203_new_n1709_), .B(w_mem_inst__abc_21203_new_n1688_), .Y(w_mem_inst__abc_21203_new_n1710_));
OR2X2 OR2X2_1904 ( .A(w_mem_inst__abc_21203_new_n1712_), .B(w_mem_inst_w_mem_8__1_), .Y(w_mem_inst__abc_21203_new_n1713_));
OR2X2 OR2X2_1905 ( .A(w_mem_inst__abc_21203_new_n1714_), .B(w_mem_inst_w_mem_13__1_), .Y(w_mem_inst__abc_21203_new_n1715_));
OR2X2 OR2X2_1906 ( .A(w_mem_inst_w_mem_2__1_), .B(w_mem_inst_w_mem_0__1_), .Y(w_mem_inst__abc_21203_new_n1718_));
OR2X2 OR2X2_1907 ( .A(w_mem_inst__abc_21203_new_n1717_), .B(w_mem_inst__abc_21203_new_n1721_), .Y(w_mem_inst__abc_21203_new_n1722_));
OR2X2 OR2X2_1908 ( .A(w_mem_inst__abc_21203_new_n1723_), .B(w_mem_inst__abc_21203_new_n1716_), .Y(w_mem_inst__abc_21203_new_n1724_));
OR2X2 OR2X2_1909 ( .A(w_mem_inst__abc_21203_new_n1725_), .B(w_mem_inst__abc_21203_new_n1587_), .Y(w_mem_inst__abc_21203_new_n1726_));
OR2X2 OR2X2_191 ( .A(_abc_15497_new_n1299_), .B(_abc_15497_new_n1303_), .Y(_abc_15497_new_n1304_));
OR2X2 OR2X2_1910 ( .A(w_mem_inst__abc_21203_new_n1727_), .B(w_mem_inst__abc_21203_new_n1586_), .Y(w_mem_inst__abc_21203_new_n1728_));
OR2X2 OR2X2_1911 ( .A(w_mem_inst__abc_21203_new_n1729_), .B(w_mem_inst__abc_21203_new_n1730_), .Y(w_mem_inst__abc_21203_new_n1731_));
OR2X2 OR2X2_1912 ( .A(w_mem_inst__abc_21203_new_n1731_), .B(w_mem_inst__abc_21203_new_n1728_), .Y(w_mem_inst__abc_21203_new_n1732_));
OR2X2 OR2X2_1913 ( .A(w_mem_inst__abc_21203_new_n1733_), .B(w_mem_inst__abc_21203_new_n1734_), .Y(w_mem_inst__abc_21203_new_n1735_));
OR2X2 OR2X2_1914 ( .A(w_mem_inst__abc_21203_new_n1732_), .B(w_mem_inst__abc_21203_new_n1735_), .Y(w_mem_inst__abc_21203_new_n1736_));
OR2X2 OR2X2_1915 ( .A(w_mem_inst__abc_21203_new_n1738_), .B(w_mem_inst__abc_21203_new_n1739_), .Y(w_mem_inst__abc_21203_new_n1740_));
OR2X2 OR2X2_1916 ( .A(w_mem_inst__abc_21203_new_n1740_), .B(w_mem_inst__abc_21203_new_n1737_), .Y(w_mem_inst__abc_21203_new_n1741_));
OR2X2 OR2X2_1917 ( .A(w_mem_inst__abc_21203_new_n1742_), .B(w_mem_inst__abc_21203_new_n1743_), .Y(w_mem_inst__abc_21203_new_n1744_));
OR2X2 OR2X2_1918 ( .A(w_mem_inst__abc_21203_new_n1745_), .B(w_mem_inst__abc_21203_new_n1746_), .Y(w_mem_inst__abc_21203_new_n1747_));
OR2X2 OR2X2_1919 ( .A(w_mem_inst__abc_21203_new_n1744_), .B(w_mem_inst__abc_21203_new_n1747_), .Y(w_mem_inst__abc_21203_new_n1748_));
OR2X2 OR2X2_192 ( .A(_abc_15497_new_n1298_), .B(_abc_15497_new_n1305_), .Y(_abc_15497_new_n1306_));
OR2X2 OR2X2_1920 ( .A(w_mem_inst__abc_21203_new_n1749_), .B(w_mem_inst__abc_21203_new_n1750_), .Y(w_mem_inst__abc_21203_new_n1751_));
OR2X2 OR2X2_1921 ( .A(w_mem_inst__abc_21203_new_n1752_), .B(w_mem_inst__abc_21203_new_n1753_), .Y(w_mem_inst__abc_21203_new_n1754_));
OR2X2 OR2X2_1922 ( .A(w_mem_inst__abc_21203_new_n1751_), .B(w_mem_inst__abc_21203_new_n1754_), .Y(w_mem_inst__abc_21203_new_n1755_));
OR2X2 OR2X2_1923 ( .A(w_mem_inst__abc_21203_new_n1748_), .B(w_mem_inst__abc_21203_new_n1755_), .Y(w_mem_inst__abc_21203_new_n1756_));
OR2X2 OR2X2_1924 ( .A(w_mem_inst__abc_21203_new_n1756_), .B(w_mem_inst__abc_21203_new_n1741_), .Y(w_mem_inst__abc_21203_new_n1757_));
OR2X2 OR2X2_1925 ( .A(w_mem_inst__abc_21203_new_n1757_), .B(w_mem_inst__abc_21203_new_n1736_), .Y(w_mem_inst__abc_21203_new_n1758_));
OR2X2 OR2X2_1926 ( .A(w_mem_inst__abc_21203_new_n1760_), .B(w_mem_inst_w_mem_8__2_), .Y(w_mem_inst__abc_21203_new_n1761_));
OR2X2 OR2X2_1927 ( .A(w_mem_inst__abc_21203_new_n1762_), .B(w_mem_inst_w_mem_13__2_), .Y(w_mem_inst__abc_21203_new_n1763_));
OR2X2 OR2X2_1928 ( .A(w_mem_inst_w_mem_2__2_), .B(w_mem_inst_w_mem_0__2_), .Y(w_mem_inst__abc_21203_new_n1766_));
OR2X2 OR2X2_1929 ( .A(w_mem_inst__abc_21203_new_n1765_), .B(w_mem_inst__abc_21203_new_n1769_), .Y(w_mem_inst__abc_21203_new_n1770_));
OR2X2 OR2X2_193 ( .A(_abc_15497_new_n1308_), .B(_abc_15497_new_n1297_), .Y(_0H4_reg_31_0__19_));
OR2X2 OR2X2_1930 ( .A(w_mem_inst__abc_21203_new_n1771_), .B(w_mem_inst__abc_21203_new_n1764_), .Y(w_mem_inst__abc_21203_new_n1772_));
OR2X2 OR2X2_1931 ( .A(w_mem_inst__abc_21203_new_n1773_), .B(w_mem_inst__abc_21203_new_n1587_), .Y(w_mem_inst__abc_21203_new_n1774_));
OR2X2 OR2X2_1932 ( .A(w_mem_inst__abc_21203_new_n1775_), .B(w_mem_inst__abc_21203_new_n1586_), .Y(w_mem_inst__abc_21203_new_n1776_));
OR2X2 OR2X2_1933 ( .A(w_mem_inst__abc_21203_new_n1777_), .B(w_mem_inst__abc_21203_new_n1778_), .Y(w_mem_inst__abc_21203_new_n1779_));
OR2X2 OR2X2_1934 ( .A(w_mem_inst__abc_21203_new_n1779_), .B(w_mem_inst__abc_21203_new_n1776_), .Y(w_mem_inst__abc_21203_new_n1780_));
OR2X2 OR2X2_1935 ( .A(w_mem_inst__abc_21203_new_n1781_), .B(w_mem_inst__abc_21203_new_n1782_), .Y(w_mem_inst__abc_21203_new_n1783_));
OR2X2 OR2X2_1936 ( .A(w_mem_inst__abc_21203_new_n1780_), .B(w_mem_inst__abc_21203_new_n1783_), .Y(w_mem_inst__abc_21203_new_n1784_));
OR2X2 OR2X2_1937 ( .A(w_mem_inst__abc_21203_new_n1786_), .B(w_mem_inst__abc_21203_new_n1787_), .Y(w_mem_inst__abc_21203_new_n1788_));
OR2X2 OR2X2_1938 ( .A(w_mem_inst__abc_21203_new_n1788_), .B(w_mem_inst__abc_21203_new_n1785_), .Y(w_mem_inst__abc_21203_new_n1789_));
OR2X2 OR2X2_1939 ( .A(w_mem_inst__abc_21203_new_n1790_), .B(w_mem_inst__abc_21203_new_n1791_), .Y(w_mem_inst__abc_21203_new_n1792_));
OR2X2 OR2X2_194 ( .A(_abc_15497_new_n1310_), .B(_abc_15497_new_n1301_), .Y(_abc_15497_new_n1311_));
OR2X2 OR2X2_1940 ( .A(w_mem_inst__abc_21203_new_n1793_), .B(w_mem_inst__abc_21203_new_n1794_), .Y(w_mem_inst__abc_21203_new_n1795_));
OR2X2 OR2X2_1941 ( .A(w_mem_inst__abc_21203_new_n1792_), .B(w_mem_inst__abc_21203_new_n1795_), .Y(w_mem_inst__abc_21203_new_n1796_));
OR2X2 OR2X2_1942 ( .A(w_mem_inst__abc_21203_new_n1797_), .B(w_mem_inst__abc_21203_new_n1798_), .Y(w_mem_inst__abc_21203_new_n1799_));
OR2X2 OR2X2_1943 ( .A(w_mem_inst__abc_21203_new_n1800_), .B(w_mem_inst__abc_21203_new_n1801_), .Y(w_mem_inst__abc_21203_new_n1802_));
OR2X2 OR2X2_1944 ( .A(w_mem_inst__abc_21203_new_n1799_), .B(w_mem_inst__abc_21203_new_n1802_), .Y(w_mem_inst__abc_21203_new_n1803_));
OR2X2 OR2X2_1945 ( .A(w_mem_inst__abc_21203_new_n1796_), .B(w_mem_inst__abc_21203_new_n1803_), .Y(w_mem_inst__abc_21203_new_n1804_));
OR2X2 OR2X2_1946 ( .A(w_mem_inst__abc_21203_new_n1804_), .B(w_mem_inst__abc_21203_new_n1789_), .Y(w_mem_inst__abc_21203_new_n1805_));
OR2X2 OR2X2_1947 ( .A(w_mem_inst__abc_21203_new_n1805_), .B(w_mem_inst__abc_21203_new_n1784_), .Y(w_mem_inst__abc_21203_new_n1806_));
OR2X2 OR2X2_1948 ( .A(w_mem_inst__abc_21203_new_n1808_), .B(w_mem_inst_w_mem_8__3_), .Y(w_mem_inst__abc_21203_new_n1809_));
OR2X2 OR2X2_1949 ( .A(w_mem_inst__abc_21203_new_n1810_), .B(w_mem_inst_w_mem_13__3_), .Y(w_mem_inst__abc_21203_new_n1811_));
OR2X2 OR2X2_195 ( .A(_abc_15497_new_n1287_), .B(_abc_15497_new_n1286_), .Y(_abc_15497_new_n1313_));
OR2X2 OR2X2_1950 ( .A(w_mem_inst_w_mem_2__3_), .B(w_mem_inst_w_mem_0__3_), .Y(w_mem_inst__abc_21203_new_n1814_));
OR2X2 OR2X2_1951 ( .A(w_mem_inst__abc_21203_new_n1813_), .B(w_mem_inst__abc_21203_new_n1817_), .Y(w_mem_inst__abc_21203_new_n1818_));
OR2X2 OR2X2_1952 ( .A(w_mem_inst__abc_21203_new_n1819_), .B(w_mem_inst__abc_21203_new_n1812_), .Y(w_mem_inst__abc_21203_new_n1820_));
OR2X2 OR2X2_1953 ( .A(w_mem_inst__abc_21203_new_n1821_), .B(w_mem_inst__abc_21203_new_n1587_), .Y(w_mem_inst__abc_21203_new_n1822_));
OR2X2 OR2X2_1954 ( .A(w_mem_inst__abc_21203_new_n1823_), .B(w_mem_inst__abc_21203_new_n1586_), .Y(w_mem_inst__abc_21203_new_n1824_));
OR2X2 OR2X2_1955 ( .A(w_mem_inst__abc_21203_new_n1825_), .B(w_mem_inst__abc_21203_new_n1826_), .Y(w_mem_inst__abc_21203_new_n1827_));
OR2X2 OR2X2_1956 ( .A(w_mem_inst__abc_21203_new_n1827_), .B(w_mem_inst__abc_21203_new_n1824_), .Y(w_mem_inst__abc_21203_new_n1828_));
OR2X2 OR2X2_1957 ( .A(w_mem_inst__abc_21203_new_n1829_), .B(w_mem_inst__abc_21203_new_n1830_), .Y(w_mem_inst__abc_21203_new_n1831_));
OR2X2 OR2X2_1958 ( .A(w_mem_inst__abc_21203_new_n1828_), .B(w_mem_inst__abc_21203_new_n1831_), .Y(w_mem_inst__abc_21203_new_n1832_));
OR2X2 OR2X2_1959 ( .A(w_mem_inst__abc_21203_new_n1834_), .B(w_mem_inst__abc_21203_new_n1835_), .Y(w_mem_inst__abc_21203_new_n1836_));
OR2X2 OR2X2_196 ( .A(_abc_15497_new_n1315_), .B(_abc_15497_new_n1313_), .Y(_abc_15497_new_n1316_));
OR2X2 OR2X2_1960 ( .A(w_mem_inst__abc_21203_new_n1836_), .B(w_mem_inst__abc_21203_new_n1833_), .Y(w_mem_inst__abc_21203_new_n1837_));
OR2X2 OR2X2_1961 ( .A(w_mem_inst__abc_21203_new_n1838_), .B(w_mem_inst__abc_21203_new_n1839_), .Y(w_mem_inst__abc_21203_new_n1840_));
OR2X2 OR2X2_1962 ( .A(w_mem_inst__abc_21203_new_n1841_), .B(w_mem_inst__abc_21203_new_n1842_), .Y(w_mem_inst__abc_21203_new_n1843_));
OR2X2 OR2X2_1963 ( .A(w_mem_inst__abc_21203_new_n1840_), .B(w_mem_inst__abc_21203_new_n1843_), .Y(w_mem_inst__abc_21203_new_n1844_));
OR2X2 OR2X2_1964 ( .A(w_mem_inst__abc_21203_new_n1845_), .B(w_mem_inst__abc_21203_new_n1846_), .Y(w_mem_inst__abc_21203_new_n1847_));
OR2X2 OR2X2_1965 ( .A(w_mem_inst__abc_21203_new_n1848_), .B(w_mem_inst__abc_21203_new_n1849_), .Y(w_mem_inst__abc_21203_new_n1850_));
OR2X2 OR2X2_1966 ( .A(w_mem_inst__abc_21203_new_n1847_), .B(w_mem_inst__abc_21203_new_n1850_), .Y(w_mem_inst__abc_21203_new_n1851_));
OR2X2 OR2X2_1967 ( .A(w_mem_inst__abc_21203_new_n1844_), .B(w_mem_inst__abc_21203_new_n1851_), .Y(w_mem_inst__abc_21203_new_n1852_));
OR2X2 OR2X2_1968 ( .A(w_mem_inst__abc_21203_new_n1852_), .B(w_mem_inst__abc_21203_new_n1837_), .Y(w_mem_inst__abc_21203_new_n1853_));
OR2X2 OR2X2_1969 ( .A(w_mem_inst__abc_21203_new_n1853_), .B(w_mem_inst__abc_21203_new_n1832_), .Y(w_mem_inst__abc_21203_new_n1854_));
OR2X2 OR2X2_197 ( .A(_abc_15497_new_n1321_), .B(_abc_15497_new_n1318_), .Y(_abc_15497_new_n1322_));
OR2X2 OR2X2_1970 ( .A(w_mem_inst__abc_21203_new_n1856_), .B(w_mem_inst_w_mem_8__4_), .Y(w_mem_inst__abc_21203_new_n1857_));
OR2X2 OR2X2_1971 ( .A(w_mem_inst__abc_21203_new_n1858_), .B(w_mem_inst_w_mem_13__4_), .Y(w_mem_inst__abc_21203_new_n1859_));
OR2X2 OR2X2_1972 ( .A(w_mem_inst_w_mem_2__4_), .B(w_mem_inst_w_mem_0__4_), .Y(w_mem_inst__abc_21203_new_n1862_));
OR2X2 OR2X2_1973 ( .A(w_mem_inst__abc_21203_new_n1861_), .B(w_mem_inst__abc_21203_new_n1865_), .Y(w_mem_inst__abc_21203_new_n1866_));
OR2X2 OR2X2_1974 ( .A(w_mem_inst__abc_21203_new_n1867_), .B(w_mem_inst__abc_21203_new_n1860_), .Y(w_mem_inst__abc_21203_new_n1868_));
OR2X2 OR2X2_1975 ( .A(w_mem_inst__abc_21203_new_n1869_), .B(w_mem_inst__abc_21203_new_n1587_), .Y(w_mem_inst__abc_21203_new_n1870_));
OR2X2 OR2X2_1976 ( .A(w_mem_inst__abc_21203_new_n1871_), .B(w_mem_inst__abc_21203_new_n1586_), .Y(w_mem_inst__abc_21203_new_n1872_));
OR2X2 OR2X2_1977 ( .A(w_mem_inst__abc_21203_new_n1873_), .B(w_mem_inst__abc_21203_new_n1874_), .Y(w_mem_inst__abc_21203_new_n1875_));
OR2X2 OR2X2_1978 ( .A(w_mem_inst__abc_21203_new_n1875_), .B(w_mem_inst__abc_21203_new_n1872_), .Y(w_mem_inst__abc_21203_new_n1876_));
OR2X2 OR2X2_1979 ( .A(w_mem_inst__abc_21203_new_n1877_), .B(w_mem_inst__abc_21203_new_n1878_), .Y(w_mem_inst__abc_21203_new_n1879_));
OR2X2 OR2X2_198 ( .A(e_reg_20_), .B(\digest[20] ), .Y(_abc_15497_new_n1323_));
OR2X2 OR2X2_1980 ( .A(w_mem_inst__abc_21203_new_n1876_), .B(w_mem_inst__abc_21203_new_n1879_), .Y(w_mem_inst__abc_21203_new_n1880_));
OR2X2 OR2X2_1981 ( .A(w_mem_inst__abc_21203_new_n1882_), .B(w_mem_inst__abc_21203_new_n1883_), .Y(w_mem_inst__abc_21203_new_n1884_));
OR2X2 OR2X2_1982 ( .A(w_mem_inst__abc_21203_new_n1884_), .B(w_mem_inst__abc_21203_new_n1881_), .Y(w_mem_inst__abc_21203_new_n1885_));
OR2X2 OR2X2_1983 ( .A(w_mem_inst__abc_21203_new_n1886_), .B(w_mem_inst__abc_21203_new_n1887_), .Y(w_mem_inst__abc_21203_new_n1888_));
OR2X2 OR2X2_1984 ( .A(w_mem_inst__abc_21203_new_n1889_), .B(w_mem_inst__abc_21203_new_n1890_), .Y(w_mem_inst__abc_21203_new_n1891_));
OR2X2 OR2X2_1985 ( .A(w_mem_inst__abc_21203_new_n1888_), .B(w_mem_inst__abc_21203_new_n1891_), .Y(w_mem_inst__abc_21203_new_n1892_));
OR2X2 OR2X2_1986 ( .A(w_mem_inst__abc_21203_new_n1893_), .B(w_mem_inst__abc_21203_new_n1894_), .Y(w_mem_inst__abc_21203_new_n1895_));
OR2X2 OR2X2_1987 ( .A(w_mem_inst__abc_21203_new_n1896_), .B(w_mem_inst__abc_21203_new_n1897_), .Y(w_mem_inst__abc_21203_new_n1898_));
OR2X2 OR2X2_1988 ( .A(w_mem_inst__abc_21203_new_n1895_), .B(w_mem_inst__abc_21203_new_n1898_), .Y(w_mem_inst__abc_21203_new_n1899_));
OR2X2 OR2X2_1989 ( .A(w_mem_inst__abc_21203_new_n1892_), .B(w_mem_inst__abc_21203_new_n1899_), .Y(w_mem_inst__abc_21203_new_n1900_));
OR2X2 OR2X2_199 ( .A(_abc_15497_new_n1322_), .B(_abc_15497_new_n1326_), .Y(_abc_15497_new_n1327_));
OR2X2 OR2X2_1990 ( .A(w_mem_inst__abc_21203_new_n1900_), .B(w_mem_inst__abc_21203_new_n1885_), .Y(w_mem_inst__abc_21203_new_n1901_));
OR2X2 OR2X2_1991 ( .A(w_mem_inst__abc_21203_new_n1901_), .B(w_mem_inst__abc_21203_new_n1880_), .Y(w_mem_inst__abc_21203_new_n1902_));
OR2X2 OR2X2_1992 ( .A(w_mem_inst__abc_21203_new_n1904_), .B(w_mem_inst_w_mem_8__5_), .Y(w_mem_inst__abc_21203_new_n1905_));
OR2X2 OR2X2_1993 ( .A(w_mem_inst__abc_21203_new_n1906_), .B(w_mem_inst_w_mem_13__5_), .Y(w_mem_inst__abc_21203_new_n1907_));
OR2X2 OR2X2_1994 ( .A(w_mem_inst_w_mem_2__5_), .B(w_mem_inst_w_mem_0__5_), .Y(w_mem_inst__abc_21203_new_n1910_));
OR2X2 OR2X2_1995 ( .A(w_mem_inst__abc_21203_new_n1909_), .B(w_mem_inst__abc_21203_new_n1913_), .Y(w_mem_inst__abc_21203_new_n1914_));
OR2X2 OR2X2_1996 ( .A(w_mem_inst__abc_21203_new_n1915_), .B(w_mem_inst__abc_21203_new_n1908_), .Y(w_mem_inst__abc_21203_new_n1916_));
OR2X2 OR2X2_1997 ( .A(w_mem_inst__abc_21203_new_n1917_), .B(w_mem_inst__abc_21203_new_n1587_), .Y(w_mem_inst__abc_21203_new_n1918_));
OR2X2 OR2X2_1998 ( .A(w_mem_inst__abc_21203_new_n1919_), .B(w_mem_inst__abc_21203_new_n1586_), .Y(w_mem_inst__abc_21203_new_n1920_));
OR2X2 OR2X2_1999 ( .A(w_mem_inst__abc_21203_new_n1921_), .B(w_mem_inst__abc_21203_new_n1922_), .Y(w_mem_inst__abc_21203_new_n1923_));
OR2X2 OR2X2_2 ( .A(c_reg_22_), .B(\digest[86] ), .Y(_abc_15497_new_n709_));
OR2X2 OR2X2_20 ( .A(c_reg_12_), .B(\digest[76] ), .Y(_abc_15497_new_n781_));
OR2X2 OR2X2_200 ( .A(_abc_15497_new_n699_), .B(\digest[20] ), .Y(_abc_15497_new_n1332_));
OR2X2 OR2X2_2000 ( .A(w_mem_inst__abc_21203_new_n1923_), .B(w_mem_inst__abc_21203_new_n1920_), .Y(w_mem_inst__abc_21203_new_n1924_));
OR2X2 OR2X2_2001 ( .A(w_mem_inst__abc_21203_new_n1925_), .B(w_mem_inst__abc_21203_new_n1926_), .Y(w_mem_inst__abc_21203_new_n1927_));
OR2X2 OR2X2_2002 ( .A(w_mem_inst__abc_21203_new_n1924_), .B(w_mem_inst__abc_21203_new_n1927_), .Y(w_mem_inst__abc_21203_new_n1928_));
OR2X2 OR2X2_2003 ( .A(w_mem_inst__abc_21203_new_n1930_), .B(w_mem_inst__abc_21203_new_n1931_), .Y(w_mem_inst__abc_21203_new_n1932_));
OR2X2 OR2X2_2004 ( .A(w_mem_inst__abc_21203_new_n1932_), .B(w_mem_inst__abc_21203_new_n1929_), .Y(w_mem_inst__abc_21203_new_n1933_));
OR2X2 OR2X2_2005 ( .A(w_mem_inst__abc_21203_new_n1934_), .B(w_mem_inst__abc_21203_new_n1935_), .Y(w_mem_inst__abc_21203_new_n1936_));
OR2X2 OR2X2_2006 ( .A(w_mem_inst__abc_21203_new_n1937_), .B(w_mem_inst__abc_21203_new_n1938_), .Y(w_mem_inst__abc_21203_new_n1939_));
OR2X2 OR2X2_2007 ( .A(w_mem_inst__abc_21203_new_n1936_), .B(w_mem_inst__abc_21203_new_n1939_), .Y(w_mem_inst__abc_21203_new_n1940_));
OR2X2 OR2X2_2008 ( .A(w_mem_inst__abc_21203_new_n1941_), .B(w_mem_inst__abc_21203_new_n1942_), .Y(w_mem_inst__abc_21203_new_n1943_));
OR2X2 OR2X2_2009 ( .A(w_mem_inst__abc_21203_new_n1944_), .B(w_mem_inst__abc_21203_new_n1945_), .Y(w_mem_inst__abc_21203_new_n1946_));
OR2X2 OR2X2_201 ( .A(_abc_15497_new_n1331_), .B(_abc_15497_new_n1333_), .Y(_0H4_reg_31_0__20_));
OR2X2 OR2X2_2010 ( .A(w_mem_inst__abc_21203_new_n1943_), .B(w_mem_inst__abc_21203_new_n1946_), .Y(w_mem_inst__abc_21203_new_n1947_));
OR2X2 OR2X2_2011 ( .A(w_mem_inst__abc_21203_new_n1940_), .B(w_mem_inst__abc_21203_new_n1947_), .Y(w_mem_inst__abc_21203_new_n1948_));
OR2X2 OR2X2_2012 ( .A(w_mem_inst__abc_21203_new_n1948_), .B(w_mem_inst__abc_21203_new_n1933_), .Y(w_mem_inst__abc_21203_new_n1949_));
OR2X2 OR2X2_2013 ( .A(w_mem_inst__abc_21203_new_n1949_), .B(w_mem_inst__abc_21203_new_n1928_), .Y(w_mem_inst__abc_21203_new_n1950_));
OR2X2 OR2X2_2014 ( .A(w_mem_inst__abc_21203_new_n1952_), .B(w_mem_inst_w_mem_8__6_), .Y(w_mem_inst__abc_21203_new_n1953_));
OR2X2 OR2X2_2015 ( .A(w_mem_inst__abc_21203_new_n1954_), .B(w_mem_inst_w_mem_13__6_), .Y(w_mem_inst__abc_21203_new_n1955_));
OR2X2 OR2X2_2016 ( .A(w_mem_inst_w_mem_2__6_), .B(w_mem_inst_w_mem_0__6_), .Y(w_mem_inst__abc_21203_new_n1958_));
OR2X2 OR2X2_2017 ( .A(w_mem_inst__abc_21203_new_n1957_), .B(w_mem_inst__abc_21203_new_n1961_), .Y(w_mem_inst__abc_21203_new_n1962_));
OR2X2 OR2X2_2018 ( .A(w_mem_inst__abc_21203_new_n1963_), .B(w_mem_inst__abc_21203_new_n1956_), .Y(w_mem_inst__abc_21203_new_n1964_));
OR2X2 OR2X2_2019 ( .A(w_mem_inst__abc_21203_new_n1965_), .B(w_mem_inst__abc_21203_new_n1587_), .Y(w_mem_inst__abc_21203_new_n1966_));
OR2X2 OR2X2_202 ( .A(e_reg_21_), .B(\digest[21] ), .Y(_abc_15497_new_n1336_));
OR2X2 OR2X2_2020 ( .A(w_mem_inst__abc_21203_new_n1967_), .B(w_mem_inst__abc_21203_new_n1586_), .Y(w_mem_inst__abc_21203_new_n1968_));
OR2X2 OR2X2_2021 ( .A(w_mem_inst__abc_21203_new_n1969_), .B(w_mem_inst__abc_21203_new_n1970_), .Y(w_mem_inst__abc_21203_new_n1971_));
OR2X2 OR2X2_2022 ( .A(w_mem_inst__abc_21203_new_n1971_), .B(w_mem_inst__abc_21203_new_n1968_), .Y(w_mem_inst__abc_21203_new_n1972_));
OR2X2 OR2X2_2023 ( .A(w_mem_inst__abc_21203_new_n1973_), .B(w_mem_inst__abc_21203_new_n1974_), .Y(w_mem_inst__abc_21203_new_n1975_));
OR2X2 OR2X2_2024 ( .A(w_mem_inst__abc_21203_new_n1972_), .B(w_mem_inst__abc_21203_new_n1975_), .Y(w_mem_inst__abc_21203_new_n1976_));
OR2X2 OR2X2_2025 ( .A(w_mem_inst__abc_21203_new_n1978_), .B(w_mem_inst__abc_21203_new_n1979_), .Y(w_mem_inst__abc_21203_new_n1980_));
OR2X2 OR2X2_2026 ( .A(w_mem_inst__abc_21203_new_n1980_), .B(w_mem_inst__abc_21203_new_n1977_), .Y(w_mem_inst__abc_21203_new_n1981_));
OR2X2 OR2X2_2027 ( .A(w_mem_inst__abc_21203_new_n1982_), .B(w_mem_inst__abc_21203_new_n1983_), .Y(w_mem_inst__abc_21203_new_n1984_));
OR2X2 OR2X2_2028 ( .A(w_mem_inst__abc_21203_new_n1985_), .B(w_mem_inst__abc_21203_new_n1986_), .Y(w_mem_inst__abc_21203_new_n1987_));
OR2X2 OR2X2_2029 ( .A(w_mem_inst__abc_21203_new_n1984_), .B(w_mem_inst__abc_21203_new_n1987_), .Y(w_mem_inst__abc_21203_new_n1988_));
OR2X2 OR2X2_203 ( .A(_abc_15497_new_n1339_), .B(_abc_15497_new_n1324_), .Y(_abc_15497_new_n1340_));
OR2X2 OR2X2_2030 ( .A(w_mem_inst__abc_21203_new_n1989_), .B(w_mem_inst__abc_21203_new_n1990_), .Y(w_mem_inst__abc_21203_new_n1991_));
OR2X2 OR2X2_2031 ( .A(w_mem_inst__abc_21203_new_n1992_), .B(w_mem_inst__abc_21203_new_n1993_), .Y(w_mem_inst__abc_21203_new_n1994_));
OR2X2 OR2X2_2032 ( .A(w_mem_inst__abc_21203_new_n1991_), .B(w_mem_inst__abc_21203_new_n1994_), .Y(w_mem_inst__abc_21203_new_n1995_));
OR2X2 OR2X2_2033 ( .A(w_mem_inst__abc_21203_new_n1988_), .B(w_mem_inst__abc_21203_new_n1995_), .Y(w_mem_inst__abc_21203_new_n1996_));
OR2X2 OR2X2_2034 ( .A(w_mem_inst__abc_21203_new_n1996_), .B(w_mem_inst__abc_21203_new_n1981_), .Y(w_mem_inst__abc_21203_new_n1997_));
OR2X2 OR2X2_2035 ( .A(w_mem_inst__abc_21203_new_n1997_), .B(w_mem_inst__abc_21203_new_n1976_), .Y(w_mem_inst__abc_21203_new_n1998_));
OR2X2 OR2X2_2036 ( .A(w_mem_inst__abc_21203_new_n2000_), .B(w_mem_inst_w_mem_8__7_), .Y(w_mem_inst__abc_21203_new_n2001_));
OR2X2 OR2X2_2037 ( .A(w_mem_inst__abc_21203_new_n2002_), .B(w_mem_inst_w_mem_13__7_), .Y(w_mem_inst__abc_21203_new_n2003_));
OR2X2 OR2X2_2038 ( .A(w_mem_inst_w_mem_2__7_), .B(w_mem_inst_w_mem_0__7_), .Y(w_mem_inst__abc_21203_new_n2006_));
OR2X2 OR2X2_2039 ( .A(w_mem_inst__abc_21203_new_n2005_), .B(w_mem_inst__abc_21203_new_n2009_), .Y(w_mem_inst__abc_21203_new_n2010_));
OR2X2 OR2X2_204 ( .A(_abc_15497_new_n1328_), .B(_abc_15497_new_n1340_), .Y(_abc_15497_new_n1341_));
OR2X2 OR2X2_2040 ( .A(w_mem_inst__abc_21203_new_n2011_), .B(w_mem_inst__abc_21203_new_n2004_), .Y(w_mem_inst__abc_21203_new_n2012_));
OR2X2 OR2X2_2041 ( .A(w_mem_inst__abc_21203_new_n2013_), .B(w_mem_inst__abc_21203_new_n1587_), .Y(w_mem_inst__abc_21203_new_n2014_));
OR2X2 OR2X2_2042 ( .A(w_mem_inst__abc_21203_new_n2015_), .B(w_mem_inst__abc_21203_new_n1586_), .Y(w_mem_inst__abc_21203_new_n2016_));
OR2X2 OR2X2_2043 ( .A(w_mem_inst__abc_21203_new_n2017_), .B(w_mem_inst__abc_21203_new_n2018_), .Y(w_mem_inst__abc_21203_new_n2019_));
OR2X2 OR2X2_2044 ( .A(w_mem_inst__abc_21203_new_n2019_), .B(w_mem_inst__abc_21203_new_n2016_), .Y(w_mem_inst__abc_21203_new_n2020_));
OR2X2 OR2X2_2045 ( .A(w_mem_inst__abc_21203_new_n2021_), .B(w_mem_inst__abc_21203_new_n2022_), .Y(w_mem_inst__abc_21203_new_n2023_));
OR2X2 OR2X2_2046 ( .A(w_mem_inst__abc_21203_new_n2020_), .B(w_mem_inst__abc_21203_new_n2023_), .Y(w_mem_inst__abc_21203_new_n2024_));
OR2X2 OR2X2_2047 ( .A(w_mem_inst__abc_21203_new_n2026_), .B(w_mem_inst__abc_21203_new_n2027_), .Y(w_mem_inst__abc_21203_new_n2028_));
OR2X2 OR2X2_2048 ( .A(w_mem_inst__abc_21203_new_n2028_), .B(w_mem_inst__abc_21203_new_n2025_), .Y(w_mem_inst__abc_21203_new_n2029_));
OR2X2 OR2X2_2049 ( .A(w_mem_inst__abc_21203_new_n2030_), .B(w_mem_inst__abc_21203_new_n2031_), .Y(w_mem_inst__abc_21203_new_n2032_));
OR2X2 OR2X2_205 ( .A(_abc_15497_new_n1349_), .B(_abc_15497_new_n1335_), .Y(_0H4_reg_31_0__21_));
OR2X2 OR2X2_2050 ( .A(w_mem_inst__abc_21203_new_n2033_), .B(w_mem_inst__abc_21203_new_n2034_), .Y(w_mem_inst__abc_21203_new_n2035_));
OR2X2 OR2X2_2051 ( .A(w_mem_inst__abc_21203_new_n2032_), .B(w_mem_inst__abc_21203_new_n2035_), .Y(w_mem_inst__abc_21203_new_n2036_));
OR2X2 OR2X2_2052 ( .A(w_mem_inst__abc_21203_new_n2037_), .B(w_mem_inst__abc_21203_new_n2038_), .Y(w_mem_inst__abc_21203_new_n2039_));
OR2X2 OR2X2_2053 ( .A(w_mem_inst__abc_21203_new_n2040_), .B(w_mem_inst__abc_21203_new_n2041_), .Y(w_mem_inst__abc_21203_new_n2042_));
OR2X2 OR2X2_2054 ( .A(w_mem_inst__abc_21203_new_n2039_), .B(w_mem_inst__abc_21203_new_n2042_), .Y(w_mem_inst__abc_21203_new_n2043_));
OR2X2 OR2X2_2055 ( .A(w_mem_inst__abc_21203_new_n2036_), .B(w_mem_inst__abc_21203_new_n2043_), .Y(w_mem_inst__abc_21203_new_n2044_));
OR2X2 OR2X2_2056 ( .A(w_mem_inst__abc_21203_new_n2044_), .B(w_mem_inst__abc_21203_new_n2029_), .Y(w_mem_inst__abc_21203_new_n2045_));
OR2X2 OR2X2_2057 ( .A(w_mem_inst__abc_21203_new_n2045_), .B(w_mem_inst__abc_21203_new_n2024_), .Y(w_mem_inst__abc_21203_new_n2046_));
OR2X2 OR2X2_2058 ( .A(w_mem_inst__abc_21203_new_n2048_), .B(w_mem_inst_w_mem_8__8_), .Y(w_mem_inst__abc_21203_new_n2049_));
OR2X2 OR2X2_2059 ( .A(w_mem_inst__abc_21203_new_n2050_), .B(w_mem_inst_w_mem_13__8_), .Y(w_mem_inst__abc_21203_new_n2051_));
OR2X2 OR2X2_206 ( .A(e_reg_22_), .B(\digest[22] ), .Y(_abc_15497_new_n1354_));
OR2X2 OR2X2_2060 ( .A(w_mem_inst_w_mem_2__8_), .B(w_mem_inst_w_mem_0__8_), .Y(w_mem_inst__abc_21203_new_n2054_));
OR2X2 OR2X2_2061 ( .A(w_mem_inst__abc_21203_new_n2053_), .B(w_mem_inst__abc_21203_new_n2057_), .Y(w_mem_inst__abc_21203_new_n2058_));
OR2X2 OR2X2_2062 ( .A(w_mem_inst__abc_21203_new_n2059_), .B(w_mem_inst__abc_21203_new_n2052_), .Y(w_mem_inst__abc_21203_new_n2060_));
OR2X2 OR2X2_2063 ( .A(w_mem_inst__abc_21203_new_n2061_), .B(w_mem_inst__abc_21203_new_n1587_), .Y(w_mem_inst__abc_21203_new_n2062_));
OR2X2 OR2X2_2064 ( .A(w_mem_inst__abc_21203_new_n2063_), .B(w_mem_inst__abc_21203_new_n1586_), .Y(w_mem_inst__abc_21203_new_n2064_));
OR2X2 OR2X2_2065 ( .A(w_mem_inst__abc_21203_new_n2065_), .B(w_mem_inst__abc_21203_new_n2066_), .Y(w_mem_inst__abc_21203_new_n2067_));
OR2X2 OR2X2_2066 ( .A(w_mem_inst__abc_21203_new_n2067_), .B(w_mem_inst__abc_21203_new_n2064_), .Y(w_mem_inst__abc_21203_new_n2068_));
OR2X2 OR2X2_2067 ( .A(w_mem_inst__abc_21203_new_n2069_), .B(w_mem_inst__abc_21203_new_n2070_), .Y(w_mem_inst__abc_21203_new_n2071_));
OR2X2 OR2X2_2068 ( .A(w_mem_inst__abc_21203_new_n2068_), .B(w_mem_inst__abc_21203_new_n2071_), .Y(w_mem_inst__abc_21203_new_n2072_));
OR2X2 OR2X2_2069 ( .A(w_mem_inst__abc_21203_new_n2074_), .B(w_mem_inst__abc_21203_new_n2075_), .Y(w_mem_inst__abc_21203_new_n2076_));
OR2X2 OR2X2_207 ( .A(_abc_15497_new_n1353_), .B(_abc_15497_new_n1357_), .Y(_abc_15497_new_n1358_));
OR2X2 OR2X2_2070 ( .A(w_mem_inst__abc_21203_new_n2076_), .B(w_mem_inst__abc_21203_new_n2073_), .Y(w_mem_inst__abc_21203_new_n2077_));
OR2X2 OR2X2_2071 ( .A(w_mem_inst__abc_21203_new_n2078_), .B(w_mem_inst__abc_21203_new_n2079_), .Y(w_mem_inst__abc_21203_new_n2080_));
OR2X2 OR2X2_2072 ( .A(w_mem_inst__abc_21203_new_n2081_), .B(w_mem_inst__abc_21203_new_n2082_), .Y(w_mem_inst__abc_21203_new_n2083_));
OR2X2 OR2X2_2073 ( .A(w_mem_inst__abc_21203_new_n2080_), .B(w_mem_inst__abc_21203_new_n2083_), .Y(w_mem_inst__abc_21203_new_n2084_));
OR2X2 OR2X2_2074 ( .A(w_mem_inst__abc_21203_new_n2085_), .B(w_mem_inst__abc_21203_new_n2086_), .Y(w_mem_inst__abc_21203_new_n2087_));
OR2X2 OR2X2_2075 ( .A(w_mem_inst__abc_21203_new_n2088_), .B(w_mem_inst__abc_21203_new_n2089_), .Y(w_mem_inst__abc_21203_new_n2090_));
OR2X2 OR2X2_2076 ( .A(w_mem_inst__abc_21203_new_n2087_), .B(w_mem_inst__abc_21203_new_n2090_), .Y(w_mem_inst__abc_21203_new_n2091_));
OR2X2 OR2X2_2077 ( .A(w_mem_inst__abc_21203_new_n2084_), .B(w_mem_inst__abc_21203_new_n2091_), .Y(w_mem_inst__abc_21203_new_n2092_));
OR2X2 OR2X2_2078 ( .A(w_mem_inst__abc_21203_new_n2092_), .B(w_mem_inst__abc_21203_new_n2077_), .Y(w_mem_inst__abc_21203_new_n2093_));
OR2X2 OR2X2_2079 ( .A(w_mem_inst__abc_21203_new_n2093_), .B(w_mem_inst__abc_21203_new_n2072_), .Y(w_mem_inst__abc_21203_new_n2094_));
OR2X2 OR2X2_208 ( .A(_abc_15497_new_n699_), .B(\digest[22] ), .Y(_abc_15497_new_n1363_));
OR2X2 OR2X2_2080 ( .A(w_mem_inst__abc_21203_new_n2096_), .B(w_mem_inst_w_mem_8__9_), .Y(w_mem_inst__abc_21203_new_n2097_));
OR2X2 OR2X2_2081 ( .A(w_mem_inst__abc_21203_new_n2098_), .B(w_mem_inst_w_mem_13__9_), .Y(w_mem_inst__abc_21203_new_n2099_));
OR2X2 OR2X2_2082 ( .A(w_mem_inst_w_mem_2__9_), .B(w_mem_inst_w_mem_0__9_), .Y(w_mem_inst__abc_21203_new_n2102_));
OR2X2 OR2X2_2083 ( .A(w_mem_inst__abc_21203_new_n2101_), .B(w_mem_inst__abc_21203_new_n2105_), .Y(w_mem_inst__abc_21203_new_n2106_));
OR2X2 OR2X2_2084 ( .A(w_mem_inst__abc_21203_new_n2107_), .B(w_mem_inst__abc_21203_new_n2100_), .Y(w_mem_inst__abc_21203_new_n2108_));
OR2X2 OR2X2_2085 ( .A(w_mem_inst__abc_21203_new_n2109_), .B(w_mem_inst__abc_21203_new_n1587_), .Y(w_mem_inst__abc_21203_new_n2110_));
OR2X2 OR2X2_2086 ( .A(w_mem_inst__abc_21203_new_n2111_), .B(w_mem_inst__abc_21203_new_n1586_), .Y(w_mem_inst__abc_21203_new_n2112_));
OR2X2 OR2X2_2087 ( .A(w_mem_inst__abc_21203_new_n2113_), .B(w_mem_inst__abc_21203_new_n2114_), .Y(w_mem_inst__abc_21203_new_n2115_));
OR2X2 OR2X2_2088 ( .A(w_mem_inst__abc_21203_new_n2115_), .B(w_mem_inst__abc_21203_new_n2112_), .Y(w_mem_inst__abc_21203_new_n2116_));
OR2X2 OR2X2_2089 ( .A(w_mem_inst__abc_21203_new_n2117_), .B(w_mem_inst__abc_21203_new_n2118_), .Y(w_mem_inst__abc_21203_new_n2119_));
OR2X2 OR2X2_209 ( .A(_abc_15497_new_n1362_), .B(_abc_15497_new_n1364_), .Y(_0H4_reg_31_0__22_));
OR2X2 OR2X2_2090 ( .A(w_mem_inst__abc_21203_new_n2116_), .B(w_mem_inst__abc_21203_new_n2119_), .Y(w_mem_inst__abc_21203_new_n2120_));
OR2X2 OR2X2_2091 ( .A(w_mem_inst__abc_21203_new_n2122_), .B(w_mem_inst__abc_21203_new_n2123_), .Y(w_mem_inst__abc_21203_new_n2124_));
OR2X2 OR2X2_2092 ( .A(w_mem_inst__abc_21203_new_n2124_), .B(w_mem_inst__abc_21203_new_n2121_), .Y(w_mem_inst__abc_21203_new_n2125_));
OR2X2 OR2X2_2093 ( .A(w_mem_inst__abc_21203_new_n2126_), .B(w_mem_inst__abc_21203_new_n2127_), .Y(w_mem_inst__abc_21203_new_n2128_));
OR2X2 OR2X2_2094 ( .A(w_mem_inst__abc_21203_new_n2129_), .B(w_mem_inst__abc_21203_new_n2130_), .Y(w_mem_inst__abc_21203_new_n2131_));
OR2X2 OR2X2_2095 ( .A(w_mem_inst__abc_21203_new_n2128_), .B(w_mem_inst__abc_21203_new_n2131_), .Y(w_mem_inst__abc_21203_new_n2132_));
OR2X2 OR2X2_2096 ( .A(w_mem_inst__abc_21203_new_n2133_), .B(w_mem_inst__abc_21203_new_n2134_), .Y(w_mem_inst__abc_21203_new_n2135_));
OR2X2 OR2X2_2097 ( .A(w_mem_inst__abc_21203_new_n2136_), .B(w_mem_inst__abc_21203_new_n2137_), .Y(w_mem_inst__abc_21203_new_n2138_));
OR2X2 OR2X2_2098 ( .A(w_mem_inst__abc_21203_new_n2135_), .B(w_mem_inst__abc_21203_new_n2138_), .Y(w_mem_inst__abc_21203_new_n2139_));
OR2X2 OR2X2_2099 ( .A(w_mem_inst__abc_21203_new_n2132_), .B(w_mem_inst__abc_21203_new_n2139_), .Y(w_mem_inst__abc_21203_new_n2140_));
OR2X2 OR2X2_21 ( .A(c_reg_11_), .B(\digest[75] ), .Y(_abc_15497_new_n786_));
OR2X2 OR2X2_210 ( .A(e_reg_23_), .B(\digest[23] ), .Y(_abc_15497_new_n1367_));
OR2X2 OR2X2_2100 ( .A(w_mem_inst__abc_21203_new_n2140_), .B(w_mem_inst__abc_21203_new_n2125_), .Y(w_mem_inst__abc_21203_new_n2141_));
OR2X2 OR2X2_2101 ( .A(w_mem_inst__abc_21203_new_n2141_), .B(w_mem_inst__abc_21203_new_n2120_), .Y(w_mem_inst__abc_21203_new_n2142_));
OR2X2 OR2X2_2102 ( .A(w_mem_inst__abc_21203_new_n2144_), .B(w_mem_inst_w_mem_8__10_), .Y(w_mem_inst__abc_21203_new_n2145_));
OR2X2 OR2X2_2103 ( .A(w_mem_inst__abc_21203_new_n2146_), .B(w_mem_inst_w_mem_13__10_), .Y(w_mem_inst__abc_21203_new_n2147_));
OR2X2 OR2X2_2104 ( .A(w_mem_inst_w_mem_2__10_), .B(w_mem_inst_w_mem_0__10_), .Y(w_mem_inst__abc_21203_new_n2150_));
OR2X2 OR2X2_2105 ( .A(w_mem_inst__abc_21203_new_n2149_), .B(w_mem_inst__abc_21203_new_n2153_), .Y(w_mem_inst__abc_21203_new_n2154_));
OR2X2 OR2X2_2106 ( .A(w_mem_inst__abc_21203_new_n2155_), .B(w_mem_inst__abc_21203_new_n2148_), .Y(w_mem_inst__abc_21203_new_n2156_));
OR2X2 OR2X2_2107 ( .A(w_mem_inst__abc_21203_new_n2157_), .B(w_mem_inst__abc_21203_new_n1587_), .Y(w_mem_inst__abc_21203_new_n2158_));
OR2X2 OR2X2_2108 ( .A(w_mem_inst__abc_21203_new_n2159_), .B(w_mem_inst__abc_21203_new_n1586_), .Y(w_mem_inst__abc_21203_new_n2160_));
OR2X2 OR2X2_2109 ( .A(w_mem_inst__abc_21203_new_n2161_), .B(w_mem_inst__abc_21203_new_n2162_), .Y(w_mem_inst__abc_21203_new_n2163_));
OR2X2 OR2X2_211 ( .A(_abc_15497_new_n1374_), .B(_abc_15497_new_n1371_), .Y(_abc_15497_new_n1375_));
OR2X2 OR2X2_2110 ( .A(w_mem_inst__abc_21203_new_n2163_), .B(w_mem_inst__abc_21203_new_n2160_), .Y(w_mem_inst__abc_21203_new_n2164_));
OR2X2 OR2X2_2111 ( .A(w_mem_inst__abc_21203_new_n2165_), .B(w_mem_inst__abc_21203_new_n2166_), .Y(w_mem_inst__abc_21203_new_n2167_));
OR2X2 OR2X2_2112 ( .A(w_mem_inst__abc_21203_new_n2164_), .B(w_mem_inst__abc_21203_new_n2167_), .Y(w_mem_inst__abc_21203_new_n2168_));
OR2X2 OR2X2_2113 ( .A(w_mem_inst__abc_21203_new_n2170_), .B(w_mem_inst__abc_21203_new_n2171_), .Y(w_mem_inst__abc_21203_new_n2172_));
OR2X2 OR2X2_2114 ( .A(w_mem_inst__abc_21203_new_n2172_), .B(w_mem_inst__abc_21203_new_n2169_), .Y(w_mem_inst__abc_21203_new_n2173_));
OR2X2 OR2X2_2115 ( .A(w_mem_inst__abc_21203_new_n2174_), .B(w_mem_inst__abc_21203_new_n2175_), .Y(w_mem_inst__abc_21203_new_n2176_));
OR2X2 OR2X2_2116 ( .A(w_mem_inst__abc_21203_new_n2177_), .B(w_mem_inst__abc_21203_new_n2178_), .Y(w_mem_inst__abc_21203_new_n2179_));
OR2X2 OR2X2_2117 ( .A(w_mem_inst__abc_21203_new_n2176_), .B(w_mem_inst__abc_21203_new_n2179_), .Y(w_mem_inst__abc_21203_new_n2180_));
OR2X2 OR2X2_2118 ( .A(w_mem_inst__abc_21203_new_n2181_), .B(w_mem_inst__abc_21203_new_n2182_), .Y(w_mem_inst__abc_21203_new_n2183_));
OR2X2 OR2X2_2119 ( .A(w_mem_inst__abc_21203_new_n2184_), .B(w_mem_inst__abc_21203_new_n2185_), .Y(w_mem_inst__abc_21203_new_n2186_));
OR2X2 OR2X2_212 ( .A(_abc_15497_new_n699_), .B(\digest[23] ), .Y(_abc_15497_new_n1377_));
OR2X2 OR2X2_2120 ( .A(w_mem_inst__abc_21203_new_n2183_), .B(w_mem_inst__abc_21203_new_n2186_), .Y(w_mem_inst__abc_21203_new_n2187_));
OR2X2 OR2X2_2121 ( .A(w_mem_inst__abc_21203_new_n2180_), .B(w_mem_inst__abc_21203_new_n2187_), .Y(w_mem_inst__abc_21203_new_n2188_));
OR2X2 OR2X2_2122 ( .A(w_mem_inst__abc_21203_new_n2188_), .B(w_mem_inst__abc_21203_new_n2173_), .Y(w_mem_inst__abc_21203_new_n2189_));
OR2X2 OR2X2_2123 ( .A(w_mem_inst__abc_21203_new_n2189_), .B(w_mem_inst__abc_21203_new_n2168_), .Y(w_mem_inst__abc_21203_new_n2190_));
OR2X2 OR2X2_2124 ( .A(w_mem_inst__abc_21203_new_n2192_), .B(w_mem_inst_w_mem_8__11_), .Y(w_mem_inst__abc_21203_new_n2193_));
OR2X2 OR2X2_2125 ( .A(w_mem_inst__abc_21203_new_n2194_), .B(w_mem_inst_w_mem_13__11_), .Y(w_mem_inst__abc_21203_new_n2195_));
OR2X2 OR2X2_2126 ( .A(w_mem_inst_w_mem_2__11_), .B(w_mem_inst_w_mem_0__11_), .Y(w_mem_inst__abc_21203_new_n2198_));
OR2X2 OR2X2_2127 ( .A(w_mem_inst__abc_21203_new_n2197_), .B(w_mem_inst__abc_21203_new_n2201_), .Y(w_mem_inst__abc_21203_new_n2202_));
OR2X2 OR2X2_2128 ( .A(w_mem_inst__abc_21203_new_n2203_), .B(w_mem_inst__abc_21203_new_n2196_), .Y(w_mem_inst__abc_21203_new_n2204_));
OR2X2 OR2X2_2129 ( .A(w_mem_inst__abc_21203_new_n2205_), .B(w_mem_inst__abc_21203_new_n1587_), .Y(w_mem_inst__abc_21203_new_n2206_));
OR2X2 OR2X2_213 ( .A(_abc_15497_new_n1376_), .B(_abc_15497_new_n1378_), .Y(_0H4_reg_31_0__23_));
OR2X2 OR2X2_2130 ( .A(w_mem_inst__abc_21203_new_n2207_), .B(w_mem_inst__abc_21203_new_n1586_), .Y(w_mem_inst__abc_21203_new_n2208_));
OR2X2 OR2X2_2131 ( .A(w_mem_inst__abc_21203_new_n2209_), .B(w_mem_inst__abc_21203_new_n2210_), .Y(w_mem_inst__abc_21203_new_n2211_));
OR2X2 OR2X2_2132 ( .A(w_mem_inst__abc_21203_new_n2211_), .B(w_mem_inst__abc_21203_new_n2208_), .Y(w_mem_inst__abc_21203_new_n2212_));
OR2X2 OR2X2_2133 ( .A(w_mem_inst__abc_21203_new_n2213_), .B(w_mem_inst__abc_21203_new_n2214_), .Y(w_mem_inst__abc_21203_new_n2215_));
OR2X2 OR2X2_2134 ( .A(w_mem_inst__abc_21203_new_n2212_), .B(w_mem_inst__abc_21203_new_n2215_), .Y(w_mem_inst__abc_21203_new_n2216_));
OR2X2 OR2X2_2135 ( .A(w_mem_inst__abc_21203_new_n2218_), .B(w_mem_inst__abc_21203_new_n2219_), .Y(w_mem_inst__abc_21203_new_n2220_));
OR2X2 OR2X2_2136 ( .A(w_mem_inst__abc_21203_new_n2220_), .B(w_mem_inst__abc_21203_new_n2217_), .Y(w_mem_inst__abc_21203_new_n2221_));
OR2X2 OR2X2_2137 ( .A(w_mem_inst__abc_21203_new_n2222_), .B(w_mem_inst__abc_21203_new_n2223_), .Y(w_mem_inst__abc_21203_new_n2224_));
OR2X2 OR2X2_2138 ( .A(w_mem_inst__abc_21203_new_n2225_), .B(w_mem_inst__abc_21203_new_n2226_), .Y(w_mem_inst__abc_21203_new_n2227_));
OR2X2 OR2X2_2139 ( .A(w_mem_inst__abc_21203_new_n2224_), .B(w_mem_inst__abc_21203_new_n2227_), .Y(w_mem_inst__abc_21203_new_n2228_));
OR2X2 OR2X2_214 ( .A(_abc_15497_new_n1383_), .B(_abc_15497_new_n1368_), .Y(_abc_15497_new_n1384_));
OR2X2 OR2X2_2140 ( .A(w_mem_inst__abc_21203_new_n2229_), .B(w_mem_inst__abc_21203_new_n2230_), .Y(w_mem_inst__abc_21203_new_n2231_));
OR2X2 OR2X2_2141 ( .A(w_mem_inst__abc_21203_new_n2232_), .B(w_mem_inst__abc_21203_new_n2233_), .Y(w_mem_inst__abc_21203_new_n2234_));
OR2X2 OR2X2_2142 ( .A(w_mem_inst__abc_21203_new_n2231_), .B(w_mem_inst__abc_21203_new_n2234_), .Y(w_mem_inst__abc_21203_new_n2235_));
OR2X2 OR2X2_2143 ( .A(w_mem_inst__abc_21203_new_n2228_), .B(w_mem_inst__abc_21203_new_n2235_), .Y(w_mem_inst__abc_21203_new_n2236_));
OR2X2 OR2X2_2144 ( .A(w_mem_inst__abc_21203_new_n2236_), .B(w_mem_inst__abc_21203_new_n2221_), .Y(w_mem_inst__abc_21203_new_n2237_));
OR2X2 OR2X2_2145 ( .A(w_mem_inst__abc_21203_new_n2237_), .B(w_mem_inst__abc_21203_new_n2216_), .Y(w_mem_inst__abc_21203_new_n2238_));
OR2X2 OR2X2_2146 ( .A(w_mem_inst__abc_21203_new_n2240_), .B(w_mem_inst_w_mem_8__12_), .Y(w_mem_inst__abc_21203_new_n2241_));
OR2X2 OR2X2_2147 ( .A(w_mem_inst__abc_21203_new_n2242_), .B(w_mem_inst_w_mem_13__12_), .Y(w_mem_inst__abc_21203_new_n2243_));
OR2X2 OR2X2_2148 ( .A(w_mem_inst_w_mem_2__12_), .B(w_mem_inst_w_mem_0__12_), .Y(w_mem_inst__abc_21203_new_n2246_));
OR2X2 OR2X2_2149 ( .A(w_mem_inst__abc_21203_new_n2245_), .B(w_mem_inst__abc_21203_new_n2249_), .Y(w_mem_inst__abc_21203_new_n2250_));
OR2X2 OR2X2_215 ( .A(_abc_15497_new_n1386_), .B(_abc_15497_new_n1384_), .Y(_abc_15497_new_n1387_));
OR2X2 OR2X2_2150 ( .A(w_mem_inst__abc_21203_new_n2251_), .B(w_mem_inst__abc_21203_new_n2244_), .Y(w_mem_inst__abc_21203_new_n2252_));
OR2X2 OR2X2_2151 ( .A(w_mem_inst__abc_21203_new_n2253_), .B(w_mem_inst__abc_21203_new_n1587_), .Y(w_mem_inst__abc_21203_new_n2254_));
OR2X2 OR2X2_2152 ( .A(w_mem_inst__abc_21203_new_n2255_), .B(w_mem_inst__abc_21203_new_n1586_), .Y(w_mem_inst__abc_21203_new_n2256_));
OR2X2 OR2X2_2153 ( .A(w_mem_inst__abc_21203_new_n2257_), .B(w_mem_inst__abc_21203_new_n2258_), .Y(w_mem_inst__abc_21203_new_n2259_));
OR2X2 OR2X2_2154 ( .A(w_mem_inst__abc_21203_new_n2259_), .B(w_mem_inst__abc_21203_new_n2256_), .Y(w_mem_inst__abc_21203_new_n2260_));
OR2X2 OR2X2_2155 ( .A(w_mem_inst__abc_21203_new_n2261_), .B(w_mem_inst__abc_21203_new_n2262_), .Y(w_mem_inst__abc_21203_new_n2263_));
OR2X2 OR2X2_2156 ( .A(w_mem_inst__abc_21203_new_n2260_), .B(w_mem_inst__abc_21203_new_n2263_), .Y(w_mem_inst__abc_21203_new_n2264_));
OR2X2 OR2X2_2157 ( .A(w_mem_inst__abc_21203_new_n2266_), .B(w_mem_inst__abc_21203_new_n2267_), .Y(w_mem_inst__abc_21203_new_n2268_));
OR2X2 OR2X2_2158 ( .A(w_mem_inst__abc_21203_new_n2268_), .B(w_mem_inst__abc_21203_new_n2265_), .Y(w_mem_inst__abc_21203_new_n2269_));
OR2X2 OR2X2_2159 ( .A(w_mem_inst__abc_21203_new_n2270_), .B(w_mem_inst__abc_21203_new_n2271_), .Y(w_mem_inst__abc_21203_new_n2272_));
OR2X2 OR2X2_216 ( .A(_abc_15497_new_n1382_), .B(_abc_15497_new_n1387_), .Y(_abc_15497_new_n1388_));
OR2X2 OR2X2_2160 ( .A(w_mem_inst__abc_21203_new_n2273_), .B(w_mem_inst__abc_21203_new_n2274_), .Y(w_mem_inst__abc_21203_new_n2275_));
OR2X2 OR2X2_2161 ( .A(w_mem_inst__abc_21203_new_n2272_), .B(w_mem_inst__abc_21203_new_n2275_), .Y(w_mem_inst__abc_21203_new_n2276_));
OR2X2 OR2X2_2162 ( .A(w_mem_inst__abc_21203_new_n2277_), .B(w_mem_inst__abc_21203_new_n2278_), .Y(w_mem_inst__abc_21203_new_n2279_));
OR2X2 OR2X2_2163 ( .A(w_mem_inst__abc_21203_new_n2280_), .B(w_mem_inst__abc_21203_new_n2281_), .Y(w_mem_inst__abc_21203_new_n2282_));
OR2X2 OR2X2_2164 ( .A(w_mem_inst__abc_21203_new_n2279_), .B(w_mem_inst__abc_21203_new_n2282_), .Y(w_mem_inst__abc_21203_new_n2283_));
OR2X2 OR2X2_2165 ( .A(w_mem_inst__abc_21203_new_n2276_), .B(w_mem_inst__abc_21203_new_n2283_), .Y(w_mem_inst__abc_21203_new_n2284_));
OR2X2 OR2X2_2166 ( .A(w_mem_inst__abc_21203_new_n2284_), .B(w_mem_inst__abc_21203_new_n2269_), .Y(w_mem_inst__abc_21203_new_n2285_));
OR2X2 OR2X2_2167 ( .A(w_mem_inst__abc_21203_new_n2285_), .B(w_mem_inst__abc_21203_new_n2264_), .Y(w_mem_inst__abc_21203_new_n2286_));
OR2X2 OR2X2_2168 ( .A(w_mem_inst__abc_21203_new_n2288_), .B(w_mem_inst_w_mem_8__13_), .Y(w_mem_inst__abc_21203_new_n2289_));
OR2X2 OR2X2_2169 ( .A(w_mem_inst__abc_21203_new_n2290_), .B(w_mem_inst_w_mem_13__13_), .Y(w_mem_inst__abc_21203_new_n2291_));
OR2X2 OR2X2_217 ( .A(_abc_15497_new_n1390_), .B(_abc_15497_new_n1388_), .Y(_abc_15497_new_n1391_));
OR2X2 OR2X2_2170 ( .A(w_mem_inst_w_mem_2__13_), .B(w_mem_inst_w_mem_0__13_), .Y(w_mem_inst__abc_21203_new_n2294_));
OR2X2 OR2X2_2171 ( .A(w_mem_inst__abc_21203_new_n2293_), .B(w_mem_inst__abc_21203_new_n2297_), .Y(w_mem_inst__abc_21203_new_n2298_));
OR2X2 OR2X2_2172 ( .A(w_mem_inst__abc_21203_new_n2299_), .B(w_mem_inst__abc_21203_new_n2292_), .Y(w_mem_inst__abc_21203_new_n2300_));
OR2X2 OR2X2_2173 ( .A(w_mem_inst__abc_21203_new_n2301_), .B(w_mem_inst__abc_21203_new_n1587_), .Y(w_mem_inst__abc_21203_new_n2302_));
OR2X2 OR2X2_2174 ( .A(w_mem_inst__abc_21203_new_n2303_), .B(w_mem_inst__abc_21203_new_n1586_), .Y(w_mem_inst__abc_21203_new_n2304_));
OR2X2 OR2X2_2175 ( .A(w_mem_inst__abc_21203_new_n2305_), .B(w_mem_inst__abc_21203_new_n2306_), .Y(w_mem_inst__abc_21203_new_n2307_));
OR2X2 OR2X2_2176 ( .A(w_mem_inst__abc_21203_new_n2307_), .B(w_mem_inst__abc_21203_new_n2304_), .Y(w_mem_inst__abc_21203_new_n2308_));
OR2X2 OR2X2_2177 ( .A(w_mem_inst__abc_21203_new_n2309_), .B(w_mem_inst__abc_21203_new_n2310_), .Y(w_mem_inst__abc_21203_new_n2311_));
OR2X2 OR2X2_2178 ( .A(w_mem_inst__abc_21203_new_n2308_), .B(w_mem_inst__abc_21203_new_n2311_), .Y(w_mem_inst__abc_21203_new_n2312_));
OR2X2 OR2X2_2179 ( .A(w_mem_inst__abc_21203_new_n2314_), .B(w_mem_inst__abc_21203_new_n2315_), .Y(w_mem_inst__abc_21203_new_n2316_));
OR2X2 OR2X2_218 ( .A(e_reg_24_), .B(\digest[24] ), .Y(_abc_15497_new_n1392_));
OR2X2 OR2X2_2180 ( .A(w_mem_inst__abc_21203_new_n2316_), .B(w_mem_inst__abc_21203_new_n2313_), .Y(w_mem_inst__abc_21203_new_n2317_));
OR2X2 OR2X2_2181 ( .A(w_mem_inst__abc_21203_new_n2318_), .B(w_mem_inst__abc_21203_new_n2319_), .Y(w_mem_inst__abc_21203_new_n2320_));
OR2X2 OR2X2_2182 ( .A(w_mem_inst__abc_21203_new_n2321_), .B(w_mem_inst__abc_21203_new_n2322_), .Y(w_mem_inst__abc_21203_new_n2323_));
OR2X2 OR2X2_2183 ( .A(w_mem_inst__abc_21203_new_n2320_), .B(w_mem_inst__abc_21203_new_n2323_), .Y(w_mem_inst__abc_21203_new_n2324_));
OR2X2 OR2X2_2184 ( .A(w_mem_inst__abc_21203_new_n2325_), .B(w_mem_inst__abc_21203_new_n2326_), .Y(w_mem_inst__abc_21203_new_n2327_));
OR2X2 OR2X2_2185 ( .A(w_mem_inst__abc_21203_new_n2328_), .B(w_mem_inst__abc_21203_new_n2329_), .Y(w_mem_inst__abc_21203_new_n2330_));
OR2X2 OR2X2_2186 ( .A(w_mem_inst__abc_21203_new_n2327_), .B(w_mem_inst__abc_21203_new_n2330_), .Y(w_mem_inst__abc_21203_new_n2331_));
OR2X2 OR2X2_2187 ( .A(w_mem_inst__abc_21203_new_n2324_), .B(w_mem_inst__abc_21203_new_n2331_), .Y(w_mem_inst__abc_21203_new_n2332_));
OR2X2 OR2X2_2188 ( .A(w_mem_inst__abc_21203_new_n2332_), .B(w_mem_inst__abc_21203_new_n2317_), .Y(w_mem_inst__abc_21203_new_n2333_));
OR2X2 OR2X2_2189 ( .A(w_mem_inst__abc_21203_new_n2333_), .B(w_mem_inst__abc_21203_new_n2312_), .Y(w_mem_inst__abc_21203_new_n2334_));
OR2X2 OR2X2_219 ( .A(_abc_15497_new_n1391_), .B(_abc_15497_new_n1395_), .Y(_abc_15497_new_n1396_));
OR2X2 OR2X2_2190 ( .A(w_mem_inst__abc_21203_new_n2336_), .B(w_mem_inst_w_mem_8__14_), .Y(w_mem_inst__abc_21203_new_n2337_));
OR2X2 OR2X2_2191 ( .A(w_mem_inst__abc_21203_new_n2338_), .B(w_mem_inst_w_mem_13__14_), .Y(w_mem_inst__abc_21203_new_n2339_));
OR2X2 OR2X2_2192 ( .A(w_mem_inst_w_mem_2__14_), .B(w_mem_inst_w_mem_0__14_), .Y(w_mem_inst__abc_21203_new_n2342_));
OR2X2 OR2X2_2193 ( .A(w_mem_inst__abc_21203_new_n2341_), .B(w_mem_inst__abc_21203_new_n2345_), .Y(w_mem_inst__abc_21203_new_n2346_));
OR2X2 OR2X2_2194 ( .A(w_mem_inst__abc_21203_new_n2347_), .B(w_mem_inst__abc_21203_new_n2340_), .Y(w_mem_inst__abc_21203_new_n2348_));
OR2X2 OR2X2_2195 ( .A(w_mem_inst__abc_21203_new_n2349_), .B(w_mem_inst__abc_21203_new_n1587_), .Y(w_mem_inst__abc_21203_new_n2350_));
OR2X2 OR2X2_2196 ( .A(w_mem_inst__abc_21203_new_n2351_), .B(w_mem_inst__abc_21203_new_n1586_), .Y(w_mem_inst__abc_21203_new_n2352_));
OR2X2 OR2X2_2197 ( .A(w_mem_inst__abc_21203_new_n2353_), .B(w_mem_inst__abc_21203_new_n2354_), .Y(w_mem_inst__abc_21203_new_n2355_));
OR2X2 OR2X2_2198 ( .A(w_mem_inst__abc_21203_new_n2355_), .B(w_mem_inst__abc_21203_new_n2352_), .Y(w_mem_inst__abc_21203_new_n2356_));
OR2X2 OR2X2_2199 ( .A(w_mem_inst__abc_21203_new_n2357_), .B(w_mem_inst__abc_21203_new_n2358_), .Y(w_mem_inst__abc_21203_new_n2359_));
OR2X2 OR2X2_22 ( .A(_abc_15497_new_n788_), .B(_abc_15497_new_n785_), .Y(_abc_15497_new_n789_));
OR2X2 OR2X2_220 ( .A(_abc_15497_new_n699_), .B(\digest[24] ), .Y(_abc_15497_new_n1401_));
OR2X2 OR2X2_2200 ( .A(w_mem_inst__abc_21203_new_n2356_), .B(w_mem_inst__abc_21203_new_n2359_), .Y(w_mem_inst__abc_21203_new_n2360_));
OR2X2 OR2X2_2201 ( .A(w_mem_inst__abc_21203_new_n2362_), .B(w_mem_inst__abc_21203_new_n2363_), .Y(w_mem_inst__abc_21203_new_n2364_));
OR2X2 OR2X2_2202 ( .A(w_mem_inst__abc_21203_new_n2364_), .B(w_mem_inst__abc_21203_new_n2361_), .Y(w_mem_inst__abc_21203_new_n2365_));
OR2X2 OR2X2_2203 ( .A(w_mem_inst__abc_21203_new_n2366_), .B(w_mem_inst__abc_21203_new_n2367_), .Y(w_mem_inst__abc_21203_new_n2368_));
OR2X2 OR2X2_2204 ( .A(w_mem_inst__abc_21203_new_n2369_), .B(w_mem_inst__abc_21203_new_n2370_), .Y(w_mem_inst__abc_21203_new_n2371_));
OR2X2 OR2X2_2205 ( .A(w_mem_inst__abc_21203_new_n2368_), .B(w_mem_inst__abc_21203_new_n2371_), .Y(w_mem_inst__abc_21203_new_n2372_));
OR2X2 OR2X2_2206 ( .A(w_mem_inst__abc_21203_new_n2373_), .B(w_mem_inst__abc_21203_new_n2374_), .Y(w_mem_inst__abc_21203_new_n2375_));
OR2X2 OR2X2_2207 ( .A(w_mem_inst__abc_21203_new_n2376_), .B(w_mem_inst__abc_21203_new_n2377_), .Y(w_mem_inst__abc_21203_new_n2378_));
OR2X2 OR2X2_2208 ( .A(w_mem_inst__abc_21203_new_n2375_), .B(w_mem_inst__abc_21203_new_n2378_), .Y(w_mem_inst__abc_21203_new_n2379_));
OR2X2 OR2X2_2209 ( .A(w_mem_inst__abc_21203_new_n2372_), .B(w_mem_inst__abc_21203_new_n2379_), .Y(w_mem_inst__abc_21203_new_n2380_));
OR2X2 OR2X2_221 ( .A(_abc_15497_new_n1400_), .B(_abc_15497_new_n1402_), .Y(_0H4_reg_31_0__24_));
OR2X2 OR2X2_2210 ( .A(w_mem_inst__abc_21203_new_n2380_), .B(w_mem_inst__abc_21203_new_n2365_), .Y(w_mem_inst__abc_21203_new_n2381_));
OR2X2 OR2X2_2211 ( .A(w_mem_inst__abc_21203_new_n2381_), .B(w_mem_inst__abc_21203_new_n2360_), .Y(w_mem_inst__abc_21203_new_n2382_));
OR2X2 OR2X2_2212 ( .A(w_mem_inst__abc_21203_new_n2384_), .B(w_mem_inst_w_mem_8__15_), .Y(w_mem_inst__abc_21203_new_n2385_));
OR2X2 OR2X2_2213 ( .A(w_mem_inst__abc_21203_new_n2386_), .B(w_mem_inst_w_mem_13__15_), .Y(w_mem_inst__abc_21203_new_n2387_));
OR2X2 OR2X2_2214 ( .A(w_mem_inst_w_mem_2__15_), .B(w_mem_inst_w_mem_0__15_), .Y(w_mem_inst__abc_21203_new_n2390_));
OR2X2 OR2X2_2215 ( .A(w_mem_inst__abc_21203_new_n2389_), .B(w_mem_inst__abc_21203_new_n2393_), .Y(w_mem_inst__abc_21203_new_n2394_));
OR2X2 OR2X2_2216 ( .A(w_mem_inst__abc_21203_new_n2395_), .B(w_mem_inst__abc_21203_new_n2388_), .Y(w_mem_inst__abc_21203_new_n2396_));
OR2X2 OR2X2_2217 ( .A(w_mem_inst__abc_21203_new_n2397_), .B(w_mem_inst__abc_21203_new_n1587_), .Y(w_mem_inst__abc_21203_new_n2398_));
OR2X2 OR2X2_2218 ( .A(w_mem_inst__abc_21203_new_n2399_), .B(w_mem_inst__abc_21203_new_n1586_), .Y(w_mem_inst__abc_21203_new_n2400_));
OR2X2 OR2X2_2219 ( .A(w_mem_inst__abc_21203_new_n2401_), .B(w_mem_inst__abc_21203_new_n2402_), .Y(w_mem_inst__abc_21203_new_n2403_));
OR2X2 OR2X2_222 ( .A(e_reg_25_), .B(\digest[25] ), .Y(_abc_15497_new_n1406_));
OR2X2 OR2X2_2220 ( .A(w_mem_inst__abc_21203_new_n2403_), .B(w_mem_inst__abc_21203_new_n2400_), .Y(w_mem_inst__abc_21203_new_n2404_));
OR2X2 OR2X2_2221 ( .A(w_mem_inst__abc_21203_new_n2405_), .B(w_mem_inst__abc_21203_new_n2406_), .Y(w_mem_inst__abc_21203_new_n2407_));
OR2X2 OR2X2_2222 ( .A(w_mem_inst__abc_21203_new_n2404_), .B(w_mem_inst__abc_21203_new_n2407_), .Y(w_mem_inst__abc_21203_new_n2408_));
OR2X2 OR2X2_2223 ( .A(w_mem_inst__abc_21203_new_n2410_), .B(w_mem_inst__abc_21203_new_n2411_), .Y(w_mem_inst__abc_21203_new_n2412_));
OR2X2 OR2X2_2224 ( .A(w_mem_inst__abc_21203_new_n2412_), .B(w_mem_inst__abc_21203_new_n2409_), .Y(w_mem_inst__abc_21203_new_n2413_));
OR2X2 OR2X2_2225 ( .A(w_mem_inst__abc_21203_new_n2414_), .B(w_mem_inst__abc_21203_new_n2415_), .Y(w_mem_inst__abc_21203_new_n2416_));
OR2X2 OR2X2_2226 ( .A(w_mem_inst__abc_21203_new_n2417_), .B(w_mem_inst__abc_21203_new_n2418_), .Y(w_mem_inst__abc_21203_new_n2419_));
OR2X2 OR2X2_2227 ( .A(w_mem_inst__abc_21203_new_n2416_), .B(w_mem_inst__abc_21203_new_n2419_), .Y(w_mem_inst__abc_21203_new_n2420_));
OR2X2 OR2X2_2228 ( .A(w_mem_inst__abc_21203_new_n2421_), .B(w_mem_inst__abc_21203_new_n2422_), .Y(w_mem_inst__abc_21203_new_n2423_));
OR2X2 OR2X2_2229 ( .A(w_mem_inst__abc_21203_new_n2424_), .B(w_mem_inst__abc_21203_new_n2425_), .Y(w_mem_inst__abc_21203_new_n2426_));
OR2X2 OR2X2_223 ( .A(_abc_15497_new_n1405_), .B(_abc_15497_new_n1409_), .Y(_abc_15497_new_n1410_));
OR2X2 OR2X2_2230 ( .A(w_mem_inst__abc_21203_new_n2423_), .B(w_mem_inst__abc_21203_new_n2426_), .Y(w_mem_inst__abc_21203_new_n2427_));
OR2X2 OR2X2_2231 ( .A(w_mem_inst__abc_21203_new_n2420_), .B(w_mem_inst__abc_21203_new_n2427_), .Y(w_mem_inst__abc_21203_new_n2428_));
OR2X2 OR2X2_2232 ( .A(w_mem_inst__abc_21203_new_n2428_), .B(w_mem_inst__abc_21203_new_n2413_), .Y(w_mem_inst__abc_21203_new_n2429_));
OR2X2 OR2X2_2233 ( .A(w_mem_inst__abc_21203_new_n2429_), .B(w_mem_inst__abc_21203_new_n2408_), .Y(w_mem_inst__abc_21203_new_n2430_));
OR2X2 OR2X2_2234 ( .A(w_mem_inst__abc_21203_new_n2432_), .B(w_mem_inst_w_mem_8__16_), .Y(w_mem_inst__abc_21203_new_n2433_));
OR2X2 OR2X2_2235 ( .A(w_mem_inst__abc_21203_new_n2434_), .B(w_mem_inst_w_mem_13__16_), .Y(w_mem_inst__abc_21203_new_n2435_));
OR2X2 OR2X2_2236 ( .A(w_mem_inst_w_mem_2__16_), .B(w_mem_inst_w_mem_0__16_), .Y(w_mem_inst__abc_21203_new_n2438_));
OR2X2 OR2X2_2237 ( .A(w_mem_inst__abc_21203_new_n2437_), .B(w_mem_inst__abc_21203_new_n2441_), .Y(w_mem_inst__abc_21203_new_n2442_));
OR2X2 OR2X2_2238 ( .A(w_mem_inst__abc_21203_new_n2443_), .B(w_mem_inst__abc_21203_new_n2436_), .Y(w_mem_inst__abc_21203_new_n2444_));
OR2X2 OR2X2_2239 ( .A(w_mem_inst__abc_21203_new_n2445_), .B(w_mem_inst__abc_21203_new_n1587_), .Y(w_mem_inst__abc_21203_new_n2446_));
OR2X2 OR2X2_224 ( .A(_abc_15497_new_n1404_), .B(_abc_15497_new_n1411_), .Y(_abc_15497_new_n1412_));
OR2X2 OR2X2_2240 ( .A(w_mem_inst__abc_21203_new_n2447_), .B(w_mem_inst__abc_21203_new_n1586_), .Y(w_mem_inst__abc_21203_new_n2448_));
OR2X2 OR2X2_2241 ( .A(w_mem_inst__abc_21203_new_n2449_), .B(w_mem_inst__abc_21203_new_n2450_), .Y(w_mem_inst__abc_21203_new_n2451_));
OR2X2 OR2X2_2242 ( .A(w_mem_inst__abc_21203_new_n2451_), .B(w_mem_inst__abc_21203_new_n2448_), .Y(w_mem_inst__abc_21203_new_n2452_));
OR2X2 OR2X2_2243 ( .A(w_mem_inst__abc_21203_new_n2453_), .B(w_mem_inst__abc_21203_new_n2454_), .Y(w_mem_inst__abc_21203_new_n2455_));
OR2X2 OR2X2_2244 ( .A(w_mem_inst__abc_21203_new_n2452_), .B(w_mem_inst__abc_21203_new_n2455_), .Y(w_mem_inst__abc_21203_new_n2456_));
OR2X2 OR2X2_2245 ( .A(w_mem_inst__abc_21203_new_n2458_), .B(w_mem_inst__abc_21203_new_n2459_), .Y(w_mem_inst__abc_21203_new_n2460_));
OR2X2 OR2X2_2246 ( .A(w_mem_inst__abc_21203_new_n2460_), .B(w_mem_inst__abc_21203_new_n2457_), .Y(w_mem_inst__abc_21203_new_n2461_));
OR2X2 OR2X2_2247 ( .A(w_mem_inst__abc_21203_new_n2462_), .B(w_mem_inst__abc_21203_new_n2463_), .Y(w_mem_inst__abc_21203_new_n2464_));
OR2X2 OR2X2_2248 ( .A(w_mem_inst__abc_21203_new_n2465_), .B(w_mem_inst__abc_21203_new_n2466_), .Y(w_mem_inst__abc_21203_new_n2467_));
OR2X2 OR2X2_2249 ( .A(w_mem_inst__abc_21203_new_n2464_), .B(w_mem_inst__abc_21203_new_n2467_), .Y(w_mem_inst__abc_21203_new_n2468_));
OR2X2 OR2X2_225 ( .A(_abc_15497_new_n699_), .B(\digest[25] ), .Y(_abc_15497_new_n1415_));
OR2X2 OR2X2_2250 ( .A(w_mem_inst__abc_21203_new_n2469_), .B(w_mem_inst__abc_21203_new_n2470_), .Y(w_mem_inst__abc_21203_new_n2471_));
OR2X2 OR2X2_2251 ( .A(w_mem_inst__abc_21203_new_n2472_), .B(w_mem_inst__abc_21203_new_n2473_), .Y(w_mem_inst__abc_21203_new_n2474_));
OR2X2 OR2X2_2252 ( .A(w_mem_inst__abc_21203_new_n2471_), .B(w_mem_inst__abc_21203_new_n2474_), .Y(w_mem_inst__abc_21203_new_n2475_));
OR2X2 OR2X2_2253 ( .A(w_mem_inst__abc_21203_new_n2468_), .B(w_mem_inst__abc_21203_new_n2475_), .Y(w_mem_inst__abc_21203_new_n2476_));
OR2X2 OR2X2_2254 ( .A(w_mem_inst__abc_21203_new_n2476_), .B(w_mem_inst__abc_21203_new_n2461_), .Y(w_mem_inst__abc_21203_new_n2477_));
OR2X2 OR2X2_2255 ( .A(w_mem_inst__abc_21203_new_n2477_), .B(w_mem_inst__abc_21203_new_n2456_), .Y(w_mem_inst__abc_21203_new_n2478_));
OR2X2 OR2X2_2256 ( .A(w_mem_inst__abc_21203_new_n2480_), .B(w_mem_inst_w_mem_8__17_), .Y(w_mem_inst__abc_21203_new_n2481_));
OR2X2 OR2X2_2257 ( .A(w_mem_inst__abc_21203_new_n2482_), .B(w_mem_inst_w_mem_13__17_), .Y(w_mem_inst__abc_21203_new_n2483_));
OR2X2 OR2X2_2258 ( .A(w_mem_inst_w_mem_2__17_), .B(w_mem_inst_w_mem_0__17_), .Y(w_mem_inst__abc_21203_new_n2486_));
OR2X2 OR2X2_2259 ( .A(w_mem_inst__abc_21203_new_n2485_), .B(w_mem_inst__abc_21203_new_n2489_), .Y(w_mem_inst__abc_21203_new_n2490_));
OR2X2 OR2X2_226 ( .A(_abc_15497_new_n1414_), .B(_abc_15497_new_n1416_), .Y(_0H4_reg_31_0__25_));
OR2X2 OR2X2_2260 ( .A(w_mem_inst__abc_21203_new_n2491_), .B(w_mem_inst__abc_21203_new_n2484_), .Y(w_mem_inst__abc_21203_new_n2492_));
OR2X2 OR2X2_2261 ( .A(w_mem_inst__abc_21203_new_n2493_), .B(w_mem_inst__abc_21203_new_n1587_), .Y(w_mem_inst__abc_21203_new_n2494_));
OR2X2 OR2X2_2262 ( .A(w_mem_inst__abc_21203_new_n2495_), .B(w_mem_inst__abc_21203_new_n1586_), .Y(w_mem_inst__abc_21203_new_n2496_));
OR2X2 OR2X2_2263 ( .A(w_mem_inst__abc_21203_new_n2497_), .B(w_mem_inst__abc_21203_new_n2498_), .Y(w_mem_inst__abc_21203_new_n2499_));
OR2X2 OR2X2_2264 ( .A(w_mem_inst__abc_21203_new_n2499_), .B(w_mem_inst__abc_21203_new_n2496_), .Y(w_mem_inst__abc_21203_new_n2500_));
OR2X2 OR2X2_2265 ( .A(w_mem_inst__abc_21203_new_n2501_), .B(w_mem_inst__abc_21203_new_n2502_), .Y(w_mem_inst__abc_21203_new_n2503_));
OR2X2 OR2X2_2266 ( .A(w_mem_inst__abc_21203_new_n2500_), .B(w_mem_inst__abc_21203_new_n2503_), .Y(w_mem_inst__abc_21203_new_n2504_));
OR2X2 OR2X2_2267 ( .A(w_mem_inst__abc_21203_new_n2506_), .B(w_mem_inst__abc_21203_new_n2507_), .Y(w_mem_inst__abc_21203_new_n2508_));
OR2X2 OR2X2_2268 ( .A(w_mem_inst__abc_21203_new_n2508_), .B(w_mem_inst__abc_21203_new_n2505_), .Y(w_mem_inst__abc_21203_new_n2509_));
OR2X2 OR2X2_2269 ( .A(w_mem_inst__abc_21203_new_n2510_), .B(w_mem_inst__abc_21203_new_n2511_), .Y(w_mem_inst__abc_21203_new_n2512_));
OR2X2 OR2X2_227 ( .A(_abc_15497_new_n1421_), .B(_abc_15497_new_n1407_), .Y(_abc_15497_new_n1422_));
OR2X2 OR2X2_2270 ( .A(w_mem_inst__abc_21203_new_n2513_), .B(w_mem_inst__abc_21203_new_n2514_), .Y(w_mem_inst__abc_21203_new_n2515_));
OR2X2 OR2X2_2271 ( .A(w_mem_inst__abc_21203_new_n2512_), .B(w_mem_inst__abc_21203_new_n2515_), .Y(w_mem_inst__abc_21203_new_n2516_));
OR2X2 OR2X2_2272 ( .A(w_mem_inst__abc_21203_new_n2517_), .B(w_mem_inst__abc_21203_new_n2518_), .Y(w_mem_inst__abc_21203_new_n2519_));
OR2X2 OR2X2_2273 ( .A(w_mem_inst__abc_21203_new_n2520_), .B(w_mem_inst__abc_21203_new_n2521_), .Y(w_mem_inst__abc_21203_new_n2522_));
OR2X2 OR2X2_2274 ( .A(w_mem_inst__abc_21203_new_n2519_), .B(w_mem_inst__abc_21203_new_n2522_), .Y(w_mem_inst__abc_21203_new_n2523_));
OR2X2 OR2X2_2275 ( .A(w_mem_inst__abc_21203_new_n2516_), .B(w_mem_inst__abc_21203_new_n2523_), .Y(w_mem_inst__abc_21203_new_n2524_));
OR2X2 OR2X2_2276 ( .A(w_mem_inst__abc_21203_new_n2524_), .B(w_mem_inst__abc_21203_new_n2509_), .Y(w_mem_inst__abc_21203_new_n2525_));
OR2X2 OR2X2_2277 ( .A(w_mem_inst__abc_21203_new_n2525_), .B(w_mem_inst__abc_21203_new_n2504_), .Y(w_mem_inst__abc_21203_new_n2526_));
OR2X2 OR2X2_2278 ( .A(w_mem_inst__abc_21203_new_n2528_), .B(w_mem_inst_w_mem_8__18_), .Y(w_mem_inst__abc_21203_new_n2529_));
OR2X2 OR2X2_2279 ( .A(w_mem_inst__abc_21203_new_n2530_), .B(w_mem_inst_w_mem_13__18_), .Y(w_mem_inst__abc_21203_new_n2531_));
OR2X2 OR2X2_228 ( .A(_abc_15497_new_n1420_), .B(_abc_15497_new_n1422_), .Y(_abc_15497_new_n1423_));
OR2X2 OR2X2_2280 ( .A(w_mem_inst_w_mem_2__18_), .B(w_mem_inst_w_mem_0__18_), .Y(w_mem_inst__abc_21203_new_n2534_));
OR2X2 OR2X2_2281 ( .A(w_mem_inst__abc_21203_new_n2533_), .B(w_mem_inst__abc_21203_new_n2537_), .Y(w_mem_inst__abc_21203_new_n2538_));
OR2X2 OR2X2_2282 ( .A(w_mem_inst__abc_21203_new_n2539_), .B(w_mem_inst__abc_21203_new_n2532_), .Y(w_mem_inst__abc_21203_new_n2540_));
OR2X2 OR2X2_2283 ( .A(w_mem_inst__abc_21203_new_n2541_), .B(w_mem_inst__abc_21203_new_n1587_), .Y(w_mem_inst__abc_21203_new_n2542_));
OR2X2 OR2X2_2284 ( .A(w_mem_inst__abc_21203_new_n2543_), .B(w_mem_inst__abc_21203_new_n1586_), .Y(w_mem_inst__abc_21203_new_n2544_));
OR2X2 OR2X2_2285 ( .A(w_mem_inst__abc_21203_new_n2545_), .B(w_mem_inst__abc_21203_new_n2546_), .Y(w_mem_inst__abc_21203_new_n2547_));
OR2X2 OR2X2_2286 ( .A(w_mem_inst__abc_21203_new_n2547_), .B(w_mem_inst__abc_21203_new_n2544_), .Y(w_mem_inst__abc_21203_new_n2548_));
OR2X2 OR2X2_2287 ( .A(w_mem_inst__abc_21203_new_n2549_), .B(w_mem_inst__abc_21203_new_n2550_), .Y(w_mem_inst__abc_21203_new_n2551_));
OR2X2 OR2X2_2288 ( .A(w_mem_inst__abc_21203_new_n2548_), .B(w_mem_inst__abc_21203_new_n2551_), .Y(w_mem_inst__abc_21203_new_n2552_));
OR2X2 OR2X2_2289 ( .A(w_mem_inst__abc_21203_new_n2554_), .B(w_mem_inst__abc_21203_new_n2555_), .Y(w_mem_inst__abc_21203_new_n2556_));
OR2X2 OR2X2_229 ( .A(e_reg_26_), .B(\digest[26] ), .Y(_abc_15497_new_n1424_));
OR2X2 OR2X2_2290 ( .A(w_mem_inst__abc_21203_new_n2556_), .B(w_mem_inst__abc_21203_new_n2553_), .Y(w_mem_inst__abc_21203_new_n2557_));
OR2X2 OR2X2_2291 ( .A(w_mem_inst__abc_21203_new_n2558_), .B(w_mem_inst__abc_21203_new_n2559_), .Y(w_mem_inst__abc_21203_new_n2560_));
OR2X2 OR2X2_2292 ( .A(w_mem_inst__abc_21203_new_n2561_), .B(w_mem_inst__abc_21203_new_n2562_), .Y(w_mem_inst__abc_21203_new_n2563_));
OR2X2 OR2X2_2293 ( .A(w_mem_inst__abc_21203_new_n2560_), .B(w_mem_inst__abc_21203_new_n2563_), .Y(w_mem_inst__abc_21203_new_n2564_));
OR2X2 OR2X2_2294 ( .A(w_mem_inst__abc_21203_new_n2565_), .B(w_mem_inst__abc_21203_new_n2566_), .Y(w_mem_inst__abc_21203_new_n2567_));
OR2X2 OR2X2_2295 ( .A(w_mem_inst__abc_21203_new_n2568_), .B(w_mem_inst__abc_21203_new_n2569_), .Y(w_mem_inst__abc_21203_new_n2570_));
OR2X2 OR2X2_2296 ( .A(w_mem_inst__abc_21203_new_n2567_), .B(w_mem_inst__abc_21203_new_n2570_), .Y(w_mem_inst__abc_21203_new_n2571_));
OR2X2 OR2X2_2297 ( .A(w_mem_inst__abc_21203_new_n2564_), .B(w_mem_inst__abc_21203_new_n2571_), .Y(w_mem_inst__abc_21203_new_n2572_));
OR2X2 OR2X2_2298 ( .A(w_mem_inst__abc_21203_new_n2572_), .B(w_mem_inst__abc_21203_new_n2557_), .Y(w_mem_inst__abc_21203_new_n2573_));
OR2X2 OR2X2_2299 ( .A(w_mem_inst__abc_21203_new_n2573_), .B(w_mem_inst__abc_21203_new_n2552_), .Y(w_mem_inst__abc_21203_new_n2574_));
OR2X2 OR2X2_23 ( .A(c_reg_10_), .B(\digest[74] ), .Y(_abc_15497_new_n793_));
OR2X2 OR2X2_230 ( .A(_abc_15497_new_n1423_), .B(_abc_15497_new_n1427_), .Y(_abc_15497_new_n1428_));
OR2X2 OR2X2_2300 ( .A(w_mem_inst__abc_21203_new_n2576_), .B(w_mem_inst_w_mem_8__19_), .Y(w_mem_inst__abc_21203_new_n2577_));
OR2X2 OR2X2_2301 ( .A(w_mem_inst__abc_21203_new_n2578_), .B(w_mem_inst_w_mem_13__19_), .Y(w_mem_inst__abc_21203_new_n2579_));
OR2X2 OR2X2_2302 ( .A(w_mem_inst_w_mem_2__19_), .B(w_mem_inst_w_mem_0__19_), .Y(w_mem_inst__abc_21203_new_n2582_));
OR2X2 OR2X2_2303 ( .A(w_mem_inst__abc_21203_new_n2581_), .B(w_mem_inst__abc_21203_new_n2585_), .Y(w_mem_inst__abc_21203_new_n2586_));
OR2X2 OR2X2_2304 ( .A(w_mem_inst__abc_21203_new_n2587_), .B(w_mem_inst__abc_21203_new_n2580_), .Y(w_mem_inst__abc_21203_new_n2588_));
OR2X2 OR2X2_2305 ( .A(w_mem_inst__abc_21203_new_n2589_), .B(w_mem_inst__abc_21203_new_n1587_), .Y(w_mem_inst__abc_21203_new_n2590_));
OR2X2 OR2X2_2306 ( .A(w_mem_inst__abc_21203_new_n2591_), .B(w_mem_inst__abc_21203_new_n1586_), .Y(w_mem_inst__abc_21203_new_n2592_));
OR2X2 OR2X2_2307 ( .A(w_mem_inst__abc_21203_new_n2593_), .B(w_mem_inst__abc_21203_new_n2594_), .Y(w_mem_inst__abc_21203_new_n2595_));
OR2X2 OR2X2_2308 ( .A(w_mem_inst__abc_21203_new_n2595_), .B(w_mem_inst__abc_21203_new_n2592_), .Y(w_mem_inst__abc_21203_new_n2596_));
OR2X2 OR2X2_2309 ( .A(w_mem_inst__abc_21203_new_n2597_), .B(w_mem_inst__abc_21203_new_n2598_), .Y(w_mem_inst__abc_21203_new_n2599_));
OR2X2 OR2X2_231 ( .A(_abc_15497_new_n1432_), .B(_abc_15497_new_n1418_), .Y(_0H4_reg_31_0__26_));
OR2X2 OR2X2_2310 ( .A(w_mem_inst__abc_21203_new_n2596_), .B(w_mem_inst__abc_21203_new_n2599_), .Y(w_mem_inst__abc_21203_new_n2600_));
OR2X2 OR2X2_2311 ( .A(w_mem_inst__abc_21203_new_n2602_), .B(w_mem_inst__abc_21203_new_n2603_), .Y(w_mem_inst__abc_21203_new_n2604_));
OR2X2 OR2X2_2312 ( .A(w_mem_inst__abc_21203_new_n2604_), .B(w_mem_inst__abc_21203_new_n2601_), .Y(w_mem_inst__abc_21203_new_n2605_));
OR2X2 OR2X2_2313 ( .A(w_mem_inst__abc_21203_new_n2606_), .B(w_mem_inst__abc_21203_new_n2607_), .Y(w_mem_inst__abc_21203_new_n2608_));
OR2X2 OR2X2_2314 ( .A(w_mem_inst__abc_21203_new_n2609_), .B(w_mem_inst__abc_21203_new_n2610_), .Y(w_mem_inst__abc_21203_new_n2611_));
OR2X2 OR2X2_2315 ( .A(w_mem_inst__abc_21203_new_n2608_), .B(w_mem_inst__abc_21203_new_n2611_), .Y(w_mem_inst__abc_21203_new_n2612_));
OR2X2 OR2X2_2316 ( .A(w_mem_inst__abc_21203_new_n2613_), .B(w_mem_inst__abc_21203_new_n2614_), .Y(w_mem_inst__abc_21203_new_n2615_));
OR2X2 OR2X2_2317 ( .A(w_mem_inst__abc_21203_new_n2616_), .B(w_mem_inst__abc_21203_new_n2617_), .Y(w_mem_inst__abc_21203_new_n2618_));
OR2X2 OR2X2_2318 ( .A(w_mem_inst__abc_21203_new_n2615_), .B(w_mem_inst__abc_21203_new_n2618_), .Y(w_mem_inst__abc_21203_new_n2619_));
OR2X2 OR2X2_2319 ( .A(w_mem_inst__abc_21203_new_n2612_), .B(w_mem_inst__abc_21203_new_n2619_), .Y(w_mem_inst__abc_21203_new_n2620_));
OR2X2 OR2X2_232 ( .A(e_reg_27_), .B(\digest[27] ), .Y(_abc_15497_new_n1435_));
OR2X2 OR2X2_2320 ( .A(w_mem_inst__abc_21203_new_n2620_), .B(w_mem_inst__abc_21203_new_n2605_), .Y(w_mem_inst__abc_21203_new_n2621_));
OR2X2 OR2X2_2321 ( .A(w_mem_inst__abc_21203_new_n2621_), .B(w_mem_inst__abc_21203_new_n2600_), .Y(w_mem_inst__abc_21203_new_n2622_));
OR2X2 OR2X2_2322 ( .A(w_mem_inst__abc_21203_new_n2624_), .B(w_mem_inst_w_mem_8__20_), .Y(w_mem_inst__abc_21203_new_n2625_));
OR2X2 OR2X2_2323 ( .A(w_mem_inst__abc_21203_new_n2626_), .B(w_mem_inst_w_mem_13__20_), .Y(w_mem_inst__abc_21203_new_n2627_));
OR2X2 OR2X2_2324 ( .A(w_mem_inst_w_mem_2__20_), .B(w_mem_inst_w_mem_0__20_), .Y(w_mem_inst__abc_21203_new_n2630_));
OR2X2 OR2X2_2325 ( .A(w_mem_inst__abc_21203_new_n2629_), .B(w_mem_inst__abc_21203_new_n2633_), .Y(w_mem_inst__abc_21203_new_n2634_));
OR2X2 OR2X2_2326 ( .A(w_mem_inst__abc_21203_new_n2635_), .B(w_mem_inst__abc_21203_new_n2628_), .Y(w_mem_inst__abc_21203_new_n2636_));
OR2X2 OR2X2_2327 ( .A(w_mem_inst__abc_21203_new_n2637_), .B(w_mem_inst__abc_21203_new_n1587_), .Y(w_mem_inst__abc_21203_new_n2638_));
OR2X2 OR2X2_2328 ( .A(w_mem_inst__abc_21203_new_n2639_), .B(w_mem_inst__abc_21203_new_n1586_), .Y(w_mem_inst__abc_21203_new_n2640_));
OR2X2 OR2X2_2329 ( .A(w_mem_inst__abc_21203_new_n2641_), .B(w_mem_inst__abc_21203_new_n2642_), .Y(w_mem_inst__abc_21203_new_n2643_));
OR2X2 OR2X2_233 ( .A(_abc_15497_new_n1438_), .B(_abc_15497_new_n1425_), .Y(_abc_15497_new_n1439_));
OR2X2 OR2X2_2330 ( .A(w_mem_inst__abc_21203_new_n2643_), .B(w_mem_inst__abc_21203_new_n2640_), .Y(w_mem_inst__abc_21203_new_n2644_));
OR2X2 OR2X2_2331 ( .A(w_mem_inst__abc_21203_new_n2645_), .B(w_mem_inst__abc_21203_new_n2646_), .Y(w_mem_inst__abc_21203_new_n2647_));
OR2X2 OR2X2_2332 ( .A(w_mem_inst__abc_21203_new_n2644_), .B(w_mem_inst__abc_21203_new_n2647_), .Y(w_mem_inst__abc_21203_new_n2648_));
OR2X2 OR2X2_2333 ( .A(w_mem_inst__abc_21203_new_n2650_), .B(w_mem_inst__abc_21203_new_n2651_), .Y(w_mem_inst__abc_21203_new_n2652_));
OR2X2 OR2X2_2334 ( .A(w_mem_inst__abc_21203_new_n2652_), .B(w_mem_inst__abc_21203_new_n2649_), .Y(w_mem_inst__abc_21203_new_n2653_));
OR2X2 OR2X2_2335 ( .A(w_mem_inst__abc_21203_new_n2654_), .B(w_mem_inst__abc_21203_new_n2655_), .Y(w_mem_inst__abc_21203_new_n2656_));
OR2X2 OR2X2_2336 ( .A(w_mem_inst__abc_21203_new_n2657_), .B(w_mem_inst__abc_21203_new_n2658_), .Y(w_mem_inst__abc_21203_new_n2659_));
OR2X2 OR2X2_2337 ( .A(w_mem_inst__abc_21203_new_n2656_), .B(w_mem_inst__abc_21203_new_n2659_), .Y(w_mem_inst__abc_21203_new_n2660_));
OR2X2 OR2X2_2338 ( .A(w_mem_inst__abc_21203_new_n2661_), .B(w_mem_inst__abc_21203_new_n2662_), .Y(w_mem_inst__abc_21203_new_n2663_));
OR2X2 OR2X2_2339 ( .A(w_mem_inst__abc_21203_new_n2664_), .B(w_mem_inst__abc_21203_new_n2665_), .Y(w_mem_inst__abc_21203_new_n2666_));
OR2X2 OR2X2_234 ( .A(_abc_15497_new_n1429_), .B(_abc_15497_new_n1439_), .Y(_abc_15497_new_n1440_));
OR2X2 OR2X2_2340 ( .A(w_mem_inst__abc_21203_new_n2663_), .B(w_mem_inst__abc_21203_new_n2666_), .Y(w_mem_inst__abc_21203_new_n2667_));
OR2X2 OR2X2_2341 ( .A(w_mem_inst__abc_21203_new_n2660_), .B(w_mem_inst__abc_21203_new_n2667_), .Y(w_mem_inst__abc_21203_new_n2668_));
OR2X2 OR2X2_2342 ( .A(w_mem_inst__abc_21203_new_n2668_), .B(w_mem_inst__abc_21203_new_n2653_), .Y(w_mem_inst__abc_21203_new_n2669_));
OR2X2 OR2X2_2343 ( .A(w_mem_inst__abc_21203_new_n2669_), .B(w_mem_inst__abc_21203_new_n2648_), .Y(w_mem_inst__abc_21203_new_n2670_));
OR2X2 OR2X2_2344 ( .A(w_mem_inst__abc_21203_new_n2672_), .B(w_mem_inst_w_mem_8__21_), .Y(w_mem_inst__abc_21203_new_n2673_));
OR2X2 OR2X2_2345 ( .A(w_mem_inst__abc_21203_new_n2674_), .B(w_mem_inst_w_mem_13__21_), .Y(w_mem_inst__abc_21203_new_n2675_));
OR2X2 OR2X2_2346 ( .A(w_mem_inst_w_mem_2__21_), .B(w_mem_inst_w_mem_0__21_), .Y(w_mem_inst__abc_21203_new_n2678_));
OR2X2 OR2X2_2347 ( .A(w_mem_inst__abc_21203_new_n2677_), .B(w_mem_inst__abc_21203_new_n2681_), .Y(w_mem_inst__abc_21203_new_n2682_));
OR2X2 OR2X2_2348 ( .A(w_mem_inst__abc_21203_new_n2683_), .B(w_mem_inst__abc_21203_new_n2676_), .Y(w_mem_inst__abc_21203_new_n2684_));
OR2X2 OR2X2_2349 ( .A(w_mem_inst__abc_21203_new_n2685_), .B(w_mem_inst__abc_21203_new_n1587_), .Y(w_mem_inst__abc_21203_new_n2686_));
OR2X2 OR2X2_235 ( .A(_abc_15497_new_n1105_), .B(_abc_15497_new_n1443_), .Y(_abc_15497_new_n1444_));
OR2X2 OR2X2_2350 ( .A(w_mem_inst__abc_21203_new_n2687_), .B(w_mem_inst__abc_21203_new_n1586_), .Y(w_mem_inst__abc_21203_new_n2688_));
OR2X2 OR2X2_2351 ( .A(w_mem_inst__abc_21203_new_n2689_), .B(w_mem_inst__abc_21203_new_n2690_), .Y(w_mem_inst__abc_21203_new_n2691_));
OR2X2 OR2X2_2352 ( .A(w_mem_inst__abc_21203_new_n2691_), .B(w_mem_inst__abc_21203_new_n2688_), .Y(w_mem_inst__abc_21203_new_n2692_));
OR2X2 OR2X2_2353 ( .A(w_mem_inst__abc_21203_new_n2693_), .B(w_mem_inst__abc_21203_new_n2694_), .Y(w_mem_inst__abc_21203_new_n2695_));
OR2X2 OR2X2_2354 ( .A(w_mem_inst__abc_21203_new_n2692_), .B(w_mem_inst__abc_21203_new_n2695_), .Y(w_mem_inst__abc_21203_new_n2696_));
OR2X2 OR2X2_2355 ( .A(w_mem_inst__abc_21203_new_n2698_), .B(w_mem_inst__abc_21203_new_n2699_), .Y(w_mem_inst__abc_21203_new_n2700_));
OR2X2 OR2X2_2356 ( .A(w_mem_inst__abc_21203_new_n2700_), .B(w_mem_inst__abc_21203_new_n2697_), .Y(w_mem_inst__abc_21203_new_n2701_));
OR2X2 OR2X2_2357 ( .A(w_mem_inst__abc_21203_new_n2702_), .B(w_mem_inst__abc_21203_new_n2703_), .Y(w_mem_inst__abc_21203_new_n2704_));
OR2X2 OR2X2_2358 ( .A(w_mem_inst__abc_21203_new_n2705_), .B(w_mem_inst__abc_21203_new_n2706_), .Y(w_mem_inst__abc_21203_new_n2707_));
OR2X2 OR2X2_2359 ( .A(w_mem_inst__abc_21203_new_n2704_), .B(w_mem_inst__abc_21203_new_n2707_), .Y(w_mem_inst__abc_21203_new_n2708_));
OR2X2 OR2X2_236 ( .A(_abc_15497_new_n1445_), .B(_abc_15497_new_n1446_), .Y(_abc_15497_new_n1447_));
OR2X2 OR2X2_2360 ( .A(w_mem_inst__abc_21203_new_n2709_), .B(w_mem_inst__abc_21203_new_n2710_), .Y(w_mem_inst__abc_21203_new_n2711_));
OR2X2 OR2X2_2361 ( .A(w_mem_inst__abc_21203_new_n2712_), .B(w_mem_inst__abc_21203_new_n2713_), .Y(w_mem_inst__abc_21203_new_n2714_));
OR2X2 OR2X2_2362 ( .A(w_mem_inst__abc_21203_new_n2711_), .B(w_mem_inst__abc_21203_new_n2714_), .Y(w_mem_inst__abc_21203_new_n2715_));
OR2X2 OR2X2_2363 ( .A(w_mem_inst__abc_21203_new_n2708_), .B(w_mem_inst__abc_21203_new_n2715_), .Y(w_mem_inst__abc_21203_new_n2716_));
OR2X2 OR2X2_2364 ( .A(w_mem_inst__abc_21203_new_n2716_), .B(w_mem_inst__abc_21203_new_n2701_), .Y(w_mem_inst__abc_21203_new_n2717_));
OR2X2 OR2X2_2365 ( .A(w_mem_inst__abc_21203_new_n2717_), .B(w_mem_inst__abc_21203_new_n2696_), .Y(w_mem_inst__abc_21203_new_n2718_));
OR2X2 OR2X2_2366 ( .A(w_mem_inst__abc_21203_new_n2720_), .B(w_mem_inst_w_mem_8__22_), .Y(w_mem_inst__abc_21203_new_n2721_));
OR2X2 OR2X2_2367 ( .A(w_mem_inst__abc_21203_new_n2722_), .B(w_mem_inst_w_mem_13__22_), .Y(w_mem_inst__abc_21203_new_n2723_));
OR2X2 OR2X2_2368 ( .A(w_mem_inst_w_mem_2__22_), .B(w_mem_inst_w_mem_0__22_), .Y(w_mem_inst__abc_21203_new_n2726_));
OR2X2 OR2X2_2369 ( .A(w_mem_inst__abc_21203_new_n2725_), .B(w_mem_inst__abc_21203_new_n2729_), .Y(w_mem_inst__abc_21203_new_n2730_));
OR2X2 OR2X2_237 ( .A(_abc_15497_new_n1448_), .B(_abc_15497_new_n1449_), .Y(_abc_15497_new_n1450_));
OR2X2 OR2X2_2370 ( .A(w_mem_inst__abc_21203_new_n2731_), .B(w_mem_inst__abc_21203_new_n2724_), .Y(w_mem_inst__abc_21203_new_n2732_));
OR2X2 OR2X2_2371 ( .A(w_mem_inst__abc_21203_new_n2733_), .B(w_mem_inst__abc_21203_new_n1587_), .Y(w_mem_inst__abc_21203_new_n2734_));
OR2X2 OR2X2_2372 ( .A(w_mem_inst__abc_21203_new_n2735_), .B(w_mem_inst__abc_21203_new_n1586_), .Y(w_mem_inst__abc_21203_new_n2736_));
OR2X2 OR2X2_2373 ( .A(w_mem_inst__abc_21203_new_n2737_), .B(w_mem_inst__abc_21203_new_n2738_), .Y(w_mem_inst__abc_21203_new_n2739_));
OR2X2 OR2X2_2374 ( .A(w_mem_inst__abc_21203_new_n2739_), .B(w_mem_inst__abc_21203_new_n2736_), .Y(w_mem_inst__abc_21203_new_n2740_));
OR2X2 OR2X2_2375 ( .A(w_mem_inst__abc_21203_new_n2741_), .B(w_mem_inst__abc_21203_new_n2742_), .Y(w_mem_inst__abc_21203_new_n2743_));
OR2X2 OR2X2_2376 ( .A(w_mem_inst__abc_21203_new_n2740_), .B(w_mem_inst__abc_21203_new_n2743_), .Y(w_mem_inst__abc_21203_new_n2744_));
OR2X2 OR2X2_2377 ( .A(w_mem_inst__abc_21203_new_n2746_), .B(w_mem_inst__abc_21203_new_n2747_), .Y(w_mem_inst__abc_21203_new_n2748_));
OR2X2 OR2X2_2378 ( .A(w_mem_inst__abc_21203_new_n2748_), .B(w_mem_inst__abc_21203_new_n2745_), .Y(w_mem_inst__abc_21203_new_n2749_));
OR2X2 OR2X2_2379 ( .A(w_mem_inst__abc_21203_new_n2750_), .B(w_mem_inst__abc_21203_new_n2751_), .Y(w_mem_inst__abc_21203_new_n2752_));
OR2X2 OR2X2_238 ( .A(_abc_15497_new_n1451_), .B(_abc_15497_new_n1452_), .Y(_abc_15497_new_n1453_));
OR2X2 OR2X2_2380 ( .A(w_mem_inst__abc_21203_new_n2753_), .B(w_mem_inst__abc_21203_new_n2754_), .Y(w_mem_inst__abc_21203_new_n2755_));
OR2X2 OR2X2_2381 ( .A(w_mem_inst__abc_21203_new_n2752_), .B(w_mem_inst__abc_21203_new_n2755_), .Y(w_mem_inst__abc_21203_new_n2756_));
OR2X2 OR2X2_2382 ( .A(w_mem_inst__abc_21203_new_n2757_), .B(w_mem_inst__abc_21203_new_n2758_), .Y(w_mem_inst__abc_21203_new_n2759_));
OR2X2 OR2X2_2383 ( .A(w_mem_inst__abc_21203_new_n2760_), .B(w_mem_inst__abc_21203_new_n2761_), .Y(w_mem_inst__abc_21203_new_n2762_));
OR2X2 OR2X2_2384 ( .A(w_mem_inst__abc_21203_new_n2759_), .B(w_mem_inst__abc_21203_new_n2762_), .Y(w_mem_inst__abc_21203_new_n2763_));
OR2X2 OR2X2_2385 ( .A(w_mem_inst__abc_21203_new_n2756_), .B(w_mem_inst__abc_21203_new_n2763_), .Y(w_mem_inst__abc_21203_new_n2764_));
OR2X2 OR2X2_2386 ( .A(w_mem_inst__abc_21203_new_n2764_), .B(w_mem_inst__abc_21203_new_n2749_), .Y(w_mem_inst__abc_21203_new_n2765_));
OR2X2 OR2X2_2387 ( .A(w_mem_inst__abc_21203_new_n2765_), .B(w_mem_inst__abc_21203_new_n2744_), .Y(w_mem_inst__abc_21203_new_n2766_));
OR2X2 OR2X2_2388 ( .A(w_mem_inst__abc_21203_new_n2768_), .B(w_mem_inst_w_mem_8__23_), .Y(w_mem_inst__abc_21203_new_n2769_));
OR2X2 OR2X2_2389 ( .A(w_mem_inst__abc_21203_new_n2770_), .B(w_mem_inst_w_mem_13__23_), .Y(w_mem_inst__abc_21203_new_n2771_));
OR2X2 OR2X2_239 ( .A(_abc_15497_new_n1455_), .B(_abc_15497_new_n1457_), .Y(_abc_15497_new_n1458_));
OR2X2 OR2X2_2390 ( .A(w_mem_inst_w_mem_2__23_), .B(w_mem_inst_w_mem_0__23_), .Y(w_mem_inst__abc_21203_new_n2774_));
OR2X2 OR2X2_2391 ( .A(w_mem_inst__abc_21203_new_n2773_), .B(w_mem_inst__abc_21203_new_n2777_), .Y(w_mem_inst__abc_21203_new_n2778_));
OR2X2 OR2X2_2392 ( .A(w_mem_inst__abc_21203_new_n2779_), .B(w_mem_inst__abc_21203_new_n2772_), .Y(w_mem_inst__abc_21203_new_n2780_));
OR2X2 OR2X2_2393 ( .A(w_mem_inst__abc_21203_new_n2781_), .B(w_mem_inst__abc_21203_new_n1587_), .Y(w_mem_inst__abc_21203_new_n2782_));
OR2X2 OR2X2_2394 ( .A(w_mem_inst__abc_21203_new_n2783_), .B(w_mem_inst__abc_21203_new_n1586_), .Y(w_mem_inst__abc_21203_new_n2784_));
OR2X2 OR2X2_2395 ( .A(w_mem_inst__abc_21203_new_n2785_), .B(w_mem_inst__abc_21203_new_n2786_), .Y(w_mem_inst__abc_21203_new_n2787_));
OR2X2 OR2X2_2396 ( .A(w_mem_inst__abc_21203_new_n2787_), .B(w_mem_inst__abc_21203_new_n2784_), .Y(w_mem_inst__abc_21203_new_n2788_));
OR2X2 OR2X2_2397 ( .A(w_mem_inst__abc_21203_new_n2789_), .B(w_mem_inst__abc_21203_new_n2790_), .Y(w_mem_inst__abc_21203_new_n2791_));
OR2X2 OR2X2_2398 ( .A(w_mem_inst__abc_21203_new_n2788_), .B(w_mem_inst__abc_21203_new_n2791_), .Y(w_mem_inst__abc_21203_new_n2792_));
OR2X2 OR2X2_2399 ( .A(w_mem_inst__abc_21203_new_n2794_), .B(w_mem_inst__abc_21203_new_n2795_), .Y(w_mem_inst__abc_21203_new_n2796_));
OR2X2 OR2X2_24 ( .A(c_reg_9_), .B(\digest[73] ), .Y(_abc_15497_new_n797_));
OR2X2 OR2X2_240 ( .A(_abc_15497_new_n1463_), .B(_abc_15497_new_n1434_), .Y(_0H4_reg_31_0__27_));
OR2X2 OR2X2_2400 ( .A(w_mem_inst__abc_21203_new_n2796_), .B(w_mem_inst__abc_21203_new_n2793_), .Y(w_mem_inst__abc_21203_new_n2797_));
OR2X2 OR2X2_2401 ( .A(w_mem_inst__abc_21203_new_n2798_), .B(w_mem_inst__abc_21203_new_n2799_), .Y(w_mem_inst__abc_21203_new_n2800_));
OR2X2 OR2X2_2402 ( .A(w_mem_inst__abc_21203_new_n2801_), .B(w_mem_inst__abc_21203_new_n2802_), .Y(w_mem_inst__abc_21203_new_n2803_));
OR2X2 OR2X2_2403 ( .A(w_mem_inst__abc_21203_new_n2800_), .B(w_mem_inst__abc_21203_new_n2803_), .Y(w_mem_inst__abc_21203_new_n2804_));
OR2X2 OR2X2_2404 ( .A(w_mem_inst__abc_21203_new_n2805_), .B(w_mem_inst__abc_21203_new_n2806_), .Y(w_mem_inst__abc_21203_new_n2807_));
OR2X2 OR2X2_2405 ( .A(w_mem_inst__abc_21203_new_n2808_), .B(w_mem_inst__abc_21203_new_n2809_), .Y(w_mem_inst__abc_21203_new_n2810_));
OR2X2 OR2X2_2406 ( .A(w_mem_inst__abc_21203_new_n2807_), .B(w_mem_inst__abc_21203_new_n2810_), .Y(w_mem_inst__abc_21203_new_n2811_));
OR2X2 OR2X2_2407 ( .A(w_mem_inst__abc_21203_new_n2804_), .B(w_mem_inst__abc_21203_new_n2811_), .Y(w_mem_inst__abc_21203_new_n2812_));
OR2X2 OR2X2_2408 ( .A(w_mem_inst__abc_21203_new_n2812_), .B(w_mem_inst__abc_21203_new_n2797_), .Y(w_mem_inst__abc_21203_new_n2813_));
OR2X2 OR2X2_2409 ( .A(w_mem_inst__abc_21203_new_n2813_), .B(w_mem_inst__abc_21203_new_n2792_), .Y(w_mem_inst__abc_21203_new_n2814_));
OR2X2 OR2X2_241 ( .A(_abc_15497_new_n1466_), .B(_abc_15497_new_n1468_), .Y(_abc_15497_new_n1469_));
OR2X2 OR2X2_2410 ( .A(w_mem_inst__abc_21203_new_n2816_), .B(w_mem_inst_w_mem_8__24_), .Y(w_mem_inst__abc_21203_new_n2817_));
OR2X2 OR2X2_2411 ( .A(w_mem_inst__abc_21203_new_n2818_), .B(w_mem_inst_w_mem_13__24_), .Y(w_mem_inst__abc_21203_new_n2819_));
OR2X2 OR2X2_2412 ( .A(w_mem_inst_w_mem_2__24_), .B(w_mem_inst_w_mem_0__24_), .Y(w_mem_inst__abc_21203_new_n2822_));
OR2X2 OR2X2_2413 ( .A(w_mem_inst__abc_21203_new_n2821_), .B(w_mem_inst__abc_21203_new_n2825_), .Y(w_mem_inst__abc_21203_new_n2826_));
OR2X2 OR2X2_2414 ( .A(w_mem_inst__abc_21203_new_n2827_), .B(w_mem_inst__abc_21203_new_n2820_), .Y(w_mem_inst__abc_21203_new_n2828_));
OR2X2 OR2X2_2415 ( .A(w_mem_inst__abc_21203_new_n2829_), .B(w_mem_inst__abc_21203_new_n1587_), .Y(w_mem_inst__abc_21203_new_n2830_));
OR2X2 OR2X2_2416 ( .A(w_mem_inst__abc_21203_new_n2831_), .B(w_mem_inst__abc_21203_new_n1586_), .Y(w_mem_inst__abc_21203_new_n2832_));
OR2X2 OR2X2_2417 ( .A(w_mem_inst__abc_21203_new_n2833_), .B(w_mem_inst__abc_21203_new_n2834_), .Y(w_mem_inst__abc_21203_new_n2835_));
OR2X2 OR2X2_2418 ( .A(w_mem_inst__abc_21203_new_n2835_), .B(w_mem_inst__abc_21203_new_n2832_), .Y(w_mem_inst__abc_21203_new_n2836_));
OR2X2 OR2X2_2419 ( .A(w_mem_inst__abc_21203_new_n2837_), .B(w_mem_inst__abc_21203_new_n2838_), .Y(w_mem_inst__abc_21203_new_n2839_));
OR2X2 OR2X2_242 ( .A(e_reg_28_), .B(\digest[28] ), .Y(_abc_15497_new_n1470_));
OR2X2 OR2X2_2420 ( .A(w_mem_inst__abc_21203_new_n2836_), .B(w_mem_inst__abc_21203_new_n2839_), .Y(w_mem_inst__abc_21203_new_n2840_));
OR2X2 OR2X2_2421 ( .A(w_mem_inst__abc_21203_new_n2842_), .B(w_mem_inst__abc_21203_new_n2843_), .Y(w_mem_inst__abc_21203_new_n2844_));
OR2X2 OR2X2_2422 ( .A(w_mem_inst__abc_21203_new_n2844_), .B(w_mem_inst__abc_21203_new_n2841_), .Y(w_mem_inst__abc_21203_new_n2845_));
OR2X2 OR2X2_2423 ( .A(w_mem_inst__abc_21203_new_n2846_), .B(w_mem_inst__abc_21203_new_n2847_), .Y(w_mem_inst__abc_21203_new_n2848_));
OR2X2 OR2X2_2424 ( .A(w_mem_inst__abc_21203_new_n2849_), .B(w_mem_inst__abc_21203_new_n2850_), .Y(w_mem_inst__abc_21203_new_n2851_));
OR2X2 OR2X2_2425 ( .A(w_mem_inst__abc_21203_new_n2848_), .B(w_mem_inst__abc_21203_new_n2851_), .Y(w_mem_inst__abc_21203_new_n2852_));
OR2X2 OR2X2_2426 ( .A(w_mem_inst__abc_21203_new_n2853_), .B(w_mem_inst__abc_21203_new_n2854_), .Y(w_mem_inst__abc_21203_new_n2855_));
OR2X2 OR2X2_2427 ( .A(w_mem_inst__abc_21203_new_n2856_), .B(w_mem_inst__abc_21203_new_n2857_), .Y(w_mem_inst__abc_21203_new_n2858_));
OR2X2 OR2X2_2428 ( .A(w_mem_inst__abc_21203_new_n2855_), .B(w_mem_inst__abc_21203_new_n2858_), .Y(w_mem_inst__abc_21203_new_n2859_));
OR2X2 OR2X2_2429 ( .A(w_mem_inst__abc_21203_new_n2852_), .B(w_mem_inst__abc_21203_new_n2859_), .Y(w_mem_inst__abc_21203_new_n2860_));
OR2X2 OR2X2_243 ( .A(_abc_15497_new_n1469_), .B(_abc_15497_new_n1473_), .Y(_abc_15497_new_n1474_));
OR2X2 OR2X2_2430 ( .A(w_mem_inst__abc_21203_new_n2860_), .B(w_mem_inst__abc_21203_new_n2845_), .Y(w_mem_inst__abc_21203_new_n2861_));
OR2X2 OR2X2_2431 ( .A(w_mem_inst__abc_21203_new_n2861_), .B(w_mem_inst__abc_21203_new_n2840_), .Y(w_mem_inst__abc_21203_new_n2862_));
OR2X2 OR2X2_2432 ( .A(w_mem_inst__abc_21203_new_n2864_), .B(w_mem_inst_w_mem_8__25_), .Y(w_mem_inst__abc_21203_new_n2865_));
OR2X2 OR2X2_2433 ( .A(w_mem_inst__abc_21203_new_n2866_), .B(w_mem_inst_w_mem_13__25_), .Y(w_mem_inst__abc_21203_new_n2867_));
OR2X2 OR2X2_2434 ( .A(w_mem_inst_w_mem_2__25_), .B(w_mem_inst_w_mem_0__25_), .Y(w_mem_inst__abc_21203_new_n2870_));
OR2X2 OR2X2_2435 ( .A(w_mem_inst__abc_21203_new_n2869_), .B(w_mem_inst__abc_21203_new_n2873_), .Y(w_mem_inst__abc_21203_new_n2874_));
OR2X2 OR2X2_2436 ( .A(w_mem_inst__abc_21203_new_n2875_), .B(w_mem_inst__abc_21203_new_n2868_), .Y(w_mem_inst__abc_21203_new_n2876_));
OR2X2 OR2X2_2437 ( .A(w_mem_inst__abc_21203_new_n2877_), .B(w_mem_inst__abc_21203_new_n1587_), .Y(w_mem_inst__abc_21203_new_n2878_));
OR2X2 OR2X2_2438 ( .A(w_mem_inst__abc_21203_new_n2879_), .B(w_mem_inst__abc_21203_new_n1586_), .Y(w_mem_inst__abc_21203_new_n2880_));
OR2X2 OR2X2_2439 ( .A(w_mem_inst__abc_21203_new_n2881_), .B(w_mem_inst__abc_21203_new_n2882_), .Y(w_mem_inst__abc_21203_new_n2883_));
OR2X2 OR2X2_244 ( .A(_abc_15497_new_n1475_), .B(_abc_15497_new_n1476_), .Y(_abc_15497_new_n1477_));
OR2X2 OR2X2_2440 ( .A(w_mem_inst__abc_21203_new_n2883_), .B(w_mem_inst__abc_21203_new_n2880_), .Y(w_mem_inst__abc_21203_new_n2884_));
OR2X2 OR2X2_2441 ( .A(w_mem_inst__abc_21203_new_n2885_), .B(w_mem_inst__abc_21203_new_n2886_), .Y(w_mem_inst__abc_21203_new_n2887_));
OR2X2 OR2X2_2442 ( .A(w_mem_inst__abc_21203_new_n2884_), .B(w_mem_inst__abc_21203_new_n2887_), .Y(w_mem_inst__abc_21203_new_n2888_));
OR2X2 OR2X2_2443 ( .A(w_mem_inst__abc_21203_new_n2890_), .B(w_mem_inst__abc_21203_new_n2891_), .Y(w_mem_inst__abc_21203_new_n2892_));
OR2X2 OR2X2_2444 ( .A(w_mem_inst__abc_21203_new_n2892_), .B(w_mem_inst__abc_21203_new_n2889_), .Y(w_mem_inst__abc_21203_new_n2893_));
OR2X2 OR2X2_2445 ( .A(w_mem_inst__abc_21203_new_n2894_), .B(w_mem_inst__abc_21203_new_n2895_), .Y(w_mem_inst__abc_21203_new_n2896_));
OR2X2 OR2X2_2446 ( .A(w_mem_inst__abc_21203_new_n2897_), .B(w_mem_inst__abc_21203_new_n2898_), .Y(w_mem_inst__abc_21203_new_n2899_));
OR2X2 OR2X2_2447 ( .A(w_mem_inst__abc_21203_new_n2896_), .B(w_mem_inst__abc_21203_new_n2899_), .Y(w_mem_inst__abc_21203_new_n2900_));
OR2X2 OR2X2_2448 ( .A(w_mem_inst__abc_21203_new_n2901_), .B(w_mem_inst__abc_21203_new_n2902_), .Y(w_mem_inst__abc_21203_new_n2903_));
OR2X2 OR2X2_2449 ( .A(w_mem_inst__abc_21203_new_n2904_), .B(w_mem_inst__abc_21203_new_n2905_), .Y(w_mem_inst__abc_21203_new_n2906_));
OR2X2 OR2X2_245 ( .A(_abc_15497_new_n1479_), .B(_abc_15497_new_n1465_), .Y(_0H4_reg_31_0__28_));
OR2X2 OR2X2_2450 ( .A(w_mem_inst__abc_21203_new_n2903_), .B(w_mem_inst__abc_21203_new_n2906_), .Y(w_mem_inst__abc_21203_new_n2907_));
OR2X2 OR2X2_2451 ( .A(w_mem_inst__abc_21203_new_n2900_), .B(w_mem_inst__abc_21203_new_n2907_), .Y(w_mem_inst__abc_21203_new_n2908_));
OR2X2 OR2X2_2452 ( .A(w_mem_inst__abc_21203_new_n2908_), .B(w_mem_inst__abc_21203_new_n2893_), .Y(w_mem_inst__abc_21203_new_n2909_));
OR2X2 OR2X2_2453 ( .A(w_mem_inst__abc_21203_new_n2909_), .B(w_mem_inst__abc_21203_new_n2888_), .Y(w_mem_inst__abc_21203_new_n2910_));
OR2X2 OR2X2_2454 ( .A(w_mem_inst__abc_21203_new_n2912_), .B(w_mem_inst_w_mem_8__26_), .Y(w_mem_inst__abc_21203_new_n2913_));
OR2X2 OR2X2_2455 ( .A(w_mem_inst__abc_21203_new_n2914_), .B(w_mem_inst_w_mem_13__26_), .Y(w_mem_inst__abc_21203_new_n2915_));
OR2X2 OR2X2_2456 ( .A(w_mem_inst_w_mem_2__26_), .B(w_mem_inst_w_mem_0__26_), .Y(w_mem_inst__abc_21203_new_n2918_));
OR2X2 OR2X2_2457 ( .A(w_mem_inst__abc_21203_new_n2917_), .B(w_mem_inst__abc_21203_new_n2921_), .Y(w_mem_inst__abc_21203_new_n2922_));
OR2X2 OR2X2_2458 ( .A(w_mem_inst__abc_21203_new_n2923_), .B(w_mem_inst__abc_21203_new_n2916_), .Y(w_mem_inst__abc_21203_new_n2924_));
OR2X2 OR2X2_2459 ( .A(w_mem_inst__abc_21203_new_n2925_), .B(w_mem_inst__abc_21203_new_n1587_), .Y(w_mem_inst__abc_21203_new_n2926_));
OR2X2 OR2X2_246 ( .A(_abc_15497_new_n1481_), .B(digest_update), .Y(_abc_15497_new_n1482_));
OR2X2 OR2X2_2460 ( .A(w_mem_inst__abc_21203_new_n2927_), .B(w_mem_inst__abc_21203_new_n1586_), .Y(w_mem_inst__abc_21203_new_n2928_));
OR2X2 OR2X2_2461 ( .A(w_mem_inst__abc_21203_new_n2929_), .B(w_mem_inst__abc_21203_new_n2930_), .Y(w_mem_inst__abc_21203_new_n2931_));
OR2X2 OR2X2_2462 ( .A(w_mem_inst__abc_21203_new_n2931_), .B(w_mem_inst__abc_21203_new_n2928_), .Y(w_mem_inst__abc_21203_new_n2932_));
OR2X2 OR2X2_2463 ( .A(w_mem_inst__abc_21203_new_n2933_), .B(w_mem_inst__abc_21203_new_n2934_), .Y(w_mem_inst__abc_21203_new_n2935_));
OR2X2 OR2X2_2464 ( .A(w_mem_inst__abc_21203_new_n2932_), .B(w_mem_inst__abc_21203_new_n2935_), .Y(w_mem_inst__abc_21203_new_n2936_));
OR2X2 OR2X2_2465 ( .A(w_mem_inst__abc_21203_new_n2938_), .B(w_mem_inst__abc_21203_new_n2939_), .Y(w_mem_inst__abc_21203_new_n2940_));
OR2X2 OR2X2_2466 ( .A(w_mem_inst__abc_21203_new_n2940_), .B(w_mem_inst__abc_21203_new_n2937_), .Y(w_mem_inst__abc_21203_new_n2941_));
OR2X2 OR2X2_2467 ( .A(w_mem_inst__abc_21203_new_n2942_), .B(w_mem_inst__abc_21203_new_n2943_), .Y(w_mem_inst__abc_21203_new_n2944_));
OR2X2 OR2X2_2468 ( .A(w_mem_inst__abc_21203_new_n2945_), .B(w_mem_inst__abc_21203_new_n2946_), .Y(w_mem_inst__abc_21203_new_n2947_));
OR2X2 OR2X2_2469 ( .A(w_mem_inst__abc_21203_new_n2944_), .B(w_mem_inst__abc_21203_new_n2947_), .Y(w_mem_inst__abc_21203_new_n2948_));
OR2X2 OR2X2_247 ( .A(e_reg_29_), .B(\digest[29] ), .Y(_abc_15497_new_n1484_));
OR2X2 OR2X2_2470 ( .A(w_mem_inst__abc_21203_new_n2949_), .B(w_mem_inst__abc_21203_new_n2950_), .Y(w_mem_inst__abc_21203_new_n2951_));
OR2X2 OR2X2_2471 ( .A(w_mem_inst__abc_21203_new_n2952_), .B(w_mem_inst__abc_21203_new_n2953_), .Y(w_mem_inst__abc_21203_new_n2954_));
OR2X2 OR2X2_2472 ( .A(w_mem_inst__abc_21203_new_n2951_), .B(w_mem_inst__abc_21203_new_n2954_), .Y(w_mem_inst__abc_21203_new_n2955_));
OR2X2 OR2X2_2473 ( .A(w_mem_inst__abc_21203_new_n2948_), .B(w_mem_inst__abc_21203_new_n2955_), .Y(w_mem_inst__abc_21203_new_n2956_));
OR2X2 OR2X2_2474 ( .A(w_mem_inst__abc_21203_new_n2956_), .B(w_mem_inst__abc_21203_new_n2941_), .Y(w_mem_inst__abc_21203_new_n2957_));
OR2X2 OR2X2_2475 ( .A(w_mem_inst__abc_21203_new_n2957_), .B(w_mem_inst__abc_21203_new_n2936_), .Y(w_mem_inst__abc_21203_new_n2958_));
OR2X2 OR2X2_2476 ( .A(w_mem_inst__abc_21203_new_n2960_), .B(w_mem_inst_w_mem_8__27_), .Y(w_mem_inst__abc_21203_new_n2961_));
OR2X2 OR2X2_2477 ( .A(w_mem_inst__abc_21203_new_n2962_), .B(w_mem_inst_w_mem_13__27_), .Y(w_mem_inst__abc_21203_new_n2963_));
OR2X2 OR2X2_2478 ( .A(w_mem_inst_w_mem_2__27_), .B(w_mem_inst_w_mem_0__27_), .Y(w_mem_inst__abc_21203_new_n2966_));
OR2X2 OR2X2_2479 ( .A(w_mem_inst__abc_21203_new_n2965_), .B(w_mem_inst__abc_21203_new_n2969_), .Y(w_mem_inst__abc_21203_new_n2970_));
OR2X2 OR2X2_248 ( .A(_abc_15497_new_n1489_), .B(_abc_15497_new_n1471_), .Y(_abc_15497_new_n1490_));
OR2X2 OR2X2_2480 ( .A(w_mem_inst__abc_21203_new_n2971_), .B(w_mem_inst__abc_21203_new_n2964_), .Y(w_mem_inst__abc_21203_new_n2972_));
OR2X2 OR2X2_2481 ( .A(w_mem_inst__abc_21203_new_n2973_), .B(w_mem_inst__abc_21203_new_n1587_), .Y(w_mem_inst__abc_21203_new_n2974_));
OR2X2 OR2X2_2482 ( .A(w_mem_inst__abc_21203_new_n2975_), .B(w_mem_inst__abc_21203_new_n1586_), .Y(w_mem_inst__abc_21203_new_n2976_));
OR2X2 OR2X2_2483 ( .A(w_mem_inst__abc_21203_new_n2977_), .B(w_mem_inst__abc_21203_new_n2978_), .Y(w_mem_inst__abc_21203_new_n2979_));
OR2X2 OR2X2_2484 ( .A(w_mem_inst__abc_21203_new_n2979_), .B(w_mem_inst__abc_21203_new_n2976_), .Y(w_mem_inst__abc_21203_new_n2980_));
OR2X2 OR2X2_2485 ( .A(w_mem_inst__abc_21203_new_n2981_), .B(w_mem_inst__abc_21203_new_n2982_), .Y(w_mem_inst__abc_21203_new_n2983_));
OR2X2 OR2X2_2486 ( .A(w_mem_inst__abc_21203_new_n2980_), .B(w_mem_inst__abc_21203_new_n2983_), .Y(w_mem_inst__abc_21203_new_n2984_));
OR2X2 OR2X2_2487 ( .A(w_mem_inst__abc_21203_new_n2986_), .B(w_mem_inst__abc_21203_new_n2987_), .Y(w_mem_inst__abc_21203_new_n2988_));
OR2X2 OR2X2_2488 ( .A(w_mem_inst__abc_21203_new_n2988_), .B(w_mem_inst__abc_21203_new_n2985_), .Y(w_mem_inst__abc_21203_new_n2989_));
OR2X2 OR2X2_2489 ( .A(w_mem_inst__abc_21203_new_n2990_), .B(w_mem_inst__abc_21203_new_n2991_), .Y(w_mem_inst__abc_21203_new_n2992_));
OR2X2 OR2X2_249 ( .A(_abc_15497_new_n1492_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n1493_));
OR2X2 OR2X2_2490 ( .A(w_mem_inst__abc_21203_new_n2993_), .B(w_mem_inst__abc_21203_new_n2994_), .Y(w_mem_inst__abc_21203_new_n2995_));
OR2X2 OR2X2_2491 ( .A(w_mem_inst__abc_21203_new_n2992_), .B(w_mem_inst__abc_21203_new_n2995_), .Y(w_mem_inst__abc_21203_new_n2996_));
OR2X2 OR2X2_2492 ( .A(w_mem_inst__abc_21203_new_n2997_), .B(w_mem_inst__abc_21203_new_n2998_), .Y(w_mem_inst__abc_21203_new_n2999_));
OR2X2 OR2X2_2493 ( .A(w_mem_inst__abc_21203_new_n3000_), .B(w_mem_inst__abc_21203_new_n3001_), .Y(w_mem_inst__abc_21203_new_n3002_));
OR2X2 OR2X2_2494 ( .A(w_mem_inst__abc_21203_new_n2999_), .B(w_mem_inst__abc_21203_new_n3002_), .Y(w_mem_inst__abc_21203_new_n3003_));
OR2X2 OR2X2_2495 ( .A(w_mem_inst__abc_21203_new_n2996_), .B(w_mem_inst__abc_21203_new_n3003_), .Y(w_mem_inst__abc_21203_new_n3004_));
OR2X2 OR2X2_2496 ( .A(w_mem_inst__abc_21203_new_n3004_), .B(w_mem_inst__abc_21203_new_n2989_), .Y(w_mem_inst__abc_21203_new_n3005_));
OR2X2 OR2X2_2497 ( .A(w_mem_inst__abc_21203_new_n3005_), .B(w_mem_inst__abc_21203_new_n2984_), .Y(w_mem_inst__abc_21203_new_n3006_));
OR2X2 OR2X2_2498 ( .A(w_mem_inst__abc_21203_new_n3008_), .B(w_mem_inst_w_mem_8__28_), .Y(w_mem_inst__abc_21203_new_n3009_));
OR2X2 OR2X2_2499 ( .A(w_mem_inst__abc_21203_new_n3010_), .B(w_mem_inst_w_mem_13__28_), .Y(w_mem_inst__abc_21203_new_n3011_));
OR2X2 OR2X2_25 ( .A(_abc_15497_new_n799_), .B(_abc_15497_new_n796_), .Y(_abc_15497_new_n800_));
OR2X2 OR2X2_250 ( .A(_abc_15497_new_n1493_), .B(_abc_15497_new_n1488_), .Y(_abc_15497_new_n1494_));
OR2X2 OR2X2_2500 ( .A(w_mem_inst_w_mem_2__28_), .B(w_mem_inst_w_mem_0__28_), .Y(w_mem_inst__abc_21203_new_n3014_));
OR2X2 OR2X2_2501 ( .A(w_mem_inst__abc_21203_new_n3013_), .B(w_mem_inst__abc_21203_new_n3017_), .Y(w_mem_inst__abc_21203_new_n3018_));
OR2X2 OR2X2_2502 ( .A(w_mem_inst__abc_21203_new_n3019_), .B(w_mem_inst__abc_21203_new_n3012_), .Y(w_mem_inst__abc_21203_new_n3020_));
OR2X2 OR2X2_2503 ( .A(w_mem_inst__abc_21203_new_n3021_), .B(w_mem_inst__abc_21203_new_n1587_), .Y(w_mem_inst__abc_21203_new_n3022_));
OR2X2 OR2X2_2504 ( .A(w_mem_inst__abc_21203_new_n3023_), .B(w_mem_inst__abc_21203_new_n1586_), .Y(w_mem_inst__abc_21203_new_n3024_));
OR2X2 OR2X2_2505 ( .A(w_mem_inst__abc_21203_new_n3025_), .B(w_mem_inst__abc_21203_new_n3026_), .Y(w_mem_inst__abc_21203_new_n3027_));
OR2X2 OR2X2_2506 ( .A(w_mem_inst__abc_21203_new_n3027_), .B(w_mem_inst__abc_21203_new_n3024_), .Y(w_mem_inst__abc_21203_new_n3028_));
OR2X2 OR2X2_2507 ( .A(w_mem_inst__abc_21203_new_n3029_), .B(w_mem_inst__abc_21203_new_n3030_), .Y(w_mem_inst__abc_21203_new_n3031_));
OR2X2 OR2X2_2508 ( .A(w_mem_inst__abc_21203_new_n3028_), .B(w_mem_inst__abc_21203_new_n3031_), .Y(w_mem_inst__abc_21203_new_n3032_));
OR2X2 OR2X2_2509 ( .A(w_mem_inst__abc_21203_new_n3034_), .B(w_mem_inst__abc_21203_new_n3035_), .Y(w_mem_inst__abc_21203_new_n3036_));
OR2X2 OR2X2_251 ( .A(e_reg_30_), .B(\digest[30] ), .Y(_abc_15497_new_n1496_));
OR2X2 OR2X2_2510 ( .A(w_mem_inst__abc_21203_new_n3036_), .B(w_mem_inst__abc_21203_new_n3033_), .Y(w_mem_inst__abc_21203_new_n3037_));
OR2X2 OR2X2_2511 ( .A(w_mem_inst__abc_21203_new_n3038_), .B(w_mem_inst__abc_21203_new_n3039_), .Y(w_mem_inst__abc_21203_new_n3040_));
OR2X2 OR2X2_2512 ( .A(w_mem_inst__abc_21203_new_n3041_), .B(w_mem_inst__abc_21203_new_n3042_), .Y(w_mem_inst__abc_21203_new_n3043_));
OR2X2 OR2X2_2513 ( .A(w_mem_inst__abc_21203_new_n3040_), .B(w_mem_inst__abc_21203_new_n3043_), .Y(w_mem_inst__abc_21203_new_n3044_));
OR2X2 OR2X2_2514 ( .A(w_mem_inst__abc_21203_new_n3045_), .B(w_mem_inst__abc_21203_new_n3046_), .Y(w_mem_inst__abc_21203_new_n3047_));
OR2X2 OR2X2_2515 ( .A(w_mem_inst__abc_21203_new_n3048_), .B(w_mem_inst__abc_21203_new_n3049_), .Y(w_mem_inst__abc_21203_new_n3050_));
OR2X2 OR2X2_2516 ( .A(w_mem_inst__abc_21203_new_n3047_), .B(w_mem_inst__abc_21203_new_n3050_), .Y(w_mem_inst__abc_21203_new_n3051_));
OR2X2 OR2X2_2517 ( .A(w_mem_inst__abc_21203_new_n3044_), .B(w_mem_inst__abc_21203_new_n3051_), .Y(w_mem_inst__abc_21203_new_n3052_));
OR2X2 OR2X2_2518 ( .A(w_mem_inst__abc_21203_new_n3052_), .B(w_mem_inst__abc_21203_new_n3037_), .Y(w_mem_inst__abc_21203_new_n3053_));
OR2X2 OR2X2_2519 ( .A(w_mem_inst__abc_21203_new_n3053_), .B(w_mem_inst__abc_21203_new_n3032_), .Y(w_mem_inst__abc_21203_new_n3054_));
OR2X2 OR2X2_252 ( .A(_abc_15497_new_n1500_), .B(_abc_15497_new_n1485_), .Y(_abc_15497_new_n1501_));
OR2X2 OR2X2_2520 ( .A(w_mem_inst__abc_21203_new_n3056_), .B(w_mem_inst_w_mem_8__29_), .Y(w_mem_inst__abc_21203_new_n3057_));
OR2X2 OR2X2_2521 ( .A(w_mem_inst__abc_21203_new_n3058_), .B(w_mem_inst_w_mem_13__29_), .Y(w_mem_inst__abc_21203_new_n3059_));
OR2X2 OR2X2_2522 ( .A(w_mem_inst_w_mem_2__29_), .B(w_mem_inst_w_mem_0__29_), .Y(w_mem_inst__abc_21203_new_n3062_));
OR2X2 OR2X2_2523 ( .A(w_mem_inst__abc_21203_new_n3061_), .B(w_mem_inst__abc_21203_new_n3065_), .Y(w_mem_inst__abc_21203_new_n3066_));
OR2X2 OR2X2_2524 ( .A(w_mem_inst__abc_21203_new_n3067_), .B(w_mem_inst__abc_21203_new_n3060_), .Y(w_mem_inst__abc_21203_new_n3068_));
OR2X2 OR2X2_2525 ( .A(w_mem_inst__abc_21203_new_n3069_), .B(w_mem_inst__abc_21203_new_n1587_), .Y(w_mem_inst__abc_21203_new_n3070_));
OR2X2 OR2X2_2526 ( .A(w_mem_inst__abc_21203_new_n3071_), .B(w_mem_inst__abc_21203_new_n1586_), .Y(w_mem_inst__abc_21203_new_n3072_));
OR2X2 OR2X2_2527 ( .A(w_mem_inst__abc_21203_new_n3073_), .B(w_mem_inst__abc_21203_new_n3074_), .Y(w_mem_inst__abc_21203_new_n3075_));
OR2X2 OR2X2_2528 ( .A(w_mem_inst__abc_21203_new_n3075_), .B(w_mem_inst__abc_21203_new_n3072_), .Y(w_mem_inst__abc_21203_new_n3076_));
OR2X2 OR2X2_2529 ( .A(w_mem_inst__abc_21203_new_n3077_), .B(w_mem_inst__abc_21203_new_n3078_), .Y(w_mem_inst__abc_21203_new_n3079_));
OR2X2 OR2X2_253 ( .A(_abc_15497_new_n1501_), .B(_abc_15497_new_n1499_), .Y(_abc_15497_new_n1502_));
OR2X2 OR2X2_2530 ( .A(w_mem_inst__abc_21203_new_n3076_), .B(w_mem_inst__abc_21203_new_n3079_), .Y(w_mem_inst__abc_21203_new_n3080_));
OR2X2 OR2X2_2531 ( .A(w_mem_inst__abc_21203_new_n3082_), .B(w_mem_inst__abc_21203_new_n3083_), .Y(w_mem_inst__abc_21203_new_n3084_));
OR2X2 OR2X2_2532 ( .A(w_mem_inst__abc_21203_new_n3084_), .B(w_mem_inst__abc_21203_new_n3081_), .Y(w_mem_inst__abc_21203_new_n3085_));
OR2X2 OR2X2_2533 ( .A(w_mem_inst__abc_21203_new_n3086_), .B(w_mem_inst__abc_21203_new_n3087_), .Y(w_mem_inst__abc_21203_new_n3088_));
OR2X2 OR2X2_2534 ( .A(w_mem_inst__abc_21203_new_n3089_), .B(w_mem_inst__abc_21203_new_n3090_), .Y(w_mem_inst__abc_21203_new_n3091_));
OR2X2 OR2X2_2535 ( .A(w_mem_inst__abc_21203_new_n3088_), .B(w_mem_inst__abc_21203_new_n3091_), .Y(w_mem_inst__abc_21203_new_n3092_));
OR2X2 OR2X2_2536 ( .A(w_mem_inst__abc_21203_new_n3093_), .B(w_mem_inst__abc_21203_new_n3094_), .Y(w_mem_inst__abc_21203_new_n3095_));
OR2X2 OR2X2_2537 ( .A(w_mem_inst__abc_21203_new_n3096_), .B(w_mem_inst__abc_21203_new_n3097_), .Y(w_mem_inst__abc_21203_new_n3098_));
OR2X2 OR2X2_2538 ( .A(w_mem_inst__abc_21203_new_n3095_), .B(w_mem_inst__abc_21203_new_n3098_), .Y(w_mem_inst__abc_21203_new_n3099_));
OR2X2 OR2X2_2539 ( .A(w_mem_inst__abc_21203_new_n3092_), .B(w_mem_inst__abc_21203_new_n3099_), .Y(w_mem_inst__abc_21203_new_n3100_));
OR2X2 OR2X2_254 ( .A(_abc_15497_new_n1505_), .B(_abc_15497_new_n1504_), .Y(_abc_15497_new_n1506_));
OR2X2 OR2X2_2540 ( .A(w_mem_inst__abc_21203_new_n3100_), .B(w_mem_inst__abc_21203_new_n3085_), .Y(w_mem_inst__abc_21203_new_n3101_));
OR2X2 OR2X2_2541 ( .A(w_mem_inst__abc_21203_new_n3101_), .B(w_mem_inst__abc_21203_new_n3080_), .Y(w_mem_inst__abc_21203_new_n3102_));
OR2X2 OR2X2_2542 ( .A(w_mem_inst__abc_21203_new_n3104_), .B(w_mem_inst_w_mem_8__30_), .Y(w_mem_inst__abc_21203_new_n3105_));
OR2X2 OR2X2_2543 ( .A(w_mem_inst__abc_21203_new_n3106_), .B(w_mem_inst_w_mem_13__30_), .Y(w_mem_inst__abc_21203_new_n3107_));
OR2X2 OR2X2_2544 ( .A(w_mem_inst_w_mem_2__30_), .B(w_mem_inst_w_mem_0__30_), .Y(w_mem_inst__abc_21203_new_n3110_));
OR2X2 OR2X2_2545 ( .A(w_mem_inst__abc_21203_new_n3109_), .B(w_mem_inst__abc_21203_new_n3113_), .Y(w_mem_inst__abc_21203_new_n3114_));
OR2X2 OR2X2_2546 ( .A(w_mem_inst__abc_21203_new_n3115_), .B(w_mem_inst__abc_21203_new_n3108_), .Y(w_mem_inst__abc_21203_new_n3116_));
OR2X2 OR2X2_2547 ( .A(w_mem_inst__abc_21203_new_n3117_), .B(w_mem_inst__abc_21203_new_n1587_), .Y(w_mem_inst__abc_21203_new_n3118_));
OR2X2 OR2X2_2548 ( .A(w_mem_inst__abc_21203_new_n3119_), .B(w_mem_inst__abc_21203_new_n1586_), .Y(w_mem_inst__abc_21203_new_n3120_));
OR2X2 OR2X2_2549 ( .A(w_mem_inst__abc_21203_new_n3121_), .B(w_mem_inst__abc_21203_new_n3122_), .Y(w_mem_inst__abc_21203_new_n3123_));
OR2X2 OR2X2_255 ( .A(_abc_15497_new_n1506_), .B(_abc_15497_new_n1503_), .Y(_abc_15497_new_n1507_));
OR2X2 OR2X2_2550 ( .A(w_mem_inst__abc_21203_new_n3123_), .B(w_mem_inst__abc_21203_new_n3120_), .Y(w_mem_inst__abc_21203_new_n3124_));
OR2X2 OR2X2_2551 ( .A(w_mem_inst__abc_21203_new_n3125_), .B(w_mem_inst__abc_21203_new_n3126_), .Y(w_mem_inst__abc_21203_new_n3127_));
OR2X2 OR2X2_2552 ( .A(w_mem_inst__abc_21203_new_n3124_), .B(w_mem_inst__abc_21203_new_n3127_), .Y(w_mem_inst__abc_21203_new_n3128_));
OR2X2 OR2X2_2553 ( .A(w_mem_inst__abc_21203_new_n3130_), .B(w_mem_inst__abc_21203_new_n3131_), .Y(w_mem_inst__abc_21203_new_n3132_));
OR2X2 OR2X2_2554 ( .A(w_mem_inst__abc_21203_new_n3132_), .B(w_mem_inst__abc_21203_new_n3129_), .Y(w_mem_inst__abc_21203_new_n3133_));
OR2X2 OR2X2_2555 ( .A(w_mem_inst__abc_21203_new_n3134_), .B(w_mem_inst__abc_21203_new_n3135_), .Y(w_mem_inst__abc_21203_new_n3136_));
OR2X2 OR2X2_2556 ( .A(w_mem_inst__abc_21203_new_n3137_), .B(w_mem_inst__abc_21203_new_n3138_), .Y(w_mem_inst__abc_21203_new_n3139_));
OR2X2 OR2X2_2557 ( .A(w_mem_inst__abc_21203_new_n3136_), .B(w_mem_inst__abc_21203_new_n3139_), .Y(w_mem_inst__abc_21203_new_n3140_));
OR2X2 OR2X2_2558 ( .A(w_mem_inst__abc_21203_new_n3141_), .B(w_mem_inst__abc_21203_new_n3142_), .Y(w_mem_inst__abc_21203_new_n3143_));
OR2X2 OR2X2_2559 ( .A(w_mem_inst__abc_21203_new_n3144_), .B(w_mem_inst__abc_21203_new_n3145_), .Y(w_mem_inst__abc_21203_new_n3146_));
OR2X2 OR2X2_256 ( .A(_abc_15497_new_n699_), .B(\digest[30] ), .Y(_abc_15497_new_n1510_));
OR2X2 OR2X2_2560 ( .A(w_mem_inst__abc_21203_new_n3143_), .B(w_mem_inst__abc_21203_new_n3146_), .Y(w_mem_inst__abc_21203_new_n3147_));
OR2X2 OR2X2_2561 ( .A(w_mem_inst__abc_21203_new_n3140_), .B(w_mem_inst__abc_21203_new_n3147_), .Y(w_mem_inst__abc_21203_new_n3148_));
OR2X2 OR2X2_2562 ( .A(w_mem_inst__abc_21203_new_n3148_), .B(w_mem_inst__abc_21203_new_n3133_), .Y(w_mem_inst__abc_21203_new_n3149_));
OR2X2 OR2X2_2563 ( .A(w_mem_inst__abc_21203_new_n3149_), .B(w_mem_inst__abc_21203_new_n3128_), .Y(w_mem_inst__abc_21203_new_n3150_));
OR2X2 OR2X2_2564 ( .A(w_mem_inst__abc_21203_new_n3159_), .B(w_mem_inst__abc_21203_new_n3157_), .Y(w_mem_inst__abc_21203_new_n3160_));
OR2X2 OR2X2_2565 ( .A(w_mem_inst__abc_21203_new_n3160_), .B(w_mem_inst__abc_21203_new_n3156_), .Y(w_mem_inst__0w_mem_13__31_0__0_));
OR2X2 OR2X2_2566 ( .A(w_mem_inst__abc_21203_new_n3165_), .B(w_mem_inst__abc_21203_new_n3163_), .Y(w_mem_inst__abc_21203_new_n3166_));
OR2X2 OR2X2_2567 ( .A(w_mem_inst__abc_21203_new_n3166_), .B(w_mem_inst__abc_21203_new_n3162_), .Y(w_mem_inst__0w_mem_13__31_0__1_));
OR2X2 OR2X2_2568 ( .A(w_mem_inst__abc_21203_new_n3171_), .B(w_mem_inst__abc_21203_new_n3169_), .Y(w_mem_inst__abc_21203_new_n3172_));
OR2X2 OR2X2_2569 ( .A(w_mem_inst__abc_21203_new_n3172_), .B(w_mem_inst__abc_21203_new_n3168_), .Y(w_mem_inst__0w_mem_13__31_0__2_));
OR2X2 OR2X2_257 ( .A(_abc_15497_new_n1509_), .B(_abc_15497_new_n1511_), .Y(_0H4_reg_31_0__30_));
OR2X2 OR2X2_2570 ( .A(w_mem_inst__abc_21203_new_n3177_), .B(w_mem_inst__abc_21203_new_n3175_), .Y(w_mem_inst__abc_21203_new_n3178_));
OR2X2 OR2X2_2571 ( .A(w_mem_inst__abc_21203_new_n3178_), .B(w_mem_inst__abc_21203_new_n3174_), .Y(w_mem_inst__0w_mem_13__31_0__3_));
OR2X2 OR2X2_2572 ( .A(w_mem_inst__abc_21203_new_n3183_), .B(w_mem_inst__abc_21203_new_n3181_), .Y(w_mem_inst__abc_21203_new_n3184_));
OR2X2 OR2X2_2573 ( .A(w_mem_inst__abc_21203_new_n3184_), .B(w_mem_inst__abc_21203_new_n3180_), .Y(w_mem_inst__0w_mem_13__31_0__4_));
OR2X2 OR2X2_2574 ( .A(w_mem_inst__abc_21203_new_n3189_), .B(w_mem_inst__abc_21203_new_n3187_), .Y(w_mem_inst__abc_21203_new_n3190_));
OR2X2 OR2X2_2575 ( .A(w_mem_inst__abc_21203_new_n3190_), .B(w_mem_inst__abc_21203_new_n3186_), .Y(w_mem_inst__0w_mem_13__31_0__5_));
OR2X2 OR2X2_2576 ( .A(w_mem_inst__abc_21203_new_n3195_), .B(w_mem_inst__abc_21203_new_n3193_), .Y(w_mem_inst__abc_21203_new_n3196_));
OR2X2 OR2X2_2577 ( .A(w_mem_inst__abc_21203_new_n3196_), .B(w_mem_inst__abc_21203_new_n3192_), .Y(w_mem_inst__0w_mem_13__31_0__6_));
OR2X2 OR2X2_2578 ( .A(w_mem_inst__abc_21203_new_n3201_), .B(w_mem_inst__abc_21203_new_n3199_), .Y(w_mem_inst__abc_21203_new_n3202_));
OR2X2 OR2X2_2579 ( .A(w_mem_inst__abc_21203_new_n3202_), .B(w_mem_inst__abc_21203_new_n3198_), .Y(w_mem_inst__0w_mem_13__31_0__7_));
OR2X2 OR2X2_258 ( .A(_abc_15497_new_n1513_), .B(_abc_15497_new_n1497_), .Y(_abc_15497_new_n1514_));
OR2X2 OR2X2_2580 ( .A(w_mem_inst__abc_21203_new_n3207_), .B(w_mem_inst__abc_21203_new_n3205_), .Y(w_mem_inst__abc_21203_new_n3208_));
OR2X2 OR2X2_2581 ( .A(w_mem_inst__abc_21203_new_n3208_), .B(w_mem_inst__abc_21203_new_n3204_), .Y(w_mem_inst__0w_mem_13__31_0__8_));
OR2X2 OR2X2_2582 ( .A(w_mem_inst__abc_21203_new_n3213_), .B(w_mem_inst__abc_21203_new_n3211_), .Y(w_mem_inst__abc_21203_new_n3214_));
OR2X2 OR2X2_2583 ( .A(w_mem_inst__abc_21203_new_n3214_), .B(w_mem_inst__abc_21203_new_n3210_), .Y(w_mem_inst__0w_mem_13__31_0__9_));
OR2X2 OR2X2_2584 ( .A(w_mem_inst__abc_21203_new_n3219_), .B(w_mem_inst__abc_21203_new_n3217_), .Y(w_mem_inst__abc_21203_new_n3220_));
OR2X2 OR2X2_2585 ( .A(w_mem_inst__abc_21203_new_n3220_), .B(w_mem_inst__abc_21203_new_n3216_), .Y(w_mem_inst__0w_mem_13__31_0__10_));
OR2X2 OR2X2_2586 ( .A(w_mem_inst__abc_21203_new_n3225_), .B(w_mem_inst__abc_21203_new_n3223_), .Y(w_mem_inst__abc_21203_new_n3226_));
OR2X2 OR2X2_2587 ( .A(w_mem_inst__abc_21203_new_n3226_), .B(w_mem_inst__abc_21203_new_n3222_), .Y(w_mem_inst__0w_mem_13__31_0__11_));
OR2X2 OR2X2_2588 ( .A(w_mem_inst__abc_21203_new_n3231_), .B(w_mem_inst__abc_21203_new_n3229_), .Y(w_mem_inst__abc_21203_new_n3232_));
OR2X2 OR2X2_2589 ( .A(w_mem_inst__abc_21203_new_n3232_), .B(w_mem_inst__abc_21203_new_n3228_), .Y(w_mem_inst__0w_mem_13__31_0__12_));
OR2X2 OR2X2_259 ( .A(_abc_15497_new_n1515_), .B(\digest[31] ), .Y(_abc_15497_new_n1516_));
OR2X2 OR2X2_2590 ( .A(w_mem_inst__abc_21203_new_n3237_), .B(w_mem_inst__abc_21203_new_n3235_), .Y(w_mem_inst__abc_21203_new_n3238_));
OR2X2 OR2X2_2591 ( .A(w_mem_inst__abc_21203_new_n3238_), .B(w_mem_inst__abc_21203_new_n3234_), .Y(w_mem_inst__0w_mem_13__31_0__13_));
OR2X2 OR2X2_2592 ( .A(w_mem_inst__abc_21203_new_n3243_), .B(w_mem_inst__abc_21203_new_n3241_), .Y(w_mem_inst__abc_21203_new_n3244_));
OR2X2 OR2X2_2593 ( .A(w_mem_inst__abc_21203_new_n3244_), .B(w_mem_inst__abc_21203_new_n3240_), .Y(w_mem_inst__0w_mem_13__31_0__14_));
OR2X2 OR2X2_2594 ( .A(w_mem_inst__abc_21203_new_n3249_), .B(w_mem_inst__abc_21203_new_n3247_), .Y(w_mem_inst__abc_21203_new_n3250_));
OR2X2 OR2X2_2595 ( .A(w_mem_inst__abc_21203_new_n3250_), .B(w_mem_inst__abc_21203_new_n3246_), .Y(w_mem_inst__0w_mem_13__31_0__15_));
OR2X2 OR2X2_2596 ( .A(w_mem_inst__abc_21203_new_n3255_), .B(w_mem_inst__abc_21203_new_n3253_), .Y(w_mem_inst__abc_21203_new_n3256_));
OR2X2 OR2X2_2597 ( .A(w_mem_inst__abc_21203_new_n3256_), .B(w_mem_inst__abc_21203_new_n3252_), .Y(w_mem_inst__0w_mem_13__31_0__16_));
OR2X2 OR2X2_2598 ( .A(w_mem_inst__abc_21203_new_n3261_), .B(w_mem_inst__abc_21203_new_n3259_), .Y(w_mem_inst__abc_21203_new_n3262_));
OR2X2 OR2X2_2599 ( .A(w_mem_inst__abc_21203_new_n3262_), .B(w_mem_inst__abc_21203_new_n3258_), .Y(w_mem_inst__0w_mem_13__31_0__17_));
OR2X2 OR2X2_26 ( .A(c_reg_7_), .B(\digest[71] ), .Y(_abc_15497_new_n802_));
OR2X2 OR2X2_260 ( .A(_abc_15497_new_n1517_), .B(e_reg_31_), .Y(_abc_15497_new_n1518_));
OR2X2 OR2X2_2600 ( .A(w_mem_inst__abc_21203_new_n3267_), .B(w_mem_inst__abc_21203_new_n3265_), .Y(w_mem_inst__abc_21203_new_n3268_));
OR2X2 OR2X2_2601 ( .A(w_mem_inst__abc_21203_new_n3268_), .B(w_mem_inst__abc_21203_new_n3264_), .Y(w_mem_inst__0w_mem_13__31_0__18_));
OR2X2 OR2X2_2602 ( .A(w_mem_inst__abc_21203_new_n3273_), .B(w_mem_inst__abc_21203_new_n3271_), .Y(w_mem_inst__abc_21203_new_n3274_));
OR2X2 OR2X2_2603 ( .A(w_mem_inst__abc_21203_new_n3274_), .B(w_mem_inst__abc_21203_new_n3270_), .Y(w_mem_inst__0w_mem_13__31_0__19_));
OR2X2 OR2X2_2604 ( .A(w_mem_inst__abc_21203_new_n3279_), .B(w_mem_inst__abc_21203_new_n3277_), .Y(w_mem_inst__abc_21203_new_n3280_));
OR2X2 OR2X2_2605 ( .A(w_mem_inst__abc_21203_new_n3280_), .B(w_mem_inst__abc_21203_new_n3276_), .Y(w_mem_inst__0w_mem_13__31_0__20_));
OR2X2 OR2X2_2606 ( .A(w_mem_inst__abc_21203_new_n3285_), .B(w_mem_inst__abc_21203_new_n3283_), .Y(w_mem_inst__abc_21203_new_n3286_));
OR2X2 OR2X2_2607 ( .A(w_mem_inst__abc_21203_new_n3286_), .B(w_mem_inst__abc_21203_new_n3282_), .Y(w_mem_inst__0w_mem_13__31_0__21_));
OR2X2 OR2X2_2608 ( .A(w_mem_inst__abc_21203_new_n3291_), .B(w_mem_inst__abc_21203_new_n3289_), .Y(w_mem_inst__abc_21203_new_n3292_));
OR2X2 OR2X2_2609 ( .A(w_mem_inst__abc_21203_new_n3292_), .B(w_mem_inst__abc_21203_new_n3288_), .Y(w_mem_inst__0w_mem_13__31_0__22_));
OR2X2 OR2X2_261 ( .A(_abc_15497_new_n1514_), .B(_abc_15497_new_n1520_), .Y(_abc_15497_new_n1521_));
OR2X2 OR2X2_2610 ( .A(w_mem_inst__abc_21203_new_n3297_), .B(w_mem_inst__abc_21203_new_n3295_), .Y(w_mem_inst__abc_21203_new_n3298_));
OR2X2 OR2X2_2611 ( .A(w_mem_inst__abc_21203_new_n3298_), .B(w_mem_inst__abc_21203_new_n3294_), .Y(w_mem_inst__0w_mem_13__31_0__23_));
OR2X2 OR2X2_2612 ( .A(w_mem_inst__abc_21203_new_n3303_), .B(w_mem_inst__abc_21203_new_n3301_), .Y(w_mem_inst__abc_21203_new_n3304_));
OR2X2 OR2X2_2613 ( .A(w_mem_inst__abc_21203_new_n3304_), .B(w_mem_inst__abc_21203_new_n3300_), .Y(w_mem_inst__0w_mem_13__31_0__24_));
OR2X2 OR2X2_2614 ( .A(w_mem_inst__abc_21203_new_n3309_), .B(w_mem_inst__abc_21203_new_n3307_), .Y(w_mem_inst__abc_21203_new_n3310_));
OR2X2 OR2X2_2615 ( .A(w_mem_inst__abc_21203_new_n3310_), .B(w_mem_inst__abc_21203_new_n3306_), .Y(w_mem_inst__0w_mem_13__31_0__25_));
OR2X2 OR2X2_2616 ( .A(w_mem_inst__abc_21203_new_n3315_), .B(w_mem_inst__abc_21203_new_n3313_), .Y(w_mem_inst__abc_21203_new_n3316_));
OR2X2 OR2X2_2617 ( .A(w_mem_inst__abc_21203_new_n3316_), .B(w_mem_inst__abc_21203_new_n3312_), .Y(w_mem_inst__0w_mem_13__31_0__26_));
OR2X2 OR2X2_2618 ( .A(w_mem_inst__abc_21203_new_n3321_), .B(w_mem_inst__abc_21203_new_n3319_), .Y(w_mem_inst__abc_21203_new_n3322_));
OR2X2 OR2X2_2619 ( .A(w_mem_inst__abc_21203_new_n3322_), .B(w_mem_inst__abc_21203_new_n3318_), .Y(w_mem_inst__0w_mem_13__31_0__27_));
OR2X2 OR2X2_262 ( .A(_abc_15497_new_n1522_), .B(_abc_15497_new_n1519_), .Y(_abc_15497_new_n1523_));
OR2X2 OR2X2_2620 ( .A(w_mem_inst__abc_21203_new_n3327_), .B(w_mem_inst__abc_21203_new_n3325_), .Y(w_mem_inst__abc_21203_new_n3328_));
OR2X2 OR2X2_2621 ( .A(w_mem_inst__abc_21203_new_n3328_), .B(w_mem_inst__abc_21203_new_n3324_), .Y(w_mem_inst__0w_mem_13__31_0__28_));
OR2X2 OR2X2_2622 ( .A(w_mem_inst__abc_21203_new_n3333_), .B(w_mem_inst__abc_21203_new_n3331_), .Y(w_mem_inst__abc_21203_new_n3334_));
OR2X2 OR2X2_2623 ( .A(w_mem_inst__abc_21203_new_n3334_), .B(w_mem_inst__abc_21203_new_n3330_), .Y(w_mem_inst__0w_mem_13__31_0__29_));
OR2X2 OR2X2_2624 ( .A(w_mem_inst__abc_21203_new_n3339_), .B(w_mem_inst__abc_21203_new_n3337_), .Y(w_mem_inst__abc_21203_new_n3340_));
OR2X2 OR2X2_2625 ( .A(w_mem_inst__abc_21203_new_n3340_), .B(w_mem_inst__abc_21203_new_n3336_), .Y(w_mem_inst__0w_mem_13__31_0__30_));
OR2X2 OR2X2_2626 ( .A(w_mem_inst__abc_21203_new_n3345_), .B(w_mem_inst__abc_21203_new_n3343_), .Y(w_mem_inst__abc_21203_new_n3346_));
OR2X2 OR2X2_2627 ( .A(w_mem_inst__abc_21203_new_n3346_), .B(w_mem_inst__abc_21203_new_n3342_), .Y(w_mem_inst__0w_mem_13__31_0__31_));
OR2X2 OR2X2_2628 ( .A(w_mem_inst__abc_21203_new_n3350_), .B(w_mem_inst__abc_21203_new_n3349_), .Y(w_mem_inst__abc_21203_new_n3351_));
OR2X2 OR2X2_2629 ( .A(w_mem_inst__abc_21203_new_n3348_), .B(w_mem_inst__abc_21203_new_n3352_), .Y(w_mem_inst__0w_mem_15__31_0__0_));
OR2X2 OR2X2_263 ( .A(_abc_15497_new_n699_), .B(\digest[31] ), .Y(_abc_15497_new_n1526_));
OR2X2 OR2X2_2630 ( .A(w_mem_inst__abc_21203_new_n3355_), .B(w_mem_inst__abc_21203_new_n3354_), .Y(w_mem_inst__abc_21203_new_n3356_));
OR2X2 OR2X2_2631 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst__abc_21203_new_n3356_), .Y(w_mem_inst__abc_21203_new_n3357_));
OR2X2 OR2X2_2632 ( .A(w_mem_inst__abc_21203_new_n1677_), .B(w_mem_inst__abc_21203_new_n3154_), .Y(w_mem_inst__abc_21203_new_n3358_));
OR2X2 OR2X2_2633 ( .A(w_mem_inst__abc_21203_new_n3361_), .B(w_mem_inst__abc_21203_new_n3360_), .Y(w_mem_inst__abc_21203_new_n3362_));
OR2X2 OR2X2_2634 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst__abc_21203_new_n3362_), .Y(w_mem_inst__abc_21203_new_n3363_));
OR2X2 OR2X2_2635 ( .A(w_mem_inst__abc_21203_new_n1725_), .B(w_mem_inst__abc_21203_new_n3154_), .Y(w_mem_inst__abc_21203_new_n3364_));
OR2X2 OR2X2_2636 ( .A(w_mem_inst__abc_21203_new_n3368_), .B(w_mem_inst__abc_21203_new_n3367_), .Y(w_mem_inst__abc_21203_new_n3369_));
OR2X2 OR2X2_2637 ( .A(w_mem_inst__abc_21203_new_n3366_), .B(w_mem_inst__abc_21203_new_n3370_), .Y(w_mem_inst__0w_mem_15__31_0__3_));
OR2X2 OR2X2_2638 ( .A(w_mem_inst__abc_21203_new_n3373_), .B(w_mem_inst__abc_21203_new_n3372_), .Y(w_mem_inst__abc_21203_new_n3374_));
OR2X2 OR2X2_2639 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst__abc_21203_new_n3374_), .Y(w_mem_inst__abc_21203_new_n3375_));
OR2X2 OR2X2_264 ( .A(_abc_15497_new_n1525_), .B(_abc_15497_new_n1527_), .Y(_0H4_reg_31_0__31_));
OR2X2 OR2X2_2640 ( .A(w_mem_inst__abc_21203_new_n1821_), .B(w_mem_inst__abc_21203_new_n3154_), .Y(w_mem_inst__abc_21203_new_n3376_));
OR2X2 OR2X2_2641 ( .A(w_mem_inst__abc_21203_new_n3380_), .B(w_mem_inst__abc_21203_new_n3379_), .Y(w_mem_inst__abc_21203_new_n3381_));
OR2X2 OR2X2_2642 ( .A(w_mem_inst__abc_21203_new_n3378_), .B(w_mem_inst__abc_21203_new_n3382_), .Y(w_mem_inst__0w_mem_15__31_0__5_));
OR2X2 OR2X2_2643 ( .A(w_mem_inst__abc_21203_new_n3386_), .B(w_mem_inst__abc_21203_new_n3385_), .Y(w_mem_inst__abc_21203_new_n3387_));
OR2X2 OR2X2_2644 ( .A(w_mem_inst__abc_21203_new_n3384_), .B(w_mem_inst__abc_21203_new_n3388_), .Y(w_mem_inst__0w_mem_15__31_0__6_));
OR2X2 OR2X2_2645 ( .A(w_mem_inst__abc_21203_new_n3392_), .B(w_mem_inst__abc_21203_new_n3391_), .Y(w_mem_inst__abc_21203_new_n3393_));
OR2X2 OR2X2_2646 ( .A(w_mem_inst__abc_21203_new_n3390_), .B(w_mem_inst__abc_21203_new_n3394_), .Y(w_mem_inst__0w_mem_15__31_0__7_));
OR2X2 OR2X2_2647 ( .A(w_mem_inst__abc_21203_new_n3397_), .B(w_mem_inst__abc_21203_new_n3396_), .Y(w_mem_inst__abc_21203_new_n3398_));
OR2X2 OR2X2_2648 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst__abc_21203_new_n3398_), .Y(w_mem_inst__abc_21203_new_n3399_));
OR2X2 OR2X2_2649 ( .A(w_mem_inst__abc_21203_new_n2013_), .B(w_mem_inst__abc_21203_new_n3154_), .Y(w_mem_inst__abc_21203_new_n3400_));
OR2X2 OR2X2_265 ( .A(\digest[32] ), .B(d_reg_0_), .Y(_abc_15497_new_n1531_));
OR2X2 OR2X2_2650 ( .A(w_mem_inst__abc_21203_new_n3403_), .B(w_mem_inst__abc_21203_new_n3402_), .Y(w_mem_inst__abc_21203_new_n3404_));
OR2X2 OR2X2_2651 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst__abc_21203_new_n3404_), .Y(w_mem_inst__abc_21203_new_n3405_));
OR2X2 OR2X2_2652 ( .A(w_mem_inst__abc_21203_new_n2061_), .B(w_mem_inst__abc_21203_new_n3154_), .Y(w_mem_inst__abc_21203_new_n3406_));
OR2X2 OR2X2_2653 ( .A(w_mem_inst__abc_21203_new_n3410_), .B(w_mem_inst__abc_21203_new_n3409_), .Y(w_mem_inst__abc_21203_new_n3411_));
OR2X2 OR2X2_2654 ( .A(w_mem_inst__abc_21203_new_n3408_), .B(w_mem_inst__abc_21203_new_n3412_), .Y(w_mem_inst__0w_mem_15__31_0__10_));
OR2X2 OR2X2_2655 ( .A(w_mem_inst__abc_21203_new_n3416_), .B(w_mem_inst__abc_21203_new_n3415_), .Y(w_mem_inst__abc_21203_new_n3417_));
OR2X2 OR2X2_2656 ( .A(w_mem_inst__abc_21203_new_n3414_), .B(w_mem_inst__abc_21203_new_n3418_), .Y(w_mem_inst__0w_mem_15__31_0__11_));
OR2X2 OR2X2_2657 ( .A(w_mem_inst__abc_21203_new_n3421_), .B(w_mem_inst__abc_21203_new_n3420_), .Y(w_mem_inst__abc_21203_new_n3422_));
OR2X2 OR2X2_2658 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst__abc_21203_new_n3422_), .Y(w_mem_inst__abc_21203_new_n3423_));
OR2X2 OR2X2_2659 ( .A(w_mem_inst__abc_21203_new_n2205_), .B(w_mem_inst__abc_21203_new_n3154_), .Y(w_mem_inst__abc_21203_new_n3424_));
OR2X2 OR2X2_266 ( .A(_abc_15497_new_n1534_), .B(_abc_15497_new_n1533_), .Y(_0H3_reg_31_0__0_));
OR2X2 OR2X2_2660 ( .A(w_mem_inst__abc_21203_new_n3428_), .B(w_mem_inst__abc_21203_new_n3427_), .Y(w_mem_inst__abc_21203_new_n3429_));
OR2X2 OR2X2_2661 ( .A(w_mem_inst__abc_21203_new_n3426_), .B(w_mem_inst__abc_21203_new_n3430_), .Y(w_mem_inst__0w_mem_15__31_0__13_));
OR2X2 OR2X2_2662 ( .A(w_mem_inst__abc_21203_new_n3434_), .B(w_mem_inst__abc_21203_new_n3433_), .Y(w_mem_inst__abc_21203_new_n3435_));
OR2X2 OR2X2_2663 ( .A(w_mem_inst__abc_21203_new_n3432_), .B(w_mem_inst__abc_21203_new_n3436_), .Y(w_mem_inst__0w_mem_15__31_0__14_));
OR2X2 OR2X2_2664 ( .A(w_mem_inst__abc_21203_new_n3439_), .B(w_mem_inst__abc_21203_new_n3438_), .Y(w_mem_inst__abc_21203_new_n3440_));
OR2X2 OR2X2_2665 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst__abc_21203_new_n3440_), .Y(w_mem_inst__abc_21203_new_n3441_));
OR2X2 OR2X2_2666 ( .A(w_mem_inst__abc_21203_new_n2349_), .B(w_mem_inst__abc_21203_new_n3154_), .Y(w_mem_inst__abc_21203_new_n3442_));
OR2X2 OR2X2_2667 ( .A(w_mem_inst__abc_21203_new_n3446_), .B(w_mem_inst__abc_21203_new_n3445_), .Y(w_mem_inst__abc_21203_new_n3447_));
OR2X2 OR2X2_2668 ( .A(w_mem_inst__abc_21203_new_n3444_), .B(w_mem_inst__abc_21203_new_n3448_), .Y(w_mem_inst__0w_mem_15__31_0__16_));
OR2X2 OR2X2_2669 ( .A(w_mem_inst__abc_21203_new_n3452_), .B(w_mem_inst__abc_21203_new_n3451_), .Y(w_mem_inst__abc_21203_new_n3453_));
OR2X2 OR2X2_267 ( .A(\digest[33] ), .B(d_reg_1_), .Y(_abc_15497_new_n1536_));
OR2X2 OR2X2_2670 ( .A(w_mem_inst__abc_21203_new_n3450_), .B(w_mem_inst__abc_21203_new_n3454_), .Y(w_mem_inst__0w_mem_15__31_0__17_));
OR2X2 OR2X2_2671 ( .A(w_mem_inst__abc_21203_new_n3458_), .B(w_mem_inst__abc_21203_new_n3457_), .Y(w_mem_inst__abc_21203_new_n3459_));
OR2X2 OR2X2_2672 ( .A(w_mem_inst__abc_21203_new_n3456_), .B(w_mem_inst__abc_21203_new_n3460_), .Y(w_mem_inst__0w_mem_15__31_0__18_));
OR2X2 OR2X2_2673 ( .A(w_mem_inst__abc_21203_new_n3464_), .B(w_mem_inst__abc_21203_new_n3463_), .Y(w_mem_inst__abc_21203_new_n3465_));
OR2X2 OR2X2_2674 ( .A(w_mem_inst__abc_21203_new_n3462_), .B(w_mem_inst__abc_21203_new_n3466_), .Y(w_mem_inst__0w_mem_15__31_0__19_));
OR2X2 OR2X2_2675 ( .A(w_mem_inst__abc_21203_new_n3470_), .B(w_mem_inst__abc_21203_new_n3469_), .Y(w_mem_inst__abc_21203_new_n3471_));
OR2X2 OR2X2_2676 ( .A(w_mem_inst__abc_21203_new_n3468_), .B(w_mem_inst__abc_21203_new_n3472_), .Y(w_mem_inst__0w_mem_15__31_0__20_));
OR2X2 OR2X2_2677 ( .A(w_mem_inst__abc_21203_new_n3476_), .B(w_mem_inst__abc_21203_new_n3475_), .Y(w_mem_inst__abc_21203_new_n3477_));
OR2X2 OR2X2_2678 ( .A(w_mem_inst__abc_21203_new_n3474_), .B(w_mem_inst__abc_21203_new_n3478_), .Y(w_mem_inst__0w_mem_15__31_0__21_));
OR2X2 OR2X2_2679 ( .A(w_mem_inst__abc_21203_new_n3482_), .B(w_mem_inst__abc_21203_new_n3481_), .Y(w_mem_inst__abc_21203_new_n3483_));
OR2X2 OR2X2_268 ( .A(_abc_15497_new_n1539_), .B(_abc_15497_new_n1529_), .Y(_abc_15497_new_n1542_));
OR2X2 OR2X2_2680 ( .A(w_mem_inst__abc_21203_new_n3480_), .B(w_mem_inst__abc_21203_new_n3484_), .Y(w_mem_inst__0w_mem_15__31_0__22_));
OR2X2 OR2X2_2681 ( .A(w_mem_inst__abc_21203_new_n3488_), .B(w_mem_inst__abc_21203_new_n3487_), .Y(w_mem_inst__abc_21203_new_n3489_));
OR2X2 OR2X2_2682 ( .A(w_mem_inst__abc_21203_new_n3486_), .B(w_mem_inst__abc_21203_new_n3490_), .Y(w_mem_inst__0w_mem_15__31_0__23_));
OR2X2 OR2X2_2683 ( .A(w_mem_inst__abc_21203_new_n3493_), .B(w_mem_inst__abc_21203_new_n3492_), .Y(w_mem_inst__abc_21203_new_n3494_));
OR2X2 OR2X2_2684 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst__abc_21203_new_n3494_), .Y(w_mem_inst__abc_21203_new_n3495_));
OR2X2 OR2X2_2685 ( .A(w_mem_inst__abc_21203_new_n2781_), .B(w_mem_inst__abc_21203_new_n3154_), .Y(w_mem_inst__abc_21203_new_n3496_));
OR2X2 OR2X2_2686 ( .A(w_mem_inst__abc_21203_new_n3499_), .B(w_mem_inst__abc_21203_new_n3498_), .Y(w_mem_inst__abc_21203_new_n3500_));
OR2X2 OR2X2_2687 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst__abc_21203_new_n3500_), .Y(w_mem_inst__abc_21203_new_n3501_));
OR2X2 OR2X2_2688 ( .A(w_mem_inst__abc_21203_new_n2829_), .B(w_mem_inst__abc_21203_new_n3154_), .Y(w_mem_inst__abc_21203_new_n3502_));
OR2X2 OR2X2_2689 ( .A(w_mem_inst__abc_21203_new_n3506_), .B(w_mem_inst__abc_21203_new_n3505_), .Y(w_mem_inst__abc_21203_new_n3507_));
OR2X2 OR2X2_269 ( .A(_abc_15497_new_n1543_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n1544_));
OR2X2 OR2X2_2690 ( .A(w_mem_inst__abc_21203_new_n3504_), .B(w_mem_inst__abc_21203_new_n3508_), .Y(w_mem_inst__0w_mem_15__31_0__26_));
OR2X2 OR2X2_2691 ( .A(w_mem_inst__abc_21203_new_n3512_), .B(w_mem_inst__abc_21203_new_n3511_), .Y(w_mem_inst__abc_21203_new_n3513_));
OR2X2 OR2X2_2692 ( .A(w_mem_inst__abc_21203_new_n3510_), .B(w_mem_inst__abc_21203_new_n3514_), .Y(w_mem_inst__0w_mem_15__31_0__27_));
OR2X2 OR2X2_2693 ( .A(w_mem_inst__abc_21203_new_n3517_), .B(w_mem_inst__abc_21203_new_n3516_), .Y(w_mem_inst__abc_21203_new_n3518_));
OR2X2 OR2X2_2694 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst__abc_21203_new_n3518_), .Y(w_mem_inst__abc_21203_new_n3519_));
OR2X2 OR2X2_2695 ( .A(w_mem_inst__abc_21203_new_n2973_), .B(w_mem_inst__abc_21203_new_n3154_), .Y(w_mem_inst__abc_21203_new_n3520_));
OR2X2 OR2X2_2696 ( .A(w_mem_inst__abc_21203_new_n3524_), .B(w_mem_inst__abc_21203_new_n3523_), .Y(w_mem_inst__abc_21203_new_n3525_));
OR2X2 OR2X2_2697 ( .A(w_mem_inst__abc_21203_new_n3522_), .B(w_mem_inst__abc_21203_new_n3526_), .Y(w_mem_inst__0w_mem_15__31_0__29_));
OR2X2 OR2X2_2698 ( .A(w_mem_inst__abc_21203_new_n3530_), .B(w_mem_inst__abc_21203_new_n3529_), .Y(w_mem_inst__abc_21203_new_n3531_));
OR2X2 OR2X2_2699 ( .A(w_mem_inst__abc_21203_new_n3528_), .B(w_mem_inst__abc_21203_new_n3532_), .Y(w_mem_inst__0w_mem_15__31_0__30_));
OR2X2 OR2X2_27 ( .A(_abc_15497_new_n804_), .B(_abc_15497_new_n801_), .Y(_abc_15497_new_n805_));
OR2X2 OR2X2_270 ( .A(_abc_15497_new_n699_), .B(\digest[33] ), .Y(_abc_15497_new_n1545_));
OR2X2 OR2X2_2700 ( .A(w_mem_inst__abc_21203_new_n3535_), .B(w_mem_inst__abc_21203_new_n3534_), .Y(w_mem_inst__abc_21203_new_n3536_));
OR2X2 OR2X2_2701 ( .A(w_mem_inst__abc_21203_new_n3153_), .B(w_mem_inst__abc_21203_new_n3536_), .Y(w_mem_inst__abc_21203_new_n3537_));
OR2X2 OR2X2_2702 ( .A(w_mem_inst__abc_21203_new_n3117_), .B(w_mem_inst__abc_21203_new_n3154_), .Y(w_mem_inst__abc_21203_new_n3538_));
OR2X2 OR2X2_2703 ( .A(w_mem_inst__abc_21203_new_n3543_), .B(w_mem_inst__abc_21203_new_n3541_), .Y(w_mem_inst__abc_21203_new_n3544_));
OR2X2 OR2X2_2704 ( .A(w_mem_inst__abc_21203_new_n3544_), .B(w_mem_inst__abc_21203_new_n3540_), .Y(w_mem_inst__0w_mem_14__31_0__0_));
OR2X2 OR2X2_2705 ( .A(w_mem_inst__abc_21203_new_n3549_), .B(w_mem_inst__abc_21203_new_n3547_), .Y(w_mem_inst__abc_21203_new_n3550_));
OR2X2 OR2X2_2706 ( .A(w_mem_inst__abc_21203_new_n3550_), .B(w_mem_inst__abc_21203_new_n3546_), .Y(w_mem_inst__0w_mem_14__31_0__1_));
OR2X2 OR2X2_2707 ( .A(w_mem_inst__abc_21203_new_n3555_), .B(w_mem_inst__abc_21203_new_n3553_), .Y(w_mem_inst__abc_21203_new_n3556_));
OR2X2 OR2X2_2708 ( .A(w_mem_inst__abc_21203_new_n3556_), .B(w_mem_inst__abc_21203_new_n3552_), .Y(w_mem_inst__0w_mem_14__31_0__2_));
OR2X2 OR2X2_2709 ( .A(w_mem_inst__abc_21203_new_n3561_), .B(w_mem_inst__abc_21203_new_n3559_), .Y(w_mem_inst__abc_21203_new_n3562_));
OR2X2 OR2X2_271 ( .A(_abc_15497_new_n1545_), .B(digest_update), .Y(_abc_15497_new_n1546_));
OR2X2 OR2X2_2710 ( .A(w_mem_inst__abc_21203_new_n3562_), .B(w_mem_inst__abc_21203_new_n3558_), .Y(w_mem_inst__0w_mem_14__31_0__3_));
OR2X2 OR2X2_2711 ( .A(w_mem_inst__abc_21203_new_n3567_), .B(w_mem_inst__abc_21203_new_n3565_), .Y(w_mem_inst__abc_21203_new_n3568_));
OR2X2 OR2X2_2712 ( .A(w_mem_inst__abc_21203_new_n3568_), .B(w_mem_inst__abc_21203_new_n3564_), .Y(w_mem_inst__0w_mem_14__31_0__4_));
OR2X2 OR2X2_2713 ( .A(w_mem_inst__abc_21203_new_n3573_), .B(w_mem_inst__abc_21203_new_n3571_), .Y(w_mem_inst__abc_21203_new_n3574_));
OR2X2 OR2X2_2714 ( .A(w_mem_inst__abc_21203_new_n3574_), .B(w_mem_inst__abc_21203_new_n3570_), .Y(w_mem_inst__0w_mem_14__31_0__5_));
OR2X2 OR2X2_2715 ( .A(w_mem_inst__abc_21203_new_n3579_), .B(w_mem_inst__abc_21203_new_n3577_), .Y(w_mem_inst__abc_21203_new_n3580_));
OR2X2 OR2X2_2716 ( .A(w_mem_inst__abc_21203_new_n3580_), .B(w_mem_inst__abc_21203_new_n3576_), .Y(w_mem_inst__0w_mem_14__31_0__6_));
OR2X2 OR2X2_2717 ( .A(w_mem_inst__abc_21203_new_n3585_), .B(w_mem_inst__abc_21203_new_n3583_), .Y(w_mem_inst__abc_21203_new_n3586_));
OR2X2 OR2X2_2718 ( .A(w_mem_inst__abc_21203_new_n3586_), .B(w_mem_inst__abc_21203_new_n3582_), .Y(w_mem_inst__0w_mem_14__31_0__7_));
OR2X2 OR2X2_2719 ( .A(w_mem_inst__abc_21203_new_n3591_), .B(w_mem_inst__abc_21203_new_n3589_), .Y(w_mem_inst__abc_21203_new_n3592_));
OR2X2 OR2X2_272 ( .A(_abc_15497_new_n1540_), .B(_abc_15497_new_n1537_), .Y(_abc_15497_new_n1548_));
OR2X2 OR2X2_2720 ( .A(w_mem_inst__abc_21203_new_n3592_), .B(w_mem_inst__abc_21203_new_n3588_), .Y(w_mem_inst__0w_mem_14__31_0__8_));
OR2X2 OR2X2_2721 ( .A(w_mem_inst__abc_21203_new_n3597_), .B(w_mem_inst__abc_21203_new_n3595_), .Y(w_mem_inst__abc_21203_new_n3598_));
OR2X2 OR2X2_2722 ( .A(w_mem_inst__abc_21203_new_n3598_), .B(w_mem_inst__abc_21203_new_n3594_), .Y(w_mem_inst__0w_mem_14__31_0__9_));
OR2X2 OR2X2_2723 ( .A(w_mem_inst__abc_21203_new_n3603_), .B(w_mem_inst__abc_21203_new_n3601_), .Y(w_mem_inst__abc_21203_new_n3604_));
OR2X2 OR2X2_2724 ( .A(w_mem_inst__abc_21203_new_n3604_), .B(w_mem_inst__abc_21203_new_n3600_), .Y(w_mem_inst__0w_mem_14__31_0__10_));
OR2X2 OR2X2_2725 ( .A(w_mem_inst__abc_21203_new_n3609_), .B(w_mem_inst__abc_21203_new_n3607_), .Y(w_mem_inst__abc_21203_new_n3610_));
OR2X2 OR2X2_2726 ( .A(w_mem_inst__abc_21203_new_n3610_), .B(w_mem_inst__abc_21203_new_n3606_), .Y(w_mem_inst__0w_mem_14__31_0__11_));
OR2X2 OR2X2_2727 ( .A(w_mem_inst__abc_21203_new_n3615_), .B(w_mem_inst__abc_21203_new_n3613_), .Y(w_mem_inst__abc_21203_new_n3616_));
OR2X2 OR2X2_2728 ( .A(w_mem_inst__abc_21203_new_n3616_), .B(w_mem_inst__abc_21203_new_n3612_), .Y(w_mem_inst__0w_mem_14__31_0__12_));
OR2X2 OR2X2_2729 ( .A(w_mem_inst__abc_21203_new_n3621_), .B(w_mem_inst__abc_21203_new_n3619_), .Y(w_mem_inst__abc_21203_new_n3622_));
OR2X2 OR2X2_273 ( .A(\digest[34] ), .B(d_reg_2_), .Y(_abc_15497_new_n1549_));
OR2X2 OR2X2_2730 ( .A(w_mem_inst__abc_21203_new_n3622_), .B(w_mem_inst__abc_21203_new_n3618_), .Y(w_mem_inst__0w_mem_14__31_0__13_));
OR2X2 OR2X2_2731 ( .A(w_mem_inst__abc_21203_new_n3627_), .B(w_mem_inst__abc_21203_new_n3625_), .Y(w_mem_inst__abc_21203_new_n3628_));
OR2X2 OR2X2_2732 ( .A(w_mem_inst__abc_21203_new_n3628_), .B(w_mem_inst__abc_21203_new_n3624_), .Y(w_mem_inst__0w_mem_14__31_0__14_));
OR2X2 OR2X2_2733 ( .A(w_mem_inst__abc_21203_new_n3633_), .B(w_mem_inst__abc_21203_new_n3631_), .Y(w_mem_inst__abc_21203_new_n3634_));
OR2X2 OR2X2_2734 ( .A(w_mem_inst__abc_21203_new_n3634_), .B(w_mem_inst__abc_21203_new_n3630_), .Y(w_mem_inst__0w_mem_14__31_0__15_));
OR2X2 OR2X2_2735 ( .A(w_mem_inst__abc_21203_new_n3639_), .B(w_mem_inst__abc_21203_new_n3637_), .Y(w_mem_inst__abc_21203_new_n3640_));
OR2X2 OR2X2_2736 ( .A(w_mem_inst__abc_21203_new_n3640_), .B(w_mem_inst__abc_21203_new_n3636_), .Y(w_mem_inst__0w_mem_14__31_0__16_));
OR2X2 OR2X2_2737 ( .A(w_mem_inst__abc_21203_new_n3645_), .B(w_mem_inst__abc_21203_new_n3643_), .Y(w_mem_inst__abc_21203_new_n3646_));
OR2X2 OR2X2_2738 ( .A(w_mem_inst__abc_21203_new_n3646_), .B(w_mem_inst__abc_21203_new_n3642_), .Y(w_mem_inst__0w_mem_14__31_0__17_));
OR2X2 OR2X2_2739 ( .A(w_mem_inst__abc_21203_new_n3651_), .B(w_mem_inst__abc_21203_new_n3649_), .Y(w_mem_inst__abc_21203_new_n3652_));
OR2X2 OR2X2_274 ( .A(_abc_15497_new_n1548_), .B(_abc_15497_new_n1552_), .Y(_abc_15497_new_n1555_));
OR2X2 OR2X2_2740 ( .A(w_mem_inst__abc_21203_new_n3652_), .B(w_mem_inst__abc_21203_new_n3648_), .Y(w_mem_inst__0w_mem_14__31_0__18_));
OR2X2 OR2X2_2741 ( .A(w_mem_inst__abc_21203_new_n3657_), .B(w_mem_inst__abc_21203_new_n3655_), .Y(w_mem_inst__abc_21203_new_n3658_));
OR2X2 OR2X2_2742 ( .A(w_mem_inst__abc_21203_new_n3658_), .B(w_mem_inst__abc_21203_new_n3654_), .Y(w_mem_inst__0w_mem_14__31_0__19_));
OR2X2 OR2X2_2743 ( .A(w_mem_inst__abc_21203_new_n3663_), .B(w_mem_inst__abc_21203_new_n3661_), .Y(w_mem_inst__abc_21203_new_n3664_));
OR2X2 OR2X2_2744 ( .A(w_mem_inst__abc_21203_new_n3664_), .B(w_mem_inst__abc_21203_new_n3660_), .Y(w_mem_inst__0w_mem_14__31_0__20_));
OR2X2 OR2X2_2745 ( .A(w_mem_inst__abc_21203_new_n3669_), .B(w_mem_inst__abc_21203_new_n3667_), .Y(w_mem_inst__abc_21203_new_n3670_));
OR2X2 OR2X2_2746 ( .A(w_mem_inst__abc_21203_new_n3670_), .B(w_mem_inst__abc_21203_new_n3666_), .Y(w_mem_inst__0w_mem_14__31_0__21_));
OR2X2 OR2X2_2747 ( .A(w_mem_inst__abc_21203_new_n3675_), .B(w_mem_inst__abc_21203_new_n3673_), .Y(w_mem_inst__abc_21203_new_n3676_));
OR2X2 OR2X2_2748 ( .A(w_mem_inst__abc_21203_new_n3676_), .B(w_mem_inst__abc_21203_new_n3672_), .Y(w_mem_inst__0w_mem_14__31_0__22_));
OR2X2 OR2X2_2749 ( .A(w_mem_inst__abc_21203_new_n3681_), .B(w_mem_inst__abc_21203_new_n3679_), .Y(w_mem_inst__abc_21203_new_n3682_));
OR2X2 OR2X2_275 ( .A(_abc_15497_new_n1556_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n1557_));
OR2X2 OR2X2_2750 ( .A(w_mem_inst__abc_21203_new_n3682_), .B(w_mem_inst__abc_21203_new_n3678_), .Y(w_mem_inst__0w_mem_14__31_0__23_));
OR2X2 OR2X2_2751 ( .A(w_mem_inst__abc_21203_new_n3687_), .B(w_mem_inst__abc_21203_new_n3685_), .Y(w_mem_inst__abc_21203_new_n3688_));
OR2X2 OR2X2_2752 ( .A(w_mem_inst__abc_21203_new_n3688_), .B(w_mem_inst__abc_21203_new_n3684_), .Y(w_mem_inst__0w_mem_14__31_0__24_));
OR2X2 OR2X2_2753 ( .A(w_mem_inst__abc_21203_new_n3693_), .B(w_mem_inst__abc_21203_new_n3691_), .Y(w_mem_inst__abc_21203_new_n3694_));
OR2X2 OR2X2_2754 ( .A(w_mem_inst__abc_21203_new_n3694_), .B(w_mem_inst__abc_21203_new_n3690_), .Y(w_mem_inst__0w_mem_14__31_0__25_));
OR2X2 OR2X2_2755 ( .A(w_mem_inst__abc_21203_new_n3699_), .B(w_mem_inst__abc_21203_new_n3697_), .Y(w_mem_inst__abc_21203_new_n3700_));
OR2X2 OR2X2_2756 ( .A(w_mem_inst__abc_21203_new_n3700_), .B(w_mem_inst__abc_21203_new_n3696_), .Y(w_mem_inst__0w_mem_14__31_0__26_));
OR2X2 OR2X2_2757 ( .A(w_mem_inst__abc_21203_new_n3705_), .B(w_mem_inst__abc_21203_new_n3703_), .Y(w_mem_inst__abc_21203_new_n3706_));
OR2X2 OR2X2_2758 ( .A(w_mem_inst__abc_21203_new_n3706_), .B(w_mem_inst__abc_21203_new_n3702_), .Y(w_mem_inst__0w_mem_14__31_0__27_));
OR2X2 OR2X2_2759 ( .A(w_mem_inst__abc_21203_new_n3711_), .B(w_mem_inst__abc_21203_new_n3709_), .Y(w_mem_inst__abc_21203_new_n3712_));
OR2X2 OR2X2_276 ( .A(_abc_15497_new_n699_), .B(\digest[34] ), .Y(_abc_15497_new_n1558_));
OR2X2 OR2X2_2760 ( .A(w_mem_inst__abc_21203_new_n3712_), .B(w_mem_inst__abc_21203_new_n3708_), .Y(w_mem_inst__0w_mem_14__31_0__28_));
OR2X2 OR2X2_2761 ( .A(w_mem_inst__abc_21203_new_n3717_), .B(w_mem_inst__abc_21203_new_n3715_), .Y(w_mem_inst__abc_21203_new_n3718_));
OR2X2 OR2X2_2762 ( .A(w_mem_inst__abc_21203_new_n3718_), .B(w_mem_inst__abc_21203_new_n3714_), .Y(w_mem_inst__0w_mem_14__31_0__29_));
OR2X2 OR2X2_2763 ( .A(w_mem_inst__abc_21203_new_n3723_), .B(w_mem_inst__abc_21203_new_n3721_), .Y(w_mem_inst__abc_21203_new_n3724_));
OR2X2 OR2X2_2764 ( .A(w_mem_inst__abc_21203_new_n3724_), .B(w_mem_inst__abc_21203_new_n3720_), .Y(w_mem_inst__0w_mem_14__31_0__30_));
OR2X2 OR2X2_2765 ( .A(w_mem_inst__abc_21203_new_n3729_), .B(w_mem_inst__abc_21203_new_n3727_), .Y(w_mem_inst__abc_21203_new_n3730_));
OR2X2 OR2X2_2766 ( .A(w_mem_inst__abc_21203_new_n3730_), .B(w_mem_inst__abc_21203_new_n3726_), .Y(w_mem_inst__0w_mem_14__31_0__31_));
OR2X2 OR2X2_2767 ( .A(w_mem_inst__abc_21203_new_n3735_), .B(w_mem_inst__abc_21203_new_n3733_), .Y(w_mem_inst__abc_21203_new_n3736_));
OR2X2 OR2X2_2768 ( .A(w_mem_inst__abc_21203_new_n3736_), .B(w_mem_inst__abc_21203_new_n3732_), .Y(w_mem_inst__0w_mem_10__31_0__0_));
OR2X2 OR2X2_2769 ( .A(w_mem_inst__abc_21203_new_n3741_), .B(w_mem_inst__abc_21203_new_n3739_), .Y(w_mem_inst__abc_21203_new_n3742_));
OR2X2 OR2X2_277 ( .A(_abc_15497_new_n1558_), .B(digest_update), .Y(_abc_15497_new_n1559_));
OR2X2 OR2X2_2770 ( .A(w_mem_inst__abc_21203_new_n3742_), .B(w_mem_inst__abc_21203_new_n3738_), .Y(w_mem_inst__0w_mem_10__31_0__1_));
OR2X2 OR2X2_2771 ( .A(w_mem_inst__abc_21203_new_n3747_), .B(w_mem_inst__abc_21203_new_n3745_), .Y(w_mem_inst__abc_21203_new_n3748_));
OR2X2 OR2X2_2772 ( .A(w_mem_inst__abc_21203_new_n3748_), .B(w_mem_inst__abc_21203_new_n3744_), .Y(w_mem_inst__0w_mem_10__31_0__2_));
OR2X2 OR2X2_2773 ( .A(w_mem_inst__abc_21203_new_n3753_), .B(w_mem_inst__abc_21203_new_n3751_), .Y(w_mem_inst__abc_21203_new_n3754_));
OR2X2 OR2X2_2774 ( .A(w_mem_inst__abc_21203_new_n3754_), .B(w_mem_inst__abc_21203_new_n3750_), .Y(w_mem_inst__0w_mem_10__31_0__3_));
OR2X2 OR2X2_2775 ( .A(w_mem_inst__abc_21203_new_n3759_), .B(w_mem_inst__abc_21203_new_n3757_), .Y(w_mem_inst__abc_21203_new_n3760_));
OR2X2 OR2X2_2776 ( .A(w_mem_inst__abc_21203_new_n3760_), .B(w_mem_inst__abc_21203_new_n3756_), .Y(w_mem_inst__0w_mem_10__31_0__4_));
OR2X2 OR2X2_2777 ( .A(w_mem_inst__abc_21203_new_n3765_), .B(w_mem_inst__abc_21203_new_n3763_), .Y(w_mem_inst__abc_21203_new_n3766_));
OR2X2 OR2X2_2778 ( .A(w_mem_inst__abc_21203_new_n3766_), .B(w_mem_inst__abc_21203_new_n3762_), .Y(w_mem_inst__0w_mem_10__31_0__5_));
OR2X2 OR2X2_2779 ( .A(w_mem_inst__abc_21203_new_n3771_), .B(w_mem_inst__abc_21203_new_n3769_), .Y(w_mem_inst__abc_21203_new_n3772_));
OR2X2 OR2X2_278 ( .A(_abc_15497_new_n1553_), .B(_abc_15497_new_n1550_), .Y(_abc_15497_new_n1562_));
OR2X2 OR2X2_2780 ( .A(w_mem_inst__abc_21203_new_n3772_), .B(w_mem_inst__abc_21203_new_n3768_), .Y(w_mem_inst__0w_mem_10__31_0__6_));
OR2X2 OR2X2_2781 ( .A(w_mem_inst__abc_21203_new_n3777_), .B(w_mem_inst__abc_21203_new_n3775_), .Y(w_mem_inst__abc_21203_new_n3778_));
OR2X2 OR2X2_2782 ( .A(w_mem_inst__abc_21203_new_n3778_), .B(w_mem_inst__abc_21203_new_n3774_), .Y(w_mem_inst__0w_mem_10__31_0__7_));
OR2X2 OR2X2_2783 ( .A(w_mem_inst__abc_21203_new_n3783_), .B(w_mem_inst__abc_21203_new_n3781_), .Y(w_mem_inst__abc_21203_new_n3784_));
OR2X2 OR2X2_2784 ( .A(w_mem_inst__abc_21203_new_n3784_), .B(w_mem_inst__abc_21203_new_n3780_), .Y(w_mem_inst__0w_mem_10__31_0__8_));
OR2X2 OR2X2_2785 ( .A(w_mem_inst__abc_21203_new_n3789_), .B(w_mem_inst__abc_21203_new_n3787_), .Y(w_mem_inst__abc_21203_new_n3790_));
OR2X2 OR2X2_2786 ( .A(w_mem_inst__abc_21203_new_n3790_), .B(w_mem_inst__abc_21203_new_n3786_), .Y(w_mem_inst__0w_mem_10__31_0__9_));
OR2X2 OR2X2_2787 ( .A(w_mem_inst__abc_21203_new_n3795_), .B(w_mem_inst__abc_21203_new_n3793_), .Y(w_mem_inst__abc_21203_new_n3796_));
OR2X2 OR2X2_2788 ( .A(w_mem_inst__abc_21203_new_n3796_), .B(w_mem_inst__abc_21203_new_n3792_), .Y(w_mem_inst__0w_mem_10__31_0__10_));
OR2X2 OR2X2_2789 ( .A(w_mem_inst__abc_21203_new_n3801_), .B(w_mem_inst__abc_21203_new_n3799_), .Y(w_mem_inst__abc_21203_new_n3802_));
OR2X2 OR2X2_279 ( .A(\digest[35] ), .B(d_reg_3_), .Y(_abc_15497_new_n1563_));
OR2X2 OR2X2_2790 ( .A(w_mem_inst__abc_21203_new_n3802_), .B(w_mem_inst__abc_21203_new_n3798_), .Y(w_mem_inst__0w_mem_10__31_0__11_));
OR2X2 OR2X2_2791 ( .A(w_mem_inst__abc_21203_new_n3807_), .B(w_mem_inst__abc_21203_new_n3805_), .Y(w_mem_inst__abc_21203_new_n3808_));
OR2X2 OR2X2_2792 ( .A(w_mem_inst__abc_21203_new_n3808_), .B(w_mem_inst__abc_21203_new_n3804_), .Y(w_mem_inst__0w_mem_10__31_0__12_));
OR2X2 OR2X2_2793 ( .A(w_mem_inst__abc_21203_new_n3813_), .B(w_mem_inst__abc_21203_new_n3811_), .Y(w_mem_inst__abc_21203_new_n3814_));
OR2X2 OR2X2_2794 ( .A(w_mem_inst__abc_21203_new_n3814_), .B(w_mem_inst__abc_21203_new_n3810_), .Y(w_mem_inst__0w_mem_10__31_0__13_));
OR2X2 OR2X2_2795 ( .A(w_mem_inst__abc_21203_new_n3819_), .B(w_mem_inst__abc_21203_new_n3817_), .Y(w_mem_inst__abc_21203_new_n3820_));
OR2X2 OR2X2_2796 ( .A(w_mem_inst__abc_21203_new_n3820_), .B(w_mem_inst__abc_21203_new_n3816_), .Y(w_mem_inst__0w_mem_10__31_0__14_));
OR2X2 OR2X2_2797 ( .A(w_mem_inst__abc_21203_new_n3825_), .B(w_mem_inst__abc_21203_new_n3823_), .Y(w_mem_inst__abc_21203_new_n3826_));
OR2X2 OR2X2_2798 ( .A(w_mem_inst__abc_21203_new_n3826_), .B(w_mem_inst__abc_21203_new_n3822_), .Y(w_mem_inst__0w_mem_10__31_0__15_));
OR2X2 OR2X2_2799 ( .A(w_mem_inst__abc_21203_new_n3831_), .B(w_mem_inst__abc_21203_new_n3829_), .Y(w_mem_inst__abc_21203_new_n3832_));
OR2X2 OR2X2_28 ( .A(c_reg_6_), .B(\digest[70] ), .Y(_abc_15497_new_n809_));
OR2X2 OR2X2_280 ( .A(_abc_15497_new_n1562_), .B(_abc_15497_new_n1566_), .Y(_abc_15497_new_n1567_));
OR2X2 OR2X2_2800 ( .A(w_mem_inst__abc_21203_new_n3832_), .B(w_mem_inst__abc_21203_new_n3828_), .Y(w_mem_inst__0w_mem_10__31_0__16_));
OR2X2 OR2X2_2801 ( .A(w_mem_inst__abc_21203_new_n3837_), .B(w_mem_inst__abc_21203_new_n3835_), .Y(w_mem_inst__abc_21203_new_n3838_));
OR2X2 OR2X2_2802 ( .A(w_mem_inst__abc_21203_new_n3838_), .B(w_mem_inst__abc_21203_new_n3834_), .Y(w_mem_inst__0w_mem_10__31_0__17_));
OR2X2 OR2X2_2803 ( .A(w_mem_inst__abc_21203_new_n3843_), .B(w_mem_inst__abc_21203_new_n3841_), .Y(w_mem_inst__abc_21203_new_n3844_));
OR2X2 OR2X2_2804 ( .A(w_mem_inst__abc_21203_new_n3844_), .B(w_mem_inst__abc_21203_new_n3840_), .Y(w_mem_inst__0w_mem_10__31_0__18_));
OR2X2 OR2X2_2805 ( .A(w_mem_inst__abc_21203_new_n3849_), .B(w_mem_inst__abc_21203_new_n3847_), .Y(w_mem_inst__abc_21203_new_n3850_));
OR2X2 OR2X2_2806 ( .A(w_mem_inst__abc_21203_new_n3850_), .B(w_mem_inst__abc_21203_new_n3846_), .Y(w_mem_inst__0w_mem_10__31_0__19_));
OR2X2 OR2X2_2807 ( .A(w_mem_inst__abc_21203_new_n3855_), .B(w_mem_inst__abc_21203_new_n3853_), .Y(w_mem_inst__abc_21203_new_n3856_));
OR2X2 OR2X2_2808 ( .A(w_mem_inst__abc_21203_new_n3856_), .B(w_mem_inst__abc_21203_new_n3852_), .Y(w_mem_inst__0w_mem_10__31_0__20_));
OR2X2 OR2X2_2809 ( .A(w_mem_inst__abc_21203_new_n3861_), .B(w_mem_inst__abc_21203_new_n3859_), .Y(w_mem_inst__abc_21203_new_n3862_));
OR2X2 OR2X2_281 ( .A(_abc_15497_new_n1568_), .B(_abc_15497_new_n1569_), .Y(_abc_15497_new_n1570_));
OR2X2 OR2X2_2810 ( .A(w_mem_inst__abc_21203_new_n3862_), .B(w_mem_inst__abc_21203_new_n3858_), .Y(w_mem_inst__0w_mem_10__31_0__21_));
OR2X2 OR2X2_2811 ( .A(w_mem_inst__abc_21203_new_n3867_), .B(w_mem_inst__abc_21203_new_n3865_), .Y(w_mem_inst__abc_21203_new_n3868_));
OR2X2 OR2X2_2812 ( .A(w_mem_inst__abc_21203_new_n3868_), .B(w_mem_inst__abc_21203_new_n3864_), .Y(w_mem_inst__0w_mem_10__31_0__22_));
OR2X2 OR2X2_2813 ( .A(w_mem_inst__abc_21203_new_n3873_), .B(w_mem_inst__abc_21203_new_n3871_), .Y(w_mem_inst__abc_21203_new_n3874_));
OR2X2 OR2X2_2814 ( .A(w_mem_inst__abc_21203_new_n3874_), .B(w_mem_inst__abc_21203_new_n3870_), .Y(w_mem_inst__0w_mem_10__31_0__23_));
OR2X2 OR2X2_2815 ( .A(w_mem_inst__abc_21203_new_n3879_), .B(w_mem_inst__abc_21203_new_n3877_), .Y(w_mem_inst__abc_21203_new_n3880_));
OR2X2 OR2X2_2816 ( .A(w_mem_inst__abc_21203_new_n3880_), .B(w_mem_inst__abc_21203_new_n3876_), .Y(w_mem_inst__0w_mem_10__31_0__24_));
OR2X2 OR2X2_2817 ( .A(w_mem_inst__abc_21203_new_n3885_), .B(w_mem_inst__abc_21203_new_n3883_), .Y(w_mem_inst__abc_21203_new_n3886_));
OR2X2 OR2X2_2818 ( .A(w_mem_inst__abc_21203_new_n3886_), .B(w_mem_inst__abc_21203_new_n3882_), .Y(w_mem_inst__0w_mem_10__31_0__25_));
OR2X2 OR2X2_2819 ( .A(w_mem_inst__abc_21203_new_n3891_), .B(w_mem_inst__abc_21203_new_n3889_), .Y(w_mem_inst__abc_21203_new_n3892_));
OR2X2 OR2X2_282 ( .A(_abc_15497_new_n1572_), .B(_abc_15497_new_n1561_), .Y(_0H3_reg_31_0__3_));
OR2X2 OR2X2_2820 ( .A(w_mem_inst__abc_21203_new_n3892_), .B(w_mem_inst__abc_21203_new_n3888_), .Y(w_mem_inst__0w_mem_10__31_0__26_));
OR2X2 OR2X2_2821 ( .A(w_mem_inst__abc_21203_new_n3897_), .B(w_mem_inst__abc_21203_new_n3895_), .Y(w_mem_inst__abc_21203_new_n3898_));
OR2X2 OR2X2_2822 ( .A(w_mem_inst__abc_21203_new_n3898_), .B(w_mem_inst__abc_21203_new_n3894_), .Y(w_mem_inst__0w_mem_10__31_0__27_));
OR2X2 OR2X2_2823 ( .A(w_mem_inst__abc_21203_new_n3903_), .B(w_mem_inst__abc_21203_new_n3901_), .Y(w_mem_inst__abc_21203_new_n3904_));
OR2X2 OR2X2_2824 ( .A(w_mem_inst__abc_21203_new_n3904_), .B(w_mem_inst__abc_21203_new_n3900_), .Y(w_mem_inst__0w_mem_10__31_0__28_));
OR2X2 OR2X2_2825 ( .A(w_mem_inst__abc_21203_new_n3909_), .B(w_mem_inst__abc_21203_new_n3907_), .Y(w_mem_inst__abc_21203_new_n3910_));
OR2X2 OR2X2_2826 ( .A(w_mem_inst__abc_21203_new_n3910_), .B(w_mem_inst__abc_21203_new_n3906_), .Y(w_mem_inst__0w_mem_10__31_0__29_));
OR2X2 OR2X2_2827 ( .A(w_mem_inst__abc_21203_new_n3915_), .B(w_mem_inst__abc_21203_new_n3913_), .Y(w_mem_inst__abc_21203_new_n3916_));
OR2X2 OR2X2_2828 ( .A(w_mem_inst__abc_21203_new_n3916_), .B(w_mem_inst__abc_21203_new_n3912_), .Y(w_mem_inst__0w_mem_10__31_0__30_));
OR2X2 OR2X2_2829 ( .A(w_mem_inst__abc_21203_new_n3921_), .B(w_mem_inst__abc_21203_new_n3919_), .Y(w_mem_inst__abc_21203_new_n3922_));
OR2X2 OR2X2_283 ( .A(\digest[36] ), .B(d_reg_4_), .Y(_abc_15497_new_n1574_));
OR2X2 OR2X2_2830 ( .A(w_mem_inst__abc_21203_new_n3922_), .B(w_mem_inst__abc_21203_new_n3918_), .Y(w_mem_inst__0w_mem_10__31_0__31_));
OR2X2 OR2X2_2831 ( .A(w_mem_inst__abc_21203_new_n3927_), .B(w_mem_inst__abc_21203_new_n3925_), .Y(w_mem_inst__abc_21203_new_n3928_));
OR2X2 OR2X2_2832 ( .A(w_mem_inst__abc_21203_new_n3928_), .B(w_mem_inst__abc_21203_new_n3924_), .Y(w_mem_inst__0w_mem_12__31_0__0_));
OR2X2 OR2X2_2833 ( .A(w_mem_inst__abc_21203_new_n3933_), .B(w_mem_inst__abc_21203_new_n3931_), .Y(w_mem_inst__abc_21203_new_n3934_));
OR2X2 OR2X2_2834 ( .A(w_mem_inst__abc_21203_new_n3934_), .B(w_mem_inst__abc_21203_new_n3930_), .Y(w_mem_inst__0w_mem_12__31_0__1_));
OR2X2 OR2X2_2835 ( .A(w_mem_inst__abc_21203_new_n3939_), .B(w_mem_inst__abc_21203_new_n3937_), .Y(w_mem_inst__abc_21203_new_n3940_));
OR2X2 OR2X2_2836 ( .A(w_mem_inst__abc_21203_new_n3940_), .B(w_mem_inst__abc_21203_new_n3936_), .Y(w_mem_inst__0w_mem_12__31_0__2_));
OR2X2 OR2X2_2837 ( .A(w_mem_inst__abc_21203_new_n3945_), .B(w_mem_inst__abc_21203_new_n3943_), .Y(w_mem_inst__abc_21203_new_n3946_));
OR2X2 OR2X2_2838 ( .A(w_mem_inst__abc_21203_new_n3946_), .B(w_mem_inst__abc_21203_new_n3942_), .Y(w_mem_inst__0w_mem_12__31_0__3_));
OR2X2 OR2X2_2839 ( .A(w_mem_inst__abc_21203_new_n3951_), .B(w_mem_inst__abc_21203_new_n3949_), .Y(w_mem_inst__abc_21203_new_n3952_));
OR2X2 OR2X2_284 ( .A(_abc_15497_new_n1578_), .B(_abc_15497_new_n1564_), .Y(_abc_15497_new_n1579_));
OR2X2 OR2X2_2840 ( .A(w_mem_inst__abc_21203_new_n3952_), .B(w_mem_inst__abc_21203_new_n3948_), .Y(w_mem_inst__0w_mem_12__31_0__4_));
OR2X2 OR2X2_2841 ( .A(w_mem_inst__abc_21203_new_n3957_), .B(w_mem_inst__abc_21203_new_n3955_), .Y(w_mem_inst__abc_21203_new_n3958_));
OR2X2 OR2X2_2842 ( .A(w_mem_inst__abc_21203_new_n3958_), .B(w_mem_inst__abc_21203_new_n3954_), .Y(w_mem_inst__0w_mem_12__31_0__5_));
OR2X2 OR2X2_2843 ( .A(w_mem_inst__abc_21203_new_n3963_), .B(w_mem_inst__abc_21203_new_n3961_), .Y(w_mem_inst__abc_21203_new_n3964_));
OR2X2 OR2X2_2844 ( .A(w_mem_inst__abc_21203_new_n3964_), .B(w_mem_inst__abc_21203_new_n3960_), .Y(w_mem_inst__0w_mem_12__31_0__6_));
OR2X2 OR2X2_2845 ( .A(w_mem_inst__abc_21203_new_n3969_), .B(w_mem_inst__abc_21203_new_n3967_), .Y(w_mem_inst__abc_21203_new_n3970_));
OR2X2 OR2X2_2846 ( .A(w_mem_inst__abc_21203_new_n3970_), .B(w_mem_inst__abc_21203_new_n3966_), .Y(w_mem_inst__0w_mem_12__31_0__7_));
OR2X2 OR2X2_2847 ( .A(w_mem_inst__abc_21203_new_n3975_), .B(w_mem_inst__abc_21203_new_n3973_), .Y(w_mem_inst__abc_21203_new_n3976_));
OR2X2 OR2X2_2848 ( .A(w_mem_inst__abc_21203_new_n3976_), .B(w_mem_inst__abc_21203_new_n3972_), .Y(w_mem_inst__0w_mem_12__31_0__8_));
OR2X2 OR2X2_2849 ( .A(w_mem_inst__abc_21203_new_n3981_), .B(w_mem_inst__abc_21203_new_n3979_), .Y(w_mem_inst__abc_21203_new_n3982_));
OR2X2 OR2X2_285 ( .A(_abc_15497_new_n1579_), .B(_abc_15497_new_n1577_), .Y(_abc_15497_new_n1582_));
OR2X2 OR2X2_2850 ( .A(w_mem_inst__abc_21203_new_n3982_), .B(w_mem_inst__abc_21203_new_n3978_), .Y(w_mem_inst__0w_mem_12__31_0__9_));
OR2X2 OR2X2_2851 ( .A(w_mem_inst__abc_21203_new_n3987_), .B(w_mem_inst__abc_21203_new_n3985_), .Y(w_mem_inst__abc_21203_new_n3988_));
OR2X2 OR2X2_2852 ( .A(w_mem_inst__abc_21203_new_n3988_), .B(w_mem_inst__abc_21203_new_n3984_), .Y(w_mem_inst__0w_mem_12__31_0__10_));
OR2X2 OR2X2_2853 ( .A(w_mem_inst__abc_21203_new_n3993_), .B(w_mem_inst__abc_21203_new_n3991_), .Y(w_mem_inst__abc_21203_new_n3994_));
OR2X2 OR2X2_2854 ( .A(w_mem_inst__abc_21203_new_n3994_), .B(w_mem_inst__abc_21203_new_n3990_), .Y(w_mem_inst__0w_mem_12__31_0__11_));
OR2X2 OR2X2_2855 ( .A(w_mem_inst__abc_21203_new_n3999_), .B(w_mem_inst__abc_21203_new_n3997_), .Y(w_mem_inst__abc_21203_new_n4000_));
OR2X2 OR2X2_2856 ( .A(w_mem_inst__abc_21203_new_n4000_), .B(w_mem_inst__abc_21203_new_n3996_), .Y(w_mem_inst__0w_mem_12__31_0__12_));
OR2X2 OR2X2_2857 ( .A(w_mem_inst__abc_21203_new_n4005_), .B(w_mem_inst__abc_21203_new_n4003_), .Y(w_mem_inst__abc_21203_new_n4006_));
OR2X2 OR2X2_2858 ( .A(w_mem_inst__abc_21203_new_n4006_), .B(w_mem_inst__abc_21203_new_n4002_), .Y(w_mem_inst__0w_mem_12__31_0__13_));
OR2X2 OR2X2_2859 ( .A(w_mem_inst__abc_21203_new_n4011_), .B(w_mem_inst__abc_21203_new_n4009_), .Y(w_mem_inst__abc_21203_new_n4012_));
OR2X2 OR2X2_286 ( .A(_abc_15497_new_n1583_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n1584_));
OR2X2 OR2X2_2860 ( .A(w_mem_inst__abc_21203_new_n4012_), .B(w_mem_inst__abc_21203_new_n4008_), .Y(w_mem_inst__0w_mem_12__31_0__14_));
OR2X2 OR2X2_2861 ( .A(w_mem_inst__abc_21203_new_n4017_), .B(w_mem_inst__abc_21203_new_n4015_), .Y(w_mem_inst__abc_21203_new_n4018_));
OR2X2 OR2X2_2862 ( .A(w_mem_inst__abc_21203_new_n4018_), .B(w_mem_inst__abc_21203_new_n4014_), .Y(w_mem_inst__0w_mem_12__31_0__15_));
OR2X2 OR2X2_2863 ( .A(w_mem_inst__abc_21203_new_n4023_), .B(w_mem_inst__abc_21203_new_n4021_), .Y(w_mem_inst__abc_21203_new_n4024_));
OR2X2 OR2X2_2864 ( .A(w_mem_inst__abc_21203_new_n4024_), .B(w_mem_inst__abc_21203_new_n4020_), .Y(w_mem_inst__0w_mem_12__31_0__16_));
OR2X2 OR2X2_2865 ( .A(w_mem_inst__abc_21203_new_n4029_), .B(w_mem_inst__abc_21203_new_n4027_), .Y(w_mem_inst__abc_21203_new_n4030_));
OR2X2 OR2X2_2866 ( .A(w_mem_inst__abc_21203_new_n4030_), .B(w_mem_inst__abc_21203_new_n4026_), .Y(w_mem_inst__0w_mem_12__31_0__17_));
OR2X2 OR2X2_2867 ( .A(w_mem_inst__abc_21203_new_n4035_), .B(w_mem_inst__abc_21203_new_n4033_), .Y(w_mem_inst__abc_21203_new_n4036_));
OR2X2 OR2X2_2868 ( .A(w_mem_inst__abc_21203_new_n4036_), .B(w_mem_inst__abc_21203_new_n4032_), .Y(w_mem_inst__0w_mem_12__31_0__18_));
OR2X2 OR2X2_2869 ( .A(w_mem_inst__abc_21203_new_n4041_), .B(w_mem_inst__abc_21203_new_n4039_), .Y(w_mem_inst__abc_21203_new_n4042_));
OR2X2 OR2X2_287 ( .A(_abc_15497_new_n699_), .B(\digest[36] ), .Y(_abc_15497_new_n1585_));
OR2X2 OR2X2_2870 ( .A(w_mem_inst__abc_21203_new_n4042_), .B(w_mem_inst__abc_21203_new_n4038_), .Y(w_mem_inst__0w_mem_12__31_0__19_));
OR2X2 OR2X2_2871 ( .A(w_mem_inst__abc_21203_new_n4047_), .B(w_mem_inst__abc_21203_new_n4045_), .Y(w_mem_inst__abc_21203_new_n4048_));
OR2X2 OR2X2_2872 ( .A(w_mem_inst__abc_21203_new_n4048_), .B(w_mem_inst__abc_21203_new_n4044_), .Y(w_mem_inst__0w_mem_12__31_0__20_));
OR2X2 OR2X2_2873 ( .A(w_mem_inst__abc_21203_new_n4053_), .B(w_mem_inst__abc_21203_new_n4051_), .Y(w_mem_inst__abc_21203_new_n4054_));
OR2X2 OR2X2_2874 ( .A(w_mem_inst__abc_21203_new_n4054_), .B(w_mem_inst__abc_21203_new_n4050_), .Y(w_mem_inst__0w_mem_12__31_0__21_));
OR2X2 OR2X2_2875 ( .A(w_mem_inst__abc_21203_new_n4059_), .B(w_mem_inst__abc_21203_new_n4057_), .Y(w_mem_inst__abc_21203_new_n4060_));
OR2X2 OR2X2_2876 ( .A(w_mem_inst__abc_21203_new_n4060_), .B(w_mem_inst__abc_21203_new_n4056_), .Y(w_mem_inst__0w_mem_12__31_0__22_));
OR2X2 OR2X2_2877 ( .A(w_mem_inst__abc_21203_new_n4065_), .B(w_mem_inst__abc_21203_new_n4063_), .Y(w_mem_inst__abc_21203_new_n4066_));
OR2X2 OR2X2_2878 ( .A(w_mem_inst__abc_21203_new_n4066_), .B(w_mem_inst__abc_21203_new_n4062_), .Y(w_mem_inst__0w_mem_12__31_0__23_));
OR2X2 OR2X2_2879 ( .A(w_mem_inst__abc_21203_new_n4071_), .B(w_mem_inst__abc_21203_new_n4069_), .Y(w_mem_inst__abc_21203_new_n4072_));
OR2X2 OR2X2_288 ( .A(_abc_15497_new_n1585_), .B(digest_update), .Y(_abc_15497_new_n1586_));
OR2X2 OR2X2_2880 ( .A(w_mem_inst__abc_21203_new_n4072_), .B(w_mem_inst__abc_21203_new_n4068_), .Y(w_mem_inst__0w_mem_12__31_0__24_));
OR2X2 OR2X2_2881 ( .A(w_mem_inst__abc_21203_new_n4077_), .B(w_mem_inst__abc_21203_new_n4075_), .Y(w_mem_inst__abc_21203_new_n4078_));
OR2X2 OR2X2_2882 ( .A(w_mem_inst__abc_21203_new_n4078_), .B(w_mem_inst__abc_21203_new_n4074_), .Y(w_mem_inst__0w_mem_12__31_0__25_));
OR2X2 OR2X2_2883 ( .A(w_mem_inst__abc_21203_new_n4083_), .B(w_mem_inst__abc_21203_new_n4081_), .Y(w_mem_inst__abc_21203_new_n4084_));
OR2X2 OR2X2_2884 ( .A(w_mem_inst__abc_21203_new_n4084_), .B(w_mem_inst__abc_21203_new_n4080_), .Y(w_mem_inst__0w_mem_12__31_0__26_));
OR2X2 OR2X2_2885 ( .A(w_mem_inst__abc_21203_new_n4089_), .B(w_mem_inst__abc_21203_new_n4087_), .Y(w_mem_inst__abc_21203_new_n4090_));
OR2X2 OR2X2_2886 ( .A(w_mem_inst__abc_21203_new_n4090_), .B(w_mem_inst__abc_21203_new_n4086_), .Y(w_mem_inst__0w_mem_12__31_0__27_));
OR2X2 OR2X2_2887 ( .A(w_mem_inst__abc_21203_new_n4095_), .B(w_mem_inst__abc_21203_new_n4093_), .Y(w_mem_inst__abc_21203_new_n4096_));
OR2X2 OR2X2_2888 ( .A(w_mem_inst__abc_21203_new_n4096_), .B(w_mem_inst__abc_21203_new_n4092_), .Y(w_mem_inst__0w_mem_12__31_0__28_));
OR2X2 OR2X2_2889 ( .A(w_mem_inst__abc_21203_new_n4101_), .B(w_mem_inst__abc_21203_new_n4099_), .Y(w_mem_inst__abc_21203_new_n4102_));
OR2X2 OR2X2_289 ( .A(_abc_15497_new_n1580_), .B(_abc_15497_new_n1575_), .Y(_abc_15497_new_n1588_));
OR2X2 OR2X2_2890 ( .A(w_mem_inst__abc_21203_new_n4102_), .B(w_mem_inst__abc_21203_new_n4098_), .Y(w_mem_inst__0w_mem_12__31_0__29_));
OR2X2 OR2X2_2891 ( .A(w_mem_inst__abc_21203_new_n4107_), .B(w_mem_inst__abc_21203_new_n4105_), .Y(w_mem_inst__abc_21203_new_n4108_));
OR2X2 OR2X2_2892 ( .A(w_mem_inst__abc_21203_new_n4108_), .B(w_mem_inst__abc_21203_new_n4104_), .Y(w_mem_inst__0w_mem_12__31_0__30_));
OR2X2 OR2X2_2893 ( .A(w_mem_inst__abc_21203_new_n4113_), .B(w_mem_inst__abc_21203_new_n4111_), .Y(w_mem_inst__abc_21203_new_n4114_));
OR2X2 OR2X2_2894 ( .A(w_mem_inst__abc_21203_new_n4114_), .B(w_mem_inst__abc_21203_new_n4110_), .Y(w_mem_inst__0w_mem_12__31_0__31_));
OR2X2 OR2X2_2895 ( .A(w_mem_inst__abc_21203_new_n4119_), .B(w_mem_inst__abc_21203_new_n4117_), .Y(w_mem_inst__abc_21203_new_n4120_));
OR2X2 OR2X2_2896 ( .A(w_mem_inst__abc_21203_new_n4120_), .B(w_mem_inst__abc_21203_new_n4116_), .Y(w_mem_inst__0w_mem_11__31_0__0_));
OR2X2 OR2X2_2897 ( .A(w_mem_inst__abc_21203_new_n4125_), .B(w_mem_inst__abc_21203_new_n4123_), .Y(w_mem_inst__abc_21203_new_n4126_));
OR2X2 OR2X2_2898 ( .A(w_mem_inst__abc_21203_new_n4126_), .B(w_mem_inst__abc_21203_new_n4122_), .Y(w_mem_inst__0w_mem_11__31_0__1_));
OR2X2 OR2X2_2899 ( .A(w_mem_inst__abc_21203_new_n4131_), .B(w_mem_inst__abc_21203_new_n4129_), .Y(w_mem_inst__abc_21203_new_n4132_));
OR2X2 OR2X2_29 ( .A(c_reg_5_), .B(\digest[69] ), .Y(_abc_15497_new_n813_));
OR2X2 OR2X2_290 ( .A(\digest[37] ), .B(d_reg_5_), .Y(_abc_15497_new_n1589_));
OR2X2 OR2X2_2900 ( .A(w_mem_inst__abc_21203_new_n4132_), .B(w_mem_inst__abc_21203_new_n4128_), .Y(w_mem_inst__0w_mem_11__31_0__2_));
OR2X2 OR2X2_2901 ( .A(w_mem_inst__abc_21203_new_n4137_), .B(w_mem_inst__abc_21203_new_n4135_), .Y(w_mem_inst__abc_21203_new_n4138_));
OR2X2 OR2X2_2902 ( .A(w_mem_inst__abc_21203_new_n4138_), .B(w_mem_inst__abc_21203_new_n4134_), .Y(w_mem_inst__0w_mem_11__31_0__3_));
OR2X2 OR2X2_2903 ( .A(w_mem_inst__abc_21203_new_n4143_), .B(w_mem_inst__abc_21203_new_n4141_), .Y(w_mem_inst__abc_21203_new_n4144_));
OR2X2 OR2X2_2904 ( .A(w_mem_inst__abc_21203_new_n4144_), .B(w_mem_inst__abc_21203_new_n4140_), .Y(w_mem_inst__0w_mem_11__31_0__4_));
OR2X2 OR2X2_2905 ( .A(w_mem_inst__abc_21203_new_n4149_), .B(w_mem_inst__abc_21203_new_n4147_), .Y(w_mem_inst__abc_21203_new_n4150_));
OR2X2 OR2X2_2906 ( .A(w_mem_inst__abc_21203_new_n4150_), .B(w_mem_inst__abc_21203_new_n4146_), .Y(w_mem_inst__0w_mem_11__31_0__5_));
OR2X2 OR2X2_2907 ( .A(w_mem_inst__abc_21203_new_n4155_), .B(w_mem_inst__abc_21203_new_n4153_), .Y(w_mem_inst__abc_21203_new_n4156_));
OR2X2 OR2X2_2908 ( .A(w_mem_inst__abc_21203_new_n4156_), .B(w_mem_inst__abc_21203_new_n4152_), .Y(w_mem_inst__0w_mem_11__31_0__6_));
OR2X2 OR2X2_2909 ( .A(w_mem_inst__abc_21203_new_n4161_), .B(w_mem_inst__abc_21203_new_n4159_), .Y(w_mem_inst__abc_21203_new_n4162_));
OR2X2 OR2X2_291 ( .A(_abc_15497_new_n1588_), .B(_abc_15497_new_n1592_), .Y(_abc_15497_new_n1593_));
OR2X2 OR2X2_2910 ( .A(w_mem_inst__abc_21203_new_n4162_), .B(w_mem_inst__abc_21203_new_n4158_), .Y(w_mem_inst__0w_mem_11__31_0__7_));
OR2X2 OR2X2_2911 ( .A(w_mem_inst__abc_21203_new_n4167_), .B(w_mem_inst__abc_21203_new_n4165_), .Y(w_mem_inst__abc_21203_new_n4168_));
OR2X2 OR2X2_2912 ( .A(w_mem_inst__abc_21203_new_n4168_), .B(w_mem_inst__abc_21203_new_n4164_), .Y(w_mem_inst__0w_mem_11__31_0__8_));
OR2X2 OR2X2_2913 ( .A(w_mem_inst__abc_21203_new_n4173_), .B(w_mem_inst__abc_21203_new_n4171_), .Y(w_mem_inst__abc_21203_new_n4174_));
OR2X2 OR2X2_2914 ( .A(w_mem_inst__abc_21203_new_n4174_), .B(w_mem_inst__abc_21203_new_n4170_), .Y(w_mem_inst__0w_mem_11__31_0__9_));
OR2X2 OR2X2_2915 ( .A(w_mem_inst__abc_21203_new_n4179_), .B(w_mem_inst__abc_21203_new_n4177_), .Y(w_mem_inst__abc_21203_new_n4180_));
OR2X2 OR2X2_2916 ( .A(w_mem_inst__abc_21203_new_n4180_), .B(w_mem_inst__abc_21203_new_n4176_), .Y(w_mem_inst__0w_mem_11__31_0__10_));
OR2X2 OR2X2_2917 ( .A(w_mem_inst__abc_21203_new_n4185_), .B(w_mem_inst__abc_21203_new_n4183_), .Y(w_mem_inst__abc_21203_new_n4186_));
OR2X2 OR2X2_2918 ( .A(w_mem_inst__abc_21203_new_n4186_), .B(w_mem_inst__abc_21203_new_n4182_), .Y(w_mem_inst__0w_mem_11__31_0__11_));
OR2X2 OR2X2_2919 ( .A(w_mem_inst__abc_21203_new_n4191_), .B(w_mem_inst__abc_21203_new_n4189_), .Y(w_mem_inst__abc_21203_new_n4192_));
OR2X2 OR2X2_292 ( .A(_abc_15497_new_n699_), .B(\digest[37] ), .Y(_abc_15497_new_n1598_));
OR2X2 OR2X2_2920 ( .A(w_mem_inst__abc_21203_new_n4192_), .B(w_mem_inst__abc_21203_new_n4188_), .Y(w_mem_inst__0w_mem_11__31_0__12_));
OR2X2 OR2X2_2921 ( .A(w_mem_inst__abc_21203_new_n4197_), .B(w_mem_inst__abc_21203_new_n4195_), .Y(w_mem_inst__abc_21203_new_n4198_));
OR2X2 OR2X2_2922 ( .A(w_mem_inst__abc_21203_new_n4198_), .B(w_mem_inst__abc_21203_new_n4194_), .Y(w_mem_inst__0w_mem_11__31_0__13_));
OR2X2 OR2X2_2923 ( .A(w_mem_inst__abc_21203_new_n4203_), .B(w_mem_inst__abc_21203_new_n4201_), .Y(w_mem_inst__abc_21203_new_n4204_));
OR2X2 OR2X2_2924 ( .A(w_mem_inst__abc_21203_new_n4204_), .B(w_mem_inst__abc_21203_new_n4200_), .Y(w_mem_inst__0w_mem_11__31_0__14_));
OR2X2 OR2X2_2925 ( .A(w_mem_inst__abc_21203_new_n4209_), .B(w_mem_inst__abc_21203_new_n4207_), .Y(w_mem_inst__abc_21203_new_n4210_));
OR2X2 OR2X2_2926 ( .A(w_mem_inst__abc_21203_new_n4210_), .B(w_mem_inst__abc_21203_new_n4206_), .Y(w_mem_inst__0w_mem_11__31_0__15_));
OR2X2 OR2X2_2927 ( .A(w_mem_inst__abc_21203_new_n4215_), .B(w_mem_inst__abc_21203_new_n4213_), .Y(w_mem_inst__abc_21203_new_n4216_));
OR2X2 OR2X2_2928 ( .A(w_mem_inst__abc_21203_new_n4216_), .B(w_mem_inst__abc_21203_new_n4212_), .Y(w_mem_inst__0w_mem_11__31_0__16_));
OR2X2 OR2X2_2929 ( .A(w_mem_inst__abc_21203_new_n4221_), .B(w_mem_inst__abc_21203_new_n4219_), .Y(w_mem_inst__abc_21203_new_n4222_));
OR2X2 OR2X2_293 ( .A(_abc_15497_new_n1597_), .B(_abc_15497_new_n1599_), .Y(_0H3_reg_31_0__5_));
OR2X2 OR2X2_2930 ( .A(w_mem_inst__abc_21203_new_n4222_), .B(w_mem_inst__abc_21203_new_n4218_), .Y(w_mem_inst__0w_mem_11__31_0__17_));
OR2X2 OR2X2_2931 ( .A(w_mem_inst__abc_21203_new_n4227_), .B(w_mem_inst__abc_21203_new_n4225_), .Y(w_mem_inst__abc_21203_new_n4228_));
OR2X2 OR2X2_2932 ( .A(w_mem_inst__abc_21203_new_n4228_), .B(w_mem_inst__abc_21203_new_n4224_), .Y(w_mem_inst__0w_mem_11__31_0__18_));
OR2X2 OR2X2_2933 ( .A(w_mem_inst__abc_21203_new_n4233_), .B(w_mem_inst__abc_21203_new_n4231_), .Y(w_mem_inst__abc_21203_new_n4234_));
OR2X2 OR2X2_2934 ( .A(w_mem_inst__abc_21203_new_n4234_), .B(w_mem_inst__abc_21203_new_n4230_), .Y(w_mem_inst__0w_mem_11__31_0__19_));
OR2X2 OR2X2_2935 ( .A(w_mem_inst__abc_21203_new_n4239_), .B(w_mem_inst__abc_21203_new_n4237_), .Y(w_mem_inst__abc_21203_new_n4240_));
OR2X2 OR2X2_2936 ( .A(w_mem_inst__abc_21203_new_n4240_), .B(w_mem_inst__abc_21203_new_n4236_), .Y(w_mem_inst__0w_mem_11__31_0__20_));
OR2X2 OR2X2_2937 ( .A(w_mem_inst__abc_21203_new_n4245_), .B(w_mem_inst__abc_21203_new_n4243_), .Y(w_mem_inst__abc_21203_new_n4246_));
OR2X2 OR2X2_2938 ( .A(w_mem_inst__abc_21203_new_n4246_), .B(w_mem_inst__abc_21203_new_n4242_), .Y(w_mem_inst__0w_mem_11__31_0__21_));
OR2X2 OR2X2_2939 ( .A(w_mem_inst__abc_21203_new_n4251_), .B(w_mem_inst__abc_21203_new_n4249_), .Y(w_mem_inst__abc_21203_new_n4252_));
OR2X2 OR2X2_294 ( .A(_abc_15497_new_n1594_), .B(_abc_15497_new_n1590_), .Y(_abc_15497_new_n1601_));
OR2X2 OR2X2_2940 ( .A(w_mem_inst__abc_21203_new_n4252_), .B(w_mem_inst__abc_21203_new_n4248_), .Y(w_mem_inst__0w_mem_11__31_0__22_));
OR2X2 OR2X2_2941 ( .A(w_mem_inst__abc_21203_new_n4257_), .B(w_mem_inst__abc_21203_new_n4255_), .Y(w_mem_inst__abc_21203_new_n4258_));
OR2X2 OR2X2_2942 ( .A(w_mem_inst__abc_21203_new_n4258_), .B(w_mem_inst__abc_21203_new_n4254_), .Y(w_mem_inst__0w_mem_11__31_0__23_));
OR2X2 OR2X2_2943 ( .A(w_mem_inst__abc_21203_new_n4263_), .B(w_mem_inst__abc_21203_new_n4261_), .Y(w_mem_inst__abc_21203_new_n4264_));
OR2X2 OR2X2_2944 ( .A(w_mem_inst__abc_21203_new_n4264_), .B(w_mem_inst__abc_21203_new_n4260_), .Y(w_mem_inst__0w_mem_11__31_0__24_));
OR2X2 OR2X2_2945 ( .A(w_mem_inst__abc_21203_new_n4269_), .B(w_mem_inst__abc_21203_new_n4267_), .Y(w_mem_inst__abc_21203_new_n4270_));
OR2X2 OR2X2_2946 ( .A(w_mem_inst__abc_21203_new_n4270_), .B(w_mem_inst__abc_21203_new_n4266_), .Y(w_mem_inst__0w_mem_11__31_0__25_));
OR2X2 OR2X2_2947 ( .A(w_mem_inst__abc_21203_new_n4275_), .B(w_mem_inst__abc_21203_new_n4273_), .Y(w_mem_inst__abc_21203_new_n4276_));
OR2X2 OR2X2_2948 ( .A(w_mem_inst__abc_21203_new_n4276_), .B(w_mem_inst__abc_21203_new_n4272_), .Y(w_mem_inst__0w_mem_11__31_0__26_));
OR2X2 OR2X2_2949 ( .A(w_mem_inst__abc_21203_new_n4281_), .B(w_mem_inst__abc_21203_new_n4279_), .Y(w_mem_inst__abc_21203_new_n4282_));
OR2X2 OR2X2_295 ( .A(\digest[38] ), .B(d_reg_6_), .Y(_abc_15497_new_n1602_));
OR2X2 OR2X2_2950 ( .A(w_mem_inst__abc_21203_new_n4282_), .B(w_mem_inst__abc_21203_new_n4278_), .Y(w_mem_inst__0w_mem_11__31_0__27_));
OR2X2 OR2X2_2951 ( .A(w_mem_inst__abc_21203_new_n4287_), .B(w_mem_inst__abc_21203_new_n4285_), .Y(w_mem_inst__abc_21203_new_n4288_));
OR2X2 OR2X2_2952 ( .A(w_mem_inst__abc_21203_new_n4288_), .B(w_mem_inst__abc_21203_new_n4284_), .Y(w_mem_inst__0w_mem_11__31_0__28_));
OR2X2 OR2X2_2953 ( .A(w_mem_inst__abc_21203_new_n4293_), .B(w_mem_inst__abc_21203_new_n4291_), .Y(w_mem_inst__abc_21203_new_n4294_));
OR2X2 OR2X2_2954 ( .A(w_mem_inst__abc_21203_new_n4294_), .B(w_mem_inst__abc_21203_new_n4290_), .Y(w_mem_inst__0w_mem_11__31_0__29_));
OR2X2 OR2X2_2955 ( .A(w_mem_inst__abc_21203_new_n4299_), .B(w_mem_inst__abc_21203_new_n4297_), .Y(w_mem_inst__abc_21203_new_n4300_));
OR2X2 OR2X2_2956 ( .A(w_mem_inst__abc_21203_new_n4300_), .B(w_mem_inst__abc_21203_new_n4296_), .Y(w_mem_inst__0w_mem_11__31_0__30_));
OR2X2 OR2X2_2957 ( .A(w_mem_inst__abc_21203_new_n4305_), .B(w_mem_inst__abc_21203_new_n4303_), .Y(w_mem_inst__abc_21203_new_n4306_));
OR2X2 OR2X2_2958 ( .A(w_mem_inst__abc_21203_new_n4306_), .B(w_mem_inst__abc_21203_new_n4302_), .Y(w_mem_inst__0w_mem_11__31_0__31_));
OR2X2 OR2X2_2959 ( .A(w_mem_inst__abc_21203_new_n4311_), .B(w_mem_inst__abc_21203_new_n4309_), .Y(w_mem_inst__abc_21203_new_n4312_));
OR2X2 OR2X2_296 ( .A(_abc_15497_new_n1601_), .B(_abc_15497_new_n1605_), .Y(_abc_15497_new_n1606_));
OR2X2 OR2X2_2960 ( .A(w_mem_inst__abc_21203_new_n4312_), .B(w_mem_inst__abc_21203_new_n4308_), .Y(w_mem_inst__0w_mem_7__31_0__0_));
OR2X2 OR2X2_2961 ( .A(w_mem_inst__abc_21203_new_n4317_), .B(w_mem_inst__abc_21203_new_n4315_), .Y(w_mem_inst__abc_21203_new_n4318_));
OR2X2 OR2X2_2962 ( .A(w_mem_inst__abc_21203_new_n4318_), .B(w_mem_inst__abc_21203_new_n4314_), .Y(w_mem_inst__0w_mem_7__31_0__1_));
OR2X2 OR2X2_2963 ( .A(w_mem_inst__abc_21203_new_n4323_), .B(w_mem_inst__abc_21203_new_n4321_), .Y(w_mem_inst__abc_21203_new_n4324_));
OR2X2 OR2X2_2964 ( .A(w_mem_inst__abc_21203_new_n4324_), .B(w_mem_inst__abc_21203_new_n4320_), .Y(w_mem_inst__0w_mem_7__31_0__2_));
OR2X2 OR2X2_2965 ( .A(w_mem_inst__abc_21203_new_n4329_), .B(w_mem_inst__abc_21203_new_n4327_), .Y(w_mem_inst__abc_21203_new_n4330_));
OR2X2 OR2X2_2966 ( .A(w_mem_inst__abc_21203_new_n4330_), .B(w_mem_inst__abc_21203_new_n4326_), .Y(w_mem_inst__0w_mem_7__31_0__3_));
OR2X2 OR2X2_2967 ( .A(w_mem_inst__abc_21203_new_n4335_), .B(w_mem_inst__abc_21203_new_n4333_), .Y(w_mem_inst__abc_21203_new_n4336_));
OR2X2 OR2X2_2968 ( .A(w_mem_inst__abc_21203_new_n4336_), .B(w_mem_inst__abc_21203_new_n4332_), .Y(w_mem_inst__0w_mem_7__31_0__4_));
OR2X2 OR2X2_2969 ( .A(w_mem_inst__abc_21203_new_n4341_), .B(w_mem_inst__abc_21203_new_n4339_), .Y(w_mem_inst__abc_21203_new_n4342_));
OR2X2 OR2X2_297 ( .A(_abc_15497_new_n699_), .B(\digest[38] ), .Y(_abc_15497_new_n1611_));
OR2X2 OR2X2_2970 ( .A(w_mem_inst__abc_21203_new_n4342_), .B(w_mem_inst__abc_21203_new_n4338_), .Y(w_mem_inst__0w_mem_7__31_0__5_));
OR2X2 OR2X2_2971 ( .A(w_mem_inst__abc_21203_new_n4347_), .B(w_mem_inst__abc_21203_new_n4345_), .Y(w_mem_inst__abc_21203_new_n4348_));
OR2X2 OR2X2_2972 ( .A(w_mem_inst__abc_21203_new_n4348_), .B(w_mem_inst__abc_21203_new_n4344_), .Y(w_mem_inst__0w_mem_7__31_0__6_));
OR2X2 OR2X2_2973 ( .A(w_mem_inst__abc_21203_new_n4353_), .B(w_mem_inst__abc_21203_new_n4351_), .Y(w_mem_inst__abc_21203_new_n4354_));
OR2X2 OR2X2_2974 ( .A(w_mem_inst__abc_21203_new_n4354_), .B(w_mem_inst__abc_21203_new_n4350_), .Y(w_mem_inst__0w_mem_7__31_0__7_));
OR2X2 OR2X2_2975 ( .A(w_mem_inst__abc_21203_new_n4359_), .B(w_mem_inst__abc_21203_new_n4357_), .Y(w_mem_inst__abc_21203_new_n4360_));
OR2X2 OR2X2_2976 ( .A(w_mem_inst__abc_21203_new_n4360_), .B(w_mem_inst__abc_21203_new_n4356_), .Y(w_mem_inst__0w_mem_7__31_0__8_));
OR2X2 OR2X2_2977 ( .A(w_mem_inst__abc_21203_new_n4365_), .B(w_mem_inst__abc_21203_new_n4363_), .Y(w_mem_inst__abc_21203_new_n4366_));
OR2X2 OR2X2_2978 ( .A(w_mem_inst__abc_21203_new_n4366_), .B(w_mem_inst__abc_21203_new_n4362_), .Y(w_mem_inst__0w_mem_7__31_0__9_));
OR2X2 OR2X2_2979 ( .A(w_mem_inst__abc_21203_new_n4371_), .B(w_mem_inst__abc_21203_new_n4369_), .Y(w_mem_inst__abc_21203_new_n4372_));
OR2X2 OR2X2_298 ( .A(_abc_15497_new_n1610_), .B(_abc_15497_new_n1612_), .Y(_0H3_reg_31_0__6_));
OR2X2 OR2X2_2980 ( .A(w_mem_inst__abc_21203_new_n4372_), .B(w_mem_inst__abc_21203_new_n4368_), .Y(w_mem_inst__0w_mem_7__31_0__10_));
OR2X2 OR2X2_2981 ( .A(w_mem_inst__abc_21203_new_n4377_), .B(w_mem_inst__abc_21203_new_n4375_), .Y(w_mem_inst__abc_21203_new_n4378_));
OR2X2 OR2X2_2982 ( .A(w_mem_inst__abc_21203_new_n4378_), .B(w_mem_inst__abc_21203_new_n4374_), .Y(w_mem_inst__0w_mem_7__31_0__11_));
OR2X2 OR2X2_2983 ( .A(w_mem_inst__abc_21203_new_n4383_), .B(w_mem_inst__abc_21203_new_n4381_), .Y(w_mem_inst__abc_21203_new_n4384_));
OR2X2 OR2X2_2984 ( .A(w_mem_inst__abc_21203_new_n4384_), .B(w_mem_inst__abc_21203_new_n4380_), .Y(w_mem_inst__0w_mem_7__31_0__12_));
OR2X2 OR2X2_2985 ( .A(w_mem_inst__abc_21203_new_n4389_), .B(w_mem_inst__abc_21203_new_n4387_), .Y(w_mem_inst__abc_21203_new_n4390_));
OR2X2 OR2X2_2986 ( .A(w_mem_inst__abc_21203_new_n4390_), .B(w_mem_inst__abc_21203_new_n4386_), .Y(w_mem_inst__0w_mem_7__31_0__13_));
OR2X2 OR2X2_2987 ( .A(w_mem_inst__abc_21203_new_n4395_), .B(w_mem_inst__abc_21203_new_n4393_), .Y(w_mem_inst__abc_21203_new_n4396_));
OR2X2 OR2X2_2988 ( .A(w_mem_inst__abc_21203_new_n4396_), .B(w_mem_inst__abc_21203_new_n4392_), .Y(w_mem_inst__0w_mem_7__31_0__14_));
OR2X2 OR2X2_2989 ( .A(w_mem_inst__abc_21203_new_n4401_), .B(w_mem_inst__abc_21203_new_n4399_), .Y(w_mem_inst__abc_21203_new_n4402_));
OR2X2 OR2X2_299 ( .A(\digest[39] ), .B(d_reg_7_), .Y(_abc_15497_new_n1615_));
OR2X2 OR2X2_2990 ( .A(w_mem_inst__abc_21203_new_n4402_), .B(w_mem_inst__abc_21203_new_n4398_), .Y(w_mem_inst__0w_mem_7__31_0__15_));
OR2X2 OR2X2_2991 ( .A(w_mem_inst__abc_21203_new_n4407_), .B(w_mem_inst__abc_21203_new_n4405_), .Y(w_mem_inst__abc_21203_new_n4408_));
OR2X2 OR2X2_2992 ( .A(w_mem_inst__abc_21203_new_n4408_), .B(w_mem_inst__abc_21203_new_n4404_), .Y(w_mem_inst__0w_mem_7__31_0__16_));
OR2X2 OR2X2_2993 ( .A(w_mem_inst__abc_21203_new_n4413_), .B(w_mem_inst__abc_21203_new_n4411_), .Y(w_mem_inst__abc_21203_new_n4414_));
OR2X2 OR2X2_2994 ( .A(w_mem_inst__abc_21203_new_n4414_), .B(w_mem_inst__abc_21203_new_n4410_), .Y(w_mem_inst__0w_mem_7__31_0__17_));
OR2X2 OR2X2_2995 ( .A(w_mem_inst__abc_21203_new_n4419_), .B(w_mem_inst__abc_21203_new_n4417_), .Y(w_mem_inst__abc_21203_new_n4420_));
OR2X2 OR2X2_2996 ( .A(w_mem_inst__abc_21203_new_n4420_), .B(w_mem_inst__abc_21203_new_n4416_), .Y(w_mem_inst__0w_mem_7__31_0__18_));
OR2X2 OR2X2_2997 ( .A(w_mem_inst__abc_21203_new_n4425_), .B(w_mem_inst__abc_21203_new_n4423_), .Y(w_mem_inst__abc_21203_new_n4426_));
OR2X2 OR2X2_2998 ( .A(w_mem_inst__abc_21203_new_n4426_), .B(w_mem_inst__abc_21203_new_n4422_), .Y(w_mem_inst__0w_mem_7__31_0__19_));
OR2X2 OR2X2_2999 ( .A(w_mem_inst__abc_21203_new_n4431_), .B(w_mem_inst__abc_21203_new_n4429_), .Y(w_mem_inst__abc_21203_new_n4432_));
OR2X2 OR2X2_3 ( .A(c_reg_21_), .B(\digest[85] ), .Y(_abc_15497_new_n717_));
OR2X2 OR2X2_30 ( .A(c_reg_3_), .B(\digest[67] ), .Y(_abc_15497_new_n816_));
OR2X2 OR2X2_300 ( .A(_abc_15497_new_n1607_), .B(_abc_15497_new_n1603_), .Y(_abc_15497_new_n1619_));
OR2X2 OR2X2_3000 ( .A(w_mem_inst__abc_21203_new_n4432_), .B(w_mem_inst__abc_21203_new_n4428_), .Y(w_mem_inst__0w_mem_7__31_0__20_));
OR2X2 OR2X2_3001 ( .A(w_mem_inst__abc_21203_new_n4437_), .B(w_mem_inst__abc_21203_new_n4435_), .Y(w_mem_inst__abc_21203_new_n4438_));
OR2X2 OR2X2_3002 ( .A(w_mem_inst__abc_21203_new_n4438_), .B(w_mem_inst__abc_21203_new_n4434_), .Y(w_mem_inst__0w_mem_7__31_0__21_));
OR2X2 OR2X2_3003 ( .A(w_mem_inst__abc_21203_new_n4443_), .B(w_mem_inst__abc_21203_new_n4441_), .Y(w_mem_inst__abc_21203_new_n4444_));
OR2X2 OR2X2_3004 ( .A(w_mem_inst__abc_21203_new_n4444_), .B(w_mem_inst__abc_21203_new_n4440_), .Y(w_mem_inst__0w_mem_7__31_0__22_));
OR2X2 OR2X2_3005 ( .A(w_mem_inst__abc_21203_new_n4449_), .B(w_mem_inst__abc_21203_new_n4447_), .Y(w_mem_inst__abc_21203_new_n4450_));
OR2X2 OR2X2_3006 ( .A(w_mem_inst__abc_21203_new_n4450_), .B(w_mem_inst__abc_21203_new_n4446_), .Y(w_mem_inst__0w_mem_7__31_0__23_));
OR2X2 OR2X2_3007 ( .A(w_mem_inst__abc_21203_new_n4455_), .B(w_mem_inst__abc_21203_new_n4453_), .Y(w_mem_inst__abc_21203_new_n4456_));
OR2X2 OR2X2_3008 ( .A(w_mem_inst__abc_21203_new_n4456_), .B(w_mem_inst__abc_21203_new_n4452_), .Y(w_mem_inst__0w_mem_7__31_0__24_));
OR2X2 OR2X2_3009 ( .A(w_mem_inst__abc_21203_new_n4461_), .B(w_mem_inst__abc_21203_new_n4459_), .Y(w_mem_inst__abc_21203_new_n4462_));
OR2X2 OR2X2_301 ( .A(_abc_15497_new_n1619_), .B(_abc_15497_new_n1618_), .Y(_abc_15497_new_n1620_));
OR2X2 OR2X2_3010 ( .A(w_mem_inst__abc_21203_new_n4462_), .B(w_mem_inst__abc_21203_new_n4458_), .Y(w_mem_inst__0w_mem_7__31_0__25_));
OR2X2 OR2X2_3011 ( .A(w_mem_inst__abc_21203_new_n4467_), .B(w_mem_inst__abc_21203_new_n4465_), .Y(w_mem_inst__abc_21203_new_n4468_));
OR2X2 OR2X2_3012 ( .A(w_mem_inst__abc_21203_new_n4468_), .B(w_mem_inst__abc_21203_new_n4464_), .Y(w_mem_inst__0w_mem_7__31_0__26_));
OR2X2 OR2X2_3013 ( .A(w_mem_inst__abc_21203_new_n4473_), .B(w_mem_inst__abc_21203_new_n4471_), .Y(w_mem_inst__abc_21203_new_n4474_));
OR2X2 OR2X2_3014 ( .A(w_mem_inst__abc_21203_new_n4474_), .B(w_mem_inst__abc_21203_new_n4470_), .Y(w_mem_inst__0w_mem_7__31_0__27_));
OR2X2 OR2X2_3015 ( .A(w_mem_inst__abc_21203_new_n4479_), .B(w_mem_inst__abc_21203_new_n4477_), .Y(w_mem_inst__abc_21203_new_n4480_));
OR2X2 OR2X2_3016 ( .A(w_mem_inst__abc_21203_new_n4480_), .B(w_mem_inst__abc_21203_new_n4476_), .Y(w_mem_inst__0w_mem_7__31_0__28_));
OR2X2 OR2X2_3017 ( .A(w_mem_inst__abc_21203_new_n4485_), .B(w_mem_inst__abc_21203_new_n4483_), .Y(w_mem_inst__abc_21203_new_n4486_));
OR2X2 OR2X2_3018 ( .A(w_mem_inst__abc_21203_new_n4486_), .B(w_mem_inst__abc_21203_new_n4482_), .Y(w_mem_inst__0w_mem_7__31_0__29_));
OR2X2 OR2X2_3019 ( .A(w_mem_inst__abc_21203_new_n4491_), .B(w_mem_inst__abc_21203_new_n4489_), .Y(w_mem_inst__abc_21203_new_n4492_));
OR2X2 OR2X2_302 ( .A(_abc_15497_new_n1624_), .B(_abc_15497_new_n1614_), .Y(_0H3_reg_31_0__7_));
OR2X2 OR2X2_3020 ( .A(w_mem_inst__abc_21203_new_n4492_), .B(w_mem_inst__abc_21203_new_n4488_), .Y(w_mem_inst__0w_mem_7__31_0__30_));
OR2X2 OR2X2_3021 ( .A(w_mem_inst__abc_21203_new_n4497_), .B(w_mem_inst__abc_21203_new_n4495_), .Y(w_mem_inst__abc_21203_new_n4498_));
OR2X2 OR2X2_3022 ( .A(w_mem_inst__abc_21203_new_n4498_), .B(w_mem_inst__abc_21203_new_n4494_), .Y(w_mem_inst__0w_mem_7__31_0__31_));
OR2X2 OR2X2_3023 ( .A(w_mem_inst__abc_21203_new_n4503_), .B(w_mem_inst__abc_21203_new_n4501_), .Y(w_mem_inst__abc_21203_new_n4504_));
OR2X2 OR2X2_3024 ( .A(w_mem_inst__abc_21203_new_n4504_), .B(w_mem_inst__abc_21203_new_n4500_), .Y(w_mem_inst__0w_mem_9__31_0__0_));
OR2X2 OR2X2_3025 ( .A(w_mem_inst__abc_21203_new_n4509_), .B(w_mem_inst__abc_21203_new_n4507_), .Y(w_mem_inst__abc_21203_new_n4510_));
OR2X2 OR2X2_3026 ( .A(w_mem_inst__abc_21203_new_n4510_), .B(w_mem_inst__abc_21203_new_n4506_), .Y(w_mem_inst__0w_mem_9__31_0__1_));
OR2X2 OR2X2_3027 ( .A(w_mem_inst__abc_21203_new_n4515_), .B(w_mem_inst__abc_21203_new_n4513_), .Y(w_mem_inst__abc_21203_new_n4516_));
OR2X2 OR2X2_3028 ( .A(w_mem_inst__abc_21203_new_n4516_), .B(w_mem_inst__abc_21203_new_n4512_), .Y(w_mem_inst__0w_mem_9__31_0__2_));
OR2X2 OR2X2_3029 ( .A(w_mem_inst__abc_21203_new_n4521_), .B(w_mem_inst__abc_21203_new_n4519_), .Y(w_mem_inst__abc_21203_new_n4522_));
OR2X2 OR2X2_303 ( .A(_abc_15497_new_n1621_), .B(_abc_15497_new_n1616_), .Y(_abc_15497_new_n1627_));
OR2X2 OR2X2_3030 ( .A(w_mem_inst__abc_21203_new_n4522_), .B(w_mem_inst__abc_21203_new_n4518_), .Y(w_mem_inst__0w_mem_9__31_0__3_));
OR2X2 OR2X2_3031 ( .A(w_mem_inst__abc_21203_new_n4527_), .B(w_mem_inst__abc_21203_new_n4525_), .Y(w_mem_inst__abc_21203_new_n4528_));
OR2X2 OR2X2_3032 ( .A(w_mem_inst__abc_21203_new_n4528_), .B(w_mem_inst__abc_21203_new_n4524_), .Y(w_mem_inst__0w_mem_9__31_0__4_));
OR2X2 OR2X2_3033 ( .A(w_mem_inst__abc_21203_new_n4533_), .B(w_mem_inst__abc_21203_new_n4531_), .Y(w_mem_inst__abc_21203_new_n4534_));
OR2X2 OR2X2_3034 ( .A(w_mem_inst__abc_21203_new_n4534_), .B(w_mem_inst__abc_21203_new_n4530_), .Y(w_mem_inst__0w_mem_9__31_0__5_));
OR2X2 OR2X2_3035 ( .A(w_mem_inst__abc_21203_new_n4539_), .B(w_mem_inst__abc_21203_new_n4537_), .Y(w_mem_inst__abc_21203_new_n4540_));
OR2X2 OR2X2_3036 ( .A(w_mem_inst__abc_21203_new_n4540_), .B(w_mem_inst__abc_21203_new_n4536_), .Y(w_mem_inst__0w_mem_9__31_0__6_));
OR2X2 OR2X2_3037 ( .A(w_mem_inst__abc_21203_new_n4545_), .B(w_mem_inst__abc_21203_new_n4543_), .Y(w_mem_inst__abc_21203_new_n4546_));
OR2X2 OR2X2_3038 ( .A(w_mem_inst__abc_21203_new_n4546_), .B(w_mem_inst__abc_21203_new_n4542_), .Y(w_mem_inst__0w_mem_9__31_0__7_));
OR2X2 OR2X2_3039 ( .A(w_mem_inst__abc_21203_new_n4551_), .B(w_mem_inst__abc_21203_new_n4549_), .Y(w_mem_inst__abc_21203_new_n4552_));
OR2X2 OR2X2_304 ( .A(\digest[40] ), .B(d_reg_8_), .Y(_abc_15497_new_n1628_));
OR2X2 OR2X2_3040 ( .A(w_mem_inst__abc_21203_new_n4552_), .B(w_mem_inst__abc_21203_new_n4548_), .Y(w_mem_inst__0w_mem_9__31_0__8_));
OR2X2 OR2X2_3041 ( .A(w_mem_inst__abc_21203_new_n4557_), .B(w_mem_inst__abc_21203_new_n4555_), .Y(w_mem_inst__abc_21203_new_n4558_));
OR2X2 OR2X2_3042 ( .A(w_mem_inst__abc_21203_new_n4558_), .B(w_mem_inst__abc_21203_new_n4554_), .Y(w_mem_inst__0w_mem_9__31_0__9_));
OR2X2 OR2X2_3043 ( .A(w_mem_inst__abc_21203_new_n4563_), .B(w_mem_inst__abc_21203_new_n4561_), .Y(w_mem_inst__abc_21203_new_n4564_));
OR2X2 OR2X2_3044 ( .A(w_mem_inst__abc_21203_new_n4564_), .B(w_mem_inst__abc_21203_new_n4560_), .Y(w_mem_inst__0w_mem_9__31_0__10_));
OR2X2 OR2X2_3045 ( .A(w_mem_inst__abc_21203_new_n4569_), .B(w_mem_inst__abc_21203_new_n4567_), .Y(w_mem_inst__abc_21203_new_n4570_));
OR2X2 OR2X2_3046 ( .A(w_mem_inst__abc_21203_new_n4570_), .B(w_mem_inst__abc_21203_new_n4566_), .Y(w_mem_inst__0w_mem_9__31_0__11_));
OR2X2 OR2X2_3047 ( .A(w_mem_inst__abc_21203_new_n4575_), .B(w_mem_inst__abc_21203_new_n4573_), .Y(w_mem_inst__abc_21203_new_n4576_));
OR2X2 OR2X2_3048 ( .A(w_mem_inst__abc_21203_new_n4576_), .B(w_mem_inst__abc_21203_new_n4572_), .Y(w_mem_inst__0w_mem_9__31_0__12_));
OR2X2 OR2X2_3049 ( .A(w_mem_inst__abc_21203_new_n4581_), .B(w_mem_inst__abc_21203_new_n4579_), .Y(w_mem_inst__abc_21203_new_n4582_));
OR2X2 OR2X2_305 ( .A(_abc_15497_new_n1627_), .B(_abc_15497_new_n1631_), .Y(_abc_15497_new_n1632_));
OR2X2 OR2X2_3050 ( .A(w_mem_inst__abc_21203_new_n4582_), .B(w_mem_inst__abc_21203_new_n4578_), .Y(w_mem_inst__0w_mem_9__31_0__13_));
OR2X2 OR2X2_3051 ( .A(w_mem_inst__abc_21203_new_n4587_), .B(w_mem_inst__abc_21203_new_n4585_), .Y(w_mem_inst__abc_21203_new_n4588_));
OR2X2 OR2X2_3052 ( .A(w_mem_inst__abc_21203_new_n4588_), .B(w_mem_inst__abc_21203_new_n4584_), .Y(w_mem_inst__0w_mem_9__31_0__14_));
OR2X2 OR2X2_3053 ( .A(w_mem_inst__abc_21203_new_n4593_), .B(w_mem_inst__abc_21203_new_n4591_), .Y(w_mem_inst__abc_21203_new_n4594_));
OR2X2 OR2X2_3054 ( .A(w_mem_inst__abc_21203_new_n4594_), .B(w_mem_inst__abc_21203_new_n4590_), .Y(w_mem_inst__0w_mem_9__31_0__15_));
OR2X2 OR2X2_3055 ( .A(w_mem_inst__abc_21203_new_n4599_), .B(w_mem_inst__abc_21203_new_n4597_), .Y(w_mem_inst__abc_21203_new_n4600_));
OR2X2 OR2X2_3056 ( .A(w_mem_inst__abc_21203_new_n4600_), .B(w_mem_inst__abc_21203_new_n4596_), .Y(w_mem_inst__0w_mem_9__31_0__16_));
OR2X2 OR2X2_3057 ( .A(w_mem_inst__abc_21203_new_n4605_), .B(w_mem_inst__abc_21203_new_n4603_), .Y(w_mem_inst__abc_21203_new_n4606_));
OR2X2 OR2X2_3058 ( .A(w_mem_inst__abc_21203_new_n4606_), .B(w_mem_inst__abc_21203_new_n4602_), .Y(w_mem_inst__0w_mem_9__31_0__17_));
OR2X2 OR2X2_3059 ( .A(w_mem_inst__abc_21203_new_n4611_), .B(w_mem_inst__abc_21203_new_n4609_), .Y(w_mem_inst__abc_21203_new_n4612_));
OR2X2 OR2X2_306 ( .A(_abc_15497_new_n1636_), .B(_abc_15497_new_n1626_), .Y(_0H3_reg_31_0__8_));
OR2X2 OR2X2_3060 ( .A(w_mem_inst__abc_21203_new_n4612_), .B(w_mem_inst__abc_21203_new_n4608_), .Y(w_mem_inst__0w_mem_9__31_0__18_));
OR2X2 OR2X2_3061 ( .A(w_mem_inst__abc_21203_new_n4617_), .B(w_mem_inst__abc_21203_new_n4615_), .Y(w_mem_inst__abc_21203_new_n4618_));
OR2X2 OR2X2_3062 ( .A(w_mem_inst__abc_21203_new_n4618_), .B(w_mem_inst__abc_21203_new_n4614_), .Y(w_mem_inst__0w_mem_9__31_0__19_));
OR2X2 OR2X2_3063 ( .A(w_mem_inst__abc_21203_new_n4623_), .B(w_mem_inst__abc_21203_new_n4621_), .Y(w_mem_inst__abc_21203_new_n4624_));
OR2X2 OR2X2_3064 ( .A(w_mem_inst__abc_21203_new_n4624_), .B(w_mem_inst__abc_21203_new_n4620_), .Y(w_mem_inst__0w_mem_9__31_0__20_));
OR2X2 OR2X2_3065 ( .A(w_mem_inst__abc_21203_new_n4629_), .B(w_mem_inst__abc_21203_new_n4627_), .Y(w_mem_inst__abc_21203_new_n4630_));
OR2X2 OR2X2_3066 ( .A(w_mem_inst__abc_21203_new_n4630_), .B(w_mem_inst__abc_21203_new_n4626_), .Y(w_mem_inst__0w_mem_9__31_0__21_));
OR2X2 OR2X2_3067 ( .A(w_mem_inst__abc_21203_new_n4635_), .B(w_mem_inst__abc_21203_new_n4633_), .Y(w_mem_inst__abc_21203_new_n4636_));
OR2X2 OR2X2_3068 ( .A(w_mem_inst__abc_21203_new_n4636_), .B(w_mem_inst__abc_21203_new_n4632_), .Y(w_mem_inst__0w_mem_9__31_0__22_));
OR2X2 OR2X2_3069 ( .A(w_mem_inst__abc_21203_new_n4641_), .B(w_mem_inst__abc_21203_new_n4639_), .Y(w_mem_inst__abc_21203_new_n4642_));
OR2X2 OR2X2_307 ( .A(\digest[41] ), .B(d_reg_9_), .Y(_abc_15497_new_n1639_));
OR2X2 OR2X2_3070 ( .A(w_mem_inst__abc_21203_new_n4642_), .B(w_mem_inst__abc_21203_new_n4638_), .Y(w_mem_inst__0w_mem_9__31_0__23_));
OR2X2 OR2X2_3071 ( .A(w_mem_inst__abc_21203_new_n4647_), .B(w_mem_inst__abc_21203_new_n4645_), .Y(w_mem_inst__abc_21203_new_n4648_));
OR2X2 OR2X2_3072 ( .A(w_mem_inst__abc_21203_new_n4648_), .B(w_mem_inst__abc_21203_new_n4644_), .Y(w_mem_inst__0w_mem_9__31_0__24_));
OR2X2 OR2X2_3073 ( .A(w_mem_inst__abc_21203_new_n4653_), .B(w_mem_inst__abc_21203_new_n4651_), .Y(w_mem_inst__abc_21203_new_n4654_));
OR2X2 OR2X2_3074 ( .A(w_mem_inst__abc_21203_new_n4654_), .B(w_mem_inst__abc_21203_new_n4650_), .Y(w_mem_inst__0w_mem_9__31_0__25_));
OR2X2 OR2X2_3075 ( .A(w_mem_inst__abc_21203_new_n4659_), .B(w_mem_inst__abc_21203_new_n4657_), .Y(w_mem_inst__abc_21203_new_n4660_));
OR2X2 OR2X2_3076 ( .A(w_mem_inst__abc_21203_new_n4660_), .B(w_mem_inst__abc_21203_new_n4656_), .Y(w_mem_inst__0w_mem_9__31_0__26_));
OR2X2 OR2X2_3077 ( .A(w_mem_inst__abc_21203_new_n4665_), .B(w_mem_inst__abc_21203_new_n4663_), .Y(w_mem_inst__abc_21203_new_n4666_));
OR2X2 OR2X2_3078 ( .A(w_mem_inst__abc_21203_new_n4666_), .B(w_mem_inst__abc_21203_new_n4662_), .Y(w_mem_inst__0w_mem_9__31_0__27_));
OR2X2 OR2X2_3079 ( .A(w_mem_inst__abc_21203_new_n4671_), .B(w_mem_inst__abc_21203_new_n4669_), .Y(w_mem_inst__abc_21203_new_n4672_));
OR2X2 OR2X2_308 ( .A(_abc_15497_new_n1642_), .B(_abc_15497_new_n1629_), .Y(_abc_15497_new_n1643_));
OR2X2 OR2X2_3080 ( .A(w_mem_inst__abc_21203_new_n4672_), .B(w_mem_inst__abc_21203_new_n4668_), .Y(w_mem_inst__0w_mem_9__31_0__28_));
OR2X2 OR2X2_3081 ( .A(w_mem_inst__abc_21203_new_n4677_), .B(w_mem_inst__abc_21203_new_n4675_), .Y(w_mem_inst__abc_21203_new_n4678_));
OR2X2 OR2X2_3082 ( .A(w_mem_inst__abc_21203_new_n4678_), .B(w_mem_inst__abc_21203_new_n4674_), .Y(w_mem_inst__0w_mem_9__31_0__29_));
OR2X2 OR2X2_3083 ( .A(w_mem_inst__abc_21203_new_n4683_), .B(w_mem_inst__abc_21203_new_n4681_), .Y(w_mem_inst__abc_21203_new_n4684_));
OR2X2 OR2X2_3084 ( .A(w_mem_inst__abc_21203_new_n4684_), .B(w_mem_inst__abc_21203_new_n4680_), .Y(w_mem_inst__0w_mem_9__31_0__30_));
OR2X2 OR2X2_3085 ( .A(w_mem_inst__abc_21203_new_n4689_), .B(w_mem_inst__abc_21203_new_n4687_), .Y(w_mem_inst__abc_21203_new_n4690_));
OR2X2 OR2X2_3086 ( .A(w_mem_inst__abc_21203_new_n4690_), .B(w_mem_inst__abc_21203_new_n4686_), .Y(w_mem_inst__0w_mem_9__31_0__31_));
OR2X2 OR2X2_3087 ( .A(w_mem_inst__abc_21203_new_n4695_), .B(w_mem_inst__abc_21203_new_n4693_), .Y(w_mem_inst__abc_21203_new_n4696_));
OR2X2 OR2X2_3088 ( .A(w_mem_inst__abc_21203_new_n4696_), .B(w_mem_inst__abc_21203_new_n4692_), .Y(w_mem_inst__0w_mem_8__31_0__0_));
OR2X2 OR2X2_3089 ( .A(w_mem_inst__abc_21203_new_n4701_), .B(w_mem_inst__abc_21203_new_n4699_), .Y(w_mem_inst__abc_21203_new_n4702_));
OR2X2 OR2X2_309 ( .A(_abc_15497_new_n1633_), .B(_abc_15497_new_n1643_), .Y(_abc_15497_new_n1644_));
OR2X2 OR2X2_3090 ( .A(w_mem_inst__abc_21203_new_n4702_), .B(w_mem_inst__abc_21203_new_n4698_), .Y(w_mem_inst__0w_mem_8__31_0__1_));
OR2X2 OR2X2_3091 ( .A(w_mem_inst__abc_21203_new_n4707_), .B(w_mem_inst__abc_21203_new_n4705_), .Y(w_mem_inst__abc_21203_new_n4708_));
OR2X2 OR2X2_3092 ( .A(w_mem_inst__abc_21203_new_n4708_), .B(w_mem_inst__abc_21203_new_n4704_), .Y(w_mem_inst__0w_mem_8__31_0__2_));
OR2X2 OR2X2_3093 ( .A(w_mem_inst__abc_21203_new_n4713_), .B(w_mem_inst__abc_21203_new_n4711_), .Y(w_mem_inst__abc_21203_new_n4714_));
OR2X2 OR2X2_3094 ( .A(w_mem_inst__abc_21203_new_n4714_), .B(w_mem_inst__abc_21203_new_n4710_), .Y(w_mem_inst__0w_mem_8__31_0__3_));
OR2X2 OR2X2_3095 ( .A(w_mem_inst__abc_21203_new_n4719_), .B(w_mem_inst__abc_21203_new_n4717_), .Y(w_mem_inst__abc_21203_new_n4720_));
OR2X2 OR2X2_3096 ( .A(w_mem_inst__abc_21203_new_n4720_), .B(w_mem_inst__abc_21203_new_n4716_), .Y(w_mem_inst__0w_mem_8__31_0__4_));
OR2X2 OR2X2_3097 ( .A(w_mem_inst__abc_21203_new_n4725_), .B(w_mem_inst__abc_21203_new_n4723_), .Y(w_mem_inst__abc_21203_new_n4726_));
OR2X2 OR2X2_3098 ( .A(w_mem_inst__abc_21203_new_n4726_), .B(w_mem_inst__abc_21203_new_n4722_), .Y(w_mem_inst__0w_mem_8__31_0__5_));
OR2X2 OR2X2_3099 ( .A(w_mem_inst__abc_21203_new_n4731_), .B(w_mem_inst__abc_21203_new_n4729_), .Y(w_mem_inst__abc_21203_new_n4732_));
OR2X2 OR2X2_31 ( .A(c_reg_1_), .B(\digest[65] ), .Y(_abc_15497_new_n821_));
OR2X2 OR2X2_310 ( .A(_abc_15497_new_n1652_), .B(_abc_15497_new_n1638_), .Y(_0H3_reg_31_0__9_));
OR2X2 OR2X2_3100 ( .A(w_mem_inst__abc_21203_new_n4732_), .B(w_mem_inst__abc_21203_new_n4728_), .Y(w_mem_inst__0w_mem_8__31_0__6_));
OR2X2 OR2X2_3101 ( .A(w_mem_inst__abc_21203_new_n4737_), .B(w_mem_inst__abc_21203_new_n4735_), .Y(w_mem_inst__abc_21203_new_n4738_));
OR2X2 OR2X2_3102 ( .A(w_mem_inst__abc_21203_new_n4738_), .B(w_mem_inst__abc_21203_new_n4734_), .Y(w_mem_inst__0w_mem_8__31_0__7_));
OR2X2 OR2X2_3103 ( .A(w_mem_inst__abc_21203_new_n4743_), .B(w_mem_inst__abc_21203_new_n4741_), .Y(w_mem_inst__abc_21203_new_n4744_));
OR2X2 OR2X2_3104 ( .A(w_mem_inst__abc_21203_new_n4744_), .B(w_mem_inst__abc_21203_new_n4740_), .Y(w_mem_inst__0w_mem_8__31_0__8_));
OR2X2 OR2X2_3105 ( .A(w_mem_inst__abc_21203_new_n4749_), .B(w_mem_inst__abc_21203_new_n4747_), .Y(w_mem_inst__abc_21203_new_n4750_));
OR2X2 OR2X2_3106 ( .A(w_mem_inst__abc_21203_new_n4750_), .B(w_mem_inst__abc_21203_new_n4746_), .Y(w_mem_inst__0w_mem_8__31_0__9_));
OR2X2 OR2X2_3107 ( .A(w_mem_inst__abc_21203_new_n4755_), .B(w_mem_inst__abc_21203_new_n4753_), .Y(w_mem_inst__abc_21203_new_n4756_));
OR2X2 OR2X2_3108 ( .A(w_mem_inst__abc_21203_new_n4756_), .B(w_mem_inst__abc_21203_new_n4752_), .Y(w_mem_inst__0w_mem_8__31_0__10_));
OR2X2 OR2X2_3109 ( .A(w_mem_inst__abc_21203_new_n4761_), .B(w_mem_inst__abc_21203_new_n4759_), .Y(w_mem_inst__abc_21203_new_n4762_));
OR2X2 OR2X2_311 ( .A(\digest[42] ), .B(d_reg_10_), .Y(_abc_15497_new_n1657_));
OR2X2 OR2X2_3110 ( .A(w_mem_inst__abc_21203_new_n4762_), .B(w_mem_inst__abc_21203_new_n4758_), .Y(w_mem_inst__0w_mem_8__31_0__11_));
OR2X2 OR2X2_3111 ( .A(w_mem_inst__abc_21203_new_n4767_), .B(w_mem_inst__abc_21203_new_n4765_), .Y(w_mem_inst__abc_21203_new_n4768_));
OR2X2 OR2X2_3112 ( .A(w_mem_inst__abc_21203_new_n4768_), .B(w_mem_inst__abc_21203_new_n4764_), .Y(w_mem_inst__0w_mem_8__31_0__12_));
OR2X2 OR2X2_3113 ( .A(w_mem_inst__abc_21203_new_n4773_), .B(w_mem_inst__abc_21203_new_n4771_), .Y(w_mem_inst__abc_21203_new_n4774_));
OR2X2 OR2X2_3114 ( .A(w_mem_inst__abc_21203_new_n4774_), .B(w_mem_inst__abc_21203_new_n4770_), .Y(w_mem_inst__0w_mem_8__31_0__13_));
OR2X2 OR2X2_3115 ( .A(w_mem_inst__abc_21203_new_n4779_), .B(w_mem_inst__abc_21203_new_n4777_), .Y(w_mem_inst__abc_21203_new_n4780_));
OR2X2 OR2X2_3116 ( .A(w_mem_inst__abc_21203_new_n4780_), .B(w_mem_inst__abc_21203_new_n4776_), .Y(w_mem_inst__0w_mem_8__31_0__14_));
OR2X2 OR2X2_3117 ( .A(w_mem_inst__abc_21203_new_n4785_), .B(w_mem_inst__abc_21203_new_n4783_), .Y(w_mem_inst__abc_21203_new_n4786_));
OR2X2 OR2X2_3118 ( .A(w_mem_inst__abc_21203_new_n4786_), .B(w_mem_inst__abc_21203_new_n4782_), .Y(w_mem_inst__0w_mem_8__31_0__15_));
OR2X2 OR2X2_3119 ( .A(w_mem_inst__abc_21203_new_n4791_), .B(w_mem_inst__abc_21203_new_n4789_), .Y(w_mem_inst__abc_21203_new_n4792_));
OR2X2 OR2X2_312 ( .A(_abc_15497_new_n1656_), .B(_abc_15497_new_n1660_), .Y(_abc_15497_new_n1661_));
OR2X2 OR2X2_3120 ( .A(w_mem_inst__abc_21203_new_n4792_), .B(w_mem_inst__abc_21203_new_n4788_), .Y(w_mem_inst__0w_mem_8__31_0__16_));
OR2X2 OR2X2_3121 ( .A(w_mem_inst__abc_21203_new_n4797_), .B(w_mem_inst__abc_21203_new_n4795_), .Y(w_mem_inst__abc_21203_new_n4798_));
OR2X2 OR2X2_3122 ( .A(w_mem_inst__abc_21203_new_n4798_), .B(w_mem_inst__abc_21203_new_n4794_), .Y(w_mem_inst__0w_mem_8__31_0__17_));
OR2X2 OR2X2_3123 ( .A(w_mem_inst__abc_21203_new_n4803_), .B(w_mem_inst__abc_21203_new_n4801_), .Y(w_mem_inst__abc_21203_new_n4804_));
OR2X2 OR2X2_3124 ( .A(w_mem_inst__abc_21203_new_n4804_), .B(w_mem_inst__abc_21203_new_n4800_), .Y(w_mem_inst__0w_mem_8__31_0__18_));
OR2X2 OR2X2_3125 ( .A(w_mem_inst__abc_21203_new_n4809_), .B(w_mem_inst__abc_21203_new_n4807_), .Y(w_mem_inst__abc_21203_new_n4810_));
OR2X2 OR2X2_3126 ( .A(w_mem_inst__abc_21203_new_n4810_), .B(w_mem_inst__abc_21203_new_n4806_), .Y(w_mem_inst__0w_mem_8__31_0__19_));
OR2X2 OR2X2_3127 ( .A(w_mem_inst__abc_21203_new_n4815_), .B(w_mem_inst__abc_21203_new_n4813_), .Y(w_mem_inst__abc_21203_new_n4816_));
OR2X2 OR2X2_3128 ( .A(w_mem_inst__abc_21203_new_n4816_), .B(w_mem_inst__abc_21203_new_n4812_), .Y(w_mem_inst__0w_mem_8__31_0__20_));
OR2X2 OR2X2_3129 ( .A(w_mem_inst__abc_21203_new_n4821_), .B(w_mem_inst__abc_21203_new_n4819_), .Y(w_mem_inst__abc_21203_new_n4822_));
OR2X2 OR2X2_313 ( .A(_abc_15497_new_n699_), .B(\digest[42] ), .Y(_abc_15497_new_n1666_));
OR2X2 OR2X2_3130 ( .A(w_mem_inst__abc_21203_new_n4822_), .B(w_mem_inst__abc_21203_new_n4818_), .Y(w_mem_inst__0w_mem_8__31_0__21_));
OR2X2 OR2X2_3131 ( .A(w_mem_inst__abc_21203_new_n4827_), .B(w_mem_inst__abc_21203_new_n4825_), .Y(w_mem_inst__abc_21203_new_n4828_));
OR2X2 OR2X2_3132 ( .A(w_mem_inst__abc_21203_new_n4828_), .B(w_mem_inst__abc_21203_new_n4824_), .Y(w_mem_inst__0w_mem_8__31_0__22_));
OR2X2 OR2X2_3133 ( .A(w_mem_inst__abc_21203_new_n4833_), .B(w_mem_inst__abc_21203_new_n4831_), .Y(w_mem_inst__abc_21203_new_n4834_));
OR2X2 OR2X2_3134 ( .A(w_mem_inst__abc_21203_new_n4834_), .B(w_mem_inst__abc_21203_new_n4830_), .Y(w_mem_inst__0w_mem_8__31_0__23_));
OR2X2 OR2X2_3135 ( .A(w_mem_inst__abc_21203_new_n4839_), .B(w_mem_inst__abc_21203_new_n4837_), .Y(w_mem_inst__abc_21203_new_n4840_));
OR2X2 OR2X2_3136 ( .A(w_mem_inst__abc_21203_new_n4840_), .B(w_mem_inst__abc_21203_new_n4836_), .Y(w_mem_inst__0w_mem_8__31_0__24_));
OR2X2 OR2X2_3137 ( .A(w_mem_inst__abc_21203_new_n4845_), .B(w_mem_inst__abc_21203_new_n4843_), .Y(w_mem_inst__abc_21203_new_n4846_));
OR2X2 OR2X2_3138 ( .A(w_mem_inst__abc_21203_new_n4846_), .B(w_mem_inst__abc_21203_new_n4842_), .Y(w_mem_inst__0w_mem_8__31_0__25_));
OR2X2 OR2X2_3139 ( .A(w_mem_inst__abc_21203_new_n4851_), .B(w_mem_inst__abc_21203_new_n4849_), .Y(w_mem_inst__abc_21203_new_n4852_));
OR2X2 OR2X2_314 ( .A(_abc_15497_new_n1665_), .B(_abc_15497_new_n1667_), .Y(_0H3_reg_31_0__10_));
OR2X2 OR2X2_3140 ( .A(w_mem_inst__abc_21203_new_n4852_), .B(w_mem_inst__abc_21203_new_n4848_), .Y(w_mem_inst__0w_mem_8__31_0__26_));
OR2X2 OR2X2_3141 ( .A(w_mem_inst__abc_21203_new_n4857_), .B(w_mem_inst__abc_21203_new_n4855_), .Y(w_mem_inst__abc_21203_new_n4858_));
OR2X2 OR2X2_3142 ( .A(w_mem_inst__abc_21203_new_n4858_), .B(w_mem_inst__abc_21203_new_n4854_), .Y(w_mem_inst__0w_mem_8__31_0__27_));
OR2X2 OR2X2_3143 ( .A(w_mem_inst__abc_21203_new_n4863_), .B(w_mem_inst__abc_21203_new_n4861_), .Y(w_mem_inst__abc_21203_new_n4864_));
OR2X2 OR2X2_3144 ( .A(w_mem_inst__abc_21203_new_n4864_), .B(w_mem_inst__abc_21203_new_n4860_), .Y(w_mem_inst__0w_mem_8__31_0__28_));
OR2X2 OR2X2_3145 ( .A(w_mem_inst__abc_21203_new_n4869_), .B(w_mem_inst__abc_21203_new_n4867_), .Y(w_mem_inst__abc_21203_new_n4870_));
OR2X2 OR2X2_3146 ( .A(w_mem_inst__abc_21203_new_n4870_), .B(w_mem_inst__abc_21203_new_n4866_), .Y(w_mem_inst__0w_mem_8__31_0__29_));
OR2X2 OR2X2_3147 ( .A(w_mem_inst__abc_21203_new_n4875_), .B(w_mem_inst__abc_21203_new_n4873_), .Y(w_mem_inst__abc_21203_new_n4876_));
OR2X2 OR2X2_3148 ( .A(w_mem_inst__abc_21203_new_n4876_), .B(w_mem_inst__abc_21203_new_n4872_), .Y(w_mem_inst__0w_mem_8__31_0__30_));
OR2X2 OR2X2_3149 ( .A(w_mem_inst__abc_21203_new_n4881_), .B(w_mem_inst__abc_21203_new_n4879_), .Y(w_mem_inst__abc_21203_new_n4882_));
OR2X2 OR2X2_315 ( .A(\digest[43] ), .B(d_reg_11_), .Y(_abc_15497_new_n1672_));
OR2X2 OR2X2_3150 ( .A(w_mem_inst__abc_21203_new_n4882_), .B(w_mem_inst__abc_21203_new_n4878_), .Y(w_mem_inst__0w_mem_8__31_0__31_));
OR2X2 OR2X2_3151 ( .A(w_mem_inst__abc_21203_new_n4887_), .B(w_mem_inst__abc_21203_new_n4885_), .Y(w_mem_inst__abc_21203_new_n4888_));
OR2X2 OR2X2_3152 ( .A(w_mem_inst__abc_21203_new_n4888_), .B(w_mem_inst__abc_21203_new_n4884_), .Y(w_mem_inst__0w_mem_4__31_0__0_));
OR2X2 OR2X2_3153 ( .A(w_mem_inst__abc_21203_new_n4893_), .B(w_mem_inst__abc_21203_new_n4891_), .Y(w_mem_inst__abc_21203_new_n4894_));
OR2X2 OR2X2_3154 ( .A(w_mem_inst__abc_21203_new_n4894_), .B(w_mem_inst__abc_21203_new_n4890_), .Y(w_mem_inst__0w_mem_4__31_0__1_));
OR2X2 OR2X2_3155 ( .A(w_mem_inst__abc_21203_new_n4899_), .B(w_mem_inst__abc_21203_new_n4897_), .Y(w_mem_inst__abc_21203_new_n4900_));
OR2X2 OR2X2_3156 ( .A(w_mem_inst__abc_21203_new_n4900_), .B(w_mem_inst__abc_21203_new_n4896_), .Y(w_mem_inst__0w_mem_4__31_0__2_));
OR2X2 OR2X2_3157 ( .A(w_mem_inst__abc_21203_new_n4905_), .B(w_mem_inst__abc_21203_new_n4903_), .Y(w_mem_inst__abc_21203_new_n4906_));
OR2X2 OR2X2_3158 ( .A(w_mem_inst__abc_21203_new_n4906_), .B(w_mem_inst__abc_21203_new_n4902_), .Y(w_mem_inst__0w_mem_4__31_0__3_));
OR2X2 OR2X2_3159 ( .A(w_mem_inst__abc_21203_new_n4911_), .B(w_mem_inst__abc_21203_new_n4909_), .Y(w_mem_inst__abc_21203_new_n4912_));
OR2X2 OR2X2_316 ( .A(_abc_15497_new_n1671_), .B(_abc_15497_new_n1675_), .Y(_abc_15497_new_n1676_));
OR2X2 OR2X2_3160 ( .A(w_mem_inst__abc_21203_new_n4912_), .B(w_mem_inst__abc_21203_new_n4908_), .Y(w_mem_inst__0w_mem_4__31_0__4_));
OR2X2 OR2X2_3161 ( .A(w_mem_inst__abc_21203_new_n4917_), .B(w_mem_inst__abc_21203_new_n4915_), .Y(w_mem_inst__abc_21203_new_n4918_));
OR2X2 OR2X2_3162 ( .A(w_mem_inst__abc_21203_new_n4918_), .B(w_mem_inst__abc_21203_new_n4914_), .Y(w_mem_inst__0w_mem_4__31_0__5_));
OR2X2 OR2X2_3163 ( .A(w_mem_inst__abc_21203_new_n4923_), .B(w_mem_inst__abc_21203_new_n4921_), .Y(w_mem_inst__abc_21203_new_n4924_));
OR2X2 OR2X2_3164 ( .A(w_mem_inst__abc_21203_new_n4924_), .B(w_mem_inst__abc_21203_new_n4920_), .Y(w_mem_inst__0w_mem_4__31_0__6_));
OR2X2 OR2X2_3165 ( .A(w_mem_inst__abc_21203_new_n4929_), .B(w_mem_inst__abc_21203_new_n4927_), .Y(w_mem_inst__abc_21203_new_n4930_));
OR2X2 OR2X2_3166 ( .A(w_mem_inst__abc_21203_new_n4930_), .B(w_mem_inst__abc_21203_new_n4926_), .Y(w_mem_inst__0w_mem_4__31_0__7_));
OR2X2 OR2X2_3167 ( .A(w_mem_inst__abc_21203_new_n4935_), .B(w_mem_inst__abc_21203_new_n4933_), .Y(w_mem_inst__abc_21203_new_n4936_));
OR2X2 OR2X2_3168 ( .A(w_mem_inst__abc_21203_new_n4936_), .B(w_mem_inst__abc_21203_new_n4932_), .Y(w_mem_inst__0w_mem_4__31_0__8_));
OR2X2 OR2X2_3169 ( .A(w_mem_inst__abc_21203_new_n4941_), .B(w_mem_inst__abc_21203_new_n4939_), .Y(w_mem_inst__abc_21203_new_n4942_));
OR2X2 OR2X2_317 ( .A(_abc_15497_new_n1670_), .B(_abc_15497_new_n1677_), .Y(_abc_15497_new_n1678_));
OR2X2 OR2X2_3170 ( .A(w_mem_inst__abc_21203_new_n4942_), .B(w_mem_inst__abc_21203_new_n4938_), .Y(w_mem_inst__0w_mem_4__31_0__9_));
OR2X2 OR2X2_3171 ( .A(w_mem_inst__abc_21203_new_n4947_), .B(w_mem_inst__abc_21203_new_n4945_), .Y(w_mem_inst__abc_21203_new_n4948_));
OR2X2 OR2X2_3172 ( .A(w_mem_inst__abc_21203_new_n4948_), .B(w_mem_inst__abc_21203_new_n4944_), .Y(w_mem_inst__0w_mem_4__31_0__10_));
OR2X2 OR2X2_3173 ( .A(w_mem_inst__abc_21203_new_n4953_), .B(w_mem_inst__abc_21203_new_n4951_), .Y(w_mem_inst__abc_21203_new_n4954_));
OR2X2 OR2X2_3174 ( .A(w_mem_inst__abc_21203_new_n4954_), .B(w_mem_inst__abc_21203_new_n4950_), .Y(w_mem_inst__0w_mem_4__31_0__11_));
OR2X2 OR2X2_3175 ( .A(w_mem_inst__abc_21203_new_n4959_), .B(w_mem_inst__abc_21203_new_n4957_), .Y(w_mem_inst__abc_21203_new_n4960_));
OR2X2 OR2X2_3176 ( .A(w_mem_inst__abc_21203_new_n4960_), .B(w_mem_inst__abc_21203_new_n4956_), .Y(w_mem_inst__0w_mem_4__31_0__12_));
OR2X2 OR2X2_3177 ( .A(w_mem_inst__abc_21203_new_n4965_), .B(w_mem_inst__abc_21203_new_n4963_), .Y(w_mem_inst__abc_21203_new_n4966_));
OR2X2 OR2X2_3178 ( .A(w_mem_inst__abc_21203_new_n4966_), .B(w_mem_inst__abc_21203_new_n4962_), .Y(w_mem_inst__0w_mem_4__31_0__13_));
OR2X2 OR2X2_3179 ( .A(w_mem_inst__abc_21203_new_n4971_), .B(w_mem_inst__abc_21203_new_n4969_), .Y(w_mem_inst__abc_21203_new_n4972_));
OR2X2 OR2X2_318 ( .A(_abc_15497_new_n1680_), .B(_abc_15497_new_n1669_), .Y(_0H3_reg_31_0__11_));
OR2X2 OR2X2_3180 ( .A(w_mem_inst__abc_21203_new_n4972_), .B(w_mem_inst__abc_21203_new_n4968_), .Y(w_mem_inst__0w_mem_4__31_0__14_));
OR2X2 OR2X2_3181 ( .A(w_mem_inst__abc_21203_new_n4977_), .B(w_mem_inst__abc_21203_new_n4975_), .Y(w_mem_inst__abc_21203_new_n4978_));
OR2X2 OR2X2_3182 ( .A(w_mem_inst__abc_21203_new_n4978_), .B(w_mem_inst__abc_21203_new_n4974_), .Y(w_mem_inst__0w_mem_4__31_0__15_));
OR2X2 OR2X2_3183 ( .A(w_mem_inst__abc_21203_new_n4983_), .B(w_mem_inst__abc_21203_new_n4981_), .Y(w_mem_inst__abc_21203_new_n4984_));
OR2X2 OR2X2_3184 ( .A(w_mem_inst__abc_21203_new_n4984_), .B(w_mem_inst__abc_21203_new_n4980_), .Y(w_mem_inst__0w_mem_4__31_0__16_));
OR2X2 OR2X2_3185 ( .A(w_mem_inst__abc_21203_new_n4989_), .B(w_mem_inst__abc_21203_new_n4987_), .Y(w_mem_inst__abc_21203_new_n4990_));
OR2X2 OR2X2_3186 ( .A(w_mem_inst__abc_21203_new_n4990_), .B(w_mem_inst__abc_21203_new_n4986_), .Y(w_mem_inst__0w_mem_4__31_0__17_));
OR2X2 OR2X2_3187 ( .A(w_mem_inst__abc_21203_new_n4995_), .B(w_mem_inst__abc_21203_new_n4993_), .Y(w_mem_inst__abc_21203_new_n4996_));
OR2X2 OR2X2_3188 ( .A(w_mem_inst__abc_21203_new_n4996_), .B(w_mem_inst__abc_21203_new_n4992_), .Y(w_mem_inst__0w_mem_4__31_0__18_));
OR2X2 OR2X2_3189 ( .A(w_mem_inst__abc_21203_new_n5001_), .B(w_mem_inst__abc_21203_new_n4999_), .Y(w_mem_inst__abc_21203_new_n5002_));
OR2X2 OR2X2_319 ( .A(_abc_15497_new_n1687_), .B(_abc_15497_new_n1673_), .Y(_abc_15497_new_n1688_));
OR2X2 OR2X2_3190 ( .A(w_mem_inst__abc_21203_new_n5002_), .B(w_mem_inst__abc_21203_new_n4998_), .Y(w_mem_inst__0w_mem_4__31_0__19_));
OR2X2 OR2X2_3191 ( .A(w_mem_inst__abc_21203_new_n5007_), .B(w_mem_inst__abc_21203_new_n5005_), .Y(w_mem_inst__abc_21203_new_n5008_));
OR2X2 OR2X2_3192 ( .A(w_mem_inst__abc_21203_new_n5008_), .B(w_mem_inst__abc_21203_new_n5004_), .Y(w_mem_inst__0w_mem_4__31_0__20_));
OR2X2 OR2X2_3193 ( .A(w_mem_inst__abc_21203_new_n5013_), .B(w_mem_inst__abc_21203_new_n5011_), .Y(w_mem_inst__abc_21203_new_n5014_));
OR2X2 OR2X2_3194 ( .A(w_mem_inst__abc_21203_new_n5014_), .B(w_mem_inst__abc_21203_new_n5010_), .Y(w_mem_inst__0w_mem_4__31_0__21_));
OR2X2 OR2X2_3195 ( .A(w_mem_inst__abc_21203_new_n5019_), .B(w_mem_inst__abc_21203_new_n5017_), .Y(w_mem_inst__abc_21203_new_n5020_));
OR2X2 OR2X2_3196 ( .A(w_mem_inst__abc_21203_new_n5020_), .B(w_mem_inst__abc_21203_new_n5016_), .Y(w_mem_inst__0w_mem_4__31_0__22_));
OR2X2 OR2X2_3197 ( .A(w_mem_inst__abc_21203_new_n5025_), .B(w_mem_inst__abc_21203_new_n5023_), .Y(w_mem_inst__abc_21203_new_n5026_));
OR2X2 OR2X2_3198 ( .A(w_mem_inst__abc_21203_new_n5026_), .B(w_mem_inst__abc_21203_new_n5022_), .Y(w_mem_inst__0w_mem_4__31_0__23_));
OR2X2 OR2X2_3199 ( .A(w_mem_inst__abc_21203_new_n5031_), .B(w_mem_inst__abc_21203_new_n5029_), .Y(w_mem_inst__abc_21203_new_n5032_));
OR2X2 OR2X2_32 ( .A(_abc_15497_new_n823_), .B(_abc_15497_new_n818_), .Y(_abc_15497_new_n824_));
OR2X2 OR2X2_320 ( .A(_abc_15497_new_n1686_), .B(_abc_15497_new_n1688_), .Y(_abc_15497_new_n1689_));
OR2X2 OR2X2_3200 ( .A(w_mem_inst__abc_21203_new_n5032_), .B(w_mem_inst__abc_21203_new_n5028_), .Y(w_mem_inst__0w_mem_4__31_0__24_));
OR2X2 OR2X2_3201 ( .A(w_mem_inst__abc_21203_new_n5037_), .B(w_mem_inst__abc_21203_new_n5035_), .Y(w_mem_inst__abc_21203_new_n5038_));
OR2X2 OR2X2_3202 ( .A(w_mem_inst__abc_21203_new_n5038_), .B(w_mem_inst__abc_21203_new_n5034_), .Y(w_mem_inst__0w_mem_4__31_0__25_));
OR2X2 OR2X2_3203 ( .A(w_mem_inst__abc_21203_new_n5043_), .B(w_mem_inst__abc_21203_new_n5041_), .Y(w_mem_inst__abc_21203_new_n5044_));
OR2X2 OR2X2_3204 ( .A(w_mem_inst__abc_21203_new_n5044_), .B(w_mem_inst__abc_21203_new_n5040_), .Y(w_mem_inst__0w_mem_4__31_0__26_));
OR2X2 OR2X2_3205 ( .A(w_mem_inst__abc_21203_new_n5049_), .B(w_mem_inst__abc_21203_new_n5047_), .Y(w_mem_inst__abc_21203_new_n5050_));
OR2X2 OR2X2_3206 ( .A(w_mem_inst__abc_21203_new_n5050_), .B(w_mem_inst__abc_21203_new_n5046_), .Y(w_mem_inst__0w_mem_4__31_0__27_));
OR2X2 OR2X2_3207 ( .A(w_mem_inst__abc_21203_new_n5055_), .B(w_mem_inst__abc_21203_new_n5053_), .Y(w_mem_inst__abc_21203_new_n5056_));
OR2X2 OR2X2_3208 ( .A(w_mem_inst__abc_21203_new_n5056_), .B(w_mem_inst__abc_21203_new_n5052_), .Y(w_mem_inst__0w_mem_4__31_0__28_));
OR2X2 OR2X2_3209 ( .A(w_mem_inst__abc_21203_new_n5061_), .B(w_mem_inst__abc_21203_new_n5059_), .Y(w_mem_inst__abc_21203_new_n5062_));
OR2X2 OR2X2_321 ( .A(_abc_15497_new_n1684_), .B(_abc_15497_new_n1689_), .Y(_abc_15497_new_n1690_));
OR2X2 OR2X2_3210 ( .A(w_mem_inst__abc_21203_new_n5062_), .B(w_mem_inst__abc_21203_new_n5058_), .Y(w_mem_inst__0w_mem_4__31_0__29_));
OR2X2 OR2X2_3211 ( .A(w_mem_inst__abc_21203_new_n5067_), .B(w_mem_inst__abc_21203_new_n5065_), .Y(w_mem_inst__abc_21203_new_n5068_));
OR2X2 OR2X2_3212 ( .A(w_mem_inst__abc_21203_new_n5068_), .B(w_mem_inst__abc_21203_new_n5064_), .Y(w_mem_inst__0w_mem_4__31_0__30_));
OR2X2 OR2X2_3213 ( .A(w_mem_inst__abc_21203_new_n5073_), .B(w_mem_inst__abc_21203_new_n5071_), .Y(w_mem_inst__abc_21203_new_n5074_));
OR2X2 OR2X2_3214 ( .A(w_mem_inst__abc_21203_new_n5074_), .B(w_mem_inst__abc_21203_new_n5070_), .Y(w_mem_inst__0w_mem_4__31_0__31_));
OR2X2 OR2X2_3215 ( .A(w_mem_inst__abc_21203_new_n5079_), .B(w_mem_inst__abc_21203_new_n5077_), .Y(w_mem_inst__abc_21203_new_n5080_));
OR2X2 OR2X2_3216 ( .A(w_mem_inst__abc_21203_new_n5080_), .B(w_mem_inst__abc_21203_new_n5076_), .Y(w_mem_inst__0w_mem_6__31_0__0_));
OR2X2 OR2X2_3217 ( .A(w_mem_inst__abc_21203_new_n5085_), .B(w_mem_inst__abc_21203_new_n5083_), .Y(w_mem_inst__abc_21203_new_n5086_));
OR2X2 OR2X2_3218 ( .A(w_mem_inst__abc_21203_new_n5086_), .B(w_mem_inst__abc_21203_new_n5082_), .Y(w_mem_inst__0w_mem_6__31_0__1_));
OR2X2 OR2X2_3219 ( .A(w_mem_inst__abc_21203_new_n5091_), .B(w_mem_inst__abc_21203_new_n5089_), .Y(w_mem_inst__abc_21203_new_n5092_));
OR2X2 OR2X2_322 ( .A(\digest[44] ), .B(d_reg_12_), .Y(_abc_15497_new_n1691_));
OR2X2 OR2X2_3220 ( .A(w_mem_inst__abc_21203_new_n5092_), .B(w_mem_inst__abc_21203_new_n5088_), .Y(w_mem_inst__0w_mem_6__31_0__2_));
OR2X2 OR2X2_3221 ( .A(w_mem_inst__abc_21203_new_n5097_), .B(w_mem_inst__abc_21203_new_n5095_), .Y(w_mem_inst__abc_21203_new_n5098_));
OR2X2 OR2X2_3222 ( .A(w_mem_inst__abc_21203_new_n5098_), .B(w_mem_inst__abc_21203_new_n5094_), .Y(w_mem_inst__0w_mem_6__31_0__3_));
OR2X2 OR2X2_3223 ( .A(w_mem_inst__abc_21203_new_n5103_), .B(w_mem_inst__abc_21203_new_n5101_), .Y(w_mem_inst__abc_21203_new_n5104_));
OR2X2 OR2X2_3224 ( .A(w_mem_inst__abc_21203_new_n5104_), .B(w_mem_inst__abc_21203_new_n5100_), .Y(w_mem_inst__0w_mem_6__31_0__4_));
OR2X2 OR2X2_3225 ( .A(w_mem_inst__abc_21203_new_n5109_), .B(w_mem_inst__abc_21203_new_n5107_), .Y(w_mem_inst__abc_21203_new_n5110_));
OR2X2 OR2X2_3226 ( .A(w_mem_inst__abc_21203_new_n5110_), .B(w_mem_inst__abc_21203_new_n5106_), .Y(w_mem_inst__0w_mem_6__31_0__5_));
OR2X2 OR2X2_3227 ( .A(w_mem_inst__abc_21203_new_n5115_), .B(w_mem_inst__abc_21203_new_n5113_), .Y(w_mem_inst__abc_21203_new_n5116_));
OR2X2 OR2X2_3228 ( .A(w_mem_inst__abc_21203_new_n5116_), .B(w_mem_inst__abc_21203_new_n5112_), .Y(w_mem_inst__0w_mem_6__31_0__6_));
OR2X2 OR2X2_3229 ( .A(w_mem_inst__abc_21203_new_n5121_), .B(w_mem_inst__abc_21203_new_n5119_), .Y(w_mem_inst__abc_21203_new_n5122_));
OR2X2 OR2X2_323 ( .A(_abc_15497_new_n1690_), .B(_abc_15497_new_n1694_), .Y(_abc_15497_new_n1695_));
OR2X2 OR2X2_3230 ( .A(w_mem_inst__abc_21203_new_n5122_), .B(w_mem_inst__abc_21203_new_n5118_), .Y(w_mem_inst__0w_mem_6__31_0__7_));
OR2X2 OR2X2_3231 ( .A(w_mem_inst__abc_21203_new_n5127_), .B(w_mem_inst__abc_21203_new_n5125_), .Y(w_mem_inst__abc_21203_new_n5128_));
OR2X2 OR2X2_3232 ( .A(w_mem_inst__abc_21203_new_n5128_), .B(w_mem_inst__abc_21203_new_n5124_), .Y(w_mem_inst__0w_mem_6__31_0__8_));
OR2X2 OR2X2_3233 ( .A(w_mem_inst__abc_21203_new_n5133_), .B(w_mem_inst__abc_21203_new_n5131_), .Y(w_mem_inst__abc_21203_new_n5134_));
OR2X2 OR2X2_3234 ( .A(w_mem_inst__abc_21203_new_n5134_), .B(w_mem_inst__abc_21203_new_n5130_), .Y(w_mem_inst__0w_mem_6__31_0__9_));
OR2X2 OR2X2_3235 ( .A(w_mem_inst__abc_21203_new_n5139_), .B(w_mem_inst__abc_21203_new_n5137_), .Y(w_mem_inst__abc_21203_new_n5140_));
OR2X2 OR2X2_3236 ( .A(w_mem_inst__abc_21203_new_n5140_), .B(w_mem_inst__abc_21203_new_n5136_), .Y(w_mem_inst__0w_mem_6__31_0__10_));
OR2X2 OR2X2_3237 ( .A(w_mem_inst__abc_21203_new_n5145_), .B(w_mem_inst__abc_21203_new_n5143_), .Y(w_mem_inst__abc_21203_new_n5146_));
OR2X2 OR2X2_3238 ( .A(w_mem_inst__abc_21203_new_n5146_), .B(w_mem_inst__abc_21203_new_n5142_), .Y(w_mem_inst__0w_mem_6__31_0__11_));
OR2X2 OR2X2_3239 ( .A(w_mem_inst__abc_21203_new_n5151_), .B(w_mem_inst__abc_21203_new_n5149_), .Y(w_mem_inst__abc_21203_new_n5152_));
OR2X2 OR2X2_324 ( .A(_abc_15497_new_n699_), .B(\digest[44] ), .Y(_abc_15497_new_n1700_));
OR2X2 OR2X2_3240 ( .A(w_mem_inst__abc_21203_new_n5152_), .B(w_mem_inst__abc_21203_new_n5148_), .Y(w_mem_inst__0w_mem_6__31_0__12_));
OR2X2 OR2X2_3241 ( .A(w_mem_inst__abc_21203_new_n5157_), .B(w_mem_inst__abc_21203_new_n5155_), .Y(w_mem_inst__abc_21203_new_n5158_));
OR2X2 OR2X2_3242 ( .A(w_mem_inst__abc_21203_new_n5158_), .B(w_mem_inst__abc_21203_new_n5154_), .Y(w_mem_inst__0w_mem_6__31_0__13_));
OR2X2 OR2X2_3243 ( .A(w_mem_inst__abc_21203_new_n5163_), .B(w_mem_inst__abc_21203_new_n5161_), .Y(w_mem_inst__abc_21203_new_n5164_));
OR2X2 OR2X2_3244 ( .A(w_mem_inst__abc_21203_new_n5164_), .B(w_mem_inst__abc_21203_new_n5160_), .Y(w_mem_inst__0w_mem_6__31_0__14_));
OR2X2 OR2X2_3245 ( .A(w_mem_inst__abc_21203_new_n5169_), .B(w_mem_inst__abc_21203_new_n5167_), .Y(w_mem_inst__abc_21203_new_n5170_));
OR2X2 OR2X2_3246 ( .A(w_mem_inst__abc_21203_new_n5170_), .B(w_mem_inst__abc_21203_new_n5166_), .Y(w_mem_inst__0w_mem_6__31_0__15_));
OR2X2 OR2X2_3247 ( .A(w_mem_inst__abc_21203_new_n5175_), .B(w_mem_inst__abc_21203_new_n5173_), .Y(w_mem_inst__abc_21203_new_n5176_));
OR2X2 OR2X2_3248 ( .A(w_mem_inst__abc_21203_new_n5176_), .B(w_mem_inst__abc_21203_new_n5172_), .Y(w_mem_inst__0w_mem_6__31_0__16_));
OR2X2 OR2X2_3249 ( .A(w_mem_inst__abc_21203_new_n5181_), .B(w_mem_inst__abc_21203_new_n5179_), .Y(w_mem_inst__abc_21203_new_n5182_));
OR2X2 OR2X2_325 ( .A(_abc_15497_new_n1699_), .B(_abc_15497_new_n1701_), .Y(_0H3_reg_31_0__12_));
OR2X2 OR2X2_3250 ( .A(w_mem_inst__abc_21203_new_n5182_), .B(w_mem_inst__abc_21203_new_n5178_), .Y(w_mem_inst__0w_mem_6__31_0__17_));
OR2X2 OR2X2_3251 ( .A(w_mem_inst__abc_21203_new_n5187_), .B(w_mem_inst__abc_21203_new_n5185_), .Y(w_mem_inst__abc_21203_new_n5188_));
OR2X2 OR2X2_3252 ( .A(w_mem_inst__abc_21203_new_n5188_), .B(w_mem_inst__abc_21203_new_n5184_), .Y(w_mem_inst__0w_mem_6__31_0__18_));
OR2X2 OR2X2_3253 ( .A(w_mem_inst__abc_21203_new_n5193_), .B(w_mem_inst__abc_21203_new_n5191_), .Y(w_mem_inst__abc_21203_new_n5194_));
OR2X2 OR2X2_3254 ( .A(w_mem_inst__abc_21203_new_n5194_), .B(w_mem_inst__abc_21203_new_n5190_), .Y(w_mem_inst__0w_mem_6__31_0__19_));
OR2X2 OR2X2_3255 ( .A(w_mem_inst__abc_21203_new_n5199_), .B(w_mem_inst__abc_21203_new_n5197_), .Y(w_mem_inst__abc_21203_new_n5200_));
OR2X2 OR2X2_3256 ( .A(w_mem_inst__abc_21203_new_n5200_), .B(w_mem_inst__abc_21203_new_n5196_), .Y(w_mem_inst__0w_mem_6__31_0__20_));
OR2X2 OR2X2_3257 ( .A(w_mem_inst__abc_21203_new_n5205_), .B(w_mem_inst__abc_21203_new_n5203_), .Y(w_mem_inst__abc_21203_new_n5206_));
OR2X2 OR2X2_3258 ( .A(w_mem_inst__abc_21203_new_n5206_), .B(w_mem_inst__abc_21203_new_n5202_), .Y(w_mem_inst__0w_mem_6__31_0__21_));
OR2X2 OR2X2_3259 ( .A(w_mem_inst__abc_21203_new_n5211_), .B(w_mem_inst__abc_21203_new_n5209_), .Y(w_mem_inst__abc_21203_new_n5212_));
OR2X2 OR2X2_326 ( .A(\digest[45] ), .B(d_reg_13_), .Y(_abc_15497_new_n1704_));
OR2X2 OR2X2_3260 ( .A(w_mem_inst__abc_21203_new_n5212_), .B(w_mem_inst__abc_21203_new_n5208_), .Y(w_mem_inst__0w_mem_6__31_0__22_));
OR2X2 OR2X2_3261 ( .A(w_mem_inst__abc_21203_new_n5217_), .B(w_mem_inst__abc_21203_new_n5215_), .Y(w_mem_inst__abc_21203_new_n5218_));
OR2X2 OR2X2_3262 ( .A(w_mem_inst__abc_21203_new_n5218_), .B(w_mem_inst__abc_21203_new_n5214_), .Y(w_mem_inst__0w_mem_6__31_0__23_));
OR2X2 OR2X2_3263 ( .A(w_mem_inst__abc_21203_new_n5223_), .B(w_mem_inst__abc_21203_new_n5221_), .Y(w_mem_inst__abc_21203_new_n5224_));
OR2X2 OR2X2_3264 ( .A(w_mem_inst__abc_21203_new_n5224_), .B(w_mem_inst__abc_21203_new_n5220_), .Y(w_mem_inst__0w_mem_6__31_0__24_));
OR2X2 OR2X2_3265 ( .A(w_mem_inst__abc_21203_new_n5229_), .B(w_mem_inst__abc_21203_new_n5227_), .Y(w_mem_inst__abc_21203_new_n5230_));
OR2X2 OR2X2_3266 ( .A(w_mem_inst__abc_21203_new_n5230_), .B(w_mem_inst__abc_21203_new_n5226_), .Y(w_mem_inst__0w_mem_6__31_0__25_));
OR2X2 OR2X2_3267 ( .A(w_mem_inst__abc_21203_new_n5235_), .B(w_mem_inst__abc_21203_new_n5233_), .Y(w_mem_inst__abc_21203_new_n5236_));
OR2X2 OR2X2_3268 ( .A(w_mem_inst__abc_21203_new_n5236_), .B(w_mem_inst__abc_21203_new_n5232_), .Y(w_mem_inst__0w_mem_6__31_0__26_));
OR2X2 OR2X2_3269 ( .A(w_mem_inst__abc_21203_new_n5241_), .B(w_mem_inst__abc_21203_new_n5239_), .Y(w_mem_inst__abc_21203_new_n5242_));
OR2X2 OR2X2_327 ( .A(_abc_15497_new_n1707_), .B(_abc_15497_new_n1692_), .Y(_abc_15497_new_n1708_));
OR2X2 OR2X2_3270 ( .A(w_mem_inst__abc_21203_new_n5242_), .B(w_mem_inst__abc_21203_new_n5238_), .Y(w_mem_inst__0w_mem_6__31_0__27_));
OR2X2 OR2X2_3271 ( .A(w_mem_inst__abc_21203_new_n5247_), .B(w_mem_inst__abc_21203_new_n5245_), .Y(w_mem_inst__abc_21203_new_n5248_));
OR2X2 OR2X2_3272 ( .A(w_mem_inst__abc_21203_new_n5248_), .B(w_mem_inst__abc_21203_new_n5244_), .Y(w_mem_inst__0w_mem_6__31_0__28_));
OR2X2 OR2X2_3273 ( .A(w_mem_inst__abc_21203_new_n5253_), .B(w_mem_inst__abc_21203_new_n5251_), .Y(w_mem_inst__abc_21203_new_n5254_));
OR2X2 OR2X2_3274 ( .A(w_mem_inst__abc_21203_new_n5254_), .B(w_mem_inst__abc_21203_new_n5250_), .Y(w_mem_inst__0w_mem_6__31_0__29_));
OR2X2 OR2X2_3275 ( .A(w_mem_inst__abc_21203_new_n5259_), .B(w_mem_inst__abc_21203_new_n5257_), .Y(w_mem_inst__abc_21203_new_n5260_));
OR2X2 OR2X2_3276 ( .A(w_mem_inst__abc_21203_new_n5260_), .B(w_mem_inst__abc_21203_new_n5256_), .Y(w_mem_inst__0w_mem_6__31_0__30_));
OR2X2 OR2X2_3277 ( .A(w_mem_inst__abc_21203_new_n5265_), .B(w_mem_inst__abc_21203_new_n5263_), .Y(w_mem_inst__abc_21203_new_n5266_));
OR2X2 OR2X2_3278 ( .A(w_mem_inst__abc_21203_new_n5266_), .B(w_mem_inst__abc_21203_new_n5262_), .Y(w_mem_inst__0w_mem_6__31_0__31_));
OR2X2 OR2X2_3279 ( .A(w_mem_inst__abc_21203_new_n5271_), .B(w_mem_inst__abc_21203_new_n5269_), .Y(w_mem_inst__abc_21203_new_n5272_));
OR2X2 OR2X2_328 ( .A(_abc_15497_new_n1696_), .B(_abc_15497_new_n1708_), .Y(_abc_15497_new_n1709_));
OR2X2 OR2X2_3280 ( .A(w_mem_inst__abc_21203_new_n5272_), .B(w_mem_inst__abc_21203_new_n5268_), .Y(w_mem_inst__0w_mem_5__31_0__0_));
OR2X2 OR2X2_3281 ( .A(w_mem_inst__abc_21203_new_n5277_), .B(w_mem_inst__abc_21203_new_n5275_), .Y(w_mem_inst__abc_21203_new_n5278_));
OR2X2 OR2X2_3282 ( .A(w_mem_inst__abc_21203_new_n5278_), .B(w_mem_inst__abc_21203_new_n5274_), .Y(w_mem_inst__0w_mem_5__31_0__1_));
OR2X2 OR2X2_3283 ( .A(w_mem_inst__abc_21203_new_n5283_), .B(w_mem_inst__abc_21203_new_n5281_), .Y(w_mem_inst__abc_21203_new_n5284_));
OR2X2 OR2X2_3284 ( .A(w_mem_inst__abc_21203_new_n5284_), .B(w_mem_inst__abc_21203_new_n5280_), .Y(w_mem_inst__0w_mem_5__31_0__2_));
OR2X2 OR2X2_3285 ( .A(w_mem_inst__abc_21203_new_n5289_), .B(w_mem_inst__abc_21203_new_n5287_), .Y(w_mem_inst__abc_21203_new_n5290_));
OR2X2 OR2X2_3286 ( .A(w_mem_inst__abc_21203_new_n5290_), .B(w_mem_inst__abc_21203_new_n5286_), .Y(w_mem_inst__0w_mem_5__31_0__3_));
OR2X2 OR2X2_3287 ( .A(w_mem_inst__abc_21203_new_n5295_), .B(w_mem_inst__abc_21203_new_n5293_), .Y(w_mem_inst__abc_21203_new_n5296_));
OR2X2 OR2X2_3288 ( .A(w_mem_inst__abc_21203_new_n5296_), .B(w_mem_inst__abc_21203_new_n5292_), .Y(w_mem_inst__0w_mem_5__31_0__4_));
OR2X2 OR2X2_3289 ( .A(w_mem_inst__abc_21203_new_n5301_), .B(w_mem_inst__abc_21203_new_n5299_), .Y(w_mem_inst__abc_21203_new_n5302_));
OR2X2 OR2X2_329 ( .A(_abc_15497_new_n1717_), .B(_abc_15497_new_n1703_), .Y(_0H3_reg_31_0__13_));
OR2X2 OR2X2_3290 ( .A(w_mem_inst__abc_21203_new_n5302_), .B(w_mem_inst__abc_21203_new_n5298_), .Y(w_mem_inst__0w_mem_5__31_0__5_));
OR2X2 OR2X2_3291 ( .A(w_mem_inst__abc_21203_new_n5307_), .B(w_mem_inst__abc_21203_new_n5305_), .Y(w_mem_inst__abc_21203_new_n5308_));
OR2X2 OR2X2_3292 ( .A(w_mem_inst__abc_21203_new_n5308_), .B(w_mem_inst__abc_21203_new_n5304_), .Y(w_mem_inst__0w_mem_5__31_0__6_));
OR2X2 OR2X2_3293 ( .A(w_mem_inst__abc_21203_new_n5313_), .B(w_mem_inst__abc_21203_new_n5311_), .Y(w_mem_inst__abc_21203_new_n5314_));
OR2X2 OR2X2_3294 ( .A(w_mem_inst__abc_21203_new_n5314_), .B(w_mem_inst__abc_21203_new_n5310_), .Y(w_mem_inst__0w_mem_5__31_0__7_));
OR2X2 OR2X2_3295 ( .A(w_mem_inst__abc_21203_new_n5319_), .B(w_mem_inst__abc_21203_new_n5317_), .Y(w_mem_inst__abc_21203_new_n5320_));
OR2X2 OR2X2_3296 ( .A(w_mem_inst__abc_21203_new_n5320_), .B(w_mem_inst__abc_21203_new_n5316_), .Y(w_mem_inst__0w_mem_5__31_0__8_));
OR2X2 OR2X2_3297 ( .A(w_mem_inst__abc_21203_new_n5325_), .B(w_mem_inst__abc_21203_new_n5323_), .Y(w_mem_inst__abc_21203_new_n5326_));
OR2X2 OR2X2_3298 ( .A(w_mem_inst__abc_21203_new_n5326_), .B(w_mem_inst__abc_21203_new_n5322_), .Y(w_mem_inst__0w_mem_5__31_0__9_));
OR2X2 OR2X2_3299 ( .A(w_mem_inst__abc_21203_new_n5331_), .B(w_mem_inst__abc_21203_new_n5329_), .Y(w_mem_inst__abc_21203_new_n5332_));
OR2X2 OR2X2_33 ( .A(c_reg_2_), .B(\digest[66] ), .Y(_abc_15497_new_n826_));
OR2X2 OR2X2_330 ( .A(\digest[46] ), .B(d_reg_14_), .Y(_abc_15497_new_n1722_));
OR2X2 OR2X2_3300 ( .A(w_mem_inst__abc_21203_new_n5332_), .B(w_mem_inst__abc_21203_new_n5328_), .Y(w_mem_inst__0w_mem_5__31_0__10_));
OR2X2 OR2X2_3301 ( .A(w_mem_inst__abc_21203_new_n5337_), .B(w_mem_inst__abc_21203_new_n5335_), .Y(w_mem_inst__abc_21203_new_n5338_));
OR2X2 OR2X2_3302 ( .A(w_mem_inst__abc_21203_new_n5338_), .B(w_mem_inst__abc_21203_new_n5334_), .Y(w_mem_inst__0w_mem_5__31_0__11_));
OR2X2 OR2X2_3303 ( .A(w_mem_inst__abc_21203_new_n5343_), .B(w_mem_inst__abc_21203_new_n5341_), .Y(w_mem_inst__abc_21203_new_n5344_));
OR2X2 OR2X2_3304 ( .A(w_mem_inst__abc_21203_new_n5344_), .B(w_mem_inst__abc_21203_new_n5340_), .Y(w_mem_inst__0w_mem_5__31_0__12_));
OR2X2 OR2X2_3305 ( .A(w_mem_inst__abc_21203_new_n5349_), .B(w_mem_inst__abc_21203_new_n5347_), .Y(w_mem_inst__abc_21203_new_n5350_));
OR2X2 OR2X2_3306 ( .A(w_mem_inst__abc_21203_new_n5350_), .B(w_mem_inst__abc_21203_new_n5346_), .Y(w_mem_inst__0w_mem_5__31_0__13_));
OR2X2 OR2X2_3307 ( .A(w_mem_inst__abc_21203_new_n5355_), .B(w_mem_inst__abc_21203_new_n5353_), .Y(w_mem_inst__abc_21203_new_n5356_));
OR2X2 OR2X2_3308 ( .A(w_mem_inst__abc_21203_new_n5356_), .B(w_mem_inst__abc_21203_new_n5352_), .Y(w_mem_inst__0w_mem_5__31_0__14_));
OR2X2 OR2X2_3309 ( .A(w_mem_inst__abc_21203_new_n5361_), .B(w_mem_inst__abc_21203_new_n5359_), .Y(w_mem_inst__abc_21203_new_n5362_));
OR2X2 OR2X2_331 ( .A(_abc_15497_new_n1721_), .B(_abc_15497_new_n1725_), .Y(_abc_15497_new_n1726_));
OR2X2 OR2X2_3310 ( .A(w_mem_inst__abc_21203_new_n5362_), .B(w_mem_inst__abc_21203_new_n5358_), .Y(w_mem_inst__0w_mem_5__31_0__15_));
OR2X2 OR2X2_3311 ( .A(w_mem_inst__abc_21203_new_n5367_), .B(w_mem_inst__abc_21203_new_n5365_), .Y(w_mem_inst__abc_21203_new_n5368_));
OR2X2 OR2X2_3312 ( .A(w_mem_inst__abc_21203_new_n5368_), .B(w_mem_inst__abc_21203_new_n5364_), .Y(w_mem_inst__0w_mem_5__31_0__16_));
OR2X2 OR2X2_3313 ( .A(w_mem_inst__abc_21203_new_n5373_), .B(w_mem_inst__abc_21203_new_n5371_), .Y(w_mem_inst__abc_21203_new_n5374_));
OR2X2 OR2X2_3314 ( .A(w_mem_inst__abc_21203_new_n5374_), .B(w_mem_inst__abc_21203_new_n5370_), .Y(w_mem_inst__0w_mem_5__31_0__17_));
OR2X2 OR2X2_3315 ( .A(w_mem_inst__abc_21203_new_n5379_), .B(w_mem_inst__abc_21203_new_n5377_), .Y(w_mem_inst__abc_21203_new_n5380_));
OR2X2 OR2X2_3316 ( .A(w_mem_inst__abc_21203_new_n5380_), .B(w_mem_inst__abc_21203_new_n5376_), .Y(w_mem_inst__0w_mem_5__31_0__18_));
OR2X2 OR2X2_3317 ( .A(w_mem_inst__abc_21203_new_n5385_), .B(w_mem_inst__abc_21203_new_n5383_), .Y(w_mem_inst__abc_21203_new_n5386_));
OR2X2 OR2X2_3318 ( .A(w_mem_inst__abc_21203_new_n5386_), .B(w_mem_inst__abc_21203_new_n5382_), .Y(w_mem_inst__0w_mem_5__31_0__19_));
OR2X2 OR2X2_3319 ( .A(w_mem_inst__abc_21203_new_n5391_), .B(w_mem_inst__abc_21203_new_n5389_), .Y(w_mem_inst__abc_21203_new_n5392_));
OR2X2 OR2X2_332 ( .A(_abc_15497_new_n699_), .B(\digest[46] ), .Y(_abc_15497_new_n1731_));
OR2X2 OR2X2_3320 ( .A(w_mem_inst__abc_21203_new_n5392_), .B(w_mem_inst__abc_21203_new_n5388_), .Y(w_mem_inst__0w_mem_5__31_0__20_));
OR2X2 OR2X2_3321 ( .A(w_mem_inst__abc_21203_new_n5397_), .B(w_mem_inst__abc_21203_new_n5395_), .Y(w_mem_inst__abc_21203_new_n5398_));
OR2X2 OR2X2_3322 ( .A(w_mem_inst__abc_21203_new_n5398_), .B(w_mem_inst__abc_21203_new_n5394_), .Y(w_mem_inst__0w_mem_5__31_0__21_));
OR2X2 OR2X2_3323 ( .A(w_mem_inst__abc_21203_new_n5403_), .B(w_mem_inst__abc_21203_new_n5401_), .Y(w_mem_inst__abc_21203_new_n5404_));
OR2X2 OR2X2_3324 ( .A(w_mem_inst__abc_21203_new_n5404_), .B(w_mem_inst__abc_21203_new_n5400_), .Y(w_mem_inst__0w_mem_5__31_0__22_));
OR2X2 OR2X2_3325 ( .A(w_mem_inst__abc_21203_new_n5409_), .B(w_mem_inst__abc_21203_new_n5407_), .Y(w_mem_inst__abc_21203_new_n5410_));
OR2X2 OR2X2_3326 ( .A(w_mem_inst__abc_21203_new_n5410_), .B(w_mem_inst__abc_21203_new_n5406_), .Y(w_mem_inst__0w_mem_5__31_0__23_));
OR2X2 OR2X2_3327 ( .A(w_mem_inst__abc_21203_new_n5415_), .B(w_mem_inst__abc_21203_new_n5413_), .Y(w_mem_inst__abc_21203_new_n5416_));
OR2X2 OR2X2_3328 ( .A(w_mem_inst__abc_21203_new_n5416_), .B(w_mem_inst__abc_21203_new_n5412_), .Y(w_mem_inst__0w_mem_5__31_0__24_));
OR2X2 OR2X2_3329 ( .A(w_mem_inst__abc_21203_new_n5421_), .B(w_mem_inst__abc_21203_new_n5419_), .Y(w_mem_inst__abc_21203_new_n5422_));
OR2X2 OR2X2_333 ( .A(_abc_15497_new_n1730_), .B(_abc_15497_new_n1732_), .Y(_0H3_reg_31_0__14_));
OR2X2 OR2X2_3330 ( .A(w_mem_inst__abc_21203_new_n5422_), .B(w_mem_inst__abc_21203_new_n5418_), .Y(w_mem_inst__0w_mem_5__31_0__25_));
OR2X2 OR2X2_3331 ( .A(w_mem_inst__abc_21203_new_n5427_), .B(w_mem_inst__abc_21203_new_n5425_), .Y(w_mem_inst__abc_21203_new_n5428_));
OR2X2 OR2X2_3332 ( .A(w_mem_inst__abc_21203_new_n5428_), .B(w_mem_inst__abc_21203_new_n5424_), .Y(w_mem_inst__0w_mem_5__31_0__26_));
OR2X2 OR2X2_3333 ( .A(w_mem_inst__abc_21203_new_n5433_), .B(w_mem_inst__abc_21203_new_n5431_), .Y(w_mem_inst__abc_21203_new_n5434_));
OR2X2 OR2X2_3334 ( .A(w_mem_inst__abc_21203_new_n5434_), .B(w_mem_inst__abc_21203_new_n5430_), .Y(w_mem_inst__0w_mem_5__31_0__27_));
OR2X2 OR2X2_3335 ( .A(w_mem_inst__abc_21203_new_n5439_), .B(w_mem_inst__abc_21203_new_n5437_), .Y(w_mem_inst__abc_21203_new_n5440_));
OR2X2 OR2X2_3336 ( .A(w_mem_inst__abc_21203_new_n5440_), .B(w_mem_inst__abc_21203_new_n5436_), .Y(w_mem_inst__0w_mem_5__31_0__28_));
OR2X2 OR2X2_3337 ( .A(w_mem_inst__abc_21203_new_n5445_), .B(w_mem_inst__abc_21203_new_n5443_), .Y(w_mem_inst__abc_21203_new_n5446_));
OR2X2 OR2X2_3338 ( .A(w_mem_inst__abc_21203_new_n5446_), .B(w_mem_inst__abc_21203_new_n5442_), .Y(w_mem_inst__0w_mem_5__31_0__29_));
OR2X2 OR2X2_3339 ( .A(w_mem_inst__abc_21203_new_n5451_), .B(w_mem_inst__abc_21203_new_n5449_), .Y(w_mem_inst__abc_21203_new_n5452_));
OR2X2 OR2X2_334 ( .A(\digest[47] ), .B(d_reg_15_), .Y(_abc_15497_new_n1737_));
OR2X2 OR2X2_3340 ( .A(w_mem_inst__abc_21203_new_n5452_), .B(w_mem_inst__abc_21203_new_n5448_), .Y(w_mem_inst__0w_mem_5__31_0__30_));
OR2X2 OR2X2_3341 ( .A(w_mem_inst__abc_21203_new_n5457_), .B(w_mem_inst__abc_21203_new_n5455_), .Y(w_mem_inst__abc_21203_new_n5458_));
OR2X2 OR2X2_3342 ( .A(w_mem_inst__abc_21203_new_n5458_), .B(w_mem_inst__abc_21203_new_n5454_), .Y(w_mem_inst__0w_mem_5__31_0__31_));
OR2X2 OR2X2_3343 ( .A(w_mem_inst__abc_21203_new_n5463_), .B(w_mem_inst__abc_21203_new_n5461_), .Y(w_mem_inst__abc_21203_new_n5464_));
OR2X2 OR2X2_3344 ( .A(w_mem_inst__abc_21203_new_n5464_), .B(w_mem_inst__abc_21203_new_n5460_), .Y(w_mem_inst__0w_mem_1__31_0__0_));
OR2X2 OR2X2_3345 ( .A(w_mem_inst__abc_21203_new_n5469_), .B(w_mem_inst__abc_21203_new_n5467_), .Y(w_mem_inst__abc_21203_new_n5470_));
OR2X2 OR2X2_3346 ( .A(w_mem_inst__abc_21203_new_n5470_), .B(w_mem_inst__abc_21203_new_n5466_), .Y(w_mem_inst__0w_mem_1__31_0__1_));
OR2X2 OR2X2_3347 ( .A(w_mem_inst__abc_21203_new_n5475_), .B(w_mem_inst__abc_21203_new_n5473_), .Y(w_mem_inst__abc_21203_new_n5476_));
OR2X2 OR2X2_3348 ( .A(w_mem_inst__abc_21203_new_n5476_), .B(w_mem_inst__abc_21203_new_n5472_), .Y(w_mem_inst__0w_mem_1__31_0__2_));
OR2X2 OR2X2_3349 ( .A(w_mem_inst__abc_21203_new_n5481_), .B(w_mem_inst__abc_21203_new_n5479_), .Y(w_mem_inst__abc_21203_new_n5482_));
OR2X2 OR2X2_335 ( .A(_abc_15497_new_n1736_), .B(_abc_15497_new_n1740_), .Y(_abc_15497_new_n1741_));
OR2X2 OR2X2_3350 ( .A(w_mem_inst__abc_21203_new_n5482_), .B(w_mem_inst__abc_21203_new_n5478_), .Y(w_mem_inst__0w_mem_1__31_0__3_));
OR2X2 OR2X2_3351 ( .A(w_mem_inst__abc_21203_new_n5487_), .B(w_mem_inst__abc_21203_new_n5485_), .Y(w_mem_inst__abc_21203_new_n5488_));
OR2X2 OR2X2_3352 ( .A(w_mem_inst__abc_21203_new_n5488_), .B(w_mem_inst__abc_21203_new_n5484_), .Y(w_mem_inst__0w_mem_1__31_0__4_));
OR2X2 OR2X2_3353 ( .A(w_mem_inst__abc_21203_new_n5493_), .B(w_mem_inst__abc_21203_new_n5491_), .Y(w_mem_inst__abc_21203_new_n5494_));
OR2X2 OR2X2_3354 ( .A(w_mem_inst__abc_21203_new_n5494_), .B(w_mem_inst__abc_21203_new_n5490_), .Y(w_mem_inst__0w_mem_1__31_0__5_));
OR2X2 OR2X2_3355 ( .A(w_mem_inst__abc_21203_new_n5499_), .B(w_mem_inst__abc_21203_new_n5497_), .Y(w_mem_inst__abc_21203_new_n5500_));
OR2X2 OR2X2_3356 ( .A(w_mem_inst__abc_21203_new_n5500_), .B(w_mem_inst__abc_21203_new_n5496_), .Y(w_mem_inst__0w_mem_1__31_0__6_));
OR2X2 OR2X2_3357 ( .A(w_mem_inst__abc_21203_new_n5505_), .B(w_mem_inst__abc_21203_new_n5503_), .Y(w_mem_inst__abc_21203_new_n5506_));
OR2X2 OR2X2_3358 ( .A(w_mem_inst__abc_21203_new_n5506_), .B(w_mem_inst__abc_21203_new_n5502_), .Y(w_mem_inst__0w_mem_1__31_0__7_));
OR2X2 OR2X2_3359 ( .A(w_mem_inst__abc_21203_new_n5511_), .B(w_mem_inst__abc_21203_new_n5509_), .Y(w_mem_inst__abc_21203_new_n5512_));
OR2X2 OR2X2_336 ( .A(_abc_15497_new_n1735_), .B(_abc_15497_new_n1742_), .Y(_abc_15497_new_n1743_));
OR2X2 OR2X2_3360 ( .A(w_mem_inst__abc_21203_new_n5512_), .B(w_mem_inst__abc_21203_new_n5508_), .Y(w_mem_inst__0w_mem_1__31_0__8_));
OR2X2 OR2X2_3361 ( .A(w_mem_inst__abc_21203_new_n5517_), .B(w_mem_inst__abc_21203_new_n5515_), .Y(w_mem_inst__abc_21203_new_n5518_));
OR2X2 OR2X2_3362 ( .A(w_mem_inst__abc_21203_new_n5518_), .B(w_mem_inst__abc_21203_new_n5514_), .Y(w_mem_inst__0w_mem_1__31_0__9_));
OR2X2 OR2X2_3363 ( .A(w_mem_inst__abc_21203_new_n5523_), .B(w_mem_inst__abc_21203_new_n5521_), .Y(w_mem_inst__abc_21203_new_n5524_));
OR2X2 OR2X2_3364 ( .A(w_mem_inst__abc_21203_new_n5524_), .B(w_mem_inst__abc_21203_new_n5520_), .Y(w_mem_inst__0w_mem_1__31_0__10_));
OR2X2 OR2X2_3365 ( .A(w_mem_inst__abc_21203_new_n5529_), .B(w_mem_inst__abc_21203_new_n5527_), .Y(w_mem_inst__abc_21203_new_n5530_));
OR2X2 OR2X2_3366 ( .A(w_mem_inst__abc_21203_new_n5530_), .B(w_mem_inst__abc_21203_new_n5526_), .Y(w_mem_inst__0w_mem_1__31_0__11_));
OR2X2 OR2X2_3367 ( .A(w_mem_inst__abc_21203_new_n5535_), .B(w_mem_inst__abc_21203_new_n5533_), .Y(w_mem_inst__abc_21203_new_n5536_));
OR2X2 OR2X2_3368 ( .A(w_mem_inst__abc_21203_new_n5536_), .B(w_mem_inst__abc_21203_new_n5532_), .Y(w_mem_inst__0w_mem_1__31_0__12_));
OR2X2 OR2X2_3369 ( .A(w_mem_inst__abc_21203_new_n5541_), .B(w_mem_inst__abc_21203_new_n5539_), .Y(w_mem_inst__abc_21203_new_n5542_));
OR2X2 OR2X2_337 ( .A(_abc_15497_new_n1745_), .B(_abc_15497_new_n1734_), .Y(_0H3_reg_31_0__15_));
OR2X2 OR2X2_3370 ( .A(w_mem_inst__abc_21203_new_n5542_), .B(w_mem_inst__abc_21203_new_n5538_), .Y(w_mem_inst__0w_mem_1__31_0__13_));
OR2X2 OR2X2_3371 ( .A(w_mem_inst__abc_21203_new_n5547_), .B(w_mem_inst__abc_21203_new_n5545_), .Y(w_mem_inst__abc_21203_new_n5548_));
OR2X2 OR2X2_3372 ( .A(w_mem_inst__abc_21203_new_n5548_), .B(w_mem_inst__abc_21203_new_n5544_), .Y(w_mem_inst__0w_mem_1__31_0__14_));
OR2X2 OR2X2_3373 ( .A(w_mem_inst__abc_21203_new_n5553_), .B(w_mem_inst__abc_21203_new_n5551_), .Y(w_mem_inst__abc_21203_new_n5554_));
OR2X2 OR2X2_3374 ( .A(w_mem_inst__abc_21203_new_n5554_), .B(w_mem_inst__abc_21203_new_n5550_), .Y(w_mem_inst__0w_mem_1__31_0__15_));
OR2X2 OR2X2_3375 ( .A(w_mem_inst__abc_21203_new_n5559_), .B(w_mem_inst__abc_21203_new_n5557_), .Y(w_mem_inst__abc_21203_new_n5560_));
OR2X2 OR2X2_3376 ( .A(w_mem_inst__abc_21203_new_n5560_), .B(w_mem_inst__abc_21203_new_n5556_), .Y(w_mem_inst__0w_mem_1__31_0__16_));
OR2X2 OR2X2_3377 ( .A(w_mem_inst__abc_21203_new_n5565_), .B(w_mem_inst__abc_21203_new_n5563_), .Y(w_mem_inst__abc_21203_new_n5566_));
OR2X2 OR2X2_3378 ( .A(w_mem_inst__abc_21203_new_n5566_), .B(w_mem_inst__abc_21203_new_n5562_), .Y(w_mem_inst__0w_mem_1__31_0__17_));
OR2X2 OR2X2_3379 ( .A(w_mem_inst__abc_21203_new_n5571_), .B(w_mem_inst__abc_21203_new_n5569_), .Y(w_mem_inst__abc_21203_new_n5572_));
OR2X2 OR2X2_338 ( .A(_abc_15497_new_n1719_), .B(_abc_15497_new_n1749_), .Y(_abc_15497_new_n1750_));
OR2X2 OR2X2_3380 ( .A(w_mem_inst__abc_21203_new_n5572_), .B(w_mem_inst__abc_21203_new_n5568_), .Y(w_mem_inst__0w_mem_1__31_0__18_));
OR2X2 OR2X2_3381 ( .A(w_mem_inst__abc_21203_new_n5577_), .B(w_mem_inst__abc_21203_new_n5575_), .Y(w_mem_inst__abc_21203_new_n5578_));
OR2X2 OR2X2_3382 ( .A(w_mem_inst__abc_21203_new_n5578_), .B(w_mem_inst__abc_21203_new_n5574_), .Y(w_mem_inst__0w_mem_1__31_0__19_));
OR2X2 OR2X2_3383 ( .A(w_mem_inst__abc_21203_new_n5583_), .B(w_mem_inst__abc_21203_new_n5581_), .Y(w_mem_inst__abc_21203_new_n5584_));
OR2X2 OR2X2_3384 ( .A(w_mem_inst__abc_21203_new_n5584_), .B(w_mem_inst__abc_21203_new_n5580_), .Y(w_mem_inst__0w_mem_1__31_0__20_));
OR2X2 OR2X2_3385 ( .A(w_mem_inst__abc_21203_new_n5589_), .B(w_mem_inst__abc_21203_new_n5587_), .Y(w_mem_inst__abc_21203_new_n5590_));
OR2X2 OR2X2_3386 ( .A(w_mem_inst__abc_21203_new_n5590_), .B(w_mem_inst__abc_21203_new_n5586_), .Y(w_mem_inst__0w_mem_1__31_0__21_));
OR2X2 OR2X2_3387 ( .A(w_mem_inst__abc_21203_new_n5595_), .B(w_mem_inst__abc_21203_new_n5593_), .Y(w_mem_inst__abc_21203_new_n5596_));
OR2X2 OR2X2_3388 ( .A(w_mem_inst__abc_21203_new_n5596_), .B(w_mem_inst__abc_21203_new_n5592_), .Y(w_mem_inst__0w_mem_1__31_0__22_));
OR2X2 OR2X2_3389 ( .A(w_mem_inst__abc_21203_new_n5601_), .B(w_mem_inst__abc_21203_new_n5599_), .Y(w_mem_inst__abc_21203_new_n5602_));
OR2X2 OR2X2_339 ( .A(_abc_15497_new_n1751_), .B(_abc_15497_new_n1738_), .Y(_abc_15497_new_n1752_));
OR2X2 OR2X2_3390 ( .A(w_mem_inst__abc_21203_new_n5602_), .B(w_mem_inst__abc_21203_new_n5598_), .Y(w_mem_inst__0w_mem_1__31_0__23_));
OR2X2 OR2X2_3391 ( .A(w_mem_inst__abc_21203_new_n5607_), .B(w_mem_inst__abc_21203_new_n5605_), .Y(w_mem_inst__abc_21203_new_n5608_));
OR2X2 OR2X2_3392 ( .A(w_mem_inst__abc_21203_new_n5608_), .B(w_mem_inst__abc_21203_new_n5604_), .Y(w_mem_inst__0w_mem_1__31_0__24_));
OR2X2 OR2X2_3393 ( .A(w_mem_inst__abc_21203_new_n5613_), .B(w_mem_inst__abc_21203_new_n5611_), .Y(w_mem_inst__abc_21203_new_n5614_));
OR2X2 OR2X2_3394 ( .A(w_mem_inst__abc_21203_new_n5614_), .B(w_mem_inst__abc_21203_new_n5610_), .Y(w_mem_inst__0w_mem_1__31_0__25_));
OR2X2 OR2X2_3395 ( .A(w_mem_inst__abc_21203_new_n5619_), .B(w_mem_inst__abc_21203_new_n5617_), .Y(w_mem_inst__abc_21203_new_n5620_));
OR2X2 OR2X2_3396 ( .A(w_mem_inst__abc_21203_new_n5620_), .B(w_mem_inst__abc_21203_new_n5616_), .Y(w_mem_inst__0w_mem_1__31_0__26_));
OR2X2 OR2X2_3397 ( .A(w_mem_inst__abc_21203_new_n5625_), .B(w_mem_inst__abc_21203_new_n5623_), .Y(w_mem_inst__abc_21203_new_n5626_));
OR2X2 OR2X2_3398 ( .A(w_mem_inst__abc_21203_new_n5626_), .B(w_mem_inst__abc_21203_new_n5622_), .Y(w_mem_inst__0w_mem_1__31_0__27_));
OR2X2 OR2X2_3399 ( .A(w_mem_inst__abc_21203_new_n5631_), .B(w_mem_inst__abc_21203_new_n5629_), .Y(w_mem_inst__abc_21203_new_n5632_));
OR2X2 OR2X2_34 ( .A(_abc_15497_new_n828_), .B(_abc_15497_new_n817_), .Y(_abc_15497_new_n829_));
OR2X2 OR2X2_340 ( .A(_abc_15497_new_n1757_), .B(_abc_15497_new_n1755_), .Y(_abc_15497_new_n1758_));
OR2X2 OR2X2_3400 ( .A(w_mem_inst__abc_21203_new_n5632_), .B(w_mem_inst__abc_21203_new_n5628_), .Y(w_mem_inst__0w_mem_1__31_0__28_));
OR2X2 OR2X2_3401 ( .A(w_mem_inst__abc_21203_new_n5637_), .B(w_mem_inst__abc_21203_new_n5635_), .Y(w_mem_inst__abc_21203_new_n5638_));
OR2X2 OR2X2_3402 ( .A(w_mem_inst__abc_21203_new_n5638_), .B(w_mem_inst__abc_21203_new_n5634_), .Y(w_mem_inst__0w_mem_1__31_0__29_));
OR2X2 OR2X2_3403 ( .A(w_mem_inst__abc_21203_new_n5643_), .B(w_mem_inst__abc_21203_new_n5641_), .Y(w_mem_inst__abc_21203_new_n5644_));
OR2X2 OR2X2_3404 ( .A(w_mem_inst__abc_21203_new_n5644_), .B(w_mem_inst__abc_21203_new_n5640_), .Y(w_mem_inst__0w_mem_1__31_0__30_));
OR2X2 OR2X2_3405 ( .A(w_mem_inst__abc_21203_new_n5649_), .B(w_mem_inst__abc_21203_new_n5647_), .Y(w_mem_inst__abc_21203_new_n5650_));
OR2X2 OR2X2_3406 ( .A(w_mem_inst__abc_21203_new_n5650_), .B(w_mem_inst__abc_21203_new_n5646_), .Y(w_mem_inst__0w_mem_1__31_0__31_));
OR2X2 OR2X2_3407 ( .A(w_mem_inst__abc_21203_new_n5655_), .B(w_mem_inst__abc_21203_new_n5653_), .Y(w_mem_inst__abc_21203_new_n5656_));
OR2X2 OR2X2_3408 ( .A(w_mem_inst__abc_21203_new_n5656_), .B(w_mem_inst__abc_21203_new_n5652_), .Y(w_mem_inst__0w_mem_3__31_0__0_));
OR2X2 OR2X2_3409 ( .A(w_mem_inst__abc_21203_new_n5661_), .B(w_mem_inst__abc_21203_new_n5659_), .Y(w_mem_inst__abc_21203_new_n5662_));
OR2X2 OR2X2_341 ( .A(\digest[48] ), .B(d_reg_16_), .Y(_abc_15497_new_n1759_));
OR2X2 OR2X2_3410 ( .A(w_mem_inst__abc_21203_new_n5662_), .B(w_mem_inst__abc_21203_new_n5658_), .Y(w_mem_inst__0w_mem_3__31_0__1_));
OR2X2 OR2X2_3411 ( .A(w_mem_inst__abc_21203_new_n5667_), .B(w_mem_inst__abc_21203_new_n5665_), .Y(w_mem_inst__abc_21203_new_n5668_));
OR2X2 OR2X2_3412 ( .A(w_mem_inst__abc_21203_new_n5668_), .B(w_mem_inst__abc_21203_new_n5664_), .Y(w_mem_inst__0w_mem_3__31_0__2_));
OR2X2 OR2X2_3413 ( .A(w_mem_inst__abc_21203_new_n5673_), .B(w_mem_inst__abc_21203_new_n5671_), .Y(w_mem_inst__abc_21203_new_n5674_));
OR2X2 OR2X2_3414 ( .A(w_mem_inst__abc_21203_new_n5674_), .B(w_mem_inst__abc_21203_new_n5670_), .Y(w_mem_inst__0w_mem_3__31_0__3_));
OR2X2 OR2X2_3415 ( .A(w_mem_inst__abc_21203_new_n5679_), .B(w_mem_inst__abc_21203_new_n5677_), .Y(w_mem_inst__abc_21203_new_n5680_));
OR2X2 OR2X2_3416 ( .A(w_mem_inst__abc_21203_new_n5680_), .B(w_mem_inst__abc_21203_new_n5676_), .Y(w_mem_inst__0w_mem_3__31_0__4_));
OR2X2 OR2X2_3417 ( .A(w_mem_inst__abc_21203_new_n5685_), .B(w_mem_inst__abc_21203_new_n5683_), .Y(w_mem_inst__abc_21203_new_n5686_));
OR2X2 OR2X2_3418 ( .A(w_mem_inst__abc_21203_new_n5686_), .B(w_mem_inst__abc_21203_new_n5682_), .Y(w_mem_inst__0w_mem_3__31_0__5_));
OR2X2 OR2X2_3419 ( .A(w_mem_inst__abc_21203_new_n5691_), .B(w_mem_inst__abc_21203_new_n5689_), .Y(w_mem_inst__abc_21203_new_n5692_));
OR2X2 OR2X2_342 ( .A(_abc_15497_new_n1758_), .B(_abc_15497_new_n1762_), .Y(_abc_15497_new_n1763_));
OR2X2 OR2X2_3420 ( .A(w_mem_inst__abc_21203_new_n5692_), .B(w_mem_inst__abc_21203_new_n5688_), .Y(w_mem_inst__0w_mem_3__31_0__6_));
OR2X2 OR2X2_3421 ( .A(w_mem_inst__abc_21203_new_n5697_), .B(w_mem_inst__abc_21203_new_n5695_), .Y(w_mem_inst__abc_21203_new_n5698_));
OR2X2 OR2X2_3422 ( .A(w_mem_inst__abc_21203_new_n5698_), .B(w_mem_inst__abc_21203_new_n5694_), .Y(w_mem_inst__0w_mem_3__31_0__7_));
OR2X2 OR2X2_3423 ( .A(w_mem_inst__abc_21203_new_n5703_), .B(w_mem_inst__abc_21203_new_n5701_), .Y(w_mem_inst__abc_21203_new_n5704_));
OR2X2 OR2X2_3424 ( .A(w_mem_inst__abc_21203_new_n5704_), .B(w_mem_inst__abc_21203_new_n5700_), .Y(w_mem_inst__0w_mem_3__31_0__8_));
OR2X2 OR2X2_3425 ( .A(w_mem_inst__abc_21203_new_n5709_), .B(w_mem_inst__abc_21203_new_n5707_), .Y(w_mem_inst__abc_21203_new_n5710_));
OR2X2 OR2X2_3426 ( .A(w_mem_inst__abc_21203_new_n5710_), .B(w_mem_inst__abc_21203_new_n5706_), .Y(w_mem_inst__0w_mem_3__31_0__9_));
OR2X2 OR2X2_3427 ( .A(w_mem_inst__abc_21203_new_n5715_), .B(w_mem_inst__abc_21203_new_n5713_), .Y(w_mem_inst__abc_21203_new_n5716_));
OR2X2 OR2X2_3428 ( .A(w_mem_inst__abc_21203_new_n5716_), .B(w_mem_inst__abc_21203_new_n5712_), .Y(w_mem_inst__0w_mem_3__31_0__10_));
OR2X2 OR2X2_3429 ( .A(w_mem_inst__abc_21203_new_n5721_), .B(w_mem_inst__abc_21203_new_n5719_), .Y(w_mem_inst__abc_21203_new_n5722_));
OR2X2 OR2X2_343 ( .A(_abc_15497_new_n1767_), .B(_abc_15497_new_n1747_), .Y(_0H3_reg_31_0__16_));
OR2X2 OR2X2_3430 ( .A(w_mem_inst__abc_21203_new_n5722_), .B(w_mem_inst__abc_21203_new_n5718_), .Y(w_mem_inst__0w_mem_3__31_0__11_));
OR2X2 OR2X2_3431 ( .A(w_mem_inst__abc_21203_new_n5727_), .B(w_mem_inst__abc_21203_new_n5725_), .Y(w_mem_inst__abc_21203_new_n5728_));
OR2X2 OR2X2_3432 ( .A(w_mem_inst__abc_21203_new_n5728_), .B(w_mem_inst__abc_21203_new_n5724_), .Y(w_mem_inst__0w_mem_3__31_0__12_));
OR2X2 OR2X2_3433 ( .A(w_mem_inst__abc_21203_new_n5733_), .B(w_mem_inst__abc_21203_new_n5731_), .Y(w_mem_inst__abc_21203_new_n5734_));
OR2X2 OR2X2_3434 ( .A(w_mem_inst__abc_21203_new_n5734_), .B(w_mem_inst__abc_21203_new_n5730_), .Y(w_mem_inst__0w_mem_3__31_0__13_));
OR2X2 OR2X2_3435 ( .A(w_mem_inst__abc_21203_new_n5739_), .B(w_mem_inst__abc_21203_new_n5737_), .Y(w_mem_inst__abc_21203_new_n5740_));
OR2X2 OR2X2_3436 ( .A(w_mem_inst__abc_21203_new_n5740_), .B(w_mem_inst__abc_21203_new_n5736_), .Y(w_mem_inst__0w_mem_3__31_0__14_));
OR2X2 OR2X2_3437 ( .A(w_mem_inst__abc_21203_new_n5745_), .B(w_mem_inst__abc_21203_new_n5743_), .Y(w_mem_inst__abc_21203_new_n5746_));
OR2X2 OR2X2_3438 ( .A(w_mem_inst__abc_21203_new_n5746_), .B(w_mem_inst__abc_21203_new_n5742_), .Y(w_mem_inst__0w_mem_3__31_0__15_));
OR2X2 OR2X2_3439 ( .A(w_mem_inst__abc_21203_new_n5751_), .B(w_mem_inst__abc_21203_new_n5749_), .Y(w_mem_inst__abc_21203_new_n5752_));
OR2X2 OR2X2_344 ( .A(\digest[49] ), .B(d_reg_17_), .Y(_abc_15497_new_n1770_));
OR2X2 OR2X2_3440 ( .A(w_mem_inst__abc_21203_new_n5752_), .B(w_mem_inst__abc_21203_new_n5748_), .Y(w_mem_inst__0w_mem_3__31_0__16_));
OR2X2 OR2X2_3441 ( .A(w_mem_inst__abc_21203_new_n5757_), .B(w_mem_inst__abc_21203_new_n5755_), .Y(w_mem_inst__abc_21203_new_n5758_));
OR2X2 OR2X2_3442 ( .A(w_mem_inst__abc_21203_new_n5758_), .B(w_mem_inst__abc_21203_new_n5754_), .Y(w_mem_inst__0w_mem_3__31_0__17_));
OR2X2 OR2X2_3443 ( .A(w_mem_inst__abc_21203_new_n5763_), .B(w_mem_inst__abc_21203_new_n5761_), .Y(w_mem_inst__abc_21203_new_n5764_));
OR2X2 OR2X2_3444 ( .A(w_mem_inst__abc_21203_new_n5764_), .B(w_mem_inst__abc_21203_new_n5760_), .Y(w_mem_inst__0w_mem_3__31_0__18_));
OR2X2 OR2X2_3445 ( .A(w_mem_inst__abc_21203_new_n5769_), .B(w_mem_inst__abc_21203_new_n5767_), .Y(w_mem_inst__abc_21203_new_n5770_));
OR2X2 OR2X2_3446 ( .A(w_mem_inst__abc_21203_new_n5770_), .B(w_mem_inst__abc_21203_new_n5766_), .Y(w_mem_inst__0w_mem_3__31_0__19_));
OR2X2 OR2X2_3447 ( .A(w_mem_inst__abc_21203_new_n5775_), .B(w_mem_inst__abc_21203_new_n5773_), .Y(w_mem_inst__abc_21203_new_n5776_));
OR2X2 OR2X2_3448 ( .A(w_mem_inst__abc_21203_new_n5776_), .B(w_mem_inst__abc_21203_new_n5772_), .Y(w_mem_inst__0w_mem_3__31_0__20_));
OR2X2 OR2X2_3449 ( .A(w_mem_inst__abc_21203_new_n5781_), .B(w_mem_inst__abc_21203_new_n5779_), .Y(w_mem_inst__abc_21203_new_n5782_));
OR2X2 OR2X2_345 ( .A(_abc_15497_new_n1777_), .B(_abc_15497_new_n1774_), .Y(_abc_15497_new_n1778_));
OR2X2 OR2X2_3450 ( .A(w_mem_inst__abc_21203_new_n5782_), .B(w_mem_inst__abc_21203_new_n5778_), .Y(w_mem_inst__0w_mem_3__31_0__21_));
OR2X2 OR2X2_3451 ( .A(w_mem_inst__abc_21203_new_n5787_), .B(w_mem_inst__abc_21203_new_n5785_), .Y(w_mem_inst__abc_21203_new_n5788_));
OR2X2 OR2X2_3452 ( .A(w_mem_inst__abc_21203_new_n5788_), .B(w_mem_inst__abc_21203_new_n5784_), .Y(w_mem_inst__0w_mem_3__31_0__22_));
OR2X2 OR2X2_3453 ( .A(w_mem_inst__abc_21203_new_n5793_), .B(w_mem_inst__abc_21203_new_n5791_), .Y(w_mem_inst__abc_21203_new_n5794_));
OR2X2 OR2X2_3454 ( .A(w_mem_inst__abc_21203_new_n5794_), .B(w_mem_inst__abc_21203_new_n5790_), .Y(w_mem_inst__0w_mem_3__31_0__23_));
OR2X2 OR2X2_3455 ( .A(w_mem_inst__abc_21203_new_n5799_), .B(w_mem_inst__abc_21203_new_n5797_), .Y(w_mem_inst__abc_21203_new_n5800_));
OR2X2 OR2X2_3456 ( .A(w_mem_inst__abc_21203_new_n5800_), .B(w_mem_inst__abc_21203_new_n5796_), .Y(w_mem_inst__0w_mem_3__31_0__24_));
OR2X2 OR2X2_3457 ( .A(w_mem_inst__abc_21203_new_n5805_), .B(w_mem_inst__abc_21203_new_n5803_), .Y(w_mem_inst__abc_21203_new_n5806_));
OR2X2 OR2X2_3458 ( .A(w_mem_inst__abc_21203_new_n5806_), .B(w_mem_inst__abc_21203_new_n5802_), .Y(w_mem_inst__0w_mem_3__31_0__25_));
OR2X2 OR2X2_3459 ( .A(w_mem_inst__abc_21203_new_n5811_), .B(w_mem_inst__abc_21203_new_n5809_), .Y(w_mem_inst__abc_21203_new_n5812_));
OR2X2 OR2X2_346 ( .A(_abc_15497_new_n699_), .B(\digest[49] ), .Y(_abc_15497_new_n1780_));
OR2X2 OR2X2_3460 ( .A(w_mem_inst__abc_21203_new_n5812_), .B(w_mem_inst__abc_21203_new_n5808_), .Y(w_mem_inst__0w_mem_3__31_0__26_));
OR2X2 OR2X2_3461 ( .A(w_mem_inst__abc_21203_new_n5817_), .B(w_mem_inst__abc_21203_new_n5815_), .Y(w_mem_inst__abc_21203_new_n5818_));
OR2X2 OR2X2_3462 ( .A(w_mem_inst__abc_21203_new_n5818_), .B(w_mem_inst__abc_21203_new_n5814_), .Y(w_mem_inst__0w_mem_3__31_0__27_));
OR2X2 OR2X2_3463 ( .A(w_mem_inst__abc_21203_new_n5823_), .B(w_mem_inst__abc_21203_new_n5821_), .Y(w_mem_inst__abc_21203_new_n5824_));
OR2X2 OR2X2_3464 ( .A(w_mem_inst__abc_21203_new_n5824_), .B(w_mem_inst__abc_21203_new_n5820_), .Y(w_mem_inst__0w_mem_3__31_0__28_));
OR2X2 OR2X2_3465 ( .A(w_mem_inst__abc_21203_new_n5829_), .B(w_mem_inst__abc_21203_new_n5827_), .Y(w_mem_inst__abc_21203_new_n5830_));
OR2X2 OR2X2_3466 ( .A(w_mem_inst__abc_21203_new_n5830_), .B(w_mem_inst__abc_21203_new_n5826_), .Y(w_mem_inst__0w_mem_3__31_0__29_));
OR2X2 OR2X2_3467 ( .A(w_mem_inst__abc_21203_new_n5835_), .B(w_mem_inst__abc_21203_new_n5833_), .Y(w_mem_inst__abc_21203_new_n5836_));
OR2X2 OR2X2_3468 ( .A(w_mem_inst__abc_21203_new_n5836_), .B(w_mem_inst__abc_21203_new_n5832_), .Y(w_mem_inst__0w_mem_3__31_0__30_));
OR2X2 OR2X2_3469 ( .A(w_mem_inst__abc_21203_new_n5841_), .B(w_mem_inst__abc_21203_new_n5839_), .Y(w_mem_inst__abc_21203_new_n5842_));
OR2X2 OR2X2_347 ( .A(_abc_15497_new_n1779_), .B(_abc_15497_new_n1781_), .Y(_0H3_reg_31_0__17_));
OR2X2 OR2X2_3470 ( .A(w_mem_inst__abc_21203_new_n5842_), .B(w_mem_inst__abc_21203_new_n5838_), .Y(w_mem_inst__0w_mem_3__31_0__31_));
OR2X2 OR2X2_3471 ( .A(w_mem_inst__abc_21203_new_n5847_), .B(w_mem_inst__abc_21203_new_n5845_), .Y(w_mem_inst__abc_21203_new_n5848_));
OR2X2 OR2X2_3472 ( .A(w_mem_inst__abc_21203_new_n5848_), .B(w_mem_inst__abc_21203_new_n5844_), .Y(w_mem_inst__0w_mem_2__31_0__0_));
OR2X2 OR2X2_3473 ( .A(w_mem_inst__abc_21203_new_n5853_), .B(w_mem_inst__abc_21203_new_n5851_), .Y(w_mem_inst__abc_21203_new_n5854_));
OR2X2 OR2X2_3474 ( .A(w_mem_inst__abc_21203_new_n5854_), .B(w_mem_inst__abc_21203_new_n5850_), .Y(w_mem_inst__0w_mem_2__31_0__1_));
OR2X2 OR2X2_3475 ( .A(w_mem_inst__abc_21203_new_n5859_), .B(w_mem_inst__abc_21203_new_n5857_), .Y(w_mem_inst__abc_21203_new_n5860_));
OR2X2 OR2X2_3476 ( .A(w_mem_inst__abc_21203_new_n5860_), .B(w_mem_inst__abc_21203_new_n5856_), .Y(w_mem_inst__0w_mem_2__31_0__2_));
OR2X2 OR2X2_3477 ( .A(w_mem_inst__abc_21203_new_n5865_), .B(w_mem_inst__abc_21203_new_n5863_), .Y(w_mem_inst__abc_21203_new_n5866_));
OR2X2 OR2X2_3478 ( .A(w_mem_inst__abc_21203_new_n5866_), .B(w_mem_inst__abc_21203_new_n5862_), .Y(w_mem_inst__0w_mem_2__31_0__3_));
OR2X2 OR2X2_3479 ( .A(w_mem_inst__abc_21203_new_n5871_), .B(w_mem_inst__abc_21203_new_n5869_), .Y(w_mem_inst__abc_21203_new_n5872_));
OR2X2 OR2X2_348 ( .A(_abc_15497_new_n1784_), .B(_abc_15497_new_n1771_), .Y(_abc_15497_new_n1785_));
OR2X2 OR2X2_3480 ( .A(w_mem_inst__abc_21203_new_n5872_), .B(w_mem_inst__abc_21203_new_n5868_), .Y(w_mem_inst__0w_mem_2__31_0__4_));
OR2X2 OR2X2_3481 ( .A(w_mem_inst__abc_21203_new_n5877_), .B(w_mem_inst__abc_21203_new_n5875_), .Y(w_mem_inst__abc_21203_new_n5878_));
OR2X2 OR2X2_3482 ( .A(w_mem_inst__abc_21203_new_n5878_), .B(w_mem_inst__abc_21203_new_n5874_), .Y(w_mem_inst__0w_mem_2__31_0__5_));
OR2X2 OR2X2_3483 ( .A(w_mem_inst__abc_21203_new_n5883_), .B(w_mem_inst__abc_21203_new_n5881_), .Y(w_mem_inst__abc_21203_new_n5884_));
OR2X2 OR2X2_3484 ( .A(w_mem_inst__abc_21203_new_n5884_), .B(w_mem_inst__abc_21203_new_n5880_), .Y(w_mem_inst__0w_mem_2__31_0__6_));
OR2X2 OR2X2_3485 ( .A(w_mem_inst__abc_21203_new_n5889_), .B(w_mem_inst__abc_21203_new_n5887_), .Y(w_mem_inst__abc_21203_new_n5890_));
OR2X2 OR2X2_3486 ( .A(w_mem_inst__abc_21203_new_n5890_), .B(w_mem_inst__abc_21203_new_n5886_), .Y(w_mem_inst__0w_mem_2__31_0__7_));
OR2X2 OR2X2_3487 ( .A(w_mem_inst__abc_21203_new_n5895_), .B(w_mem_inst__abc_21203_new_n5893_), .Y(w_mem_inst__abc_21203_new_n5896_));
OR2X2 OR2X2_3488 ( .A(w_mem_inst__abc_21203_new_n5896_), .B(w_mem_inst__abc_21203_new_n5892_), .Y(w_mem_inst__0w_mem_2__31_0__8_));
OR2X2 OR2X2_3489 ( .A(w_mem_inst__abc_21203_new_n5901_), .B(w_mem_inst__abc_21203_new_n5899_), .Y(w_mem_inst__abc_21203_new_n5902_));
OR2X2 OR2X2_349 ( .A(_abc_15497_new_n1787_), .B(_abc_15497_new_n1785_), .Y(_abc_15497_new_n1788_));
OR2X2 OR2X2_3490 ( .A(w_mem_inst__abc_21203_new_n5902_), .B(w_mem_inst__abc_21203_new_n5898_), .Y(w_mem_inst__0w_mem_2__31_0__9_));
OR2X2 OR2X2_3491 ( .A(w_mem_inst__abc_21203_new_n5907_), .B(w_mem_inst__abc_21203_new_n5905_), .Y(w_mem_inst__abc_21203_new_n5908_));
OR2X2 OR2X2_3492 ( .A(w_mem_inst__abc_21203_new_n5908_), .B(w_mem_inst__abc_21203_new_n5904_), .Y(w_mem_inst__0w_mem_2__31_0__10_));
OR2X2 OR2X2_3493 ( .A(w_mem_inst__abc_21203_new_n5913_), .B(w_mem_inst__abc_21203_new_n5911_), .Y(w_mem_inst__abc_21203_new_n5914_));
OR2X2 OR2X2_3494 ( .A(w_mem_inst__abc_21203_new_n5914_), .B(w_mem_inst__abc_21203_new_n5910_), .Y(w_mem_inst__0w_mem_2__31_0__11_));
OR2X2 OR2X2_3495 ( .A(w_mem_inst__abc_21203_new_n5919_), .B(w_mem_inst__abc_21203_new_n5917_), .Y(w_mem_inst__abc_21203_new_n5920_));
OR2X2 OR2X2_3496 ( .A(w_mem_inst__abc_21203_new_n5920_), .B(w_mem_inst__abc_21203_new_n5916_), .Y(w_mem_inst__0w_mem_2__31_0__12_));
OR2X2 OR2X2_3497 ( .A(w_mem_inst__abc_21203_new_n5925_), .B(w_mem_inst__abc_21203_new_n5923_), .Y(w_mem_inst__abc_21203_new_n5926_));
OR2X2 OR2X2_3498 ( .A(w_mem_inst__abc_21203_new_n5926_), .B(w_mem_inst__abc_21203_new_n5922_), .Y(w_mem_inst__0w_mem_2__31_0__13_));
OR2X2 OR2X2_3499 ( .A(w_mem_inst__abc_21203_new_n5931_), .B(w_mem_inst__abc_21203_new_n5929_), .Y(w_mem_inst__abc_21203_new_n5932_));
OR2X2 OR2X2_35 ( .A(_abc_15497_new_n830_), .B(_abc_15497_new_n815_), .Y(_abc_15497_new_n831_));
OR2X2 OR2X2_350 ( .A(\digest[50] ), .B(d_reg_18_), .Y(_abc_15497_new_n1789_));
OR2X2 OR2X2_3500 ( .A(w_mem_inst__abc_21203_new_n5932_), .B(w_mem_inst__abc_21203_new_n5928_), .Y(w_mem_inst__0w_mem_2__31_0__14_));
OR2X2 OR2X2_3501 ( .A(w_mem_inst__abc_21203_new_n5937_), .B(w_mem_inst__abc_21203_new_n5935_), .Y(w_mem_inst__abc_21203_new_n5938_));
OR2X2 OR2X2_3502 ( .A(w_mem_inst__abc_21203_new_n5938_), .B(w_mem_inst__abc_21203_new_n5934_), .Y(w_mem_inst__0w_mem_2__31_0__15_));
OR2X2 OR2X2_3503 ( .A(w_mem_inst__abc_21203_new_n5943_), .B(w_mem_inst__abc_21203_new_n5941_), .Y(w_mem_inst__abc_21203_new_n5944_));
OR2X2 OR2X2_3504 ( .A(w_mem_inst__abc_21203_new_n5944_), .B(w_mem_inst__abc_21203_new_n5940_), .Y(w_mem_inst__0w_mem_2__31_0__16_));
OR2X2 OR2X2_3505 ( .A(w_mem_inst__abc_21203_new_n5949_), .B(w_mem_inst__abc_21203_new_n5947_), .Y(w_mem_inst__abc_21203_new_n5950_));
OR2X2 OR2X2_3506 ( .A(w_mem_inst__abc_21203_new_n5950_), .B(w_mem_inst__abc_21203_new_n5946_), .Y(w_mem_inst__0w_mem_2__31_0__17_));
OR2X2 OR2X2_3507 ( .A(w_mem_inst__abc_21203_new_n5955_), .B(w_mem_inst__abc_21203_new_n5953_), .Y(w_mem_inst__abc_21203_new_n5956_));
OR2X2 OR2X2_3508 ( .A(w_mem_inst__abc_21203_new_n5956_), .B(w_mem_inst__abc_21203_new_n5952_), .Y(w_mem_inst__0w_mem_2__31_0__18_));
OR2X2 OR2X2_3509 ( .A(w_mem_inst__abc_21203_new_n5961_), .B(w_mem_inst__abc_21203_new_n5959_), .Y(w_mem_inst__abc_21203_new_n5962_));
OR2X2 OR2X2_351 ( .A(_abc_15497_new_n1788_), .B(_abc_15497_new_n1792_), .Y(_abc_15497_new_n1793_));
OR2X2 OR2X2_3510 ( .A(w_mem_inst__abc_21203_new_n5962_), .B(w_mem_inst__abc_21203_new_n5958_), .Y(w_mem_inst__0w_mem_2__31_0__19_));
OR2X2 OR2X2_3511 ( .A(w_mem_inst__abc_21203_new_n5967_), .B(w_mem_inst__abc_21203_new_n5965_), .Y(w_mem_inst__abc_21203_new_n5968_));
OR2X2 OR2X2_3512 ( .A(w_mem_inst__abc_21203_new_n5968_), .B(w_mem_inst__abc_21203_new_n5964_), .Y(w_mem_inst__0w_mem_2__31_0__20_));
OR2X2 OR2X2_3513 ( .A(w_mem_inst__abc_21203_new_n5973_), .B(w_mem_inst__abc_21203_new_n5971_), .Y(w_mem_inst__abc_21203_new_n5974_));
OR2X2 OR2X2_3514 ( .A(w_mem_inst__abc_21203_new_n5974_), .B(w_mem_inst__abc_21203_new_n5970_), .Y(w_mem_inst__0w_mem_2__31_0__21_));
OR2X2 OR2X2_3515 ( .A(w_mem_inst__abc_21203_new_n5979_), .B(w_mem_inst__abc_21203_new_n5977_), .Y(w_mem_inst__abc_21203_new_n5980_));
OR2X2 OR2X2_3516 ( .A(w_mem_inst__abc_21203_new_n5980_), .B(w_mem_inst__abc_21203_new_n5976_), .Y(w_mem_inst__0w_mem_2__31_0__22_));
OR2X2 OR2X2_3517 ( .A(w_mem_inst__abc_21203_new_n5985_), .B(w_mem_inst__abc_21203_new_n5983_), .Y(w_mem_inst__abc_21203_new_n5986_));
OR2X2 OR2X2_3518 ( .A(w_mem_inst__abc_21203_new_n5986_), .B(w_mem_inst__abc_21203_new_n5982_), .Y(w_mem_inst__0w_mem_2__31_0__23_));
OR2X2 OR2X2_3519 ( .A(w_mem_inst__abc_21203_new_n5991_), .B(w_mem_inst__abc_21203_new_n5989_), .Y(w_mem_inst__abc_21203_new_n5992_));
OR2X2 OR2X2_352 ( .A(_abc_15497_new_n1797_), .B(_abc_15497_new_n1783_), .Y(_0H3_reg_31_0__18_));
OR2X2 OR2X2_3520 ( .A(w_mem_inst__abc_21203_new_n5992_), .B(w_mem_inst__abc_21203_new_n5988_), .Y(w_mem_inst__0w_mem_2__31_0__24_));
OR2X2 OR2X2_3521 ( .A(w_mem_inst__abc_21203_new_n5997_), .B(w_mem_inst__abc_21203_new_n5995_), .Y(w_mem_inst__abc_21203_new_n5998_));
OR2X2 OR2X2_3522 ( .A(w_mem_inst__abc_21203_new_n5998_), .B(w_mem_inst__abc_21203_new_n5994_), .Y(w_mem_inst__0w_mem_2__31_0__25_));
OR2X2 OR2X2_3523 ( .A(w_mem_inst__abc_21203_new_n6003_), .B(w_mem_inst__abc_21203_new_n6001_), .Y(w_mem_inst__abc_21203_new_n6004_));
OR2X2 OR2X2_3524 ( .A(w_mem_inst__abc_21203_new_n6004_), .B(w_mem_inst__abc_21203_new_n6000_), .Y(w_mem_inst__0w_mem_2__31_0__26_));
OR2X2 OR2X2_3525 ( .A(w_mem_inst__abc_21203_new_n6009_), .B(w_mem_inst__abc_21203_new_n6007_), .Y(w_mem_inst__abc_21203_new_n6010_));
OR2X2 OR2X2_3526 ( .A(w_mem_inst__abc_21203_new_n6010_), .B(w_mem_inst__abc_21203_new_n6006_), .Y(w_mem_inst__0w_mem_2__31_0__27_));
OR2X2 OR2X2_3527 ( .A(w_mem_inst__abc_21203_new_n6015_), .B(w_mem_inst__abc_21203_new_n6013_), .Y(w_mem_inst__abc_21203_new_n6016_));
OR2X2 OR2X2_3528 ( .A(w_mem_inst__abc_21203_new_n6016_), .B(w_mem_inst__abc_21203_new_n6012_), .Y(w_mem_inst__0w_mem_2__31_0__28_));
OR2X2 OR2X2_3529 ( .A(w_mem_inst__abc_21203_new_n6021_), .B(w_mem_inst__abc_21203_new_n6019_), .Y(w_mem_inst__abc_21203_new_n6022_));
OR2X2 OR2X2_353 ( .A(\digest[51] ), .B(d_reg_19_), .Y(_abc_15497_new_n1802_));
OR2X2 OR2X2_3530 ( .A(w_mem_inst__abc_21203_new_n6022_), .B(w_mem_inst__abc_21203_new_n6018_), .Y(w_mem_inst__0w_mem_2__31_0__29_));
OR2X2 OR2X2_3531 ( .A(w_mem_inst__abc_21203_new_n6027_), .B(w_mem_inst__abc_21203_new_n6025_), .Y(w_mem_inst__abc_21203_new_n6028_));
OR2X2 OR2X2_3532 ( .A(w_mem_inst__abc_21203_new_n6028_), .B(w_mem_inst__abc_21203_new_n6024_), .Y(w_mem_inst__0w_mem_2__31_0__30_));
OR2X2 OR2X2_3533 ( .A(w_mem_inst__abc_21203_new_n6033_), .B(w_mem_inst__abc_21203_new_n6031_), .Y(w_mem_inst__abc_21203_new_n6034_));
OR2X2 OR2X2_3534 ( .A(w_mem_inst__abc_21203_new_n6034_), .B(w_mem_inst__abc_21203_new_n6030_), .Y(w_mem_inst__0w_mem_2__31_0__31_));
OR2X2 OR2X2_3535 ( .A(w_mem_inst__abc_21203_new_n6039_), .B(w_mem_inst__abc_21203_new_n6037_), .Y(w_mem_inst__abc_21203_new_n6040_));
OR2X2 OR2X2_3536 ( .A(w_mem_inst__abc_21203_new_n6040_), .B(w_mem_inst__abc_21203_new_n6036_), .Y(w_mem_inst__0w_mem_0__31_0__0_));
OR2X2 OR2X2_3537 ( .A(w_mem_inst__abc_21203_new_n6045_), .B(w_mem_inst__abc_21203_new_n6043_), .Y(w_mem_inst__abc_21203_new_n6046_));
OR2X2 OR2X2_3538 ( .A(w_mem_inst__abc_21203_new_n6046_), .B(w_mem_inst__abc_21203_new_n6042_), .Y(w_mem_inst__0w_mem_0__31_0__1_));
OR2X2 OR2X2_3539 ( .A(w_mem_inst__abc_21203_new_n6051_), .B(w_mem_inst__abc_21203_new_n6049_), .Y(w_mem_inst__abc_21203_new_n6052_));
OR2X2 OR2X2_354 ( .A(_abc_15497_new_n1801_), .B(_abc_15497_new_n1805_), .Y(_abc_15497_new_n1806_));
OR2X2 OR2X2_3540 ( .A(w_mem_inst__abc_21203_new_n6052_), .B(w_mem_inst__abc_21203_new_n6048_), .Y(w_mem_inst__0w_mem_0__31_0__2_));
OR2X2 OR2X2_3541 ( .A(w_mem_inst__abc_21203_new_n6057_), .B(w_mem_inst__abc_21203_new_n6055_), .Y(w_mem_inst__abc_21203_new_n6058_));
OR2X2 OR2X2_3542 ( .A(w_mem_inst__abc_21203_new_n6058_), .B(w_mem_inst__abc_21203_new_n6054_), .Y(w_mem_inst__0w_mem_0__31_0__3_));
OR2X2 OR2X2_3543 ( .A(w_mem_inst__abc_21203_new_n6063_), .B(w_mem_inst__abc_21203_new_n6061_), .Y(w_mem_inst__abc_21203_new_n6064_));
OR2X2 OR2X2_3544 ( .A(w_mem_inst__abc_21203_new_n6064_), .B(w_mem_inst__abc_21203_new_n6060_), .Y(w_mem_inst__0w_mem_0__31_0__4_));
OR2X2 OR2X2_3545 ( .A(w_mem_inst__abc_21203_new_n6069_), .B(w_mem_inst__abc_21203_new_n6067_), .Y(w_mem_inst__abc_21203_new_n6070_));
OR2X2 OR2X2_3546 ( .A(w_mem_inst__abc_21203_new_n6070_), .B(w_mem_inst__abc_21203_new_n6066_), .Y(w_mem_inst__0w_mem_0__31_0__5_));
OR2X2 OR2X2_3547 ( .A(w_mem_inst__abc_21203_new_n6075_), .B(w_mem_inst__abc_21203_new_n6073_), .Y(w_mem_inst__abc_21203_new_n6076_));
OR2X2 OR2X2_3548 ( .A(w_mem_inst__abc_21203_new_n6076_), .B(w_mem_inst__abc_21203_new_n6072_), .Y(w_mem_inst__0w_mem_0__31_0__6_));
OR2X2 OR2X2_3549 ( .A(w_mem_inst__abc_21203_new_n6081_), .B(w_mem_inst__abc_21203_new_n6079_), .Y(w_mem_inst__abc_21203_new_n6082_));
OR2X2 OR2X2_355 ( .A(_abc_15497_new_n1800_), .B(_abc_15497_new_n1807_), .Y(_abc_15497_new_n1808_));
OR2X2 OR2X2_3550 ( .A(w_mem_inst__abc_21203_new_n6082_), .B(w_mem_inst__abc_21203_new_n6078_), .Y(w_mem_inst__0w_mem_0__31_0__7_));
OR2X2 OR2X2_3551 ( .A(w_mem_inst__abc_21203_new_n6087_), .B(w_mem_inst__abc_21203_new_n6085_), .Y(w_mem_inst__abc_21203_new_n6088_));
OR2X2 OR2X2_3552 ( .A(w_mem_inst__abc_21203_new_n6088_), .B(w_mem_inst__abc_21203_new_n6084_), .Y(w_mem_inst__0w_mem_0__31_0__8_));
OR2X2 OR2X2_3553 ( .A(w_mem_inst__abc_21203_new_n6093_), .B(w_mem_inst__abc_21203_new_n6091_), .Y(w_mem_inst__abc_21203_new_n6094_));
OR2X2 OR2X2_3554 ( .A(w_mem_inst__abc_21203_new_n6094_), .B(w_mem_inst__abc_21203_new_n6090_), .Y(w_mem_inst__0w_mem_0__31_0__9_));
OR2X2 OR2X2_3555 ( .A(w_mem_inst__abc_21203_new_n6099_), .B(w_mem_inst__abc_21203_new_n6097_), .Y(w_mem_inst__abc_21203_new_n6100_));
OR2X2 OR2X2_3556 ( .A(w_mem_inst__abc_21203_new_n6100_), .B(w_mem_inst__abc_21203_new_n6096_), .Y(w_mem_inst__0w_mem_0__31_0__10_));
OR2X2 OR2X2_3557 ( .A(w_mem_inst__abc_21203_new_n6105_), .B(w_mem_inst__abc_21203_new_n6103_), .Y(w_mem_inst__abc_21203_new_n6106_));
OR2X2 OR2X2_3558 ( .A(w_mem_inst__abc_21203_new_n6106_), .B(w_mem_inst__abc_21203_new_n6102_), .Y(w_mem_inst__0w_mem_0__31_0__11_));
OR2X2 OR2X2_3559 ( .A(w_mem_inst__abc_21203_new_n6111_), .B(w_mem_inst__abc_21203_new_n6109_), .Y(w_mem_inst__abc_21203_new_n6112_));
OR2X2 OR2X2_356 ( .A(_abc_15497_new_n1810_), .B(_abc_15497_new_n1799_), .Y(_0H3_reg_31_0__19_));
OR2X2 OR2X2_3560 ( .A(w_mem_inst__abc_21203_new_n6112_), .B(w_mem_inst__abc_21203_new_n6108_), .Y(w_mem_inst__0w_mem_0__31_0__12_));
OR2X2 OR2X2_3561 ( .A(w_mem_inst__abc_21203_new_n6117_), .B(w_mem_inst__abc_21203_new_n6115_), .Y(w_mem_inst__abc_21203_new_n6118_));
OR2X2 OR2X2_3562 ( .A(w_mem_inst__abc_21203_new_n6118_), .B(w_mem_inst__abc_21203_new_n6114_), .Y(w_mem_inst__0w_mem_0__31_0__13_));
OR2X2 OR2X2_3563 ( .A(w_mem_inst__abc_21203_new_n6123_), .B(w_mem_inst__abc_21203_new_n6121_), .Y(w_mem_inst__abc_21203_new_n6124_));
OR2X2 OR2X2_3564 ( .A(w_mem_inst__abc_21203_new_n6124_), .B(w_mem_inst__abc_21203_new_n6120_), .Y(w_mem_inst__0w_mem_0__31_0__14_));
OR2X2 OR2X2_3565 ( .A(w_mem_inst__abc_21203_new_n6129_), .B(w_mem_inst__abc_21203_new_n6127_), .Y(w_mem_inst__abc_21203_new_n6130_));
OR2X2 OR2X2_3566 ( .A(w_mem_inst__abc_21203_new_n6130_), .B(w_mem_inst__abc_21203_new_n6126_), .Y(w_mem_inst__0w_mem_0__31_0__15_));
OR2X2 OR2X2_3567 ( .A(w_mem_inst__abc_21203_new_n6135_), .B(w_mem_inst__abc_21203_new_n6133_), .Y(w_mem_inst__abc_21203_new_n6136_));
OR2X2 OR2X2_3568 ( .A(w_mem_inst__abc_21203_new_n6136_), .B(w_mem_inst__abc_21203_new_n6132_), .Y(w_mem_inst__0w_mem_0__31_0__16_));
OR2X2 OR2X2_3569 ( .A(w_mem_inst__abc_21203_new_n6141_), .B(w_mem_inst__abc_21203_new_n6139_), .Y(w_mem_inst__abc_21203_new_n6142_));
OR2X2 OR2X2_357 ( .A(_abc_15497_new_n1816_), .B(_abc_15497_new_n1803_), .Y(_abc_15497_new_n1817_));
OR2X2 OR2X2_3570 ( .A(w_mem_inst__abc_21203_new_n6142_), .B(w_mem_inst__abc_21203_new_n6138_), .Y(w_mem_inst__0w_mem_0__31_0__17_));
OR2X2 OR2X2_3571 ( .A(w_mem_inst__abc_21203_new_n6147_), .B(w_mem_inst__abc_21203_new_n6145_), .Y(w_mem_inst__abc_21203_new_n6148_));
OR2X2 OR2X2_3572 ( .A(w_mem_inst__abc_21203_new_n6148_), .B(w_mem_inst__abc_21203_new_n6144_), .Y(w_mem_inst__0w_mem_0__31_0__18_));
OR2X2 OR2X2_3573 ( .A(w_mem_inst__abc_21203_new_n6153_), .B(w_mem_inst__abc_21203_new_n6151_), .Y(w_mem_inst__abc_21203_new_n6154_));
OR2X2 OR2X2_3574 ( .A(w_mem_inst__abc_21203_new_n6154_), .B(w_mem_inst__abc_21203_new_n6150_), .Y(w_mem_inst__0w_mem_0__31_0__19_));
OR2X2 OR2X2_3575 ( .A(w_mem_inst__abc_21203_new_n6159_), .B(w_mem_inst__abc_21203_new_n6157_), .Y(w_mem_inst__abc_21203_new_n6160_));
OR2X2 OR2X2_3576 ( .A(w_mem_inst__abc_21203_new_n6160_), .B(w_mem_inst__abc_21203_new_n6156_), .Y(w_mem_inst__0w_mem_0__31_0__20_));
OR2X2 OR2X2_3577 ( .A(w_mem_inst__abc_21203_new_n6165_), .B(w_mem_inst__abc_21203_new_n6163_), .Y(w_mem_inst__abc_21203_new_n6166_));
OR2X2 OR2X2_3578 ( .A(w_mem_inst__abc_21203_new_n6166_), .B(w_mem_inst__abc_21203_new_n6162_), .Y(w_mem_inst__0w_mem_0__31_0__21_));
OR2X2 OR2X2_3579 ( .A(w_mem_inst__abc_21203_new_n6171_), .B(w_mem_inst__abc_21203_new_n6169_), .Y(w_mem_inst__abc_21203_new_n6172_));
OR2X2 OR2X2_358 ( .A(_abc_15497_new_n1815_), .B(_abc_15497_new_n1817_), .Y(_abc_15497_new_n1818_));
OR2X2 OR2X2_3580 ( .A(w_mem_inst__abc_21203_new_n6172_), .B(w_mem_inst__abc_21203_new_n6168_), .Y(w_mem_inst__0w_mem_0__31_0__22_));
OR2X2 OR2X2_3581 ( .A(w_mem_inst__abc_21203_new_n6177_), .B(w_mem_inst__abc_21203_new_n6175_), .Y(w_mem_inst__abc_21203_new_n6178_));
OR2X2 OR2X2_3582 ( .A(w_mem_inst__abc_21203_new_n6178_), .B(w_mem_inst__abc_21203_new_n6174_), .Y(w_mem_inst__0w_mem_0__31_0__23_));
OR2X2 OR2X2_3583 ( .A(w_mem_inst__abc_21203_new_n6183_), .B(w_mem_inst__abc_21203_new_n6181_), .Y(w_mem_inst__abc_21203_new_n6184_));
OR2X2 OR2X2_3584 ( .A(w_mem_inst__abc_21203_new_n6184_), .B(w_mem_inst__abc_21203_new_n6180_), .Y(w_mem_inst__0w_mem_0__31_0__24_));
OR2X2 OR2X2_3585 ( .A(w_mem_inst__abc_21203_new_n6189_), .B(w_mem_inst__abc_21203_new_n6187_), .Y(w_mem_inst__abc_21203_new_n6190_));
OR2X2 OR2X2_3586 ( .A(w_mem_inst__abc_21203_new_n6190_), .B(w_mem_inst__abc_21203_new_n6186_), .Y(w_mem_inst__0w_mem_0__31_0__25_));
OR2X2 OR2X2_3587 ( .A(w_mem_inst__abc_21203_new_n6195_), .B(w_mem_inst__abc_21203_new_n6193_), .Y(w_mem_inst__abc_21203_new_n6196_));
OR2X2 OR2X2_3588 ( .A(w_mem_inst__abc_21203_new_n6196_), .B(w_mem_inst__abc_21203_new_n6192_), .Y(w_mem_inst__0w_mem_0__31_0__26_));
OR2X2 OR2X2_3589 ( .A(w_mem_inst__abc_21203_new_n6201_), .B(w_mem_inst__abc_21203_new_n6199_), .Y(w_mem_inst__abc_21203_new_n6202_));
OR2X2 OR2X2_359 ( .A(_abc_15497_new_n1814_), .B(_abc_15497_new_n1818_), .Y(_abc_15497_new_n1819_));
OR2X2 OR2X2_3590 ( .A(w_mem_inst__abc_21203_new_n6202_), .B(w_mem_inst__abc_21203_new_n6198_), .Y(w_mem_inst__0w_mem_0__31_0__27_));
OR2X2 OR2X2_3591 ( .A(w_mem_inst__abc_21203_new_n6207_), .B(w_mem_inst__abc_21203_new_n6205_), .Y(w_mem_inst__abc_21203_new_n6208_));
OR2X2 OR2X2_3592 ( .A(w_mem_inst__abc_21203_new_n6208_), .B(w_mem_inst__abc_21203_new_n6204_), .Y(w_mem_inst__0w_mem_0__31_0__28_));
OR2X2 OR2X2_3593 ( .A(w_mem_inst__abc_21203_new_n6213_), .B(w_mem_inst__abc_21203_new_n6211_), .Y(w_mem_inst__abc_21203_new_n6214_));
OR2X2 OR2X2_3594 ( .A(w_mem_inst__abc_21203_new_n6214_), .B(w_mem_inst__abc_21203_new_n6210_), .Y(w_mem_inst__0w_mem_0__31_0__29_));
OR2X2 OR2X2_3595 ( .A(w_mem_inst__abc_21203_new_n6219_), .B(w_mem_inst__abc_21203_new_n6217_), .Y(w_mem_inst__abc_21203_new_n6220_));
OR2X2 OR2X2_3596 ( .A(w_mem_inst__abc_21203_new_n6220_), .B(w_mem_inst__abc_21203_new_n6216_), .Y(w_mem_inst__0w_mem_0__31_0__30_));
OR2X2 OR2X2_3597 ( .A(w_mem_inst__abc_21203_new_n6225_), .B(w_mem_inst__abc_21203_new_n6223_), .Y(w_mem_inst__abc_21203_new_n6226_));
OR2X2 OR2X2_3598 ( .A(w_mem_inst__abc_21203_new_n6226_), .B(w_mem_inst__abc_21203_new_n6222_), .Y(w_mem_inst__0w_mem_0__31_0__31_));
OR2X2 OR2X2_3599 ( .A(w_mem_inst_w_ctr_reg_0_), .B(round_ctr_inc), .Y(w_mem_inst__abc_21203_new_n6228_));
OR2X2 OR2X2_36 ( .A(c_reg_4_), .B(\digest[68] ), .Y(_abc_15497_new_n833_));
OR2X2 OR2X2_360 ( .A(\digest[52] ), .B(d_reg_20_), .Y(_abc_15497_new_n1820_));
OR2X2 OR2X2_3600 ( .A(w_mem_inst__abc_21203_new_n6230_), .B(w_mem_inst__abc_21203_new_n1610_), .Y(w_mem_inst__abc_21203_new_n6231_));
OR2X2 OR2X2_3601 ( .A(w_mem_inst__abc_21203_new_n1604_), .B(w_mem_inst__abc_21203_new_n1639_), .Y(w_mem_inst__abc_21203_new_n6234_));
OR2X2 OR2X2_3602 ( .A(w_mem_inst__abc_21203_new_n6235_), .B(w_mem_inst__abc_21203_new_n6233_), .Y(w_mem_inst__0w_ctr_reg_6_0__1_));
OR2X2 OR2X2_3603 ( .A(w_mem_inst__abc_21203_new_n3152_), .B(round_ctr_inc), .Y(w_mem_inst__abc_21203_new_n6237_));
OR2X2 OR2X2_3604 ( .A(w_mem_inst__abc_21203_new_n6238_), .B(w_mem_inst__abc_21203_new_n6239_), .Y(w_mem_inst__abc_21203_new_n6240_));
OR2X2 OR2X2_3605 ( .A(w_mem_inst__abc_21203_new_n6242_), .B(w_mem_inst__abc_21203_new_n6245_), .Y(w_mem_inst__abc_21203_new_n6246_));
OR2X2 OR2X2_3606 ( .A(w_mem_inst__abc_21203_new_n6247_), .B(w_mem_inst__abc_21203_new_n6250_), .Y(w_mem_inst__abc_21203_new_n6251_));
OR2X2 OR2X2_3607 ( .A(w_mem_inst__abc_21203_new_n6252_), .B(w_mem_inst__abc_21203_new_n6255_), .Y(w_mem_inst__abc_21203_new_n6256_));
OR2X2 OR2X2_3608 ( .A(w_mem_inst__abc_21203_new_n6257_), .B(w_mem_inst__abc_21203_new_n6260_), .Y(w_mem_inst__abc_21203_new_n6261_));
OR2X2 OR2X2_361 ( .A(_abc_15497_new_n1819_), .B(_abc_15497_new_n1823_), .Y(_abc_15497_new_n1824_));
OR2X2 OR2X2_362 ( .A(_abc_15497_new_n699_), .B(\digest[52] ), .Y(_abc_15497_new_n1829_));
OR2X2 OR2X2_363 ( .A(_abc_15497_new_n1828_), .B(_abc_15497_new_n1830_), .Y(_0H3_reg_31_0__20_));
OR2X2 OR2X2_364 ( .A(\digest[53] ), .B(d_reg_21_), .Y(_abc_15497_new_n1834_));
OR2X2 OR2X2_365 ( .A(_abc_15497_new_n1833_), .B(_abc_15497_new_n1837_), .Y(_abc_15497_new_n1838_));
OR2X2 OR2X2_366 ( .A(_abc_15497_new_n1832_), .B(_abc_15497_new_n1839_), .Y(_abc_15497_new_n1840_));
OR2X2 OR2X2_367 ( .A(_abc_15497_new_n699_), .B(\digest[53] ), .Y(_abc_15497_new_n1843_));
OR2X2 OR2X2_368 ( .A(_abc_15497_new_n1842_), .B(_abc_15497_new_n1844_), .Y(_0H3_reg_31_0__21_));
OR2X2 OR2X2_369 ( .A(\digest[54] ), .B(d_reg_22_), .Y(_abc_15497_new_n1847_));
OR2X2 OR2X2_37 ( .A(_abc_15497_new_n835_), .B(_abc_15497_new_n814_), .Y(_abc_15497_new_n836_));
OR2X2 OR2X2_370 ( .A(_abc_15497_new_n1853_), .B(_abc_15497_new_n1851_), .Y(_abc_15497_new_n1854_));
OR2X2 OR2X2_371 ( .A(_abc_15497_new_n1855_), .B(_abc_15497_new_n1850_), .Y(_abc_15497_new_n1856_));
OR2X2 OR2X2_372 ( .A(_abc_15497_new_n1860_), .B(_abc_15497_new_n1846_), .Y(_0H3_reg_31_0__22_));
OR2X2 OR2X2_373 ( .A(_abc_15497_new_n1857_), .B(_abc_15497_new_n1848_), .Y(_abc_15497_new_n1863_));
OR2X2 OR2X2_374 ( .A(\digest[55] ), .B(d_reg_23_), .Y(_abc_15497_new_n1864_));
OR2X2 OR2X2_375 ( .A(_abc_15497_new_n1863_), .B(_abc_15497_new_n1867_), .Y(_abc_15497_new_n1868_));
OR2X2 OR2X2_376 ( .A(_abc_15497_new_n1869_), .B(_abc_15497_new_n1870_), .Y(_abc_15497_new_n1871_));
OR2X2 OR2X2_377 ( .A(_abc_15497_new_n1873_), .B(_abc_15497_new_n1862_), .Y(_0H3_reg_31_0__23_));
OR2X2 OR2X2_378 ( .A(_abc_15497_new_n1876_), .B(_abc_15497_new_n1865_), .Y(_abc_15497_new_n1877_));
OR2X2 OR2X2_379 ( .A(_abc_15497_new_n1852_), .B(_abc_15497_new_n1851_), .Y(_abc_15497_new_n1879_));
OR2X2 OR2X2_38 ( .A(_abc_15497_new_n837_), .B(_abc_15497_new_n812_), .Y(_abc_15497_new_n838_));
OR2X2 OR2X2_380 ( .A(_abc_15497_new_n1881_), .B(_abc_15497_new_n1879_), .Y(_abc_15497_new_n1882_));
OR2X2 OR2X2_381 ( .A(_abc_15497_new_n1887_), .B(_abc_15497_new_n1884_), .Y(_abc_15497_new_n1888_));
OR2X2 OR2X2_382 ( .A(\digest[56] ), .B(d_reg_24_), .Y(_abc_15497_new_n1889_));
OR2X2 OR2X2_383 ( .A(_abc_15497_new_n1888_), .B(_abc_15497_new_n1892_), .Y(_abc_15497_new_n1893_));
OR2X2 OR2X2_384 ( .A(_abc_15497_new_n1897_), .B(_abc_15497_new_n1875_), .Y(_0H3_reg_31_0__24_));
OR2X2 OR2X2_385 ( .A(\digest[57] ), .B(d_reg_25_), .Y(_abc_15497_new_n1900_));
OR2X2 OR2X2_386 ( .A(_abc_15497_new_n1903_), .B(_abc_15497_new_n1890_), .Y(_abc_15497_new_n1904_));
OR2X2 OR2X2_387 ( .A(_abc_15497_new_n1894_), .B(_abc_15497_new_n1904_), .Y(_abc_15497_new_n1905_));
OR2X2 OR2X2_388 ( .A(_abc_15497_new_n1913_), .B(_abc_15497_new_n1899_), .Y(_0H3_reg_31_0__25_));
OR2X2 OR2X2_389 ( .A(\digest[58] ), .B(d_reg_26_), .Y(_abc_15497_new_n1919_));
OR2X2 OR2X2_39 ( .A(_abc_15497_new_n839_), .B(_abc_15497_new_n805_), .Y(_abc_15497_new_n840_));
OR2X2 OR2X2_390 ( .A(_abc_15497_new_n1918_), .B(_abc_15497_new_n1922_), .Y(_abc_15497_new_n1923_));
OR2X2 OR2X2_391 ( .A(_abc_15497_new_n1927_), .B(_abc_15497_new_n1915_), .Y(_0H3_reg_31_0__26_));
OR2X2 OR2X2_392 ( .A(\digest[59] ), .B(d_reg_27_), .Y(_abc_15497_new_n1930_));
OR2X2 OR2X2_393 ( .A(_abc_15497_new_n1933_), .B(_abc_15497_new_n1920_), .Y(_abc_15497_new_n1934_));
OR2X2 OR2X2_394 ( .A(_abc_15497_new_n1924_), .B(_abc_15497_new_n1934_), .Y(_abc_15497_new_n1935_));
OR2X2 OR2X2_395 ( .A(_abc_15497_new_n1917_), .B(_abc_15497_new_n1937_), .Y(_abc_15497_new_n1938_));
OR2X2 OR2X2_396 ( .A(_abc_15497_new_n1943_), .B(_abc_15497_new_n1929_), .Y(_0H3_reg_31_0__27_));
OR2X2 OR2X2_397 ( .A(_abc_15497_new_n1916_), .B(_abc_15497_new_n1937_), .Y(_abc_15497_new_n1948_));
OR2X2 OR2X2_398 ( .A(_abc_15497_new_n1946_), .B(_abc_15497_new_n1950_), .Y(_abc_15497_new_n1951_));
OR2X2 OR2X2_399 ( .A(\digest[60] ), .B(d_reg_28_), .Y(_abc_15497_new_n1952_));
OR2X2 OR2X2_4 ( .A(_abc_15497_new_n719_), .B(_abc_15497_new_n716_), .Y(_abc_15497_new_n720_));
OR2X2 OR2X2_40 ( .A(c_reg_8_), .B(\digest[72] ), .Y(_abc_15497_new_n844_));
OR2X2 OR2X2_400 ( .A(_abc_15497_new_n1951_), .B(_abc_15497_new_n1955_), .Y(_abc_15497_new_n1956_));
OR2X2 OR2X2_401 ( .A(_abc_15497_new_n699_), .B(\digest[60] ), .Y(_abc_15497_new_n1961_));
OR2X2 OR2X2_402 ( .A(_abc_15497_new_n1960_), .B(_abc_15497_new_n1962_), .Y(_0H3_reg_31_0__28_));
OR2X2 OR2X2_403 ( .A(\digest[61] ), .B(d_reg_29_), .Y(_abc_15497_new_n1967_));
OR2X2 OR2X2_404 ( .A(_abc_15497_new_n1966_), .B(_abc_15497_new_n1970_), .Y(_abc_15497_new_n1971_));
OR2X2 OR2X2_405 ( .A(_abc_15497_new_n1965_), .B(_abc_15497_new_n1972_), .Y(_abc_15497_new_n1973_));
OR2X2 OR2X2_406 ( .A(_abc_15497_new_n1975_), .B(_abc_15497_new_n1964_), .Y(_0H3_reg_31_0__29_));
OR2X2 OR2X2_407 ( .A(\digest[62] ), .B(d_reg_30_), .Y(_abc_15497_new_n1980_));
OR2X2 OR2X2_408 ( .A(_abc_15497_new_n1982_), .B(_abc_15497_new_n1968_), .Y(_abc_15497_new_n1983_));
OR2X2 OR2X2_409 ( .A(_abc_15497_new_n1985_), .B(_abc_15497_new_n1983_), .Y(_abc_15497_new_n1986_));
OR2X2 OR2X2_41 ( .A(_abc_15497_new_n847_), .B(_abc_15497_new_n800_), .Y(_abc_15497_new_n848_));
OR2X2 OR2X2_410 ( .A(_abc_15497_new_n1986_), .B(_abc_15497_new_n1981_), .Y(_abc_15497_new_n1989_));
OR2X2 OR2X2_411 ( .A(_abc_15497_new_n1991_), .B(_abc_15497_new_n1977_), .Y(_0H3_reg_31_0__30_));
OR2X2 OR2X2_412 ( .A(_abc_15497_new_n1987_), .B(_abc_15497_new_n1978_), .Y(_abc_15497_new_n1994_));
OR2X2 OR2X2_413 ( .A(\digest[63] ), .B(d_reg_31_), .Y(_abc_15497_new_n1996_));
OR2X2 OR2X2_414 ( .A(_abc_15497_new_n1995_), .B(_abc_15497_new_n2000_), .Y(_abc_15497_new_n2001_));
OR2X2 OR2X2_415 ( .A(_abc_15497_new_n1994_), .B(_abc_15497_new_n1999_), .Y(_abc_15497_new_n2002_));
OR2X2 OR2X2_416 ( .A(_abc_15497_new_n2004_), .B(_abc_15497_new_n1993_), .Y(_0H3_reg_31_0__31_));
OR2X2 OR2X2_417 ( .A(next), .B(init), .Y(_abc_15497_new_n2006_));
OR2X2 OR2X2_418 ( .A(_abc_15497_new_n2014_), .B(_abc_15497_new_n2015_), .Y(_abc_15497_new_n2016_));
OR2X2 OR2X2_419 ( .A(_abc_15497_new_n2016_), .B(_abc_15497_new_n2011_), .Y(_0e_reg_31_0__0_));
OR2X2 OR2X2_42 ( .A(_abc_15497_new_n849_), .B(_abc_15497_new_n789_), .Y(_abc_15497_new_n850_));
OR2X2 OR2X2_420 ( .A(_abc_15497_new_n2020_), .B(_abc_15497_new_n2021_), .Y(_abc_15497_new_n2022_));
OR2X2 OR2X2_421 ( .A(_abc_15497_new_n2022_), .B(_abc_15497_new_n2018_), .Y(_0e_reg_31_0__1_));
OR2X2 OR2X2_422 ( .A(_abc_15497_new_n2026_), .B(_abc_15497_new_n2027_), .Y(_abc_15497_new_n2028_));
OR2X2 OR2X2_423 ( .A(_abc_15497_new_n2028_), .B(_abc_15497_new_n2024_), .Y(_0e_reg_31_0__2_));
OR2X2 OR2X2_424 ( .A(_abc_15497_new_n2032_), .B(_abc_15497_new_n2033_), .Y(_abc_15497_new_n2034_));
OR2X2 OR2X2_425 ( .A(_abc_15497_new_n2034_), .B(_abc_15497_new_n2030_), .Y(_0e_reg_31_0__3_));
OR2X2 OR2X2_426 ( .A(_abc_15497_new_n2037_), .B(_abc_15497_new_n2038_), .Y(_abc_15497_new_n2039_));
OR2X2 OR2X2_427 ( .A(_abc_15497_new_n2039_), .B(_abc_15497_new_n2036_), .Y(_0e_reg_31_0__4_));
OR2X2 OR2X2_428 ( .A(_abc_15497_new_n2042_), .B(_abc_15497_new_n2043_), .Y(_abc_15497_new_n2044_));
OR2X2 OR2X2_429 ( .A(_abc_15497_new_n2044_), .B(_abc_15497_new_n2041_), .Y(_0e_reg_31_0__5_));
OR2X2 OR2X2_43 ( .A(_abc_15497_new_n851_), .B(_abc_15497_new_n780_), .Y(_abc_15497_new_n852_));
OR2X2 OR2X2_430 ( .A(_abc_15497_new_n2047_), .B(_abc_15497_new_n2048_), .Y(_abc_15497_new_n2049_));
OR2X2 OR2X2_431 ( .A(_abc_15497_new_n2049_), .B(_abc_15497_new_n2046_), .Y(_0e_reg_31_0__6_));
OR2X2 OR2X2_432 ( .A(_abc_15497_new_n2052_), .B(_abc_15497_new_n2053_), .Y(_abc_15497_new_n2054_));
OR2X2 OR2X2_433 ( .A(_abc_15497_new_n2054_), .B(_abc_15497_new_n2051_), .Y(_0e_reg_31_0__7_));
OR2X2 OR2X2_434 ( .A(_abc_15497_new_n2057_), .B(_abc_15497_new_n2058_), .Y(_abc_15497_new_n2059_));
OR2X2 OR2X2_435 ( .A(_abc_15497_new_n2059_), .B(_abc_15497_new_n2056_), .Y(_0e_reg_31_0__8_));
OR2X2 OR2X2_436 ( .A(_abc_15497_new_n2063_), .B(_abc_15497_new_n2064_), .Y(_abc_15497_new_n2065_));
OR2X2 OR2X2_437 ( .A(_abc_15497_new_n2065_), .B(_abc_15497_new_n2061_), .Y(_0e_reg_31_0__9_));
OR2X2 OR2X2_438 ( .A(_abc_15497_new_n2069_), .B(_abc_15497_new_n2070_), .Y(_abc_15497_new_n2071_));
OR2X2 OR2X2_439 ( .A(_abc_15497_new_n2071_), .B(_abc_15497_new_n2067_), .Y(_0e_reg_31_0__10_));
OR2X2 OR2X2_44 ( .A(c_reg_16_), .B(\digest[80] ), .Y(_abc_15497_new_n853_));
OR2X2 OR2X2_440 ( .A(_abc_15497_new_n2075_), .B(_abc_15497_new_n2076_), .Y(_abc_15497_new_n2077_));
OR2X2 OR2X2_441 ( .A(_abc_15497_new_n2077_), .B(_abc_15497_new_n2073_), .Y(_0e_reg_31_0__11_));
OR2X2 OR2X2_442 ( .A(_abc_15497_new_n2081_), .B(_abc_15497_new_n2082_), .Y(_abc_15497_new_n2083_));
OR2X2 OR2X2_443 ( .A(_abc_15497_new_n2083_), .B(_abc_15497_new_n2079_), .Y(_0e_reg_31_0__12_));
OR2X2 OR2X2_444 ( .A(_abc_15497_new_n2086_), .B(_abc_15497_new_n2087_), .Y(_abc_15497_new_n2088_));
OR2X2 OR2X2_445 ( .A(_abc_15497_new_n2088_), .B(_abc_15497_new_n2085_), .Y(_0e_reg_31_0__13_));
OR2X2 OR2X2_446 ( .A(_abc_15497_new_n2091_), .B(_abc_15497_new_n2092_), .Y(_abc_15497_new_n2093_));
OR2X2 OR2X2_447 ( .A(_abc_15497_new_n2093_), .B(_abc_15497_new_n2090_), .Y(_0e_reg_31_0__14_));
OR2X2 OR2X2_448 ( .A(_abc_15497_new_n2096_), .B(_abc_15497_new_n2097_), .Y(_abc_15497_new_n2098_));
OR2X2 OR2X2_449 ( .A(_abc_15497_new_n2098_), .B(_abc_15497_new_n2095_), .Y(_0e_reg_31_0__15_));
OR2X2 OR2X2_45 ( .A(_abc_15497_new_n858_), .B(_abc_15497_new_n757_), .Y(_abc_15497_new_n859_));
OR2X2 OR2X2_450 ( .A(_abc_15497_new_n2102_), .B(_abc_15497_new_n2103_), .Y(_abc_15497_new_n2104_));
OR2X2 OR2X2_451 ( .A(_abc_15497_new_n2104_), .B(_abc_15497_new_n2100_), .Y(_0e_reg_31_0__16_));
OR2X2 OR2X2_452 ( .A(_abc_15497_new_n2107_), .B(_abc_15497_new_n2108_), .Y(_abc_15497_new_n2109_));
OR2X2 OR2X2_453 ( .A(_abc_15497_new_n2109_), .B(_abc_15497_new_n2106_), .Y(_0e_reg_31_0__17_));
OR2X2 OR2X2_454 ( .A(_abc_15497_new_n2113_), .B(_abc_15497_new_n2114_), .Y(_abc_15497_new_n2115_));
OR2X2 OR2X2_455 ( .A(_abc_15497_new_n2115_), .B(_abc_15497_new_n2111_), .Y(_0e_reg_31_0__18_));
OR2X2 OR2X2_456 ( .A(_abc_15497_new_n2119_), .B(_abc_15497_new_n2120_), .Y(_abc_15497_new_n2121_));
OR2X2 OR2X2_457 ( .A(_abc_15497_new_n2121_), .B(_abc_15497_new_n2117_), .Y(_0e_reg_31_0__19_));
OR2X2 OR2X2_458 ( .A(_abc_15497_new_n2124_), .B(_abc_15497_new_n2125_), .Y(_abc_15497_new_n2126_));
OR2X2 OR2X2_459 ( .A(_abc_15497_new_n2126_), .B(_abc_15497_new_n2123_), .Y(_0e_reg_31_0__20_));
OR2X2 OR2X2_46 ( .A(c_reg_25_), .B(\digest[89] ), .Y(_abc_15497_new_n862_));
OR2X2 OR2X2_460 ( .A(_abc_15497_new_n2130_), .B(_abc_15497_new_n2131_), .Y(_abc_15497_new_n2132_));
OR2X2 OR2X2_461 ( .A(_abc_15497_new_n2132_), .B(_abc_15497_new_n2128_), .Y(_0e_reg_31_0__21_));
OR2X2 OR2X2_462 ( .A(_abc_15497_new_n2135_), .B(_abc_15497_new_n2136_), .Y(_abc_15497_new_n2137_));
OR2X2 OR2X2_463 ( .A(_abc_15497_new_n2137_), .B(_abc_15497_new_n2134_), .Y(_0e_reg_31_0__22_));
OR2X2 OR2X2_464 ( .A(_abc_15497_new_n2140_), .B(_abc_15497_new_n2141_), .Y(_abc_15497_new_n2142_));
OR2X2 OR2X2_465 ( .A(_abc_15497_new_n2142_), .B(_abc_15497_new_n2139_), .Y(_0e_reg_31_0__23_));
OR2X2 OR2X2_466 ( .A(_abc_15497_new_n2145_), .B(_abc_15497_new_n2146_), .Y(_abc_15497_new_n2147_));
OR2X2 OR2X2_467 ( .A(_abc_15497_new_n2147_), .B(_abc_15497_new_n2144_), .Y(_0e_reg_31_0__24_));
OR2X2 OR2X2_468 ( .A(_abc_15497_new_n2150_), .B(_abc_15497_new_n2151_), .Y(_abc_15497_new_n2152_));
OR2X2 OR2X2_469 ( .A(_abc_15497_new_n2152_), .B(_abc_15497_new_n2149_), .Y(_0e_reg_31_0__25_));
OR2X2 OR2X2_47 ( .A(c_reg_24_), .B(\digest[88] ), .Y(_abc_15497_new_n866_));
OR2X2 OR2X2_470 ( .A(_abc_15497_new_n2156_), .B(_abc_15497_new_n2157_), .Y(_abc_15497_new_n2158_));
OR2X2 OR2X2_471 ( .A(_abc_15497_new_n2158_), .B(_abc_15497_new_n2154_), .Y(_0e_reg_31_0__26_));
OR2X2 OR2X2_472 ( .A(_abc_15497_new_n2162_), .B(_abc_15497_new_n2163_), .Y(_abc_15497_new_n2164_));
OR2X2 OR2X2_473 ( .A(_abc_15497_new_n2164_), .B(_abc_15497_new_n2160_), .Y(_0e_reg_31_0__27_));
OR2X2 OR2X2_474 ( .A(_abc_15497_new_n2168_), .B(_abc_15497_new_n2169_), .Y(_abc_15497_new_n2170_));
OR2X2 OR2X2_475 ( .A(_abc_15497_new_n2170_), .B(_abc_15497_new_n2166_), .Y(_0e_reg_31_0__28_));
OR2X2 OR2X2_476 ( .A(_abc_15497_new_n2173_), .B(_abc_15497_new_n2174_), .Y(_abc_15497_new_n2175_));
OR2X2 OR2X2_477 ( .A(_abc_15497_new_n2175_), .B(_abc_15497_new_n2172_), .Y(_0e_reg_31_0__29_));
OR2X2 OR2X2_478 ( .A(_abc_15497_new_n2178_), .B(_abc_15497_new_n2179_), .Y(_abc_15497_new_n2180_));
OR2X2 OR2X2_479 ( .A(_abc_15497_new_n2180_), .B(_abc_15497_new_n2177_), .Y(_0e_reg_31_0__30_));
OR2X2 OR2X2_48 ( .A(_abc_15497_new_n870_), .B(_abc_15497_new_n860_), .Y(_abc_15497_new_n871_));
OR2X2 OR2X2_480 ( .A(_abc_15497_new_n2183_), .B(_abc_15497_new_n2184_), .Y(_abc_15497_new_n2185_));
OR2X2 OR2X2_481 ( .A(_abc_15497_new_n2185_), .B(_abc_15497_new_n2182_), .Y(_0e_reg_31_0__31_));
OR2X2 OR2X2_482 ( .A(\digest[96] ), .B(b_reg_0_), .Y(_abc_15497_new_n2187_));
OR2X2 OR2X2_483 ( .A(_abc_15497_new_n699_), .B(\digest[96] ), .Y(_abc_15497_new_n2192_));
OR2X2 OR2X2_484 ( .A(_abc_15497_new_n2191_), .B(_abc_15497_new_n2193_), .Y(_0H1_reg_31_0__0_));
OR2X2 OR2X2_485 ( .A(\digest[97] ), .B(b_reg_1_), .Y(_abc_15497_new_n2195_));
OR2X2 OR2X2_486 ( .A(_abc_15497_new_n2196_), .B(_abc_15497_new_n2197_), .Y(_abc_15497_new_n2198_));
OR2X2 OR2X2_487 ( .A(_abc_15497_new_n2198_), .B(_abc_15497_new_n2189_), .Y(_abc_15497_new_n2199_));
OR2X2 OR2X2_488 ( .A(_abc_15497_new_n2201_), .B(_abc_15497_new_n2188_), .Y(_abc_15497_new_n2202_));
OR2X2 OR2X2_489 ( .A(_abc_15497_new_n2204_), .B(_abc_15497_new_n2205_), .Y(_0H1_reg_31_0__1_));
OR2X2 OR2X2_49 ( .A(_abc_15497_new_n869_), .B(_abc_15497_new_n871_), .Y(_abc_15497_new_n872_));
OR2X2 OR2X2_490 ( .A(\digest[98] ), .B(b_reg_2_), .Y(_abc_15497_new_n2208_));
OR2X2 OR2X2_491 ( .A(_abc_15497_new_n2207_), .B(_abc_15497_new_n2212_), .Y(_abc_15497_new_n2213_));
OR2X2 OR2X2_492 ( .A(_abc_15497_new_n2214_), .B(_abc_15497_new_n2197_), .Y(_abc_15497_new_n2215_));
OR2X2 OR2X2_493 ( .A(_abc_15497_new_n2215_), .B(_abc_15497_new_n2211_), .Y(_abc_15497_new_n2216_));
OR2X2 OR2X2_494 ( .A(_abc_15497_new_n2218_), .B(_abc_15497_new_n2219_), .Y(_0H1_reg_31_0__2_));
OR2X2 OR2X2_495 ( .A(_abc_15497_new_n2221_), .B(_abc_15497_new_n2209_), .Y(_abc_15497_new_n2222_));
OR2X2 OR2X2_496 ( .A(\digest[99] ), .B(b_reg_3_), .Y(_abc_15497_new_n2223_));
OR2X2 OR2X2_497 ( .A(_abc_15497_new_n2222_), .B(_abc_15497_new_n2226_), .Y(_abc_15497_new_n2227_));
OR2X2 OR2X2_498 ( .A(_abc_15497_new_n2228_), .B(_abc_15497_new_n2229_), .Y(_abc_15497_new_n2230_));
OR2X2 OR2X2_499 ( .A(_abc_15497_new_n699_), .B(\digest[99] ), .Y(_abc_15497_new_n2233_));
OR2X2 OR2X2_5 ( .A(_abc_15497_new_n721_), .B(_abc_15497_new_n712_), .Y(_abc_15497_new_n722_));
OR2X2 OR2X2_50 ( .A(\digest[90] ), .B(c_reg_26_), .Y(_abc_15497_new_n873_));
OR2X2 OR2X2_500 ( .A(_abc_15497_new_n2232_), .B(_abc_15497_new_n2234_), .Y(_0H1_reg_31_0__3_));
OR2X2 OR2X2_501 ( .A(\digest[100] ), .B(b_reg_4_), .Y(_abc_15497_new_n2236_));
OR2X2 OR2X2_502 ( .A(_abc_15497_new_n2228_), .B(_abc_15497_new_n2241_), .Y(_abc_15497_new_n2242_));
OR2X2 OR2X2_503 ( .A(_abc_15497_new_n2243_), .B(_abc_15497_new_n2240_), .Y(_abc_15497_new_n2244_));
OR2X2 OR2X2_504 ( .A(_abc_15497_new_n2245_), .B(_abc_15497_new_n2224_), .Y(_abc_15497_new_n2246_));
OR2X2 OR2X2_505 ( .A(_abc_15497_new_n2246_), .B(_abc_15497_new_n2239_), .Y(_abc_15497_new_n2247_));
OR2X2 OR2X2_506 ( .A(_abc_15497_new_n2249_), .B(_abc_15497_new_n2250_), .Y(_0H1_reg_31_0__4_));
OR2X2 OR2X2_507 ( .A(_abc_15497_new_n2253_), .B(_abc_15497_new_n2237_), .Y(_abc_15497_new_n2254_));
OR2X2 OR2X2_508 ( .A(\digest[101] ), .B(b_reg_5_), .Y(_abc_15497_new_n2255_));
OR2X2 OR2X2_509 ( .A(_abc_15497_new_n2254_), .B(_abc_15497_new_n2258_), .Y(_abc_15497_new_n2259_));
OR2X2 OR2X2_51 ( .A(_abc_15497_new_n872_), .B(_abc_15497_new_n876_), .Y(_abc_15497_new_n877_));
OR2X2 OR2X2_510 ( .A(_abc_15497_new_n2260_), .B(_abc_15497_new_n2261_), .Y(_abc_15497_new_n2262_));
OR2X2 OR2X2_511 ( .A(_abc_15497_new_n2264_), .B(_abc_15497_new_n2252_), .Y(_0H1_reg_31_0__5_));
OR2X2 OR2X2_512 ( .A(_abc_15497_new_n2267_), .B(_abc_15497_new_n2256_), .Y(_abc_15497_new_n2268_));
OR2X2 OR2X2_513 ( .A(\digest[102] ), .B(b_reg_6_), .Y(_abc_15497_new_n2269_));
OR2X2 OR2X2_514 ( .A(_abc_15497_new_n2268_), .B(_abc_15497_new_n2272_), .Y(_abc_15497_new_n2273_));
OR2X2 OR2X2_515 ( .A(_abc_15497_new_n2274_), .B(_abc_15497_new_n2275_), .Y(_abc_15497_new_n2276_));
OR2X2 OR2X2_516 ( .A(_abc_15497_new_n2278_), .B(_abc_15497_new_n2266_), .Y(_0H1_reg_31_0__6_));
OR2X2 OR2X2_517 ( .A(_abc_15497_new_n699_), .B(\digest[103] ), .Y(_abc_15497_new_n2280_));
OR2X2 OR2X2_518 ( .A(_abc_15497_new_n2280_), .B(digest_update), .Y(_abc_15497_new_n2281_));
OR2X2 OR2X2_519 ( .A(\digest[103] ), .B(b_reg_7_), .Y(_abc_15497_new_n2283_));
OR2X2 OR2X2_52 ( .A(_abc_15497_new_n881_), .B(_abc_15497_new_n702_), .Y(_0H2_reg_31_0__26_));
OR2X2 OR2X2_520 ( .A(_abc_15497_new_n2288_), .B(_abc_15497_new_n2270_), .Y(_abc_15497_new_n2289_));
OR2X2 OR2X2_521 ( .A(_abc_15497_new_n2291_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n2292_));
OR2X2 OR2X2_522 ( .A(_abc_15497_new_n2292_), .B(_abc_15497_new_n2287_), .Y(_abc_15497_new_n2293_));
OR2X2 OR2X2_523 ( .A(\digest[104] ), .B(b_reg_8_), .Y(_abc_15497_new_n2295_));
OR2X2 OR2X2_524 ( .A(_abc_15497_new_n2299_), .B(_abc_15497_new_n2284_), .Y(_abc_15497_new_n2300_));
OR2X2 OR2X2_525 ( .A(_abc_15497_new_n2300_), .B(_abc_15497_new_n2298_), .Y(_abc_15497_new_n2301_));
OR2X2 OR2X2_526 ( .A(_abc_15497_new_n699_), .B(\digest[104] ), .Y(_abc_15497_new_n2306_));
OR2X2 OR2X2_527 ( .A(_abc_15497_new_n2305_), .B(_abc_15497_new_n2307_), .Y(_0H1_reg_31_0__8_));
OR2X2 OR2X2_528 ( .A(\digest[105] ), .B(b_reg_9_), .Y(_abc_15497_new_n2311_));
OR2X2 OR2X2_529 ( .A(_abc_15497_new_n2310_), .B(_abc_15497_new_n2314_), .Y(_abc_15497_new_n2315_));
OR2X2 OR2X2_53 ( .A(\digest[91] ), .B(c_reg_27_), .Y(_abc_15497_new_n885_));
OR2X2 OR2X2_530 ( .A(_abc_15497_new_n2309_), .B(_abc_15497_new_n2316_), .Y(_abc_15497_new_n2317_));
OR2X2 OR2X2_531 ( .A(_abc_15497_new_n699_), .B(\digest[105] ), .Y(_abc_15497_new_n2320_));
OR2X2 OR2X2_532 ( .A(_abc_15497_new_n2319_), .B(_abc_15497_new_n2321_), .Y(_0H1_reg_31_0__9_));
OR2X2 OR2X2_533 ( .A(_abc_15497_new_n2316_), .B(_abc_15497_new_n2297_), .Y(_abc_15497_new_n2326_));
OR2X2 OR2X2_534 ( .A(_abc_15497_new_n2325_), .B(_abc_15497_new_n2328_), .Y(_abc_15497_new_n2329_));
OR2X2 OR2X2_535 ( .A(\digest[106] ), .B(b_reg_10_), .Y(_abc_15497_new_n2330_));
OR2X2 OR2X2_536 ( .A(_abc_15497_new_n2329_), .B(_abc_15497_new_n2333_), .Y(_abc_15497_new_n2334_));
OR2X2 OR2X2_537 ( .A(_abc_15497_new_n2338_), .B(_abc_15497_new_n2323_), .Y(_0H1_reg_31_0__10_));
OR2X2 OR2X2_538 ( .A(\digest[107] ), .B(b_reg_11_), .Y(_abc_15497_new_n2341_));
OR2X2 OR2X2_539 ( .A(_abc_15497_new_n2348_), .B(_abc_15497_new_n2345_), .Y(_abc_15497_new_n2349_));
OR2X2 OR2X2_54 ( .A(_abc_15497_new_n884_), .B(_abc_15497_new_n888_), .Y(_abc_15497_new_n889_));
OR2X2 OR2X2_540 ( .A(_abc_15497_new_n699_), .B(\digest[107] ), .Y(_abc_15497_new_n2351_));
OR2X2 OR2X2_541 ( .A(_abc_15497_new_n2350_), .B(_abc_15497_new_n2352_), .Y(_0H1_reg_31_0__11_));
OR2X2 OR2X2_542 ( .A(\digest[108] ), .B(b_reg_12_), .Y(_abc_15497_new_n2355_));
OR2X2 OR2X2_543 ( .A(_abc_15497_new_n2359_), .B(_abc_15497_new_n2342_), .Y(_abc_15497_new_n2360_));
OR2X2 OR2X2_544 ( .A(_abc_15497_new_n2362_), .B(_abc_15497_new_n2360_), .Y(_abc_15497_new_n2363_));
OR2X2 OR2X2_545 ( .A(_abc_15497_new_n2365_), .B(_abc_15497_new_n2363_), .Y(_abc_15497_new_n2366_));
OR2X2 OR2X2_546 ( .A(_abc_15497_new_n2366_), .B(_abc_15497_new_n2358_), .Y(_abc_15497_new_n2367_));
OR2X2 OR2X2_547 ( .A(_abc_15497_new_n2371_), .B(_abc_15497_new_n2354_), .Y(_0H1_reg_31_0__12_));
OR2X2 OR2X2_548 ( .A(\digest[109] ), .B(b_reg_13_), .Y(_abc_15497_new_n2375_));
OR2X2 OR2X2_549 ( .A(_abc_15497_new_n2374_), .B(_abc_15497_new_n2378_), .Y(_abc_15497_new_n2379_));
OR2X2 OR2X2_55 ( .A(_abc_15497_new_n883_), .B(_abc_15497_new_n890_), .Y(_abc_15497_new_n891_));
OR2X2 OR2X2_550 ( .A(_abc_15497_new_n2373_), .B(_abc_15497_new_n2380_), .Y(_abc_15497_new_n2381_));
OR2X2 OR2X2_551 ( .A(_abc_15497_new_n699_), .B(\digest[109] ), .Y(_abc_15497_new_n2384_));
OR2X2 OR2X2_552 ( .A(_abc_15497_new_n2383_), .B(_abc_15497_new_n2385_), .Y(_0H1_reg_31_0__13_));
OR2X2 OR2X2_553 ( .A(\digest[110] ), .B(b_reg_14_), .Y(_abc_15497_new_n2388_));
OR2X2 OR2X2_554 ( .A(_abc_15497_new_n2394_), .B(_abc_15497_new_n2392_), .Y(_abc_15497_new_n2395_));
OR2X2 OR2X2_555 ( .A(_abc_15497_new_n2396_), .B(_abc_15497_new_n2391_), .Y(_abc_15497_new_n2397_));
OR2X2 OR2X2_556 ( .A(_abc_15497_new_n2401_), .B(_abc_15497_new_n2387_), .Y(_0H1_reg_31_0__14_));
OR2X2 OR2X2_557 ( .A(\digest[111] ), .B(b_reg_15_), .Y(_abc_15497_new_n2405_));
OR2X2 OR2X2_558 ( .A(_abc_15497_new_n2404_), .B(_abc_15497_new_n2408_), .Y(_abc_15497_new_n2409_));
OR2X2 OR2X2_559 ( .A(_abc_15497_new_n2403_), .B(_abc_15497_new_n2410_), .Y(_abc_15497_new_n2411_));
OR2X2 OR2X2_56 ( .A(_abc_15497_new_n699_), .B(\digest[91] ), .Y(_abc_15497_new_n894_));
OR2X2 OR2X2_560 ( .A(_abc_15497_new_n699_), .B(\digest[111] ), .Y(_abc_15497_new_n2414_));
OR2X2 OR2X2_561 ( .A(_abc_15497_new_n2413_), .B(_abc_15497_new_n2415_), .Y(_0H1_reg_31_0__15_));
OR2X2 OR2X2_562 ( .A(_abc_15497_new_n2417_), .B(_abc_15497_new_n2406_), .Y(_abc_15497_new_n2418_));
OR2X2 OR2X2_563 ( .A(_abc_15497_new_n2393_), .B(_abc_15497_new_n2392_), .Y(_abc_15497_new_n2420_));
OR2X2 OR2X2_564 ( .A(_abc_15497_new_n2422_), .B(_abc_15497_new_n2420_), .Y(_abc_15497_new_n2423_));
OR2X2 OR2X2_565 ( .A(_abc_15497_new_n2428_), .B(_abc_15497_new_n2425_), .Y(_abc_15497_new_n2429_));
OR2X2 OR2X2_566 ( .A(\digest[112] ), .B(b_reg_16_), .Y(_abc_15497_new_n2430_));
OR2X2 OR2X2_567 ( .A(_abc_15497_new_n2429_), .B(_abc_15497_new_n2433_), .Y(_abc_15497_new_n2434_));
OR2X2 OR2X2_568 ( .A(_abc_15497_new_n699_), .B(\digest[112] ), .Y(_abc_15497_new_n2439_));
OR2X2 OR2X2_569 ( .A(_abc_15497_new_n2438_), .B(_abc_15497_new_n2440_), .Y(_0H1_reg_31_0__16_));
OR2X2 OR2X2_57 ( .A(_abc_15497_new_n893_), .B(_abc_15497_new_n895_), .Y(_0H2_reg_31_0__27_));
OR2X2 OR2X2_570 ( .A(\digest[113] ), .B(b_reg_17_), .Y(_abc_15497_new_n2443_));
OR2X2 OR2X2_571 ( .A(_abc_15497_new_n2446_), .B(_abc_15497_new_n2431_), .Y(_abc_15497_new_n2447_));
OR2X2 OR2X2_572 ( .A(_abc_15497_new_n2435_), .B(_abc_15497_new_n2447_), .Y(_abc_15497_new_n2448_));
OR2X2 OR2X2_573 ( .A(_abc_15497_new_n2456_), .B(_abc_15497_new_n2442_), .Y(_0H1_reg_31_0__17_));
OR2X2 OR2X2_574 ( .A(\digest[114] ), .B(b_reg_18_), .Y(_abc_15497_new_n2461_));
OR2X2 OR2X2_575 ( .A(_abc_15497_new_n2460_), .B(_abc_15497_new_n2464_), .Y(_abc_15497_new_n2465_));
OR2X2 OR2X2_576 ( .A(_abc_15497_new_n699_), .B(\digest[114] ), .Y(_abc_15497_new_n2470_));
OR2X2 OR2X2_577 ( .A(_abc_15497_new_n2469_), .B(_abc_15497_new_n2471_), .Y(_0H1_reg_31_0__18_));
OR2X2 OR2X2_578 ( .A(\digest[115] ), .B(b_reg_19_), .Y(_abc_15497_new_n2474_));
OR2X2 OR2X2_579 ( .A(_abc_15497_new_n2481_), .B(_abc_15497_new_n2478_), .Y(_abc_15497_new_n2482_));
OR2X2 OR2X2_58 ( .A(_abc_15497_new_n897_), .B(_abc_15497_new_n886_), .Y(_abc_15497_new_n898_));
OR2X2 OR2X2_580 ( .A(_abc_15497_new_n699_), .B(\digest[115] ), .Y(_abc_15497_new_n2484_));
OR2X2 OR2X2_581 ( .A(_abc_15497_new_n2483_), .B(_abc_15497_new_n2485_), .Y(_0H1_reg_31_0__19_));
OR2X2 OR2X2_582 ( .A(_abc_15497_new_n2458_), .B(_abc_15497_new_n2489_), .Y(_abc_15497_new_n2490_));
OR2X2 OR2X2_583 ( .A(_abc_15497_new_n2491_), .B(_abc_15497_new_n2475_), .Y(_abc_15497_new_n2492_));
OR2X2 OR2X2_584 ( .A(_abc_15497_new_n2497_), .B(_abc_15497_new_n2495_), .Y(_abc_15497_new_n2498_));
OR2X2 OR2X2_585 ( .A(\digest[116] ), .B(b_reg_20_), .Y(_abc_15497_new_n2499_));
OR2X2 OR2X2_586 ( .A(_abc_15497_new_n2498_), .B(_abc_15497_new_n2502_), .Y(_abc_15497_new_n2503_));
OR2X2 OR2X2_587 ( .A(_abc_15497_new_n2507_), .B(_abc_15497_new_n2487_), .Y(_0H1_reg_31_0__20_));
OR2X2 OR2X2_588 ( .A(\digest[117] ), .B(b_reg_21_), .Y(_abc_15497_new_n2510_));
OR2X2 OR2X2_589 ( .A(_abc_15497_new_n2513_), .B(_abc_15497_new_n2500_), .Y(_abc_15497_new_n2514_));
OR2X2 OR2X2_59 ( .A(_abc_15497_new_n900_), .B(_abc_15497_new_n898_), .Y(_abc_15497_new_n901_));
OR2X2 OR2X2_590 ( .A(_abc_15497_new_n2504_), .B(_abc_15497_new_n2514_), .Y(_abc_15497_new_n2515_));
OR2X2 OR2X2_591 ( .A(_abc_15497_new_n2517_), .B(_abc_15497_new_n2518_), .Y(_abc_15497_new_n2519_));
OR2X2 OR2X2_592 ( .A(_abc_15497_new_n2522_), .B(_abc_15497_new_n2509_), .Y(_0H1_reg_31_0__21_));
OR2X2 OR2X2_593 ( .A(\digest[118] ), .B(b_reg_22_), .Y(_abc_15497_new_n2526_));
OR2X2 OR2X2_594 ( .A(_abc_15497_new_n2525_), .B(_abc_15497_new_n2529_), .Y(_abc_15497_new_n2530_));
OR2X2 OR2X2_595 ( .A(_abc_15497_new_n699_), .B(\digest[118] ), .Y(_abc_15497_new_n2535_));
OR2X2 OR2X2_596 ( .A(_abc_15497_new_n2534_), .B(_abc_15497_new_n2536_), .Y(_0H1_reg_31_0__22_));
OR2X2 OR2X2_597 ( .A(_abc_15497_new_n2531_), .B(_abc_15497_new_n2527_), .Y(_abc_15497_new_n2538_));
OR2X2 OR2X2_598 ( .A(\digest[119] ), .B(b_reg_23_), .Y(_abc_15497_new_n2540_));
OR2X2 OR2X2_599 ( .A(_abc_15497_new_n2544_), .B(_abc_15497_new_n2546_), .Y(_abc_15497_new_n2547_));
OR2X2 OR2X2_6 ( .A(_abc_15497_new_n723_), .B(_abc_15497_new_n704_), .Y(_abc_15497_new_n724_));
OR2X2 OR2X2_60 ( .A(\digest[92] ), .B(c_reg_28_), .Y(_abc_15497_new_n902_));
OR2X2 OR2X2_600 ( .A(_abc_15497_new_n699_), .B(\digest[119] ), .Y(_abc_15497_new_n2549_));
OR2X2 OR2X2_601 ( .A(_abc_15497_new_n2548_), .B(_abc_15497_new_n2550_), .Y(_0H1_reg_31_0__23_));
OR2X2 OR2X2_602 ( .A(_abc_15497_new_n2555_), .B(_abc_15497_new_n2541_), .Y(_abc_15497_new_n2556_));
OR2X2 OR2X2_603 ( .A(_abc_15497_new_n2518_), .B(_abc_15497_new_n2511_), .Y(_abc_15497_new_n2557_));
OR2X2 OR2X2_604 ( .A(_abc_15497_new_n2558_), .B(_abc_15497_new_n2556_), .Y(_abc_15497_new_n2559_));
OR2X2 OR2X2_605 ( .A(_abc_15497_new_n2554_), .B(_abc_15497_new_n2559_), .Y(_abc_15497_new_n2560_));
OR2X2 OR2X2_606 ( .A(_abc_15497_new_n2562_), .B(_abc_15497_new_n2560_), .Y(_abc_15497_new_n2563_));
OR2X2 OR2X2_607 ( .A(\digest[120] ), .B(b_reg_24_), .Y(_abc_15497_new_n2564_));
OR2X2 OR2X2_608 ( .A(_abc_15497_new_n2563_), .B(_abc_15497_new_n2567_), .Y(_abc_15497_new_n2568_));
OR2X2 OR2X2_609 ( .A(_abc_15497_new_n699_), .B(\digest[120] ), .Y(_abc_15497_new_n2573_));
OR2X2 OR2X2_61 ( .A(_abc_15497_new_n901_), .B(_abc_15497_new_n905_), .Y(_abc_15497_new_n906_));
OR2X2 OR2X2_610 ( .A(_abc_15497_new_n2572_), .B(_abc_15497_new_n2574_), .Y(_0H1_reg_31_0__24_));
OR2X2 OR2X2_611 ( .A(\digest[121] ), .B(b_reg_25_), .Y(_abc_15497_new_n2578_));
OR2X2 OR2X2_612 ( .A(_abc_15497_new_n2577_), .B(_abc_15497_new_n2581_), .Y(_abc_15497_new_n2582_));
OR2X2 OR2X2_613 ( .A(_abc_15497_new_n2576_), .B(_abc_15497_new_n2583_), .Y(_abc_15497_new_n2584_));
OR2X2 OR2X2_614 ( .A(_abc_15497_new_n699_), .B(\digest[121] ), .Y(_abc_15497_new_n2587_));
OR2X2 OR2X2_615 ( .A(_abc_15497_new_n2586_), .B(_abc_15497_new_n2588_), .Y(_0H1_reg_31_0__25_));
OR2X2 OR2X2_616 ( .A(_abc_15497_new_n2592_), .B(_abc_15497_new_n2579_), .Y(_abc_15497_new_n2593_));
OR2X2 OR2X2_617 ( .A(_abc_15497_new_n2591_), .B(_abc_15497_new_n2593_), .Y(_abc_15497_new_n2594_));
OR2X2 OR2X2_618 ( .A(\digest[122] ), .B(b_reg_26_), .Y(_abc_15497_new_n2595_));
OR2X2 OR2X2_619 ( .A(_abc_15497_new_n2594_), .B(_abc_15497_new_n2598_), .Y(_abc_15497_new_n2599_));
OR2X2 OR2X2_62 ( .A(_abc_15497_new_n699_), .B(\digest[92] ), .Y(_abc_15497_new_n911_));
OR2X2 OR2X2_620 ( .A(_abc_15497_new_n699_), .B(\digest[122] ), .Y(_abc_15497_new_n2604_));
OR2X2 OR2X2_621 ( .A(_abc_15497_new_n2603_), .B(_abc_15497_new_n2605_), .Y(_0H1_reg_31_0__26_));
OR2X2 OR2X2_622 ( .A(\digest[123] ), .B(b_reg_27_), .Y(_abc_15497_new_n2609_));
OR2X2 OR2X2_623 ( .A(_abc_15497_new_n2608_), .B(_abc_15497_new_n2612_), .Y(_abc_15497_new_n2613_));
OR2X2 OR2X2_624 ( .A(_abc_15497_new_n2607_), .B(_abc_15497_new_n2614_), .Y(_abc_15497_new_n2615_));
OR2X2 OR2X2_625 ( .A(_abc_15497_new_n699_), .B(\digest[123] ), .Y(_abc_15497_new_n2618_));
OR2X2 OR2X2_626 ( .A(_abc_15497_new_n2617_), .B(_abc_15497_new_n2619_), .Y(_0H1_reg_31_0__27_));
OR2X2 OR2X2_627 ( .A(_abc_15497_new_n2622_), .B(_abc_15497_new_n2610_), .Y(_abc_15497_new_n2623_));
OR2X2 OR2X2_628 ( .A(_abc_15497_new_n2625_), .B(_abc_15497_new_n2623_), .Y(_abc_15497_new_n2626_));
OR2X2 OR2X2_629 ( .A(\digest[124] ), .B(b_reg_28_), .Y(_abc_15497_new_n2627_));
OR2X2 OR2X2_63 ( .A(_abc_15497_new_n910_), .B(_abc_15497_new_n912_), .Y(_0H2_reg_31_0__28_));
OR2X2 OR2X2_630 ( .A(_abc_15497_new_n2626_), .B(_abc_15497_new_n2630_), .Y(_abc_15497_new_n2631_));
OR2X2 OR2X2_631 ( .A(_abc_15497_new_n2635_), .B(_abc_15497_new_n2621_), .Y(_0H1_reg_31_0__28_));
OR2X2 OR2X2_632 ( .A(_abc_15497_new_n699_), .B(\digest[125] ), .Y(_abc_15497_new_n2637_));
OR2X2 OR2X2_633 ( .A(_abc_15497_new_n2637_), .B(digest_update), .Y(_abc_15497_new_n2638_));
OR2X2 OR2X2_634 ( .A(_abc_15497_new_n2632_), .B(_abc_15497_new_n2628_), .Y(_abc_15497_new_n2639_));
OR2X2 OR2X2_635 ( .A(\digest[125] ), .B(b_reg_29_), .Y(_abc_15497_new_n2641_));
OR2X2 OR2X2_636 ( .A(_abc_15497_new_n2647_), .B(_abc_15497_new_n698_), .Y(_abc_15497_new_n2648_));
OR2X2 OR2X2_637 ( .A(_abc_15497_new_n2648_), .B(_abc_15497_new_n2645_), .Y(_abc_15497_new_n2649_));
OR2X2 OR2X2_638 ( .A(\digest[126] ), .B(b_reg_30_), .Y(_abc_15497_new_n2651_));
OR2X2 OR2X2_639 ( .A(_abc_15497_new_n2655_), .B(_abc_15497_new_n2642_), .Y(_abc_15497_new_n2656_));
OR2X2 OR2X2_64 ( .A(\digest[93] ), .B(c_reg_29_), .Y(_abc_15497_new_n917_));
OR2X2 OR2X2_640 ( .A(_abc_15497_new_n2658_), .B(_abc_15497_new_n2656_), .Y(_abc_15497_new_n2659_));
OR2X2 OR2X2_641 ( .A(_abc_15497_new_n2659_), .B(_abc_15497_new_n2654_), .Y(_abc_15497_new_n2660_));
OR2X2 OR2X2_642 ( .A(_abc_15497_new_n2282_), .B(_abc_15497_new_n2666_), .Y(_abc_15497_new_n2667_));
OR2X2 OR2X2_643 ( .A(_abc_15497_new_n2668_), .B(_abc_15497_new_n2669_), .Y(_abc_15497_new_n2670_));
OR2X2 OR2X2_644 ( .A(_abc_15497_new_n2671_), .B(_abc_15497_new_n2672_), .Y(_abc_15497_new_n2673_));
OR2X2 OR2X2_645 ( .A(_abc_15497_new_n2674_), .B(_abc_15497_new_n2675_), .Y(_abc_15497_new_n2676_));
OR2X2 OR2X2_646 ( .A(_abc_15497_new_n2677_), .B(_abc_15497_new_n2678_), .Y(_abc_15497_new_n2679_));
OR2X2 OR2X2_647 ( .A(_abc_15497_new_n2681_), .B(_abc_15497_new_n2682_), .Y(_abc_15497_new_n2683_));
OR2X2 OR2X2_648 ( .A(_abc_15497_new_n2684_), .B(_abc_15497_new_n2685_), .Y(_abc_15497_new_n2686_));
OR2X2 OR2X2_649 ( .A(_abc_15497_new_n2687_), .B(_abc_15497_new_n2661_), .Y(_abc_15497_new_n2688_));
OR2X2 OR2X2_65 ( .A(_abc_15497_new_n916_), .B(_abc_15497_new_n920_), .Y(_abc_15497_new_n921_));
OR2X2 OR2X2_650 ( .A(_abc_15497_new_n699_), .B(\digest[126] ), .Y(_abc_15497_new_n2691_));
OR2X2 OR2X2_651 ( .A(_abc_15497_new_n2690_), .B(_abc_15497_new_n2692_), .Y(_0H1_reg_31_0__30_));
OR2X2 OR2X2_652 ( .A(_abc_15497_new_n2694_), .B(_abc_15497_new_n2652_), .Y(_abc_15497_new_n2695_));
OR2X2 OR2X2_653 ( .A(_abc_15497_new_n2696_), .B(b_reg_31_), .Y(_abc_15497_new_n2697_));
OR2X2 OR2X2_654 ( .A(_abc_15497_new_n2698_), .B(\digest[127] ), .Y(_abc_15497_new_n2699_));
OR2X2 OR2X2_655 ( .A(_abc_15497_new_n2695_), .B(_abc_15497_new_n2701_), .Y(_abc_15497_new_n2702_));
OR2X2 OR2X2_656 ( .A(_abc_15497_new_n2703_), .B(_abc_15497_new_n2700_), .Y(_abc_15497_new_n2704_));
OR2X2 OR2X2_657 ( .A(_abc_15497_new_n699_), .B(\digest[127] ), .Y(_abc_15497_new_n2707_));
OR2X2 OR2X2_658 ( .A(_abc_15497_new_n2706_), .B(_abc_15497_new_n2708_), .Y(_0H1_reg_31_0__31_));
OR2X2 OR2X2_659 ( .A(\digest[128] ), .B(a_reg_0_), .Y(_abc_15497_new_n2710_));
OR2X2 OR2X2_66 ( .A(_abc_15497_new_n915_), .B(_abc_15497_new_n922_), .Y(_abc_15497_new_n923_));
OR2X2 OR2X2_660 ( .A(_abc_15497_new_n699_), .B(\digest[128] ), .Y(_abc_15497_new_n2715_));
OR2X2 OR2X2_661 ( .A(_abc_15497_new_n2714_), .B(_abc_15497_new_n2716_), .Y(_0H0_reg_31_0__0_));
OR2X2 OR2X2_662 ( .A(\digest[129] ), .B(a_reg_1_), .Y(_abc_15497_new_n2718_));
OR2X2 OR2X2_663 ( .A(_abc_15497_new_n2721_), .B(_abc_15497_new_n2711_), .Y(_abc_15497_new_n2724_));
OR2X2 OR2X2_664 ( .A(_abc_15497_new_n2726_), .B(_abc_15497_new_n2727_), .Y(_0H0_reg_31_0__1_));
OR2X2 OR2X2_665 ( .A(\digest[130] ), .B(a_reg_2_), .Y(_abc_15497_new_n2731_));
OR2X2 OR2X2_666 ( .A(_abc_15497_new_n2730_), .B(_abc_15497_new_n2734_), .Y(_abc_15497_new_n2735_));
OR2X2 OR2X2_667 ( .A(_abc_15497_new_n2729_), .B(_abc_15497_new_n2736_), .Y(_abc_15497_new_n2737_));
OR2X2 OR2X2_668 ( .A(_abc_15497_new_n2739_), .B(_abc_15497_new_n2740_), .Y(_0H0_reg_31_0__2_));
OR2X2 OR2X2_669 ( .A(\digest[131] ), .B(a_reg_3_), .Y(_abc_15497_new_n2745_));
OR2X2 OR2X2_67 ( .A(_abc_15497_new_n925_), .B(_abc_15497_new_n914_), .Y(_0H2_reg_31_0__29_));
OR2X2 OR2X2_670 ( .A(_abc_15497_new_n2744_), .B(_abc_15497_new_n2748_), .Y(_abc_15497_new_n2749_));
OR2X2 OR2X2_671 ( .A(_abc_15497_new_n2743_), .B(_abc_15497_new_n2750_), .Y(_abc_15497_new_n2751_));
OR2X2 OR2X2_672 ( .A(_abc_15497_new_n2753_), .B(_abc_15497_new_n2742_), .Y(_0H0_reg_31_0__3_));
OR2X2 OR2X2_673 ( .A(\digest[132] ), .B(a_reg_4_), .Y(_abc_15497_new_n2755_));
OR2X2 OR2X2_674 ( .A(_abc_15497_new_n2743_), .B(_abc_15497_new_n2759_), .Y(_abc_15497_new_n2760_));
OR2X2 OR2X2_675 ( .A(_abc_15497_new_n2762_), .B(_abc_15497_new_n2758_), .Y(_abc_15497_new_n2763_));
OR2X2 OR2X2_676 ( .A(_abc_15497_new_n2761_), .B(_abc_15497_new_n2764_), .Y(_abc_15497_new_n2765_));
OR2X2 OR2X2_677 ( .A(_abc_15497_new_n2767_), .B(_abc_15497_new_n2768_), .Y(_0H0_reg_31_0__4_));
OR2X2 OR2X2_678 ( .A(\digest[133] ), .B(a_reg_5_), .Y(_abc_15497_new_n2773_));
OR2X2 OR2X2_679 ( .A(_abc_15497_new_n2772_), .B(_abc_15497_new_n2776_), .Y(_abc_15497_new_n2777_));
OR2X2 OR2X2_68 ( .A(\digest[94] ), .B(c_reg_30_), .Y(_abc_15497_new_n930_));
OR2X2 OR2X2_680 ( .A(_abc_15497_new_n2771_), .B(_abc_15497_new_n2778_), .Y(_abc_15497_new_n2779_));
OR2X2 OR2X2_681 ( .A(_abc_15497_new_n2781_), .B(_abc_15497_new_n2770_), .Y(_0H0_reg_31_0__5_));
OR2X2 OR2X2_682 ( .A(\digest[134] ), .B(a_reg_6_), .Y(_abc_15497_new_n2786_));
OR2X2 OR2X2_683 ( .A(_abc_15497_new_n2785_), .B(_abc_15497_new_n2789_), .Y(_abc_15497_new_n2790_));
OR2X2 OR2X2_684 ( .A(_abc_15497_new_n2784_), .B(_abc_15497_new_n2791_), .Y(_abc_15497_new_n2792_));
OR2X2 OR2X2_685 ( .A(_abc_15497_new_n2794_), .B(_abc_15497_new_n2783_), .Y(_0H0_reg_31_0__6_));
OR2X2 OR2X2_686 ( .A(\digest[135] ), .B(a_reg_7_), .Y(_abc_15497_new_n2798_));
OR2X2 OR2X2_687 ( .A(_abc_15497_new_n2801_), .B(_abc_15497_new_n2787_), .Y(_abc_15497_new_n2802_));
OR2X2 OR2X2_688 ( .A(_abc_15497_new_n2797_), .B(_abc_15497_new_n2802_), .Y(_abc_15497_new_n2803_));
OR2X2 OR2X2_689 ( .A(_abc_15497_new_n2792_), .B(_abc_15497_new_n2804_), .Y(_abc_15497_new_n2805_));
OR2X2 OR2X2_69 ( .A(_abc_15497_new_n933_), .B(_abc_15497_new_n918_), .Y(_abc_15497_new_n934_));
OR2X2 OR2X2_690 ( .A(_abc_15497_new_n2810_), .B(_abc_15497_new_n2796_), .Y(_0H0_reg_31_0__7_));
OR2X2 OR2X2_691 ( .A(_abc_15497_new_n2806_), .B(_abc_15497_new_n2799_), .Y(_abc_15497_new_n2813_));
OR2X2 OR2X2_692 ( .A(_abc_15497_new_n2812_), .B(_abc_15497_new_n2813_), .Y(_abc_15497_new_n2814_));
OR2X2 OR2X2_693 ( .A(\digest[136] ), .B(a_reg_8_), .Y(_abc_15497_new_n2815_));
OR2X2 OR2X2_694 ( .A(_abc_15497_new_n2814_), .B(_abc_15497_new_n2818_), .Y(_abc_15497_new_n2819_));
OR2X2 OR2X2_695 ( .A(_abc_15497_new_n699_), .B(\digest[136] ), .Y(_abc_15497_new_n2824_));
OR2X2 OR2X2_696 ( .A(_abc_15497_new_n2823_), .B(_abc_15497_new_n2825_), .Y(_0H0_reg_31_0__8_));
OR2X2 OR2X2_697 ( .A(\digest[137] ), .B(a_reg_9_), .Y(_abc_15497_new_n2829_));
OR2X2 OR2X2_698 ( .A(_abc_15497_new_n2828_), .B(_abc_15497_new_n2832_), .Y(_abc_15497_new_n2833_));
OR2X2 OR2X2_699 ( .A(_abc_15497_new_n2827_), .B(_abc_15497_new_n2834_), .Y(_abc_15497_new_n2835_));
OR2X2 OR2X2_7 ( .A(c_reg_20_), .B(\digest[84] ), .Y(_abc_15497_new_n727_));
OR2X2 OR2X2_70 ( .A(_abc_15497_new_n949_), .B(_abc_15497_new_n818_), .Y(_abc_15497_new_n950_));
OR2X2 OR2X2_700 ( .A(_abc_15497_new_n699_), .B(\digest[137] ), .Y(_abc_15497_new_n2838_));
OR2X2 OR2X2_701 ( .A(_abc_15497_new_n2837_), .B(_abc_15497_new_n2839_), .Y(_0H0_reg_31_0__9_));
OR2X2 OR2X2_702 ( .A(\digest[138] ), .B(a_reg_10_), .Y(_abc_15497_new_n2842_));
OR2X2 OR2X2_703 ( .A(_abc_15497_new_n2834_), .B(_abc_15497_new_n2817_), .Y(_abc_15497_new_n2846_));
OR2X2 OR2X2_704 ( .A(_abc_15497_new_n2850_), .B(_abc_15497_new_n2848_), .Y(_abc_15497_new_n2851_));
OR2X2 OR2X2_705 ( .A(_abc_15497_new_n2851_), .B(_abc_15497_new_n2845_), .Y(_abc_15497_new_n2852_));
OR2X2 OR2X2_706 ( .A(_abc_15497_new_n2856_), .B(_abc_15497_new_n2841_), .Y(_0H0_reg_31_0__10_));
OR2X2 OR2X2_707 ( .A(\digest[139] ), .B(a_reg_11_), .Y(_abc_15497_new_n2861_));
OR2X2 OR2X2_708 ( .A(_abc_15497_new_n2860_), .B(_abc_15497_new_n2864_), .Y(_abc_15497_new_n2865_));
OR2X2 OR2X2_709 ( .A(_abc_15497_new_n2859_), .B(_abc_15497_new_n2866_), .Y(_abc_15497_new_n2867_));
OR2X2 OR2X2_71 ( .A(_abc_15497_new_n950_), .B(_abc_15497_new_n948_), .Y(_abc_15497_new_n951_));
OR2X2 OR2X2_710 ( .A(_abc_15497_new_n2869_), .B(_abc_15497_new_n2858_), .Y(_0H0_reg_31_0__11_));
OR2X2 OR2X2_711 ( .A(_abc_15497_new_n2866_), .B(_abc_15497_new_n2844_), .Y(_abc_15497_new_n2877_));
OR2X2 OR2X2_712 ( .A(_abc_15497_new_n2874_), .B(_abc_15497_new_n2880_), .Y(_abc_15497_new_n2881_));
OR2X2 OR2X2_713 ( .A(\digest[140] ), .B(a_reg_12_), .Y(_abc_15497_new_n2882_));
OR2X2 OR2X2_714 ( .A(_abc_15497_new_n2881_), .B(_abc_15497_new_n2885_), .Y(_abc_15497_new_n2886_));
OR2X2 OR2X2_715 ( .A(_abc_15497_new_n2890_), .B(_abc_15497_new_n2871_), .Y(_0H0_reg_31_0__12_));
OR2X2 OR2X2_716 ( .A(\digest[141] ), .B(a_reg_13_), .Y(_abc_15497_new_n2894_));
OR2X2 OR2X2_717 ( .A(_abc_15497_new_n2893_), .B(_abc_15497_new_n2897_), .Y(_abc_15497_new_n2898_));
OR2X2 OR2X2_718 ( .A(_abc_15497_new_n2892_), .B(_abc_15497_new_n2899_), .Y(_abc_15497_new_n2900_));
OR2X2 OR2X2_719 ( .A(_abc_15497_new_n699_), .B(\digest[141] ), .Y(_abc_15497_new_n2903_));
OR2X2 OR2X2_72 ( .A(_abc_15497_new_n952_), .B(_abc_15497_new_n953_), .Y(_abc_15497_new_n954_));
OR2X2 OR2X2_720 ( .A(_abc_15497_new_n2902_), .B(_abc_15497_new_n2904_), .Y(_0H0_reg_31_0__13_));
OR2X2 OR2X2_721 ( .A(\digest[142] ), .B(a_reg_14_), .Y(_abc_15497_new_n2907_));
OR2X2 OR2X2_722 ( .A(_abc_15497_new_n2913_), .B(_abc_15497_new_n2911_), .Y(_abc_15497_new_n2914_));
OR2X2 OR2X2_723 ( .A(_abc_15497_new_n2915_), .B(_abc_15497_new_n2910_), .Y(_abc_15497_new_n2916_));
OR2X2 OR2X2_724 ( .A(_abc_15497_new_n2920_), .B(_abc_15497_new_n2906_), .Y(_0H0_reg_31_0__14_));
OR2X2 OR2X2_725 ( .A(\digest[143] ), .B(a_reg_15_), .Y(_abc_15497_new_n2925_));
OR2X2 OR2X2_726 ( .A(_abc_15497_new_n2924_), .B(_abc_15497_new_n2928_), .Y(_abc_15497_new_n2929_));
OR2X2 OR2X2_727 ( .A(_abc_15497_new_n2923_), .B(_abc_15497_new_n2930_), .Y(_abc_15497_new_n2931_));
OR2X2 OR2X2_728 ( .A(_abc_15497_new_n2933_), .B(_abc_15497_new_n2922_), .Y(_0H0_reg_31_0__15_));
OR2X2 OR2X2_729 ( .A(_abc_15497_new_n2935_), .B(_abc_15497_new_n2926_), .Y(_abc_15497_new_n2936_));
OR2X2 OR2X2_73 ( .A(_abc_15497_new_n955_), .B(_abc_15497_new_n947_), .Y(_abc_15497_new_n956_));
OR2X2 OR2X2_730 ( .A(_abc_15497_new_n2912_), .B(_abc_15497_new_n2911_), .Y(_abc_15497_new_n2938_));
OR2X2 OR2X2_731 ( .A(_abc_15497_new_n2940_), .B(_abc_15497_new_n2938_), .Y(_abc_15497_new_n2941_));
OR2X2 OR2X2_732 ( .A(_abc_15497_new_n2946_), .B(_abc_15497_new_n2943_), .Y(_abc_15497_new_n2947_));
OR2X2 OR2X2_733 ( .A(\digest[144] ), .B(a_reg_16_), .Y(_abc_15497_new_n2948_));
OR2X2 OR2X2_734 ( .A(_abc_15497_new_n2947_), .B(_abc_15497_new_n2951_), .Y(_abc_15497_new_n2952_));
OR2X2 OR2X2_735 ( .A(_abc_15497_new_n699_), .B(\digest[144] ), .Y(_abc_15497_new_n2957_));
OR2X2 OR2X2_736 ( .A(_abc_15497_new_n2956_), .B(_abc_15497_new_n2958_), .Y(_0H0_reg_31_0__16_));
OR2X2 OR2X2_737 ( .A(\digest[145] ), .B(a_reg_17_), .Y(_abc_15497_new_n2961_));
OR2X2 OR2X2_738 ( .A(_abc_15497_new_n2964_), .B(_abc_15497_new_n2949_), .Y(_abc_15497_new_n2965_));
OR2X2 OR2X2_739 ( .A(_abc_15497_new_n2953_), .B(_abc_15497_new_n2965_), .Y(_abc_15497_new_n2966_));
OR2X2 OR2X2_74 ( .A(_abc_15497_new_n957_), .B(_abc_15497_new_n958_), .Y(_abc_15497_new_n959_));
OR2X2 OR2X2_740 ( .A(_abc_15497_new_n2974_), .B(_abc_15497_new_n2960_), .Y(_0H0_reg_31_0__17_));
OR2X2 OR2X2_741 ( .A(\digest[146] ), .B(a_reg_18_), .Y(_abc_15497_new_n2979_));
OR2X2 OR2X2_742 ( .A(_abc_15497_new_n2978_), .B(_abc_15497_new_n2982_), .Y(_abc_15497_new_n2983_));
OR2X2 OR2X2_743 ( .A(_abc_15497_new_n699_), .B(\digest[146] ), .Y(_abc_15497_new_n2988_));
OR2X2 OR2X2_744 ( .A(_abc_15497_new_n2987_), .B(_abc_15497_new_n2989_), .Y(_0H0_reg_31_0__18_));
OR2X2 OR2X2_745 ( .A(\digest[147] ), .B(a_reg_19_), .Y(_abc_15497_new_n2994_));
OR2X2 OR2X2_746 ( .A(_abc_15497_new_n2993_), .B(_abc_15497_new_n2997_), .Y(_abc_15497_new_n2998_));
OR2X2 OR2X2_747 ( .A(_abc_15497_new_n2992_), .B(_abc_15497_new_n2999_), .Y(_abc_15497_new_n3000_));
OR2X2 OR2X2_748 ( .A(_abc_15497_new_n3002_), .B(_abc_15497_new_n2991_), .Y(_0H0_reg_31_0__19_));
OR2X2 OR2X2_749 ( .A(_abc_15497_new_n3010_), .B(_abc_15497_new_n2995_), .Y(_abc_15497_new_n3011_));
OR2X2 OR2X2_75 ( .A(_abc_15497_new_n960_), .B(_abc_15497_new_n945_), .Y(_abc_15497_new_n961_));
OR2X2 OR2X2_750 ( .A(_abc_15497_new_n3009_), .B(_abc_15497_new_n3011_), .Y(_abc_15497_new_n3012_));
OR2X2 OR2X2_751 ( .A(_abc_15497_new_n3007_), .B(_abc_15497_new_n3012_), .Y(_abc_15497_new_n3013_));
OR2X2 OR2X2_752 ( .A(\digest[148] ), .B(a_reg_20_), .Y(_abc_15497_new_n3014_));
OR2X2 OR2X2_753 ( .A(_abc_15497_new_n3013_), .B(_abc_15497_new_n3017_), .Y(_abc_15497_new_n3018_));
OR2X2 OR2X2_754 ( .A(_abc_15497_new_n3022_), .B(_abc_15497_new_n3004_), .Y(_0H0_reg_31_0__20_));
OR2X2 OR2X2_755 ( .A(\digest[149] ), .B(a_reg_21_), .Y(_abc_15497_new_n3025_));
OR2X2 OR2X2_756 ( .A(_abc_15497_new_n3028_), .B(_abc_15497_new_n3015_), .Y(_abc_15497_new_n3029_));
OR2X2 OR2X2_757 ( .A(_abc_15497_new_n3019_), .B(_abc_15497_new_n3029_), .Y(_abc_15497_new_n3030_));
OR2X2 OR2X2_758 ( .A(_abc_15497_new_n3032_), .B(_abc_15497_new_n3033_), .Y(_abc_15497_new_n3034_));
OR2X2 OR2X2_759 ( .A(_abc_15497_new_n3037_), .B(_abc_15497_new_n3024_), .Y(_0H0_reg_31_0__21_));
OR2X2 OR2X2_76 ( .A(_abc_15497_new_n962_), .B(_abc_15497_new_n943_), .Y(_abc_15497_new_n963_));
OR2X2 OR2X2_760 ( .A(\digest[150] ), .B(a_reg_22_), .Y(_abc_15497_new_n3041_));
OR2X2 OR2X2_761 ( .A(_abc_15497_new_n3040_), .B(_abc_15497_new_n3044_), .Y(_abc_15497_new_n3045_));
OR2X2 OR2X2_762 ( .A(_abc_15497_new_n699_), .B(\digest[150] ), .Y(_abc_15497_new_n3050_));
OR2X2 OR2X2_763 ( .A(_abc_15497_new_n3049_), .B(_abc_15497_new_n3051_), .Y(_0H0_reg_31_0__22_));
OR2X2 OR2X2_764 ( .A(\digest[151] ), .B(a_reg_23_), .Y(_abc_15497_new_n3056_));
OR2X2 OR2X2_765 ( .A(_abc_15497_new_n3055_), .B(_abc_15497_new_n3059_), .Y(_abc_15497_new_n3060_));
OR2X2 OR2X2_766 ( .A(_abc_15497_new_n3054_), .B(_abc_15497_new_n3061_), .Y(_abc_15497_new_n3062_));
OR2X2 OR2X2_767 ( .A(_abc_15497_new_n3064_), .B(_abc_15497_new_n3053_), .Y(_0H0_reg_31_0__23_));
OR2X2 OR2X2_768 ( .A(_abc_15497_new_n3033_), .B(_abc_15497_new_n3026_), .Y(_abc_15497_new_n3066_));
OR2X2 OR2X2_769 ( .A(_abc_15497_new_n3069_), .B(_abc_15497_new_n3057_), .Y(_abc_15497_new_n3070_));
OR2X2 OR2X2_77 ( .A(_abc_15497_new_n964_), .B(_abc_15497_new_n965_), .Y(_abc_15497_new_n966_));
OR2X2 OR2X2_770 ( .A(_abc_15497_new_n3068_), .B(_abc_15497_new_n3070_), .Y(_abc_15497_new_n3071_));
OR2X2 OR2X2_771 ( .A(_abc_15497_new_n3073_), .B(_abc_15497_new_n3071_), .Y(_abc_15497_new_n3074_));
OR2X2 OR2X2_772 ( .A(\digest[152] ), .B(a_reg_24_), .Y(_abc_15497_new_n3075_));
OR2X2 OR2X2_773 ( .A(_abc_15497_new_n3074_), .B(_abc_15497_new_n3078_), .Y(_abc_15497_new_n3079_));
OR2X2 OR2X2_774 ( .A(_abc_15497_new_n699_), .B(\digest[152] ), .Y(_abc_15497_new_n3084_));
OR2X2 OR2X2_775 ( .A(_abc_15497_new_n3083_), .B(_abc_15497_new_n3085_), .Y(_0H0_reg_31_0__24_));
OR2X2 OR2X2_776 ( .A(\digest[153] ), .B(a_reg_25_), .Y(_abc_15497_new_n3089_));
OR2X2 OR2X2_777 ( .A(_abc_15497_new_n3088_), .B(_abc_15497_new_n3092_), .Y(_abc_15497_new_n3093_));
OR2X2 OR2X2_778 ( .A(_abc_15497_new_n3087_), .B(_abc_15497_new_n3094_), .Y(_abc_15497_new_n3095_));
OR2X2 OR2X2_779 ( .A(_abc_15497_new_n699_), .B(\digest[153] ), .Y(_abc_15497_new_n3098_));
OR2X2 OR2X2_78 ( .A(_abc_15497_new_n967_), .B(_abc_15497_new_n940_), .Y(_abc_15497_new_n968_));
OR2X2 OR2X2_780 ( .A(_abc_15497_new_n3097_), .B(_abc_15497_new_n3099_), .Y(_0H0_reg_31_0__25_));
OR2X2 OR2X2_781 ( .A(_abc_15497_new_n3103_), .B(_abc_15497_new_n3090_), .Y(_abc_15497_new_n3104_));
OR2X2 OR2X2_782 ( .A(_abc_15497_new_n3102_), .B(_abc_15497_new_n3104_), .Y(_abc_15497_new_n3105_));
OR2X2 OR2X2_783 ( .A(\digest[154] ), .B(a_reg_26_), .Y(_abc_15497_new_n3106_));
OR2X2 OR2X2_784 ( .A(_abc_15497_new_n3105_), .B(_abc_15497_new_n3109_), .Y(_abc_15497_new_n3110_));
OR2X2 OR2X2_785 ( .A(_abc_15497_new_n699_), .B(\digest[154] ), .Y(_abc_15497_new_n3115_));
OR2X2 OR2X2_786 ( .A(_abc_15497_new_n3114_), .B(_abc_15497_new_n3116_), .Y(_0H0_reg_31_0__26_));
OR2X2 OR2X2_787 ( .A(\digest[155] ), .B(a_reg_27_), .Y(_abc_15497_new_n3119_));
OR2X2 OR2X2_788 ( .A(_abc_15497_new_n3122_), .B(_abc_15497_new_n3107_), .Y(_abc_15497_new_n3123_));
OR2X2 OR2X2_789 ( .A(_abc_15497_new_n3111_), .B(_abc_15497_new_n3123_), .Y(_abc_15497_new_n3124_));
OR2X2 OR2X2_79 ( .A(_abc_15497_new_n969_), .B(_abc_15497_new_n938_), .Y(_abc_15497_new_n970_));
OR2X2 OR2X2_790 ( .A(_abc_15497_new_n3126_), .B(_abc_15497_new_n3125_), .Y(_abc_15497_new_n3127_));
OR2X2 OR2X2_791 ( .A(_abc_15497_new_n3129_), .B(_abc_15497_new_n3118_), .Y(_0H0_reg_31_0__27_));
OR2X2 OR2X2_792 ( .A(_abc_15497_new_n3134_), .B(_abc_15497_new_n3141_), .Y(_abc_15497_new_n3142_));
OR2X2 OR2X2_793 ( .A(\digest[156] ), .B(a_reg_28_), .Y(_abc_15497_new_n3143_));
OR2X2 OR2X2_794 ( .A(_abc_15497_new_n3142_), .B(_abc_15497_new_n3146_), .Y(_abc_15497_new_n3147_));
OR2X2 OR2X2_795 ( .A(_abc_15497_new_n3151_), .B(_abc_15497_new_n3131_), .Y(_0H0_reg_31_0__28_));
OR2X2 OR2X2_796 ( .A(\digest[157] ), .B(a_reg_29_), .Y(_abc_15497_new_n3154_));
OR2X2 OR2X2_797 ( .A(_abc_15497_new_n3153_), .B(_abc_15497_new_n3158_), .Y(_abc_15497_new_n3159_));
OR2X2 OR2X2_798 ( .A(_abc_15497_new_n3160_), .B(_abc_15497_new_n3157_), .Y(_abc_15497_new_n3161_));
OR2X2 OR2X2_799 ( .A(_abc_15497_new_n699_), .B(\digest[157] ), .Y(_abc_15497_new_n3164_));
OR2X2 OR2X2_8 ( .A(c_reg_19_), .B(\digest[83] ), .Y(_abc_15497_new_n733_));
OR2X2 OR2X2_80 ( .A(_abc_15497_new_n971_), .B(_abc_15497_new_n972_), .Y(_abc_15497_new_n973_));
OR2X2 OR2X2_800 ( .A(_abc_15497_new_n3163_), .B(_abc_15497_new_n3165_), .Y(_0H0_reg_31_0__29_));
OR2X2 OR2X2_801 ( .A(\digest[158] ), .B(a_reg_30_), .Y(_abc_15497_new_n3167_));
OR2X2 OR2X2_802 ( .A(_abc_15497_new_n3171_), .B(_abc_15497_new_n3155_), .Y(_abc_15497_new_n3172_));
OR2X2 OR2X2_803 ( .A(_abc_15497_new_n3174_), .B(_abc_15497_new_n3172_), .Y(_abc_15497_new_n3175_));
OR2X2 OR2X2_804 ( .A(_abc_15497_new_n3175_), .B(_abc_15497_new_n3170_), .Y(_abc_15497_new_n3176_));
OR2X2 OR2X2_805 ( .A(_abc_15497_new_n699_), .B(\digest[158] ), .Y(_abc_15497_new_n3181_));
OR2X2 OR2X2_806 ( .A(_abc_15497_new_n3180_), .B(_abc_15497_new_n3182_), .Y(_0H0_reg_31_0__30_));
OR2X2 OR2X2_807 ( .A(_abc_15497_new_n3177_), .B(_abc_15497_new_n3168_), .Y(_abc_15497_new_n3185_));
OR2X2 OR2X2_808 ( .A(\digest[159] ), .B(a_reg_31_), .Y(_abc_15497_new_n3187_));
OR2X2 OR2X2_809 ( .A(_abc_15497_new_n3186_), .B(_abc_15497_new_n3191_), .Y(_abc_15497_new_n3192_));
OR2X2 OR2X2_81 ( .A(_abc_15497_new_n974_), .B(_abc_15497_new_n975_), .Y(_abc_15497_new_n976_));
OR2X2 OR2X2_810 ( .A(_abc_15497_new_n3185_), .B(_abc_15497_new_n3190_), .Y(_abc_15497_new_n3193_));
OR2X2 OR2X2_811 ( .A(_abc_15497_new_n3195_), .B(_abc_15497_new_n3184_), .Y(_0H0_reg_31_0__31_));
OR2X2 OR2X2_812 ( .A(_abc_15497_new_n3198_), .B(_abc_15497_new_n3199_), .Y(_abc_15497_new_n3200_));
OR2X2 OR2X2_813 ( .A(_abc_15497_new_n3200_), .B(_abc_15497_new_n3197_), .Y(_0b_reg_31_0__0_));
OR2X2 OR2X2_814 ( .A(_abc_15497_new_n3204_), .B(_abc_15497_new_n3205_), .Y(_abc_15497_new_n3206_));
OR2X2 OR2X2_815 ( .A(_abc_15497_new_n3206_), .B(_abc_15497_new_n3202_), .Y(_0b_reg_31_0__1_));
OR2X2 OR2X2_816 ( .A(_abc_15497_new_n3210_), .B(_abc_15497_new_n3211_), .Y(_abc_15497_new_n3212_));
OR2X2 OR2X2_817 ( .A(_abc_15497_new_n3212_), .B(_abc_15497_new_n3208_), .Y(_0b_reg_31_0__2_));
OR2X2 OR2X2_818 ( .A(_abc_15497_new_n3215_), .B(_abc_15497_new_n3216_), .Y(_abc_15497_new_n3217_));
OR2X2 OR2X2_819 ( .A(_abc_15497_new_n3217_), .B(_abc_15497_new_n3214_), .Y(_0b_reg_31_0__3_));
OR2X2 OR2X2_82 ( .A(_abc_15497_new_n978_), .B(_abc_15497_new_n979_), .Y(_abc_15497_new_n980_));
OR2X2 OR2X2_820 ( .A(_abc_15497_new_n3221_), .B(_abc_15497_new_n3222_), .Y(_abc_15497_new_n3223_));
OR2X2 OR2X2_821 ( .A(_abc_15497_new_n3223_), .B(_abc_15497_new_n3219_), .Y(_0b_reg_31_0__4_));
OR2X2 OR2X2_822 ( .A(_abc_15497_new_n3227_), .B(_abc_15497_new_n3228_), .Y(_abc_15497_new_n3229_));
OR2X2 OR2X2_823 ( .A(_abc_15497_new_n3229_), .B(_abc_15497_new_n3225_), .Y(_0b_reg_31_0__5_));
OR2X2 OR2X2_824 ( .A(_abc_15497_new_n3233_), .B(_abc_15497_new_n3234_), .Y(_abc_15497_new_n3235_));
OR2X2 OR2X2_825 ( .A(_abc_15497_new_n3235_), .B(_abc_15497_new_n3231_), .Y(_0b_reg_31_0__6_));
OR2X2 OR2X2_826 ( .A(_abc_15497_new_n3238_), .B(_abc_15497_new_n3239_), .Y(_abc_15497_new_n3240_));
OR2X2 OR2X2_827 ( .A(_abc_15497_new_n3240_), .B(_abc_15497_new_n3237_), .Y(_0b_reg_31_0__7_));
OR2X2 OR2X2_828 ( .A(_abc_15497_new_n3243_), .B(_abc_15497_new_n3244_), .Y(_abc_15497_new_n3245_));
OR2X2 OR2X2_829 ( .A(_abc_15497_new_n3245_), .B(_abc_15497_new_n3242_), .Y(_0b_reg_31_0__8_));
OR2X2 OR2X2_83 ( .A(_abc_15497_new_n981_), .B(_abc_15497_new_n983_), .Y(_abc_15497_new_n984_));
OR2X2 OR2X2_830 ( .A(_abc_15497_new_n3248_), .B(_abc_15497_new_n3249_), .Y(_abc_15497_new_n3250_));
OR2X2 OR2X2_831 ( .A(_abc_15497_new_n3250_), .B(_abc_15497_new_n3247_), .Y(_0b_reg_31_0__9_));
OR2X2 OR2X2_832 ( .A(_abc_15497_new_n3254_), .B(_abc_15497_new_n3255_), .Y(_abc_15497_new_n3256_));
OR2X2 OR2X2_833 ( .A(_abc_15497_new_n3256_), .B(_abc_15497_new_n3252_), .Y(_0b_reg_31_0__10_));
OR2X2 OR2X2_834 ( .A(_abc_15497_new_n3259_), .B(_abc_15497_new_n3260_), .Y(_abc_15497_new_n3261_));
OR2X2 OR2X2_835 ( .A(_abc_15497_new_n3261_), .B(_abc_15497_new_n3258_), .Y(_0b_reg_31_0__11_));
OR2X2 OR2X2_836 ( .A(_abc_15497_new_n3265_), .B(_abc_15497_new_n3266_), .Y(_abc_15497_new_n3267_));
OR2X2 OR2X2_837 ( .A(_abc_15497_new_n3267_), .B(_abc_15497_new_n3263_), .Y(_0b_reg_31_0__12_));
OR2X2 OR2X2_838 ( .A(_abc_15497_new_n3270_), .B(_abc_15497_new_n3271_), .Y(_abc_15497_new_n3272_));
OR2X2 OR2X2_839 ( .A(_abc_15497_new_n3272_), .B(_abc_15497_new_n3269_), .Y(_0b_reg_31_0__13_));
OR2X2 OR2X2_84 ( .A(_abc_15497_new_n985_), .B(_abc_15497_new_n932_), .Y(_abc_15497_new_n986_));
OR2X2 OR2X2_840 ( .A(_abc_15497_new_n3276_), .B(_abc_15497_new_n3277_), .Y(_abc_15497_new_n3278_));
OR2X2 OR2X2_841 ( .A(_abc_15497_new_n3278_), .B(_abc_15497_new_n3274_), .Y(_0b_reg_31_0__14_));
OR2X2 OR2X2_842 ( .A(_abc_15497_new_n3281_), .B(_abc_15497_new_n3282_), .Y(_abc_15497_new_n3283_));
OR2X2 OR2X2_843 ( .A(_abc_15497_new_n3283_), .B(_abc_15497_new_n3280_), .Y(_0b_reg_31_0__15_));
OR2X2 OR2X2_844 ( .A(_abc_15497_new_n3286_), .B(_abc_15497_new_n3287_), .Y(_abc_15497_new_n3288_));
OR2X2 OR2X2_845 ( .A(_abc_15497_new_n3288_), .B(_abc_15497_new_n3285_), .Y(_0b_reg_31_0__16_));
OR2X2 OR2X2_846 ( .A(_abc_15497_new_n3292_), .B(_abc_15497_new_n3293_), .Y(_abc_15497_new_n3294_));
OR2X2 OR2X2_847 ( .A(_abc_15497_new_n3294_), .B(_abc_15497_new_n3290_), .Y(_0b_reg_31_0__17_));
OR2X2 OR2X2_848 ( .A(_abc_15497_new_n3297_), .B(_abc_15497_new_n3298_), .Y(_abc_15497_new_n3299_));
OR2X2 OR2X2_849 ( .A(_abc_15497_new_n3299_), .B(_abc_15497_new_n3296_), .Y(_0b_reg_31_0__18_));
OR2X2 OR2X2_85 ( .A(_abc_15497_new_n987_), .B(_abc_15497_new_n934_), .Y(_abc_15497_new_n988_));
OR2X2 OR2X2_850 ( .A(_abc_15497_new_n3302_), .B(_abc_15497_new_n3303_), .Y(_abc_15497_new_n3304_));
OR2X2 OR2X2_851 ( .A(_abc_15497_new_n3304_), .B(_abc_15497_new_n3301_), .Y(_0b_reg_31_0__19_));
OR2X2 OR2X2_852 ( .A(_abc_15497_new_n3308_), .B(_abc_15497_new_n3309_), .Y(_abc_15497_new_n3310_));
OR2X2 OR2X2_853 ( .A(_abc_15497_new_n3310_), .B(_abc_15497_new_n3306_), .Y(_0b_reg_31_0__20_));
OR2X2 OR2X2_854 ( .A(_abc_15497_new_n3314_), .B(_abc_15497_new_n3315_), .Y(_abc_15497_new_n3316_));
OR2X2 OR2X2_855 ( .A(_abc_15497_new_n3316_), .B(_abc_15497_new_n3312_), .Y(_0b_reg_31_0__21_));
OR2X2 OR2X2_856 ( .A(_abc_15497_new_n3319_), .B(_abc_15497_new_n3320_), .Y(_abc_15497_new_n3321_));
OR2X2 OR2X2_857 ( .A(_abc_15497_new_n3321_), .B(_abc_15497_new_n3318_), .Y(_0b_reg_31_0__22_));
OR2X2 OR2X2_858 ( .A(_abc_15497_new_n3324_), .B(_abc_15497_new_n3325_), .Y(_abc_15497_new_n3326_));
OR2X2 OR2X2_859 ( .A(_abc_15497_new_n3326_), .B(_abc_15497_new_n3323_), .Y(_0b_reg_31_0__23_));
OR2X2 OR2X2_86 ( .A(_abc_15497_new_n988_), .B(_abc_15497_new_n931_), .Y(_abc_15497_new_n989_));
OR2X2 OR2X2_860 ( .A(_abc_15497_new_n3329_), .B(_abc_15497_new_n3330_), .Y(_abc_15497_new_n3331_));
OR2X2 OR2X2_861 ( .A(_abc_15497_new_n3331_), .B(_abc_15497_new_n3328_), .Y(_0b_reg_31_0__24_));
OR2X2 OR2X2_862 ( .A(_abc_15497_new_n3334_), .B(_abc_15497_new_n3335_), .Y(_abc_15497_new_n3336_));
OR2X2 OR2X2_863 ( .A(_abc_15497_new_n3336_), .B(_abc_15497_new_n3333_), .Y(_0b_reg_31_0__25_));
OR2X2 OR2X2_864 ( .A(_abc_15497_new_n3339_), .B(_abc_15497_new_n3340_), .Y(_abc_15497_new_n3341_));
OR2X2 OR2X2_865 ( .A(_abc_15497_new_n3341_), .B(_abc_15497_new_n3338_), .Y(_0b_reg_31_0__26_));
OR2X2 OR2X2_866 ( .A(_abc_15497_new_n3344_), .B(_abc_15497_new_n3345_), .Y(_abc_15497_new_n3346_));
OR2X2 OR2X2_867 ( .A(_abc_15497_new_n3346_), .B(_abc_15497_new_n3343_), .Y(_0b_reg_31_0__27_));
OR2X2 OR2X2_868 ( .A(_abc_15497_new_n3350_), .B(_abc_15497_new_n3351_), .Y(_abc_15497_new_n3352_));
OR2X2 OR2X2_869 ( .A(_abc_15497_new_n3352_), .B(_abc_15497_new_n3348_), .Y(_0b_reg_31_0__28_));
OR2X2 OR2X2_87 ( .A(_abc_15497_new_n991_), .B(_abc_15497_new_n927_), .Y(_0H2_reg_31_0__30_));
OR2X2 OR2X2_870 ( .A(_abc_15497_new_n3355_), .B(_abc_15497_new_n3356_), .Y(_abc_15497_new_n3357_));
OR2X2 OR2X2_871 ( .A(_abc_15497_new_n3357_), .B(_abc_15497_new_n3354_), .Y(_0b_reg_31_0__29_));
OR2X2 OR2X2_872 ( .A(_abc_15497_new_n3360_), .B(_abc_15497_new_n3361_), .Y(_abc_15497_new_n3362_));
OR2X2 OR2X2_873 ( .A(_abc_15497_new_n3362_), .B(_abc_15497_new_n3359_), .Y(_0b_reg_31_0__30_));
OR2X2 OR2X2_874 ( .A(_abc_15497_new_n3365_), .B(_abc_15497_new_n3366_), .Y(_abc_15497_new_n3367_));
OR2X2 OR2X2_875 ( .A(_abc_15497_new_n3367_), .B(_abc_15497_new_n3364_), .Y(_0b_reg_31_0__31_));
OR2X2 OR2X2_876 ( .A(_abc_15497_new_n3371_), .B(_abc_15497_new_n3372_), .Y(_abc_15497_new_n3373_));
OR2X2 OR2X2_877 ( .A(_abc_15497_new_n3373_), .B(_abc_15497_new_n3369_), .Y(_0d_reg_31_0__0_));
OR2X2 OR2X2_878 ( .A(_abc_15497_new_n3376_), .B(_abc_15497_new_n3377_), .Y(_abc_15497_new_n3378_));
OR2X2 OR2X2_879 ( .A(_abc_15497_new_n3378_), .B(_abc_15497_new_n3375_), .Y(_0d_reg_31_0__1_));
OR2X2 OR2X2_88 ( .A(_abc_15497_new_n993_), .B(_abc_15497_new_n928_), .Y(_abc_15497_new_n994_));
OR2X2 OR2X2_880 ( .A(_abc_15497_new_n3381_), .B(_abc_15497_new_n3382_), .Y(_abc_15497_new_n3383_));
OR2X2 OR2X2_881 ( .A(_abc_15497_new_n3383_), .B(_abc_15497_new_n3380_), .Y(_0d_reg_31_0__2_));
OR2X2 OR2X2_882 ( .A(_abc_15497_new_n3387_), .B(_abc_15497_new_n3388_), .Y(_abc_15497_new_n3389_));
OR2X2 OR2X2_883 ( .A(_abc_15497_new_n3389_), .B(_abc_15497_new_n3385_), .Y(_0d_reg_31_0__3_));
OR2X2 OR2X2_884 ( .A(_abc_15497_new_n3392_), .B(_abc_15497_new_n3393_), .Y(_abc_15497_new_n3394_));
OR2X2 OR2X2_885 ( .A(_abc_15497_new_n3394_), .B(_abc_15497_new_n3391_), .Y(_0d_reg_31_0__4_));
OR2X2 OR2X2_886 ( .A(_abc_15497_new_n3397_), .B(_abc_15497_new_n3398_), .Y(_abc_15497_new_n3399_));
OR2X2 OR2X2_887 ( .A(_abc_15497_new_n3399_), .B(_abc_15497_new_n3396_), .Y(_0d_reg_31_0__5_));
OR2X2 OR2X2_888 ( .A(_abc_15497_new_n3402_), .B(_abc_15497_new_n3403_), .Y(_abc_15497_new_n3404_));
OR2X2 OR2X2_889 ( .A(_abc_15497_new_n3404_), .B(_abc_15497_new_n3401_), .Y(_0d_reg_31_0__6_));
OR2X2 OR2X2_89 ( .A(_abc_15497_new_n995_), .B(c_reg_31_), .Y(_abc_15497_new_n996_));
OR2X2 OR2X2_890 ( .A(_abc_15497_new_n3408_), .B(_abc_15497_new_n3409_), .Y(_abc_15497_new_n3410_));
OR2X2 OR2X2_891 ( .A(_abc_15497_new_n3410_), .B(_abc_15497_new_n3406_), .Y(_0d_reg_31_0__7_));
OR2X2 OR2X2_892 ( .A(_abc_15497_new_n3414_), .B(_abc_15497_new_n3415_), .Y(_abc_15497_new_n3416_));
OR2X2 OR2X2_893 ( .A(_abc_15497_new_n3416_), .B(_abc_15497_new_n3412_), .Y(_0d_reg_31_0__8_));
OR2X2 OR2X2_894 ( .A(_abc_15497_new_n3420_), .B(_abc_15497_new_n3421_), .Y(_abc_15497_new_n3422_));
OR2X2 OR2X2_895 ( .A(_abc_15497_new_n3422_), .B(_abc_15497_new_n3418_), .Y(_0d_reg_31_0__9_));
OR2X2 OR2X2_896 ( .A(_abc_15497_new_n3425_), .B(_abc_15497_new_n3426_), .Y(_abc_15497_new_n3427_));
OR2X2 OR2X2_897 ( .A(_abc_15497_new_n3427_), .B(_abc_15497_new_n3424_), .Y(_0d_reg_31_0__10_));
OR2X2 OR2X2_898 ( .A(_abc_15497_new_n3431_), .B(_abc_15497_new_n3432_), .Y(_abc_15497_new_n3433_));
OR2X2 OR2X2_899 ( .A(_abc_15497_new_n3433_), .B(_abc_15497_new_n3429_), .Y(_0d_reg_31_0__11_));
OR2X2 OR2X2_9 ( .A(c_reg_18_), .B(\digest[82] ), .Y(_abc_15497_new_n737_));
OR2X2 OR2X2_90 ( .A(_abc_15497_new_n997_), .B(\digest[95] ), .Y(_abc_15497_new_n998_));
OR2X2 OR2X2_900 ( .A(_abc_15497_new_n3436_), .B(_abc_15497_new_n3437_), .Y(_abc_15497_new_n3438_));
OR2X2 OR2X2_901 ( .A(_abc_15497_new_n3438_), .B(_abc_15497_new_n3435_), .Y(_0d_reg_31_0__12_));
OR2X2 OR2X2_902 ( .A(_abc_15497_new_n3442_), .B(_abc_15497_new_n3443_), .Y(_abc_15497_new_n3444_));
OR2X2 OR2X2_903 ( .A(_abc_15497_new_n3444_), .B(_abc_15497_new_n3440_), .Y(_0d_reg_31_0__13_));
OR2X2 OR2X2_904 ( .A(_abc_15497_new_n3447_), .B(_abc_15497_new_n3448_), .Y(_abc_15497_new_n3449_));
OR2X2 OR2X2_905 ( .A(_abc_15497_new_n3449_), .B(_abc_15497_new_n3446_), .Y(_0d_reg_31_0__14_));
OR2X2 OR2X2_906 ( .A(_abc_15497_new_n3453_), .B(_abc_15497_new_n3454_), .Y(_abc_15497_new_n3455_));
OR2X2 OR2X2_907 ( .A(_abc_15497_new_n3455_), .B(_abc_15497_new_n3451_), .Y(_0d_reg_31_0__15_));
OR2X2 OR2X2_908 ( .A(_abc_15497_new_n3459_), .B(_abc_15497_new_n3460_), .Y(_abc_15497_new_n3461_));
OR2X2 OR2X2_909 ( .A(_abc_15497_new_n3461_), .B(_abc_15497_new_n3457_), .Y(_0d_reg_31_0__16_));
OR2X2 OR2X2_91 ( .A(_abc_15497_new_n994_), .B(_abc_15497_new_n1000_), .Y(_abc_15497_new_n1001_));
OR2X2 OR2X2_910 ( .A(_abc_15497_new_n3464_), .B(_abc_15497_new_n3465_), .Y(_abc_15497_new_n3466_));
OR2X2 OR2X2_911 ( .A(_abc_15497_new_n3466_), .B(_abc_15497_new_n3463_), .Y(_0d_reg_31_0__17_));
OR2X2 OR2X2_912 ( .A(_abc_15497_new_n3470_), .B(_abc_15497_new_n3471_), .Y(_abc_15497_new_n3472_));
OR2X2 OR2X2_913 ( .A(_abc_15497_new_n3472_), .B(_abc_15497_new_n3468_), .Y(_0d_reg_31_0__18_));
OR2X2 OR2X2_914 ( .A(_abc_15497_new_n3476_), .B(_abc_15497_new_n3477_), .Y(_abc_15497_new_n3478_));
OR2X2 OR2X2_915 ( .A(_abc_15497_new_n3478_), .B(_abc_15497_new_n3474_), .Y(_0d_reg_31_0__19_));
OR2X2 OR2X2_916 ( .A(_abc_15497_new_n3481_), .B(_abc_15497_new_n3482_), .Y(_abc_15497_new_n3483_));
OR2X2 OR2X2_917 ( .A(_abc_15497_new_n3483_), .B(_abc_15497_new_n3480_), .Y(_0d_reg_31_0__20_));
OR2X2 OR2X2_918 ( .A(_abc_15497_new_n3486_), .B(_abc_15497_new_n3487_), .Y(_abc_15497_new_n3488_));
OR2X2 OR2X2_919 ( .A(_abc_15497_new_n3488_), .B(_abc_15497_new_n3485_), .Y(_0d_reg_31_0__21_));
OR2X2 OR2X2_92 ( .A(_abc_15497_new_n1002_), .B(_abc_15497_new_n999_), .Y(_abc_15497_new_n1003_));
OR2X2 OR2X2_920 ( .A(_abc_15497_new_n3492_), .B(_abc_15497_new_n3493_), .Y(_abc_15497_new_n3494_));
OR2X2 OR2X2_921 ( .A(_abc_15497_new_n3494_), .B(_abc_15497_new_n3490_), .Y(_0d_reg_31_0__22_));
OR2X2 OR2X2_922 ( .A(_abc_15497_new_n3498_), .B(_abc_15497_new_n3499_), .Y(_abc_15497_new_n3500_));
OR2X2 OR2X2_923 ( .A(_abc_15497_new_n3500_), .B(_abc_15497_new_n3496_), .Y(_0d_reg_31_0__23_));
OR2X2 OR2X2_924 ( .A(_abc_15497_new_n3504_), .B(_abc_15497_new_n3505_), .Y(_abc_15497_new_n3506_));
OR2X2 OR2X2_925 ( .A(_abc_15497_new_n3506_), .B(_abc_15497_new_n3502_), .Y(_0d_reg_31_0__24_));
OR2X2 OR2X2_926 ( .A(_abc_15497_new_n3510_), .B(_abc_15497_new_n3511_), .Y(_abc_15497_new_n3512_));
OR2X2 OR2X2_927 ( .A(_abc_15497_new_n3512_), .B(_abc_15497_new_n3508_), .Y(_0d_reg_31_0__25_));
OR2X2 OR2X2_928 ( .A(_abc_15497_new_n3516_), .B(_abc_15497_new_n3517_), .Y(_abc_15497_new_n3518_));
OR2X2 OR2X2_929 ( .A(_abc_15497_new_n3518_), .B(_abc_15497_new_n3514_), .Y(_0d_reg_31_0__26_));
OR2X2 OR2X2_93 ( .A(_abc_15497_new_n699_), .B(\digest[95] ), .Y(_abc_15497_new_n1006_));
OR2X2 OR2X2_930 ( .A(_abc_15497_new_n3522_), .B(_abc_15497_new_n3523_), .Y(_abc_15497_new_n3524_));
OR2X2 OR2X2_931 ( .A(_abc_15497_new_n3524_), .B(_abc_15497_new_n3520_), .Y(_0d_reg_31_0__27_));
OR2X2 OR2X2_932 ( .A(_abc_15497_new_n3527_), .B(_abc_15497_new_n3528_), .Y(_abc_15497_new_n3529_));
OR2X2 OR2X2_933 ( .A(_abc_15497_new_n3529_), .B(_abc_15497_new_n3526_), .Y(_0d_reg_31_0__28_));
OR2X2 OR2X2_934 ( .A(_abc_15497_new_n3533_), .B(_abc_15497_new_n3534_), .Y(_abc_15497_new_n3535_));
OR2X2 OR2X2_935 ( .A(_abc_15497_new_n3535_), .B(_abc_15497_new_n3531_), .Y(_0d_reg_31_0__29_));
OR2X2 OR2X2_936 ( .A(_abc_15497_new_n3539_), .B(_abc_15497_new_n3540_), .Y(_abc_15497_new_n3541_));
OR2X2 OR2X2_937 ( .A(_abc_15497_new_n3541_), .B(_abc_15497_new_n3537_), .Y(_0d_reg_31_0__30_));
OR2X2 OR2X2_938 ( .A(_abc_15497_new_n3545_), .B(_abc_15497_new_n3546_), .Y(_abc_15497_new_n3547_));
OR2X2 OR2X2_939 ( .A(_abc_15497_new_n3547_), .B(_abc_15497_new_n3543_), .Y(_0d_reg_31_0__31_));
OR2X2 OR2X2_94 ( .A(_abc_15497_new_n1005_), .B(_abc_15497_new_n1007_), .Y(_0H2_reg_31_0__31_));
OR2X2 OR2X2_940 ( .A(_abc_15497_new_n3551_), .B(_abc_15497_new_n3552_), .Y(_abc_15497_new_n3553_));
OR2X2 OR2X2_941 ( .A(_abc_15497_new_n3553_), .B(_abc_15497_new_n3549_), .Y(_0c_reg_31_0__0_));
OR2X2 OR2X2_942 ( .A(_abc_15497_new_n699_), .B(\digest[65] ), .Y(_abc_15497_new_n3556_));
OR2X2 OR2X2_943 ( .A(_abc_15497_new_n3557_), .B(_abc_15497_new_n3558_), .Y(_abc_15497_new_n3559_));
OR2X2 OR2X2_944 ( .A(_abc_15497_new_n3559_), .B(_abc_15497_new_n3555_), .Y(_0c_reg_31_0__1_));
OR2X2 OR2X2_945 ( .A(_abc_15497_new_n699_), .B(\digest[66] ), .Y(_abc_15497_new_n3562_));
OR2X2 OR2X2_946 ( .A(_abc_15497_new_n3563_), .B(_abc_15497_new_n3564_), .Y(_abc_15497_new_n3565_));
OR2X2 OR2X2_947 ( .A(_abc_15497_new_n3565_), .B(_abc_15497_new_n3561_), .Y(_0c_reg_31_0__2_));
OR2X2 OR2X2_948 ( .A(_abc_15497_new_n699_), .B(\digest[67] ), .Y(_abc_15497_new_n3568_));
OR2X2 OR2X2_949 ( .A(_abc_15497_new_n3569_), .B(_abc_15497_new_n3570_), .Y(_abc_15497_new_n3571_));
OR2X2 OR2X2_95 ( .A(e_reg_0_), .B(\digest[0] ), .Y(_abc_15497_new_n1011_));
OR2X2 OR2X2_950 ( .A(_abc_15497_new_n3571_), .B(_abc_15497_new_n3567_), .Y(_0c_reg_31_0__3_));
OR2X2 OR2X2_951 ( .A(_abc_15497_new_n699_), .B(\digest[68] ), .Y(_abc_15497_new_n3574_));
OR2X2 OR2X2_952 ( .A(_abc_15497_new_n3575_), .B(_abc_15497_new_n3576_), .Y(_abc_15497_new_n3577_));
OR2X2 OR2X2_953 ( .A(_abc_15497_new_n3577_), .B(_abc_15497_new_n3573_), .Y(_0c_reg_31_0__4_));
OR2X2 OR2X2_954 ( .A(_abc_15497_new_n699_), .B(\digest[69] ), .Y(_abc_15497_new_n3580_));
OR2X2 OR2X2_955 ( .A(_abc_15497_new_n3581_), .B(_abc_15497_new_n3582_), .Y(_abc_15497_new_n3583_));
OR2X2 OR2X2_956 ( .A(_abc_15497_new_n3583_), .B(_abc_15497_new_n3579_), .Y(_0c_reg_31_0__5_));
OR2X2 OR2X2_957 ( .A(_abc_15497_new_n699_), .B(\digest[70] ), .Y(_abc_15497_new_n3586_));
OR2X2 OR2X2_958 ( .A(_abc_15497_new_n3587_), .B(_abc_15497_new_n3588_), .Y(_abc_15497_new_n3589_));
OR2X2 OR2X2_959 ( .A(_abc_15497_new_n3589_), .B(_abc_15497_new_n3585_), .Y(_0c_reg_31_0__6_));
OR2X2 OR2X2_96 ( .A(_abc_15497_new_n1014_), .B(_abc_15497_new_n1013_), .Y(_0H4_reg_31_0__0_));
OR2X2 OR2X2_960 ( .A(_abc_15497_new_n699_), .B(\digest[71] ), .Y(_abc_15497_new_n3592_));
OR2X2 OR2X2_961 ( .A(_abc_15497_new_n3593_), .B(_abc_15497_new_n3594_), .Y(_abc_15497_new_n3595_));
OR2X2 OR2X2_962 ( .A(_abc_15497_new_n3595_), .B(_abc_15497_new_n3591_), .Y(_0c_reg_31_0__7_));
OR2X2 OR2X2_963 ( .A(_abc_15497_new_n3599_), .B(_abc_15497_new_n3600_), .Y(_abc_15497_new_n3601_));
OR2X2 OR2X2_964 ( .A(_abc_15497_new_n3601_), .B(_abc_15497_new_n3597_), .Y(_0c_reg_31_0__8_));
OR2X2 OR2X2_965 ( .A(_abc_15497_new_n3605_), .B(_abc_15497_new_n3606_), .Y(_abc_15497_new_n3607_));
OR2X2 OR2X2_966 ( .A(_abc_15497_new_n3607_), .B(_abc_15497_new_n3603_), .Y(_0c_reg_31_0__9_));
OR2X2 OR2X2_967 ( .A(_abc_15497_new_n699_), .B(\digest[74] ), .Y(_abc_15497_new_n3610_));
OR2X2 OR2X2_968 ( .A(_abc_15497_new_n3611_), .B(_abc_15497_new_n3612_), .Y(_abc_15497_new_n3613_));
OR2X2 OR2X2_969 ( .A(_abc_15497_new_n3613_), .B(_abc_15497_new_n3609_), .Y(_0c_reg_31_0__10_));
OR2X2 OR2X2_97 ( .A(e_reg_1_), .B(\digest[1] ), .Y(_abc_15497_new_n1016_));
OR2X2 OR2X2_970 ( .A(_abc_15497_new_n699_), .B(\digest[75] ), .Y(_abc_15497_new_n3616_));
OR2X2 OR2X2_971 ( .A(_abc_15497_new_n3617_), .B(_abc_15497_new_n3618_), .Y(_abc_15497_new_n3619_));
OR2X2 OR2X2_972 ( .A(_abc_15497_new_n3619_), .B(_abc_15497_new_n3615_), .Y(_0c_reg_31_0__11_));
OR2X2 OR2X2_973 ( .A(_abc_15497_new_n699_), .B(\digest[76] ), .Y(_abc_15497_new_n3622_));
OR2X2 OR2X2_974 ( .A(_abc_15497_new_n3623_), .B(_abc_15497_new_n3624_), .Y(_abc_15497_new_n3625_));
OR2X2 OR2X2_975 ( .A(_abc_15497_new_n3625_), .B(_abc_15497_new_n3621_), .Y(_0c_reg_31_0__12_));
OR2X2 OR2X2_976 ( .A(_abc_15497_new_n3629_), .B(_abc_15497_new_n3630_), .Y(_abc_15497_new_n3631_));
OR2X2 OR2X2_977 ( .A(_abc_15497_new_n3631_), .B(_abc_15497_new_n3627_), .Y(_0c_reg_31_0__13_));
OR2X2 OR2X2_978 ( .A(_abc_15497_new_n699_), .B(\digest[78] ), .Y(_abc_15497_new_n3634_));
OR2X2 OR2X2_979 ( .A(_abc_15497_new_n3635_), .B(_abc_15497_new_n3636_), .Y(_abc_15497_new_n3637_));
OR2X2 OR2X2_98 ( .A(_abc_15497_new_n1017_), .B(_abc_15497_new_n1018_), .Y(_abc_15497_new_n1019_));
OR2X2 OR2X2_980 ( .A(_abc_15497_new_n3637_), .B(_abc_15497_new_n3633_), .Y(_0c_reg_31_0__14_));
OR2X2 OR2X2_981 ( .A(_abc_15497_new_n699_), .B(\digest[79] ), .Y(_abc_15497_new_n3640_));
OR2X2 OR2X2_982 ( .A(_abc_15497_new_n3641_), .B(_abc_15497_new_n3642_), .Y(_abc_15497_new_n3643_));
OR2X2 OR2X2_983 ( .A(_abc_15497_new_n3643_), .B(_abc_15497_new_n3639_), .Y(_0c_reg_31_0__15_));
OR2X2 OR2X2_984 ( .A(_abc_15497_new_n3647_), .B(_abc_15497_new_n3648_), .Y(_abc_15497_new_n3649_));
OR2X2 OR2X2_985 ( .A(_abc_15497_new_n3649_), .B(_abc_15497_new_n3645_), .Y(_0c_reg_31_0__16_));
OR2X2 OR2X2_986 ( .A(_abc_15497_new_n699_), .B(\digest[81] ), .Y(_abc_15497_new_n3652_));
OR2X2 OR2X2_987 ( .A(_abc_15497_new_n3653_), .B(_abc_15497_new_n3654_), .Y(_abc_15497_new_n3655_));
OR2X2 OR2X2_988 ( .A(_abc_15497_new_n3655_), .B(_abc_15497_new_n3651_), .Y(_0c_reg_31_0__17_));
OR2X2 OR2X2_989 ( .A(_abc_15497_new_n3659_), .B(_abc_15497_new_n3660_), .Y(_abc_15497_new_n3661_));
OR2X2 OR2X2_99 ( .A(_abc_15497_new_n1019_), .B(_abc_15497_new_n1010_), .Y(_abc_15497_new_n1020_));
OR2X2 OR2X2_990 ( .A(_abc_15497_new_n3661_), .B(_abc_15497_new_n3657_), .Y(_0c_reg_31_0__18_));
OR2X2 OR2X2_991 ( .A(_abc_15497_new_n699_), .B(\digest[83] ), .Y(_abc_15497_new_n3664_));
OR2X2 OR2X2_992 ( .A(_abc_15497_new_n3665_), .B(_abc_15497_new_n3666_), .Y(_abc_15497_new_n3667_));
OR2X2 OR2X2_993 ( .A(_abc_15497_new_n3667_), .B(_abc_15497_new_n3663_), .Y(_0c_reg_31_0__19_));
OR2X2 OR2X2_994 ( .A(_abc_15497_new_n699_), .B(\digest[84] ), .Y(_abc_15497_new_n3670_));
OR2X2 OR2X2_995 ( .A(_abc_15497_new_n3671_), .B(_abc_15497_new_n3672_), .Y(_abc_15497_new_n3673_));
OR2X2 OR2X2_996 ( .A(_abc_15497_new_n3673_), .B(_abc_15497_new_n3669_), .Y(_0c_reg_31_0__20_));
OR2X2 OR2X2_997 ( .A(_abc_15497_new_n699_), .B(\digest[85] ), .Y(_abc_15497_new_n3676_));
OR2X2 OR2X2_998 ( .A(_abc_15497_new_n3677_), .B(_abc_15497_new_n3678_), .Y(_abc_15497_new_n3679_));
OR2X2 OR2X2_999 ( .A(_abc_15497_new_n3679_), .B(_abc_15497_new_n3675_), .Y(_0c_reg_31_0__21_));


endmodule