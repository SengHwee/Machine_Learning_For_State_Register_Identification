
module mc_top(clk_i, rst_i, \wb_data_i[0] , \wb_data_i[1] , \wb_data_i[2] , \wb_data_i[3] , \wb_data_i[4] , \wb_data_i[5] , \wb_data_i[6] , \wb_data_i[7] , \wb_data_i[8] , \wb_data_i[9] , \wb_data_i[10] , \wb_data_i[11] , \wb_data_i[12] , \wb_data_i[13] , \wb_data_i[14] , \wb_data_i[15] , \wb_data_i[16] , \wb_data_i[17] , \wb_data_i[18] , \wb_data_i[19] , \wb_data_i[20] , \wb_data_i[21] , \wb_data_i[22] , \wb_data_i[23] , \wb_data_i[24] , \wb_data_i[25] , \wb_data_i[26] , \wb_data_i[27] , \wb_data_i[28] , \wb_data_i[29] , \wb_data_i[30] , \wb_data_i[31] , \wb_addr_i[0] , \wb_addr_i[1] , \wb_addr_i[2] , \wb_addr_i[3] , \wb_addr_i[4] , \wb_addr_i[5] , \wb_addr_i[6] , \wb_addr_i[7] , \wb_addr_i[8] , \wb_addr_i[9] , \wb_addr_i[10] , \wb_addr_i[11] , \wb_addr_i[12] , \wb_addr_i[13] , \wb_addr_i[14] , \wb_addr_i[15] , \wb_addr_i[16] , \wb_addr_i[17] , \wb_addr_i[18] , \wb_addr_i[19] , \wb_addr_i[20] , \wb_addr_i[21] , \wb_addr_i[22] , \wb_addr_i[23] , \wb_addr_i[24] , \wb_addr_i[25] , \wb_addr_i[26] , \wb_addr_i[27] , \wb_addr_i[28] , \wb_addr_i[29] , \wb_addr_i[30] , \wb_addr_i[31] , \wb_sel_i[0] , \wb_sel_i[1] , \wb_sel_i[2] , \wb_sel_i[3] , wb_we_i, wb_cyc_i, wb_stb_i, susp_req_i, resume_req_i, mc_clk_i, mc_br_pad_i, mc_ack_pad_i, \mc_data_pad_i[0] , \mc_data_pad_i[1] , \mc_data_pad_i[2] , \mc_data_pad_i[3] , \mc_data_pad_i[4] , \mc_data_pad_i[5] , \mc_data_pad_i[6] , \mc_data_pad_i[7] , \mc_data_pad_i[8] , \mc_data_pad_i[9] , \mc_data_pad_i[10] , \mc_data_pad_i[11] , \mc_data_pad_i[12] , \mc_data_pad_i[13] , \mc_data_pad_i[14] , \mc_data_pad_i[15] , \mc_data_pad_i[16] , \mc_data_pad_i[17] , \mc_data_pad_i[18] , \mc_data_pad_i[19] , \mc_data_pad_i[20] , \mc_data_pad_i[21] , \mc_data_pad_i[22] , \mc_data_pad_i[23] , \mc_data_pad_i[24] , \mc_data_pad_i[25] , \mc_data_pad_i[26] , \mc_data_pad_i[27] , \mc_data_pad_i[28] , \mc_data_pad_i[29] , \mc_data_pad_i[30] , \mc_data_pad_i[31] , \mc_dp_pad_i[0] , \mc_dp_pad_i[1] , \mc_dp_pad_i[2] , \mc_dp_pad_i[3] , mc_sts_pad_i, \wb_data_o[0] , \wb_data_o[1] , \wb_data_o[2] , \wb_data_o[3] , \wb_data_o[4] , \wb_data_o[5] , \wb_data_o[6] , \wb_data_o[7] , \wb_data_o[8] , \wb_data_o[9] , \wb_data_o[10] , \wb_data_o[11] , \wb_data_o[12] , \wb_data_o[13] , \wb_data_o[14] , \wb_data_o[15] , \wb_data_o[16] , \wb_data_o[17] , \wb_data_o[18] , \wb_data_o[19] , \wb_data_o[20] , \wb_data_o[21] , \wb_data_o[22] , \wb_data_o[23] , \wb_data_o[24] , \wb_data_o[25] , \wb_data_o[26] , \wb_data_o[27] , \wb_data_o[28] , \wb_data_o[29] , \wb_data_o[30] , \wb_data_o[31] , wb_ack_o, wb_err_o, suspended_o, \poc_o[0] , \poc_o[1] , \poc_o[2] , \poc_o[3] , \poc_o[4] , \poc_o[5] , \poc_o[6] , \poc_o[7] , \poc_o[8] , \poc_o[9] , \poc_o[10] , \poc_o[11] , \poc_o[12] , \poc_o[13] , \poc_o[14] , \poc_o[15] , \poc_o[16] , \poc_o[17] , \poc_o[18] , \poc_o[19] , \poc_o[20] , \poc_o[21] , \poc_o[22] , \poc_o[23] , \poc_o[24] , \poc_o[25] , \poc_o[26] , \poc_o[27] , \poc_o[28] , \poc_o[29] , \poc_o[30] , \poc_o[31] , mc_bg_pad_o, \mc_addr_pad_o[0] , \mc_addr_pad_o[1] , \mc_addr_pad_o[2] , \mc_addr_pad_o[3] , \mc_addr_pad_o[4] , \mc_addr_pad_o[5] , \mc_addr_pad_o[6] , \mc_addr_pad_o[7] , \mc_addr_pad_o[8] , \mc_addr_pad_o[9] , \mc_addr_pad_o[10] , \mc_addr_pad_o[11] , \mc_addr_pad_o[12] , \mc_addr_pad_o[13] , \mc_addr_pad_o[14] , \mc_addr_pad_o[15] , \mc_addr_pad_o[16] , \mc_addr_pad_o[17] , \mc_addr_pad_o[18] , \mc_addr_pad_o[19] , \mc_addr_pad_o[20] , \mc_addr_pad_o[21] , \mc_addr_pad_o[22] , \mc_addr_pad_o[23] , \mc_data_pad_o[0] , \mc_data_pad_o[1] , \mc_data_pad_o[2] , \mc_data_pad_o[3] , \mc_data_pad_o[4] , \mc_data_pad_o[5] , \mc_data_pad_o[6] , \mc_data_pad_o[7] , \mc_data_pad_o[8] , \mc_data_pad_o[9] , \mc_data_pad_o[10] , \mc_data_pad_o[11] , \mc_data_pad_o[12] , \mc_data_pad_o[13] , \mc_data_pad_o[14] , \mc_data_pad_o[15] , \mc_data_pad_o[16] , \mc_data_pad_o[17] , \mc_data_pad_o[18] , \mc_data_pad_o[19] , \mc_data_pad_o[20] , \mc_data_pad_o[21] , \mc_data_pad_o[22] , \mc_data_pad_o[23] , \mc_data_pad_o[24] , \mc_data_pad_o[25] , \mc_data_pad_o[26] , \mc_data_pad_o[27] , \mc_data_pad_o[28] , \mc_data_pad_o[29] , \mc_data_pad_o[30] , \mc_data_pad_o[31] , \mc_dp_pad_o[0] , \mc_dp_pad_o[1] , \mc_dp_pad_o[2] , \mc_dp_pad_o[3] , mc_doe_pad_doe_o, \mc_dqm_pad_o[0] , \mc_dqm_pad_o[1] , \mc_dqm_pad_o[2] , \mc_dqm_pad_o[3] , mc_oe_pad_o_, mc_we_pad_o_, mc_cas_pad_o_, mc_ras_pad_o_, mc_cke_pad_o_, \mc_cs_pad_o_[0] , \mc_cs_pad_o_[1] , \mc_cs_pad_o_[2] , \mc_cs_pad_o_[3] , \mc_cs_pad_o_[4] , \mc_cs_pad_o_[5] , \mc_cs_pad_o_[6] , \mc_cs_pad_o_[7] , mc_rp_pad_o_, mc_vpen_pad_o, mc_adsc_pad_o_, mc_adv_pad_o_, mc_zz_pad_o, mc_coe_pad_coe_o);
  wire _abc_55805_n237_1;
  wire _abc_55805_n238_1;
  wire _abc_55805_n239_1;
  wire _abc_55805_n240;
  wire _abc_55805_n240_bF_buf0;
  wire _abc_55805_n240_bF_buf1;
  wire _abc_55805_n240_bF_buf2;
  wire _abc_55805_n240_bF_buf3;
  wire _abc_55805_n240_bF_buf4;
  wire _abc_55805_n240_bF_buf5;
  wire _abc_55805_n241_1;
  wire _abc_55805_n242_1;
  wire _abc_55805_n243;
  wire _abc_55805_n244_1;
  wire _abc_55805_n245_1;
  wire _abc_55805_n246;
  wire _abc_55805_n248;
  wire _abc_55805_n249;
  wire _abc_55805_n250;
  wire _abc_55805_n251;
  wire _abc_55805_n252;
  wire _abc_55805_n254;
  wire _abc_55805_n255;
  wire _abc_55805_n256;
  wire _abc_55805_n257;
  wire _abc_55805_n258;
  wire _abc_55805_n260;
  wire _abc_55805_n261;
  wire _abc_55805_n262;
  wire _abc_55805_n263;
  wire _abc_55805_n264;
  wire _abc_55805_n266;
  wire _abc_55805_n267;
  wire _abc_55805_n268;
  wire _abc_55805_n269;
  wire _abc_55805_n270;
  wire _abc_55805_n272;
  wire _abc_55805_n273;
  wire _abc_55805_n274;
  wire _abc_55805_n275;
  wire _abc_55805_n276;
  wire _abc_55805_n278;
  wire _abc_55805_n279;
  wire _abc_55805_n280;
  wire _abc_55805_n281;
  wire _abc_55805_n282;
  wire _abc_55805_n284;
  wire _abc_55805_n285;
  wire _abc_55805_n286;
  wire _abc_55805_n287;
  wire _abc_55805_n288;
  wire _abc_55805_n290;
  wire _abc_55805_n291;
  wire _abc_55805_n293;
  wire _abc_55805_n294;
  wire _abc_55805_n296;
  wire _abc_55805_n297;
  wire _abc_55805_n299;
  wire _abc_55805_n300;
  wire _abc_55805_n302;
  wire _abc_55805_n303;
  wire _abc_55805_n305;
  wire _abc_55805_n306;
  wire _abc_55805_n308;
  wire _abc_55805_n309;
  wire _abc_55805_n311;
  wire _abc_55805_n312;
  wire _abc_55805_n314;
  wire _abc_55805_n315;
  wire _abc_55805_n317;
  wire _abc_55805_n318;
  wire _abc_55805_n320;
  wire _abc_55805_n321;
  wire _abc_55805_n323;
  wire _abc_55805_n324;
  wire _abc_55805_n326;
  wire _abc_55805_n327;
  wire _abc_55805_n329;
  wire _abc_55805_n330;
  wire _abc_55805_n332;
  wire _abc_55805_n333;
  wire _abc_55805_n335;
  wire _abc_55805_n336;
  wire _abc_55805_n338;
  wire _abc_55805_n339;
  wire _abc_55805_n341;
  wire _abc_55805_n342;
  wire _abc_55805_n344;
  wire _abc_55805_n345;
  wire _abc_55805_n347;
  wire _abc_55805_n348;
  wire _abc_55805_n350;
  wire _abc_55805_n351;
  wire _abc_55805_n353;
  wire _abc_55805_n354;
  wire _abc_55805_n356;
  wire _abc_55805_n357;
  wire _abc_55805_n359;
  wire _abc_55805_n360;
  wire _abc_55805_n362;
  wire _abc_55805_n363;
  wire _abc_55805_n365;
  wire _abc_55805_n366;
  wire _abc_55805_n368;
  wire _abc_55805_n369;
  wire _abc_55805_n371;
  wire _abc_55805_n372;
  wire _abc_55805_n389;
  wire _abc_55805_n390;
  wire _abc_55805_n392;
  wire _abc_55805_n393;
  wire _abc_55805_n395;
  wire _abc_55805_n396;
  wire _abc_55805_n398;
  wire _abc_55805_n399;
  wire _abc_55805_n401;
  wire _abc_55805_n402;
  wire _abc_55805_n404;
  wire _abc_55805_n405;
  wire _abc_55805_n407;
  wire _abc_55805_n408;
  wire _abc_55805_n413;
  wire _abc_55805_n414;
  wire _abc_55805_n416;
  wire _abc_55805_n417;
  wire _abc_55805_n482;
  wire _abc_55805_n483;
  wire _abc_55805_n484;
  wire _auto_iopadmap_cc_313_execute_56218_0_;
  wire _auto_iopadmap_cc_313_execute_56218_10_;
  wire _auto_iopadmap_cc_313_execute_56218_11_;
  wire _auto_iopadmap_cc_313_execute_56218_12_;
  wire _auto_iopadmap_cc_313_execute_56218_13_;
  wire _auto_iopadmap_cc_313_execute_56218_14_;
  wire _auto_iopadmap_cc_313_execute_56218_15_;
  wire _auto_iopadmap_cc_313_execute_56218_16_;
  wire _auto_iopadmap_cc_313_execute_56218_17_;
  wire _auto_iopadmap_cc_313_execute_56218_18_;
  wire _auto_iopadmap_cc_313_execute_56218_19_;
  wire _auto_iopadmap_cc_313_execute_56218_1_;
  wire _auto_iopadmap_cc_313_execute_56218_20_;
  wire _auto_iopadmap_cc_313_execute_56218_21_;
  wire _auto_iopadmap_cc_313_execute_56218_22_;
  wire _auto_iopadmap_cc_313_execute_56218_23_;
  wire _auto_iopadmap_cc_313_execute_56218_2_;
  wire _auto_iopadmap_cc_313_execute_56218_3_;
  wire _auto_iopadmap_cc_313_execute_56218_4_;
  wire _auto_iopadmap_cc_313_execute_56218_5_;
  wire _auto_iopadmap_cc_313_execute_56218_6_;
  wire _auto_iopadmap_cc_313_execute_56218_7_;
  wire _auto_iopadmap_cc_313_execute_56218_8_;
  wire _auto_iopadmap_cc_313_execute_56218_9_;
  wire _auto_iopadmap_cc_313_execute_56243;
  wire _auto_iopadmap_cc_313_execute_56245;
  wire _auto_iopadmap_cc_313_execute_56247;
  wire _auto_iopadmap_cc_313_execute_56249;
  wire _auto_iopadmap_cc_313_execute_56251;
  wire _auto_iopadmap_cc_313_execute_56253;
  wire _auto_iopadmap_cc_313_execute_56255_0_;
  wire _auto_iopadmap_cc_313_execute_56255_1_;
  wire _auto_iopadmap_cc_313_execute_56255_2_;
  wire _auto_iopadmap_cc_313_execute_56255_3_;
  wire _auto_iopadmap_cc_313_execute_56255_4_;
  wire _auto_iopadmap_cc_313_execute_56255_5_;
  wire _auto_iopadmap_cc_313_execute_56255_6_;
  wire _auto_iopadmap_cc_313_execute_56255_7_;
  wire _auto_iopadmap_cc_313_execute_56264_0_;
  wire _auto_iopadmap_cc_313_execute_56264_10_;
  wire _auto_iopadmap_cc_313_execute_56264_11_;
  wire _auto_iopadmap_cc_313_execute_56264_12_;
  wire _auto_iopadmap_cc_313_execute_56264_13_;
  wire _auto_iopadmap_cc_313_execute_56264_14_;
  wire _auto_iopadmap_cc_313_execute_56264_15_;
  wire _auto_iopadmap_cc_313_execute_56264_16_;
  wire _auto_iopadmap_cc_313_execute_56264_17_;
  wire _auto_iopadmap_cc_313_execute_56264_18_;
  wire _auto_iopadmap_cc_313_execute_56264_19_;
  wire _auto_iopadmap_cc_313_execute_56264_1_;
  wire _auto_iopadmap_cc_313_execute_56264_20_;
  wire _auto_iopadmap_cc_313_execute_56264_21_;
  wire _auto_iopadmap_cc_313_execute_56264_22_;
  wire _auto_iopadmap_cc_313_execute_56264_23_;
  wire _auto_iopadmap_cc_313_execute_56264_24_;
  wire _auto_iopadmap_cc_313_execute_56264_25_;
  wire _auto_iopadmap_cc_313_execute_56264_26_;
  wire _auto_iopadmap_cc_313_execute_56264_27_;
  wire _auto_iopadmap_cc_313_execute_56264_28_;
  wire _auto_iopadmap_cc_313_execute_56264_29_;
  wire _auto_iopadmap_cc_313_execute_56264_2_;
  wire _auto_iopadmap_cc_313_execute_56264_30_;
  wire _auto_iopadmap_cc_313_execute_56264_31_;
  wire _auto_iopadmap_cc_313_execute_56264_3_;
  wire _auto_iopadmap_cc_313_execute_56264_4_;
  wire _auto_iopadmap_cc_313_execute_56264_5_;
  wire _auto_iopadmap_cc_313_execute_56264_6_;
  wire _auto_iopadmap_cc_313_execute_56264_7_;
  wire _auto_iopadmap_cc_313_execute_56264_8_;
  wire _auto_iopadmap_cc_313_execute_56264_9_;
  wire _auto_iopadmap_cc_313_execute_56297;
  wire _auto_iopadmap_cc_313_execute_56299_0_;
  wire _auto_iopadmap_cc_313_execute_56299_1_;
  wire _auto_iopadmap_cc_313_execute_56299_2_;
  wire _auto_iopadmap_cc_313_execute_56299_3_;
  wire _auto_iopadmap_cc_313_execute_56304_0_;
  wire _auto_iopadmap_cc_313_execute_56304_1_;
  wire _auto_iopadmap_cc_313_execute_56304_2_;
  wire _auto_iopadmap_cc_313_execute_56304_3_;
  wire _auto_iopadmap_cc_313_execute_56309;
  wire _auto_iopadmap_cc_313_execute_56311;
  wire _auto_iopadmap_cc_313_execute_56313;
  wire _auto_iopadmap_cc_313_execute_56315;
  wire _auto_iopadmap_cc_313_execute_56317;
  wire _auto_iopadmap_cc_313_execute_56319;
  wire _auto_iopadmap_cc_313_execute_56321_0_;
  wire _auto_iopadmap_cc_313_execute_56321_10_;
  wire _auto_iopadmap_cc_313_execute_56321_11_;
  wire _auto_iopadmap_cc_313_execute_56321_12_;
  wire _auto_iopadmap_cc_313_execute_56321_13_;
  wire _auto_iopadmap_cc_313_execute_56321_14_;
  wire _auto_iopadmap_cc_313_execute_56321_15_;
  wire _auto_iopadmap_cc_313_execute_56321_16_;
  wire _auto_iopadmap_cc_313_execute_56321_17_;
  wire _auto_iopadmap_cc_313_execute_56321_18_;
  wire _auto_iopadmap_cc_313_execute_56321_19_;
  wire _auto_iopadmap_cc_313_execute_56321_1_;
  wire _auto_iopadmap_cc_313_execute_56321_20_;
  wire _auto_iopadmap_cc_313_execute_56321_21_;
  wire _auto_iopadmap_cc_313_execute_56321_22_;
  wire _auto_iopadmap_cc_313_execute_56321_23_;
  wire _auto_iopadmap_cc_313_execute_56321_24_;
  wire _auto_iopadmap_cc_313_execute_56321_25_;
  wire _auto_iopadmap_cc_313_execute_56321_26_;
  wire _auto_iopadmap_cc_313_execute_56321_27_;
  wire _auto_iopadmap_cc_313_execute_56321_28_;
  wire _auto_iopadmap_cc_313_execute_56321_29_;
  wire _auto_iopadmap_cc_313_execute_56321_2_;
  wire _auto_iopadmap_cc_313_execute_56321_30_;
  wire _auto_iopadmap_cc_313_execute_56321_31_;
  wire _auto_iopadmap_cc_313_execute_56321_3_;
  wire _auto_iopadmap_cc_313_execute_56321_4_;
  wire _auto_iopadmap_cc_313_execute_56321_5_;
  wire _auto_iopadmap_cc_313_execute_56321_6_;
  wire _auto_iopadmap_cc_313_execute_56321_7_;
  wire _auto_iopadmap_cc_313_execute_56321_8_;
  wire _auto_iopadmap_cc_313_execute_56321_9_;
  wire _auto_iopadmap_cc_313_execute_56354;
  wire _auto_iopadmap_cc_313_execute_56356;
  wire _auto_iopadmap_cc_313_execute_56358_0_;
  wire _auto_iopadmap_cc_313_execute_56358_10_;
  wire _auto_iopadmap_cc_313_execute_56358_11_;
  wire _auto_iopadmap_cc_313_execute_56358_12_;
  wire _auto_iopadmap_cc_313_execute_56358_13_;
  wire _auto_iopadmap_cc_313_execute_56358_14_;
  wire _auto_iopadmap_cc_313_execute_56358_15_;
  wire _auto_iopadmap_cc_313_execute_56358_16_;
  wire _auto_iopadmap_cc_313_execute_56358_17_;
  wire _auto_iopadmap_cc_313_execute_56358_18_;
  wire _auto_iopadmap_cc_313_execute_56358_19_;
  wire _auto_iopadmap_cc_313_execute_56358_1_;
  wire _auto_iopadmap_cc_313_execute_56358_20_;
  wire _auto_iopadmap_cc_313_execute_56358_21_;
  wire _auto_iopadmap_cc_313_execute_56358_22_;
  wire _auto_iopadmap_cc_313_execute_56358_23_;
  wire _auto_iopadmap_cc_313_execute_56358_24_;
  wire _auto_iopadmap_cc_313_execute_56358_25_;
  wire _auto_iopadmap_cc_313_execute_56358_26_;
  wire _auto_iopadmap_cc_313_execute_56358_27_;
  wire _auto_iopadmap_cc_313_execute_56358_28_;
  wire _auto_iopadmap_cc_313_execute_56358_29_;
  wire _auto_iopadmap_cc_313_execute_56358_2_;
  wire _auto_iopadmap_cc_313_execute_56358_30_;
  wire _auto_iopadmap_cc_313_execute_56358_31_;
  wire _auto_iopadmap_cc_313_execute_56358_3_;
  wire _auto_iopadmap_cc_313_execute_56358_4_;
  wire _auto_iopadmap_cc_313_execute_56358_5_;
  wire _auto_iopadmap_cc_313_execute_56358_6_;
  wire _auto_iopadmap_cc_313_execute_56358_7_;
  wire _auto_iopadmap_cc_313_execute_56358_8_;
  wire _auto_iopadmap_cc_313_execute_56358_9_;
  wire _auto_iopadmap_cc_313_execute_56391;
  wire bank_adr_0_;
  wire bank_adr_0_bF_buf0;
  wire bank_adr_0_bF_buf1;
  wire bank_adr_0_bF_buf2;
  wire bank_adr_0_bF_buf3;
  wire bank_adr_1_;
  wire bank_adr_1_bF_buf0;
  wire bank_adr_1_bF_buf1;
  wire bank_adr_1_bF_buf2;
  wire bank_adr_1_bF_buf3;
  wire bank_clr;
  wire bank_clr_all;
  wire bank_open;
  wire bank_set;
  wire cas_;
  input clk_i;
  wire clk_i_bF_buf0;
  wire clk_i_bF_buf1;
  wire clk_i_bF_buf10;
  wire clk_i_bF_buf100;
  wire clk_i_bF_buf101;
  wire clk_i_bF_buf102;
  wire clk_i_bF_buf103;
  wire clk_i_bF_buf104;
  wire clk_i_bF_buf105;
  wire clk_i_bF_buf106;
  wire clk_i_bF_buf107;
  wire clk_i_bF_buf108;
  wire clk_i_bF_buf109;
  wire clk_i_bF_buf11;
  wire clk_i_bF_buf110;
  wire clk_i_bF_buf111;
  wire clk_i_bF_buf112;
  wire clk_i_bF_buf113;
  wire clk_i_bF_buf114;
  wire clk_i_bF_buf115;
  wire clk_i_bF_buf116;
  wire clk_i_bF_buf117;
  wire clk_i_bF_buf118;
  wire clk_i_bF_buf119;
  wire clk_i_bF_buf12;
  wire clk_i_bF_buf120;
  wire clk_i_bF_buf121;
  wire clk_i_bF_buf122;
  wire clk_i_bF_buf123;
  wire clk_i_bF_buf124;
  wire clk_i_bF_buf125;
  wire clk_i_bF_buf13;
  wire clk_i_bF_buf14;
  wire clk_i_bF_buf15;
  wire clk_i_bF_buf16;
  wire clk_i_bF_buf17;
  wire clk_i_bF_buf18;
  wire clk_i_bF_buf19;
  wire clk_i_bF_buf2;
  wire clk_i_bF_buf20;
  wire clk_i_bF_buf21;
  wire clk_i_bF_buf22;
  wire clk_i_bF_buf23;
  wire clk_i_bF_buf24;
  wire clk_i_bF_buf25;
  wire clk_i_bF_buf26;
  wire clk_i_bF_buf27;
  wire clk_i_bF_buf28;
  wire clk_i_bF_buf29;
  wire clk_i_bF_buf3;
  wire clk_i_bF_buf30;
  wire clk_i_bF_buf31;
  wire clk_i_bF_buf32;
  wire clk_i_bF_buf33;
  wire clk_i_bF_buf34;
  wire clk_i_bF_buf35;
  wire clk_i_bF_buf36;
  wire clk_i_bF_buf37;
  wire clk_i_bF_buf38;
  wire clk_i_bF_buf39;
  wire clk_i_bF_buf4;
  wire clk_i_bF_buf40;
  wire clk_i_bF_buf41;
  wire clk_i_bF_buf42;
  wire clk_i_bF_buf43;
  wire clk_i_bF_buf44;
  wire clk_i_bF_buf45;
  wire clk_i_bF_buf46;
  wire clk_i_bF_buf47;
  wire clk_i_bF_buf48;
  wire clk_i_bF_buf49;
  wire clk_i_bF_buf5;
  wire clk_i_bF_buf50;
  wire clk_i_bF_buf51;
  wire clk_i_bF_buf52;
  wire clk_i_bF_buf53;
  wire clk_i_bF_buf54;
  wire clk_i_bF_buf55;
  wire clk_i_bF_buf56;
  wire clk_i_bF_buf57;
  wire clk_i_bF_buf58;
  wire clk_i_bF_buf59;
  wire clk_i_bF_buf6;
  wire clk_i_bF_buf60;
  wire clk_i_bF_buf61;
  wire clk_i_bF_buf62;
  wire clk_i_bF_buf63;
  wire clk_i_bF_buf64;
  wire clk_i_bF_buf65;
  wire clk_i_bF_buf66;
  wire clk_i_bF_buf67;
  wire clk_i_bF_buf68;
  wire clk_i_bF_buf69;
  wire clk_i_bF_buf7;
  wire clk_i_bF_buf70;
  wire clk_i_bF_buf71;
  wire clk_i_bF_buf72;
  wire clk_i_bF_buf73;
  wire clk_i_bF_buf74;
  wire clk_i_bF_buf75;
  wire clk_i_bF_buf76;
  wire clk_i_bF_buf77;
  wire clk_i_bF_buf78;
  wire clk_i_bF_buf79;
  wire clk_i_bF_buf8;
  wire clk_i_bF_buf80;
  wire clk_i_bF_buf81;
  wire clk_i_bF_buf82;
  wire clk_i_bF_buf83;
  wire clk_i_bF_buf84;
  wire clk_i_bF_buf85;
  wire clk_i_bF_buf86;
  wire clk_i_bF_buf87;
  wire clk_i_bF_buf88;
  wire clk_i_bF_buf89;
  wire clk_i_bF_buf9;
  wire clk_i_bF_buf90;
  wire clk_i_bF_buf91;
  wire clk_i_bF_buf92;
  wire clk_i_bF_buf93;
  wire clk_i_bF_buf94;
  wire clk_i_bF_buf95;
  wire clk_i_bF_buf96;
  wire clk_i_bF_buf97;
  wire clk_i_bF_buf98;
  wire clk_i_bF_buf99;
  wire clk_i_hier0_bF_buf0;
  wire clk_i_hier0_bF_buf1;
  wire clk_i_hier0_bF_buf10;
  wire clk_i_hier0_bF_buf2;
  wire clk_i_hier0_bF_buf3;
  wire clk_i_hier0_bF_buf4;
  wire clk_i_hier0_bF_buf5;
  wire clk_i_hier0_bF_buf6;
  wire clk_i_hier0_bF_buf7;
  wire clk_i_hier0_bF_buf8;
  wire clk_i_hier0_bF_buf9;
  wire cmd_a10;
  wire cs_0_;
  wire cs_1_;
  wire cs_2_;
  wire cs_3_;
  wire cs_4_;
  wire cs_5_;
  wire cs_6_;
  wire cs_7_;
  wire cs_en;
  wire cs_le;
  wire cs_le_bF_buf0;
  wire cs_le_bF_buf1;
  wire cs_le_bF_buf2;
  wire cs_le_bF_buf3;
  wire cs_le_bF_buf4;
  wire cs_le_d;
  wire cs_need_rfr_0_;
  wire cs_need_rfr_1_;
  wire cs_need_rfr_2_;
  wire cs_need_rfr_3_;
  wire cs_need_rfr_4_;
  wire cs_need_rfr_5_;
  wire cs_need_rfr_6_;
  wire cs_need_rfr_7_;
  wire csc_10_;
  wire csc_1_;
  wire csc_2_;
  wire csc_3_;
  wire csc_4_;
  wire csc_5_;
  wire csc_5_bF_buf0;
  wire csc_5_bF_buf1;
  wire csc_5_bF_buf2;
  wire csc_5_bF_buf3;
  wire csc_5_bF_buf4;
  wire csc_6_;
  wire csc_7_;
  wire csc_9_;
  wire csc_s_1_;
  wire csc_s_2_;
  wire csc_s_2_bF_buf0;
  wire csc_s_2_bF_buf1;
  wire csc_s_2_bF_buf2;
  wire csc_s_2_bF_buf3;
  wire csc_s_2_bF_buf4;
  wire csc_s_3_;
  wire csc_s_4_;
  wire csc_s_5_;
  wire csc_s_5_bF_buf0;
  wire csc_s_5_bF_buf1;
  wire csc_s_5_bF_buf2;
  wire csc_s_5_bF_buf3;
  wire csc_s_5_bF_buf4;
  wire csc_s_6_;
  wire csc_s_7_;
  wire data_oe;
  wire dv;
  wire err;
  wire fs;
  wire init_ack;
  wire init_req;
  wire lmr_ack;
  wire lmr_req;
  wire lmr_sel;
  wire lmr_sel_bF_buf0;
  wire lmr_sel_bF_buf1;
  wire lmr_sel_bF_buf2;
  wire lmr_sel_bF_buf3;
  wire lmr_sel_bF_buf4;
  wire lmr_sel_bF_buf5;
  wire lmr_sel_bF_buf6;
  input mc_ack_pad_i;
  wire mc_ack_r;
  wire mc_addr_d_0_;
  wire mc_addr_d_10_;
  wire mc_addr_d_11_;
  wire mc_addr_d_12_;
  wire mc_addr_d_13_;
  wire mc_addr_d_14_;
  wire mc_addr_d_15_;
  wire mc_addr_d_16_;
  wire mc_addr_d_17_;
  wire mc_addr_d_18_;
  wire mc_addr_d_19_;
  wire mc_addr_d_1_;
  wire mc_addr_d_20_;
  wire mc_addr_d_21_;
  wire mc_addr_d_22_;
  wire mc_addr_d_23_;
  wire mc_addr_d_2_;
  wire mc_addr_d_3_;
  wire mc_addr_d_4_;
  wire mc_addr_d_5_;
  wire mc_addr_d_6_;
  wire mc_addr_d_7_;
  wire mc_addr_d_8_;
  wire mc_addr_d_9_;
  output \mc_addr_pad_o[0] ;
  output \mc_addr_pad_o[10] ;
  output \mc_addr_pad_o[11] ;
  output \mc_addr_pad_o[12] ;
  output \mc_addr_pad_o[13] ;
  output \mc_addr_pad_o[14] ;
  output \mc_addr_pad_o[15] ;
  output \mc_addr_pad_o[16] ;
  output \mc_addr_pad_o[17] ;
  output \mc_addr_pad_o[18] ;
  output \mc_addr_pad_o[19] ;
  output \mc_addr_pad_o[1] ;
  output \mc_addr_pad_o[20] ;
  output \mc_addr_pad_o[21] ;
  output \mc_addr_pad_o[22] ;
  output \mc_addr_pad_o[23] ;
  output \mc_addr_pad_o[2] ;
  output \mc_addr_pad_o[3] ;
  output \mc_addr_pad_o[4] ;
  output \mc_addr_pad_o[5] ;
  output \mc_addr_pad_o[6] ;
  output \mc_addr_pad_o[7] ;
  output \mc_addr_pad_o[8] ;
  output \mc_addr_pad_o[9] ;
  wire mc_adsc_d;
  output mc_adsc_pad_o_;
  wire mc_adv_d;
  output mc_adv_pad_o_;
  wire mc_bg_d;
  output mc_bg_pad_o;
  input mc_br_pad_i;
  wire mc_br_r;
  wire mc_c_oe_d;
  output mc_cas_pad_o_;
  output mc_cke_pad_o_;
  input mc_clk_i;
  wire mc_clk_i_bF_buf0;
  wire mc_clk_i_bF_buf1;
  wire mc_clk_i_bF_buf10;
  wire mc_clk_i_bF_buf2;
  wire mc_clk_i_bF_buf3;
  wire mc_clk_i_bF_buf4;
  wire mc_clk_i_bF_buf5;
  wire mc_clk_i_bF_buf6;
  wire mc_clk_i_bF_buf7;
  wire mc_clk_i_bF_buf8;
  wire mc_clk_i_bF_buf9;
  output mc_coe_pad_coe_o;
  output \mc_cs_pad_o_[0] ;
  output \mc_cs_pad_o_[1] ;
  output \mc_cs_pad_o_[2] ;
  output \mc_cs_pad_o_[3] ;
  output \mc_cs_pad_o_[4] ;
  output \mc_cs_pad_o_[5] ;
  output \mc_cs_pad_o_[6] ;
  output \mc_cs_pad_o_[7] ;
  wire mc_data_ir_0_;
  wire mc_data_ir_10_;
  wire mc_data_ir_11_;
  wire mc_data_ir_12_;
  wire mc_data_ir_13_;
  wire mc_data_ir_14_;
  wire mc_data_ir_15_;
  wire mc_data_ir_16_;
  wire mc_data_ir_17_;
  wire mc_data_ir_18_;
  wire mc_data_ir_19_;
  wire mc_data_ir_1_;
  wire mc_data_ir_20_;
  wire mc_data_ir_21_;
  wire mc_data_ir_22_;
  wire mc_data_ir_23_;
  wire mc_data_ir_24_;
  wire mc_data_ir_25_;
  wire mc_data_ir_26_;
  wire mc_data_ir_27_;
  wire mc_data_ir_28_;
  wire mc_data_ir_29_;
  wire mc_data_ir_2_;
  wire mc_data_ir_30_;
  wire mc_data_ir_31_;
  wire mc_data_ir_32_;
  wire mc_data_ir_33_;
  wire mc_data_ir_34_;
  wire mc_data_ir_35_;
  wire mc_data_ir_3_;
  wire mc_data_ir_4_;
  wire mc_data_ir_5_;
  wire mc_data_ir_6_;
  wire mc_data_ir_7_;
  wire mc_data_ir_8_;
  wire mc_data_ir_9_;
  wire mc_data_od_0_;
  wire mc_data_od_10_;
  wire mc_data_od_11_;
  wire mc_data_od_12_;
  wire mc_data_od_13_;
  wire mc_data_od_14_;
  wire mc_data_od_15_;
  wire mc_data_od_16_;
  wire mc_data_od_17_;
  wire mc_data_od_18_;
  wire mc_data_od_19_;
  wire mc_data_od_1_;
  wire mc_data_od_20_;
  wire mc_data_od_21_;
  wire mc_data_od_22_;
  wire mc_data_od_23_;
  wire mc_data_od_24_;
  wire mc_data_od_25_;
  wire mc_data_od_26_;
  wire mc_data_od_27_;
  wire mc_data_od_28_;
  wire mc_data_od_29_;
  wire mc_data_od_2_;
  wire mc_data_od_30_;
  wire mc_data_od_31_;
  wire mc_data_od_3_;
  wire mc_data_od_4_;
  wire mc_data_od_5_;
  wire mc_data_od_6_;
  wire mc_data_od_7_;
  wire mc_data_od_8_;
  wire mc_data_od_9_;
  input \mc_data_pad_i[0] ;
  input \mc_data_pad_i[10] ;
  input \mc_data_pad_i[11] ;
  input \mc_data_pad_i[12] ;
  input \mc_data_pad_i[13] ;
  input \mc_data_pad_i[14] ;
  input \mc_data_pad_i[15] ;
  input \mc_data_pad_i[16] ;
  input \mc_data_pad_i[17] ;
  input \mc_data_pad_i[18] ;
  input \mc_data_pad_i[19] ;
  input \mc_data_pad_i[1] ;
  input \mc_data_pad_i[20] ;
  input \mc_data_pad_i[21] ;
  input \mc_data_pad_i[22] ;
  input \mc_data_pad_i[23] ;
  input \mc_data_pad_i[24] ;
  input \mc_data_pad_i[25] ;
  input \mc_data_pad_i[26] ;
  input \mc_data_pad_i[27] ;
  input \mc_data_pad_i[28] ;
  input \mc_data_pad_i[29] ;
  input \mc_data_pad_i[2] ;
  input \mc_data_pad_i[30] ;
  input \mc_data_pad_i[31] ;
  input \mc_data_pad_i[3] ;
  input \mc_data_pad_i[4] ;
  input \mc_data_pad_i[5] ;
  input \mc_data_pad_i[6] ;
  input \mc_data_pad_i[7] ;
  input \mc_data_pad_i[8] ;
  input \mc_data_pad_i[9] ;
  output \mc_data_pad_o[0] ;
  output \mc_data_pad_o[10] ;
  output \mc_data_pad_o[11] ;
  output \mc_data_pad_o[12] ;
  output \mc_data_pad_o[13] ;
  output \mc_data_pad_o[14] ;
  output \mc_data_pad_o[15] ;
  output \mc_data_pad_o[16] ;
  output \mc_data_pad_o[17] ;
  output \mc_data_pad_o[18] ;
  output \mc_data_pad_o[19] ;
  output \mc_data_pad_o[1] ;
  output \mc_data_pad_o[20] ;
  output \mc_data_pad_o[21] ;
  output \mc_data_pad_o[22] ;
  output \mc_data_pad_o[23] ;
  output \mc_data_pad_o[24] ;
  output \mc_data_pad_o[25] ;
  output \mc_data_pad_o[26] ;
  output \mc_data_pad_o[27] ;
  output \mc_data_pad_o[28] ;
  output \mc_data_pad_o[29] ;
  output \mc_data_pad_o[2] ;
  output \mc_data_pad_o[30] ;
  output \mc_data_pad_o[31] ;
  output \mc_data_pad_o[3] ;
  output \mc_data_pad_o[4] ;
  output \mc_data_pad_o[5] ;
  output \mc_data_pad_o[6] ;
  output \mc_data_pad_o[7] ;
  output \mc_data_pad_o[8] ;
  output \mc_data_pad_o[9] ;
  output mc_doe_pad_doe_o;
  wire mc_dp_od_0_;
  wire mc_dp_od_1_;
  wire mc_dp_od_2_;
  wire mc_dp_od_3_;
  input \mc_dp_pad_i[0] ;
  input \mc_dp_pad_i[1] ;
  input \mc_dp_pad_i[2] ;
  input \mc_dp_pad_i[3] ;
  output \mc_dp_pad_o[0] ;
  output \mc_dp_pad_o[1] ;
  output \mc_dp_pad_o[2] ;
  output \mc_dp_pad_o[3] ;
  output \mc_dqm_pad_o[0] ;
  output \mc_dqm_pad_o[1] ;
  output \mc_dqm_pad_o[2] ;
  output \mc_dqm_pad_o[3] ;
  output mc_oe_pad_o_;
  output mc_ras_pad_o_;
  output mc_rp_pad_o_;
  wire mc_sts_ir;
  input mc_sts_pad_i;
  output mc_vpen_pad_o;
  output mc_we_pad_o_;
  output mc_zz_pad_o;
  wire mem_ack;
  wire mem_ack_r;
  wire mem_dout_0_;
  wire mem_dout_10_;
  wire mem_dout_11_;
  wire mem_dout_12_;
  wire mem_dout_13_;
  wire mem_dout_14_;
  wire mem_dout_15_;
  wire mem_dout_16_;
  wire mem_dout_17_;
  wire mem_dout_18_;
  wire mem_dout_19_;
  wire mem_dout_1_;
  wire mem_dout_20_;
  wire mem_dout_21_;
  wire mem_dout_22_;
  wire mem_dout_23_;
  wire mem_dout_24_;
  wire mem_dout_25_;
  wire mem_dout_26_;
  wire mem_dout_27_;
  wire mem_dout_28_;
  wire mem_dout_29_;
  wire mem_dout_2_;
  wire mem_dout_30_;
  wire mem_dout_31_;
  wire mem_dout_3_;
  wire mem_dout_4_;
  wire mem_dout_5_;
  wire mem_dout_6_;
  wire mem_dout_7_;
  wire mem_dout_8_;
  wire mem_dout_9_;
  wire next_adr;
  wire next_adr_bF_buf0;
  wire next_adr_bF_buf1;
  wire next_adr_bF_buf2;
  wire next_adr_bF_buf3;
  wire next_adr_bF_buf4;
  wire not_mem_cyc;
  wire obct_cs_0_;
  wire obct_cs_1_;
  wire obct_cs_2_;
  wire obct_cs_3_;
  wire obct_cs_4_;
  wire obct_cs_5_;
  wire obct_cs_6_;
  wire obct_cs_7_;
  wire oe_;
  wire pack_le0;
  wire pack_le1;
  wire pack_le2;
  wire page_size_10_;
  wire page_size_10_bF_buf0;
  wire page_size_10_bF_buf1;
  wire page_size_10_bF_buf2;
  wire page_size_10_bF_buf3;
  wire page_size_8_;
  wire page_size_9_;
  wire par_err;
  output \poc_o[0] ;
  output \poc_o[10] ;
  output \poc_o[11] ;
  output \poc_o[12] ;
  output \poc_o[13] ;
  output \poc_o[14] ;
  output \poc_o[15] ;
  output \poc_o[16] ;
  output \poc_o[17] ;
  output \poc_o[18] ;
  output \poc_o[19] ;
  output \poc_o[1] ;
  output \poc_o[20] ;
  output \poc_o[21] ;
  output \poc_o[22] ;
  output \poc_o[23] ;
  output \poc_o[24] ;
  output \poc_o[25] ;
  output \poc_o[26] ;
  output \poc_o[27] ;
  output \poc_o[28] ;
  output \poc_o[29] ;
  output \poc_o[2] ;
  output \poc_o[30] ;
  output \poc_o[31] ;
  output \poc_o[3] ;
  output \poc_o[4] ;
  output \poc_o[5] ;
  output \poc_o[6] ;
  output \poc_o[7] ;
  output \poc_o[8] ;
  output \poc_o[9] ;
  wire ras_;
  wire ref_int_0_;
  wire ref_int_1_;
  wire ref_int_2_;
  input resume_req_i;
  wire rf_dout_0_;
  wire rf_dout_10_;
  wire rf_dout_11_;
  wire rf_dout_12_;
  wire rf_dout_13_;
  wire rf_dout_14_;
  wire rf_dout_15_;
  wire rf_dout_16_;
  wire rf_dout_17_;
  wire rf_dout_18_;
  wire rf_dout_19_;
  wire rf_dout_1_;
  wire rf_dout_20_;
  wire rf_dout_21_;
  wire rf_dout_22_;
  wire rf_dout_23_;
  wire rf_dout_24_;
  wire rf_dout_25_;
  wire rf_dout_26_;
  wire rf_dout_27_;
  wire rf_dout_28_;
  wire rf_dout_29_;
  wire rf_dout_2_;
  wire rf_dout_30_;
  wire rf_dout_31_;
  wire rf_dout_3_;
  wire rf_dout_4_;
  wire rf_dout_5_;
  wire rf_dout_6_;
  wire rf_dout_7_;
  wire rf_dout_8_;
  wire rf_dout_9_;
  wire rfr_ack;
  wire rfr_ps_val_0_;
  wire rfr_ps_val_1_;
  wire rfr_ps_val_2_;
  wire rfr_ps_val_3_;
  wire rfr_ps_val_4_;
  wire rfr_ps_val_5_;
  wire rfr_ps_val_6_;
  wire rfr_ps_val_7_;
  wire rfr_req;
  wire row_adr_0_;
  wire row_adr_0_bF_buf0;
  wire row_adr_0_bF_buf1;
  wire row_adr_0_bF_buf2;
  wire row_adr_0_bF_buf3;
  wire row_adr_0_bF_buf4;
  wire row_adr_0_bF_buf5;
  wire row_adr_0_bF_buf6;
  wire row_adr_10_;
  wire row_adr_10_bF_buf0;
  wire row_adr_10_bF_buf1;
  wire row_adr_10_bF_buf2;
  wire row_adr_10_bF_buf3;
  wire row_adr_10_bF_buf4;
  wire row_adr_10_bF_buf5;
  wire row_adr_10_bF_buf6;
  wire row_adr_11_;
  wire row_adr_11_bF_buf0;
  wire row_adr_11_bF_buf1;
  wire row_adr_11_bF_buf2;
  wire row_adr_11_bF_buf3;
  wire row_adr_11_bF_buf4;
  wire row_adr_11_bF_buf5;
  wire row_adr_11_bF_buf6;
  wire row_adr_12_;
  wire row_adr_12_bF_buf0;
  wire row_adr_12_bF_buf1;
  wire row_adr_12_bF_buf2;
  wire row_adr_12_bF_buf3;
  wire row_adr_12_bF_buf4;
  wire row_adr_12_bF_buf5;
  wire row_adr_12_bF_buf6;
  wire row_adr_1_;
  wire row_adr_1_bF_buf0;
  wire row_adr_1_bF_buf1;
  wire row_adr_1_bF_buf2;
  wire row_adr_1_bF_buf3;
  wire row_adr_1_bF_buf4;
  wire row_adr_1_bF_buf5;
  wire row_adr_1_bF_buf6;
  wire row_adr_2_;
  wire row_adr_2_bF_buf0;
  wire row_adr_2_bF_buf1;
  wire row_adr_2_bF_buf2;
  wire row_adr_2_bF_buf3;
  wire row_adr_2_bF_buf4;
  wire row_adr_2_bF_buf5;
  wire row_adr_2_bF_buf6;
  wire row_adr_3_;
  wire row_adr_3_bF_buf0;
  wire row_adr_3_bF_buf1;
  wire row_adr_3_bF_buf2;
  wire row_adr_3_bF_buf3;
  wire row_adr_3_bF_buf4;
  wire row_adr_3_bF_buf5;
  wire row_adr_3_bF_buf6;
  wire row_adr_4_;
  wire row_adr_4_bF_buf0;
  wire row_adr_4_bF_buf1;
  wire row_adr_4_bF_buf2;
  wire row_adr_4_bF_buf3;
  wire row_adr_4_bF_buf4;
  wire row_adr_4_bF_buf5;
  wire row_adr_4_bF_buf6;
  wire row_adr_5_;
  wire row_adr_5_bF_buf0;
  wire row_adr_5_bF_buf1;
  wire row_adr_5_bF_buf2;
  wire row_adr_5_bF_buf3;
  wire row_adr_5_bF_buf4;
  wire row_adr_5_bF_buf5;
  wire row_adr_5_bF_buf6;
  wire row_adr_6_;
  wire row_adr_6_bF_buf0;
  wire row_adr_6_bF_buf1;
  wire row_adr_6_bF_buf2;
  wire row_adr_6_bF_buf3;
  wire row_adr_6_bF_buf4;
  wire row_adr_6_bF_buf5;
  wire row_adr_6_bF_buf6;
  wire row_adr_7_;
  wire row_adr_7_bF_buf0;
  wire row_adr_7_bF_buf1;
  wire row_adr_7_bF_buf2;
  wire row_adr_7_bF_buf3;
  wire row_adr_7_bF_buf4;
  wire row_adr_7_bF_buf5;
  wire row_adr_7_bF_buf6;
  wire row_adr_8_;
  wire row_adr_8_bF_buf0;
  wire row_adr_8_bF_buf1;
  wire row_adr_8_bF_buf2;
  wire row_adr_8_bF_buf3;
  wire row_adr_8_bF_buf4;
  wire row_adr_8_bF_buf5;
  wire row_adr_8_bF_buf6;
  wire row_adr_9_;
  wire row_adr_9_bF_buf0;
  wire row_adr_9_bF_buf1;
  wire row_adr_9_bF_buf2;
  wire row_adr_9_bF_buf3;
  wire row_adr_9_bF_buf4;
  wire row_adr_9_bF_buf5;
  wire row_adr_9_bF_buf6;
  wire row_same;
  wire row_sel;
  input rst_i;
  wire rst_i_bF_buf0;
  wire rst_i_bF_buf1;
  wire rst_i_bF_buf2;
  wire rst_i_bF_buf3;
  wire sp_csc_10_;
  wire sp_csc_1_;
  wire sp_csc_2_;
  wire sp_csc_3_;
  wire sp_csc_4_;
  wire sp_csc_5_;
  wire sp_csc_6_;
  wire sp_csc_7_;
  wire sp_csc_9_;
  wire sp_tms_0_;
  wire sp_tms_10_;
  wire sp_tms_11_;
  wire sp_tms_12_;
  wire sp_tms_13_;
  wire sp_tms_14_;
  wire sp_tms_15_;
  wire sp_tms_16_;
  wire sp_tms_17_;
  wire sp_tms_18_;
  wire sp_tms_19_;
  wire sp_tms_1_;
  wire sp_tms_20_;
  wire sp_tms_21_;
  wire sp_tms_22_;
  wire sp_tms_23_;
  wire sp_tms_24_;
  wire sp_tms_25_;
  wire sp_tms_26_;
  wire sp_tms_27_;
  wire sp_tms_2_;
  wire sp_tms_3_;
  wire sp_tms_4_;
  wire sp_tms_5_;
  wire sp_tms_6_;
  wire sp_tms_7_;
  wire sp_tms_8_;
  wire sp_tms_9_;
  wire spec_req_cs_0_;
  wire spec_req_cs_0_bF_buf0;
  wire spec_req_cs_0_bF_buf1;
  wire spec_req_cs_0_bF_buf2;
  wire spec_req_cs_0_bF_buf3;
  wire spec_req_cs_0_bF_buf4;
  wire spec_req_cs_0_bF_buf5;
  wire spec_req_cs_1_;
  wire spec_req_cs_1_bF_buf0;
  wire spec_req_cs_1_bF_buf1;
  wire spec_req_cs_1_bF_buf2;
  wire spec_req_cs_1_bF_buf3;
  wire spec_req_cs_1_bF_buf4;
  wire spec_req_cs_1_bF_buf5;
  wire spec_req_cs_2_;
  wire spec_req_cs_2_bF_buf0;
  wire spec_req_cs_2_bF_buf1;
  wire spec_req_cs_2_bF_buf2;
  wire spec_req_cs_2_bF_buf3;
  wire spec_req_cs_2_bF_buf4;
  wire spec_req_cs_2_bF_buf5;
  wire spec_req_cs_3_;
  wire spec_req_cs_3_bF_buf0;
  wire spec_req_cs_3_bF_buf1;
  wire spec_req_cs_3_bF_buf2;
  wire spec_req_cs_3_bF_buf3;
  wire spec_req_cs_3_bF_buf4;
  wire spec_req_cs_3_bF_buf5;
  wire spec_req_cs_4_;
  wire spec_req_cs_4_bF_buf0;
  wire spec_req_cs_4_bF_buf1;
  wire spec_req_cs_4_bF_buf2;
  wire spec_req_cs_4_bF_buf3;
  wire spec_req_cs_4_bF_buf4;
  wire spec_req_cs_4_bF_buf5;
  wire spec_req_cs_5_;
  wire spec_req_cs_5_bF_buf0;
  wire spec_req_cs_5_bF_buf1;
  wire spec_req_cs_5_bF_buf2;
  wire spec_req_cs_5_bF_buf3;
  wire spec_req_cs_5_bF_buf4;
  wire spec_req_cs_5_bF_buf5;
  wire spec_req_cs_6_;
  wire spec_req_cs_6_bF_buf0;
  wire spec_req_cs_6_bF_buf1;
  wire spec_req_cs_6_bF_buf2;
  wire spec_req_cs_6_bF_buf3;
  wire spec_req_cs_6_bF_buf4;
  wire spec_req_cs_6_bF_buf5;
  wire spec_req_cs_7_;
  input susp_req_i;
  wire susp_sel;
  output suspended_o;
  wire tms_0_;
  wire tms_10_;
  wire tms_11_;
  wire tms_12_;
  wire tms_13_;
  wire tms_14_;
  wire tms_15_;
  wire tms_16_;
  wire tms_17_;
  wire tms_18_;
  wire tms_19_;
  wire tms_1_;
  wire tms_20_;
  wire tms_21_;
  wire tms_22_;
  wire tms_23_;
  wire tms_24_;
  wire tms_25_;
  wire tms_26_;
  wire tms_27_;
  wire tms_2_;
  wire tms_3_;
  wire tms_4_;
  wire tms_5_;
  wire tms_6_;
  wire tms_7_;
  wire tms_8_;
  wire tms_9_;
  wire tms_s_0_;
  wire tms_s_10_;
  wire tms_s_11_;
  wire tms_s_12_;
  wire tms_s_13_;
  wire tms_s_14_;
  wire tms_s_15_;
  wire tms_s_16_;
  wire tms_s_17_;
  wire tms_s_18_;
  wire tms_s_19_;
  wire tms_s_1_;
  wire tms_s_20_;
  wire tms_s_21_;
  wire tms_s_22_;
  wire tms_s_23_;
  wire tms_s_24_;
  wire tms_s_25_;
  wire tms_s_26_;
  wire tms_s_27_;
  wire tms_s_2_;
  wire tms_s_3_;
  wire tms_s_4_;
  wire tms_s_5_;
  wire tms_s_6_;
  wire tms_s_7_;
  wire tms_s_8_;
  wire tms_s_9_;
  wire u0__abc_49347_n1100_1;
  wire u0__abc_49347_n1101_1;
  wire u0__abc_49347_n1102;
  wire u0__abc_49347_n1103_1;
  wire u0__abc_49347_n1104;
  wire u0__abc_49347_n1105_1;
  wire u0__abc_49347_n1106;
  wire u0__abc_49347_n1107_1;
  wire u0__abc_49347_n1109_1;
  wire u0__abc_49347_n1110;
  wire u0__abc_49347_n1111_1;
  wire u0__abc_49347_n1112;
  wire u0__abc_49347_n1113_1;
  wire u0__abc_49347_n1114;
  wire u0__abc_49347_n1116_1;
  wire u0__abc_49347_n1117_1;
  wire u0__abc_49347_n1118_1;
  wire u0__abc_49347_n1119;
  wire u0__abc_49347_n1120_1;
  wire u0__abc_49347_n1121;
  wire u0__abc_49347_n1122_1;
  wire u0__abc_49347_n1124_1;
  wire u0__abc_49347_n1125;
  wire u0__abc_49347_n1126_1;
  wire u0__abc_49347_n1127;
  wire u0__abc_49347_n1128_1;
  wire u0__abc_49347_n1129;
  wire u0__abc_49347_n1130_1;
  wire u0__abc_49347_n1131;
  wire u0__abc_49347_n1133_1;
  wire u0__abc_49347_n1134_1;
  wire u0__abc_49347_n1135_1;
  wire u0__abc_49347_n1136;
  wire u0__abc_49347_n1137_1;
  wire u0__abc_49347_n1138;
  wire u0__abc_49347_n1139_1;
  wire u0__abc_49347_n1140;
  wire u0__abc_49347_n1141_1;
  wire u0__abc_49347_n1143_1;
  wire u0__abc_49347_n1144;
  wire u0__abc_49347_n1145_1;
  wire u0__abc_49347_n1146;
  wire u0__abc_49347_n1147_1;
  wire u0__abc_49347_n1148;
  wire u0__abc_49347_n1149_1;
  wire u0__abc_49347_n1150_1;
  wire u0__abc_49347_n1151_1;
  wire u0__abc_49347_n1153;
  wire u0__abc_49347_n1154_1;
  wire u0__abc_49347_n1155;
  wire u0__abc_49347_n1156_1;
  wire u0__abc_49347_n1157;
  wire u0__abc_49347_n1158_1;
  wire u0__abc_49347_n1159;
  wire u0__abc_49347_n1160_1;
  wire u0__abc_49347_n1161;
  wire u0__abc_49347_n1163;
  wire u0__abc_49347_n1164_1;
  wire u0__abc_49347_n1165;
  wire u0__abc_49347_n1166_1;
  wire u0__abc_49347_n1167_1;
  wire u0__abc_49347_n1168_1;
  wire u0__abc_49347_n1169;
  wire u0__abc_49347_n1170_1;
  wire u0__abc_49347_n1171;
  wire u0__abc_49347_n1173;
  wire u0__abc_49347_n1174_1;
  wire u0__abc_49347_n1175;
  wire u0__abc_49347_n1175_bF_buf0;
  wire u0__abc_49347_n1175_bF_buf1;
  wire u0__abc_49347_n1175_bF_buf2;
  wire u0__abc_49347_n1175_bF_buf3;
  wire u0__abc_49347_n1175_bF_buf4;
  wire u0__abc_49347_n1175_bF_buf5;
  wire u0__abc_49347_n1175_bF_buf6;
  wire u0__abc_49347_n1176_1;
  wire u0__abc_49347_n1176_1_bF_buf0;
  wire u0__abc_49347_n1176_1_bF_buf1;
  wire u0__abc_49347_n1176_1_bF_buf2;
  wire u0__abc_49347_n1176_1_bF_buf3;
  wire u0__abc_49347_n1176_1_bF_buf4;
  wire u0__abc_49347_n1176_1_bF_buf5;
  wire u0__abc_49347_n1176_1_bF_buf6;
  wire u0__abc_49347_n1177;
  wire u0__abc_49347_n1178_1;
  wire u0__abc_49347_n1178_1_bF_buf0;
  wire u0__abc_49347_n1178_1_bF_buf1;
  wire u0__abc_49347_n1178_1_bF_buf2;
  wire u0__abc_49347_n1178_1_bF_buf3;
  wire u0__abc_49347_n1178_1_bF_buf4;
  wire u0__abc_49347_n1178_1_bF_buf5;
  wire u0__abc_49347_n1179;
  wire u0__abc_49347_n1179_bF_buf0;
  wire u0__abc_49347_n1179_bF_buf1;
  wire u0__abc_49347_n1179_bF_buf2;
  wire u0__abc_49347_n1179_bF_buf3;
  wire u0__abc_49347_n1179_bF_buf4;
  wire u0__abc_49347_n1179_bF_buf5;
  wire u0__abc_49347_n1180_1;
  wire u0__abc_49347_n1180_1_bF_buf0;
  wire u0__abc_49347_n1180_1_bF_buf1;
  wire u0__abc_49347_n1180_1_bF_buf2;
  wire u0__abc_49347_n1180_1_bF_buf3;
  wire u0__abc_49347_n1180_1_bF_buf4;
  wire u0__abc_49347_n1180_1_bF_buf5;
  wire u0__abc_49347_n1181;
  wire u0__abc_49347_n1181_bF_buf0;
  wire u0__abc_49347_n1181_bF_buf1;
  wire u0__abc_49347_n1181_bF_buf2;
  wire u0__abc_49347_n1181_bF_buf3;
  wire u0__abc_49347_n1181_bF_buf4;
  wire u0__abc_49347_n1181_bF_buf5;
  wire u0__abc_49347_n1182_1;
  wire u0__abc_49347_n1183_1;
  wire u0__abc_49347_n1183_1_bF_buf0;
  wire u0__abc_49347_n1183_1_bF_buf1;
  wire u0__abc_49347_n1183_1_bF_buf2;
  wire u0__abc_49347_n1183_1_bF_buf3;
  wire u0__abc_49347_n1183_1_bF_buf4;
  wire u0__abc_49347_n1183_1_bF_buf5;
  wire u0__abc_49347_n1184;
  wire u0__abc_49347_n1185;
  wire u0__abc_49347_n1185_bF_buf0;
  wire u0__abc_49347_n1185_bF_buf1;
  wire u0__abc_49347_n1185_bF_buf2;
  wire u0__abc_49347_n1185_bF_buf3;
  wire u0__abc_49347_n1185_bF_buf4;
  wire u0__abc_49347_n1185_bF_buf5;
  wire u0__abc_49347_n1186;
  wire u0__abc_49347_n1187;
  wire u0__abc_49347_n1188;
  wire u0__abc_49347_n1189;
  wire u0__abc_49347_n1190;
  wire u0__abc_49347_n1191_1;
  wire u0__abc_49347_n1192_1;
  wire u0__abc_49347_n1193;
  wire u0__abc_49347_n1194;
  wire u0__abc_49347_n1195;
  wire u0__abc_49347_n1196;
  wire u0__abc_49347_n1197;
  wire u0__abc_49347_n1198;
  wire u0__abc_49347_n1199;
  wire u0__abc_49347_n1200_1;
  wire u0__abc_49347_n1201_1;
  wire u0__abc_49347_n1202;
  wire u0__abc_49347_n1203;
  wire u0__abc_49347_n1203_bF_buf0;
  wire u0__abc_49347_n1203_bF_buf1;
  wire u0__abc_49347_n1203_bF_buf2;
  wire u0__abc_49347_n1203_bF_buf3;
  wire u0__abc_49347_n1203_bF_buf4;
  wire u0__abc_49347_n1203_bF_buf5;
  wire u0__abc_49347_n1204;
  wire u0__abc_49347_n1205;
  wire u0__abc_49347_n1206;
  wire u0__abc_49347_n1208;
  wire u0__abc_49347_n1209_1;
  wire u0__abc_49347_n1210_1;
  wire u0__abc_49347_n1211;
  wire u0__abc_49347_n1212;
  wire u0__abc_49347_n1213;
  wire u0__abc_49347_n1214;
  wire u0__abc_49347_n1215;
  wire u0__abc_49347_n1216;
  wire u0__abc_49347_n1217;
  wire u0__abc_49347_n1218_1;
  wire u0__abc_49347_n1219_1;
  wire u0__abc_49347_n1220;
  wire u0__abc_49347_n1221;
  wire u0__abc_49347_n1222;
  wire u0__abc_49347_n1223;
  wire u0__abc_49347_n1224;
  wire u0__abc_49347_n1225;
  wire u0__abc_49347_n1226;
  wire u0__abc_49347_n1227_1;
  wire u0__abc_49347_n1228_1;
  wire u0__abc_49347_n1229;
  wire u0__abc_49347_n1230;
  wire u0__abc_49347_n1232;
  wire u0__abc_49347_n1233;
  wire u0__abc_49347_n1234;
  wire u0__abc_49347_n1235;
  wire u0__abc_49347_n1236_1;
  wire u0__abc_49347_n1237_1;
  wire u0__abc_49347_n1238;
  wire u0__abc_49347_n1239;
  wire u0__abc_49347_n1240;
  wire u0__abc_49347_n1241;
  wire u0__abc_49347_n1242;
  wire u0__abc_49347_n1243;
  wire u0__abc_49347_n1244;
  wire u0__abc_49347_n1245_1;
  wire u0__abc_49347_n1246_1;
  wire u0__abc_49347_n1247;
  wire u0__abc_49347_n1248;
  wire u0__abc_49347_n1249;
  wire u0__abc_49347_n1250;
  wire u0__abc_49347_n1251;
  wire u0__abc_49347_n1252;
  wire u0__abc_49347_n1253;
  wire u0__abc_49347_n1254_1;
  wire u0__abc_49347_n1256;
  wire u0__abc_49347_n1257;
  wire u0__abc_49347_n1258;
  wire u0__abc_49347_n1259;
  wire u0__abc_49347_n1260;
  wire u0__abc_49347_n1261;
  wire u0__abc_49347_n1262;
  wire u0__abc_49347_n1263_1;
  wire u0__abc_49347_n1264_1;
  wire u0__abc_49347_n1265;
  wire u0__abc_49347_n1266;
  wire u0__abc_49347_n1267;
  wire u0__abc_49347_n1268;
  wire u0__abc_49347_n1269;
  wire u0__abc_49347_n1270;
  wire u0__abc_49347_n1271;
  wire u0__abc_49347_n1272_1;
  wire u0__abc_49347_n1273_1;
  wire u0__abc_49347_n1274;
  wire u0__abc_49347_n1275;
  wire u0__abc_49347_n1276;
  wire u0__abc_49347_n1277;
  wire u0__abc_49347_n1278;
  wire u0__abc_49347_n1280;
  wire u0__abc_49347_n1281_1;
  wire u0__abc_49347_n1282_1;
  wire u0__abc_49347_n1283;
  wire u0__abc_49347_n1284;
  wire u0__abc_49347_n1285;
  wire u0__abc_49347_n1286;
  wire u0__abc_49347_n1287;
  wire u0__abc_49347_n1288;
  wire u0__abc_49347_n1289;
  wire u0__abc_49347_n1290_1;
  wire u0__abc_49347_n1291_1;
  wire u0__abc_49347_n1292;
  wire u0__abc_49347_n1293;
  wire u0__abc_49347_n1294;
  wire u0__abc_49347_n1295;
  wire u0__abc_49347_n1296;
  wire u0__abc_49347_n1297;
  wire u0__abc_49347_n1298;
  wire u0__abc_49347_n1299_1;
  wire u0__abc_49347_n1300_1;
  wire u0__abc_49347_n1301;
  wire u0__abc_49347_n1302;
  wire u0__abc_49347_n1304;
  wire u0__abc_49347_n1305;
  wire u0__abc_49347_n1306;
  wire u0__abc_49347_n1307;
  wire u0__abc_49347_n1308_1;
  wire u0__abc_49347_n1309_1;
  wire u0__abc_49347_n1310;
  wire u0__abc_49347_n1311;
  wire u0__abc_49347_n1312;
  wire u0__abc_49347_n1313;
  wire u0__abc_49347_n1314;
  wire u0__abc_49347_n1315;
  wire u0__abc_49347_n1316;
  wire u0__abc_49347_n1317_1;
  wire u0__abc_49347_n1318_1;
  wire u0__abc_49347_n1319;
  wire u0__abc_49347_n1320;
  wire u0__abc_49347_n1321;
  wire u0__abc_49347_n1322;
  wire u0__abc_49347_n1323;
  wire u0__abc_49347_n1324;
  wire u0__abc_49347_n1325;
  wire u0__abc_49347_n1326_1;
  wire u0__abc_49347_n1328;
  wire u0__abc_49347_n1329;
  wire u0__abc_49347_n1330;
  wire u0__abc_49347_n1331;
  wire u0__abc_49347_n1332;
  wire u0__abc_49347_n1333;
  wire u0__abc_49347_n1334;
  wire u0__abc_49347_n1335_1;
  wire u0__abc_49347_n1336_1;
  wire u0__abc_49347_n1337;
  wire u0__abc_49347_n1338;
  wire u0__abc_49347_n1339;
  wire u0__abc_49347_n1340;
  wire u0__abc_49347_n1341;
  wire u0__abc_49347_n1342;
  wire u0__abc_49347_n1343;
  wire u0__abc_49347_n1344_1;
  wire u0__abc_49347_n1345_1;
  wire u0__abc_49347_n1346;
  wire u0__abc_49347_n1347;
  wire u0__abc_49347_n1348;
  wire u0__abc_49347_n1349;
  wire u0__abc_49347_n1350;
  wire u0__abc_49347_n1352;
  wire u0__abc_49347_n1353_1;
  wire u0__abc_49347_n1354_1;
  wire u0__abc_49347_n1355;
  wire u0__abc_49347_n1356;
  wire u0__abc_49347_n1357;
  wire u0__abc_49347_n1358;
  wire u0__abc_49347_n1359;
  wire u0__abc_49347_n1360;
  wire u0__abc_49347_n1361;
  wire u0__abc_49347_n1362_1;
  wire u0__abc_49347_n1363_1;
  wire u0__abc_49347_n1364;
  wire u0__abc_49347_n1365;
  wire u0__abc_49347_n1366;
  wire u0__abc_49347_n1367;
  wire u0__abc_49347_n1368;
  wire u0__abc_49347_n1369;
  wire u0__abc_49347_n1370;
  wire u0__abc_49347_n1371_1;
  wire u0__abc_49347_n1372_1;
  wire u0__abc_49347_n1373;
  wire u0__abc_49347_n1374;
  wire u0__abc_49347_n1376;
  wire u0__abc_49347_n1377;
  wire u0__abc_49347_n1378;
  wire u0__abc_49347_n1379;
  wire u0__abc_49347_n1380_1;
  wire u0__abc_49347_n1381_1;
  wire u0__abc_49347_n1382;
  wire u0__abc_49347_n1383;
  wire u0__abc_49347_n1384;
  wire u0__abc_49347_n1385;
  wire u0__abc_49347_n1386;
  wire u0__abc_49347_n1387;
  wire u0__abc_49347_n1388;
  wire u0__abc_49347_n1389_1;
  wire u0__abc_49347_n1390_1;
  wire u0__abc_49347_n1391;
  wire u0__abc_49347_n1392;
  wire u0__abc_49347_n1393;
  wire u0__abc_49347_n1394;
  wire u0__abc_49347_n1395;
  wire u0__abc_49347_n1396;
  wire u0__abc_49347_n1397;
  wire u0__abc_49347_n1398_1;
  wire u0__abc_49347_n1400;
  wire u0__abc_49347_n1401;
  wire u0__abc_49347_n1402;
  wire u0__abc_49347_n1403;
  wire u0__abc_49347_n1404;
  wire u0__abc_49347_n1405;
  wire u0__abc_49347_n1406;
  wire u0__abc_49347_n1407_1;
  wire u0__abc_49347_n1408_1;
  wire u0__abc_49347_n1409;
  wire u0__abc_49347_n1410;
  wire u0__abc_49347_n1411;
  wire u0__abc_49347_n1412;
  wire u0__abc_49347_n1413;
  wire u0__abc_49347_n1414;
  wire u0__abc_49347_n1415;
  wire u0__abc_49347_n1416_1;
  wire u0__abc_49347_n1417_1;
  wire u0__abc_49347_n1418;
  wire u0__abc_49347_n1419;
  wire u0__abc_49347_n1420;
  wire u0__abc_49347_n1421;
  wire u0__abc_49347_n1422;
  wire u0__abc_49347_n1424;
  wire u0__abc_49347_n1425_1;
  wire u0__abc_49347_n1426_1;
  wire u0__abc_49347_n1427;
  wire u0__abc_49347_n1428;
  wire u0__abc_49347_n1429;
  wire u0__abc_49347_n1430;
  wire u0__abc_49347_n1431;
  wire u0__abc_49347_n1432;
  wire u0__abc_49347_n1433;
  wire u0__abc_49347_n1434_1;
  wire u0__abc_49347_n1435_1;
  wire u0__abc_49347_n1436;
  wire u0__abc_49347_n1437;
  wire u0__abc_49347_n1438;
  wire u0__abc_49347_n1439;
  wire u0__abc_49347_n1440;
  wire u0__abc_49347_n1441;
  wire u0__abc_49347_n1442;
  wire u0__abc_49347_n1443_1;
  wire u0__abc_49347_n1444_1;
  wire u0__abc_49347_n1445;
  wire u0__abc_49347_n1446;
  wire u0__abc_49347_n1448;
  wire u0__abc_49347_n1449;
  wire u0__abc_49347_n1450;
  wire u0__abc_49347_n1451;
  wire u0__abc_49347_n1452_1;
  wire u0__abc_49347_n1453_1;
  wire u0__abc_49347_n1454;
  wire u0__abc_49347_n1455;
  wire u0__abc_49347_n1456;
  wire u0__abc_49347_n1457;
  wire u0__abc_49347_n1458;
  wire u0__abc_49347_n1459;
  wire u0__abc_49347_n1460;
  wire u0__abc_49347_n1461_1;
  wire u0__abc_49347_n1462_1;
  wire u0__abc_49347_n1463;
  wire u0__abc_49347_n1464;
  wire u0__abc_49347_n1465;
  wire u0__abc_49347_n1466;
  wire u0__abc_49347_n1467;
  wire u0__abc_49347_n1468;
  wire u0__abc_49347_n1469;
  wire u0__abc_49347_n1470_1;
  wire u0__abc_49347_n1472;
  wire u0__abc_49347_n1473;
  wire u0__abc_49347_n1474;
  wire u0__abc_49347_n1475;
  wire u0__abc_49347_n1476;
  wire u0__abc_49347_n1477;
  wire u0__abc_49347_n1478;
  wire u0__abc_49347_n1479_1;
  wire u0__abc_49347_n1480_1;
  wire u0__abc_49347_n1481;
  wire u0__abc_49347_n1482;
  wire u0__abc_49347_n1483;
  wire u0__abc_49347_n1484;
  wire u0__abc_49347_n1485;
  wire u0__abc_49347_n1486;
  wire u0__abc_49347_n1487;
  wire u0__abc_49347_n1488_1;
  wire u0__abc_49347_n1489_1;
  wire u0__abc_49347_n1490;
  wire u0__abc_49347_n1491;
  wire u0__abc_49347_n1492;
  wire u0__abc_49347_n1493;
  wire u0__abc_49347_n1494;
  wire u0__abc_49347_n1496;
  wire u0__abc_49347_n1497_1;
  wire u0__abc_49347_n1498_1;
  wire u0__abc_49347_n1499;
  wire u0__abc_49347_n1500;
  wire u0__abc_49347_n1501;
  wire u0__abc_49347_n1502;
  wire u0__abc_49347_n1503;
  wire u0__abc_49347_n1504;
  wire u0__abc_49347_n1505;
  wire u0__abc_49347_n1506_1;
  wire u0__abc_49347_n1507_1;
  wire u0__abc_49347_n1508;
  wire u0__abc_49347_n1509;
  wire u0__abc_49347_n1510;
  wire u0__abc_49347_n1511;
  wire u0__abc_49347_n1512;
  wire u0__abc_49347_n1513;
  wire u0__abc_49347_n1514;
  wire u0__abc_49347_n1515_1;
  wire u0__abc_49347_n1516_1;
  wire u0__abc_49347_n1517;
  wire u0__abc_49347_n1518;
  wire u0__abc_49347_n1520;
  wire u0__abc_49347_n1521;
  wire u0__abc_49347_n1522;
  wire u0__abc_49347_n1523;
  wire u0__abc_49347_n1524_1;
  wire u0__abc_49347_n1525_1;
  wire u0__abc_49347_n1526;
  wire u0__abc_49347_n1527;
  wire u0__abc_49347_n1528;
  wire u0__abc_49347_n1529;
  wire u0__abc_49347_n1530;
  wire u0__abc_49347_n1531;
  wire u0__abc_49347_n1532;
  wire u0__abc_49347_n1533_1;
  wire u0__abc_49347_n1534_1;
  wire u0__abc_49347_n1535;
  wire u0__abc_49347_n1536;
  wire u0__abc_49347_n1537;
  wire u0__abc_49347_n1538;
  wire u0__abc_49347_n1539;
  wire u0__abc_49347_n1540;
  wire u0__abc_49347_n1541;
  wire u0__abc_49347_n1542_1;
  wire u0__abc_49347_n1544;
  wire u0__abc_49347_n1545;
  wire u0__abc_49347_n1546;
  wire u0__abc_49347_n1547;
  wire u0__abc_49347_n1548;
  wire u0__abc_49347_n1549;
  wire u0__abc_49347_n1550;
  wire u0__abc_49347_n1551_1;
  wire u0__abc_49347_n1552_1;
  wire u0__abc_49347_n1553;
  wire u0__abc_49347_n1554;
  wire u0__abc_49347_n1555;
  wire u0__abc_49347_n1556;
  wire u0__abc_49347_n1557;
  wire u0__abc_49347_n1558;
  wire u0__abc_49347_n1559;
  wire u0__abc_49347_n1560_1;
  wire u0__abc_49347_n1561_1;
  wire u0__abc_49347_n1562;
  wire u0__abc_49347_n1563;
  wire u0__abc_49347_n1564;
  wire u0__abc_49347_n1565;
  wire u0__abc_49347_n1566;
  wire u0__abc_49347_n1568;
  wire u0__abc_49347_n1569_1;
  wire u0__abc_49347_n1570_1;
  wire u0__abc_49347_n1571;
  wire u0__abc_49347_n1572;
  wire u0__abc_49347_n1573;
  wire u0__abc_49347_n1574;
  wire u0__abc_49347_n1575;
  wire u0__abc_49347_n1576;
  wire u0__abc_49347_n1577;
  wire u0__abc_49347_n1578_1;
  wire u0__abc_49347_n1579_1;
  wire u0__abc_49347_n1580;
  wire u0__abc_49347_n1581;
  wire u0__abc_49347_n1582;
  wire u0__abc_49347_n1583;
  wire u0__abc_49347_n1584;
  wire u0__abc_49347_n1585;
  wire u0__abc_49347_n1586;
  wire u0__abc_49347_n1587_1;
  wire u0__abc_49347_n1588_1;
  wire u0__abc_49347_n1589;
  wire u0__abc_49347_n1590;
  wire u0__abc_49347_n1592;
  wire u0__abc_49347_n1593;
  wire u0__abc_49347_n1594;
  wire u0__abc_49347_n1595;
  wire u0__abc_49347_n1596_1;
  wire u0__abc_49347_n1597_1;
  wire u0__abc_49347_n1598;
  wire u0__abc_49347_n1599;
  wire u0__abc_49347_n1600;
  wire u0__abc_49347_n1601;
  wire u0__abc_49347_n1602;
  wire u0__abc_49347_n1603;
  wire u0__abc_49347_n1604;
  wire u0__abc_49347_n1605_1;
  wire u0__abc_49347_n1606_1;
  wire u0__abc_49347_n1607;
  wire u0__abc_49347_n1608;
  wire u0__abc_49347_n1609;
  wire u0__abc_49347_n1610;
  wire u0__abc_49347_n1611;
  wire u0__abc_49347_n1612;
  wire u0__abc_49347_n1613;
  wire u0__abc_49347_n1614_1;
  wire u0__abc_49347_n1616;
  wire u0__abc_49347_n1617;
  wire u0__abc_49347_n1618;
  wire u0__abc_49347_n1619;
  wire u0__abc_49347_n1620;
  wire u0__abc_49347_n1621;
  wire u0__abc_49347_n1622;
  wire u0__abc_49347_n1623_1;
  wire u0__abc_49347_n1624_1;
  wire u0__abc_49347_n1625;
  wire u0__abc_49347_n1626;
  wire u0__abc_49347_n1627;
  wire u0__abc_49347_n1628;
  wire u0__abc_49347_n1629;
  wire u0__abc_49347_n1630;
  wire u0__abc_49347_n1631;
  wire u0__abc_49347_n1632_1;
  wire u0__abc_49347_n1633_1;
  wire u0__abc_49347_n1634;
  wire u0__abc_49347_n1635;
  wire u0__abc_49347_n1636;
  wire u0__abc_49347_n1637;
  wire u0__abc_49347_n1638;
  wire u0__abc_49347_n1640;
  wire u0__abc_49347_n1641_1;
  wire u0__abc_49347_n1642_1;
  wire u0__abc_49347_n1643;
  wire u0__abc_49347_n1644;
  wire u0__abc_49347_n1645;
  wire u0__abc_49347_n1646;
  wire u0__abc_49347_n1647;
  wire u0__abc_49347_n1648;
  wire u0__abc_49347_n1649;
  wire u0__abc_49347_n1650_1;
  wire u0__abc_49347_n1651_1;
  wire u0__abc_49347_n1652;
  wire u0__abc_49347_n1653;
  wire u0__abc_49347_n1654;
  wire u0__abc_49347_n1655;
  wire u0__abc_49347_n1656;
  wire u0__abc_49347_n1657;
  wire u0__abc_49347_n1658;
  wire u0__abc_49347_n1659_1;
  wire u0__abc_49347_n1660_1;
  wire u0__abc_49347_n1661;
  wire u0__abc_49347_n1662;
  wire u0__abc_49347_n1664;
  wire u0__abc_49347_n1665;
  wire u0__abc_49347_n1666;
  wire u0__abc_49347_n1667;
  wire u0__abc_49347_n1668_1;
  wire u0__abc_49347_n1669_1;
  wire u0__abc_49347_n1670;
  wire u0__abc_49347_n1671;
  wire u0__abc_49347_n1672;
  wire u0__abc_49347_n1673;
  wire u0__abc_49347_n1674;
  wire u0__abc_49347_n1675;
  wire u0__abc_49347_n1676;
  wire u0__abc_49347_n1677_1;
  wire u0__abc_49347_n1678_1;
  wire u0__abc_49347_n1679;
  wire u0__abc_49347_n1680;
  wire u0__abc_49347_n1681;
  wire u0__abc_49347_n1682;
  wire u0__abc_49347_n1683;
  wire u0__abc_49347_n1684;
  wire u0__abc_49347_n1685;
  wire u0__abc_49347_n1686_1;
  wire u0__abc_49347_n1688;
  wire u0__abc_49347_n1689;
  wire u0__abc_49347_n1690;
  wire u0__abc_49347_n1691;
  wire u0__abc_49347_n1692;
  wire u0__abc_49347_n1693;
  wire u0__abc_49347_n1694;
  wire u0__abc_49347_n1695_1;
  wire u0__abc_49347_n1696_1;
  wire u0__abc_49347_n1697;
  wire u0__abc_49347_n1698;
  wire u0__abc_49347_n1699;
  wire u0__abc_49347_n1700;
  wire u0__abc_49347_n1701;
  wire u0__abc_49347_n1702;
  wire u0__abc_49347_n1703;
  wire u0__abc_49347_n1704_1;
  wire u0__abc_49347_n1705_1;
  wire u0__abc_49347_n1706;
  wire u0__abc_49347_n1707;
  wire u0__abc_49347_n1708;
  wire u0__abc_49347_n1709;
  wire u0__abc_49347_n1710;
  wire u0__abc_49347_n1712;
  wire u0__abc_49347_n1713_1;
  wire u0__abc_49347_n1714_1;
  wire u0__abc_49347_n1715;
  wire u0__abc_49347_n1716;
  wire u0__abc_49347_n1717;
  wire u0__abc_49347_n1718;
  wire u0__abc_49347_n1719;
  wire u0__abc_49347_n1720;
  wire u0__abc_49347_n1721;
  wire u0__abc_49347_n1722_1;
  wire u0__abc_49347_n1723_1;
  wire u0__abc_49347_n1724;
  wire u0__abc_49347_n1725;
  wire u0__abc_49347_n1726;
  wire u0__abc_49347_n1727;
  wire u0__abc_49347_n1728;
  wire u0__abc_49347_n1729;
  wire u0__abc_49347_n1730;
  wire u0__abc_49347_n1731_1;
  wire u0__abc_49347_n1732_1;
  wire u0__abc_49347_n1733;
  wire u0__abc_49347_n1734;
  wire u0__abc_49347_n1736;
  wire u0__abc_49347_n1737;
  wire u0__abc_49347_n1738;
  wire u0__abc_49347_n1739;
  wire u0__abc_49347_n1740_1;
  wire u0__abc_49347_n1741_1;
  wire u0__abc_49347_n1742;
  wire u0__abc_49347_n1743;
  wire u0__abc_49347_n1744;
  wire u0__abc_49347_n1745;
  wire u0__abc_49347_n1746;
  wire u0__abc_49347_n1747;
  wire u0__abc_49347_n1748;
  wire u0__abc_49347_n1749_1;
  wire u0__abc_49347_n1750_1;
  wire u0__abc_49347_n1751_1;
  wire u0__abc_49347_n1752;
  wire u0__abc_49347_n1753;
  wire u0__abc_49347_n1754_1;
  wire u0__abc_49347_n1755;
  wire u0__abc_49347_n1756_1;
  wire u0__abc_49347_n1757_1;
  wire u0__abc_49347_n1758;
  wire u0__abc_49347_n1760_1;
  wire u0__abc_49347_n1761;
  wire u0__abc_49347_n1762;
  wire u0__abc_49347_n1763_1;
  wire u0__abc_49347_n1764_1;
  wire u0__abc_49347_n1765;
  wire u0__abc_49347_n1766_1;
  wire u0__abc_49347_n1767_1;
  wire u0__abc_49347_n1768;
  wire u0__abc_49347_n1769;
  wire u0__abc_49347_n1770;
  wire u0__abc_49347_n1771_1;
  wire u0__abc_49347_n1772_1;
  wire u0__abc_49347_n1773_1;
  wire u0__abc_49347_n1774_1;
  wire u0__abc_49347_n1775_1;
  wire u0__abc_49347_n1776_1;
  wire u0__abc_49347_n1777_1;
  wire u0__abc_49347_n1778_1;
  wire u0__abc_49347_n1779_1;
  wire u0__abc_49347_n1780_1;
  wire u0__abc_49347_n1781_1;
  wire u0__abc_49347_n1782_1;
  wire u0__abc_49347_n1784_1;
  wire u0__abc_49347_n1785_1;
  wire u0__abc_49347_n1786_1;
  wire u0__abc_49347_n1787_1;
  wire u0__abc_49347_n1788_1;
  wire u0__abc_49347_n1789_1;
  wire u0__abc_49347_n1790_1;
  wire u0__abc_49347_n1791_1;
  wire u0__abc_49347_n1792_1;
  wire u0__abc_49347_n1793_1;
  wire u0__abc_49347_n1794_1;
  wire u0__abc_49347_n1795_1;
  wire u0__abc_49347_n1796_1;
  wire u0__abc_49347_n1797_1;
  wire u0__abc_49347_n1798_1;
  wire u0__abc_49347_n1799_1;
  wire u0__abc_49347_n1800_1;
  wire u0__abc_49347_n1801_1;
  wire u0__abc_49347_n1802_1;
  wire u0__abc_49347_n1803_1;
  wire u0__abc_49347_n1804_1;
  wire u0__abc_49347_n1805_1;
  wire u0__abc_49347_n1806_1;
  wire u0__abc_49347_n1808_1;
  wire u0__abc_49347_n1809_1;
  wire u0__abc_49347_n1810_1;
  wire u0__abc_49347_n1811_1;
  wire u0__abc_49347_n1812_1;
  wire u0__abc_49347_n1813_1;
  wire u0__abc_49347_n1814_1;
  wire u0__abc_49347_n1815_1;
  wire u0__abc_49347_n1816_1;
  wire u0__abc_49347_n1817_1;
  wire u0__abc_49347_n1818_1;
  wire u0__abc_49347_n1819_1;
  wire u0__abc_49347_n1820_1;
  wire u0__abc_49347_n1821_1;
  wire u0__abc_49347_n1822_1;
  wire u0__abc_49347_n1823_1;
  wire u0__abc_49347_n1824_1;
  wire u0__abc_49347_n1825_1;
  wire u0__abc_49347_n1826_1;
  wire u0__abc_49347_n1827_1;
  wire u0__abc_49347_n1828_1;
  wire u0__abc_49347_n1829_1;
  wire u0__abc_49347_n1830_1;
  wire u0__abc_49347_n1832_1;
  wire u0__abc_49347_n1833_1;
  wire u0__abc_49347_n1834_1;
  wire u0__abc_49347_n1835_1;
  wire u0__abc_49347_n1836_1;
  wire u0__abc_49347_n1837_1;
  wire u0__abc_49347_n1838_1;
  wire u0__abc_49347_n1839_1;
  wire u0__abc_49347_n1840_1;
  wire u0__abc_49347_n1841_1;
  wire u0__abc_49347_n1842_1;
  wire u0__abc_49347_n1843_1;
  wire u0__abc_49347_n1844_1;
  wire u0__abc_49347_n1845_1;
  wire u0__abc_49347_n1846_1;
  wire u0__abc_49347_n1847_1;
  wire u0__abc_49347_n1848_1;
  wire u0__abc_49347_n1849_1;
  wire u0__abc_49347_n1850_1;
  wire u0__abc_49347_n1851_1;
  wire u0__abc_49347_n1852_1;
  wire u0__abc_49347_n1853_1;
  wire u0__abc_49347_n1854_1;
  wire u0__abc_49347_n1952_1;
  wire u0__abc_49347_n1952_1_bF_buf0;
  wire u0__abc_49347_n1952_1_bF_buf1;
  wire u0__abc_49347_n1952_1_bF_buf2;
  wire u0__abc_49347_n1952_1_bF_buf3;
  wire u0__abc_49347_n1953_1;
  wire u0__abc_49347_n1953_1_bF_buf0;
  wire u0__abc_49347_n1953_1_bF_buf1;
  wire u0__abc_49347_n1953_1_bF_buf2;
  wire u0__abc_49347_n1953_1_bF_buf3;
  wire u0__abc_49347_n1978;
  wire u0__abc_49347_n1979_1;
  wire u0__abc_49347_n1980;
  wire u0__abc_49347_n1981_1;
  wire u0__abc_49347_n1982;
  wire u0__abc_49347_n1983_1;
  wire u0__abc_49347_n1984_1;
  wire u0__abc_49347_n1985;
  wire u0__abc_49347_n1986;
  wire u0__abc_49347_n1987;
  wire u0__abc_49347_n1988;
  wire u0__abc_49347_n1989;
  wire u0__abc_49347_n1990;
  wire u0__abc_49347_n1991;
  wire u0__abc_49347_n1992;
  wire u0__abc_49347_n1993;
  wire u0__abc_49347_n1994;
  wire u0__abc_49347_n1995;
  wire u0__abc_49347_n1996;
  wire u0__abc_49347_n1997;
  wire u0__abc_49347_n1998;
  wire u0__abc_49347_n1999;
  wire u0__abc_49347_n2000;
  wire u0__abc_49347_n2002;
  wire u0__abc_49347_n2003;
  wire u0__abc_49347_n2004;
  wire u0__abc_49347_n2005;
  wire u0__abc_49347_n2006;
  wire u0__abc_49347_n2007;
  wire u0__abc_49347_n2008;
  wire u0__abc_49347_n2009;
  wire u0__abc_49347_n2010;
  wire u0__abc_49347_n2011;
  wire u0__abc_49347_n2012;
  wire u0__abc_49347_n2013;
  wire u0__abc_49347_n2014;
  wire u0__abc_49347_n2015;
  wire u0__abc_49347_n2016;
  wire u0__abc_49347_n2017;
  wire u0__abc_49347_n2018;
  wire u0__abc_49347_n2019;
  wire u0__abc_49347_n2020;
  wire u0__abc_49347_n2021;
  wire u0__abc_49347_n2022;
  wire u0__abc_49347_n2023;
  wire u0__abc_49347_n2024;
  wire u0__abc_49347_n2026;
  wire u0__abc_49347_n2027;
  wire u0__abc_49347_n2028;
  wire u0__abc_49347_n2029;
  wire u0__abc_49347_n2030;
  wire u0__abc_49347_n2031;
  wire u0__abc_49347_n2032;
  wire u0__abc_49347_n2033;
  wire u0__abc_49347_n2034;
  wire u0__abc_49347_n2035;
  wire u0__abc_49347_n2036;
  wire u0__abc_49347_n2037;
  wire u0__abc_49347_n2038;
  wire u0__abc_49347_n2039;
  wire u0__abc_49347_n2040;
  wire u0__abc_49347_n2041;
  wire u0__abc_49347_n2042;
  wire u0__abc_49347_n2043;
  wire u0__abc_49347_n2044;
  wire u0__abc_49347_n2045;
  wire u0__abc_49347_n2046;
  wire u0__abc_49347_n2047;
  wire u0__abc_49347_n2048;
  wire u0__abc_49347_n2050;
  wire u0__abc_49347_n2051_1;
  wire u0__abc_49347_n2052;
  wire u0__abc_49347_n2053;
  wire u0__abc_49347_n2054;
  wire u0__abc_49347_n2055;
  wire u0__abc_49347_n2056;
  wire u0__abc_49347_n2057;
  wire u0__abc_49347_n2058;
  wire u0__abc_49347_n2059;
  wire u0__abc_49347_n2060;
  wire u0__abc_49347_n2061;
  wire u0__abc_49347_n2062;
  wire u0__abc_49347_n2063;
  wire u0__abc_49347_n2064;
  wire u0__abc_49347_n2065;
  wire u0__abc_49347_n2066;
  wire u0__abc_49347_n2067;
  wire u0__abc_49347_n2068;
  wire u0__abc_49347_n2069;
  wire u0__abc_49347_n2070;
  wire u0__abc_49347_n2071;
  wire u0__abc_49347_n2072_1;
  wire u0__abc_49347_n2074;
  wire u0__abc_49347_n2075;
  wire u0__abc_49347_n2076;
  wire u0__abc_49347_n2077;
  wire u0__abc_49347_n2078;
  wire u0__abc_49347_n2079;
  wire u0__abc_49347_n2080;
  wire u0__abc_49347_n2081;
  wire u0__abc_49347_n2082;
  wire u0__abc_49347_n2083;
  wire u0__abc_49347_n2084;
  wire u0__abc_49347_n2085;
  wire u0__abc_49347_n2086;
  wire u0__abc_49347_n2087;
  wire u0__abc_49347_n2088;
  wire u0__abc_49347_n2089;
  wire u0__abc_49347_n2090;
  wire u0__abc_49347_n2091;
  wire u0__abc_49347_n2092;
  wire u0__abc_49347_n2093;
  wire u0__abc_49347_n2094;
  wire u0__abc_49347_n2095;
  wire u0__abc_49347_n2096;
  wire u0__abc_49347_n2098;
  wire u0__abc_49347_n2099;
  wire u0__abc_49347_n2100;
  wire u0__abc_49347_n2101;
  wire u0__abc_49347_n2102;
  wire u0__abc_49347_n2103;
  wire u0__abc_49347_n2104;
  wire u0__abc_49347_n2105;
  wire u0__abc_49347_n2106;
  wire u0__abc_49347_n2107;
  wire u0__abc_49347_n2108_1;
  wire u0__abc_49347_n2109;
  wire u0__abc_49347_n2110;
  wire u0__abc_49347_n2111;
  wire u0__abc_49347_n2112;
  wire u0__abc_49347_n2113;
  wire u0__abc_49347_n2114;
  wire u0__abc_49347_n2115;
  wire u0__abc_49347_n2116;
  wire u0__abc_49347_n2117;
  wire u0__abc_49347_n2118;
  wire u0__abc_49347_n2119;
  wire u0__abc_49347_n2120;
  wire u0__abc_49347_n2122;
  wire u0__abc_49347_n2123;
  wire u0__abc_49347_n2124;
  wire u0__abc_49347_n2125;
  wire u0__abc_49347_n2126;
  wire u0__abc_49347_n2127;
  wire u0__abc_49347_n2128;
  wire u0__abc_49347_n2129;
  wire u0__abc_49347_n2130;
  wire u0__abc_49347_n2131;
  wire u0__abc_49347_n2132;
  wire u0__abc_49347_n2133;
  wire u0__abc_49347_n2134;
  wire u0__abc_49347_n2135;
  wire u0__abc_49347_n2136;
  wire u0__abc_49347_n2137;
  wire u0__abc_49347_n2138;
  wire u0__abc_49347_n2139;
  wire u0__abc_49347_n2140;
  wire u0__abc_49347_n2141;
  wire u0__abc_49347_n2142;
  wire u0__abc_49347_n2143;
  wire u0__abc_49347_n2144_1;
  wire u0__abc_49347_n2170;
  wire u0__abc_49347_n2171;
  wire u0__abc_49347_n2172;
  wire u0__abc_49347_n2173;
  wire u0__abc_49347_n2174;
  wire u0__abc_49347_n2175;
  wire u0__abc_49347_n2176;
  wire u0__abc_49347_n2177;
  wire u0__abc_49347_n2178;
  wire u0__abc_49347_n2179;
  wire u0__abc_49347_n2180_1;
  wire u0__abc_49347_n2181;
  wire u0__abc_49347_n2182;
  wire u0__abc_49347_n2183;
  wire u0__abc_49347_n2184;
  wire u0__abc_49347_n2185;
  wire u0__abc_49347_n2186;
  wire u0__abc_49347_n2187;
  wire u0__abc_49347_n2188;
  wire u0__abc_49347_n2189;
  wire u0__abc_49347_n2190;
  wire u0__abc_49347_n2191;
  wire u0__abc_49347_n2192;
  wire u0__abc_49347_n2194;
  wire u0__abc_49347_n2195;
  wire u0__abc_49347_n2196;
  wire u0__abc_49347_n2197;
  wire u0__abc_49347_n2198;
  wire u0__abc_49347_n2199;
  wire u0__abc_49347_n2200;
  wire u0__abc_49347_n2201;
  wire u0__abc_49347_n2202;
  wire u0__abc_49347_n2203;
  wire u0__abc_49347_n2204;
  wire u0__abc_49347_n2205;
  wire u0__abc_49347_n2206;
  wire u0__abc_49347_n2207;
  wire u0__abc_49347_n2208;
  wire u0__abc_49347_n2209;
  wire u0__abc_49347_n2210;
  wire u0__abc_49347_n2211;
  wire u0__abc_49347_n2212;
  wire u0__abc_49347_n2213;
  wire u0__abc_49347_n2214;
  wire u0__abc_49347_n2215;
  wire u0__abc_49347_n2216_1;
  wire u0__abc_49347_n2722;
  wire u0__abc_49347_n2723;
  wire u0__abc_49347_n2723_bF_buf0;
  wire u0__abc_49347_n2723_bF_buf1;
  wire u0__abc_49347_n2723_bF_buf2;
  wire u0__abc_49347_n2723_bF_buf3;
  wire u0__abc_49347_n2723_bF_buf4;
  wire u0__abc_49347_n2723_bF_buf5;
  wire u0__abc_49347_n2724;
  wire u0__abc_49347_n2724_bF_buf0;
  wire u0__abc_49347_n2724_bF_buf1;
  wire u0__abc_49347_n2724_bF_buf2;
  wire u0__abc_49347_n2724_bF_buf3;
  wire u0__abc_49347_n2724_bF_buf4;
  wire u0__abc_49347_n2724_bF_buf5;
  wire u0__abc_49347_n2725;
  wire u0__abc_49347_n2725_bF_buf0;
  wire u0__abc_49347_n2725_bF_buf1;
  wire u0__abc_49347_n2725_bF_buf2;
  wire u0__abc_49347_n2725_bF_buf3;
  wire u0__abc_49347_n2725_bF_buf4;
  wire u0__abc_49347_n2725_bF_buf5;
  wire u0__abc_49347_n2726;
  wire u0__abc_49347_n2726_bF_buf0;
  wire u0__abc_49347_n2726_bF_buf1;
  wire u0__abc_49347_n2726_bF_buf2;
  wire u0__abc_49347_n2726_bF_buf3;
  wire u0__abc_49347_n2726_bF_buf4;
  wire u0__abc_49347_n2726_bF_buf5;
  wire u0__abc_49347_n2727;
  wire u0__abc_49347_n2728;
  wire u0__abc_49347_n2728_bF_buf0;
  wire u0__abc_49347_n2728_bF_buf1;
  wire u0__abc_49347_n2728_bF_buf2;
  wire u0__abc_49347_n2728_bF_buf3;
  wire u0__abc_49347_n2728_bF_buf4;
  wire u0__abc_49347_n2728_bF_buf5;
  wire u0__abc_49347_n2729;
  wire u0__abc_49347_n2730;
  wire u0__abc_49347_n2730_bF_buf0;
  wire u0__abc_49347_n2730_bF_buf1;
  wire u0__abc_49347_n2730_bF_buf2;
  wire u0__abc_49347_n2730_bF_buf3;
  wire u0__abc_49347_n2730_bF_buf4;
  wire u0__abc_49347_n2730_bF_buf5;
  wire u0__abc_49347_n2731;
  wire u0__abc_49347_n2732;
  wire u0__abc_49347_n2733;
  wire u0__abc_49347_n2734;
  wire u0__abc_49347_n2735;
  wire u0__abc_49347_n2736;
  wire u0__abc_49347_n2737;
  wire u0__abc_49347_n2738;
  wire u0__abc_49347_n2739;
  wire u0__abc_49347_n2740;
  wire u0__abc_49347_n2741;
  wire u0__abc_49347_n2742;
  wire u0__abc_49347_n2743;
  wire u0__abc_49347_n2744;
  wire u0__abc_49347_n2745;
  wire u0__abc_49347_n2746;
  wire u0__abc_49347_n2747;
  wire u0__abc_49347_n2748;
  wire u0__abc_49347_n2748_bF_buf0;
  wire u0__abc_49347_n2748_bF_buf1;
  wire u0__abc_49347_n2748_bF_buf2;
  wire u0__abc_49347_n2748_bF_buf3;
  wire u0__abc_49347_n2748_bF_buf4;
  wire u0__abc_49347_n2748_bF_buf5;
  wire u0__abc_49347_n2749;
  wire u0__abc_49347_n2750;
  wire u0__abc_49347_n2751;
  wire u0__abc_49347_n2753;
  wire u0__abc_49347_n2754;
  wire u0__abc_49347_n2755;
  wire u0__abc_49347_n2756;
  wire u0__abc_49347_n2757;
  wire u0__abc_49347_n2758;
  wire u0__abc_49347_n2759;
  wire u0__abc_49347_n2760;
  wire u0__abc_49347_n2761;
  wire u0__abc_49347_n2762;
  wire u0__abc_49347_n2763;
  wire u0__abc_49347_n2764;
  wire u0__abc_49347_n2765;
  wire u0__abc_49347_n2766;
  wire u0__abc_49347_n2767;
  wire u0__abc_49347_n2768;
  wire u0__abc_49347_n2769;
  wire u0__abc_49347_n2770;
  wire u0__abc_49347_n2771;
  wire u0__abc_49347_n2772;
  wire u0__abc_49347_n2773;
  wire u0__abc_49347_n2774;
  wire u0__abc_49347_n2775;
  wire u0__abc_49347_n2777;
  wire u0__abc_49347_n2778;
  wire u0__abc_49347_n2779;
  wire u0__abc_49347_n2780;
  wire u0__abc_49347_n2781;
  wire u0__abc_49347_n2782;
  wire u0__abc_49347_n2783;
  wire u0__abc_49347_n2784_1;
  wire u0__abc_49347_n2785;
  wire u0__abc_49347_n2786;
  wire u0__abc_49347_n2787;
  wire u0__abc_49347_n2788;
  wire u0__abc_49347_n2789;
  wire u0__abc_49347_n2790;
  wire u0__abc_49347_n2791;
  wire u0__abc_49347_n2792;
  wire u0__abc_49347_n2793;
  wire u0__abc_49347_n2794;
  wire u0__abc_49347_n2795;
  wire u0__abc_49347_n2796;
  wire u0__abc_49347_n2797;
  wire u0__abc_49347_n2798;
  wire u0__abc_49347_n2799;
  wire u0__abc_49347_n2801;
  wire u0__abc_49347_n2802;
  wire u0__abc_49347_n2803;
  wire u0__abc_49347_n2804;
  wire u0__abc_49347_n2805;
  wire u0__abc_49347_n2806;
  wire u0__abc_49347_n2807;
  wire u0__abc_49347_n2808;
  wire u0__abc_49347_n2809;
  wire u0__abc_49347_n2810;
  wire u0__abc_49347_n2811;
  wire u0__abc_49347_n2812;
  wire u0__abc_49347_n2813;
  wire u0__abc_49347_n2814;
  wire u0__abc_49347_n2815;
  wire u0__abc_49347_n2816_1;
  wire u0__abc_49347_n2817;
  wire u0__abc_49347_n2818;
  wire u0__abc_49347_n2819;
  wire u0__abc_49347_n2820;
  wire u0__abc_49347_n2821;
  wire u0__abc_49347_n2822;
  wire u0__abc_49347_n2823;
  wire u0__abc_49347_n2825;
  wire u0__abc_49347_n2826;
  wire u0__abc_49347_n2827;
  wire u0__abc_49347_n2828;
  wire u0__abc_49347_n2829;
  wire u0__abc_49347_n2830;
  wire u0__abc_49347_n2831;
  wire u0__abc_49347_n2832;
  wire u0__abc_49347_n2833;
  wire u0__abc_49347_n2834;
  wire u0__abc_49347_n2835;
  wire u0__abc_49347_n2836;
  wire u0__abc_49347_n2837;
  wire u0__abc_49347_n2838;
  wire u0__abc_49347_n2839;
  wire u0__abc_49347_n2840;
  wire u0__abc_49347_n2841;
  wire u0__abc_49347_n2842;
  wire u0__abc_49347_n2843;
  wire u0__abc_49347_n2844;
  wire u0__abc_49347_n2845;
  wire u0__abc_49347_n2846;
  wire u0__abc_49347_n2847;
  wire u0__abc_49347_n2849;
  wire u0__abc_49347_n2850;
  wire u0__abc_49347_n2851;
  wire u0__abc_49347_n2852;
  wire u0__abc_49347_n2853;
  wire u0__abc_49347_n2854;
  wire u0__abc_49347_n2855;
  wire u0__abc_49347_n2856;
  wire u0__abc_49347_n2857;
  wire u0__abc_49347_n2858;
  wire u0__abc_49347_n2859;
  wire u0__abc_49347_n2860;
  wire u0__abc_49347_n2861;
  wire u0__abc_49347_n2862;
  wire u0__abc_49347_n2863;
  wire u0__abc_49347_n2864;
  wire u0__abc_49347_n2865;
  wire u0__abc_49347_n2866;
  wire u0__abc_49347_n2867;
  wire u0__abc_49347_n2868;
  wire u0__abc_49347_n2869;
  wire u0__abc_49347_n2870;
  wire u0__abc_49347_n2871;
  wire u0__abc_49347_n2873;
  wire u0__abc_49347_n2874;
  wire u0__abc_49347_n2875;
  wire u0__abc_49347_n2876;
  wire u0__abc_49347_n2877;
  wire u0__abc_49347_n2878;
  wire u0__abc_49347_n2879;
  wire u0__abc_49347_n2880;
  wire u0__abc_49347_n2881_1;
  wire u0__abc_49347_n2882;
  wire u0__abc_49347_n2883;
  wire u0__abc_49347_n2884;
  wire u0__abc_49347_n2885;
  wire u0__abc_49347_n2886;
  wire u0__abc_49347_n2887;
  wire u0__abc_49347_n2888;
  wire u0__abc_49347_n2889;
  wire u0__abc_49347_n2890;
  wire u0__abc_49347_n2891;
  wire u0__abc_49347_n2892;
  wire u0__abc_49347_n2893;
  wire u0__abc_49347_n2894;
  wire u0__abc_49347_n2895;
  wire u0__abc_49347_n2897;
  wire u0__abc_49347_n2898;
  wire u0__abc_49347_n2899;
  wire u0__abc_49347_n2900;
  wire u0__abc_49347_n2901;
  wire u0__abc_49347_n2902;
  wire u0__abc_49347_n2903;
  wire u0__abc_49347_n2904;
  wire u0__abc_49347_n2905;
  wire u0__abc_49347_n2906;
  wire u0__abc_49347_n2907;
  wire u0__abc_49347_n2908;
  wire u0__abc_49347_n2909;
  wire u0__abc_49347_n2910;
  wire u0__abc_49347_n2911;
  wire u0__abc_49347_n2912;
  wire u0__abc_49347_n2913_1;
  wire u0__abc_49347_n2914;
  wire u0__abc_49347_n2915;
  wire u0__abc_49347_n2916;
  wire u0__abc_49347_n2917;
  wire u0__abc_49347_n2918;
  wire u0__abc_49347_n2919;
  wire u0__abc_49347_n2921;
  wire u0__abc_49347_n2922;
  wire u0__abc_49347_n2923;
  wire u0__abc_49347_n2924;
  wire u0__abc_49347_n2925;
  wire u0__abc_49347_n2926;
  wire u0__abc_49347_n2927;
  wire u0__abc_49347_n2928;
  wire u0__abc_49347_n2929;
  wire u0__abc_49347_n2930;
  wire u0__abc_49347_n2931;
  wire u0__abc_49347_n2932;
  wire u0__abc_49347_n2933;
  wire u0__abc_49347_n2934;
  wire u0__abc_49347_n2935;
  wire u0__abc_49347_n2936;
  wire u0__abc_49347_n2937;
  wire u0__abc_49347_n2938;
  wire u0__abc_49347_n2939;
  wire u0__abc_49347_n2940;
  wire u0__abc_49347_n2941;
  wire u0__abc_49347_n2942;
  wire u0__abc_49347_n2943;
  wire u0__abc_49347_n2945_1;
  wire u0__abc_49347_n2946;
  wire u0__abc_49347_n2947;
  wire u0__abc_49347_n2948;
  wire u0__abc_49347_n2949;
  wire u0__abc_49347_n2950;
  wire u0__abc_49347_n2951;
  wire u0__abc_49347_n2952;
  wire u0__abc_49347_n2953;
  wire u0__abc_49347_n2954;
  wire u0__abc_49347_n2955;
  wire u0__abc_49347_n2956;
  wire u0__abc_49347_n2957;
  wire u0__abc_49347_n2958;
  wire u0__abc_49347_n2959;
  wire u0__abc_49347_n2960;
  wire u0__abc_49347_n2961;
  wire u0__abc_49347_n2962;
  wire u0__abc_49347_n2963;
  wire u0__abc_49347_n2964;
  wire u0__abc_49347_n2965;
  wire u0__abc_49347_n2966;
  wire u0__abc_49347_n2967;
  wire u0__abc_49347_n2969;
  wire u0__abc_49347_n2970;
  wire u0__abc_49347_n2971;
  wire u0__abc_49347_n2972;
  wire u0__abc_49347_n2973;
  wire u0__abc_49347_n2974;
  wire u0__abc_49347_n2975;
  wire u0__abc_49347_n2976;
  wire u0__abc_49347_n2977_1;
  wire u0__abc_49347_n2978;
  wire u0__abc_49347_n2979;
  wire u0__abc_49347_n2980;
  wire u0__abc_49347_n2981;
  wire u0__abc_49347_n2982;
  wire u0__abc_49347_n2983;
  wire u0__abc_49347_n2984;
  wire u0__abc_49347_n2985;
  wire u0__abc_49347_n2986;
  wire u0__abc_49347_n2987;
  wire u0__abc_49347_n2988;
  wire u0__abc_49347_n2989;
  wire u0__abc_49347_n2990;
  wire u0__abc_49347_n2991;
  wire u0__abc_49347_n2993;
  wire u0__abc_49347_n2994;
  wire u0__abc_49347_n2995;
  wire u0__abc_49347_n2996;
  wire u0__abc_49347_n2997;
  wire u0__abc_49347_n2998;
  wire u0__abc_49347_n2999;
  wire u0__abc_49347_n3000;
  wire u0__abc_49347_n3001;
  wire u0__abc_49347_n3002;
  wire u0__abc_49347_n3003;
  wire u0__abc_49347_n3004;
  wire u0__abc_49347_n3005;
  wire u0__abc_49347_n3006;
  wire u0__abc_49347_n3007;
  wire u0__abc_49347_n3008;
  wire u0__abc_49347_n3009_1;
  wire u0__abc_49347_n3010;
  wire u0__abc_49347_n3011;
  wire u0__abc_49347_n3012;
  wire u0__abc_49347_n3013;
  wire u0__abc_49347_n3014;
  wire u0__abc_49347_n3015;
  wire u0__abc_49347_n3017;
  wire u0__abc_49347_n3018;
  wire u0__abc_49347_n3019;
  wire u0__abc_49347_n3020;
  wire u0__abc_49347_n3021;
  wire u0__abc_49347_n3022;
  wire u0__abc_49347_n3023;
  wire u0__abc_49347_n3024;
  wire u0__abc_49347_n3025;
  wire u0__abc_49347_n3026;
  wire u0__abc_49347_n3027;
  wire u0__abc_49347_n3028;
  wire u0__abc_49347_n3029;
  wire u0__abc_49347_n3030;
  wire u0__abc_49347_n3031;
  wire u0__abc_49347_n3032;
  wire u0__abc_49347_n3033;
  wire u0__abc_49347_n3034;
  wire u0__abc_49347_n3035;
  wire u0__abc_49347_n3036;
  wire u0__abc_49347_n3037;
  wire u0__abc_49347_n3038;
  wire u0__abc_49347_n3039;
  wire u0__abc_49347_n3041_1;
  wire u0__abc_49347_n3042;
  wire u0__abc_49347_n3043;
  wire u0__abc_49347_n3044;
  wire u0__abc_49347_n3045;
  wire u0__abc_49347_n3046;
  wire u0__abc_49347_n3047;
  wire u0__abc_49347_n3048;
  wire u0__abc_49347_n3049;
  wire u0__abc_49347_n3050;
  wire u0__abc_49347_n3051;
  wire u0__abc_49347_n3052;
  wire u0__abc_49347_n3053;
  wire u0__abc_49347_n3054;
  wire u0__abc_49347_n3055;
  wire u0__abc_49347_n3056;
  wire u0__abc_49347_n3057;
  wire u0__abc_49347_n3058;
  wire u0__abc_49347_n3059;
  wire u0__abc_49347_n3060;
  wire u0__abc_49347_n3061;
  wire u0__abc_49347_n3062;
  wire u0__abc_49347_n3063;
  wire u0__abc_49347_n3065;
  wire u0__abc_49347_n3066;
  wire u0__abc_49347_n3067;
  wire u0__abc_49347_n3068;
  wire u0__abc_49347_n3069;
  wire u0__abc_49347_n3070;
  wire u0__abc_49347_n3071;
  wire u0__abc_49347_n3072;
  wire u0__abc_49347_n3073_1;
  wire u0__abc_49347_n3074;
  wire u0__abc_49347_n3075;
  wire u0__abc_49347_n3076;
  wire u0__abc_49347_n3077;
  wire u0__abc_49347_n3078;
  wire u0__abc_49347_n3079;
  wire u0__abc_49347_n3080;
  wire u0__abc_49347_n3081;
  wire u0__abc_49347_n3082;
  wire u0__abc_49347_n3083;
  wire u0__abc_49347_n3084;
  wire u0__abc_49347_n3085;
  wire u0__abc_49347_n3086;
  wire u0__abc_49347_n3087;
  wire u0__abc_49347_n3089;
  wire u0__abc_49347_n3090;
  wire u0__abc_49347_n3091;
  wire u0__abc_49347_n3092;
  wire u0__abc_49347_n3093;
  wire u0__abc_49347_n3094;
  wire u0__abc_49347_n3095;
  wire u0__abc_49347_n3096;
  wire u0__abc_49347_n3097;
  wire u0__abc_49347_n3098;
  wire u0__abc_49347_n3099;
  wire u0__abc_49347_n3100;
  wire u0__abc_49347_n3101;
  wire u0__abc_49347_n3102;
  wire u0__abc_49347_n3103;
  wire u0__abc_49347_n3104;
  wire u0__abc_49347_n3105_1;
  wire u0__abc_49347_n3106_1;
  wire u0__abc_49347_n3107;
  wire u0__abc_49347_n3108_1;
  wire u0__abc_49347_n3109;
  wire u0__abc_49347_n3110_1;
  wire u0__abc_49347_n3111;
  wire u0__abc_49347_n3113;
  wire u0__abc_49347_n3114;
  wire u0__abc_49347_n3115_1;
  wire u0__abc_49347_n3116_1;
  wire u0__abc_49347_n3117;
  wire u0__abc_49347_n3118;
  wire u0__abc_49347_n3119;
  wire u0__abc_49347_n3120_1;
  wire u0__abc_49347_n3121;
  wire u0__abc_49347_n3122;
  wire u0__abc_49347_n3123_1;
  wire u0__abc_49347_n3124;
  wire u0__abc_49347_n3125;
  wire u0__abc_49347_n3126_1;
  wire u0__abc_49347_n3127;
  wire u0__abc_49347_n3128;
  wire u0__abc_49347_n3129_1;
  wire u0__abc_49347_n3130;
  wire u0__abc_49347_n3131;
  wire u0__abc_49347_n3132_1;
  wire u0__abc_49347_n3133;
  wire u0__abc_49347_n3134;
  wire u0__abc_49347_n3135_1;
  wire u0__abc_49347_n3137;
  wire u0__abc_49347_n3138_1;
  wire u0__abc_49347_n3139;
  wire u0__abc_49347_n3140;
  wire u0__abc_49347_n3141_1;
  wire u0__abc_49347_n3142;
  wire u0__abc_49347_n3143;
  wire u0__abc_49347_n3144_1;
  wire u0__abc_49347_n3145_1;
  wire u0__abc_49347_n3146;
  wire u0__abc_49347_n3147_1;
  wire u0__abc_49347_n3148;
  wire u0__abc_49347_n3149_1;
  wire u0__abc_49347_n3150;
  wire u0__abc_49347_n3151_1;
  wire u0__abc_49347_n3152;
  wire u0__abc_49347_n3153_1;
  wire u0__abc_49347_n3154;
  wire u0__abc_49347_n3155;
  wire u0__abc_49347_n3156_1;
  wire u0__abc_49347_n3157;
  wire u0__abc_49347_n3158;
  wire u0__abc_49347_n3159;
  wire u0__abc_49347_n3161;
  wire u0__abc_49347_n3162;
  wire u0__abc_49347_n3163_1;
  wire u0__abc_49347_n3164;
  wire u0__abc_49347_n3165;
  wire u0__abc_49347_n3166;
  wire u0__abc_49347_n3167;
  wire u0__abc_49347_n3168;
  wire u0__abc_49347_n3169;
  wire u0__abc_49347_n3170_1;
  wire u0__abc_49347_n3171_1;
  wire u0__abc_49347_n3172_1;
  wire u0__abc_49347_n3173_1;
  wire u0__abc_49347_n3174_1;
  wire u0__abc_49347_n3175_1;
  wire u0__abc_49347_n3176_1;
  wire u0__abc_49347_n3177_1;
  wire u0__abc_49347_n3178_1;
  wire u0__abc_49347_n3179_1;
  wire u0__abc_49347_n3180_1;
  wire u0__abc_49347_n3181_1;
  wire u0__abc_49347_n3182_1;
  wire u0__abc_49347_n3183_1;
  wire u0__abc_49347_n3185_1;
  wire u0__abc_49347_n3186_1;
  wire u0__abc_49347_n3187_1;
  wire u0__abc_49347_n3188;
  wire u0__abc_49347_n3188_1;
  wire u0__abc_49347_n3188_bF_buf0;
  wire u0__abc_49347_n3188_bF_buf1;
  wire u0__abc_49347_n3188_bF_buf10;
  wire u0__abc_49347_n3188_bF_buf2;
  wire u0__abc_49347_n3188_bF_buf3;
  wire u0__abc_49347_n3188_bF_buf4;
  wire u0__abc_49347_n3188_bF_buf5;
  wire u0__abc_49347_n3188_bF_buf6;
  wire u0__abc_49347_n3188_bF_buf7;
  wire u0__abc_49347_n3188_bF_buf8;
  wire u0__abc_49347_n3188_bF_buf9;
  wire u0__abc_49347_n3189;
  wire u0__abc_49347_n3190;
  wire u0__abc_49347_n3191;
  wire u0__abc_49347_n3192;
  wire u0__abc_49347_n3193;
  wire u0__abc_49347_n3194;
  wire u0__abc_49347_n3195;
  wire u0__abc_49347_n3196;
  wire u0__abc_49347_n3197;
  wire u0__abc_49347_n3198;
  wire u0__abc_49347_n3199;
  wire u0__abc_49347_n3200;
  wire u0__abc_49347_n3201;
  wire u0__abc_49347_n3202;
  wire u0__abc_49347_n3203;
  wire u0__abc_49347_n3204;
  wire u0__abc_49347_n3205;
  wire u0__abc_49347_n3206;
  wire u0__abc_49347_n3207;
  wire u0__abc_49347_n3209;
  wire u0__abc_49347_n3210;
  wire u0__abc_49347_n3211;
  wire u0__abc_49347_n3212;
  wire u0__abc_49347_n3213;
  wire u0__abc_49347_n3214;
  wire u0__abc_49347_n3215;
  wire u0__abc_49347_n3216;
  wire u0__abc_49347_n3217;
  wire u0__abc_49347_n3218;
  wire u0__abc_49347_n3219;
  wire u0__abc_49347_n3220;
  wire u0__abc_49347_n3221;
  wire u0__abc_49347_n3222;
  wire u0__abc_49347_n3223;
  wire u0__abc_49347_n3224;
  wire u0__abc_49347_n3225;
  wire u0__abc_49347_n3226;
  wire u0__abc_49347_n3227;
  wire u0__abc_49347_n3228;
  wire u0__abc_49347_n3229;
  wire u0__abc_49347_n3230;
  wire u0__abc_49347_n3231;
  wire u0__abc_49347_n3233;
  wire u0__abc_49347_n3234;
  wire u0__abc_49347_n3235;
  wire u0__abc_49347_n3236;
  wire u0__abc_49347_n3237;
  wire u0__abc_49347_n3238;
  wire u0__abc_49347_n3239;
  wire u0__abc_49347_n3240;
  wire u0__abc_49347_n3241;
  wire u0__abc_49347_n3242;
  wire u0__abc_49347_n3243;
  wire u0__abc_49347_n3244;
  wire u0__abc_49347_n3245;
  wire u0__abc_49347_n3246;
  wire u0__abc_49347_n3247;
  wire u0__abc_49347_n3248;
  wire u0__abc_49347_n3249;
  wire u0__abc_49347_n3250;
  wire u0__abc_49347_n3251;
  wire u0__abc_49347_n3252;
  wire u0__abc_49347_n3253;
  wire u0__abc_49347_n3254;
  wire u0__abc_49347_n3255;
  wire u0__abc_49347_n3257;
  wire u0__abc_49347_n3258;
  wire u0__abc_49347_n3259;
  wire u0__abc_49347_n3260;
  wire u0__abc_49347_n3261;
  wire u0__abc_49347_n3262;
  wire u0__abc_49347_n3263;
  wire u0__abc_49347_n3264;
  wire u0__abc_49347_n3265;
  wire u0__abc_49347_n3266;
  wire u0__abc_49347_n3267;
  wire u0__abc_49347_n3268;
  wire u0__abc_49347_n3269;
  wire u0__abc_49347_n3270;
  wire u0__abc_49347_n3271;
  wire u0__abc_49347_n3272;
  wire u0__abc_49347_n3273;
  wire u0__abc_49347_n3274;
  wire u0__abc_49347_n3275;
  wire u0__abc_49347_n3276;
  wire u0__abc_49347_n3277;
  wire u0__abc_49347_n3278;
  wire u0__abc_49347_n3279;
  wire u0__abc_49347_n3281;
  wire u0__abc_49347_n3282;
  wire u0__abc_49347_n3283;
  wire u0__abc_49347_n3284;
  wire u0__abc_49347_n3285;
  wire u0__abc_49347_n3286;
  wire u0__abc_49347_n3287;
  wire u0__abc_49347_n3288;
  wire u0__abc_49347_n3289;
  wire u0__abc_49347_n3290;
  wire u0__abc_49347_n3291;
  wire u0__abc_49347_n3292;
  wire u0__abc_49347_n3293;
  wire u0__abc_49347_n3294;
  wire u0__abc_49347_n3295;
  wire u0__abc_49347_n3296;
  wire u0__abc_49347_n3297;
  wire u0__abc_49347_n3298;
  wire u0__abc_49347_n3299;
  wire u0__abc_49347_n3300;
  wire u0__abc_49347_n3301;
  wire u0__abc_49347_n3302;
  wire u0__abc_49347_n3303;
  wire u0__abc_49347_n3305;
  wire u0__abc_49347_n3306;
  wire u0__abc_49347_n3307;
  wire u0__abc_49347_n3308;
  wire u0__abc_49347_n3309;
  wire u0__abc_49347_n3310;
  wire u0__abc_49347_n3311;
  wire u0__abc_49347_n3312;
  wire u0__abc_49347_n3313;
  wire u0__abc_49347_n3314;
  wire u0__abc_49347_n3315;
  wire u0__abc_49347_n3316;
  wire u0__abc_49347_n3317;
  wire u0__abc_49347_n3318;
  wire u0__abc_49347_n3319;
  wire u0__abc_49347_n3320;
  wire u0__abc_49347_n3321;
  wire u0__abc_49347_n3322;
  wire u0__abc_49347_n3323;
  wire u0__abc_49347_n3324;
  wire u0__abc_49347_n3325;
  wire u0__abc_49347_n3326;
  wire u0__abc_49347_n3327;
  wire u0__abc_49347_n3329;
  wire u0__abc_49347_n3330;
  wire u0__abc_49347_n3331;
  wire u0__abc_49347_n3332;
  wire u0__abc_49347_n3333;
  wire u0__abc_49347_n3334;
  wire u0__abc_49347_n3335;
  wire u0__abc_49347_n3336;
  wire u0__abc_49347_n3337;
  wire u0__abc_49347_n3338;
  wire u0__abc_49347_n3339;
  wire u0__abc_49347_n3340;
  wire u0__abc_49347_n3341;
  wire u0__abc_49347_n3342;
  wire u0__abc_49347_n3343;
  wire u0__abc_49347_n3344;
  wire u0__abc_49347_n3345;
  wire u0__abc_49347_n3346;
  wire u0__abc_49347_n3347;
  wire u0__abc_49347_n3348;
  wire u0__abc_49347_n3349;
  wire u0__abc_49347_n3350;
  wire u0__abc_49347_n3351;
  wire u0__abc_49347_n3353;
  wire u0__abc_49347_n3354;
  wire u0__abc_49347_n3355;
  wire u0__abc_49347_n3356;
  wire u0__abc_49347_n3357;
  wire u0__abc_49347_n3358;
  wire u0__abc_49347_n3359;
  wire u0__abc_49347_n3360;
  wire u0__abc_49347_n3361;
  wire u0__abc_49347_n3362;
  wire u0__abc_49347_n3363;
  wire u0__abc_49347_n3364;
  wire u0__abc_49347_n3365;
  wire u0__abc_49347_n3366;
  wire u0__abc_49347_n3367;
  wire u0__abc_49347_n3368;
  wire u0__abc_49347_n3369;
  wire u0__abc_49347_n3370;
  wire u0__abc_49347_n3371;
  wire u0__abc_49347_n3372;
  wire u0__abc_49347_n3373;
  wire u0__abc_49347_n3374;
  wire u0__abc_49347_n3375;
  wire u0__abc_49347_n3377;
  wire u0__abc_49347_n3378;
  wire u0__abc_49347_n3379;
  wire u0__abc_49347_n3380;
  wire u0__abc_49347_n3381;
  wire u0__abc_49347_n3382;
  wire u0__abc_49347_n3383;
  wire u0__abc_49347_n3384;
  wire u0__abc_49347_n3385;
  wire u0__abc_49347_n3386;
  wire u0__abc_49347_n3387;
  wire u0__abc_49347_n3388;
  wire u0__abc_49347_n3389;
  wire u0__abc_49347_n3390;
  wire u0__abc_49347_n3391;
  wire u0__abc_49347_n3392;
  wire u0__abc_49347_n3393;
  wire u0__abc_49347_n3394;
  wire u0__abc_49347_n3395;
  wire u0__abc_49347_n3396;
  wire u0__abc_49347_n3397;
  wire u0__abc_49347_n3398;
  wire u0__abc_49347_n3399;
  wire u0__abc_49347_n3521;
  wire u0__abc_49347_n3522;
  wire u0__abc_49347_n3523;
  wire u0__abc_49347_n3524;
  wire u0__abc_49347_n3525;
  wire u0__abc_49347_n3526;
  wire u0__abc_49347_n3527;
  wire u0__abc_49347_n3528;
  wire u0__abc_49347_n3529;
  wire u0__abc_49347_n3530;
  wire u0__abc_49347_n3531;
  wire u0__abc_49347_n3532;
  wire u0__abc_49347_n3533;
  wire u0__abc_49347_n3534;
  wire u0__abc_49347_n3535;
  wire u0__abc_49347_n3536;
  wire u0__abc_49347_n3537;
  wire u0__abc_49347_n3538;
  wire u0__abc_49347_n3539;
  wire u0__abc_49347_n3540;
  wire u0__abc_49347_n3541;
  wire u0__abc_49347_n3542;
  wire u0__abc_49347_n3543;
  wire u0__abc_49347_n3545;
  wire u0__abc_49347_n3546;
  wire u0__abc_49347_n3547;
  wire u0__abc_49347_n3548;
  wire u0__abc_49347_n3549;
  wire u0__abc_49347_n3550;
  wire u0__abc_49347_n3551;
  wire u0__abc_49347_n3552;
  wire u0__abc_49347_n3553;
  wire u0__abc_49347_n3554;
  wire u0__abc_49347_n3555;
  wire u0__abc_49347_n3556;
  wire u0__abc_49347_n3557;
  wire u0__abc_49347_n3558;
  wire u0__abc_49347_n3559;
  wire u0__abc_49347_n3560;
  wire u0__abc_49347_n3561;
  wire u0__abc_49347_n3562;
  wire u0__abc_49347_n3563;
  wire u0__abc_49347_n3564;
  wire u0__abc_49347_n3565;
  wire u0__abc_49347_n3566;
  wire u0__abc_49347_n3567;
  wire u0__abc_49347_n3569;
  wire u0__abc_49347_n3570;
  wire u0__abc_49347_n3571;
  wire u0__abc_49347_n3572;
  wire u0__abc_49347_n3573;
  wire u0__abc_49347_n3574;
  wire u0__abc_49347_n3575;
  wire u0__abc_49347_n3576;
  wire u0__abc_49347_n3577;
  wire u0__abc_49347_n3578;
  wire u0__abc_49347_n3579;
  wire u0__abc_49347_n3580;
  wire u0__abc_49347_n3581;
  wire u0__abc_49347_n3582;
  wire u0__abc_49347_n3583;
  wire u0__abc_49347_n3584;
  wire u0__abc_49347_n3585;
  wire u0__abc_49347_n3586;
  wire u0__abc_49347_n3587;
  wire u0__abc_49347_n3588;
  wire u0__abc_49347_n3589;
  wire u0__abc_49347_n3590;
  wire u0__abc_49347_n3591;
  wire u0__abc_49347_n3593;
  wire u0__abc_49347_n3594;
  wire u0__abc_49347_n3595;
  wire u0__abc_49347_n3596;
  wire u0__abc_49347_n3597;
  wire u0__abc_49347_n3598;
  wire u0__abc_49347_n3599;
  wire u0__abc_49347_n3600;
  wire u0__abc_49347_n3601;
  wire u0__abc_49347_n3602;
  wire u0__abc_49347_n3603;
  wire u0__abc_49347_n3604;
  wire u0__abc_49347_n3605;
  wire u0__abc_49347_n3606;
  wire u0__abc_49347_n3607;
  wire u0__abc_49347_n3608;
  wire u0__abc_49347_n3609;
  wire u0__abc_49347_n3610;
  wire u0__abc_49347_n3611;
  wire u0__abc_49347_n3612;
  wire u0__abc_49347_n3613;
  wire u0__abc_49347_n3614;
  wire u0__abc_49347_n3615;
  wire u0__abc_49347_n3617;
  wire u0__abc_49347_n3618;
  wire u0__abc_49347_n3619;
  wire u0__abc_49347_n3620;
  wire u0__abc_49347_n3621;
  wire u0__abc_49347_n3622;
  wire u0__abc_49347_n3623;
  wire u0__abc_49347_n3624;
  wire u0__abc_49347_n3625;
  wire u0__abc_49347_n3626;
  wire u0__abc_49347_n3627;
  wire u0__abc_49347_n3628;
  wire u0__abc_49347_n3629;
  wire u0__abc_49347_n3630;
  wire u0__abc_49347_n3631;
  wire u0__abc_49347_n3632;
  wire u0__abc_49347_n3633;
  wire u0__abc_49347_n3634;
  wire u0__abc_49347_n3635;
  wire u0__abc_49347_n3636;
  wire u0__abc_49347_n3637;
  wire u0__abc_49347_n3638;
  wire u0__abc_49347_n3639;
  wire u0__abc_49347_n3641;
  wire u0__abc_49347_n3642;
  wire u0__abc_49347_n3643;
  wire u0__abc_49347_n3644;
  wire u0__abc_49347_n3645;
  wire u0__abc_49347_n3646;
  wire u0__abc_49347_n3647;
  wire u0__abc_49347_n3648;
  wire u0__abc_49347_n3649;
  wire u0__abc_49347_n3650;
  wire u0__abc_49347_n3651;
  wire u0__abc_49347_n3652;
  wire u0__abc_49347_n3653;
  wire u0__abc_49347_n3654;
  wire u0__abc_49347_n3655;
  wire u0__abc_49347_n3656;
  wire u0__abc_49347_n3657;
  wire u0__abc_49347_n3658;
  wire u0__abc_49347_n3659;
  wire u0__abc_49347_n3660;
  wire u0__abc_49347_n3661;
  wire u0__abc_49347_n3662;
  wire u0__abc_49347_n3663;
  wire u0__abc_49347_n3665;
  wire u0__abc_49347_n3666;
  wire u0__abc_49347_n3667;
  wire u0__abc_49347_n3668;
  wire u0__abc_49347_n3669;
  wire u0__abc_49347_n3670;
  wire u0__abc_49347_n3671;
  wire u0__abc_49347_n3672;
  wire u0__abc_49347_n3673;
  wire u0__abc_49347_n3674;
  wire u0__abc_49347_n3675;
  wire u0__abc_49347_n3676;
  wire u0__abc_49347_n3677;
  wire u0__abc_49347_n3678;
  wire u0__abc_49347_n3679;
  wire u0__abc_49347_n3680;
  wire u0__abc_49347_n3681;
  wire u0__abc_49347_n3682;
  wire u0__abc_49347_n3683;
  wire u0__abc_49347_n3684;
  wire u0__abc_49347_n3685;
  wire u0__abc_49347_n3686;
  wire u0__abc_49347_n3687;
  wire u0__abc_49347_n3713;
  wire u0__abc_49347_n3714;
  wire u0__abc_49347_n3715;
  wire u0__abc_49347_n3716;
  wire u0__abc_49347_n3717;
  wire u0__abc_49347_n3718;
  wire u0__abc_49347_n3719;
  wire u0__abc_49347_n3720;
  wire u0__abc_49347_n3721;
  wire u0__abc_49347_n3722;
  wire u0__abc_49347_n3723;
  wire u0__abc_49347_n3724;
  wire u0__abc_49347_n3725;
  wire u0__abc_49347_n3726;
  wire u0__abc_49347_n3727;
  wire u0__abc_49347_n3728;
  wire u0__abc_49347_n3729;
  wire u0__abc_49347_n3730;
  wire u0__abc_49347_n3731;
  wire u0__abc_49347_n3732;
  wire u0__abc_49347_n3733;
  wire u0__abc_49347_n3734;
  wire u0__abc_49347_n3735;
  wire u0__abc_49347_n3737;
  wire u0__abc_49347_n3738;
  wire u0__abc_49347_n3739;
  wire u0__abc_49347_n3740;
  wire u0__abc_49347_n3741;
  wire u0__abc_49347_n3742;
  wire u0__abc_49347_n3743;
  wire u0__abc_49347_n3744;
  wire u0__abc_49347_n3745;
  wire u0__abc_49347_n3746;
  wire u0__abc_49347_n3747;
  wire u0__abc_49347_n3748;
  wire u0__abc_49347_n3749;
  wire u0__abc_49347_n3750;
  wire u0__abc_49347_n3751;
  wire u0__abc_49347_n3752;
  wire u0__abc_49347_n3753;
  wire u0__abc_49347_n3754;
  wire u0__abc_49347_n3755;
  wire u0__abc_49347_n3756;
  wire u0__abc_49347_n3757;
  wire u0__abc_49347_n3758;
  wire u0__abc_49347_n3759;
  wire u0__abc_49347_n3761;
  wire u0__abc_49347_n3762;
  wire u0__abc_49347_n3763;
  wire u0__abc_49347_n3764;
  wire u0__abc_49347_n3765;
  wire u0__abc_49347_n3766;
  wire u0__abc_49347_n3767;
  wire u0__abc_49347_n3768;
  wire u0__abc_49347_n3769;
  wire u0__abc_49347_n3770;
  wire u0__abc_49347_n3771;
  wire u0__abc_49347_n3772;
  wire u0__abc_49347_n3773;
  wire u0__abc_49347_n3774;
  wire u0__abc_49347_n3775;
  wire u0__abc_49347_n3776;
  wire u0__abc_49347_n3777;
  wire u0__abc_49347_n3778;
  wire u0__abc_49347_n3779;
  wire u0__abc_49347_n3780;
  wire u0__abc_49347_n3781;
  wire u0__abc_49347_n3782;
  wire u0__abc_49347_n3783;
  wire u0__abc_49347_n4265;
  wire u0__abc_49347_n4266;
  wire u0__abc_49347_n4267;
  wire u0__abc_49347_n4268;
  wire u0__abc_49347_n4269;
  wire u0__abc_49347_n4270;
  wire u0__abc_49347_n4271;
  wire u0__abc_49347_n4272;
  wire u0__abc_49347_n4273;
  wire u0__abc_49347_n4274;
  wire u0__abc_49347_n4275;
  wire u0__abc_49347_n4276;
  wire u0__abc_49347_n4278;
  wire u0__abc_49347_n4279;
  wire u0__abc_49347_n4280;
  wire u0__abc_49347_n4282;
  wire u0__abc_49347_n4283;
  wire u0__abc_49347_n4285;
  wire u0__abc_49347_n4286;
  wire u0__abc_49347_n4288;
  wire u0__abc_49347_n4289;
  wire u0__abc_49347_n4291;
  wire u0__abc_49347_n4292;
  wire u0__abc_49347_n4294;
  wire u0__abc_49347_n4295;
  wire u0__abc_49347_n4297;
  wire u0__abc_49347_n4298;
  wire u0__abc_49347_n4300;
  wire u0__abc_49347_n4301;
  wire u0__abc_49347_n4303;
  wire u0__abc_49347_n4304;
  wire u0__abc_49347_n4304_bF_buf0;
  wire u0__abc_49347_n4304_bF_buf1;
  wire u0__abc_49347_n4304_bF_buf2;
  wire u0__abc_49347_n4304_bF_buf3;
  wire u0__abc_49347_n4304_bF_buf4;
  wire u0__abc_49347_n4305;
  wire u0__abc_49347_n4307;
  wire u0__abc_49347_n4308;
  wire u0__abc_49347_n4310;
  wire u0__abc_49347_n4311;
  wire u0__abc_49347_n4313;
  wire u0__abc_49347_n4314;
  wire u0__abc_49347_n4316;
  wire u0__abc_49347_n4317;
  wire u0__abc_49347_n4319;
  wire u0__abc_49347_n4320;
  wire u0__abc_49347_n4322;
  wire u0__abc_49347_n4323;
  wire u0__abc_49347_n4325;
  wire u0__abc_49347_n4326;
  wire u0__abc_49347_n4328;
  wire u0__abc_49347_n4329;
  wire u0__abc_49347_n4331;
  wire u0__abc_49347_n4332;
  wire u0__abc_49347_n4334;
  wire u0__abc_49347_n4335;
  wire u0__abc_49347_n4337;
  wire u0__abc_49347_n4338;
  wire u0__abc_49347_n4340;
  wire u0__abc_49347_n4341;
  wire u0__abc_49347_n4343;
  wire u0__abc_49347_n4344;
  wire u0__abc_49347_n4346;
  wire u0__abc_49347_n4347;
  wire u0__abc_49347_n4349;
  wire u0__abc_49347_n4350;
  wire u0__abc_49347_n4352;
  wire u0__abc_49347_n4353;
  wire u0__abc_49347_n4355;
  wire u0__abc_49347_n4356;
  wire u0__abc_49347_n4358;
  wire u0__abc_49347_n4359;
  wire u0__abc_49347_n4361;
  wire u0__abc_49347_n4362;
  wire u0__abc_49347_n4364;
  wire u0__abc_49347_n4365;
  wire u0__abc_49347_n4367;
  wire u0__abc_49347_n4368;
  wire u0__abc_49347_n4370;
  wire u0__abc_49347_n4371;
  wire u0__abc_49347_n4373;
  wire u0__abc_49347_n4374;
  wire u0__abc_49347_n4376;
  wire u0__abc_49347_n4377;
  wire u0__abc_49347_n4379;
  wire u0__abc_49347_n4380;
  wire u0__abc_49347_n4382;
  wire u0__abc_49347_n4383;
  wire u0__abc_49347_n4385;
  wire u0__abc_49347_n4386;
  wire u0__abc_49347_n4388;
  wire u0__abc_49347_n4389;
  wire u0__abc_49347_n4391;
  wire u0__abc_49347_n4392;
  wire u0__abc_49347_n4394;
  wire u0__abc_49347_n4395;
  wire u0__abc_49347_n4397;
  wire u0__abc_49347_n4398;
  wire u0__abc_49347_n4400;
  wire u0__abc_49347_n4401;
  wire u0__abc_49347_n4402;
  wire u0__abc_49347_n4403;
  wire u0__abc_49347_n4404;
  wire u0__abc_49347_n4405;
  wire u0__abc_49347_n4406;
  wire u0__abc_49347_n4407;
  wire u0__abc_49347_n4408;
  wire u0__abc_49347_n4409;
  wire u0__abc_49347_n4410;
  wire u0__abc_49347_n4412;
  wire u0__abc_49347_n4413;
  wire u0__abc_49347_n4415;
  wire u0__abc_49347_n4416;
  wire u0__abc_49347_n4418;
  wire u0__abc_49347_n4419;
  wire u0__abc_49347_n4421;
  wire u0__abc_49347_n4422;
  wire u0__abc_49347_n4424;
  wire u0__abc_49347_n4425;
  wire u0__abc_49347_n4427;
  wire u0__abc_49347_n4428;
  wire u0__abc_49347_n4430;
  wire u0__abc_49347_n4431;
  wire u0__abc_49347_n4433;
  wire u0__abc_49347_n4434;
  wire u0__abc_49347_n4436;
  wire u0__abc_49347_n4437;
  wire u0__abc_49347_n4439;
  wire u0__abc_49347_n4440;
  wire u0__abc_49347_n4442;
  wire u0__abc_49347_n4443;
  wire u0__abc_49347_n4443_bF_buf0;
  wire u0__abc_49347_n4443_bF_buf1;
  wire u0__abc_49347_n4443_bF_buf2;
  wire u0__abc_49347_n4443_bF_buf3;
  wire u0__abc_49347_n4444;
  wire u0__abc_49347_n4444_bF_buf0;
  wire u0__abc_49347_n4444_bF_buf1;
  wire u0__abc_49347_n4444_bF_buf2;
  wire u0__abc_49347_n4444_bF_buf3;
  wire u0__abc_49347_n4445;
  wire u0__abc_49347_n4446;
  wire u0__abc_49347_n4448;
  wire u0__abc_49347_n4449;
  wire u0__abc_49347_n4451;
  wire u0__abc_49347_n4452;
  wire u0__abc_49347_n4454;
  wire u0__abc_49347_n4455;
  wire u0__abc_49347_n4457;
  wire u0__abc_49347_n4458;
  wire u0__abc_49347_n4460;
  wire u0__abc_49347_n4461;
  wire u0__abc_49347_n4463;
  wire u0__abc_49347_n4464;
  wire u0__abc_49347_n4466;
  wire u0__abc_49347_n4467;
  wire u0__abc_49347_n4469;
  wire u0__abc_49347_n4470;
  wire u0__abc_49347_n4472;
  wire u0__abc_49347_n4473;
  wire u0__abc_49347_n4475;
  wire u0__abc_49347_n4476;
  wire u0__abc_49347_n4478;
  wire u0__abc_49347_n4479;
  wire u0__abc_49347_n4481;
  wire u0__abc_49347_n4482;
  wire u0__abc_49347_n4484;
  wire u0__abc_49347_n4485;
  wire u0__abc_49347_n4487;
  wire u0__abc_49347_n4488;
  wire u0__abc_49347_n4490;
  wire u0__abc_49347_n4491;
  wire u0__abc_49347_n4493;
  wire u0__abc_49347_n4494;
  wire u0__abc_49347_n4496;
  wire u0__abc_49347_n4497;
  wire u0__abc_49347_n4499;
  wire u0__abc_49347_n4500;
  wire u0__abc_49347_n4501;
  wire u0__abc_49347_n4502;
  wire u0__abc_49347_n4503;
  wire u0__abc_49347_n4504;
  wire u0__abc_49347_n4505;
  wire u0__abc_49347_n4506;
  wire u0__abc_49347_n4507;
  wire u0__abc_49347_n4507_bF_buf0;
  wire u0__abc_49347_n4507_bF_buf1;
  wire u0__abc_49347_n4507_bF_buf2;
  wire u0__abc_49347_n4507_bF_buf3;
  wire u0__abc_49347_n4508;
  wire u0__abc_49347_n4509;
  wire u0__abc_49347_n4510;
  wire u0__abc_49347_n4511;
  wire u0__abc_49347_n4511_bF_buf0;
  wire u0__abc_49347_n4511_bF_buf1;
  wire u0__abc_49347_n4511_bF_buf2;
  wire u0__abc_49347_n4511_bF_buf3;
  wire u0__abc_49347_n4511_bF_buf4;
  wire u0__abc_49347_n4512;
  wire u0__abc_49347_n4513;
  wire u0__abc_49347_n4514;
  wire u0__abc_49347_n4515;
  wire u0__abc_49347_n4516;
  wire u0__abc_49347_n4516_bF_buf0;
  wire u0__abc_49347_n4516_bF_buf1;
  wire u0__abc_49347_n4516_bF_buf2;
  wire u0__abc_49347_n4516_bF_buf3;
  wire u0__abc_49347_n4516_bF_buf4;
  wire u0__abc_49347_n4517;
  wire u0__abc_49347_n4518;
  wire u0__abc_49347_n4519;
  wire u0__abc_49347_n4519_bF_buf0;
  wire u0__abc_49347_n4519_bF_buf1;
  wire u0__abc_49347_n4519_bF_buf2;
  wire u0__abc_49347_n4519_bF_buf3;
  wire u0__abc_49347_n4519_bF_buf4;
  wire u0__abc_49347_n4520;
  wire u0__abc_49347_n4521;
  wire u0__abc_49347_n4522;
  wire u0__abc_49347_n4523;
  wire u0__abc_49347_n4524;
  wire u0__abc_49347_n4525;
  wire u0__abc_49347_n4526;
  wire u0__abc_49347_n4526_bF_buf0;
  wire u0__abc_49347_n4526_bF_buf1;
  wire u0__abc_49347_n4526_bF_buf2;
  wire u0__abc_49347_n4526_bF_buf3;
  wire u0__abc_49347_n4526_bF_buf4;
  wire u0__abc_49347_n4527;
  wire u0__abc_49347_n4528;
  wire u0__abc_49347_n4528_bF_buf0;
  wire u0__abc_49347_n4528_bF_buf1;
  wire u0__abc_49347_n4528_bF_buf2;
  wire u0__abc_49347_n4528_bF_buf3;
  wire u0__abc_49347_n4528_bF_buf4;
  wire u0__abc_49347_n4529;
  wire u0__abc_49347_n4530;
  wire u0__abc_49347_n4531;
  wire u0__abc_49347_n4531_bF_buf0;
  wire u0__abc_49347_n4531_bF_buf1;
  wire u0__abc_49347_n4531_bF_buf2;
  wire u0__abc_49347_n4531_bF_buf3;
  wire u0__abc_49347_n4531_bF_buf4;
  wire u0__abc_49347_n4532;
  wire u0__abc_49347_n4533;
  wire u0__abc_49347_n4534;
  wire u0__abc_49347_n4535;
  wire u0__abc_49347_n4535_bF_buf0;
  wire u0__abc_49347_n4535_bF_buf1;
  wire u0__abc_49347_n4535_bF_buf2;
  wire u0__abc_49347_n4535_bF_buf3;
  wire u0__abc_49347_n4535_bF_buf4;
  wire u0__abc_49347_n4536;
  wire u0__abc_49347_n4537;
  wire u0__abc_49347_n4537_bF_buf0;
  wire u0__abc_49347_n4537_bF_buf1;
  wire u0__abc_49347_n4537_bF_buf2;
  wire u0__abc_49347_n4537_bF_buf3;
  wire u0__abc_49347_n4537_bF_buf4;
  wire u0__abc_49347_n4538;
  wire u0__abc_49347_n4539;
  wire u0__abc_49347_n4539_bF_buf0;
  wire u0__abc_49347_n4539_bF_buf1;
  wire u0__abc_49347_n4539_bF_buf2;
  wire u0__abc_49347_n4539_bF_buf3;
  wire u0__abc_49347_n4539_bF_buf4;
  wire u0__abc_49347_n4540;
  wire u0__abc_49347_n4541;
  wire u0__abc_49347_n4542;
  wire u0__abc_49347_n4543;
  wire u0__abc_49347_n4544;
  wire u0__abc_49347_n4545;
  wire u0__abc_49347_n4546;
  wire u0__abc_49347_n4547;
  wire u0__abc_49347_n4548;
  wire u0__abc_49347_n4549;
  wire u0__abc_49347_n4550;
  wire u0__abc_49347_n4551;
  wire u0__abc_49347_n4552;
  wire u0__abc_49347_n4553;
  wire u0__abc_49347_n4554;
  wire u0__abc_49347_n4555;
  wire u0__abc_49347_n4556;
  wire u0__abc_49347_n4557;
  wire u0__abc_49347_n4558;
  wire u0__abc_49347_n4559;
  wire u0__abc_49347_n4560;
  wire u0__abc_49347_n4560_bF_buf0;
  wire u0__abc_49347_n4560_bF_buf1;
  wire u0__abc_49347_n4560_bF_buf2;
  wire u0__abc_49347_n4560_bF_buf3;
  wire u0__abc_49347_n4560_bF_buf4;
  wire u0__abc_49347_n4561;
  wire u0__abc_49347_n4562;
  wire u0__abc_49347_n4562_bF_buf0;
  wire u0__abc_49347_n4562_bF_buf1;
  wire u0__abc_49347_n4562_bF_buf2;
  wire u0__abc_49347_n4562_bF_buf3;
  wire u0__abc_49347_n4562_bF_buf4;
  wire u0__abc_49347_n4563;
  wire u0__abc_49347_n4564;
  wire u0__abc_49347_n4565;
  wire u0__abc_49347_n4566;
  wire u0__abc_49347_n4567;
  wire u0__abc_49347_n4567_bF_buf0;
  wire u0__abc_49347_n4567_bF_buf1;
  wire u0__abc_49347_n4567_bF_buf2;
  wire u0__abc_49347_n4567_bF_buf3;
  wire u0__abc_49347_n4567_bF_buf4;
  wire u0__abc_49347_n4568;
  wire u0__abc_49347_n4569;
  wire u0__abc_49347_n4570;
  wire u0__abc_49347_n4571;
  wire u0__abc_49347_n4571_bF_buf0;
  wire u0__abc_49347_n4571_bF_buf1;
  wire u0__abc_49347_n4571_bF_buf2;
  wire u0__abc_49347_n4571_bF_buf3;
  wire u0__abc_49347_n4571_bF_buf4;
  wire u0__abc_49347_n4572;
  wire u0__abc_49347_n4573;
  wire u0__abc_49347_n4574;
  wire u0__abc_49347_n4575;
  wire u0__abc_49347_n4576;
  wire u0__abc_49347_n4577;
  wire u0__abc_49347_n4578;
  wire u0__abc_49347_n4579;
  wire u0__abc_49347_n4580;
  wire u0__abc_49347_n4581;
  wire u0__abc_49347_n4582;
  wire u0__abc_49347_n4582_bF_buf0;
  wire u0__abc_49347_n4582_bF_buf1;
  wire u0__abc_49347_n4582_bF_buf2;
  wire u0__abc_49347_n4582_bF_buf3;
  wire u0__abc_49347_n4582_bF_buf4;
  wire u0__abc_49347_n4583;
  wire u0__abc_49347_n4584;
  wire u0__abc_49347_n4584_bF_buf0;
  wire u0__abc_49347_n4584_bF_buf1;
  wire u0__abc_49347_n4584_bF_buf2;
  wire u0__abc_49347_n4584_bF_buf3;
  wire u0__abc_49347_n4584_bF_buf4;
  wire u0__abc_49347_n4585;
  wire u0__abc_49347_n4586;
  wire u0__abc_49347_n4586_bF_buf0;
  wire u0__abc_49347_n4586_bF_buf1;
  wire u0__abc_49347_n4586_bF_buf2;
  wire u0__abc_49347_n4586_bF_buf3;
  wire u0__abc_49347_n4586_bF_buf4;
  wire u0__abc_49347_n4587;
  wire u0__abc_49347_n4588;
  wire u0__abc_49347_n4589;
  wire u0__abc_49347_n4589_bF_buf0;
  wire u0__abc_49347_n4589_bF_buf1;
  wire u0__abc_49347_n4589_bF_buf2;
  wire u0__abc_49347_n4589_bF_buf3;
  wire u0__abc_49347_n4589_bF_buf4;
  wire u0__abc_49347_n4590;
  wire u0__abc_49347_n4591;
  wire u0__abc_49347_n4592;
  wire u0__abc_49347_n4593;
  wire u0__abc_49347_n4594;
  wire u0__abc_49347_n4595;
  wire u0__abc_49347_n4596;
  wire u0__abc_49347_n4597;
  wire u0__abc_49347_n4598;
  wire u0__abc_49347_n4599;
  wire u0__abc_49347_n4600;
  wire u0__abc_49347_n4601;
  wire u0__abc_49347_n4602;
  wire u0__abc_49347_n4604;
  wire u0__abc_49347_n4605;
  wire u0__abc_49347_n4606;
  wire u0__abc_49347_n4607;
  wire u0__abc_49347_n4608;
  wire u0__abc_49347_n4609;
  wire u0__abc_49347_n4610;
  wire u0__abc_49347_n4611;
  wire u0__abc_49347_n4612;
  wire u0__abc_49347_n4613;
  wire u0__abc_49347_n4614;
  wire u0__abc_49347_n4615;
  wire u0__abc_49347_n4616;
  wire u0__abc_49347_n4617;
  wire u0__abc_49347_n4618;
  wire u0__abc_49347_n4619;
  wire u0__abc_49347_n4620;
  wire u0__abc_49347_n4621;
  wire u0__abc_49347_n4622;
  wire u0__abc_49347_n4623;
  wire u0__abc_49347_n4624;
  wire u0__abc_49347_n4625;
  wire u0__abc_49347_n4626;
  wire u0__abc_49347_n4627;
  wire u0__abc_49347_n4628;
  wire u0__abc_49347_n4629;
  wire u0__abc_49347_n4630;
  wire u0__abc_49347_n4631;
  wire u0__abc_49347_n4632;
  wire u0__abc_49347_n4633;
  wire u0__abc_49347_n4634;
  wire u0__abc_49347_n4635;
  wire u0__abc_49347_n4636;
  wire u0__abc_49347_n4637;
  wire u0__abc_49347_n4638;
  wire u0__abc_49347_n4639;
  wire u0__abc_49347_n4641;
  wire u0__abc_49347_n4642;
  wire u0__abc_49347_n4643;
  wire u0__abc_49347_n4644;
  wire u0__abc_49347_n4645;
  wire u0__abc_49347_n4646;
  wire u0__abc_49347_n4647;
  wire u0__abc_49347_n4648;
  wire u0__abc_49347_n4649;
  wire u0__abc_49347_n4650;
  wire u0__abc_49347_n4651;
  wire u0__abc_49347_n4652;
  wire u0__abc_49347_n4653;
  wire u0__abc_49347_n4654;
  wire u0__abc_49347_n4655;
  wire u0__abc_49347_n4656;
  wire u0__abc_49347_n4657;
  wire u0__abc_49347_n4658;
  wire u0__abc_49347_n4659;
  wire u0__abc_49347_n4660;
  wire u0__abc_49347_n4661;
  wire u0__abc_49347_n4662;
  wire u0__abc_49347_n4663;
  wire u0__abc_49347_n4664;
  wire u0__abc_49347_n4665;
  wire u0__abc_49347_n4666;
  wire u0__abc_49347_n4667;
  wire u0__abc_49347_n4668;
  wire u0__abc_49347_n4669;
  wire u0__abc_49347_n4670;
  wire u0__abc_49347_n4671;
  wire u0__abc_49347_n4672;
  wire u0__abc_49347_n4673;
  wire u0__abc_49347_n4674;
  wire u0__abc_49347_n4675;
  wire u0__abc_49347_n4676;
  wire u0__abc_49347_n4678;
  wire u0__abc_49347_n4679;
  wire u0__abc_49347_n4680;
  wire u0__abc_49347_n4681;
  wire u0__abc_49347_n4682;
  wire u0__abc_49347_n4683;
  wire u0__abc_49347_n4684;
  wire u0__abc_49347_n4685;
  wire u0__abc_49347_n4686;
  wire u0__abc_49347_n4687;
  wire u0__abc_49347_n4688;
  wire u0__abc_49347_n4689;
  wire u0__abc_49347_n4690;
  wire u0__abc_49347_n4691;
  wire u0__abc_49347_n4692;
  wire u0__abc_49347_n4693;
  wire u0__abc_49347_n4694;
  wire u0__abc_49347_n4695;
  wire u0__abc_49347_n4696;
  wire u0__abc_49347_n4697;
  wire u0__abc_49347_n4698;
  wire u0__abc_49347_n4699;
  wire u0__abc_49347_n4700;
  wire u0__abc_49347_n4701;
  wire u0__abc_49347_n4702;
  wire u0__abc_49347_n4703;
  wire u0__abc_49347_n4704;
  wire u0__abc_49347_n4705;
  wire u0__abc_49347_n4706;
  wire u0__abc_49347_n4707;
  wire u0__abc_49347_n4708;
  wire u0__abc_49347_n4709;
  wire u0__abc_49347_n4710;
  wire u0__abc_49347_n4711;
  wire u0__abc_49347_n4712;
  wire u0__abc_49347_n4713;
  wire u0__abc_49347_n4715;
  wire u0__abc_49347_n4716;
  wire u0__abc_49347_n4717;
  wire u0__abc_49347_n4718;
  wire u0__abc_49347_n4719;
  wire u0__abc_49347_n4720;
  wire u0__abc_49347_n4721;
  wire u0__abc_49347_n4722;
  wire u0__abc_49347_n4723;
  wire u0__abc_49347_n4724;
  wire u0__abc_49347_n4725;
  wire u0__abc_49347_n4726;
  wire u0__abc_49347_n4727;
  wire u0__abc_49347_n4728;
  wire u0__abc_49347_n4729;
  wire u0__abc_49347_n4730;
  wire u0__abc_49347_n4731;
  wire u0__abc_49347_n4732;
  wire u0__abc_49347_n4733;
  wire u0__abc_49347_n4734;
  wire u0__abc_49347_n4735;
  wire u0__abc_49347_n4736;
  wire u0__abc_49347_n4737;
  wire u0__abc_49347_n4738;
  wire u0__abc_49347_n4739;
  wire u0__abc_49347_n4740;
  wire u0__abc_49347_n4741;
  wire u0__abc_49347_n4742;
  wire u0__abc_49347_n4743;
  wire u0__abc_49347_n4744;
  wire u0__abc_49347_n4745;
  wire u0__abc_49347_n4746;
  wire u0__abc_49347_n4747;
  wire u0__abc_49347_n4748;
  wire u0__abc_49347_n4749;
  wire u0__abc_49347_n4750;
  wire u0__abc_49347_n4752;
  wire u0__abc_49347_n4753;
  wire u0__abc_49347_n4754;
  wire u0__abc_49347_n4755;
  wire u0__abc_49347_n4756;
  wire u0__abc_49347_n4757;
  wire u0__abc_49347_n4758;
  wire u0__abc_49347_n4759;
  wire u0__abc_49347_n4760;
  wire u0__abc_49347_n4761;
  wire u0__abc_49347_n4762;
  wire u0__abc_49347_n4763;
  wire u0__abc_49347_n4764;
  wire u0__abc_49347_n4765;
  wire u0__abc_49347_n4766;
  wire u0__abc_49347_n4767;
  wire u0__abc_49347_n4768;
  wire u0__abc_49347_n4769;
  wire u0__abc_49347_n4770;
  wire u0__abc_49347_n4771;
  wire u0__abc_49347_n4772;
  wire u0__abc_49347_n4773;
  wire u0__abc_49347_n4774;
  wire u0__abc_49347_n4775;
  wire u0__abc_49347_n4776;
  wire u0__abc_49347_n4777;
  wire u0__abc_49347_n4778;
  wire u0__abc_49347_n4779;
  wire u0__abc_49347_n4780;
  wire u0__abc_49347_n4781;
  wire u0__abc_49347_n4782;
  wire u0__abc_49347_n4783;
  wire u0__abc_49347_n4784;
  wire u0__abc_49347_n4785;
  wire u0__abc_49347_n4786;
  wire u0__abc_49347_n4787;
  wire u0__abc_49347_n4789;
  wire u0__abc_49347_n4790;
  wire u0__abc_49347_n4791;
  wire u0__abc_49347_n4792;
  wire u0__abc_49347_n4793;
  wire u0__abc_49347_n4794;
  wire u0__abc_49347_n4795;
  wire u0__abc_49347_n4796;
  wire u0__abc_49347_n4797;
  wire u0__abc_49347_n4798;
  wire u0__abc_49347_n4799;
  wire u0__abc_49347_n4800;
  wire u0__abc_49347_n4801;
  wire u0__abc_49347_n4802;
  wire u0__abc_49347_n4803;
  wire u0__abc_49347_n4804;
  wire u0__abc_49347_n4805;
  wire u0__abc_49347_n4806;
  wire u0__abc_49347_n4807;
  wire u0__abc_49347_n4808;
  wire u0__abc_49347_n4809;
  wire u0__abc_49347_n4810;
  wire u0__abc_49347_n4811;
  wire u0__abc_49347_n4812;
  wire u0__abc_49347_n4813;
  wire u0__abc_49347_n4814;
  wire u0__abc_49347_n4815;
  wire u0__abc_49347_n4816;
  wire u0__abc_49347_n4817;
  wire u0__abc_49347_n4818;
  wire u0__abc_49347_n4819;
  wire u0__abc_49347_n4820;
  wire u0__abc_49347_n4821;
  wire u0__abc_49347_n4822;
  wire u0__abc_49347_n4823;
  wire u0__abc_49347_n4824;
  wire u0__abc_49347_n4826;
  wire u0__abc_49347_n4827;
  wire u0__abc_49347_n4828;
  wire u0__abc_49347_n4829;
  wire u0__abc_49347_n4830;
  wire u0__abc_49347_n4831;
  wire u0__abc_49347_n4832;
  wire u0__abc_49347_n4833;
  wire u0__abc_49347_n4834;
  wire u0__abc_49347_n4835;
  wire u0__abc_49347_n4836;
  wire u0__abc_49347_n4837;
  wire u0__abc_49347_n4838;
  wire u0__abc_49347_n4839;
  wire u0__abc_49347_n4840;
  wire u0__abc_49347_n4841;
  wire u0__abc_49347_n4842;
  wire u0__abc_49347_n4843;
  wire u0__abc_49347_n4844;
  wire u0__abc_49347_n4845;
  wire u0__abc_49347_n4846;
  wire u0__abc_49347_n4847;
  wire u0__abc_49347_n4848;
  wire u0__abc_49347_n4849;
  wire u0__abc_49347_n4850;
  wire u0__abc_49347_n4851;
  wire u0__abc_49347_n4852;
  wire u0__abc_49347_n4853;
  wire u0__abc_49347_n4854;
  wire u0__abc_49347_n4855;
  wire u0__abc_49347_n4856;
  wire u0__abc_49347_n4857;
  wire u0__abc_49347_n4858;
  wire u0__abc_49347_n4859;
  wire u0__abc_49347_n4860;
  wire u0__abc_49347_n4861;
  wire u0__abc_49347_n4863;
  wire u0__abc_49347_n4864;
  wire u0__abc_49347_n4865;
  wire u0__abc_49347_n4866;
  wire u0__abc_49347_n4867;
  wire u0__abc_49347_n4868;
  wire u0__abc_49347_n4869;
  wire u0__abc_49347_n4870;
  wire u0__abc_49347_n4871;
  wire u0__abc_49347_n4872;
  wire u0__abc_49347_n4873;
  wire u0__abc_49347_n4874;
  wire u0__abc_49347_n4875;
  wire u0__abc_49347_n4876;
  wire u0__abc_49347_n4877;
  wire u0__abc_49347_n4878;
  wire u0__abc_49347_n4879;
  wire u0__abc_49347_n4880;
  wire u0__abc_49347_n4881;
  wire u0__abc_49347_n4882;
  wire u0__abc_49347_n4883;
  wire u0__abc_49347_n4884;
  wire u0__abc_49347_n4885;
  wire u0__abc_49347_n4886;
  wire u0__abc_49347_n4887;
  wire u0__abc_49347_n4888;
  wire u0__abc_49347_n4889;
  wire u0__abc_49347_n4890;
  wire u0__abc_49347_n4891;
  wire u0__abc_49347_n4892;
  wire u0__abc_49347_n4893;
  wire u0__abc_49347_n4894;
  wire u0__abc_49347_n4895;
  wire u0__abc_49347_n4896;
  wire u0__abc_49347_n4897;
  wire u0__abc_49347_n4898;
  wire u0__abc_49347_n4900;
  wire u0__abc_49347_n4901;
  wire u0__abc_49347_n4902;
  wire u0__abc_49347_n4903;
  wire u0__abc_49347_n4904;
  wire u0__abc_49347_n4905;
  wire u0__abc_49347_n4906;
  wire u0__abc_49347_n4907;
  wire u0__abc_49347_n4908;
  wire u0__abc_49347_n4909;
  wire u0__abc_49347_n4910;
  wire u0__abc_49347_n4911;
  wire u0__abc_49347_n4912;
  wire u0__abc_49347_n4913;
  wire u0__abc_49347_n4914;
  wire u0__abc_49347_n4915;
  wire u0__abc_49347_n4916;
  wire u0__abc_49347_n4917;
  wire u0__abc_49347_n4918;
  wire u0__abc_49347_n4919;
  wire u0__abc_49347_n4920;
  wire u0__abc_49347_n4921;
  wire u0__abc_49347_n4922;
  wire u0__abc_49347_n4923;
  wire u0__abc_49347_n4924;
  wire u0__abc_49347_n4925;
  wire u0__abc_49347_n4926;
  wire u0__abc_49347_n4927;
  wire u0__abc_49347_n4928;
  wire u0__abc_49347_n4929;
  wire u0__abc_49347_n4930;
  wire u0__abc_49347_n4931;
  wire u0__abc_49347_n4932;
  wire u0__abc_49347_n4933;
  wire u0__abc_49347_n4934;
  wire u0__abc_49347_n4935;
  wire u0__abc_49347_n4937;
  wire u0__abc_49347_n4938;
  wire u0__abc_49347_n4939;
  wire u0__abc_49347_n4940;
  wire u0__abc_49347_n4941;
  wire u0__abc_49347_n4942;
  wire u0__abc_49347_n4943;
  wire u0__abc_49347_n4944;
  wire u0__abc_49347_n4945;
  wire u0__abc_49347_n4946;
  wire u0__abc_49347_n4947;
  wire u0__abc_49347_n4948;
  wire u0__abc_49347_n4949;
  wire u0__abc_49347_n4950;
  wire u0__abc_49347_n4951;
  wire u0__abc_49347_n4952;
  wire u0__abc_49347_n4953;
  wire u0__abc_49347_n4954;
  wire u0__abc_49347_n4955;
  wire u0__abc_49347_n4956;
  wire u0__abc_49347_n4957;
  wire u0__abc_49347_n4958;
  wire u0__abc_49347_n4959;
  wire u0__abc_49347_n4960;
  wire u0__abc_49347_n4961;
  wire u0__abc_49347_n4962;
  wire u0__abc_49347_n4963;
  wire u0__abc_49347_n4964;
  wire u0__abc_49347_n4965;
  wire u0__abc_49347_n4966;
  wire u0__abc_49347_n4967;
  wire u0__abc_49347_n4968;
  wire u0__abc_49347_n4969;
  wire u0__abc_49347_n4970;
  wire u0__abc_49347_n4971;
  wire u0__abc_49347_n4972;
  wire u0__abc_49347_n4974;
  wire u0__abc_49347_n4975;
  wire u0__abc_49347_n4976;
  wire u0__abc_49347_n4977;
  wire u0__abc_49347_n4978;
  wire u0__abc_49347_n4979;
  wire u0__abc_49347_n4980;
  wire u0__abc_49347_n4981;
  wire u0__abc_49347_n4982;
  wire u0__abc_49347_n4983;
  wire u0__abc_49347_n4984;
  wire u0__abc_49347_n4985;
  wire u0__abc_49347_n4986;
  wire u0__abc_49347_n4987;
  wire u0__abc_49347_n4988;
  wire u0__abc_49347_n4989;
  wire u0__abc_49347_n4990;
  wire u0__abc_49347_n4991;
  wire u0__abc_49347_n4992;
  wire u0__abc_49347_n4993;
  wire u0__abc_49347_n4994;
  wire u0__abc_49347_n4995;
  wire u0__abc_49347_n4996;
  wire u0__abc_49347_n4997;
  wire u0__abc_49347_n4998;
  wire u0__abc_49347_n4999;
  wire u0__abc_49347_n5000;
  wire u0__abc_49347_n5001;
  wire u0__abc_49347_n5002;
  wire u0__abc_49347_n5003;
  wire u0__abc_49347_n5004;
  wire u0__abc_49347_n5005;
  wire u0__abc_49347_n5007;
  wire u0__abc_49347_n5008;
  wire u0__abc_49347_n5009;
  wire u0__abc_49347_n5010;
  wire u0__abc_49347_n5011;
  wire u0__abc_49347_n5012;
  wire u0__abc_49347_n5013;
  wire u0__abc_49347_n5014;
  wire u0__abc_49347_n5015;
  wire u0__abc_49347_n5016;
  wire u0__abc_49347_n5017;
  wire u0__abc_49347_n5018;
  wire u0__abc_49347_n5019;
  wire u0__abc_49347_n5020;
  wire u0__abc_49347_n5021;
  wire u0__abc_49347_n5022;
  wire u0__abc_49347_n5023;
  wire u0__abc_49347_n5024;
  wire u0__abc_49347_n5025;
  wire u0__abc_49347_n5026;
  wire u0__abc_49347_n5027;
  wire u0__abc_49347_n5028;
  wire u0__abc_49347_n5029;
  wire u0__abc_49347_n5030;
  wire u0__abc_49347_n5031;
  wire u0__abc_49347_n5032;
  wire u0__abc_49347_n5033;
  wire u0__abc_49347_n5034;
  wire u0__abc_49347_n5035;
  wire u0__abc_49347_n5036;
  wire u0__abc_49347_n5037;
  wire u0__abc_49347_n5038;
  wire u0__abc_49347_n5040;
  wire u0__abc_49347_n5041;
  wire u0__abc_49347_n5042;
  wire u0__abc_49347_n5043;
  wire u0__abc_49347_n5044;
  wire u0__abc_49347_n5045;
  wire u0__abc_49347_n5046;
  wire u0__abc_49347_n5047;
  wire u0__abc_49347_n5048;
  wire u0__abc_49347_n5049;
  wire u0__abc_49347_n5050;
  wire u0__abc_49347_n5051;
  wire u0__abc_49347_n5052;
  wire u0__abc_49347_n5053;
  wire u0__abc_49347_n5054;
  wire u0__abc_49347_n5055;
  wire u0__abc_49347_n5056;
  wire u0__abc_49347_n5057;
  wire u0__abc_49347_n5058;
  wire u0__abc_49347_n5059;
  wire u0__abc_49347_n5060;
  wire u0__abc_49347_n5061;
  wire u0__abc_49347_n5062;
  wire u0__abc_49347_n5063;
  wire u0__abc_49347_n5064;
  wire u0__abc_49347_n5065;
  wire u0__abc_49347_n5066;
  wire u0__abc_49347_n5067;
  wire u0__abc_49347_n5068;
  wire u0__abc_49347_n5069;
  wire u0__abc_49347_n5070;
  wire u0__abc_49347_n5071;
  wire u0__abc_49347_n5073;
  wire u0__abc_49347_n5074;
  wire u0__abc_49347_n5075;
  wire u0__abc_49347_n5076;
  wire u0__abc_49347_n5077;
  wire u0__abc_49347_n5078;
  wire u0__abc_49347_n5079;
  wire u0__abc_49347_n5080;
  wire u0__abc_49347_n5081;
  wire u0__abc_49347_n5082;
  wire u0__abc_49347_n5083;
  wire u0__abc_49347_n5084;
  wire u0__abc_49347_n5085;
  wire u0__abc_49347_n5086;
  wire u0__abc_49347_n5087;
  wire u0__abc_49347_n5088;
  wire u0__abc_49347_n5089;
  wire u0__abc_49347_n5090;
  wire u0__abc_49347_n5091;
  wire u0__abc_49347_n5092;
  wire u0__abc_49347_n5093;
  wire u0__abc_49347_n5094;
  wire u0__abc_49347_n5095;
  wire u0__abc_49347_n5096;
  wire u0__abc_49347_n5097;
  wire u0__abc_49347_n5098;
  wire u0__abc_49347_n5099;
  wire u0__abc_49347_n5100;
  wire u0__abc_49347_n5101;
  wire u0__abc_49347_n5102;
  wire u0__abc_49347_n5103;
  wire u0__abc_49347_n5104;
  wire u0__abc_49347_n5106;
  wire u0__abc_49347_n5107;
  wire u0__abc_49347_n5108;
  wire u0__abc_49347_n5109;
  wire u0__abc_49347_n5110;
  wire u0__abc_49347_n5111;
  wire u0__abc_49347_n5112;
  wire u0__abc_49347_n5113;
  wire u0__abc_49347_n5114;
  wire u0__abc_49347_n5115;
  wire u0__abc_49347_n5116;
  wire u0__abc_49347_n5117;
  wire u0__abc_49347_n5118;
  wire u0__abc_49347_n5119;
  wire u0__abc_49347_n5120;
  wire u0__abc_49347_n5121;
  wire u0__abc_49347_n5122;
  wire u0__abc_49347_n5123;
  wire u0__abc_49347_n5124;
  wire u0__abc_49347_n5125;
  wire u0__abc_49347_n5126;
  wire u0__abc_49347_n5127;
  wire u0__abc_49347_n5128;
  wire u0__abc_49347_n5129;
  wire u0__abc_49347_n5130;
  wire u0__abc_49347_n5131;
  wire u0__abc_49347_n5132;
  wire u0__abc_49347_n5133;
  wire u0__abc_49347_n5134;
  wire u0__abc_49347_n5135;
  wire u0__abc_49347_n5136;
  wire u0__abc_49347_n5137;
  wire u0__abc_49347_n5139;
  wire u0__abc_49347_n5140;
  wire u0__abc_49347_n5141;
  wire u0__abc_49347_n5142;
  wire u0__abc_49347_n5143;
  wire u0__abc_49347_n5144;
  wire u0__abc_49347_n5145;
  wire u0__abc_49347_n5146;
  wire u0__abc_49347_n5147;
  wire u0__abc_49347_n5148;
  wire u0__abc_49347_n5149;
  wire u0__abc_49347_n5150;
  wire u0__abc_49347_n5151;
  wire u0__abc_49347_n5152;
  wire u0__abc_49347_n5153;
  wire u0__abc_49347_n5154;
  wire u0__abc_49347_n5155;
  wire u0__abc_49347_n5156;
  wire u0__abc_49347_n5157;
  wire u0__abc_49347_n5158;
  wire u0__abc_49347_n5159;
  wire u0__abc_49347_n5160;
  wire u0__abc_49347_n5161;
  wire u0__abc_49347_n5162;
  wire u0__abc_49347_n5163;
  wire u0__abc_49347_n5164;
  wire u0__abc_49347_n5165;
  wire u0__abc_49347_n5166;
  wire u0__abc_49347_n5167;
  wire u0__abc_49347_n5168;
  wire u0__abc_49347_n5169;
  wire u0__abc_49347_n5170;
  wire u0__abc_49347_n5172;
  wire u0__abc_49347_n5173;
  wire u0__abc_49347_n5174;
  wire u0__abc_49347_n5175;
  wire u0__abc_49347_n5176;
  wire u0__abc_49347_n5177;
  wire u0__abc_49347_n5178;
  wire u0__abc_49347_n5179;
  wire u0__abc_49347_n5180;
  wire u0__abc_49347_n5181;
  wire u0__abc_49347_n5182;
  wire u0__abc_49347_n5183;
  wire u0__abc_49347_n5184;
  wire u0__abc_49347_n5185;
  wire u0__abc_49347_n5186;
  wire u0__abc_49347_n5187;
  wire u0__abc_49347_n5188;
  wire u0__abc_49347_n5189;
  wire u0__abc_49347_n5190;
  wire u0__abc_49347_n5191;
  wire u0__abc_49347_n5192;
  wire u0__abc_49347_n5193;
  wire u0__abc_49347_n5194;
  wire u0__abc_49347_n5195;
  wire u0__abc_49347_n5196;
  wire u0__abc_49347_n5197;
  wire u0__abc_49347_n5198;
  wire u0__abc_49347_n5199;
  wire u0__abc_49347_n5200;
  wire u0__abc_49347_n5201;
  wire u0__abc_49347_n5202;
  wire u0__abc_49347_n5203;
  wire u0__abc_49347_n5205;
  wire u0__abc_49347_n5206;
  wire u0__abc_49347_n5207;
  wire u0__abc_49347_n5208;
  wire u0__abc_49347_n5209;
  wire u0__abc_49347_n5210;
  wire u0__abc_49347_n5211;
  wire u0__abc_49347_n5212;
  wire u0__abc_49347_n5213;
  wire u0__abc_49347_n5214;
  wire u0__abc_49347_n5215;
  wire u0__abc_49347_n5216;
  wire u0__abc_49347_n5217;
  wire u0__abc_49347_n5218;
  wire u0__abc_49347_n5219;
  wire u0__abc_49347_n5220;
  wire u0__abc_49347_n5221;
  wire u0__abc_49347_n5222;
  wire u0__abc_49347_n5223;
  wire u0__abc_49347_n5224;
  wire u0__abc_49347_n5225;
  wire u0__abc_49347_n5226;
  wire u0__abc_49347_n5227;
  wire u0__abc_49347_n5228;
  wire u0__abc_49347_n5229;
  wire u0__abc_49347_n5230;
  wire u0__abc_49347_n5231;
  wire u0__abc_49347_n5232;
  wire u0__abc_49347_n5233;
  wire u0__abc_49347_n5234;
  wire u0__abc_49347_n5235;
  wire u0__abc_49347_n5236;
  wire u0__abc_49347_n5238;
  wire u0__abc_49347_n5239;
  wire u0__abc_49347_n5240;
  wire u0__abc_49347_n5241;
  wire u0__abc_49347_n5242;
  wire u0__abc_49347_n5243;
  wire u0__abc_49347_n5244;
  wire u0__abc_49347_n5245;
  wire u0__abc_49347_n5246;
  wire u0__abc_49347_n5247;
  wire u0__abc_49347_n5248;
  wire u0__abc_49347_n5249;
  wire u0__abc_49347_n5250;
  wire u0__abc_49347_n5251;
  wire u0__abc_49347_n5252;
  wire u0__abc_49347_n5253;
  wire u0__abc_49347_n5254;
  wire u0__abc_49347_n5255;
  wire u0__abc_49347_n5256;
  wire u0__abc_49347_n5257;
  wire u0__abc_49347_n5258;
  wire u0__abc_49347_n5259;
  wire u0__abc_49347_n5260;
  wire u0__abc_49347_n5261;
  wire u0__abc_49347_n5262;
  wire u0__abc_49347_n5263;
  wire u0__abc_49347_n5264;
  wire u0__abc_49347_n5265;
  wire u0__abc_49347_n5266;
  wire u0__abc_49347_n5267;
  wire u0__abc_49347_n5268;
  wire u0__abc_49347_n5269;
  wire u0__abc_49347_n5271;
  wire u0__abc_49347_n5272;
  wire u0__abc_49347_n5273;
  wire u0__abc_49347_n5274;
  wire u0__abc_49347_n5275;
  wire u0__abc_49347_n5276;
  wire u0__abc_49347_n5277;
  wire u0__abc_49347_n5278;
  wire u0__abc_49347_n5279;
  wire u0__abc_49347_n5280;
  wire u0__abc_49347_n5281;
  wire u0__abc_49347_n5282;
  wire u0__abc_49347_n5283;
  wire u0__abc_49347_n5284;
  wire u0__abc_49347_n5285;
  wire u0__abc_49347_n5286;
  wire u0__abc_49347_n5287;
  wire u0__abc_49347_n5288;
  wire u0__abc_49347_n5289;
  wire u0__abc_49347_n5290;
  wire u0__abc_49347_n5291;
  wire u0__abc_49347_n5292;
  wire u0__abc_49347_n5293;
  wire u0__abc_49347_n5294;
  wire u0__abc_49347_n5295;
  wire u0__abc_49347_n5296;
  wire u0__abc_49347_n5297;
  wire u0__abc_49347_n5298;
  wire u0__abc_49347_n5299;
  wire u0__abc_49347_n5300;
  wire u0__abc_49347_n5301;
  wire u0__abc_49347_n5302;
  wire u0__abc_49347_n5304;
  wire u0__abc_49347_n5305;
  wire u0__abc_49347_n5306;
  wire u0__abc_49347_n5307;
  wire u0__abc_49347_n5308;
  wire u0__abc_49347_n5309;
  wire u0__abc_49347_n5310;
  wire u0__abc_49347_n5311;
  wire u0__abc_49347_n5312;
  wire u0__abc_49347_n5313;
  wire u0__abc_49347_n5314;
  wire u0__abc_49347_n5315;
  wire u0__abc_49347_n5316;
  wire u0__abc_49347_n5317;
  wire u0__abc_49347_n5318;
  wire u0__abc_49347_n5319;
  wire u0__abc_49347_n5320;
  wire u0__abc_49347_n5321;
  wire u0__abc_49347_n5322;
  wire u0__abc_49347_n5323;
  wire u0__abc_49347_n5324;
  wire u0__abc_49347_n5325;
  wire u0__abc_49347_n5326;
  wire u0__abc_49347_n5327;
  wire u0__abc_49347_n5328;
  wire u0__abc_49347_n5329;
  wire u0__abc_49347_n5330;
  wire u0__abc_49347_n5331;
  wire u0__abc_49347_n5332;
  wire u0__abc_49347_n5333;
  wire u0__abc_49347_n5334;
  wire u0__abc_49347_n5335;
  wire u0__abc_49347_n5337;
  wire u0__abc_49347_n5338;
  wire u0__abc_49347_n5339;
  wire u0__abc_49347_n5340;
  wire u0__abc_49347_n5341;
  wire u0__abc_49347_n5342;
  wire u0__abc_49347_n5343;
  wire u0__abc_49347_n5344;
  wire u0__abc_49347_n5345;
  wire u0__abc_49347_n5346;
  wire u0__abc_49347_n5347;
  wire u0__abc_49347_n5348;
  wire u0__abc_49347_n5349;
  wire u0__abc_49347_n5350;
  wire u0__abc_49347_n5351;
  wire u0__abc_49347_n5352;
  wire u0__abc_49347_n5353;
  wire u0__abc_49347_n5354;
  wire u0__abc_49347_n5355;
  wire u0__abc_49347_n5356;
  wire u0__abc_49347_n5357;
  wire u0__abc_49347_n5358;
  wire u0__abc_49347_n5359;
  wire u0__abc_49347_n5360;
  wire u0__abc_49347_n5361;
  wire u0__abc_49347_n5362;
  wire u0__abc_49347_n5363;
  wire u0__abc_49347_n5364;
  wire u0__abc_49347_n5365;
  wire u0__abc_49347_n5366;
  wire u0__abc_49347_n5367;
  wire u0__abc_49347_n5368;
  wire u0__abc_49347_n5370;
  wire u0__abc_49347_n5371;
  wire u0__abc_49347_n5372;
  wire u0__abc_49347_n5373;
  wire u0__abc_49347_n5374;
  wire u0__abc_49347_n5375;
  wire u0__abc_49347_n5376;
  wire u0__abc_49347_n5377;
  wire u0__abc_49347_n5378;
  wire u0__abc_49347_n5379;
  wire u0__abc_49347_n5380;
  wire u0__abc_49347_n5381;
  wire u0__abc_49347_n5382;
  wire u0__abc_49347_n5383;
  wire u0__abc_49347_n5384;
  wire u0__abc_49347_n5385;
  wire u0__abc_49347_n5386;
  wire u0__abc_49347_n5387;
  wire u0__abc_49347_n5388;
  wire u0__abc_49347_n5389;
  wire u0__abc_49347_n5390;
  wire u0__abc_49347_n5391;
  wire u0__abc_49347_n5392;
  wire u0__abc_49347_n5393;
  wire u0__abc_49347_n5394;
  wire u0__abc_49347_n5395;
  wire u0__abc_49347_n5396;
  wire u0__abc_49347_n5397;
  wire u0__abc_49347_n5398;
  wire u0__abc_49347_n5399;
  wire u0__abc_49347_n5400;
  wire u0__abc_49347_n5401;
  wire u0__abc_49347_n5403;
  wire u0__abc_49347_n5404;
  wire u0__abc_49347_n5405;
  wire u0__abc_49347_n5406;
  wire u0__abc_49347_n5407;
  wire u0__abc_49347_n5408;
  wire u0__abc_49347_n5409;
  wire u0__abc_49347_n5410;
  wire u0__abc_49347_n5411;
  wire u0__abc_49347_n5412;
  wire u0__abc_49347_n5413;
  wire u0__abc_49347_n5414;
  wire u0__abc_49347_n5415;
  wire u0__abc_49347_n5416;
  wire u0__abc_49347_n5417;
  wire u0__abc_49347_n5418;
  wire u0__abc_49347_n5419;
  wire u0__abc_49347_n5420;
  wire u0__abc_49347_n5421;
  wire u0__abc_49347_n5422;
  wire u0__abc_49347_n5423;
  wire u0__abc_49347_n5424;
  wire u0__abc_49347_n5425;
  wire u0__abc_49347_n5426;
  wire u0__abc_49347_n5427;
  wire u0__abc_49347_n5428;
  wire u0__abc_49347_n5429;
  wire u0__abc_49347_n5430;
  wire u0__abc_49347_n5431;
  wire u0__abc_49347_n5432;
  wire u0__abc_49347_n5433;
  wire u0__abc_49347_n5434;
  wire u0__abc_49347_n5435;
  wire u0__abc_49347_n5436;
  wire u0__abc_49347_n5438;
  wire u0__abc_49347_n5439;
  wire u0__abc_49347_n5440;
  wire u0__abc_49347_n5441;
  wire u0__abc_49347_n5442;
  wire u0__abc_49347_n5443;
  wire u0__abc_49347_n5444;
  wire u0__abc_49347_n5445;
  wire u0__abc_49347_n5446;
  wire u0__abc_49347_n5447;
  wire u0__abc_49347_n5448;
  wire u0__abc_49347_n5449;
  wire u0__abc_49347_n5450;
  wire u0__abc_49347_n5451;
  wire u0__abc_49347_n5452;
  wire u0__abc_49347_n5453;
  wire u0__abc_49347_n5454;
  wire u0__abc_49347_n5455;
  wire u0__abc_49347_n5456;
  wire u0__abc_49347_n5457;
  wire u0__abc_49347_n5458;
  wire u0__abc_49347_n5459;
  wire u0__abc_49347_n5460;
  wire u0__abc_49347_n5461;
  wire u0__abc_49347_n5462;
  wire u0__abc_49347_n5463;
  wire u0__abc_49347_n5464;
  wire u0__abc_49347_n5465;
  wire u0__abc_49347_n5466;
  wire u0__abc_49347_n5467;
  wire u0__abc_49347_n5468;
  wire u0__abc_49347_n5469;
  wire u0__abc_49347_n5470;
  wire u0__abc_49347_n5471;
  wire u0__abc_49347_n5473;
  wire u0__abc_49347_n5474;
  wire u0__abc_49347_n5475;
  wire u0__abc_49347_n5476;
  wire u0__abc_49347_n5477;
  wire u0__abc_49347_n5478;
  wire u0__abc_49347_n5479;
  wire u0__abc_49347_n5480;
  wire u0__abc_49347_n5481;
  wire u0__abc_49347_n5482;
  wire u0__abc_49347_n5483;
  wire u0__abc_49347_n5484;
  wire u0__abc_49347_n5485;
  wire u0__abc_49347_n5486;
  wire u0__abc_49347_n5487;
  wire u0__abc_49347_n5488;
  wire u0__abc_49347_n5489;
  wire u0__abc_49347_n5490;
  wire u0__abc_49347_n5491;
  wire u0__abc_49347_n5492;
  wire u0__abc_49347_n5493;
  wire u0__abc_49347_n5494;
  wire u0__abc_49347_n5495;
  wire u0__abc_49347_n5496;
  wire u0__abc_49347_n5497;
  wire u0__abc_49347_n5498;
  wire u0__abc_49347_n5499;
  wire u0__abc_49347_n5500;
  wire u0__abc_49347_n5501;
  wire u0__abc_49347_n5502;
  wire u0__abc_49347_n5503;
  wire u0__abc_49347_n5504;
  wire u0__abc_49347_n5505;
  wire u0__abc_49347_n5506;
  wire u0__abc_49347_n5508;
  wire u0__abc_49347_n5509;
  wire u0__abc_49347_n5510;
  wire u0__abc_49347_n5511;
  wire u0__abc_49347_n5512;
  wire u0__abc_49347_n5513;
  wire u0__abc_49347_n5514;
  wire u0__abc_49347_n5515;
  wire u0__abc_49347_n5516;
  wire u0__abc_49347_n5517;
  wire u0__abc_49347_n5518;
  wire u0__abc_49347_n5519;
  wire u0__abc_49347_n5520;
  wire u0__abc_49347_n5521;
  wire u0__abc_49347_n5522;
  wire u0__abc_49347_n5523;
  wire u0__abc_49347_n5524;
  wire u0__abc_49347_n5525;
  wire u0__abc_49347_n5526;
  wire u0__abc_49347_n5527;
  wire u0__abc_49347_n5528;
  wire u0__abc_49347_n5529;
  wire u0__abc_49347_n5530;
  wire u0__abc_49347_n5531;
  wire u0__abc_49347_n5532;
  wire u0__abc_49347_n5533;
  wire u0__abc_49347_n5534;
  wire u0__abc_49347_n5535;
  wire u0__abc_49347_n5536;
  wire u0__abc_49347_n5537;
  wire u0__abc_49347_n5538;
  wire u0__abc_49347_n5539;
  wire u0__abc_49347_n5540;
  wire u0__abc_49347_n5541;
  wire u0__abc_49347_n5543;
  wire u0__abc_49347_n5544;
  wire u0__abc_49347_n5545;
  wire u0__abc_49347_n5546;
  wire u0__abc_49347_n5547;
  wire u0__abc_49347_n5548;
  wire u0__abc_49347_n5549;
  wire u0__abc_49347_n5550;
  wire u0__abc_49347_n5551;
  wire u0__abc_49347_n5552;
  wire u0__abc_49347_n5553;
  wire u0__abc_49347_n5554;
  wire u0__abc_49347_n5555;
  wire u0__abc_49347_n5556;
  wire u0__abc_49347_n5557;
  wire u0__abc_49347_n5558;
  wire u0__abc_49347_n5559;
  wire u0__abc_49347_n5560;
  wire u0__abc_49347_n5561;
  wire u0__abc_49347_n5562;
  wire u0__abc_49347_n5563;
  wire u0__abc_49347_n5564;
  wire u0__abc_49347_n5565;
  wire u0__abc_49347_n5566;
  wire u0__abc_49347_n5567;
  wire u0__abc_49347_n5568;
  wire u0__abc_49347_n5569;
  wire u0__abc_49347_n5570;
  wire u0__abc_49347_n5571;
  wire u0__abc_49347_n5572;
  wire u0__abc_49347_n5573;
  wire u0__abc_49347_n5574;
  wire u0__abc_49347_n5575;
  wire u0__abc_49347_n5576;
  wire u0__abc_49347_n5578;
  wire u0__abc_49347_n5579;
  wire u0__abc_49347_n5580;
  wire u0__abc_49347_n5581;
  wire u0__abc_49347_n5582;
  wire u0__abc_49347_n5583;
  wire u0__abc_49347_n5584;
  wire u0__abc_49347_n5585;
  wire u0__abc_49347_n5586;
  wire u0__abc_49347_n5587;
  wire u0__abc_49347_n5588;
  wire u0__abc_49347_n5589;
  wire u0__abc_49347_n5590;
  wire u0__abc_49347_n5591;
  wire u0__abc_49347_n5592;
  wire u0__abc_49347_n5593;
  wire u0__abc_49347_n5594;
  wire u0__abc_49347_n5595;
  wire u0__abc_49347_n5596;
  wire u0__abc_49347_n5597;
  wire u0__abc_49347_n5598;
  wire u0__abc_49347_n5599;
  wire u0__abc_49347_n5600;
  wire u0__abc_49347_n5601;
  wire u0__abc_49347_n5602;
  wire u0__abc_49347_n5603;
  wire u0__abc_49347_n5604;
  wire u0__abc_49347_n5605;
  wire u0__abc_49347_n5606;
  wire u0__abc_49347_n5607;
  wire u0__abc_49347_n5608;
  wire u0__abc_49347_n5609;
  wire u0__abc_49347_n5610;
  wire u0__abc_49347_n5611;
  wire u0__abc_49347_n5613;
  wire u0__abc_49347_n5614;
  wire u0__abc_49347_n5615;
  wire u0__abc_49347_n5616;
  wire u0__abc_49347_n5617;
  wire u0__abc_49347_n5618;
  wire u0__abc_49347_n5619;
  wire u0__abc_49347_n5620;
  wire u0__abc_49347_n5621;
  wire u0__abc_49347_n5622;
  wire u0__abc_49347_n5623;
  wire u0__abc_49347_n5624;
  wire u0__abc_49347_n5625;
  wire u0__abc_49347_n5626;
  wire u0__abc_49347_n5627;
  wire u0__abc_49347_n5628;
  wire u0__abc_49347_n5629;
  wire u0__abc_49347_n5630;
  wire u0__abc_49347_n5631;
  wire u0__abc_49347_n5632;
  wire u0__abc_49347_n5633;
  wire u0__abc_49347_n5634;
  wire u0__abc_49347_n5635;
  wire u0__abc_49347_n5636;
  wire u0__abc_49347_n5637;
  wire u0__abc_49347_n5638;
  wire u0__abc_49347_n5639;
  wire u0__abc_49347_n5640;
  wire u0__abc_49347_n5641;
  wire u0__abc_49347_n5642;
  wire u0__abc_49347_n5643;
  wire u0__abc_49347_n5644;
  wire u0__abc_49347_n5645;
  wire u0__abc_49347_n5646;
  wire u0__abc_49347_n5648;
  wire u0__abc_49347_n5649;
  wire u0__abc_49347_n5650;
  wire u0__abc_49347_n5651;
  wire u0__abc_49347_n5652;
  wire u0__abc_49347_n5653;
  wire u0__abc_49347_n5654;
  wire u0__abc_49347_n5655;
  wire u0__abc_49347_n5656;
  wire u0__abc_49347_n5657;
  wire u0__abc_49347_n5658;
  wire u0__abc_49347_n5659;
  wire u0__abc_49347_n5660;
  wire u0__abc_49347_n5661;
  wire u0__abc_49347_n5662;
  wire u0__abc_49347_n5663;
  wire u0__abc_49347_n5664;
  wire u0__abc_49347_n5665;
  wire u0__abc_49347_n5666;
  wire u0__abc_49347_n5667;
  wire u0__abc_49347_n5668;
  wire u0__abc_49347_n5669;
  wire u0__abc_49347_n5670;
  wire u0__abc_49347_n5671;
  wire u0__abc_49347_n5672;
  wire u0__abc_49347_n5673;
  wire u0__abc_49347_n5674;
  wire u0__abc_49347_n5675;
  wire u0__abc_49347_n5676;
  wire u0__abc_49347_n5677;
  wire u0__abc_49347_n5678;
  wire u0__abc_49347_n5679;
  wire u0__abc_49347_n5680;
  wire u0__abc_49347_n5681;
  wire u0__abc_49347_n5683;
  wire u0__abc_49347_n5684;
  wire u0__abc_49347_n5685;
  wire u0__abc_49347_n5686;
  wire u0__abc_49347_n5687;
  wire u0__abc_49347_n5692;
  wire u0__abc_49347_n5693;
  wire u0__abc_49347_n5694;
  wire u0__abc_49347_n5695;
  wire u0__abc_49347_n5696;
  wire u0__abc_49347_n5698;
  wire u0__abc_49347_n5699;
  wire u0__abc_49347_n5700;
  wire u0__abc_49347_n5701;
  wire u0__abc_49347_n5702;
  wire u0__abc_49347_n5704;
  wire u0__abc_49347_n5705;
  wire u0__abc_49347_n5706;
  wire u0__abc_49347_n5707;
  wire u0__abc_49347_n5708;
  wire u0__abc_49347_n5710;
  wire u0__abc_49347_n5711;
  wire u0__abc_49347_n5712;
  wire u0__abc_49347_n5713;
  wire u0__abc_49347_n5714;
  wire u0__abc_49347_n5716;
  wire u0__abc_49347_n5717;
  wire u0__abc_49347_n5718;
  wire u0__abc_49347_n5719;
  wire u0__abc_49347_n5720;
  wire u0__abc_49347_n5722;
  wire u0__abc_49347_n5723;
  wire u0__abc_49347_n5724;
  wire u0__abc_49347_n5725;
  wire u0__abc_49347_n5726;
  wire u0__abc_49347_n5728;
  wire u0__abc_49347_n5729;
  wire u0__abc_49347_n5730;
  wire u0__abc_49347_n5731;
  wire u0__abc_49347_n5732;
  wire u0__abc_49347_n5734;
  wire u0__abc_49347_n5735;
  wire u0__abc_49347_n5736;
  wire u0__abc_49347_n5737;
  wire u0__abc_49347_n5738;
  wire u0__abc_49347_n5740;
  wire u0__abc_49347_n5741;
  wire u0__abc_49347_n5742;
  wire u0__abc_49347_n5743;
  wire u0__abc_49347_n5744;
  wire u0__abc_49347_n5745;
  wire u0__abc_49347_n5746;
  wire u0__abc_49347_n5748;
  wire u0__abc_49347_n5749;
  wire u0__abc_49347_n5750;
  wire u0__abc_49347_n5751;
  wire u0__abc_49347_n5752;
  wire u0__abc_49347_n5753;
  wire u0__abc_49347_n5755;
  wire u0__abc_49347_n5756;
  wire u0__abc_49347_n5757;
  wire u0__abc_49347_n5758;
  wire u0__abc_49347_n5759;
  wire u0__abc_49347_n5760;
  wire u0_cs0;
  wire u0_cs0_bF_buf0;
  wire u0_cs0_bF_buf1;
  wire u0_cs0_bF_buf2;
  wire u0_cs0_bF_buf3;
  wire u0_cs0_bF_buf4;
  wire u0_cs0_bF_buf5;
  wire u0_cs1;
  wire u0_cs1_bF_buf0;
  wire u0_cs1_bF_buf1;
  wire u0_cs1_bF_buf2;
  wire u0_cs1_bF_buf3;
  wire u0_cs1_bF_buf4;
  wire u0_cs1_bF_buf5;
  wire u0_cs2;
  wire u0_cs2_bF_buf0;
  wire u0_cs2_bF_buf1;
  wire u0_cs2_bF_buf2;
  wire u0_cs2_bF_buf3;
  wire u0_cs2_bF_buf4;
  wire u0_cs2_bF_buf5;
  wire u0_cs3;
  wire u0_cs3_bF_buf0;
  wire u0_cs3_bF_buf1;
  wire u0_cs3_bF_buf2;
  wire u0_cs3_bF_buf3;
  wire u0_cs3_bF_buf4;
  wire u0_cs3_bF_buf5;
  wire u0_cs4;
  wire u0_cs4_bF_buf0;
  wire u0_cs4_bF_buf1;
  wire u0_cs4_bF_buf2;
  wire u0_cs4_bF_buf3;
  wire u0_cs4_bF_buf4;
  wire u0_cs4_bF_buf5;
  wire u0_cs5;
  wire u0_cs5_bF_buf0;
  wire u0_cs5_bF_buf1;
  wire u0_cs5_bF_buf2;
  wire u0_cs5_bF_buf3;
  wire u0_cs5_bF_buf4;
  wire u0_cs5_bF_buf5;
  wire u0_cs_0__FF_INPUT;
  wire u0_cs_1__FF_INPUT;
  wire u0_cs_2__FF_INPUT;
  wire u0_cs_3__FF_INPUT;
  wire u0_cs_4__FF_INPUT;
  wire u0_cs_5__FF_INPUT;
  wire u0_cs_6__FF_INPUT;
  wire u0_cs_7__FF_INPUT;
  wire u0_csc0_0_;
  wire u0_csc0_10_;
  wire u0_csc0_11_;
  wire u0_csc0_12_;
  wire u0_csc0_13_;
  wire u0_csc0_14_;
  wire u0_csc0_15_;
  wire u0_csc0_16_;
  wire u0_csc0_17_;
  wire u0_csc0_18_;
  wire u0_csc0_19_;
  wire u0_csc0_1_;
  wire u0_csc0_20_;
  wire u0_csc0_21_;
  wire u0_csc0_22_;
  wire u0_csc0_23_;
  wire u0_csc0_24_;
  wire u0_csc0_25_;
  wire u0_csc0_26_;
  wire u0_csc0_27_;
  wire u0_csc0_28_;
  wire u0_csc0_29_;
  wire u0_csc0_2_;
  wire u0_csc0_30_;
  wire u0_csc0_31_;
  wire u0_csc0_3_;
  wire u0_csc0_4_;
  wire u0_csc0_5_;
  wire u0_csc0_6_;
  wire u0_csc0_7_;
  wire u0_csc0_8_;
  wire u0_csc0_9_;
  wire u0_csc1_0_;
  wire u0_csc1_10_;
  wire u0_csc1_11_;
  wire u0_csc1_12_;
  wire u0_csc1_13_;
  wire u0_csc1_14_;
  wire u0_csc1_15_;
  wire u0_csc1_16_;
  wire u0_csc1_17_;
  wire u0_csc1_18_;
  wire u0_csc1_19_;
  wire u0_csc1_1_;
  wire u0_csc1_20_;
  wire u0_csc1_21_;
  wire u0_csc1_22_;
  wire u0_csc1_23_;
  wire u0_csc1_24_;
  wire u0_csc1_25_;
  wire u0_csc1_26_;
  wire u0_csc1_27_;
  wire u0_csc1_28_;
  wire u0_csc1_29_;
  wire u0_csc1_2_;
  wire u0_csc1_30_;
  wire u0_csc1_31_;
  wire u0_csc1_3_;
  wire u0_csc1_4_;
  wire u0_csc1_5_;
  wire u0_csc1_6_;
  wire u0_csc1_7_;
  wire u0_csc1_8_;
  wire u0_csc1_9_;
  wire u0_csc2_0_;
  wire u0_csc2_10_;
  wire u0_csc2_11_;
  wire u0_csc2_12_;
  wire u0_csc2_13_;
  wire u0_csc2_14_;
  wire u0_csc2_15_;
  wire u0_csc2_16_;
  wire u0_csc2_17_;
  wire u0_csc2_18_;
  wire u0_csc2_19_;
  wire u0_csc2_1_;
  wire u0_csc2_20_;
  wire u0_csc2_21_;
  wire u0_csc2_22_;
  wire u0_csc2_23_;
  wire u0_csc2_24_;
  wire u0_csc2_25_;
  wire u0_csc2_26_;
  wire u0_csc2_27_;
  wire u0_csc2_28_;
  wire u0_csc2_29_;
  wire u0_csc2_2_;
  wire u0_csc2_30_;
  wire u0_csc2_31_;
  wire u0_csc2_3_;
  wire u0_csc2_4_;
  wire u0_csc2_5_;
  wire u0_csc2_6_;
  wire u0_csc2_7_;
  wire u0_csc2_8_;
  wire u0_csc2_9_;
  wire u0_csc3_0_;
  wire u0_csc3_10_;
  wire u0_csc3_11_;
  wire u0_csc3_12_;
  wire u0_csc3_13_;
  wire u0_csc3_14_;
  wire u0_csc3_15_;
  wire u0_csc3_16_;
  wire u0_csc3_17_;
  wire u0_csc3_18_;
  wire u0_csc3_19_;
  wire u0_csc3_1_;
  wire u0_csc3_20_;
  wire u0_csc3_21_;
  wire u0_csc3_22_;
  wire u0_csc3_23_;
  wire u0_csc3_24_;
  wire u0_csc3_25_;
  wire u0_csc3_26_;
  wire u0_csc3_27_;
  wire u0_csc3_28_;
  wire u0_csc3_29_;
  wire u0_csc3_2_;
  wire u0_csc3_30_;
  wire u0_csc3_31_;
  wire u0_csc3_3_;
  wire u0_csc3_4_;
  wire u0_csc3_5_;
  wire u0_csc3_6_;
  wire u0_csc3_7_;
  wire u0_csc3_8_;
  wire u0_csc3_9_;
  wire u0_csc4_0_;
  wire u0_csc4_10_;
  wire u0_csc4_11_;
  wire u0_csc4_12_;
  wire u0_csc4_13_;
  wire u0_csc4_14_;
  wire u0_csc4_15_;
  wire u0_csc4_16_;
  wire u0_csc4_17_;
  wire u0_csc4_18_;
  wire u0_csc4_19_;
  wire u0_csc4_1_;
  wire u0_csc4_20_;
  wire u0_csc4_21_;
  wire u0_csc4_22_;
  wire u0_csc4_23_;
  wire u0_csc4_24_;
  wire u0_csc4_25_;
  wire u0_csc4_26_;
  wire u0_csc4_27_;
  wire u0_csc4_28_;
  wire u0_csc4_29_;
  wire u0_csc4_2_;
  wire u0_csc4_30_;
  wire u0_csc4_31_;
  wire u0_csc4_3_;
  wire u0_csc4_4_;
  wire u0_csc4_5_;
  wire u0_csc4_6_;
  wire u0_csc4_7_;
  wire u0_csc4_8_;
  wire u0_csc4_9_;
  wire u0_csc5_0_;
  wire u0_csc5_10_;
  wire u0_csc5_11_;
  wire u0_csc5_12_;
  wire u0_csc5_13_;
  wire u0_csc5_14_;
  wire u0_csc5_15_;
  wire u0_csc5_16_;
  wire u0_csc5_17_;
  wire u0_csc5_18_;
  wire u0_csc5_19_;
  wire u0_csc5_1_;
  wire u0_csc5_20_;
  wire u0_csc5_21_;
  wire u0_csc5_22_;
  wire u0_csc5_23_;
  wire u0_csc5_24_;
  wire u0_csc5_25_;
  wire u0_csc5_26_;
  wire u0_csc5_27_;
  wire u0_csc5_28_;
  wire u0_csc5_29_;
  wire u0_csc5_2_;
  wire u0_csc5_30_;
  wire u0_csc5_31_;
  wire u0_csc5_3_;
  wire u0_csc5_4_;
  wire u0_csc5_5_;
  wire u0_csc5_6_;
  wire u0_csc5_7_;
  wire u0_csc5_8_;
  wire u0_csc5_9_;
  wire u0_csc_10__FF_INPUT;
  wire u0_csc_11__FF_INPUT;
  wire u0_csc_1__FF_INPUT;
  wire u0_csc_2__FF_INPUT;
  wire u0_csc_3__FF_INPUT;
  wire u0_csc_4__FF_INPUT;
  wire u0_csc_5__FF_INPUT;
  wire u0_csc_6__FF_INPUT;
  wire u0_csc_7__FF_INPUT;
  wire u0_csc_9__FF_INPUT;
  wire u0_csc_mask_0_;
  wire u0_csc_mask_10_;
  wire u0_csc_mask_1_;
  wire u0_csc_mask_2_;
  wire u0_csc_mask_3_;
  wire u0_csc_mask_4_;
  wire u0_csc_mask_5_;
  wire u0_csc_mask_6_;
  wire u0_csc_mask_7_;
  wire u0_csc_mask_8_;
  wire u0_csc_mask_9_;
  wire u0_csc_mask_r_0__FF_INPUT;
  wire u0_csc_mask_r_10__FF_INPUT;
  wire u0_csc_mask_r_1__FF_INPUT;
  wire u0_csc_mask_r_2__FF_INPUT;
  wire u0_csc_mask_r_3__FF_INPUT;
  wire u0_csc_mask_r_4__FF_INPUT;
  wire u0_csc_mask_r_5__FF_INPUT;
  wire u0_csc_mask_r_6__FF_INPUT;
  wire u0_csc_mask_r_7__FF_INPUT;
  wire u0_csc_mask_r_8__FF_INPUT;
  wire u0_csc_mask_r_9__FF_INPUT;
  wire u0_csr_0_;
  wire u0_csr_3_;
  wire u0_csr_4_;
  wire u0_csr_5_;
  wire u0_csr_6_;
  wire u0_csr_7_;
  wire u0_csr_r2_0__FF_INPUT;
  wire u0_csr_r2_1__FF_INPUT;
  wire u0_csr_r2_2__FF_INPUT;
  wire u0_csr_r2_3__FF_INPUT;
  wire u0_csr_r2_4__FF_INPUT;
  wire u0_csr_r2_5__FF_INPUT;
  wire u0_csr_r2_6__FF_INPUT;
  wire u0_csr_r2_7__FF_INPUT;
  wire u0_csr_r_0__FF_INPUT;
  wire u0_csr_r_1__FF_INPUT;
  wire u0_csr_r_2__FF_INPUT;
  wire u0_csr_r_3__FF_INPUT;
  wire u0_csr_r_4__FF_INPUT;
  wire u0_csr_r_5__FF_INPUT;
  wire u0_csr_r_6__FF_INPUT;
  wire u0_csr_r_7__FF_INPUT;
  wire u0_csr_r_8__FF_INPUT;
  wire u0_csr_r_9__FF_INPUT;
  wire u0_init_ack0;
  wire u0_init_ack1;
  wire u0_init_ack2;
  wire u0_init_ack3;
  wire u0_init_ack4;
  wire u0_init_ack5;
  wire u0_init_ack_r;
  wire u0_init_req0;
  wire u0_init_req1;
  wire u0_init_req2;
  wire u0_init_req3;
  wire u0_init_req4;
  wire u0_init_req5;
  wire u0_init_req_FF_INPUT;
  wire u0_lmr_ack0;
  wire u0_lmr_ack1;
  wire u0_lmr_ack2;
  wire u0_lmr_ack3;
  wire u0_lmr_ack4;
  wire u0_lmr_ack5;
  wire u0_lmr_ack_r;
  wire u0_lmr_req0;
  wire u0_lmr_req1;
  wire u0_lmr_req2;
  wire u0_lmr_req3;
  wire u0_lmr_req4;
  wire u0_lmr_req5;
  wire u0_lmr_req_FF_INPUT;
  wire u0_poc_0__FF_INPUT;
  wire u0_poc_10__FF_INPUT;
  wire u0_poc_11__FF_INPUT;
  wire u0_poc_12__FF_INPUT;
  wire u0_poc_13__FF_INPUT;
  wire u0_poc_14__FF_INPUT;
  wire u0_poc_15__FF_INPUT;
  wire u0_poc_16__FF_INPUT;
  wire u0_poc_17__FF_INPUT;
  wire u0_poc_18__FF_INPUT;
  wire u0_poc_19__FF_INPUT;
  wire u0_poc_1__FF_INPUT;
  wire u0_poc_20__FF_INPUT;
  wire u0_poc_21__FF_INPUT;
  wire u0_poc_22__FF_INPUT;
  wire u0_poc_23__FF_INPUT;
  wire u0_poc_24__FF_INPUT;
  wire u0_poc_25__FF_INPUT;
  wire u0_poc_26__FF_INPUT;
  wire u0_poc_27__FF_INPUT;
  wire u0_poc_28__FF_INPUT;
  wire u0_poc_29__FF_INPUT;
  wire u0_poc_2__FF_INPUT;
  wire u0_poc_30__FF_INPUT;
  wire u0_poc_31__FF_INPUT;
  wire u0_poc_3__FF_INPUT;
  wire u0_poc_4__FF_INPUT;
  wire u0_poc_5__FF_INPUT;
  wire u0_poc_6__FF_INPUT;
  wire u0_poc_7__FF_INPUT;
  wire u0_poc_8__FF_INPUT;
  wire u0_poc_9__FF_INPUT;
  wire u0_rf_we;
  wire u0_rf_we_FF_INPUT;
  wire u0_rst_r1;
  wire u0_rst_r2;
  wire u0_rst_r3;
  wire u0_rst_r3_bF_buf0;
  wire u0_rst_r3_bF_buf1;
  wire u0_rst_r3_bF_buf2;
  wire u0_rst_r3_bF_buf3;
  wire u0_rst_r3_bF_buf4;
  wire u0_sp_csc_10__FF_INPUT;
  wire u0_sp_csc_1__FF_INPUT;
  wire u0_sp_csc_2__FF_INPUT;
  wire u0_sp_csc_3__FF_INPUT;
  wire u0_sp_csc_4__FF_INPUT;
  wire u0_sp_csc_5__FF_INPUT;
  wire u0_sp_csc_6__FF_INPUT;
  wire u0_sp_csc_7__FF_INPUT;
  wire u0_sp_csc_9__FF_INPUT;
  wire u0_sp_tms_0__FF_INPUT;
  wire u0_sp_tms_10__FF_INPUT;
  wire u0_sp_tms_11__FF_INPUT;
  wire u0_sp_tms_12__FF_INPUT;
  wire u0_sp_tms_13__FF_INPUT;
  wire u0_sp_tms_14__FF_INPUT;
  wire u0_sp_tms_15__FF_INPUT;
  wire u0_sp_tms_16__FF_INPUT;
  wire u0_sp_tms_17__FF_INPUT;
  wire u0_sp_tms_18__FF_INPUT;
  wire u0_sp_tms_19__FF_INPUT;
  wire u0_sp_tms_1__FF_INPUT;
  wire u0_sp_tms_20__FF_INPUT;
  wire u0_sp_tms_21__FF_INPUT;
  wire u0_sp_tms_22__FF_INPUT;
  wire u0_sp_tms_23__FF_INPUT;
  wire u0_sp_tms_24__FF_INPUT;
  wire u0_sp_tms_25__FF_INPUT;
  wire u0_sp_tms_26__FF_INPUT;
  wire u0_sp_tms_27__FF_INPUT;
  wire u0_sp_tms_2__FF_INPUT;
  wire u0_sp_tms_3__FF_INPUT;
  wire u0_sp_tms_4__FF_INPUT;
  wire u0_sp_tms_5__FF_INPUT;
  wire u0_sp_tms_6__FF_INPUT;
  wire u0_sp_tms_7__FF_INPUT;
  wire u0_sp_tms_8__FF_INPUT;
  wire u0_sp_tms_9__FF_INPUT;
  wire u0_spec_req_cs_0__FF_INPUT;
  wire u0_spec_req_cs_1__FF_INPUT;
  wire u0_spec_req_cs_2__FF_INPUT;
  wire u0_spec_req_cs_3__FF_INPUT;
  wire u0_spec_req_cs_4__FF_INPUT;
  wire u0_spec_req_cs_5__FF_INPUT;
  wire u0_spec_req_cs_6__FF_INPUT;
  wire u0_spec_req_cs_7__FF_INPUT;
  wire u0_sreq_cs_le;
  wire u0_sreq_cs_le_FF_INPUT;
  wire u0_tms0_0_;
  wire u0_tms0_10_;
  wire u0_tms0_11_;
  wire u0_tms0_12_;
  wire u0_tms0_13_;
  wire u0_tms0_14_;
  wire u0_tms0_15_;
  wire u0_tms0_16_;
  wire u0_tms0_17_;
  wire u0_tms0_18_;
  wire u0_tms0_19_;
  wire u0_tms0_1_;
  wire u0_tms0_20_;
  wire u0_tms0_21_;
  wire u0_tms0_22_;
  wire u0_tms0_23_;
  wire u0_tms0_24_;
  wire u0_tms0_25_;
  wire u0_tms0_26_;
  wire u0_tms0_27_;
  wire u0_tms0_28_;
  wire u0_tms0_29_;
  wire u0_tms0_2_;
  wire u0_tms0_30_;
  wire u0_tms0_31_;
  wire u0_tms0_3_;
  wire u0_tms0_4_;
  wire u0_tms0_5_;
  wire u0_tms0_6_;
  wire u0_tms0_7_;
  wire u0_tms0_8_;
  wire u0_tms0_9_;
  wire u0_tms1_0_;
  wire u0_tms1_10_;
  wire u0_tms1_11_;
  wire u0_tms1_12_;
  wire u0_tms1_13_;
  wire u0_tms1_14_;
  wire u0_tms1_15_;
  wire u0_tms1_16_;
  wire u0_tms1_17_;
  wire u0_tms1_18_;
  wire u0_tms1_19_;
  wire u0_tms1_1_;
  wire u0_tms1_20_;
  wire u0_tms1_21_;
  wire u0_tms1_22_;
  wire u0_tms1_23_;
  wire u0_tms1_24_;
  wire u0_tms1_25_;
  wire u0_tms1_26_;
  wire u0_tms1_27_;
  wire u0_tms1_28_;
  wire u0_tms1_29_;
  wire u0_tms1_2_;
  wire u0_tms1_30_;
  wire u0_tms1_31_;
  wire u0_tms1_3_;
  wire u0_tms1_4_;
  wire u0_tms1_5_;
  wire u0_tms1_6_;
  wire u0_tms1_7_;
  wire u0_tms1_8_;
  wire u0_tms1_9_;
  wire u0_tms2_0_;
  wire u0_tms2_10_;
  wire u0_tms2_11_;
  wire u0_tms2_12_;
  wire u0_tms2_13_;
  wire u0_tms2_14_;
  wire u0_tms2_15_;
  wire u0_tms2_16_;
  wire u0_tms2_17_;
  wire u0_tms2_18_;
  wire u0_tms2_19_;
  wire u0_tms2_1_;
  wire u0_tms2_20_;
  wire u0_tms2_21_;
  wire u0_tms2_22_;
  wire u0_tms2_23_;
  wire u0_tms2_24_;
  wire u0_tms2_25_;
  wire u0_tms2_26_;
  wire u0_tms2_27_;
  wire u0_tms2_28_;
  wire u0_tms2_29_;
  wire u0_tms2_2_;
  wire u0_tms2_30_;
  wire u0_tms2_31_;
  wire u0_tms2_3_;
  wire u0_tms2_4_;
  wire u0_tms2_5_;
  wire u0_tms2_6_;
  wire u0_tms2_7_;
  wire u0_tms2_8_;
  wire u0_tms2_9_;
  wire u0_tms3_0_;
  wire u0_tms3_10_;
  wire u0_tms3_11_;
  wire u0_tms3_12_;
  wire u0_tms3_13_;
  wire u0_tms3_14_;
  wire u0_tms3_15_;
  wire u0_tms3_16_;
  wire u0_tms3_17_;
  wire u0_tms3_18_;
  wire u0_tms3_19_;
  wire u0_tms3_1_;
  wire u0_tms3_20_;
  wire u0_tms3_21_;
  wire u0_tms3_22_;
  wire u0_tms3_23_;
  wire u0_tms3_24_;
  wire u0_tms3_25_;
  wire u0_tms3_26_;
  wire u0_tms3_27_;
  wire u0_tms3_28_;
  wire u0_tms3_29_;
  wire u0_tms3_2_;
  wire u0_tms3_30_;
  wire u0_tms3_31_;
  wire u0_tms3_3_;
  wire u0_tms3_4_;
  wire u0_tms3_5_;
  wire u0_tms3_6_;
  wire u0_tms3_7_;
  wire u0_tms3_8_;
  wire u0_tms3_9_;
  wire u0_tms4_0_;
  wire u0_tms4_10_;
  wire u0_tms4_11_;
  wire u0_tms4_12_;
  wire u0_tms4_13_;
  wire u0_tms4_14_;
  wire u0_tms4_15_;
  wire u0_tms4_16_;
  wire u0_tms4_17_;
  wire u0_tms4_18_;
  wire u0_tms4_19_;
  wire u0_tms4_1_;
  wire u0_tms4_20_;
  wire u0_tms4_21_;
  wire u0_tms4_22_;
  wire u0_tms4_23_;
  wire u0_tms4_24_;
  wire u0_tms4_25_;
  wire u0_tms4_26_;
  wire u0_tms4_27_;
  wire u0_tms4_28_;
  wire u0_tms4_29_;
  wire u0_tms4_2_;
  wire u0_tms4_30_;
  wire u0_tms4_31_;
  wire u0_tms4_3_;
  wire u0_tms4_4_;
  wire u0_tms4_5_;
  wire u0_tms4_6_;
  wire u0_tms4_7_;
  wire u0_tms4_8_;
  wire u0_tms4_9_;
  wire u0_tms5_0_;
  wire u0_tms5_10_;
  wire u0_tms5_11_;
  wire u0_tms5_12_;
  wire u0_tms5_13_;
  wire u0_tms5_14_;
  wire u0_tms5_15_;
  wire u0_tms5_16_;
  wire u0_tms5_17_;
  wire u0_tms5_18_;
  wire u0_tms5_19_;
  wire u0_tms5_1_;
  wire u0_tms5_20_;
  wire u0_tms5_21_;
  wire u0_tms5_22_;
  wire u0_tms5_23_;
  wire u0_tms5_24_;
  wire u0_tms5_25_;
  wire u0_tms5_26_;
  wire u0_tms5_27_;
  wire u0_tms5_28_;
  wire u0_tms5_29_;
  wire u0_tms5_2_;
  wire u0_tms5_30_;
  wire u0_tms5_31_;
  wire u0_tms5_3_;
  wire u0_tms5_4_;
  wire u0_tms5_5_;
  wire u0_tms5_6_;
  wire u0_tms5_7_;
  wire u0_tms5_8_;
  wire u0_tms5_9_;
  wire u0_tms_0__FF_INPUT;
  wire u0_tms_10__FF_INPUT;
  wire u0_tms_11__FF_INPUT;
  wire u0_tms_12__FF_INPUT;
  wire u0_tms_13__FF_INPUT;
  wire u0_tms_14__FF_INPUT;
  wire u0_tms_15__FF_INPUT;
  wire u0_tms_16__FF_INPUT;
  wire u0_tms_17__FF_INPUT;
  wire u0_tms_18__FF_INPUT;
  wire u0_tms_19__FF_INPUT;
  wire u0_tms_1__FF_INPUT;
  wire u0_tms_20__FF_INPUT;
  wire u0_tms_21__FF_INPUT;
  wire u0_tms_22__FF_INPUT;
  wire u0_tms_23__FF_INPUT;
  wire u0_tms_24__FF_INPUT;
  wire u0_tms_25__FF_INPUT;
  wire u0_tms_26__FF_INPUT;
  wire u0_tms_27__FF_INPUT;
  wire u0_tms_2__FF_INPUT;
  wire u0_tms_3__FF_INPUT;
  wire u0_tms_4__FF_INPUT;
  wire u0_tms_5__FF_INPUT;
  wire u0_tms_6__FF_INPUT;
  wire u0_tms_7__FF_INPUT;
  wire u0_tms_8__FF_INPUT;
  wire u0_tms_9__FF_INPUT;
  wire u0_u0__abc_43300_n201_1;
  wire u0_u0__abc_43300_n202_1;
  wire u0_u0__abc_43300_n203;
  wire u0_u0__abc_43300_n204_1;
  wire u0_u0__abc_43300_n205_1;
  wire u0_u0__abc_43300_n206;
  wire u0_u0__abc_43300_n207_1;
  wire u0_u0__abc_43300_n208_1;
  wire u0_u0__abc_43300_n209;
  wire u0_u0__abc_43300_n211_1;
  wire u0_u0__abc_43300_n212;
  wire u0_u0__abc_43300_n213_1;
  wire u0_u0__abc_43300_n214_1;
  wire u0_u0__abc_43300_n215;
  wire u0_u0__abc_43300_n217_1;
  wire u0_u0__abc_43300_n218;
  wire u0_u0__abc_43300_n218_bF_buf0;
  wire u0_u0__abc_43300_n218_bF_buf1;
  wire u0_u0__abc_43300_n218_bF_buf2;
  wire u0_u0__abc_43300_n218_bF_buf3;
  wire u0_u0__abc_43300_n218_bF_buf4;
  wire u0_u0__abc_43300_n218_bF_buf5;
  wire u0_u0__abc_43300_n218_bF_buf6;
  wire u0_u0__abc_43300_n218_bF_buf7;
  wire u0_u0__abc_43300_n219_1;
  wire u0_u0__abc_43300_n219_1_bF_buf0;
  wire u0_u0__abc_43300_n219_1_bF_buf1;
  wire u0_u0__abc_43300_n219_1_bF_buf2;
  wire u0_u0__abc_43300_n219_1_bF_buf3;
  wire u0_u0__abc_43300_n219_1_bF_buf4;
  wire u0_u0__abc_43300_n220_1;
  wire u0_u0__abc_43300_n221;
  wire u0_u0__abc_43300_n223_1;
  wire u0_u0__abc_43300_n224;
  wire u0_u0__abc_43300_n225_1;
  wire u0_u0__abc_43300_n227;
  wire u0_u0__abc_43300_n228_1;
  wire u0_u0__abc_43300_n229_1;
  wire u0_u0__abc_43300_n231_1;
  wire u0_u0__abc_43300_n232_1;
  wire u0_u0__abc_43300_n233;
  wire u0_u0__abc_43300_n235_1;
  wire u0_u0__abc_43300_n236;
  wire u0_u0__abc_43300_n237_1;
  wire u0_u0__abc_43300_n239;
  wire u0_u0__abc_43300_n240_1;
  wire u0_u0__abc_43300_n241_1;
  wire u0_u0__abc_43300_n243_1;
  wire u0_u0__abc_43300_n244_1;
  wire u0_u0__abc_43300_n245;
  wire u0_u0__abc_43300_n247_1;
  wire u0_u0__abc_43300_n248;
  wire u0_u0__abc_43300_n249_1;
  wire u0_u0__abc_43300_n251;
  wire u0_u0__abc_43300_n252_1;
  wire u0_u0__abc_43300_n253_1;
  wire u0_u0__abc_43300_n255_1;
  wire u0_u0__abc_43300_n256;
  wire u0_u0__abc_43300_n257;
  wire u0_u0__abc_43300_n259;
  wire u0_u0__abc_43300_n260_1;
  wire u0_u0__abc_43300_n261;
  wire u0_u0__abc_43300_n263;
  wire u0_u0__abc_43300_n264;
  wire u0_u0__abc_43300_n265;
  wire u0_u0__abc_43300_n267;
  wire u0_u0__abc_43300_n268_1;
  wire u0_u0__abc_43300_n269;
  wire u0_u0__abc_43300_n271;
  wire u0_u0__abc_43300_n272;
  wire u0_u0__abc_43300_n273_1;
  wire u0_u0__abc_43300_n275_1;
  wire u0_u0__abc_43300_n276;
  wire u0_u0__abc_43300_n277_1;
  wire u0_u0__abc_43300_n279_1;
  wire u0_u0__abc_43300_n280;
  wire u0_u0__abc_43300_n281;
  wire u0_u0__abc_43300_n283_1;
  wire u0_u0__abc_43300_n284;
  wire u0_u0__abc_43300_n285_1;
  wire u0_u0__abc_43300_n287_1;
  wire u0_u0__abc_43300_n288;
  wire u0_u0__abc_43300_n289_1;
  wire u0_u0__abc_43300_n291;
  wire u0_u0__abc_43300_n292;
  wire u0_u0__abc_43300_n293;
  wire u0_u0__abc_43300_n295;
  wire u0_u0__abc_43300_n296_1;
  wire u0_u0__abc_43300_n297;
  wire u0_u0__abc_43300_n299;
  wire u0_u0__abc_43300_n300;
  wire u0_u0__abc_43300_n301;
  wire u0_u0__abc_43300_n303;
  wire u0_u0__abc_43300_n304;
  wire u0_u0__abc_43300_n305;
  wire u0_u0__abc_43300_n307;
  wire u0_u0__abc_43300_n308;
  wire u0_u0__abc_43300_n309;
  wire u0_u0__abc_43300_n311;
  wire u0_u0__abc_43300_n312_1;
  wire u0_u0__abc_43300_n313;
  wire u0_u0__abc_43300_n315_1;
  wire u0_u0__abc_43300_n316_1;
  wire u0_u0__abc_43300_n317_1;
  wire u0_u0__abc_43300_n319;
  wire u0_u0__abc_43300_n320;
  wire u0_u0__abc_43300_n321_1;
  wire u0_u0__abc_43300_n323_1;
  wire u0_u0__abc_43300_n324_1;
  wire u0_u0__abc_43300_n325;
  wire u0_u0__abc_43300_n325_1;
  wire u0_u0__abc_43300_n327;
  wire u0_u0__abc_43300_n328;
  wire u0_u0__abc_43300_n329;
  wire u0_u0__abc_43300_n331;
  wire u0_u0__abc_43300_n332;
  wire u0_u0__abc_43300_n333;
  wire u0_u0__abc_43300_n335;
  wire u0_u0__abc_43300_n336;
  wire u0_u0__abc_43300_n337;
  wire u0_u0__abc_43300_n339;
  wire u0_u0__abc_43300_n340;
  wire u0_u0__abc_43300_n341;
  wire u0_u0__abc_43300_n343;
  wire u0_u0__abc_43300_n344;
  wire u0_u0__abc_43300_n345;
  wire u0_u0__abc_43300_n347;
  wire u0_u0__abc_43300_n349;
  wire u0_u0__abc_43300_n350;
  wire u0_u0__abc_43300_n350_bF_buf0;
  wire u0_u0__abc_43300_n350_bF_buf1;
  wire u0_u0__abc_43300_n350_bF_buf2;
  wire u0_u0__abc_43300_n350_bF_buf3;
  wire u0_u0__abc_43300_n350_bF_buf4;
  wire u0_u0__abc_43300_n351;
  wire u0_u0__abc_43300_n352;
  wire u0_u0__abc_43300_n354;
  wire u0_u0__abc_43300_n355;
  wire u0_u0__abc_43300_n356;
  wire u0_u0__abc_43300_n358;
  wire u0_u0__abc_43300_n359;
  wire u0_u0__abc_43300_n360;
  wire u0_u0__abc_43300_n362;
  wire u0_u0__abc_43300_n363;
  wire u0_u0__abc_43300_n364;
  wire u0_u0__abc_43300_n366;
  wire u0_u0__abc_43300_n367;
  wire u0_u0__abc_43300_n368;
  wire u0_u0__abc_43300_n370;
  wire u0_u0__abc_43300_n371;
  wire u0_u0__abc_43300_n372;
  wire u0_u0__abc_43300_n374;
  wire u0_u0__abc_43300_n375;
  wire u0_u0__abc_43300_n376;
  wire u0_u0__abc_43300_n378;
  wire u0_u0__abc_43300_n379;
  wire u0_u0__abc_43300_n380;
  wire u0_u0__abc_43300_n382;
  wire u0_u0__abc_43300_n383;
  wire u0_u0__abc_43300_n384;
  wire u0_u0__abc_43300_n386;
  wire u0_u0__abc_43300_n387;
  wire u0_u0__abc_43300_n388;
  wire u0_u0__abc_43300_n390;
  wire u0_u0__abc_43300_n391;
  wire u0_u0__abc_43300_n392;
  wire u0_u0__abc_43300_n394;
  wire u0_u0__abc_43300_n395;
  wire u0_u0__abc_43300_n396;
  wire u0_u0__abc_43300_n398;
  wire u0_u0__abc_43300_n399;
  wire u0_u0__abc_43300_n400;
  wire u0_u0__abc_43300_n402;
  wire u0_u0__abc_43300_n403;
  wire u0_u0__abc_43300_n404;
  wire u0_u0__abc_43300_n406;
  wire u0_u0__abc_43300_n407;
  wire u0_u0__abc_43300_n408;
  wire u0_u0__abc_43300_n410;
  wire u0_u0__abc_43300_n411;
  wire u0_u0__abc_43300_n412;
  wire u0_u0__abc_43300_n414;
  wire u0_u0__abc_43300_n415;
  wire u0_u0__abc_43300_n416;
  wire u0_u0__abc_43300_n418;
  wire u0_u0__abc_43300_n419;
  wire u0_u0__abc_43300_n420;
  wire u0_u0__abc_43300_n422;
  wire u0_u0__abc_43300_n423;
  wire u0_u0__abc_43300_n424;
  wire u0_u0__abc_43300_n426;
  wire u0_u0__abc_43300_n427;
  wire u0_u0__abc_43300_n428;
  wire u0_u0__abc_43300_n430;
  wire u0_u0__abc_43300_n431;
  wire u0_u0__abc_43300_n432;
  wire u0_u0__abc_43300_n434;
  wire u0_u0__abc_43300_n435;
  wire u0_u0__abc_43300_n436;
  wire u0_u0__abc_43300_n438;
  wire u0_u0__abc_43300_n439;
  wire u0_u0__abc_43300_n440;
  wire u0_u0__abc_43300_n442;
  wire u0_u0__abc_43300_n443;
  wire u0_u0__abc_43300_n444;
  wire u0_u0__abc_43300_n446;
  wire u0_u0__abc_43300_n447;
  wire u0_u0__abc_43300_n448;
  wire u0_u0__abc_43300_n450;
  wire u0_u0__abc_43300_n451;
  wire u0_u0__abc_43300_n452;
  wire u0_u0__abc_43300_n454;
  wire u0_u0__abc_43300_n455;
  wire u0_u0__abc_43300_n456;
  wire u0_u0__abc_43300_n458;
  wire u0_u0__abc_43300_n459;
  wire u0_u0__abc_43300_n460;
  wire u0_u0__abc_43300_n462;
  wire u0_u0__abc_43300_n463;
  wire u0_u0__abc_43300_n464;
  wire u0_u0__abc_43300_n466;
  wire u0_u0__abc_43300_n467;
  wire u0_u0__abc_43300_n468;
  wire u0_u0__abc_43300_n470;
  wire u0_u0__abc_43300_n471;
  wire u0_u0__abc_43300_n472;
  wire u0_u0__abc_43300_n474;
  wire u0_u0__abc_43300_n475;
  wire u0_u0__abc_43300_n476;
  wire u0_u0__abc_43300_n478;
  wire u0_u0__abc_43300_n479;
  wire u0_u0__abc_43300_n480;
  wire u0_u0__abc_43300_n481;
  wire u0_u0__abc_43300_n482;
  wire u0_u0__abc_43300_n483;
  wire u0_u0__abc_43300_n484;
  wire u0_u0__abc_43300_n485;
  wire u0_u0__abc_43300_n486;
  wire u0_u0__abc_43300_n487;
  wire u0_u0__abc_43300_n488;
  wire u0_u0__abc_43300_n489;
  wire u0_u0__abc_43300_n490;
  wire u0_u0__abc_43300_n491;
  wire u0_u0__abc_43300_n492;
  wire u0_u0__abc_43300_n493;
  wire u0_u0__abc_43300_n494;
  wire u0_u0__abc_43300_n495;
  wire u0_u0__abc_43300_n496;
  wire u0_u0__abc_43300_n497;
  wire u0_u0__abc_43300_n498;
  wire u0_u0__abc_43300_n499;
  wire u0_u0__abc_43300_n500;
  wire u0_u0__abc_43300_n501;
  wire u0_u0__abc_43300_n502;
  wire u0_u0__abc_43300_n503;
  wire u0_u0__abc_43300_n504;
  wire u0_u0__abc_43300_n505;
  wire u0_u0__abc_43300_n506;
  wire u0_u0__abc_43300_n507;
  wire u0_u0__abc_43300_n508;
  wire u0_u0__abc_43300_n509;
  wire u0_u0__abc_43300_n510;
  wire u0_u0__abc_43300_n511;
  wire u0_u0__abc_43300_n512;
  wire u0_u0__abc_43300_n513;
  wire u0_u0__abc_43300_n514;
  wire u0_u0__abc_43300_n515;
  wire u0_u0__abc_43300_n516;
  wire u0_u0__abc_43300_n517;
  wire u0_u0__abc_43300_n518;
  wire u0_u0__abc_43300_n519;
  wire u0_u0__abc_43300_n520;
  wire u0_u0__abc_43300_n521;
  wire u0_u0__abc_43300_n522;
  wire u0_u0__abc_43300_n523;
  wire u0_u0__abc_43300_n524;
  wire u0_u0__abc_43300_n525;
  wire u0_u0__abc_43300_n526;
  wire u0_u0__abc_43300_n527;
  wire u0_u0__abc_43300_n528;
  wire u0_u0__abc_43300_n529;
  wire u0_u0__abc_43300_n530;
  wire u0_u0__abc_43300_n531;
  wire u0_u0__abc_43300_n532;
  wire u0_u0__abc_43300_n533;
  wire u0_u0__abc_43300_n534;
  wire u0_u0__abc_43300_n535;
  wire u0_u0__abc_43300_n536;
  wire u0_u0__abc_43300_n537;
  wire u0_u0__abc_43300_n538;
  wire u0_u0__abc_43300_n539;
  wire u0_u0__abc_43300_n540;
  wire u0_u0__abc_43300_n541;
  wire u0_u0__abc_43300_n542;
  wire u0_u0__abc_43300_n543;
  wire u0_u0__abc_43300_n544;
  wire u0_u0__abc_43300_n546;
  wire u0_u0__abc_43300_n549;
  wire u0_u0__abc_43300_n550;
  wire u0_u0__abc_43300_n551;
  wire u0_u0__abc_43300_n552;
  wire u0_u0__abc_43300_n553;
  wire u0_u0__abc_43300_n554;
  wire u0_u0_addr_r_2_;
  wire u0_u0_addr_r_3_;
  wire u0_u0_addr_r_4_;
  wire u0_u0_addr_r_5_;
  wire u0_u0_addr_r_6_;
  wire u0_u0_csc_0__FF_INPUT;
  wire u0_u0_csc_10__FF_INPUT;
  wire u0_u0_csc_11__FF_INPUT;
  wire u0_u0_csc_12__FF_INPUT;
  wire u0_u0_csc_13__FF_INPUT;
  wire u0_u0_csc_14__FF_INPUT;
  wire u0_u0_csc_15__FF_INPUT;
  wire u0_u0_csc_16__FF_INPUT;
  wire u0_u0_csc_17__FF_INPUT;
  wire u0_u0_csc_18__FF_INPUT;
  wire u0_u0_csc_19__FF_INPUT;
  wire u0_u0_csc_1__FF_INPUT;
  wire u0_u0_csc_20__FF_INPUT;
  wire u0_u0_csc_21__FF_INPUT;
  wire u0_u0_csc_22__FF_INPUT;
  wire u0_u0_csc_23__FF_INPUT;
  wire u0_u0_csc_24__FF_INPUT;
  wire u0_u0_csc_25__FF_INPUT;
  wire u0_u0_csc_26__FF_INPUT;
  wire u0_u0_csc_27__FF_INPUT;
  wire u0_u0_csc_28__FF_INPUT;
  wire u0_u0_csc_29__FF_INPUT;
  wire u0_u0_csc_2__FF_INPUT;
  wire u0_u0_csc_30__FF_INPUT;
  wire u0_u0_csc_31__FF_INPUT;
  wire u0_u0_csc_3__FF_INPUT;
  wire u0_u0_csc_4__FF_INPUT;
  wire u0_u0_csc_5__FF_INPUT;
  wire u0_u0_csc_6__FF_INPUT;
  wire u0_u0_csc_7__FF_INPUT;
  wire u0_u0_csc_8__FF_INPUT;
  wire u0_u0_csc_9__FF_INPUT;
  wire u0_u0_init_req_FF_INPUT;
  wire u0_u0_init_req_we;
  wire u0_u0_init_req_we_FF_INPUT;
  wire u0_u0_init_req_we_FF_INPUT_bF_buf0;
  wire u0_u0_init_req_we_FF_INPUT_bF_buf1;
  wire u0_u0_init_req_we_FF_INPUT_bF_buf2;
  wire u0_u0_init_req_we_FF_INPUT_bF_buf3;
  wire u0_u0_init_req_we_FF_INPUT_bF_buf4;
  wire u0_u0_inited;
  wire u0_u0_inited_FF_INPUT;
  wire u0_u0_lmr_req_FF_INPUT;
  wire u0_u0_lmr_req_we;
  wire u0_u0_lmr_req_we_FF_INPUT;
  wire u0_u0_lmr_req_we_FF_INPUT_bF_buf0;
  wire u0_u0_lmr_req_we_FF_INPUT_bF_buf1;
  wire u0_u0_lmr_req_we_FF_INPUT_bF_buf2;
  wire u0_u0_lmr_req_we_FF_INPUT_bF_buf3;
  wire u0_u0_lmr_req_we_FF_INPUT_bF_buf4;
  wire u0_u0_rst_r1;
  wire u0_u0_rst_r2;
  wire u0_u0_tms_0__FF_INPUT;
  wire u0_u0_tms_10__FF_INPUT;
  wire u0_u0_tms_11__FF_INPUT;
  wire u0_u0_tms_12__FF_INPUT;
  wire u0_u0_tms_13__FF_INPUT;
  wire u0_u0_tms_14__FF_INPUT;
  wire u0_u0_tms_15__FF_INPUT;
  wire u0_u0_tms_16__FF_INPUT;
  wire u0_u0_tms_17__FF_INPUT;
  wire u0_u0_tms_18__FF_INPUT;
  wire u0_u0_tms_19__FF_INPUT;
  wire u0_u0_tms_1__FF_INPUT;
  wire u0_u0_tms_20__FF_INPUT;
  wire u0_u0_tms_21__FF_INPUT;
  wire u0_u0_tms_22__FF_INPUT;
  wire u0_u0_tms_23__FF_INPUT;
  wire u0_u0_tms_24__FF_INPUT;
  wire u0_u0_tms_25__FF_INPUT;
  wire u0_u0_tms_26__FF_INPUT;
  wire u0_u0_tms_27__FF_INPUT;
  wire u0_u0_tms_28__FF_INPUT;
  wire u0_u0_tms_29__FF_INPUT;
  wire u0_u0_tms_2__FF_INPUT;
  wire u0_u0_tms_30__FF_INPUT;
  wire u0_u0_tms_31__FF_INPUT;
  wire u0_u0_tms_3__FF_INPUT;
  wire u0_u0_tms_4__FF_INPUT;
  wire u0_u0_tms_5__FF_INPUT;
  wire u0_u0_tms_6__FF_INPUT;
  wire u0_u0_tms_7__FF_INPUT;
  wire u0_u0_tms_8__FF_INPUT;
  wire u0_u0_tms_9__FF_INPUT;
  wire u0_u0_wp_err;
  wire u0_u1__abc_43657_n201_1;
  wire u0_u1__abc_43657_n202;
  wire u0_u1__abc_43657_n203_1;
  wire u0_u1__abc_43657_n204_1;
  wire u0_u1__abc_43657_n205;
  wire u0_u1__abc_43657_n206_1;
  wire u0_u1__abc_43657_n207_1;
  wire u0_u1__abc_43657_n208;
  wire u0_u1__abc_43657_n209_1;
  wire u0_u1__abc_43657_n211;
  wire u0_u1__abc_43657_n212_1;
  wire u0_u1__abc_43657_n213_1;
  wire u0_u1__abc_43657_n214;
  wire u0_u1__abc_43657_n215_1;
  wire u0_u1__abc_43657_n216_1;
  wire u0_u1__abc_43657_n218_1;
  wire u0_u1__abc_43657_n219_1;
  wire u0_u1__abc_43657_n219_1_bF_buf0;
  wire u0_u1__abc_43657_n219_1_bF_buf1;
  wire u0_u1__abc_43657_n219_1_bF_buf2;
  wire u0_u1__abc_43657_n219_1_bF_buf3;
  wire u0_u1__abc_43657_n219_1_bF_buf4;
  wire u0_u1__abc_43657_n219_1_bF_buf5;
  wire u0_u1__abc_43657_n219_1_bF_buf6;
  wire u0_u1__abc_43657_n219_1_bF_buf7;
  wire u0_u1__abc_43657_n220;
  wire u0_u1__abc_43657_n221_1;
  wire u0_u1__abc_43657_n222_1;
  wire u0_u1__abc_43657_n223;
  wire u0_u1__abc_43657_n225_1;
  wire u0_u1__abc_43657_n226;
  wire u0_u1__abc_43657_n227_1;
  wire u0_u1__abc_43657_n228_1;
  wire u0_u1__abc_43657_n229;
  wire u0_u1__abc_43657_n231_1;
  wire u0_u1__abc_43657_n232;
  wire u0_u1__abc_43657_n233_1;
  wire u0_u1__abc_43657_n234_1;
  wire u0_u1__abc_43657_n235;
  wire u0_u1__abc_43657_n237_1;
  wire u0_u1__abc_43657_n238;
  wire u0_u1__abc_43657_n239_1;
  wire u0_u1__abc_43657_n240_1;
  wire u0_u1__abc_43657_n241;
  wire u0_u1__abc_43657_n243_1;
  wire u0_u1__abc_43657_n244;
  wire u0_u1__abc_43657_n245_1;
  wire u0_u1__abc_43657_n246_1;
  wire u0_u1__abc_43657_n247;
  wire u0_u1__abc_43657_n249_1;
  wire u0_u1__abc_43657_n250;
  wire u0_u1__abc_43657_n251_1;
  wire u0_u1__abc_43657_n252_1;
  wire u0_u1__abc_43657_n253;
  wire u0_u1__abc_43657_n255;
  wire u0_u1__abc_43657_n256;
  wire u0_u1__abc_43657_n257;
  wire u0_u1__abc_43657_n258;
  wire u0_u1__abc_43657_n259_1;
  wire u0_u1__abc_43657_n261_1;
  wire u0_u1__abc_43657_n262;
  wire u0_u1__abc_43657_n263;
  wire u0_u1__abc_43657_n264;
  wire u0_u1__abc_43657_n265_1;
  wire u0_u1__abc_43657_n267_1;
  wire u0_u1__abc_43657_n268;
  wire u0_u1__abc_43657_n269;
  wire u0_u1__abc_43657_n270;
  wire u0_u1__abc_43657_n271;
  wire u0_u1__abc_43657_n273;
  wire u0_u1__abc_43657_n274_1;
  wire u0_u1__abc_43657_n275;
  wire u0_u1__abc_43657_n276_1;
  wire u0_u1__abc_43657_n277;
  wire u0_u1__abc_43657_n279;
  wire u0_u1__abc_43657_n280;
  wire u0_u1__abc_43657_n281;
  wire u0_u1__abc_43657_n282_1;
  wire u0_u1__abc_43657_n283;
  wire u0_u1__abc_43657_n285;
  wire u0_u1__abc_43657_n286_1;
  wire u0_u1__abc_43657_n287;
  wire u0_u1__abc_43657_n288_1;
  wire u0_u1__abc_43657_n289;
  wire u0_u1__abc_43657_n291;
  wire u0_u1__abc_43657_n292;
  wire u0_u1__abc_43657_n293;
  wire u0_u1__abc_43657_n294;
  wire u0_u1__abc_43657_n295_1;
  wire u0_u1__abc_43657_n297_1;
  wire u0_u1__abc_43657_n298;
  wire u0_u1__abc_43657_n299;
  wire u0_u1__abc_43657_n300;
  wire u0_u1__abc_43657_n301;
  wire u0_u1__abc_43657_n303;
  wire u0_u1__abc_43657_n304;
  wire u0_u1__abc_43657_n305;
  wire u0_u1__abc_43657_n306;
  wire u0_u1__abc_43657_n307;
  wire u0_u1__abc_43657_n309_1;
  wire u0_u1__abc_43657_n310;
  wire u0_u1__abc_43657_n311_1;
  wire u0_u1__abc_43657_n312;
  wire u0_u1__abc_43657_n313_1;
  wire u0_u1__abc_43657_n315_1;
  wire u0_u1__abc_43657_n316_1;
  wire u0_u1__abc_43657_n317;
  wire u0_u1__abc_43657_n318;
  wire u0_u1__abc_43657_n319;
  wire u0_u1__abc_43657_n321;
  wire u0_u1__abc_43657_n322_1;
  wire u0_u1__abc_43657_n323_1;
  wire u0_u1__abc_43657_n324;
  wire u0_u1__abc_43657_n324_1;
  wire u0_u1__abc_43657_n325;
  wire u0_u1__abc_43657_n327;
  wire u0_u1__abc_43657_n328;
  wire u0_u1__abc_43657_n329;
  wire u0_u1__abc_43657_n330;
  wire u0_u1__abc_43657_n331;
  wire u0_u1__abc_43657_n333;
  wire u0_u1__abc_43657_n334;
  wire u0_u1__abc_43657_n335;
  wire u0_u1__abc_43657_n336;
  wire u0_u1__abc_43657_n337;
  wire u0_u1__abc_43657_n339;
  wire u0_u1__abc_43657_n340;
  wire u0_u1__abc_43657_n341;
  wire u0_u1__abc_43657_n342;
  wire u0_u1__abc_43657_n343;
  wire u0_u1__abc_43657_n345;
  wire u0_u1__abc_43657_n346;
  wire u0_u1__abc_43657_n347;
  wire u0_u1__abc_43657_n348;
  wire u0_u1__abc_43657_n349;
  wire u0_u1__abc_43657_n351;
  wire u0_u1__abc_43657_n352;
  wire u0_u1__abc_43657_n353;
  wire u0_u1__abc_43657_n354;
  wire u0_u1__abc_43657_n355;
  wire u0_u1__abc_43657_n357;
  wire u0_u1__abc_43657_n358;
  wire u0_u1__abc_43657_n359;
  wire u0_u1__abc_43657_n360;
  wire u0_u1__abc_43657_n361;
  wire u0_u1__abc_43657_n363;
  wire u0_u1__abc_43657_n364;
  wire u0_u1__abc_43657_n365;
  wire u0_u1__abc_43657_n366;
  wire u0_u1__abc_43657_n367;
  wire u0_u1__abc_43657_n369;
  wire u0_u1__abc_43657_n370;
  wire u0_u1__abc_43657_n371;
  wire u0_u1__abc_43657_n372;
  wire u0_u1__abc_43657_n373;
  wire u0_u1__abc_43657_n375;
  wire u0_u1__abc_43657_n376;
  wire u0_u1__abc_43657_n377;
  wire u0_u1__abc_43657_n378;
  wire u0_u1__abc_43657_n379;
  wire u0_u1__abc_43657_n381;
  wire u0_u1__abc_43657_n382;
  wire u0_u1__abc_43657_n383;
  wire u0_u1__abc_43657_n384;
  wire u0_u1__abc_43657_n385;
  wire u0_u1__abc_43657_n387;
  wire u0_u1__abc_43657_n388;
  wire u0_u1__abc_43657_n389;
  wire u0_u1__abc_43657_n390;
  wire u0_u1__abc_43657_n391;
  wire u0_u1__abc_43657_n393;
  wire u0_u1__abc_43657_n394;
  wire u0_u1__abc_43657_n395;
  wire u0_u1__abc_43657_n396;
  wire u0_u1__abc_43657_n397;
  wire u0_u1__abc_43657_n399;
  wire u0_u1__abc_43657_n400;
  wire u0_u1__abc_43657_n401;
  wire u0_u1__abc_43657_n402;
  wire u0_u1__abc_43657_n403;
  wire u0_u1__abc_43657_n405;
  wire u0_u1__abc_43657_n406;
  wire u0_u1__abc_43657_n407;
  wire u0_u1__abc_43657_n408;
  wire u0_u1__abc_43657_n409;
  wire u0_u1__abc_43657_n411;
  wire u0_u1__abc_43657_n413;
  wire u0_u1__abc_43657_n414;
  wire u0_u1__abc_43657_n415;
  wire u0_u1__abc_43657_n416;
  wire u0_u1__abc_43657_n418;
  wire u0_u1__abc_43657_n419;
  wire u0_u1__abc_43657_n420;
  wire u0_u1__abc_43657_n421;
  wire u0_u1__abc_43657_n423;
  wire u0_u1__abc_43657_n424;
  wire u0_u1__abc_43657_n425;
  wire u0_u1__abc_43657_n426;
  wire u0_u1__abc_43657_n428;
  wire u0_u1__abc_43657_n429;
  wire u0_u1__abc_43657_n430;
  wire u0_u1__abc_43657_n431;
  wire u0_u1__abc_43657_n433;
  wire u0_u1__abc_43657_n434;
  wire u0_u1__abc_43657_n435;
  wire u0_u1__abc_43657_n436;
  wire u0_u1__abc_43657_n438;
  wire u0_u1__abc_43657_n439;
  wire u0_u1__abc_43657_n440;
  wire u0_u1__abc_43657_n441;
  wire u0_u1__abc_43657_n443;
  wire u0_u1__abc_43657_n444;
  wire u0_u1__abc_43657_n445;
  wire u0_u1__abc_43657_n446;
  wire u0_u1__abc_43657_n448;
  wire u0_u1__abc_43657_n449;
  wire u0_u1__abc_43657_n450;
  wire u0_u1__abc_43657_n451;
  wire u0_u1__abc_43657_n453;
  wire u0_u1__abc_43657_n454;
  wire u0_u1__abc_43657_n455;
  wire u0_u1__abc_43657_n456;
  wire u0_u1__abc_43657_n458;
  wire u0_u1__abc_43657_n459;
  wire u0_u1__abc_43657_n460;
  wire u0_u1__abc_43657_n461;
  wire u0_u1__abc_43657_n463;
  wire u0_u1__abc_43657_n464;
  wire u0_u1__abc_43657_n465;
  wire u0_u1__abc_43657_n466;
  wire u0_u1__abc_43657_n468;
  wire u0_u1__abc_43657_n469;
  wire u0_u1__abc_43657_n470;
  wire u0_u1__abc_43657_n471;
  wire u0_u1__abc_43657_n473;
  wire u0_u1__abc_43657_n474;
  wire u0_u1__abc_43657_n475;
  wire u0_u1__abc_43657_n476;
  wire u0_u1__abc_43657_n478;
  wire u0_u1__abc_43657_n479;
  wire u0_u1__abc_43657_n480;
  wire u0_u1__abc_43657_n481;
  wire u0_u1__abc_43657_n483;
  wire u0_u1__abc_43657_n484;
  wire u0_u1__abc_43657_n485;
  wire u0_u1__abc_43657_n486;
  wire u0_u1__abc_43657_n488;
  wire u0_u1__abc_43657_n489;
  wire u0_u1__abc_43657_n490;
  wire u0_u1__abc_43657_n491;
  wire u0_u1__abc_43657_n493;
  wire u0_u1__abc_43657_n494;
  wire u0_u1__abc_43657_n495;
  wire u0_u1__abc_43657_n496;
  wire u0_u1__abc_43657_n498;
  wire u0_u1__abc_43657_n499;
  wire u0_u1__abc_43657_n500;
  wire u0_u1__abc_43657_n501;
  wire u0_u1__abc_43657_n503;
  wire u0_u1__abc_43657_n504;
  wire u0_u1__abc_43657_n505;
  wire u0_u1__abc_43657_n506;
  wire u0_u1__abc_43657_n508;
  wire u0_u1__abc_43657_n509;
  wire u0_u1__abc_43657_n510;
  wire u0_u1__abc_43657_n511;
  wire u0_u1__abc_43657_n513;
  wire u0_u1__abc_43657_n514;
  wire u0_u1__abc_43657_n515;
  wire u0_u1__abc_43657_n516;
  wire u0_u1__abc_43657_n518;
  wire u0_u1__abc_43657_n519;
  wire u0_u1__abc_43657_n520;
  wire u0_u1__abc_43657_n521;
  wire u0_u1__abc_43657_n523;
  wire u0_u1__abc_43657_n524;
  wire u0_u1__abc_43657_n525;
  wire u0_u1__abc_43657_n526;
  wire u0_u1__abc_43657_n528;
  wire u0_u1__abc_43657_n529;
  wire u0_u1__abc_43657_n530;
  wire u0_u1__abc_43657_n531;
  wire u0_u1__abc_43657_n533;
  wire u0_u1__abc_43657_n534;
  wire u0_u1__abc_43657_n535;
  wire u0_u1__abc_43657_n536;
  wire u0_u1__abc_43657_n538;
  wire u0_u1__abc_43657_n539;
  wire u0_u1__abc_43657_n540;
  wire u0_u1__abc_43657_n541;
  wire u0_u1__abc_43657_n543;
  wire u0_u1__abc_43657_n544;
  wire u0_u1__abc_43657_n545;
  wire u0_u1__abc_43657_n546;
  wire u0_u1__abc_43657_n548;
  wire u0_u1__abc_43657_n549;
  wire u0_u1__abc_43657_n550;
  wire u0_u1__abc_43657_n551;
  wire u0_u1__abc_43657_n553;
  wire u0_u1__abc_43657_n554;
  wire u0_u1__abc_43657_n555;
  wire u0_u1__abc_43657_n556;
  wire u0_u1__abc_43657_n558;
  wire u0_u1__abc_43657_n559;
  wire u0_u1__abc_43657_n560;
  wire u0_u1__abc_43657_n561;
  wire u0_u1__abc_43657_n563;
  wire u0_u1__abc_43657_n564;
  wire u0_u1__abc_43657_n565;
  wire u0_u1__abc_43657_n566;
  wire u0_u1__abc_43657_n568;
  wire u0_u1__abc_43657_n569;
  wire u0_u1__abc_43657_n570;
  wire u0_u1__abc_43657_n571;
  wire u0_u1__abc_43657_n573;
  wire u0_u1__abc_43657_n574;
  wire u0_u1__abc_43657_n575;
  wire u0_u1__abc_43657_n576;
  wire u0_u1__abc_43657_n577;
  wire u0_u1__abc_43657_n578;
  wire u0_u1__abc_43657_n579;
  wire u0_u1__abc_43657_n580;
  wire u0_u1__abc_43657_n581;
  wire u0_u1__abc_43657_n582;
  wire u0_u1__abc_43657_n583;
  wire u0_u1__abc_43657_n584;
  wire u0_u1__abc_43657_n585;
  wire u0_u1__abc_43657_n586;
  wire u0_u1__abc_43657_n587;
  wire u0_u1__abc_43657_n588;
  wire u0_u1__abc_43657_n589;
  wire u0_u1__abc_43657_n590;
  wire u0_u1__abc_43657_n591;
  wire u0_u1__abc_43657_n592;
  wire u0_u1__abc_43657_n593;
  wire u0_u1__abc_43657_n594;
  wire u0_u1__abc_43657_n595;
  wire u0_u1__abc_43657_n596;
  wire u0_u1__abc_43657_n597;
  wire u0_u1__abc_43657_n598;
  wire u0_u1__abc_43657_n599;
  wire u0_u1__abc_43657_n600;
  wire u0_u1__abc_43657_n601;
  wire u0_u1__abc_43657_n602;
  wire u0_u1__abc_43657_n603;
  wire u0_u1__abc_43657_n604;
  wire u0_u1__abc_43657_n605;
  wire u0_u1__abc_43657_n606;
  wire u0_u1__abc_43657_n607;
  wire u0_u1__abc_43657_n608;
  wire u0_u1__abc_43657_n609;
  wire u0_u1__abc_43657_n610;
  wire u0_u1__abc_43657_n611;
  wire u0_u1__abc_43657_n612;
  wire u0_u1__abc_43657_n613;
  wire u0_u1__abc_43657_n614;
  wire u0_u1__abc_43657_n615;
  wire u0_u1__abc_43657_n616;
  wire u0_u1__abc_43657_n617;
  wire u0_u1__abc_43657_n618;
  wire u0_u1__abc_43657_n619;
  wire u0_u1__abc_43657_n620;
  wire u0_u1__abc_43657_n621;
  wire u0_u1__abc_43657_n622;
  wire u0_u1__abc_43657_n623;
  wire u0_u1__abc_43657_n624;
  wire u0_u1__abc_43657_n625;
  wire u0_u1__abc_43657_n626;
  wire u0_u1__abc_43657_n627;
  wire u0_u1__abc_43657_n628;
  wire u0_u1__abc_43657_n629;
  wire u0_u1__abc_43657_n630;
  wire u0_u1__abc_43657_n631;
  wire u0_u1__abc_43657_n632;
  wire u0_u1__abc_43657_n633;
  wire u0_u1__abc_43657_n634;
  wire u0_u1__abc_43657_n635;
  wire u0_u1__abc_43657_n636;
  wire u0_u1__abc_43657_n637;
  wire u0_u1__abc_43657_n638;
  wire u0_u1__abc_43657_n639;
  wire u0_u1__abc_43657_n641;
  wire u0_u1__abc_43657_n644;
  wire u0_u1__abc_43657_n645;
  wire u0_u1__abc_43657_n646;
  wire u0_u1__abc_43657_n647;
  wire u0_u1__abc_43657_n648;
  wire u0_u1__abc_43657_n649;
  wire u0_u1_addr_r_2_;
  wire u0_u1_addr_r_3_;
  wire u0_u1_addr_r_4_;
  wire u0_u1_addr_r_5_;
  wire u0_u1_addr_r_6_;
  wire u0_u1_csc_0__FF_INPUT;
  wire u0_u1_csc_10__FF_INPUT;
  wire u0_u1_csc_11__FF_INPUT;
  wire u0_u1_csc_12__FF_INPUT;
  wire u0_u1_csc_13__FF_INPUT;
  wire u0_u1_csc_14__FF_INPUT;
  wire u0_u1_csc_15__FF_INPUT;
  wire u0_u1_csc_16__FF_INPUT;
  wire u0_u1_csc_17__FF_INPUT;
  wire u0_u1_csc_18__FF_INPUT;
  wire u0_u1_csc_19__FF_INPUT;
  wire u0_u1_csc_1__FF_INPUT;
  wire u0_u1_csc_20__FF_INPUT;
  wire u0_u1_csc_21__FF_INPUT;
  wire u0_u1_csc_22__FF_INPUT;
  wire u0_u1_csc_23__FF_INPUT;
  wire u0_u1_csc_24__FF_INPUT;
  wire u0_u1_csc_25__FF_INPUT;
  wire u0_u1_csc_26__FF_INPUT;
  wire u0_u1_csc_27__FF_INPUT;
  wire u0_u1_csc_28__FF_INPUT;
  wire u0_u1_csc_29__FF_INPUT;
  wire u0_u1_csc_2__FF_INPUT;
  wire u0_u1_csc_30__FF_INPUT;
  wire u0_u1_csc_31__FF_INPUT;
  wire u0_u1_csc_3__FF_INPUT;
  wire u0_u1_csc_4__FF_INPUT;
  wire u0_u1_csc_5__FF_INPUT;
  wire u0_u1_csc_6__FF_INPUT;
  wire u0_u1_csc_7__FF_INPUT;
  wire u0_u1_csc_8__FF_INPUT;
  wire u0_u1_csc_9__FF_INPUT;
  wire u0_u1_init_req_FF_INPUT;
  wire u0_u1_init_req_we;
  wire u0_u1_init_req_we_FF_INPUT;
  wire u0_u1_init_req_we_FF_INPUT_bF_buf0;
  wire u0_u1_init_req_we_FF_INPUT_bF_buf1;
  wire u0_u1_init_req_we_FF_INPUT_bF_buf2;
  wire u0_u1_init_req_we_FF_INPUT_bF_buf3;
  wire u0_u1_init_req_we_FF_INPUT_bF_buf4;
  wire u0_u1_init_req_we_FF_INPUT_bF_buf5;
  wire u0_u1_init_req_we_FF_INPUT_bF_buf6;
  wire u0_u1_init_req_we_FF_INPUT_bF_buf7;
  wire u0_u1_inited;
  wire u0_u1_inited_FF_INPUT;
  wire u0_u1_lmr_req_FF_INPUT;
  wire u0_u1_lmr_req_we;
  wire u0_u1_lmr_req_we_FF_INPUT;
  wire u0_u1_lmr_req_we_FF_INPUT_bF_buf0;
  wire u0_u1_lmr_req_we_FF_INPUT_bF_buf1;
  wire u0_u1_lmr_req_we_FF_INPUT_bF_buf2;
  wire u0_u1_lmr_req_we_FF_INPUT_bF_buf3;
  wire u0_u1_lmr_req_we_FF_INPUT_bF_buf4;
  wire u0_u1_lmr_req_we_FF_INPUT_bF_buf5;
  wire u0_u1_lmr_req_we_FF_INPUT_bF_buf6;
  wire u0_u1_lmr_req_we_FF_INPUT_bF_buf7;
  wire u0_u1_rst_r1;
  wire u0_u1_rst_r2;
  wire u0_u1_tms_0__FF_INPUT;
  wire u0_u1_tms_10__FF_INPUT;
  wire u0_u1_tms_11__FF_INPUT;
  wire u0_u1_tms_12__FF_INPUT;
  wire u0_u1_tms_13__FF_INPUT;
  wire u0_u1_tms_14__FF_INPUT;
  wire u0_u1_tms_15__FF_INPUT;
  wire u0_u1_tms_16__FF_INPUT;
  wire u0_u1_tms_17__FF_INPUT;
  wire u0_u1_tms_18__FF_INPUT;
  wire u0_u1_tms_19__FF_INPUT;
  wire u0_u1_tms_1__FF_INPUT;
  wire u0_u1_tms_20__FF_INPUT;
  wire u0_u1_tms_21__FF_INPUT;
  wire u0_u1_tms_22__FF_INPUT;
  wire u0_u1_tms_23__FF_INPUT;
  wire u0_u1_tms_24__FF_INPUT;
  wire u0_u1_tms_25__FF_INPUT;
  wire u0_u1_tms_26__FF_INPUT;
  wire u0_u1_tms_27__FF_INPUT;
  wire u0_u1_tms_28__FF_INPUT;
  wire u0_u1_tms_29__FF_INPUT;
  wire u0_u1_tms_2__FF_INPUT;
  wire u0_u1_tms_30__FF_INPUT;
  wire u0_u1_tms_31__FF_INPUT;
  wire u0_u1_tms_3__FF_INPUT;
  wire u0_u1_tms_4__FF_INPUT;
  wire u0_u1_tms_5__FF_INPUT;
  wire u0_u1_tms_6__FF_INPUT;
  wire u0_u1_tms_7__FF_INPUT;
  wire u0_u1_tms_8__FF_INPUT;
  wire u0_u1_tms_9__FF_INPUT;
  wire u0_u1_wp_err;
  wire u0_u2__abc_44109_n201_1;
  wire u0_u2__abc_44109_n202_1;
  wire u0_u2__abc_44109_n203;
  wire u0_u2__abc_44109_n204_1;
  wire u0_u2__abc_44109_n205_1;
  wire u0_u2__abc_44109_n206;
  wire u0_u2__abc_44109_n208_1;
  wire u0_u2__abc_44109_n209;
  wire u0_u2__abc_44109_n209_bF_buf0;
  wire u0_u2__abc_44109_n209_bF_buf1;
  wire u0_u2__abc_44109_n209_bF_buf2;
  wire u0_u2__abc_44109_n209_bF_buf3;
  wire u0_u2__abc_44109_n209_bF_buf4;
  wire u0_u2__abc_44109_n209_bF_buf5;
  wire u0_u2__abc_44109_n209_bF_buf6;
  wire u0_u2__abc_44109_n209_bF_buf7;
  wire u0_u2__abc_44109_n210_1;
  wire u0_u2__abc_44109_n210_1_bF_buf0;
  wire u0_u2__abc_44109_n210_1_bF_buf1;
  wire u0_u2__abc_44109_n210_1_bF_buf2;
  wire u0_u2__abc_44109_n210_1_bF_buf3;
  wire u0_u2__abc_44109_n210_1_bF_buf4;
  wire u0_u2__abc_44109_n211_1;
  wire u0_u2__abc_44109_n212;
  wire u0_u2__abc_44109_n214_1;
  wire u0_u2__abc_44109_n215;
  wire u0_u2__abc_44109_n216_1;
  wire u0_u2__abc_44109_n218;
  wire u0_u2__abc_44109_n219_1;
  wire u0_u2__abc_44109_n220_1;
  wire u0_u2__abc_44109_n222_1;
  wire u0_u2__abc_44109_n223_1;
  wire u0_u2__abc_44109_n224;
  wire u0_u2__abc_44109_n226_1;
  wire u0_u2__abc_44109_n227;
  wire u0_u2__abc_44109_n228_1;
  wire u0_u2__abc_44109_n230;
  wire u0_u2__abc_44109_n231_1;
  wire u0_u2__abc_44109_n232_1;
  wire u0_u2__abc_44109_n234_1;
  wire u0_u2__abc_44109_n235_1;
  wire u0_u2__abc_44109_n236;
  wire u0_u2__abc_44109_n238_1;
  wire u0_u2__abc_44109_n239;
  wire u0_u2__abc_44109_n240_1;
  wire u0_u2__abc_44109_n242;
  wire u0_u2__abc_44109_n243;
  wire u0_u2__abc_44109_n244;
  wire u0_u2__abc_44109_n246_1;
  wire u0_u2__abc_44109_n247;
  wire u0_u2__abc_44109_n248_1;
  wire u0_u2__abc_44109_n250_1;
  wire u0_u2__abc_44109_n251_1;
  wire u0_u2__abc_44109_n252_1;
  wire u0_u2__abc_44109_n254;
  wire u0_u2__abc_44109_n255;
  wire u0_u2__abc_44109_n256_1;
  wire u0_u2__abc_44109_n258_1;
  wire u0_u2__abc_44109_n259_1;
  wire u0_u2__abc_44109_n260_1;
  wire u0_u2__abc_44109_n262;
  wire u0_u2__abc_44109_n263_1;
  wire u0_u2__abc_44109_n264;
  wire u0_u2__abc_44109_n266;
  wire u0_u2__abc_44109_n267;
  wire u0_u2__abc_44109_n268_1;
  wire u0_u2__abc_44109_n270_1;
  wire u0_u2__abc_44109_n271;
  wire u0_u2__abc_44109_n272;
  wire u0_u2__abc_44109_n274_1;
  wire u0_u2__abc_44109_n275;
  wire u0_u2__abc_44109_n276_1;
  wire u0_u2__abc_44109_n278;
  wire u0_u2__abc_44109_n279;
  wire u0_u2__abc_44109_n280;
  wire u0_u2__abc_44109_n282;
  wire u0_u2__abc_44109_n283_1;
  wire u0_u2__abc_44109_n284;
  wire u0_u2__abc_44109_n286;
  wire u0_u2__abc_44109_n287_1;
  wire u0_u2__abc_44109_n288;
  wire u0_u2__abc_44109_n290;
  wire u0_u2__abc_44109_n291_1;
  wire u0_u2__abc_44109_n292;
  wire u0_u2__abc_44109_n294;
  wire u0_u2__abc_44109_n295_1;
  wire u0_u2__abc_44109_n296;
  wire u0_u2__abc_44109_n298;
  wire u0_u2__abc_44109_n299;
  wire u0_u2__abc_44109_n300;
  wire u0_u2__abc_44109_n302;
  wire u0_u2__abc_44109_n303;
  wire u0_u2__abc_44109_n304_1;
  wire u0_u2__abc_44109_n306_1;
  wire u0_u2__abc_44109_n307;
  wire u0_u2__abc_44109_n308;
  wire u0_u2__abc_44109_n310;
  wire u0_u2__abc_44109_n311;
  wire u0_u2__abc_44109_n312;
  wire u0_u2__abc_44109_n314;
  wire u0_u2__abc_44109_n315;
  wire u0_u2__abc_44109_n316;
  wire u0_u2__abc_44109_n318_1;
  wire u0_u2__abc_44109_n319;
  wire u0_u2__abc_44109_n320_1;
  wire u0_u2__abc_44109_n322_1;
  wire u0_u2__abc_44109_n323_1;
  wire u0_u2__abc_44109_n324;
  wire u0_u2__abc_44109_n324_1;
  wire u0_u2__abc_44109_n326;
  wire u0_u2__abc_44109_n327;
  wire u0_u2__abc_44109_n328;
  wire u0_u2__abc_44109_n330;
  wire u0_u2__abc_44109_n331;
  wire u0_u2__abc_44109_n332;
  wire u0_u2__abc_44109_n334;
  wire u0_u2__abc_44109_n335;
  wire u0_u2__abc_44109_n336;
  wire u0_u2__abc_44109_n339;
  wire u0_u2__abc_44109_n340;
  wire u0_u2__abc_44109_n340_bF_buf0;
  wire u0_u2__abc_44109_n340_bF_buf1;
  wire u0_u2__abc_44109_n340_bF_buf2;
  wire u0_u2__abc_44109_n340_bF_buf3;
  wire u0_u2__abc_44109_n340_bF_buf4;
  wire u0_u2__abc_44109_n341;
  wire u0_u2__abc_44109_n342;
  wire u0_u2__abc_44109_n344;
  wire u0_u2__abc_44109_n345;
  wire u0_u2__abc_44109_n346;
  wire u0_u2__abc_44109_n348;
  wire u0_u2__abc_44109_n349;
  wire u0_u2__abc_44109_n350;
  wire u0_u2__abc_44109_n352;
  wire u0_u2__abc_44109_n353;
  wire u0_u2__abc_44109_n354;
  wire u0_u2__abc_44109_n356;
  wire u0_u2__abc_44109_n357;
  wire u0_u2__abc_44109_n358;
  wire u0_u2__abc_44109_n360;
  wire u0_u2__abc_44109_n361;
  wire u0_u2__abc_44109_n362;
  wire u0_u2__abc_44109_n364;
  wire u0_u2__abc_44109_n365;
  wire u0_u2__abc_44109_n366;
  wire u0_u2__abc_44109_n368;
  wire u0_u2__abc_44109_n369;
  wire u0_u2__abc_44109_n370;
  wire u0_u2__abc_44109_n372;
  wire u0_u2__abc_44109_n373;
  wire u0_u2__abc_44109_n374;
  wire u0_u2__abc_44109_n376;
  wire u0_u2__abc_44109_n377;
  wire u0_u2__abc_44109_n378;
  wire u0_u2__abc_44109_n380;
  wire u0_u2__abc_44109_n381;
  wire u0_u2__abc_44109_n382;
  wire u0_u2__abc_44109_n384;
  wire u0_u2__abc_44109_n385;
  wire u0_u2__abc_44109_n386;
  wire u0_u2__abc_44109_n388;
  wire u0_u2__abc_44109_n389;
  wire u0_u2__abc_44109_n390;
  wire u0_u2__abc_44109_n392;
  wire u0_u2__abc_44109_n393;
  wire u0_u2__abc_44109_n394;
  wire u0_u2__abc_44109_n396;
  wire u0_u2__abc_44109_n397;
  wire u0_u2__abc_44109_n398;
  wire u0_u2__abc_44109_n400;
  wire u0_u2__abc_44109_n401;
  wire u0_u2__abc_44109_n402;
  wire u0_u2__abc_44109_n404;
  wire u0_u2__abc_44109_n405;
  wire u0_u2__abc_44109_n406;
  wire u0_u2__abc_44109_n408;
  wire u0_u2__abc_44109_n409;
  wire u0_u2__abc_44109_n410;
  wire u0_u2__abc_44109_n412;
  wire u0_u2__abc_44109_n413;
  wire u0_u2__abc_44109_n414;
  wire u0_u2__abc_44109_n416;
  wire u0_u2__abc_44109_n417;
  wire u0_u2__abc_44109_n418;
  wire u0_u2__abc_44109_n420;
  wire u0_u2__abc_44109_n421;
  wire u0_u2__abc_44109_n422;
  wire u0_u2__abc_44109_n424;
  wire u0_u2__abc_44109_n425;
  wire u0_u2__abc_44109_n426;
  wire u0_u2__abc_44109_n428;
  wire u0_u2__abc_44109_n429;
  wire u0_u2__abc_44109_n430;
  wire u0_u2__abc_44109_n432;
  wire u0_u2__abc_44109_n433;
  wire u0_u2__abc_44109_n434;
  wire u0_u2__abc_44109_n436;
  wire u0_u2__abc_44109_n437;
  wire u0_u2__abc_44109_n438;
  wire u0_u2__abc_44109_n440;
  wire u0_u2__abc_44109_n441;
  wire u0_u2__abc_44109_n442;
  wire u0_u2__abc_44109_n444;
  wire u0_u2__abc_44109_n445;
  wire u0_u2__abc_44109_n446;
  wire u0_u2__abc_44109_n448;
  wire u0_u2__abc_44109_n449;
  wire u0_u2__abc_44109_n450;
  wire u0_u2__abc_44109_n452;
  wire u0_u2__abc_44109_n453;
  wire u0_u2__abc_44109_n454;
  wire u0_u2__abc_44109_n456;
  wire u0_u2__abc_44109_n457;
  wire u0_u2__abc_44109_n458;
  wire u0_u2__abc_44109_n460;
  wire u0_u2__abc_44109_n461;
  wire u0_u2__abc_44109_n462;
  wire u0_u2__abc_44109_n464;
  wire u0_u2__abc_44109_n465;
  wire u0_u2__abc_44109_n466;
  wire u0_u2__abc_44109_n468;
  wire u0_u2__abc_44109_n469;
  wire u0_u2__abc_44109_n470;
  wire u0_u2__abc_44109_n471;
  wire u0_u2__abc_44109_n472;
  wire u0_u2__abc_44109_n473;
  wire u0_u2__abc_44109_n474;
  wire u0_u2__abc_44109_n475;
  wire u0_u2__abc_44109_n476;
  wire u0_u2__abc_44109_n478;
  wire u0_u2__abc_44109_n479;
  wire u0_u2__abc_44109_n480;
  wire u0_u2__abc_44109_n481;
  wire u0_u2__abc_44109_n482;
  wire u0_u2__abc_44109_n483;
  wire u0_u2__abc_44109_n486;
  wire u0_u2__abc_44109_n487;
  wire u0_u2__abc_44109_n488;
  wire u0_u2__abc_44109_n489;
  wire u0_u2__abc_44109_n490;
  wire u0_u2__abc_44109_n491;
  wire u0_u2__abc_44109_n492;
  wire u0_u2__abc_44109_n493;
  wire u0_u2__abc_44109_n494;
  wire u0_u2__abc_44109_n495;
  wire u0_u2__abc_44109_n496;
  wire u0_u2__abc_44109_n497;
  wire u0_u2__abc_44109_n498;
  wire u0_u2__abc_44109_n499;
  wire u0_u2__abc_44109_n500;
  wire u0_u2__abc_44109_n501;
  wire u0_u2__abc_44109_n502;
  wire u0_u2__abc_44109_n503;
  wire u0_u2__abc_44109_n504;
  wire u0_u2__abc_44109_n505;
  wire u0_u2__abc_44109_n506;
  wire u0_u2__abc_44109_n507;
  wire u0_u2__abc_44109_n508;
  wire u0_u2__abc_44109_n509;
  wire u0_u2__abc_44109_n510;
  wire u0_u2__abc_44109_n511;
  wire u0_u2__abc_44109_n512;
  wire u0_u2__abc_44109_n513;
  wire u0_u2__abc_44109_n514;
  wire u0_u2__abc_44109_n515;
  wire u0_u2__abc_44109_n516;
  wire u0_u2__abc_44109_n517;
  wire u0_u2__abc_44109_n518;
  wire u0_u2__abc_44109_n519;
  wire u0_u2__abc_44109_n520;
  wire u0_u2__abc_44109_n521;
  wire u0_u2__abc_44109_n522;
  wire u0_u2__abc_44109_n523;
  wire u0_u2__abc_44109_n524;
  wire u0_u2__abc_44109_n525;
  wire u0_u2__abc_44109_n526;
  wire u0_u2__abc_44109_n527;
  wire u0_u2__abc_44109_n528;
  wire u0_u2__abc_44109_n529;
  wire u0_u2__abc_44109_n530;
  wire u0_u2__abc_44109_n531;
  wire u0_u2__abc_44109_n532;
  wire u0_u2__abc_44109_n533;
  wire u0_u2__abc_44109_n534;
  wire u0_u2__abc_44109_n535;
  wire u0_u2__abc_44109_n536;
  wire u0_u2__abc_44109_n537;
  wire u0_u2__abc_44109_n538;
  wire u0_u2__abc_44109_n539;
  wire u0_u2__abc_44109_n540;
  wire u0_u2__abc_44109_n541;
  wire u0_u2__abc_44109_n542;
  wire u0_u2__abc_44109_n543;
  wire u0_u2__abc_44109_n544;
  wire u0_u2__abc_44109_n545;
  wire u0_u2__abc_44109_n546;
  wire u0_u2__abc_44109_n547;
  wire u0_u2__abc_44109_n548;
  wire u0_u2__abc_44109_n549;
  wire u0_u2__abc_44109_n550;
  wire u0_u2__abc_44109_n551;
  wire u0_u2__abc_44109_n552;
  wire u0_u2__abc_44109_n554;
  wire u0_u2_addr_r_2_;
  wire u0_u2_addr_r_3_;
  wire u0_u2_addr_r_4_;
  wire u0_u2_addr_r_5_;
  wire u0_u2_addr_r_6_;
  wire u0_u2_csc_0__FF_INPUT;
  wire u0_u2_csc_10__FF_INPUT;
  wire u0_u2_csc_11__FF_INPUT;
  wire u0_u2_csc_12__FF_INPUT;
  wire u0_u2_csc_13__FF_INPUT;
  wire u0_u2_csc_14__FF_INPUT;
  wire u0_u2_csc_15__FF_INPUT;
  wire u0_u2_csc_16__FF_INPUT;
  wire u0_u2_csc_17__FF_INPUT;
  wire u0_u2_csc_18__FF_INPUT;
  wire u0_u2_csc_19__FF_INPUT;
  wire u0_u2_csc_1__FF_INPUT;
  wire u0_u2_csc_20__FF_INPUT;
  wire u0_u2_csc_21__FF_INPUT;
  wire u0_u2_csc_22__FF_INPUT;
  wire u0_u2_csc_23__FF_INPUT;
  wire u0_u2_csc_24__FF_INPUT;
  wire u0_u2_csc_25__FF_INPUT;
  wire u0_u2_csc_26__FF_INPUT;
  wire u0_u2_csc_27__FF_INPUT;
  wire u0_u2_csc_28__FF_INPUT;
  wire u0_u2_csc_29__FF_INPUT;
  wire u0_u2_csc_2__FF_INPUT;
  wire u0_u2_csc_30__FF_INPUT;
  wire u0_u2_csc_31__FF_INPUT;
  wire u0_u2_csc_3__FF_INPUT;
  wire u0_u2_csc_4__FF_INPUT;
  wire u0_u2_csc_5__FF_INPUT;
  wire u0_u2_csc_6__FF_INPUT;
  wire u0_u2_csc_7__FF_INPUT;
  wire u0_u2_csc_8__FF_INPUT;
  wire u0_u2_csc_9__FF_INPUT;
  wire u0_u2_init_req_FF_INPUT;
  wire u0_u2_init_req_we;
  wire u0_u2_init_req_we_FF_INPUT;
  wire u0_u2_init_req_we_FF_INPUT_bF_buf0;
  wire u0_u2_init_req_we_FF_INPUT_bF_buf1;
  wire u0_u2_init_req_we_FF_INPUT_bF_buf2;
  wire u0_u2_init_req_we_FF_INPUT_bF_buf3;
  wire u0_u2_init_req_we_FF_INPUT_bF_buf4;
  wire u0_u2_inited;
  wire u0_u2_inited_FF_INPUT;
  wire u0_u2_lmr_req_FF_INPUT;
  wire u0_u2_lmr_req_we;
  wire u0_u2_lmr_req_we_FF_INPUT;
  wire u0_u2_lmr_req_we_FF_INPUT_bF_buf0;
  wire u0_u2_lmr_req_we_FF_INPUT_bF_buf1;
  wire u0_u2_lmr_req_we_FF_INPUT_bF_buf2;
  wire u0_u2_lmr_req_we_FF_INPUT_bF_buf3;
  wire u0_u2_lmr_req_we_FF_INPUT_bF_buf4;
  wire u0_u2_rst_r1;
  wire u0_u2_rst_r2;
  wire u0_u2_tms_0__FF_INPUT;
  wire u0_u2_tms_10__FF_INPUT;
  wire u0_u2_tms_11__FF_INPUT;
  wire u0_u2_tms_12__FF_INPUT;
  wire u0_u2_tms_13__FF_INPUT;
  wire u0_u2_tms_14__FF_INPUT;
  wire u0_u2_tms_15__FF_INPUT;
  wire u0_u2_tms_16__FF_INPUT;
  wire u0_u2_tms_17__FF_INPUT;
  wire u0_u2_tms_18__FF_INPUT;
  wire u0_u2_tms_19__FF_INPUT;
  wire u0_u2_tms_1__FF_INPUT;
  wire u0_u2_tms_20__FF_INPUT;
  wire u0_u2_tms_21__FF_INPUT;
  wire u0_u2_tms_22__FF_INPUT;
  wire u0_u2_tms_23__FF_INPUT;
  wire u0_u2_tms_24__FF_INPUT;
  wire u0_u2_tms_25__FF_INPUT;
  wire u0_u2_tms_26__FF_INPUT;
  wire u0_u2_tms_27__FF_INPUT;
  wire u0_u2_tms_28__FF_INPUT;
  wire u0_u2_tms_29__FF_INPUT;
  wire u0_u2_tms_2__FF_INPUT;
  wire u0_u2_tms_30__FF_INPUT;
  wire u0_u2_tms_31__FF_INPUT;
  wire u0_u2_tms_3__FF_INPUT;
  wire u0_u2_tms_4__FF_INPUT;
  wire u0_u2_tms_5__FF_INPUT;
  wire u0_u2_tms_6__FF_INPUT;
  wire u0_u2_tms_7__FF_INPUT;
  wire u0_u2_tms_8__FF_INPUT;
  wire u0_u2_tms_9__FF_INPUT;
  wire u0_u2_wp_err;
  wire u0_u3__abc_44466_n205_1;
  wire u0_u3__abc_44466_n205_1_bF_buf0;
  wire u0_u3__abc_44466_n205_1_bF_buf1;
  wire u0_u3__abc_44466_n205_1_bF_buf2;
  wire u0_u3__abc_44466_n205_1_bF_buf3;
  wire u0_u3__abc_44466_n205_1_bF_buf4;
  wire u0_u3__abc_44466_n206_1;
  wire u0_u3__abc_44466_n207;
  wire u0_u3__abc_44466_n208_1;
  wire u0_u3__abc_44466_n209_1;
  wire u0_u3__abc_44466_n210;
  wire u0_u3__abc_44466_n211_1;
  wire u0_u3__abc_44466_n212_1;
  wire u0_u3__abc_44466_n214_1;
  wire u0_u3__abc_44466_n215_1;
  wire u0_u3__abc_44466_n216;
  wire u0_u3__abc_44466_n217_1;
  wire u0_u3__abc_44466_n218_1;
  wire u0_u3__abc_44466_n219;
  wire u0_u3__abc_44466_n220_1;
  wire u0_u3__abc_44466_n221_1;
  wire u0_u3__abc_44466_n222;
  wire u0_u3__abc_44466_n224_1;
  wire u0_u3__abc_44466_n225;
  wire u0_u3__abc_44466_n226_1;
  wire u0_u3__abc_44466_n227_1;
  wire u0_u3__abc_44466_n228;
  wire u0_u3__abc_44466_n229_1;
  wire u0_u3__abc_44466_n231;
  wire u0_u3__abc_44466_n232_1;
  wire u0_u3__abc_44466_n233_1;
  wire u0_u3__abc_44466_n234;
  wire u0_u3__abc_44466_n235_1;
  wire u0_u3__abc_44466_n236_1;
  wire u0_u3__abc_44466_n238_1;
  wire u0_u3__abc_44466_n239_1;
  wire u0_u3__abc_44466_n239_1_bF_buf0;
  wire u0_u3__abc_44466_n239_1_bF_buf1;
  wire u0_u3__abc_44466_n239_1_bF_buf2;
  wire u0_u3__abc_44466_n239_1_bF_buf3;
  wire u0_u3__abc_44466_n239_1_bF_buf4;
  wire u0_u3__abc_44466_n240;
  wire u0_u3__abc_44466_n241_1;
  wire u0_u3__abc_44466_n243;
  wire u0_u3__abc_44466_n244_1;
  wire u0_u3__abc_44466_n245_1;
  wire u0_u3__abc_44466_n246;
  wire u0_u3__abc_44466_n247;
  wire u0_u3__abc_44466_n248;
  wire u0_u3__abc_44466_n249;
  wire u0_u3__abc_44466_n251;
  wire u0_u3__abc_44466_n252_1;
  wire u0_u3__abc_44466_n253;
  wire u0_u3__abc_44466_n254_1;
  wire u0_u3__abc_44466_n255_1;
  wire u0_u3__abc_44466_n256_1;
  wire u0_u3__abc_44466_n257;
  wire u0_u3__abc_44466_n259;
  wire u0_u3__abc_44466_n260_1;
  wire u0_u3__abc_44466_n261;
  wire u0_u3__abc_44466_n263_1;
  wire u0_u3__abc_44466_n264_1;
  wire u0_u3__abc_44466_n265_1;
  wire u0_u3__abc_44466_n267_1;
  wire u0_u3__abc_44466_n268;
  wire u0_u3__abc_44466_n269;
  wire u0_u3__abc_44466_n271;
  wire u0_u3__abc_44466_n272_1;
  wire u0_u3__abc_44466_n273;
  wire u0_u3__abc_44466_n275;
  wire u0_u3__abc_44466_n276;
  wire u0_u3__abc_44466_n277;
  wire u0_u3__abc_44466_n279;
  wire u0_u3__abc_44466_n280_1;
  wire u0_u3__abc_44466_n281;
  wire u0_u3__abc_44466_n283;
  wire u0_u3__abc_44466_n284;
  wire u0_u3__abc_44466_n285_1;
  wire u0_u3__abc_44466_n287_1;
  wire u0_u3__abc_44466_n288;
  wire u0_u3__abc_44466_n289_1;
  wire u0_u3__abc_44466_n291_1;
  wire u0_u3__abc_44466_n292;
  wire u0_u3__abc_44466_n293;
  wire u0_u3__abc_44466_n295_1;
  wire u0_u3__abc_44466_n296;
  wire u0_u3__abc_44466_n297_1;
  wire u0_u3__abc_44466_n299_1;
  wire u0_u3__abc_44466_n300;
  wire u0_u3__abc_44466_n301_1;
  wire u0_u3__abc_44466_n303;
  wire u0_u3__abc_44466_n304;
  wire u0_u3__abc_44466_n305;
  wire u0_u3__abc_44466_n307;
  wire u0_u3__abc_44466_n308_1;
  wire u0_u3__abc_44466_n309;
  wire u0_u3__abc_44466_n311;
  wire u0_u3__abc_44466_n312;
  wire u0_u3__abc_44466_n313;
  wire u0_u3__abc_44466_n315;
  wire u0_u3__abc_44466_n316;
  wire u0_u3__abc_44466_n317;
  wire u0_u3__abc_44466_n319;
  wire u0_u3__abc_44466_n320;
  wire u0_u3__abc_44466_n321;
  wire u0_u3__abc_44466_n323;
  wire u0_u3__abc_44466_n324_1;
  wire u0_u3__abc_44466_n325;
  wire u0_u3__abc_44466_n327_1;
  wire u0_u3__abc_44466_n328;
  wire u0_u3__abc_44466_n328_1;
  wire u0_u3__abc_44466_n329;
  wire u0_u3__abc_44466_n331;
  wire u0_u3__abc_44466_n332;
  wire u0_u3__abc_44466_n333;
  wire u0_u3__abc_44466_n335;
  wire u0_u3__abc_44466_n336;
  wire u0_u3__abc_44466_n337;
  wire u0_u3__abc_44466_n339;
  wire u0_u3__abc_44466_n340;
  wire u0_u3__abc_44466_n341;
  wire u0_u3__abc_44466_n343;
  wire u0_u3__abc_44466_n344;
  wire u0_u3__abc_44466_n345;
  wire u0_u3__abc_44466_n347;
  wire u0_u3__abc_44466_n348;
  wire u0_u3__abc_44466_n349;
  wire u0_u3__abc_44466_n351;
  wire u0_u3__abc_44466_n352;
  wire u0_u3__abc_44466_n353;
  wire u0_u3__abc_44466_n355;
  wire u0_u3__abc_44466_n356;
  wire u0_u3__abc_44466_n357;
  wire u0_u3__abc_44466_n359;
  wire u0_u3__abc_44466_n360;
  wire u0_u3__abc_44466_n361;
  wire u0_u3__abc_44466_n364;
  wire u0_u3__abc_44466_n364_bF_buf0;
  wire u0_u3__abc_44466_n364_bF_buf1;
  wire u0_u3__abc_44466_n364_bF_buf2;
  wire u0_u3__abc_44466_n364_bF_buf3;
  wire u0_u3__abc_44466_n364_bF_buf4;
  wire u0_u3__abc_44466_n365;
  wire u0_u3__abc_44466_n366;
  wire u0_u3__abc_44466_n367;
  wire u0_u3__abc_44466_n369;
  wire u0_u3__abc_44466_n370;
  wire u0_u3__abc_44466_n371;
  wire u0_u3__abc_44466_n373;
  wire u0_u3__abc_44466_n374;
  wire u0_u3__abc_44466_n375;
  wire u0_u3__abc_44466_n377;
  wire u0_u3__abc_44466_n378;
  wire u0_u3__abc_44466_n379;
  wire u0_u3__abc_44466_n381;
  wire u0_u3__abc_44466_n382;
  wire u0_u3__abc_44466_n383;
  wire u0_u3__abc_44466_n385;
  wire u0_u3__abc_44466_n386;
  wire u0_u3__abc_44466_n387;
  wire u0_u3__abc_44466_n389;
  wire u0_u3__abc_44466_n390;
  wire u0_u3__abc_44466_n391;
  wire u0_u3__abc_44466_n393;
  wire u0_u3__abc_44466_n394;
  wire u0_u3__abc_44466_n395;
  wire u0_u3__abc_44466_n397;
  wire u0_u3__abc_44466_n398;
  wire u0_u3__abc_44466_n399;
  wire u0_u3__abc_44466_n401;
  wire u0_u3__abc_44466_n402;
  wire u0_u3__abc_44466_n403;
  wire u0_u3__abc_44466_n405;
  wire u0_u3__abc_44466_n406;
  wire u0_u3__abc_44466_n407;
  wire u0_u3__abc_44466_n409;
  wire u0_u3__abc_44466_n410;
  wire u0_u3__abc_44466_n411;
  wire u0_u3__abc_44466_n413;
  wire u0_u3__abc_44466_n414;
  wire u0_u3__abc_44466_n415;
  wire u0_u3__abc_44466_n417;
  wire u0_u3__abc_44466_n418;
  wire u0_u3__abc_44466_n419;
  wire u0_u3__abc_44466_n421;
  wire u0_u3__abc_44466_n422;
  wire u0_u3__abc_44466_n423;
  wire u0_u3__abc_44466_n425;
  wire u0_u3__abc_44466_n426;
  wire u0_u3__abc_44466_n427;
  wire u0_u3__abc_44466_n429;
  wire u0_u3__abc_44466_n430;
  wire u0_u3__abc_44466_n431;
  wire u0_u3__abc_44466_n433;
  wire u0_u3__abc_44466_n434;
  wire u0_u3__abc_44466_n435;
  wire u0_u3__abc_44466_n437;
  wire u0_u3__abc_44466_n438;
  wire u0_u3__abc_44466_n439;
  wire u0_u3__abc_44466_n441;
  wire u0_u3__abc_44466_n442;
  wire u0_u3__abc_44466_n443;
  wire u0_u3__abc_44466_n445;
  wire u0_u3__abc_44466_n446;
  wire u0_u3__abc_44466_n447;
  wire u0_u3__abc_44466_n449;
  wire u0_u3__abc_44466_n450;
  wire u0_u3__abc_44466_n451;
  wire u0_u3__abc_44466_n453;
  wire u0_u3__abc_44466_n454;
  wire u0_u3__abc_44466_n455;
  wire u0_u3__abc_44466_n457;
  wire u0_u3__abc_44466_n458;
  wire u0_u3__abc_44466_n459;
  wire u0_u3__abc_44466_n461;
  wire u0_u3__abc_44466_n462;
  wire u0_u3__abc_44466_n463;
  wire u0_u3__abc_44466_n465;
  wire u0_u3__abc_44466_n466;
  wire u0_u3__abc_44466_n467;
  wire u0_u3__abc_44466_n469;
  wire u0_u3__abc_44466_n470;
  wire u0_u3__abc_44466_n471;
  wire u0_u3__abc_44466_n473;
  wire u0_u3__abc_44466_n474;
  wire u0_u3__abc_44466_n475;
  wire u0_u3__abc_44466_n477;
  wire u0_u3__abc_44466_n478;
  wire u0_u3__abc_44466_n479;
  wire u0_u3__abc_44466_n481;
  wire u0_u3__abc_44466_n482;
  wire u0_u3__abc_44466_n483;
  wire u0_u3__abc_44466_n485;
  wire u0_u3__abc_44466_n486;
  wire u0_u3__abc_44466_n487;
  wire u0_u3__abc_44466_n489;
  wire u0_u3__abc_44466_n490;
  wire u0_u3__abc_44466_n491;
  wire u0_u3__abc_44466_n493;
  wire u0_u3__abc_44466_n494;
  wire u0_u3__abc_44466_n495;
  wire u0_u3__abc_44466_n496;
  wire u0_u3__abc_44466_n497;
  wire u0_u3__abc_44466_n498;
  wire u0_u3__abc_44466_n499;
  wire u0_u3__abc_44466_n500;
  wire u0_u3__abc_44466_n501;
  wire u0_u3__abc_44466_n503;
  wire u0_u3__abc_44466_n504;
  wire u0_u3__abc_44466_n505;
  wire u0_u3__abc_44466_n506;
  wire u0_u3__abc_44466_n507;
  wire u0_u3__abc_44466_n508;
  wire u0_u3__abc_44466_n511;
  wire u0_u3__abc_44466_n512;
  wire u0_u3__abc_44466_n513;
  wire u0_u3__abc_44466_n514;
  wire u0_u3__abc_44466_n515;
  wire u0_u3__abc_44466_n516;
  wire u0_u3__abc_44466_n517;
  wire u0_u3__abc_44466_n518;
  wire u0_u3__abc_44466_n519;
  wire u0_u3__abc_44466_n520;
  wire u0_u3__abc_44466_n521;
  wire u0_u3__abc_44466_n522;
  wire u0_u3__abc_44466_n523;
  wire u0_u3__abc_44466_n524;
  wire u0_u3__abc_44466_n525;
  wire u0_u3__abc_44466_n526;
  wire u0_u3__abc_44466_n527;
  wire u0_u3__abc_44466_n528;
  wire u0_u3__abc_44466_n529;
  wire u0_u3__abc_44466_n530;
  wire u0_u3__abc_44466_n531;
  wire u0_u3__abc_44466_n532;
  wire u0_u3__abc_44466_n533;
  wire u0_u3__abc_44466_n534;
  wire u0_u3__abc_44466_n535;
  wire u0_u3__abc_44466_n536;
  wire u0_u3__abc_44466_n537;
  wire u0_u3__abc_44466_n538;
  wire u0_u3__abc_44466_n539;
  wire u0_u3__abc_44466_n540;
  wire u0_u3__abc_44466_n541;
  wire u0_u3__abc_44466_n542;
  wire u0_u3__abc_44466_n543;
  wire u0_u3__abc_44466_n544;
  wire u0_u3__abc_44466_n545;
  wire u0_u3__abc_44466_n546;
  wire u0_u3__abc_44466_n547;
  wire u0_u3__abc_44466_n548;
  wire u0_u3__abc_44466_n549;
  wire u0_u3__abc_44466_n550;
  wire u0_u3__abc_44466_n551;
  wire u0_u3__abc_44466_n552;
  wire u0_u3__abc_44466_n553;
  wire u0_u3__abc_44466_n554;
  wire u0_u3__abc_44466_n555;
  wire u0_u3__abc_44466_n556;
  wire u0_u3__abc_44466_n557;
  wire u0_u3__abc_44466_n558;
  wire u0_u3__abc_44466_n559;
  wire u0_u3__abc_44466_n560;
  wire u0_u3__abc_44466_n561;
  wire u0_u3__abc_44466_n562;
  wire u0_u3__abc_44466_n563;
  wire u0_u3__abc_44466_n564;
  wire u0_u3__abc_44466_n565;
  wire u0_u3__abc_44466_n566;
  wire u0_u3__abc_44466_n567;
  wire u0_u3__abc_44466_n568;
  wire u0_u3__abc_44466_n569;
  wire u0_u3__abc_44466_n570;
  wire u0_u3__abc_44466_n571;
  wire u0_u3__abc_44466_n572;
  wire u0_u3__abc_44466_n573;
  wire u0_u3__abc_44466_n574;
  wire u0_u3__abc_44466_n575;
  wire u0_u3__abc_44466_n576;
  wire u0_u3__abc_44466_n577;
  wire u0_u3__abc_44466_n579;
  wire u0_u3_addr_r_2_;
  wire u0_u3_addr_r_3_;
  wire u0_u3_addr_r_4_;
  wire u0_u3_addr_r_5_;
  wire u0_u3_addr_r_6_;
  wire u0_u3_csc_0__FF_INPUT;
  wire u0_u3_csc_10__FF_INPUT;
  wire u0_u3_csc_11__FF_INPUT;
  wire u0_u3_csc_12__FF_INPUT;
  wire u0_u3_csc_13__FF_INPUT;
  wire u0_u3_csc_14__FF_INPUT;
  wire u0_u3_csc_15__FF_INPUT;
  wire u0_u3_csc_16__FF_INPUT;
  wire u0_u3_csc_17__FF_INPUT;
  wire u0_u3_csc_18__FF_INPUT;
  wire u0_u3_csc_19__FF_INPUT;
  wire u0_u3_csc_1__FF_INPUT;
  wire u0_u3_csc_20__FF_INPUT;
  wire u0_u3_csc_21__FF_INPUT;
  wire u0_u3_csc_22__FF_INPUT;
  wire u0_u3_csc_23__FF_INPUT;
  wire u0_u3_csc_24__FF_INPUT;
  wire u0_u3_csc_25__FF_INPUT;
  wire u0_u3_csc_26__FF_INPUT;
  wire u0_u3_csc_27__FF_INPUT;
  wire u0_u3_csc_28__FF_INPUT;
  wire u0_u3_csc_29__FF_INPUT;
  wire u0_u3_csc_2__FF_INPUT;
  wire u0_u3_csc_30__FF_INPUT;
  wire u0_u3_csc_31__FF_INPUT;
  wire u0_u3_csc_3__FF_INPUT;
  wire u0_u3_csc_4__FF_INPUT;
  wire u0_u3_csc_5__FF_INPUT;
  wire u0_u3_csc_6__FF_INPUT;
  wire u0_u3_csc_7__FF_INPUT;
  wire u0_u3_csc_8__FF_INPUT;
  wire u0_u3_csc_9__FF_INPUT;
  wire u0_u3_init_req_FF_INPUT;
  wire u0_u3_init_req_we;
  wire u0_u3_init_req_we_FF_INPUT;
  wire u0_u3_init_req_we_FF_INPUT_bF_buf0;
  wire u0_u3_init_req_we_FF_INPUT_bF_buf1;
  wire u0_u3_init_req_we_FF_INPUT_bF_buf2;
  wire u0_u3_init_req_we_FF_INPUT_bF_buf3;
  wire u0_u3_init_req_we_FF_INPUT_bF_buf4;
  wire u0_u3_init_req_we_FF_INPUT_bF_buf5;
  wire u0_u3_inited;
  wire u0_u3_inited_FF_INPUT;
  wire u0_u3_lmr_req_FF_INPUT;
  wire u0_u3_lmr_req_we;
  wire u0_u3_lmr_req_we_FF_INPUT;
  wire u0_u3_lmr_req_we_FF_INPUT_bF_buf0;
  wire u0_u3_lmr_req_we_FF_INPUT_bF_buf1;
  wire u0_u3_lmr_req_we_FF_INPUT_bF_buf2;
  wire u0_u3_lmr_req_we_FF_INPUT_bF_buf3;
  wire u0_u3_lmr_req_we_FF_INPUT_bF_buf4;
  wire u0_u3_rst_r1;
  wire u0_u3_rst_r2;
  wire u0_u3_rst_r2_bF_buf0;
  wire u0_u3_rst_r2_bF_buf1;
  wire u0_u3_rst_r2_bF_buf2;
  wire u0_u3_rst_r2_bF_buf3;
  wire u0_u3_rst_r2_bF_buf4;
  wire u0_u3_rst_r2_bF_buf5;
  wire u0_u3_tms_0__FF_INPUT;
  wire u0_u3_tms_10__FF_INPUT;
  wire u0_u3_tms_11__FF_INPUT;
  wire u0_u3_tms_12__FF_INPUT;
  wire u0_u3_tms_13__FF_INPUT;
  wire u0_u3_tms_14__FF_INPUT;
  wire u0_u3_tms_15__FF_INPUT;
  wire u0_u3_tms_16__FF_INPUT;
  wire u0_u3_tms_17__FF_INPUT;
  wire u0_u3_tms_18__FF_INPUT;
  wire u0_u3_tms_19__FF_INPUT;
  wire u0_u3_tms_1__FF_INPUT;
  wire u0_u3_tms_20__FF_INPUT;
  wire u0_u3_tms_21__FF_INPUT;
  wire u0_u3_tms_22__FF_INPUT;
  wire u0_u3_tms_23__FF_INPUT;
  wire u0_u3_tms_24__FF_INPUT;
  wire u0_u3_tms_25__FF_INPUT;
  wire u0_u3_tms_26__FF_INPUT;
  wire u0_u3_tms_27__FF_INPUT;
  wire u0_u3_tms_28__FF_INPUT;
  wire u0_u3_tms_29__FF_INPUT;
  wire u0_u3_tms_2__FF_INPUT;
  wire u0_u3_tms_30__FF_INPUT;
  wire u0_u3_tms_31__FF_INPUT;
  wire u0_u3_tms_3__FF_INPUT;
  wire u0_u3_tms_4__FF_INPUT;
  wire u0_u3_tms_5__FF_INPUT;
  wire u0_u3_tms_6__FF_INPUT;
  wire u0_u3_tms_7__FF_INPUT;
  wire u0_u3_tms_8__FF_INPUT;
  wire u0_u3_tms_9__FF_INPUT;
  wire u0_u3_wp_err;
  wire u0_u4__abc_44844_n201_1;
  wire u0_u4__abc_44844_n202;
  wire u0_u4__abc_44844_n203_1;
  wire u0_u4__abc_44844_n204_1;
  wire u0_u4__abc_44844_n205;
  wire u0_u4__abc_44844_n206_1;
  wire u0_u4__abc_44844_n208;
  wire u0_u4__abc_44844_n209_1;
  wire u0_u4__abc_44844_n209_1_bF_buf0;
  wire u0_u4__abc_44844_n209_1_bF_buf1;
  wire u0_u4__abc_44844_n209_1_bF_buf2;
  wire u0_u4__abc_44844_n209_1_bF_buf3;
  wire u0_u4__abc_44844_n209_1_bF_buf4;
  wire u0_u4__abc_44844_n209_1_bF_buf5;
  wire u0_u4__abc_44844_n209_1_bF_buf6;
  wire u0_u4__abc_44844_n209_1_bF_buf7;
  wire u0_u4__abc_44844_n210_1;
  wire u0_u4__abc_44844_n211;
  wire u0_u4__abc_44844_n212_1;
  wire u0_u4__abc_44844_n213_1;
  wire u0_u4__abc_44844_n215_1;
  wire u0_u4__abc_44844_n216_1;
  wire u0_u4__abc_44844_n217;
  wire u0_u4__abc_44844_n218_1;
  wire u0_u4__abc_44844_n219_1;
  wire u0_u4__abc_44844_n221_1;
  wire u0_u4__abc_44844_n222_1;
  wire u0_u4__abc_44844_n223;
  wire u0_u4__abc_44844_n224_1;
  wire u0_u4__abc_44844_n225_1;
  wire u0_u4__abc_44844_n227_1;
  wire u0_u4__abc_44844_n228_1;
  wire u0_u4__abc_44844_n229;
  wire u0_u4__abc_44844_n230_1;
  wire u0_u4__abc_44844_n231_1;
  wire u0_u4__abc_44844_n233_1;
  wire u0_u4__abc_44844_n234_1;
  wire u0_u4__abc_44844_n235;
  wire u0_u4__abc_44844_n236_1;
  wire u0_u4__abc_44844_n237_1;
  wire u0_u4__abc_44844_n239_1;
  wire u0_u4__abc_44844_n240_1;
  wire u0_u4__abc_44844_n241;
  wire u0_u4__abc_44844_n242_1;
  wire u0_u4__abc_44844_n243_1;
  wire u0_u4__abc_44844_n245_1;
  wire u0_u4__abc_44844_n246_1;
  wire u0_u4__abc_44844_n247;
  wire u0_u4__abc_44844_n248_1;
  wire u0_u4__abc_44844_n249_1;
  wire u0_u4__abc_44844_n251_1;
  wire u0_u4__abc_44844_n252_1;
  wire u0_u4__abc_44844_n253;
  wire u0_u4__abc_44844_n254;
  wire u0_u4__abc_44844_n255;
  wire u0_u4__abc_44844_n257;
  wire u0_u4__abc_44844_n258_1;
  wire u0_u4__abc_44844_n259_1;
  wire u0_u4__abc_44844_n260_1;
  wire u0_u4__abc_44844_n261_1;
  wire u0_u4__abc_44844_n263_1;
  wire u0_u4__abc_44844_n264;
  wire u0_u4__abc_44844_n265;
  wire u0_u4__abc_44844_n266;
  wire u0_u4__abc_44844_n267;
  wire u0_u4__abc_44844_n269;
  wire u0_u4__abc_44844_n270_1;
  wire u0_u4__abc_44844_n271;
  wire u0_u4__abc_44844_n272;
  wire u0_u4__abc_44844_n273;
  wire u0_u4__abc_44844_n275;
  wire u0_u4__abc_44844_n276_1;
  wire u0_u4__abc_44844_n277;
  wire u0_u4__abc_44844_n278;
  wire u0_u4__abc_44844_n279;
  wire u0_u4__abc_44844_n281_1;
  wire u0_u4__abc_44844_n282;
  wire u0_u4__abc_44844_n283_1;
  wire u0_u4__abc_44844_n284;
  wire u0_u4__abc_44844_n285_1;
  wire u0_u4__abc_44844_n287_1;
  wire u0_u4__abc_44844_n288;
  wire u0_u4__abc_44844_n289;
  wire u0_u4__abc_44844_n290;
  wire u0_u4__abc_44844_n291_1;
  wire u0_u4__abc_44844_n293_1;
  wire u0_u4__abc_44844_n294;
  wire u0_u4__abc_44844_n295_1;
  wire u0_u4__abc_44844_n296;
  wire u0_u4__abc_44844_n297_1;
  wire u0_u4__abc_44844_n299;
  wire u0_u4__abc_44844_n300;
  wire u0_u4__abc_44844_n301;
  wire u0_u4__abc_44844_n302;
  wire u0_u4__abc_44844_n303;
  wire u0_u4__abc_44844_n305;
  wire u0_u4__abc_44844_n306_1;
  wire u0_u4__abc_44844_n307;
  wire u0_u4__abc_44844_n308;
  wire u0_u4__abc_44844_n309;
  wire u0_u4__abc_44844_n311;
  wire u0_u4__abc_44844_n312;
  wire u0_u4__abc_44844_n313;
  wire u0_u4__abc_44844_n314;
  wire u0_u4__abc_44844_n315;
  wire u0_u4__abc_44844_n317;
  wire u0_u4__abc_44844_n318_1;
  wire u0_u4__abc_44844_n319;
  wire u0_u4__abc_44844_n320_1;
  wire u0_u4__abc_44844_n321;
  wire u0_u4__abc_44844_n323_1;
  wire u0_u4__abc_44844_n324;
  wire u0_u4__abc_44844_n324_1;
  wire u0_u4__abc_44844_n325;
  wire u0_u4__abc_44844_n326;
  wire u0_u4__abc_44844_n327;
  wire u0_u4__abc_44844_n329;
  wire u0_u4__abc_44844_n330;
  wire u0_u4__abc_44844_n331;
  wire u0_u4__abc_44844_n332;
  wire u0_u4__abc_44844_n333;
  wire u0_u4__abc_44844_n335;
  wire u0_u4__abc_44844_n336;
  wire u0_u4__abc_44844_n337;
  wire u0_u4__abc_44844_n338;
  wire u0_u4__abc_44844_n339;
  wire u0_u4__abc_44844_n341;
  wire u0_u4__abc_44844_n342;
  wire u0_u4__abc_44844_n343;
  wire u0_u4__abc_44844_n344;
  wire u0_u4__abc_44844_n345;
  wire u0_u4__abc_44844_n347;
  wire u0_u4__abc_44844_n348;
  wire u0_u4__abc_44844_n349;
  wire u0_u4__abc_44844_n350;
  wire u0_u4__abc_44844_n351;
  wire u0_u4__abc_44844_n353;
  wire u0_u4__abc_44844_n354;
  wire u0_u4__abc_44844_n355;
  wire u0_u4__abc_44844_n356;
  wire u0_u4__abc_44844_n357;
  wire u0_u4__abc_44844_n359;
  wire u0_u4__abc_44844_n360;
  wire u0_u4__abc_44844_n361;
  wire u0_u4__abc_44844_n362;
  wire u0_u4__abc_44844_n363;
  wire u0_u4__abc_44844_n365;
  wire u0_u4__abc_44844_n366;
  wire u0_u4__abc_44844_n367;
  wire u0_u4__abc_44844_n368;
  wire u0_u4__abc_44844_n369;
  wire u0_u4__abc_44844_n371;
  wire u0_u4__abc_44844_n372;
  wire u0_u4__abc_44844_n373;
  wire u0_u4__abc_44844_n374;
  wire u0_u4__abc_44844_n375;
  wire u0_u4__abc_44844_n377;
  wire u0_u4__abc_44844_n378;
  wire u0_u4__abc_44844_n379;
  wire u0_u4__abc_44844_n380;
  wire u0_u4__abc_44844_n381;
  wire u0_u4__abc_44844_n383;
  wire u0_u4__abc_44844_n384;
  wire u0_u4__abc_44844_n385;
  wire u0_u4__abc_44844_n386;
  wire u0_u4__abc_44844_n387;
  wire u0_u4__abc_44844_n389;
  wire u0_u4__abc_44844_n390;
  wire u0_u4__abc_44844_n391;
  wire u0_u4__abc_44844_n392;
  wire u0_u4__abc_44844_n393;
  wire u0_u4__abc_44844_n395;
  wire u0_u4__abc_44844_n396;
  wire u0_u4__abc_44844_n397;
  wire u0_u4__abc_44844_n398;
  wire u0_u4__abc_44844_n399;
  wire u0_u4__abc_44844_n401;
  wire u0_u4__abc_44844_n402;
  wire u0_u4__abc_44844_n403;
  wire u0_u4__abc_44844_n404;
  wire u0_u4__abc_44844_n405;
  wire u0_u4__abc_44844_n406;
  wire u0_u4__abc_44844_n407;
  wire u0_u4__abc_44844_n408;
  wire u0_u4__abc_44844_n409;
  wire u0_u4__abc_44844_n411;
  wire u0_u4__abc_44844_n413;
  wire u0_u4__abc_44844_n414;
  wire u0_u4__abc_44844_n415;
  wire u0_u4__abc_44844_n416;
  wire u0_u4__abc_44844_n418;
  wire u0_u4__abc_44844_n419;
  wire u0_u4__abc_44844_n420;
  wire u0_u4__abc_44844_n421;
  wire u0_u4__abc_44844_n423;
  wire u0_u4__abc_44844_n424;
  wire u0_u4__abc_44844_n425;
  wire u0_u4__abc_44844_n426;
  wire u0_u4__abc_44844_n428;
  wire u0_u4__abc_44844_n429;
  wire u0_u4__abc_44844_n430;
  wire u0_u4__abc_44844_n431;
  wire u0_u4__abc_44844_n433;
  wire u0_u4__abc_44844_n434;
  wire u0_u4__abc_44844_n435;
  wire u0_u4__abc_44844_n436;
  wire u0_u4__abc_44844_n438;
  wire u0_u4__abc_44844_n439;
  wire u0_u4__abc_44844_n440;
  wire u0_u4__abc_44844_n441;
  wire u0_u4__abc_44844_n443;
  wire u0_u4__abc_44844_n444;
  wire u0_u4__abc_44844_n445;
  wire u0_u4__abc_44844_n446;
  wire u0_u4__abc_44844_n448;
  wire u0_u4__abc_44844_n449;
  wire u0_u4__abc_44844_n450;
  wire u0_u4__abc_44844_n451;
  wire u0_u4__abc_44844_n453;
  wire u0_u4__abc_44844_n454;
  wire u0_u4__abc_44844_n455;
  wire u0_u4__abc_44844_n456;
  wire u0_u4__abc_44844_n458;
  wire u0_u4__abc_44844_n459;
  wire u0_u4__abc_44844_n460;
  wire u0_u4__abc_44844_n461;
  wire u0_u4__abc_44844_n463;
  wire u0_u4__abc_44844_n464;
  wire u0_u4__abc_44844_n465;
  wire u0_u4__abc_44844_n466;
  wire u0_u4__abc_44844_n468;
  wire u0_u4__abc_44844_n469;
  wire u0_u4__abc_44844_n470;
  wire u0_u4__abc_44844_n471;
  wire u0_u4__abc_44844_n473;
  wire u0_u4__abc_44844_n474;
  wire u0_u4__abc_44844_n475;
  wire u0_u4__abc_44844_n476;
  wire u0_u4__abc_44844_n478;
  wire u0_u4__abc_44844_n479;
  wire u0_u4__abc_44844_n480;
  wire u0_u4__abc_44844_n481;
  wire u0_u4__abc_44844_n483;
  wire u0_u4__abc_44844_n484;
  wire u0_u4__abc_44844_n485;
  wire u0_u4__abc_44844_n486;
  wire u0_u4__abc_44844_n488;
  wire u0_u4__abc_44844_n489;
  wire u0_u4__abc_44844_n490;
  wire u0_u4__abc_44844_n491;
  wire u0_u4__abc_44844_n493;
  wire u0_u4__abc_44844_n494;
  wire u0_u4__abc_44844_n495;
  wire u0_u4__abc_44844_n496;
  wire u0_u4__abc_44844_n498;
  wire u0_u4__abc_44844_n499;
  wire u0_u4__abc_44844_n500;
  wire u0_u4__abc_44844_n501;
  wire u0_u4__abc_44844_n503;
  wire u0_u4__abc_44844_n504;
  wire u0_u4__abc_44844_n505;
  wire u0_u4__abc_44844_n506;
  wire u0_u4__abc_44844_n508;
  wire u0_u4__abc_44844_n509;
  wire u0_u4__abc_44844_n510;
  wire u0_u4__abc_44844_n511;
  wire u0_u4__abc_44844_n513;
  wire u0_u4__abc_44844_n514;
  wire u0_u4__abc_44844_n515;
  wire u0_u4__abc_44844_n516;
  wire u0_u4__abc_44844_n518;
  wire u0_u4__abc_44844_n519;
  wire u0_u4__abc_44844_n520;
  wire u0_u4__abc_44844_n521;
  wire u0_u4__abc_44844_n523;
  wire u0_u4__abc_44844_n524;
  wire u0_u4__abc_44844_n525;
  wire u0_u4__abc_44844_n526;
  wire u0_u4__abc_44844_n528;
  wire u0_u4__abc_44844_n529;
  wire u0_u4__abc_44844_n530;
  wire u0_u4__abc_44844_n531;
  wire u0_u4__abc_44844_n533;
  wire u0_u4__abc_44844_n534;
  wire u0_u4__abc_44844_n535;
  wire u0_u4__abc_44844_n536;
  wire u0_u4__abc_44844_n538;
  wire u0_u4__abc_44844_n539;
  wire u0_u4__abc_44844_n540;
  wire u0_u4__abc_44844_n541;
  wire u0_u4__abc_44844_n543;
  wire u0_u4__abc_44844_n544;
  wire u0_u4__abc_44844_n545;
  wire u0_u4__abc_44844_n546;
  wire u0_u4__abc_44844_n548;
  wire u0_u4__abc_44844_n549;
  wire u0_u4__abc_44844_n550;
  wire u0_u4__abc_44844_n551;
  wire u0_u4__abc_44844_n553;
  wire u0_u4__abc_44844_n554;
  wire u0_u4__abc_44844_n555;
  wire u0_u4__abc_44844_n556;
  wire u0_u4__abc_44844_n558;
  wire u0_u4__abc_44844_n559;
  wire u0_u4__abc_44844_n560;
  wire u0_u4__abc_44844_n561;
  wire u0_u4__abc_44844_n563;
  wire u0_u4__abc_44844_n564;
  wire u0_u4__abc_44844_n565;
  wire u0_u4__abc_44844_n566;
  wire u0_u4__abc_44844_n568;
  wire u0_u4__abc_44844_n569;
  wire u0_u4__abc_44844_n570;
  wire u0_u4__abc_44844_n571;
  wire u0_u4__abc_44844_n573;
  wire u0_u4__abc_44844_n574;
  wire u0_u4__abc_44844_n575;
  wire u0_u4__abc_44844_n576;
  wire u0_u4__abc_44844_n577;
  wire u0_u4__abc_44844_n578;
  wire u0_u4__abc_44844_n581;
  wire u0_u4__abc_44844_n582;
  wire u0_u4__abc_44844_n583;
  wire u0_u4__abc_44844_n584;
  wire u0_u4__abc_44844_n585;
  wire u0_u4__abc_44844_n586;
  wire u0_u4__abc_44844_n587;
  wire u0_u4__abc_44844_n588;
  wire u0_u4__abc_44844_n589;
  wire u0_u4__abc_44844_n590;
  wire u0_u4__abc_44844_n591;
  wire u0_u4__abc_44844_n592;
  wire u0_u4__abc_44844_n593;
  wire u0_u4__abc_44844_n594;
  wire u0_u4__abc_44844_n595;
  wire u0_u4__abc_44844_n596;
  wire u0_u4__abc_44844_n597;
  wire u0_u4__abc_44844_n598;
  wire u0_u4__abc_44844_n599;
  wire u0_u4__abc_44844_n600;
  wire u0_u4__abc_44844_n601;
  wire u0_u4__abc_44844_n602;
  wire u0_u4__abc_44844_n603;
  wire u0_u4__abc_44844_n604;
  wire u0_u4__abc_44844_n605;
  wire u0_u4__abc_44844_n606;
  wire u0_u4__abc_44844_n607;
  wire u0_u4__abc_44844_n608;
  wire u0_u4__abc_44844_n609;
  wire u0_u4__abc_44844_n610;
  wire u0_u4__abc_44844_n611;
  wire u0_u4__abc_44844_n612;
  wire u0_u4__abc_44844_n613;
  wire u0_u4__abc_44844_n614;
  wire u0_u4__abc_44844_n615;
  wire u0_u4__abc_44844_n616;
  wire u0_u4__abc_44844_n617;
  wire u0_u4__abc_44844_n618;
  wire u0_u4__abc_44844_n619;
  wire u0_u4__abc_44844_n620;
  wire u0_u4__abc_44844_n621;
  wire u0_u4__abc_44844_n622;
  wire u0_u4__abc_44844_n623;
  wire u0_u4__abc_44844_n624;
  wire u0_u4__abc_44844_n625;
  wire u0_u4__abc_44844_n626;
  wire u0_u4__abc_44844_n627;
  wire u0_u4__abc_44844_n628;
  wire u0_u4__abc_44844_n629;
  wire u0_u4__abc_44844_n630;
  wire u0_u4__abc_44844_n631;
  wire u0_u4__abc_44844_n632;
  wire u0_u4__abc_44844_n633;
  wire u0_u4__abc_44844_n634;
  wire u0_u4__abc_44844_n635;
  wire u0_u4__abc_44844_n636;
  wire u0_u4__abc_44844_n637;
  wire u0_u4__abc_44844_n638;
  wire u0_u4__abc_44844_n639;
  wire u0_u4__abc_44844_n640;
  wire u0_u4__abc_44844_n641;
  wire u0_u4__abc_44844_n642;
  wire u0_u4__abc_44844_n643;
  wire u0_u4__abc_44844_n644;
  wire u0_u4__abc_44844_n645;
  wire u0_u4__abc_44844_n646;
  wire u0_u4__abc_44844_n647;
  wire u0_u4__abc_44844_n649;
  wire u0_u4_addr_r_2_;
  wire u0_u4_addr_r_3_;
  wire u0_u4_addr_r_4_;
  wire u0_u4_addr_r_5_;
  wire u0_u4_addr_r_6_;
  wire u0_u4_csc_0__FF_INPUT;
  wire u0_u4_csc_10__FF_INPUT;
  wire u0_u4_csc_11__FF_INPUT;
  wire u0_u4_csc_12__FF_INPUT;
  wire u0_u4_csc_13__FF_INPUT;
  wire u0_u4_csc_14__FF_INPUT;
  wire u0_u4_csc_15__FF_INPUT;
  wire u0_u4_csc_16__FF_INPUT;
  wire u0_u4_csc_17__FF_INPUT;
  wire u0_u4_csc_18__FF_INPUT;
  wire u0_u4_csc_19__FF_INPUT;
  wire u0_u4_csc_1__FF_INPUT;
  wire u0_u4_csc_20__FF_INPUT;
  wire u0_u4_csc_21__FF_INPUT;
  wire u0_u4_csc_22__FF_INPUT;
  wire u0_u4_csc_23__FF_INPUT;
  wire u0_u4_csc_24__FF_INPUT;
  wire u0_u4_csc_25__FF_INPUT;
  wire u0_u4_csc_26__FF_INPUT;
  wire u0_u4_csc_27__FF_INPUT;
  wire u0_u4_csc_28__FF_INPUT;
  wire u0_u4_csc_29__FF_INPUT;
  wire u0_u4_csc_2__FF_INPUT;
  wire u0_u4_csc_30__FF_INPUT;
  wire u0_u4_csc_31__FF_INPUT;
  wire u0_u4_csc_3__FF_INPUT;
  wire u0_u4_csc_4__FF_INPUT;
  wire u0_u4_csc_5__FF_INPUT;
  wire u0_u4_csc_6__FF_INPUT;
  wire u0_u4_csc_7__FF_INPUT;
  wire u0_u4_csc_8__FF_INPUT;
  wire u0_u4_csc_9__FF_INPUT;
  wire u0_u4_init_req_FF_INPUT;
  wire u0_u4_init_req_we;
  wire u0_u4_init_req_we_FF_INPUT;
  wire u0_u4_init_req_we_FF_INPUT_bF_buf0;
  wire u0_u4_init_req_we_FF_INPUT_bF_buf1;
  wire u0_u4_init_req_we_FF_INPUT_bF_buf2;
  wire u0_u4_init_req_we_FF_INPUT_bF_buf3;
  wire u0_u4_init_req_we_FF_INPUT_bF_buf4;
  wire u0_u4_init_req_we_FF_INPUT_bF_buf5;
  wire u0_u4_init_req_we_FF_INPUT_bF_buf6;
  wire u0_u4_init_req_we_FF_INPUT_bF_buf7;
  wire u0_u4_inited;
  wire u0_u4_inited_FF_INPUT;
  wire u0_u4_lmr_req_FF_INPUT;
  wire u0_u4_lmr_req_we;
  wire u0_u4_lmr_req_we_FF_INPUT;
  wire u0_u4_lmr_req_we_FF_INPUT_bF_buf0;
  wire u0_u4_lmr_req_we_FF_INPUT_bF_buf1;
  wire u0_u4_lmr_req_we_FF_INPUT_bF_buf2;
  wire u0_u4_lmr_req_we_FF_INPUT_bF_buf3;
  wire u0_u4_lmr_req_we_FF_INPUT_bF_buf4;
  wire u0_u4_lmr_req_we_FF_INPUT_bF_buf5;
  wire u0_u4_lmr_req_we_FF_INPUT_bF_buf6;
  wire u0_u4_lmr_req_we_FF_INPUT_bF_buf7;
  wire u0_u4_rst_r1;
  wire u0_u4_rst_r2;
  wire u0_u4_tms_0__FF_INPUT;
  wire u0_u4_tms_10__FF_INPUT;
  wire u0_u4_tms_11__FF_INPUT;
  wire u0_u4_tms_12__FF_INPUT;
  wire u0_u4_tms_13__FF_INPUT;
  wire u0_u4_tms_14__FF_INPUT;
  wire u0_u4_tms_15__FF_INPUT;
  wire u0_u4_tms_16__FF_INPUT;
  wire u0_u4_tms_17__FF_INPUT;
  wire u0_u4_tms_18__FF_INPUT;
  wire u0_u4_tms_19__FF_INPUT;
  wire u0_u4_tms_1__FF_INPUT;
  wire u0_u4_tms_20__FF_INPUT;
  wire u0_u4_tms_21__FF_INPUT;
  wire u0_u4_tms_22__FF_INPUT;
  wire u0_u4_tms_23__FF_INPUT;
  wire u0_u4_tms_24__FF_INPUT;
  wire u0_u4_tms_25__FF_INPUT;
  wire u0_u4_tms_26__FF_INPUT;
  wire u0_u4_tms_27__FF_INPUT;
  wire u0_u4_tms_28__FF_INPUT;
  wire u0_u4_tms_29__FF_INPUT;
  wire u0_u4_tms_2__FF_INPUT;
  wire u0_u4_tms_30__FF_INPUT;
  wire u0_u4_tms_31__FF_INPUT;
  wire u0_u4_tms_3__FF_INPUT;
  wire u0_u4_tms_4__FF_INPUT;
  wire u0_u4_tms_5__FF_INPUT;
  wire u0_u4_tms_6__FF_INPUT;
  wire u0_u4_tms_7__FF_INPUT;
  wire u0_u4_tms_8__FF_INPUT;
  wire u0_u4_tms_9__FF_INPUT;
  wire u0_u4_wp_err;
  wire u0_u5__abc_45296_n201_1;
  wire u0_u5__abc_45296_n202_1;
  wire u0_u5__abc_45296_n203;
  wire u0_u5__abc_45296_n204_1;
  wire u0_u5__abc_45296_n205_1;
  wire u0_u5__abc_45296_n206;
  wire u0_u5__abc_45296_n207_1;
  wire u0_u5__abc_45296_n208_1;
  wire u0_u5__abc_45296_n209;
  wire u0_u5__abc_45296_n211_1;
  wire u0_u5__abc_45296_n212;
  wire u0_u5__abc_45296_n213_1;
  wire u0_u5__abc_45296_n214_1;
  wire u0_u5__abc_45296_n215;
  wire u0_u5__abc_45296_n217_1;
  wire u0_u5__abc_45296_n218;
  wire u0_u5__abc_45296_n218_bF_buf0;
  wire u0_u5__abc_45296_n218_bF_buf1;
  wire u0_u5__abc_45296_n218_bF_buf2;
  wire u0_u5__abc_45296_n218_bF_buf3;
  wire u0_u5__abc_45296_n218_bF_buf4;
  wire u0_u5__abc_45296_n218_bF_buf5;
  wire u0_u5__abc_45296_n218_bF_buf6;
  wire u0_u5__abc_45296_n218_bF_buf7;
  wire u0_u5__abc_45296_n219_1;
  wire u0_u5__abc_45296_n220_1;
  wire u0_u5__abc_45296_n221;
  wire u0_u5__abc_45296_n222_1;
  wire u0_u5__abc_45296_n224;
  wire u0_u5__abc_45296_n225_1;
  wire u0_u5__abc_45296_n226_1;
  wire u0_u5__abc_45296_n227;
  wire u0_u5__abc_45296_n228_1;
  wire u0_u5__abc_45296_n230;
  wire u0_u5__abc_45296_n231_1;
  wire u0_u5__abc_45296_n232_1;
  wire u0_u5__abc_45296_n233;
  wire u0_u5__abc_45296_n234_1;
  wire u0_u5__abc_45296_n236;
  wire u0_u5__abc_45296_n237_1;
  wire u0_u5__abc_45296_n238_1;
  wire u0_u5__abc_45296_n239;
  wire u0_u5__abc_45296_n240_1;
  wire u0_u5__abc_45296_n242;
  wire u0_u5__abc_45296_n243_1;
  wire u0_u5__abc_45296_n244_1;
  wire u0_u5__abc_45296_n245;
  wire u0_u5__abc_45296_n246_1;
  wire u0_u5__abc_45296_n248;
  wire u0_u5__abc_45296_n249_1;
  wire u0_u5__abc_45296_n250_1;
  wire u0_u5__abc_45296_n251;
  wire u0_u5__abc_45296_n252_1;
  wire u0_u5__abc_45296_n254;
  wire u0_u5__abc_45296_n255_1;
  wire u0_u5__abc_45296_n256;
  wire u0_u5__abc_45296_n257;
  wire u0_u5__abc_45296_n258;
  wire u0_u5__abc_45296_n260_1;
  wire u0_u5__abc_45296_n261;
  wire u0_u5__abc_45296_n262_1;
  wire u0_u5__abc_45296_n263;
  wire u0_u5__abc_45296_n264;
  wire u0_u5__abc_45296_n266_1;
  wire u0_u5__abc_45296_n267;
  wire u0_u5__abc_45296_n268_1;
  wire u0_u5__abc_45296_n269;
  wire u0_u5__abc_45296_n270;
  wire u0_u5__abc_45296_n272;
  wire u0_u5__abc_45296_n273_1;
  wire u0_u5__abc_45296_n274;
  wire u0_u5__abc_45296_n275_1;
  wire u0_u5__abc_45296_n276;
  wire u0_u5__abc_45296_n278;
  wire u0_u5__abc_45296_n279_1;
  wire u0_u5__abc_45296_n280;
  wire u0_u5__abc_45296_n281;
  wire u0_u5__abc_45296_n282;
  wire u0_u5__abc_45296_n284;
  wire u0_u5__abc_45296_n285_1;
  wire u0_u5__abc_45296_n286;
  wire u0_u5__abc_45296_n287_1;
  wire u0_u5__abc_45296_n288;
  wire u0_u5__abc_45296_n290;
  wire u0_u5__abc_45296_n291;
  wire u0_u5__abc_45296_n292;
  wire u0_u5__abc_45296_n293;
  wire u0_u5__abc_45296_n294;
  wire u0_u5__abc_45296_n296_1;
  wire u0_u5__abc_45296_n297;
  wire u0_u5__abc_45296_n298_1;
  wire u0_u5__abc_45296_n299;
  wire u0_u5__abc_45296_n300;
  wire u0_u5__abc_45296_n302;
  wire u0_u5__abc_45296_n303;
  wire u0_u5__abc_45296_n304;
  wire u0_u5__abc_45296_n305;
  wire u0_u5__abc_45296_n306;
  wire u0_u5__abc_45296_n308;
  wire u0_u5__abc_45296_n309;
  wire u0_u5__abc_45296_n310_1;
  wire u0_u5__abc_45296_n311;
  wire u0_u5__abc_45296_n312_1;
  wire u0_u5__abc_45296_n314_1;
  wire u0_u5__abc_45296_n315_1;
  wire u0_u5__abc_45296_n316_1;
  wire u0_u5__abc_45296_n317_1;
  wire u0_u5__abc_45296_n318;
  wire u0_u5__abc_45296_n320;
  wire u0_u5__abc_45296_n321_1;
  wire u0_u5__abc_45296_n322;
  wire u0_u5__abc_45296_n323_1;
  wire u0_u5__abc_45296_n324_1;
  wire u0_u5__abc_45296_n325;
  wire u0_u5__abc_45296_n326;
  wire u0_u5__abc_45296_n327;
  wire u0_u5__abc_45296_n328;
  wire u0_u5__abc_45296_n329;
  wire u0_u5__abc_45296_n330;
  wire u0_u5__abc_45296_n332;
  wire u0_u5__abc_45296_n333;
  wire u0_u5__abc_45296_n334;
  wire u0_u5__abc_45296_n335;
  wire u0_u5__abc_45296_n336;
  wire u0_u5__abc_45296_n338;
  wire u0_u5__abc_45296_n339;
  wire u0_u5__abc_45296_n340;
  wire u0_u5__abc_45296_n341;
  wire u0_u5__abc_45296_n342;
  wire u0_u5__abc_45296_n344;
  wire u0_u5__abc_45296_n345;
  wire u0_u5__abc_45296_n346;
  wire u0_u5__abc_45296_n347;
  wire u0_u5__abc_45296_n348;
  wire u0_u5__abc_45296_n350;
  wire u0_u5__abc_45296_n351;
  wire u0_u5__abc_45296_n352;
  wire u0_u5__abc_45296_n353;
  wire u0_u5__abc_45296_n354;
  wire u0_u5__abc_45296_n356;
  wire u0_u5__abc_45296_n357;
  wire u0_u5__abc_45296_n358;
  wire u0_u5__abc_45296_n359;
  wire u0_u5__abc_45296_n360;
  wire u0_u5__abc_45296_n362;
  wire u0_u5__abc_45296_n363;
  wire u0_u5__abc_45296_n364;
  wire u0_u5__abc_45296_n365;
  wire u0_u5__abc_45296_n366;
  wire u0_u5__abc_45296_n368;
  wire u0_u5__abc_45296_n369;
  wire u0_u5__abc_45296_n370;
  wire u0_u5__abc_45296_n371;
  wire u0_u5__abc_45296_n372;
  wire u0_u5__abc_45296_n374;
  wire u0_u5__abc_45296_n375;
  wire u0_u5__abc_45296_n376;
  wire u0_u5__abc_45296_n377;
  wire u0_u5__abc_45296_n378;
  wire u0_u5__abc_45296_n380;
  wire u0_u5__abc_45296_n381;
  wire u0_u5__abc_45296_n382;
  wire u0_u5__abc_45296_n383;
  wire u0_u5__abc_45296_n384;
  wire u0_u5__abc_45296_n386;
  wire u0_u5__abc_45296_n387;
  wire u0_u5__abc_45296_n388;
  wire u0_u5__abc_45296_n389;
  wire u0_u5__abc_45296_n390;
  wire u0_u5__abc_45296_n392;
  wire u0_u5__abc_45296_n393;
  wire u0_u5__abc_45296_n394;
  wire u0_u5__abc_45296_n395;
  wire u0_u5__abc_45296_n396;
  wire u0_u5__abc_45296_n398;
  wire u0_u5__abc_45296_n399;
  wire u0_u5__abc_45296_n400;
  wire u0_u5__abc_45296_n401;
  wire u0_u5__abc_45296_n402;
  wire u0_u5__abc_45296_n404;
  wire u0_u5__abc_45296_n405;
  wire u0_u5__abc_45296_n406;
  wire u0_u5__abc_45296_n407;
  wire u0_u5__abc_45296_n408;
  wire u0_u5__abc_45296_n410;
  wire u0_u5__abc_45296_n412;
  wire u0_u5__abc_45296_n413;
  wire u0_u5__abc_45296_n414;
  wire u0_u5__abc_45296_n415;
  wire u0_u5__abc_45296_n417;
  wire u0_u5__abc_45296_n418;
  wire u0_u5__abc_45296_n419;
  wire u0_u5__abc_45296_n420;
  wire u0_u5__abc_45296_n422;
  wire u0_u5__abc_45296_n423;
  wire u0_u5__abc_45296_n424;
  wire u0_u5__abc_45296_n425;
  wire u0_u5__abc_45296_n427;
  wire u0_u5__abc_45296_n428;
  wire u0_u5__abc_45296_n429;
  wire u0_u5__abc_45296_n430;
  wire u0_u5__abc_45296_n432;
  wire u0_u5__abc_45296_n433;
  wire u0_u5__abc_45296_n434;
  wire u0_u5__abc_45296_n435;
  wire u0_u5__abc_45296_n437;
  wire u0_u5__abc_45296_n438;
  wire u0_u5__abc_45296_n439;
  wire u0_u5__abc_45296_n440;
  wire u0_u5__abc_45296_n442;
  wire u0_u5__abc_45296_n443;
  wire u0_u5__abc_45296_n444;
  wire u0_u5__abc_45296_n445;
  wire u0_u5__abc_45296_n447;
  wire u0_u5__abc_45296_n448;
  wire u0_u5__abc_45296_n449;
  wire u0_u5__abc_45296_n450;
  wire u0_u5__abc_45296_n452;
  wire u0_u5__abc_45296_n453;
  wire u0_u5__abc_45296_n454;
  wire u0_u5__abc_45296_n455;
  wire u0_u5__abc_45296_n457;
  wire u0_u5__abc_45296_n458;
  wire u0_u5__abc_45296_n459;
  wire u0_u5__abc_45296_n460;
  wire u0_u5__abc_45296_n462;
  wire u0_u5__abc_45296_n463;
  wire u0_u5__abc_45296_n464;
  wire u0_u5__abc_45296_n465;
  wire u0_u5__abc_45296_n467;
  wire u0_u5__abc_45296_n468;
  wire u0_u5__abc_45296_n469;
  wire u0_u5__abc_45296_n470;
  wire u0_u5__abc_45296_n472;
  wire u0_u5__abc_45296_n473;
  wire u0_u5__abc_45296_n474;
  wire u0_u5__abc_45296_n475;
  wire u0_u5__abc_45296_n477;
  wire u0_u5__abc_45296_n478;
  wire u0_u5__abc_45296_n479;
  wire u0_u5__abc_45296_n480;
  wire u0_u5__abc_45296_n482;
  wire u0_u5__abc_45296_n483;
  wire u0_u5__abc_45296_n484;
  wire u0_u5__abc_45296_n485;
  wire u0_u5__abc_45296_n487;
  wire u0_u5__abc_45296_n488;
  wire u0_u5__abc_45296_n489;
  wire u0_u5__abc_45296_n490;
  wire u0_u5__abc_45296_n492;
  wire u0_u5__abc_45296_n493;
  wire u0_u5__abc_45296_n494;
  wire u0_u5__abc_45296_n495;
  wire u0_u5__abc_45296_n497;
  wire u0_u5__abc_45296_n498;
  wire u0_u5__abc_45296_n499;
  wire u0_u5__abc_45296_n500;
  wire u0_u5__abc_45296_n502;
  wire u0_u5__abc_45296_n503;
  wire u0_u5__abc_45296_n504;
  wire u0_u5__abc_45296_n505;
  wire u0_u5__abc_45296_n507;
  wire u0_u5__abc_45296_n508;
  wire u0_u5__abc_45296_n509;
  wire u0_u5__abc_45296_n510;
  wire u0_u5__abc_45296_n512;
  wire u0_u5__abc_45296_n513;
  wire u0_u5__abc_45296_n514;
  wire u0_u5__abc_45296_n515;
  wire u0_u5__abc_45296_n517;
  wire u0_u5__abc_45296_n518;
  wire u0_u5__abc_45296_n519;
  wire u0_u5__abc_45296_n520;
  wire u0_u5__abc_45296_n522;
  wire u0_u5__abc_45296_n523;
  wire u0_u5__abc_45296_n524;
  wire u0_u5__abc_45296_n525;
  wire u0_u5__abc_45296_n527;
  wire u0_u5__abc_45296_n528;
  wire u0_u5__abc_45296_n529;
  wire u0_u5__abc_45296_n530;
  wire u0_u5__abc_45296_n532;
  wire u0_u5__abc_45296_n533;
  wire u0_u5__abc_45296_n534;
  wire u0_u5__abc_45296_n535;
  wire u0_u5__abc_45296_n537;
  wire u0_u5__abc_45296_n538;
  wire u0_u5__abc_45296_n539;
  wire u0_u5__abc_45296_n540;
  wire u0_u5__abc_45296_n542;
  wire u0_u5__abc_45296_n543;
  wire u0_u5__abc_45296_n544;
  wire u0_u5__abc_45296_n545;
  wire u0_u5__abc_45296_n547;
  wire u0_u5__abc_45296_n548;
  wire u0_u5__abc_45296_n549;
  wire u0_u5__abc_45296_n550;
  wire u0_u5__abc_45296_n552;
  wire u0_u5__abc_45296_n553;
  wire u0_u5__abc_45296_n554;
  wire u0_u5__abc_45296_n555;
  wire u0_u5__abc_45296_n557;
  wire u0_u5__abc_45296_n558;
  wire u0_u5__abc_45296_n559;
  wire u0_u5__abc_45296_n560;
  wire u0_u5__abc_45296_n562;
  wire u0_u5__abc_45296_n563;
  wire u0_u5__abc_45296_n564;
  wire u0_u5__abc_45296_n565;
  wire u0_u5__abc_45296_n567;
  wire u0_u5__abc_45296_n568;
  wire u0_u5__abc_45296_n569;
  wire u0_u5__abc_45296_n570;
  wire u0_u5__abc_45296_n572;
  wire u0_u5__abc_45296_n573;
  wire u0_u5__abc_45296_n574;
  wire u0_u5__abc_45296_n575;
  wire u0_u5__abc_45296_n576;
  wire u0_u5__abc_45296_n577;
  wire u0_u5__abc_45296_n578;
  wire u0_u5__abc_45296_n579;
  wire u0_u5__abc_45296_n580;
  wire u0_u5__abc_45296_n581;
  wire u0_u5__abc_45296_n582;
  wire u0_u5__abc_45296_n583;
  wire u0_u5__abc_45296_n584;
  wire u0_u5__abc_45296_n585;
  wire u0_u5__abc_45296_n586;
  wire u0_u5__abc_45296_n587;
  wire u0_u5__abc_45296_n588;
  wire u0_u5__abc_45296_n589;
  wire u0_u5__abc_45296_n590;
  wire u0_u5__abc_45296_n591;
  wire u0_u5__abc_45296_n592;
  wire u0_u5__abc_45296_n593;
  wire u0_u5__abc_45296_n594;
  wire u0_u5__abc_45296_n595;
  wire u0_u5__abc_45296_n596;
  wire u0_u5__abc_45296_n597;
  wire u0_u5__abc_45296_n598;
  wire u0_u5__abc_45296_n599;
  wire u0_u5__abc_45296_n600;
  wire u0_u5__abc_45296_n601;
  wire u0_u5__abc_45296_n602;
  wire u0_u5__abc_45296_n603;
  wire u0_u5__abc_45296_n604;
  wire u0_u5__abc_45296_n605;
  wire u0_u5__abc_45296_n606;
  wire u0_u5__abc_45296_n607;
  wire u0_u5__abc_45296_n608;
  wire u0_u5__abc_45296_n609;
  wire u0_u5__abc_45296_n610;
  wire u0_u5__abc_45296_n611;
  wire u0_u5__abc_45296_n612;
  wire u0_u5__abc_45296_n613;
  wire u0_u5__abc_45296_n614;
  wire u0_u5__abc_45296_n615;
  wire u0_u5__abc_45296_n616;
  wire u0_u5__abc_45296_n617;
  wire u0_u5__abc_45296_n618;
  wire u0_u5__abc_45296_n619;
  wire u0_u5__abc_45296_n620;
  wire u0_u5__abc_45296_n621;
  wire u0_u5__abc_45296_n622;
  wire u0_u5__abc_45296_n623;
  wire u0_u5__abc_45296_n624;
  wire u0_u5__abc_45296_n625;
  wire u0_u5__abc_45296_n626;
  wire u0_u5__abc_45296_n627;
  wire u0_u5__abc_45296_n628;
  wire u0_u5__abc_45296_n629;
  wire u0_u5__abc_45296_n630;
  wire u0_u5__abc_45296_n631;
  wire u0_u5__abc_45296_n632;
  wire u0_u5__abc_45296_n633;
  wire u0_u5__abc_45296_n634;
  wire u0_u5__abc_45296_n635;
  wire u0_u5__abc_45296_n636;
  wire u0_u5__abc_45296_n637;
  wire u0_u5__abc_45296_n638;
  wire u0_u5__abc_45296_n640;
  wire u0_u5__abc_45296_n643;
  wire u0_u5__abc_45296_n644;
  wire u0_u5__abc_45296_n645;
  wire u0_u5__abc_45296_n646;
  wire u0_u5__abc_45296_n647;
  wire u0_u5__abc_45296_n648;
  wire u0_u5_addr_r_2_;
  wire u0_u5_addr_r_3_;
  wire u0_u5_addr_r_4_;
  wire u0_u5_addr_r_5_;
  wire u0_u5_addr_r_6_;
  wire u0_u5_csc_0__FF_INPUT;
  wire u0_u5_csc_10__FF_INPUT;
  wire u0_u5_csc_11__FF_INPUT;
  wire u0_u5_csc_12__FF_INPUT;
  wire u0_u5_csc_13__FF_INPUT;
  wire u0_u5_csc_14__FF_INPUT;
  wire u0_u5_csc_15__FF_INPUT;
  wire u0_u5_csc_16__FF_INPUT;
  wire u0_u5_csc_17__FF_INPUT;
  wire u0_u5_csc_18__FF_INPUT;
  wire u0_u5_csc_19__FF_INPUT;
  wire u0_u5_csc_1__FF_INPUT;
  wire u0_u5_csc_20__FF_INPUT;
  wire u0_u5_csc_21__FF_INPUT;
  wire u0_u5_csc_22__FF_INPUT;
  wire u0_u5_csc_23__FF_INPUT;
  wire u0_u5_csc_24__FF_INPUT;
  wire u0_u5_csc_25__FF_INPUT;
  wire u0_u5_csc_26__FF_INPUT;
  wire u0_u5_csc_27__FF_INPUT;
  wire u0_u5_csc_28__FF_INPUT;
  wire u0_u5_csc_29__FF_INPUT;
  wire u0_u5_csc_2__FF_INPUT;
  wire u0_u5_csc_30__FF_INPUT;
  wire u0_u5_csc_31__FF_INPUT;
  wire u0_u5_csc_3__FF_INPUT;
  wire u0_u5_csc_4__FF_INPUT;
  wire u0_u5_csc_5__FF_INPUT;
  wire u0_u5_csc_6__FF_INPUT;
  wire u0_u5_csc_7__FF_INPUT;
  wire u0_u5_csc_8__FF_INPUT;
  wire u0_u5_csc_9__FF_INPUT;
  wire u0_u5_init_req_FF_INPUT;
  wire u0_u5_init_req_we;
  wire u0_u5_init_req_we_FF_INPUT;
  wire u0_u5_init_req_we_FF_INPUT_bF_buf0;
  wire u0_u5_init_req_we_FF_INPUT_bF_buf1;
  wire u0_u5_init_req_we_FF_INPUT_bF_buf2;
  wire u0_u5_init_req_we_FF_INPUT_bF_buf3;
  wire u0_u5_init_req_we_FF_INPUT_bF_buf4;
  wire u0_u5_init_req_we_FF_INPUT_bF_buf5;
  wire u0_u5_init_req_we_FF_INPUT_bF_buf6;
  wire u0_u5_init_req_we_FF_INPUT_bF_buf7;
  wire u0_u5_inited;
  wire u0_u5_inited_FF_INPUT;
  wire u0_u5_lmr_req_FF_INPUT;
  wire u0_u5_lmr_req_we;
  wire u0_u5_lmr_req_we_FF_INPUT;
  wire u0_u5_lmr_req_we_FF_INPUT_bF_buf0;
  wire u0_u5_lmr_req_we_FF_INPUT_bF_buf1;
  wire u0_u5_lmr_req_we_FF_INPUT_bF_buf2;
  wire u0_u5_lmr_req_we_FF_INPUT_bF_buf3;
  wire u0_u5_lmr_req_we_FF_INPUT_bF_buf4;
  wire u0_u5_lmr_req_we_FF_INPUT_bF_buf5;
  wire u0_u5_lmr_req_we_FF_INPUT_bF_buf6;
  wire u0_u5_lmr_req_we_FF_INPUT_bF_buf7;
  wire u0_u5_rst_r1;
  wire u0_u5_rst_r2;
  wire u0_u5_tms_0__FF_INPUT;
  wire u0_u5_tms_10__FF_INPUT;
  wire u0_u5_tms_11__FF_INPUT;
  wire u0_u5_tms_12__FF_INPUT;
  wire u0_u5_tms_13__FF_INPUT;
  wire u0_u5_tms_14__FF_INPUT;
  wire u0_u5_tms_15__FF_INPUT;
  wire u0_u5_tms_16__FF_INPUT;
  wire u0_u5_tms_17__FF_INPUT;
  wire u0_u5_tms_18__FF_INPUT;
  wire u0_u5_tms_19__FF_INPUT;
  wire u0_u5_tms_1__FF_INPUT;
  wire u0_u5_tms_20__FF_INPUT;
  wire u0_u5_tms_21__FF_INPUT;
  wire u0_u5_tms_22__FF_INPUT;
  wire u0_u5_tms_23__FF_INPUT;
  wire u0_u5_tms_24__FF_INPUT;
  wire u0_u5_tms_25__FF_INPUT;
  wire u0_u5_tms_26__FF_INPUT;
  wire u0_u5_tms_27__FF_INPUT;
  wire u0_u5_tms_28__FF_INPUT;
  wire u0_u5_tms_29__FF_INPUT;
  wire u0_u5_tms_2__FF_INPUT;
  wire u0_u5_tms_30__FF_INPUT;
  wire u0_u5_tms_31__FF_INPUT;
  wire u0_u5_tms_3__FF_INPUT;
  wire u0_u5_tms_4__FF_INPUT;
  wire u0_u5_tms_5__FF_INPUT;
  wire u0_u5_tms_6__FF_INPUT;
  wire u0_u5_tms_7__FF_INPUT;
  wire u0_u5_tms_8__FF_INPUT;
  wire u0_u5_tms_9__FF_INPUT;
  wire u0_u5_wp_err;
  wire u0_wb_addr_r_2_;
  wire u0_wb_addr_r_3_;
  wire u0_wb_addr_r_4_;
  wire u0_wb_addr_r_5_;
  wire u0_wb_addr_r_6_;
  wire u0_wp_err;
  wire u0_wp_err_FF_INPUT;
  wire u1__abc_45852_n1000;
  wire u1__abc_45852_n1001;
  wire u1__abc_45852_n1002;
  wire u1__abc_45852_n1003;
  wire u1__abc_45852_n1004;
  wire u1__abc_45852_n1005;
  wire u1__abc_45852_n1006;
  wire u1__abc_45852_n1007;
  wire u1__abc_45852_n1008;
  wire u1__abc_45852_n1009;
  wire u1__abc_45852_n1010;
  wire u1__abc_45852_n1012;
  wire u1__abc_45852_n1013;
  wire u1__abc_45852_n1014;
  wire u1__abc_45852_n1015;
  wire u1__abc_45852_n1016;
  wire u1__abc_45852_n1017;
  wire u1__abc_45852_n1018;
  wire u1__abc_45852_n1019;
  wire u1__abc_45852_n1020;
  wire u1__abc_45852_n1021;
  wire u1__abc_45852_n1022;
  wire u1__abc_45852_n1023;
  wire u1__abc_45852_n1024;
  wire u1__abc_45852_n1025;
  wire u1__abc_45852_n1027;
  wire u1__abc_45852_n1028;
  wire u1__abc_45852_n1029;
  wire u1__abc_45852_n1030;
  wire u1__abc_45852_n1031;
  wire u1__abc_45852_n1032;
  wire u1__abc_45852_n1033;
  wire u1__abc_45852_n1034;
  wire u1__abc_45852_n1035;
  wire u1__abc_45852_n1036;
  wire u1__abc_45852_n1037;
  wire u1__abc_45852_n1038;
  wire u1__abc_45852_n1039;
  wire u1__abc_45852_n1040;
  wire u1__abc_45852_n1042;
  wire u1__abc_45852_n1043;
  wire u1__abc_45852_n1044;
  wire u1__abc_45852_n1045;
  wire u1__abc_45852_n1046;
  wire u1__abc_45852_n1047;
  wire u1__abc_45852_n1048;
  wire u1__abc_45852_n1049;
  wire u1__abc_45852_n1050;
  wire u1__abc_45852_n1051;
  wire u1__abc_45852_n1052;
  wire u1__abc_45852_n1053;
  wire u1__abc_45852_n1054;
  wire u1__abc_45852_n1055;
  wire u1__abc_45852_n1057;
  wire u1__abc_45852_n1058;
  wire u1__abc_45852_n1059;
  wire u1__abc_45852_n1060;
  wire u1__abc_45852_n1061;
  wire u1__abc_45852_n1062;
  wire u1__abc_45852_n1063;
  wire u1__abc_45852_n1064;
  wire u1__abc_45852_n1065;
  wire u1__abc_45852_n1066;
  wire u1__abc_45852_n1067;
  wire u1__abc_45852_n1068;
  wire u1__abc_45852_n1070;
  wire u1__abc_45852_n1071;
  wire u1__abc_45852_n1072;
  wire u1__abc_45852_n1073;
  wire u1__abc_45852_n1074;
  wire u1__abc_45852_n1075;
  wire u1__abc_45852_n1076;
  wire u1__abc_45852_n1077;
  wire u1__abc_45852_n1078;
  wire u1__abc_45852_n1079;
  wire u1__abc_45852_n1080;
  wire u1__abc_45852_n1081;
  wire u1__abc_45852_n1083;
  wire u1__abc_45852_n1084;
  wire u1__abc_45852_n1085;
  wire u1__abc_45852_n1086;
  wire u1__abc_45852_n1087;
  wire u1__abc_45852_n1088;
  wire u1__abc_45852_n1089;
  wire u1__abc_45852_n1090;
  wire u1__abc_45852_n1092;
  wire u1__abc_45852_n1093;
  wire u1__abc_45852_n1094;
  wire u1__abc_45852_n1095;
  wire u1__abc_45852_n1096;
  wire u1__abc_45852_n1097;
  wire u1__abc_45852_n1098;
  wire u1__abc_45852_n1099;
  wire u1__abc_45852_n1101;
  wire u1__abc_45852_n1102;
  wire u1__abc_45852_n1103;
  wire u1__abc_45852_n1104;
  wire u1__abc_45852_n1105;
  wire u1__abc_45852_n1106;
  wire u1__abc_45852_n1108;
  wire u1__abc_45852_n1109;
  wire u1__abc_45852_n1110;
  wire u1__abc_45852_n1111;
  wire u1__abc_45852_n1112;
  wire u1__abc_45852_n1113;
  wire u1__abc_45852_n1115;
  wire u1__abc_45852_n1116;
  wire u1__abc_45852_n1117;
  wire u1__abc_45852_n1118;
  wire u1__abc_45852_n1119;
  wire u1__abc_45852_n1120;
  wire u1__abc_45852_n1122;
  wire u1__abc_45852_n1123;
  wire u1__abc_45852_n1124;
  wire u1__abc_45852_n1125;
  wire u1__abc_45852_n1126;
  wire u1__abc_45852_n1127;
  wire u1__abc_45852_n1129;
  wire u1__abc_45852_n1130;
  wire u1__abc_45852_n1131;
  wire u1__abc_45852_n1132;
  wire u1__abc_45852_n1133;
  wire u1__abc_45852_n1134;
  wire u1__abc_45852_n1136;
  wire u1__abc_45852_n1137;
  wire u1__abc_45852_n1138;
  wire u1__abc_45852_n1139;
  wire u1__abc_45852_n1140;
  wire u1__abc_45852_n1141;
  wire u1__abc_45852_n1143;
  wire u1__abc_45852_n1144;
  wire u1__abc_45852_n1145;
  wire u1__abc_45852_n1146;
  wire u1__abc_45852_n1147;
  wire u1__abc_45852_n1148;
  wire u1__abc_45852_n1150;
  wire u1__abc_45852_n1151;
  wire u1__abc_45852_n1152;
  wire u1__abc_45852_n1153;
  wire u1__abc_45852_n1154;
  wire u1__abc_45852_n1155;
  wire u1__abc_45852_n1157;
  wire u1__abc_45852_n1158;
  wire u1__abc_45852_n1159;
  wire u1__abc_45852_n1160;
  wire u1__abc_45852_n1161;
  wire u1__abc_45852_n1162;
  wire u1__abc_45852_n1164;
  wire u1__abc_45852_n1165;
  wire u1__abc_45852_n1166;
  wire u1__abc_45852_n1167;
  wire u1__abc_45852_n1168;
  wire u1__abc_45852_n1169;
  wire u1__abc_45852_n1170;
  wire u1__abc_45852_n1171;
  wire u1__abc_45852_n1172;
  wire u1__abc_45852_n1173;
  wire u1__abc_45852_n1174;
  wire u1__abc_45852_n1175;
  wire u1__abc_45852_n1176;
  wire u1__abc_45852_n1177;
  wire u1__abc_45852_n1178;
  wire u1__abc_45852_n258_1;
  wire u1__abc_45852_n259_1;
  wire u1__abc_45852_n260_1;
  wire u1__abc_45852_n261;
  wire u1__abc_45852_n261_bF_buf0;
  wire u1__abc_45852_n261_bF_buf1;
  wire u1__abc_45852_n261_bF_buf2;
  wire u1__abc_45852_n261_bF_buf3;
  wire u1__abc_45852_n261_bF_buf4;
  wire u1__abc_45852_n262_1;
  wire u1__abc_45852_n263;
  wire u1__abc_45852_n264;
  wire u1__abc_45852_n265_1;
  wire u1__abc_45852_n267_1;
  wire u1__abc_45852_n268;
  wire u1__abc_45852_n269;
  wire u1__abc_45852_n270;
  wire u1__abc_45852_n271_1;
  wire u1__abc_45852_n272_1;
  wire u1__abc_45852_n273_1;
  wire u1__abc_45852_n274;
  wire u1__abc_45852_n275;
  wire u1__abc_45852_n276;
  wire u1__abc_45852_n276_bF_buf0;
  wire u1__abc_45852_n276_bF_buf1;
  wire u1__abc_45852_n276_bF_buf2;
  wire u1__abc_45852_n276_bF_buf3;
  wire u1__abc_45852_n276_bF_buf4;
  wire u1__abc_45852_n277;
  wire u1__abc_45852_n278_1;
  wire u1__abc_45852_n279_1;
  wire u1__abc_45852_n281;
  wire u1__abc_45852_n282;
  wire u1__abc_45852_n283;
  wire u1__abc_45852_n285_1;
  wire u1__abc_45852_n286_1;
  wire u1__abc_45852_n287_1;
  wire u1__abc_45852_n288;
  wire u1__abc_45852_n289;
  wire u1__abc_45852_n290;
  wire u1__abc_45852_n291;
  wire u1__abc_45852_n292_1;
  wire u1__abc_45852_n293_1;
  wire u1__abc_45852_n294_1;
  wire u1__abc_45852_n295;
  wire u1__abc_45852_n296;
  wire u1__abc_45852_n297;
  wire u1__abc_45852_n298;
  wire u1__abc_45852_n299_1;
  wire u1__abc_45852_n300_1;
  wire u1__abc_45852_n301_1;
  wire u1__abc_45852_n302;
  wire u1__abc_45852_n303;
  wire u1__abc_45852_n304;
  wire u1__abc_45852_n305;
  wire u1__abc_45852_n306_1;
  wire u1__abc_45852_n307_1;
  wire u1__abc_45852_n308_1;
  wire u1__abc_45852_n309;
  wire u1__abc_45852_n310;
  wire u1__abc_45852_n311;
  wire u1__abc_45852_n312;
  wire u1__abc_45852_n313_1;
  wire u1__abc_45852_n315_1;
  wire u1__abc_45852_n316;
  wire u1__abc_45852_n317;
  wire u1__abc_45852_n318;
  wire u1__abc_45852_n319;
  wire u1__abc_45852_n320_1;
  wire u1__abc_45852_n321_1;
  wire u1__abc_45852_n322_1;
  wire u1__abc_45852_n323;
  wire u1__abc_45852_n324;
  wire u1__abc_45852_n325;
  wire u1__abc_45852_n326;
  wire u1__abc_45852_n327_1;
  wire u1__abc_45852_n328_1;
  wire u1__abc_45852_n329_1;
  wire u1__abc_45852_n330;
  wire u1__abc_45852_n331;
  wire u1__abc_45852_n332;
  wire u1__abc_45852_n333_1;
  wire u1__abc_45852_n335_1;
  wire u1__abc_45852_n336;
  wire u1__abc_45852_n337;
  wire u1__abc_45852_n338;
  wire u1__abc_45852_n339_1;
  wire u1__abc_45852_n340_1;
  wire u1__abc_45852_n341_1;
  wire u1__abc_45852_n342;
  wire u1__abc_45852_n343;
  wire u1__abc_45852_n344;
  wire u1__abc_45852_n346_1;
  wire u1__abc_45852_n347_1;
  wire u1__abc_45852_n348;
  wire u1__abc_45852_n349;
  wire u1__abc_45852_n350;
  wire u1__abc_45852_n351_1;
  wire u1__abc_45852_n352_1;
  wire u1__abc_45852_n353_1;
  wire u1__abc_45852_n354;
  wire u1__abc_45852_n355;
  wire u1__abc_45852_n357_1;
  wire u1__abc_45852_n358_1;
  wire u1__abc_45852_n359_1;
  wire u1__abc_45852_n360;
  wire u1__abc_45852_n361;
  wire u1__abc_45852_n362;
  wire u1__abc_45852_n363_1;
  wire u1__abc_45852_n364_1;
  wire u1__abc_45852_n365_1;
  wire u1__abc_45852_n366;
  wire u1__abc_45852_n367;
  wire u1__abc_45852_n368;
  wire u1__abc_45852_n369_1;
  wire u1__abc_45852_n370_1;
  wire u1__abc_45852_n371_1;
  wire u1__abc_45852_n372;
  wire u1__abc_45852_n373;
  wire u1__abc_45852_n374;
  wire u1__abc_45852_n375_1;
  wire u1__abc_45852_n376_1;
  wire u1__abc_45852_n378;
  wire u1__abc_45852_n379;
  wire u1__abc_45852_n380;
  wire u1__abc_45852_n381_1;
  wire u1__abc_45852_n382_1;
  wire u1__abc_45852_n383_1;
  wire u1__abc_45852_n384;
  wire u1__abc_45852_n385;
  wire u1__abc_45852_n386;
  wire u1__abc_45852_n387_1;
  wire u1__abc_45852_n388_1;
  wire u1__abc_45852_n389_1;
  wire u1__abc_45852_n391;
  wire u1__abc_45852_n392;
  wire u1__abc_45852_n393_1;
  wire u1__abc_45852_n394_1;
  wire u1__abc_45852_n395_1;
  wire u1__abc_45852_n396;
  wire u1__abc_45852_n397;
  wire u1__abc_45852_n398;
  wire u1__abc_45852_n399_1;
  wire u1__abc_45852_n400_1;
  wire u1__abc_45852_n401_1;
  wire u1__abc_45852_n402;
  wire u1__abc_45852_n403;
  wire u1__abc_45852_n404;
  wire u1__abc_45852_n405_1;
  wire u1__abc_45852_n406_1;
  wire u1__abc_45852_n408;
  wire u1__abc_45852_n409;
  wire u1__abc_45852_n410;
  wire u1__abc_45852_n411_1;
  wire u1__abc_45852_n412_1;
  wire u1__abc_45852_n413_1;
  wire u1__abc_45852_n414;
  wire u1__abc_45852_n415;
  wire u1__abc_45852_n416;
  wire u1__abc_45852_n417_1;
  wire u1__abc_45852_n418_1;
  wire u1__abc_45852_n419_1;
  wire u1__abc_45852_n420_1;
  wire u1__abc_45852_n421_1;
  wire u1__abc_45852_n422_1;
  wire u1__abc_45852_n423_1;
  wire u1__abc_45852_n425_1;
  wire u1__abc_45852_n426_1;
  wire u1__abc_45852_n427_1;
  wire u1__abc_45852_n428_1;
  wire u1__abc_45852_n429_1;
  wire u1__abc_45852_n430_1;
  wire u1__abc_45852_n431_1;
  wire u1__abc_45852_n432_1;
  wire u1__abc_45852_n433_1;
  wire u1__abc_45852_n434_1;
  wire u1__abc_45852_n436_1;
  wire u1__abc_45852_n437_1;
  wire u1__abc_45852_n438_1;
  wire u1__abc_45852_n439_1;
  wire u1__abc_45852_n440_1;
  wire u1__abc_45852_n441_1;
  wire u1__abc_45852_n442_1;
  wire u1__abc_45852_n443_1;
  wire u1__abc_45852_n444_1;
  wire u1__abc_45852_n445_1;
  wire u1__abc_45852_n447_1;
  wire u1__abc_45852_n448_1;
  wire u1__abc_45852_n449_1;
  wire u1__abc_45852_n450_1;
  wire u1__abc_45852_n451_1;
  wire u1__abc_45852_n452_1;
  wire u1__abc_45852_n453_1;
  wire u1__abc_45852_n454_1;
  wire u1__abc_45852_n455_1;
  wire u1__abc_45852_n456_1;
  wire u1__abc_45852_n457_1;
  wire u1__abc_45852_n458_1;
  wire u1__abc_45852_n460_1;
  wire u1__abc_45852_n461_1;
  wire u1__abc_45852_n462_1;
  wire u1__abc_45852_n463_1;
  wire u1__abc_45852_n464_1;
  wire u1__abc_45852_n465_1;
  wire u1__abc_45852_n466_1;
  wire u1__abc_45852_n467;
  wire u1__abc_45852_n468_1;
  wire u1__abc_45852_n469;
  wire u1__abc_45852_n470_1;
  wire u1__abc_45852_n471;
  wire u1__abc_45852_n472_1;
  wire u1__abc_45852_n474_1;
  wire u1__abc_45852_n475;
  wire u1__abc_45852_n476_1;
  wire u1__abc_45852_n477_1;
  wire u1__abc_45852_n478;
  wire u1__abc_45852_n479;
  wire u1__abc_45852_n480;
  wire u1__abc_45852_n481;
  wire u1__abc_45852_n482;
  wire u1__abc_45852_n483_1;
  wire u1__abc_45852_n484;
  wire u1__abc_45852_n485;
  wire u1__abc_45852_n486;
  wire u1__abc_45852_n487;
  wire u1__abc_45852_n488_1;
  wire u1__abc_45852_n490_1;
  wire u1__abc_45852_n491;
  wire u1__abc_45852_n492;
  wire u1__abc_45852_n493;
  wire u1__abc_45852_n494_1;
  wire u1__abc_45852_n495;
  wire u1__abc_45852_n496_1;
  wire u1__abc_45852_n497;
  wire u1__abc_45852_n498;
  wire u1__abc_45852_n499;
  wire u1__abc_45852_n500_1;
  wire u1__abc_45852_n501;
  wire u1__abc_45852_n503;
  wire u1__abc_45852_n504;
  wire u1__abc_45852_n505;
  wire u1__abc_45852_n506_1;
  wire u1__abc_45852_n507;
  wire u1__abc_45852_n508_1;
  wire u1__abc_45852_n509;
  wire u1__abc_45852_n510;
  wire u1__abc_45852_n511;
  wire u1__abc_45852_n512_1;
  wire u1__abc_45852_n513;
  wire u1__abc_45852_n514_1;
  wire u1__abc_45852_n516;
  wire u1__abc_45852_n517;
  wire u1__abc_45852_n518_1;
  wire u1__abc_45852_n519;
  wire u1__abc_45852_n520_1;
  wire u1__abc_45852_n521;
  wire u1__abc_45852_n522;
  wire u1__abc_45852_n524_1;
  wire u1__abc_45852_n525;
  wire u1__abc_45852_n527;
  wire u1__abc_45852_n528;
  wire u1__abc_45852_n530_1;
  wire u1__abc_45852_n531;
  wire u1__abc_45852_n533;
  wire u1__abc_45852_n534;
  wire u1__abc_45852_n536_1;
  wire u1__abc_45852_n537;
  wire u1__abc_45852_n539;
  wire u1__abc_45852_n540;
  wire u1__abc_45852_n542_1;
  wire u1__abc_45852_n543;
  wire u1__abc_45852_n545;
  wire u1__abc_45852_n546;
  wire u1__abc_45852_n547;
  wire u1__abc_45852_n548_1;
  wire u1__abc_45852_n550_1;
  wire u1__abc_45852_n551;
  wire u1__abc_45852_n552;
  wire u1__abc_45852_n554_1;
  wire u1__abc_45852_n554_1_bF_buf0;
  wire u1__abc_45852_n554_1_bF_buf1;
  wire u1__abc_45852_n554_1_bF_buf2;
  wire u1__abc_45852_n554_1_bF_buf3;
  wire u1__abc_45852_n554_1_bF_buf4;
  wire u1__abc_45852_n555;
  wire u1__abc_45852_n556;
  wire u1__abc_45852_n556_bF_buf0;
  wire u1__abc_45852_n556_bF_buf1;
  wire u1__abc_45852_n556_bF_buf2;
  wire u1__abc_45852_n556_bF_buf3;
  wire u1__abc_45852_n557_1;
  wire u1__abc_45852_n558;
  wire u1__abc_45852_n559;
  wire u1__abc_45852_n560_1;
  wire u1__abc_45852_n561;
  wire u1__abc_45852_n562;
  wire u1__abc_45852_n562_bF_buf0;
  wire u1__abc_45852_n562_bF_buf1;
  wire u1__abc_45852_n562_bF_buf2;
  wire u1__abc_45852_n562_bF_buf3;
  wire u1__abc_45852_n563;
  wire u1__abc_45852_n564_1;
  wire u1__abc_45852_n565;
  wire u1__abc_45852_n566;
  wire u1__abc_45852_n568;
  wire u1__abc_45852_n569;
  wire u1__abc_45852_n570_1;
  wire u1__abc_45852_n571;
  wire u1__abc_45852_n572;
  wire u1__abc_45852_n573_1;
  wire u1__abc_45852_n574;
  wire u1__abc_45852_n575;
  wire u1__abc_45852_n576_1;
  wire u1__abc_45852_n577;
  wire u1__abc_45852_n579_1;
  wire u1__abc_45852_n580;
  wire u1__abc_45852_n581;
  wire u1__abc_45852_n582_1;
  wire u1__abc_45852_n583;
  wire u1__abc_45852_n584;
  wire u1__abc_45852_n585_1;
  wire u1__abc_45852_n586;
  wire u1__abc_45852_n587;
  wire u1__abc_45852_n588_1;
  wire u1__abc_45852_n590_1;
  wire u1__abc_45852_n591;
  wire u1__abc_45852_n592;
  wire u1__abc_45852_n593;
  wire u1__abc_45852_n594;
  wire u1__abc_45852_n595_1;
  wire u1__abc_45852_n596;
  wire u1__abc_45852_n597_1;
  wire u1__abc_45852_n598;
  wire u1__abc_45852_n599_1;
  wire u1__abc_45852_n601_1;
  wire u1__abc_45852_n602;
  wire u1__abc_45852_n603;
  wire u1__abc_45852_n604;
  wire u1__abc_45852_n605;
  wire u1__abc_45852_n606;
  wire u1__abc_45852_n607;
  wire u1__abc_45852_n608;
  wire u1__abc_45852_n609;
  wire u1__abc_45852_n610;
  wire u1__abc_45852_n612;
  wire u1__abc_45852_n613;
  wire u1__abc_45852_n614;
  wire u1__abc_45852_n615;
  wire u1__abc_45852_n616;
  wire u1__abc_45852_n617;
  wire u1__abc_45852_n618;
  wire u1__abc_45852_n619;
  wire u1__abc_45852_n620;
  wire u1__abc_45852_n621;
  wire u1__abc_45852_n623;
  wire u1__abc_45852_n624;
  wire u1__abc_45852_n625;
  wire u1__abc_45852_n626;
  wire u1__abc_45852_n627;
  wire u1__abc_45852_n628;
  wire u1__abc_45852_n629;
  wire u1__abc_45852_n630;
  wire u1__abc_45852_n631;
  wire u1__abc_45852_n632;
  wire u1__abc_45852_n634;
  wire u1__abc_45852_n635;
  wire u1__abc_45852_n636;
  wire u1__abc_45852_n637;
  wire u1__abc_45852_n638;
  wire u1__abc_45852_n639;
  wire u1__abc_45852_n640;
  wire u1__abc_45852_n641;
  wire u1__abc_45852_n642;
  wire u1__abc_45852_n643;
  wire u1__abc_45852_n645;
  wire u1__abc_45852_n646;
  wire u1__abc_45852_n647;
  wire u1__abc_45852_n648;
  wire u1__abc_45852_n649;
  wire u1__abc_45852_n650;
  wire u1__abc_45852_n651;
  wire u1__abc_45852_n652;
  wire u1__abc_45852_n653;
  wire u1__abc_45852_n654;
  wire u1__abc_45852_n656;
  wire u1__abc_45852_n657;
  wire u1__abc_45852_n658;
  wire u1__abc_45852_n659;
  wire u1__abc_45852_n660;
  wire u1__abc_45852_n661;
  wire u1__abc_45852_n662;
  wire u1__abc_45852_n663;
  wire u1__abc_45852_n664;
  wire u1__abc_45852_n665;
  wire u1__abc_45852_n667;
  wire u1__abc_45852_n668;
  wire u1__abc_45852_n669;
  wire u1__abc_45852_n670;
  wire u1__abc_45852_n671;
  wire u1__abc_45852_n672;
  wire u1__abc_45852_n673;
  wire u1__abc_45852_n674;
  wire u1__abc_45852_n675;
  wire u1__abc_45852_n676;
  wire u1__abc_45852_n678;
  wire u1__abc_45852_n679;
  wire u1__abc_45852_n680;
  wire u1__abc_45852_n681;
  wire u1__abc_45852_n682;
  wire u1__abc_45852_n683;
  wire u1__abc_45852_n684;
  wire u1__abc_45852_n685;
  wire u1__abc_45852_n686;
  wire u1__abc_45852_n687;
  wire u1__abc_45852_n689;
  wire u1__abc_45852_n690;
  wire u1__abc_45852_n691;
  wire u1__abc_45852_n692;
  wire u1__abc_45852_n693;
  wire u1__abc_45852_n694;
  wire u1__abc_45852_n695;
  wire u1__abc_45852_n696;
  wire u1__abc_45852_n697;
  wire u1__abc_45852_n698;
  wire u1__abc_45852_n700;
  wire u1__abc_45852_n701;
  wire u1__abc_45852_n702;
  wire u1__abc_45852_n703;
  wire u1__abc_45852_n704;
  wire u1__abc_45852_n705;
  wire u1__abc_45852_n706;
  wire u1__abc_45852_n707;
  wire u1__abc_45852_n708;
  wire u1__abc_45852_n709;
  wire u1__abc_45852_n711;
  wire u1__abc_45852_n712;
  wire u1__abc_45852_n713;
  wire u1__abc_45852_n714;
  wire u1__abc_45852_n715;
  wire u1__abc_45852_n716;
  wire u1__abc_45852_n717;
  wire u1__abc_45852_n718;
  wire u1__abc_45852_n719;
  wire u1__abc_45852_n720;
  wire u1__abc_45852_n722;
  wire u1__abc_45852_n723;
  wire u1__abc_45852_n724;
  wire u1__abc_45852_n725;
  wire u1__abc_45852_n726;
  wire u1__abc_45852_n727;
  wire u1__abc_45852_n728;
  wire u1__abc_45852_n729;
  wire u1__abc_45852_n730;
  wire u1__abc_45852_n731;
  wire u1__abc_45852_n733;
  wire u1__abc_45852_n734;
  wire u1__abc_45852_n735;
  wire u1__abc_45852_n736;
  wire u1__abc_45852_n737;
  wire u1__abc_45852_n738;
  wire u1__abc_45852_n739;
  wire u1__abc_45852_n740;
  wire u1__abc_45852_n741;
  wire u1__abc_45852_n742;
  wire u1__abc_45852_n744;
  wire u1__abc_45852_n745;
  wire u1__abc_45852_n746;
  wire u1__abc_45852_n747;
  wire u1__abc_45852_n748;
  wire u1__abc_45852_n749;
  wire u1__abc_45852_n750;
  wire u1__abc_45852_n751;
  wire u1__abc_45852_n752;
  wire u1__abc_45852_n753;
  wire u1__abc_45852_n755;
  wire u1__abc_45852_n756;
  wire u1__abc_45852_n757;
  wire u1__abc_45852_n758;
  wire u1__abc_45852_n759;
  wire u1__abc_45852_n760;
  wire u1__abc_45852_n761;
  wire u1__abc_45852_n762;
  wire u1__abc_45852_n763;
  wire u1__abc_45852_n764;
  wire u1__abc_45852_n766;
  wire u1__abc_45852_n767;
  wire u1__abc_45852_n768;
  wire u1__abc_45852_n769;
  wire u1__abc_45852_n770;
  wire u1__abc_45852_n771;
  wire u1__abc_45852_n772;
  wire u1__abc_45852_n773;
  wire u1__abc_45852_n774;
  wire u1__abc_45852_n775;
  wire u1__abc_45852_n777;
  wire u1__abc_45852_n778;
  wire u1__abc_45852_n779;
  wire u1__abc_45852_n780;
  wire u1__abc_45852_n781;
  wire u1__abc_45852_n782;
  wire u1__abc_45852_n783;
  wire u1__abc_45852_n784;
  wire u1__abc_45852_n785;
  wire u1__abc_45852_n786;
  wire u1__abc_45852_n788;
  wire u1__abc_45852_n789;
  wire u1__abc_45852_n790;
  wire u1__abc_45852_n791;
  wire u1__abc_45852_n792;
  wire u1__abc_45852_n793;
  wire u1__abc_45852_n794;
  wire u1__abc_45852_n795;
  wire u1__abc_45852_n796;
  wire u1__abc_45852_n797;
  wire u1__abc_45852_n799;
  wire u1__abc_45852_n800;
  wire u1__abc_45852_n801;
  wire u1__abc_45852_n802;
  wire u1__abc_45852_n803;
  wire u1__abc_45852_n804;
  wire u1__abc_45852_n805;
  wire u1__abc_45852_n806;
  wire u1__abc_45852_n807;
  wire u1__abc_45852_n809;
  wire u1__abc_45852_n810;
  wire u1__abc_45852_n811;
  wire u1__abc_45852_n812;
  wire u1__abc_45852_n813;
  wire u1__abc_45852_n814;
  wire u1__abc_45852_n815;
  wire u1__abc_45852_n816;
  wire u1__abc_45852_n817;
  wire u1__abc_45852_n818;
  wire u1__abc_45852_n820;
  wire u1__abc_45852_n821;
  wire u1__abc_45852_n821_bF_buf0;
  wire u1__abc_45852_n821_bF_buf1;
  wire u1__abc_45852_n821_bF_buf2;
  wire u1__abc_45852_n821_bF_buf3;
  wire u1__abc_45852_n822;
  wire u1__abc_45852_n824;
  wire u1__abc_45852_n825;
  wire u1__abc_45852_n827;
  wire u1__abc_45852_n828;
  wire u1__abc_45852_n830;
  wire u1__abc_45852_n831;
  wire u1__abc_45852_n833;
  wire u1__abc_45852_n834;
  wire u1__abc_45852_n836;
  wire u1__abc_45852_n837;
  wire u1__abc_45852_n839;
  wire u1__abc_45852_n840;
  wire u1__abc_45852_n842;
  wire u1__abc_45852_n843;
  wire u1__abc_45852_n845;
  wire u1__abc_45852_n846;
  wire u1__abc_45852_n848;
  wire u1__abc_45852_n849;
  wire u1__abc_45852_n851;
  wire u1__abc_45852_n852;
  wire u1__abc_45852_n854;
  wire u1__abc_45852_n855;
  wire u1__abc_45852_n857;
  wire u1__abc_45852_n858;
  wire u1__abc_45852_n860;
  wire u1__abc_45852_n861;
  wire u1__abc_45852_n863;
  wire u1__abc_45852_n864;
  wire u1__abc_45852_n866;
  wire u1__abc_45852_n867;
  wire u1__abc_45852_n869;
  wire u1__abc_45852_n870;
  wire u1__abc_45852_n872;
  wire u1__abc_45852_n873;
  wire u1__abc_45852_n875;
  wire u1__abc_45852_n876;
  wire u1__abc_45852_n878;
  wire u1__abc_45852_n879;
  wire u1__abc_45852_n881;
  wire u1__abc_45852_n882;
  wire u1__abc_45852_n884;
  wire u1__abc_45852_n885;
  wire u1__abc_45852_n887;
  wire u1__abc_45852_n888;
  wire u1__abc_45852_n890;
  wire u1__abc_45852_n891;
  wire u1__abc_45852_n893;
  wire u1__abc_45852_n893_bF_buf0;
  wire u1__abc_45852_n893_bF_buf1;
  wire u1__abc_45852_n893_bF_buf2;
  wire u1__abc_45852_n893_bF_buf3;
  wire u1__abc_45852_n893_bF_buf4;
  wire u1__abc_45852_n894;
  wire u1__abc_45852_n895;
  wire u1__abc_45852_n896;
  wire u1__abc_45852_n897;
  wire u1__abc_45852_n897_bF_buf0;
  wire u1__abc_45852_n897_bF_buf1;
  wire u1__abc_45852_n897_bF_buf2;
  wire u1__abc_45852_n897_bF_buf3;
  wire u1__abc_45852_n898;
  wire u1__abc_45852_n899;
  wire u1__abc_45852_n900;
  wire u1__abc_45852_n901;
  wire u1__abc_45852_n901_bF_buf0;
  wire u1__abc_45852_n901_bF_buf1;
  wire u1__abc_45852_n901_bF_buf2;
  wire u1__abc_45852_n901_bF_buf3;
  wire u1__abc_45852_n901_bF_buf4;
  wire u1__abc_45852_n902;
  wire u1__abc_45852_n903;
  wire u1__abc_45852_n903_bF_buf0;
  wire u1__abc_45852_n903_bF_buf1;
  wire u1__abc_45852_n903_bF_buf2;
  wire u1__abc_45852_n903_bF_buf3;
  wire u1__abc_45852_n904;
  wire u1__abc_45852_n905;
  wire u1__abc_45852_n906;
  wire u1__abc_45852_n907;
  wire u1__abc_45852_n908;
  wire u1__abc_45852_n909;
  wire u1__abc_45852_n910;
  wire u1__abc_45852_n911;
  wire u1__abc_45852_n912;
  wire u1__abc_45852_n913;
  wire u1__abc_45852_n914;
  wire u1__abc_45852_n915;
  wire u1__abc_45852_n916;
  wire u1__abc_45852_n917;
  wire u1__abc_45852_n918;
  wire u1__abc_45852_n919;
  wire u1__abc_45852_n920;
  wire u1__abc_45852_n922;
  wire u1__abc_45852_n923;
  wire u1__abc_45852_n924;
  wire u1__abc_45852_n925;
  wire u1__abc_45852_n926;
  wire u1__abc_45852_n927;
  wire u1__abc_45852_n928;
  wire u1__abc_45852_n929;
  wire u1__abc_45852_n930;
  wire u1__abc_45852_n931;
  wire u1__abc_45852_n932;
  wire u1__abc_45852_n933;
  wire u1__abc_45852_n934;
  wire u1__abc_45852_n935;
  wire u1__abc_45852_n937;
  wire u1__abc_45852_n938;
  wire u1__abc_45852_n939;
  wire u1__abc_45852_n940;
  wire u1__abc_45852_n941;
  wire u1__abc_45852_n942;
  wire u1__abc_45852_n943;
  wire u1__abc_45852_n944;
  wire u1__abc_45852_n945;
  wire u1__abc_45852_n946;
  wire u1__abc_45852_n947;
  wire u1__abc_45852_n948;
  wire u1__abc_45852_n949;
  wire u1__abc_45852_n950;
  wire u1__abc_45852_n952;
  wire u1__abc_45852_n953;
  wire u1__abc_45852_n954;
  wire u1__abc_45852_n955;
  wire u1__abc_45852_n956;
  wire u1__abc_45852_n957;
  wire u1__abc_45852_n958;
  wire u1__abc_45852_n959;
  wire u1__abc_45852_n960;
  wire u1__abc_45852_n961;
  wire u1__abc_45852_n962;
  wire u1__abc_45852_n963;
  wire u1__abc_45852_n964;
  wire u1__abc_45852_n965;
  wire u1__abc_45852_n967;
  wire u1__abc_45852_n968;
  wire u1__abc_45852_n969;
  wire u1__abc_45852_n970;
  wire u1__abc_45852_n971;
  wire u1__abc_45852_n972;
  wire u1__abc_45852_n973;
  wire u1__abc_45852_n974;
  wire u1__abc_45852_n975;
  wire u1__abc_45852_n976;
  wire u1__abc_45852_n977;
  wire u1__abc_45852_n978;
  wire u1__abc_45852_n979;
  wire u1__abc_45852_n980;
  wire u1__abc_45852_n982;
  wire u1__abc_45852_n983;
  wire u1__abc_45852_n984;
  wire u1__abc_45852_n985;
  wire u1__abc_45852_n986;
  wire u1__abc_45852_n987;
  wire u1__abc_45852_n988;
  wire u1__abc_45852_n989;
  wire u1__abc_45852_n990;
  wire u1__abc_45852_n991;
  wire u1__abc_45852_n992;
  wire u1__abc_45852_n993;
  wire u1__abc_45852_n994;
  wire u1__abc_45852_n995;
  wire u1__abc_45852_n997;
  wire u1__abc_45852_n998;
  wire u1__abc_45852_n999;
  wire u1_acs_addr_0_;
  wire u1_acs_addr_0__FF_INPUT;
  wire u1_acs_addr_10_;
  wire u1_acs_addr_10__FF_INPUT;
  wire u1_acs_addr_11_;
  wire u1_acs_addr_11__FF_INPUT;
  wire u1_acs_addr_12_;
  wire u1_acs_addr_12__FF_INPUT;
  wire u1_acs_addr_13_;
  wire u1_acs_addr_13__FF_INPUT;
  wire u1_acs_addr_14_;
  wire u1_acs_addr_14__FF_INPUT;
  wire u1_acs_addr_15_;
  wire u1_acs_addr_15__FF_INPUT;
  wire u1_acs_addr_16_;
  wire u1_acs_addr_16__FF_INPUT;
  wire u1_acs_addr_17_;
  wire u1_acs_addr_17__FF_INPUT;
  wire u1_acs_addr_18_;
  wire u1_acs_addr_18__FF_INPUT;
  wire u1_acs_addr_19_;
  wire u1_acs_addr_19__FF_INPUT;
  wire u1_acs_addr_1_;
  wire u1_acs_addr_1__FF_INPUT;
  wire u1_acs_addr_20_;
  wire u1_acs_addr_20__FF_INPUT;
  wire u1_acs_addr_21_;
  wire u1_acs_addr_21__FF_INPUT;
  wire u1_acs_addr_22_;
  wire u1_acs_addr_22__FF_INPUT;
  wire u1_acs_addr_23_;
  wire u1_acs_addr_23__FF_INPUT;
  wire u1_acs_addr_2_;
  wire u1_acs_addr_2__FF_INPUT;
  wire u1_acs_addr_3_;
  wire u1_acs_addr_3__FF_INPUT;
  wire u1_acs_addr_4_;
  wire u1_acs_addr_4__FF_INPUT;
  wire u1_acs_addr_5_;
  wire u1_acs_addr_5__FF_INPUT;
  wire u1_acs_addr_6_;
  wire u1_acs_addr_6__FF_INPUT;
  wire u1_acs_addr_7_;
  wire u1_acs_addr_7__FF_INPUT;
  wire u1_acs_addr_8_;
  wire u1_acs_addr_8__FF_INPUT;
  wire u1_acs_addr_9_;
  wire u1_acs_addr_9__FF_INPUT;
  wire u1_acs_addr_pl1_0_;
  wire u1_acs_addr_pl1_10_;
  wire u1_acs_addr_pl1_11_;
  wire u1_acs_addr_pl1_12_;
  wire u1_acs_addr_pl1_13_;
  wire u1_acs_addr_pl1_14_;
  wire u1_acs_addr_pl1_15_;
  wire u1_acs_addr_pl1_16_;
  wire u1_acs_addr_pl1_17_;
  wire u1_acs_addr_pl1_18_;
  wire u1_acs_addr_pl1_19_;
  wire u1_acs_addr_pl1_1_;
  wire u1_acs_addr_pl1_20_;
  wire u1_acs_addr_pl1_21_;
  wire u1_acs_addr_pl1_22_;
  wire u1_acs_addr_pl1_23_;
  wire u1_acs_addr_pl1_2_;
  wire u1_acs_addr_pl1_3_;
  wire u1_acs_addr_pl1_4_;
  wire u1_acs_addr_pl1_5_;
  wire u1_acs_addr_pl1_6_;
  wire u1_acs_addr_pl1_7_;
  wire u1_acs_addr_pl1_8_;
  wire u1_acs_addr_pl1_9_;
  wire u1_bank_adr_0__FF_INPUT;
  wire u1_bank_adr_1__FF_INPUT;
  wire u1_bas;
  wire u1_col_adr_0_;
  wire u1_col_adr_0__FF_INPUT;
  wire u1_col_adr_1_;
  wire u1_col_adr_1__FF_INPUT;
  wire u1_col_adr_2_;
  wire u1_col_adr_2__FF_INPUT;
  wire u1_col_adr_3_;
  wire u1_col_adr_3__FF_INPUT;
  wire u1_col_adr_4_;
  wire u1_col_adr_4__FF_INPUT;
  wire u1_col_adr_5_;
  wire u1_col_adr_5__FF_INPUT;
  wire u1_col_adr_6_;
  wire u1_col_adr_6__FF_INPUT;
  wire u1_col_adr_7_;
  wire u1_col_adr_7__FF_INPUT;
  wire u1_col_adr_8_;
  wire u1_col_adr_8__FF_INPUT;
  wire u1_col_adr_9_;
  wire u1_col_adr_9__FF_INPUT;
  wire u1_row_adr_0__FF_INPUT;
  wire u1_row_adr_10__FF_INPUT;
  wire u1_row_adr_11__FF_INPUT;
  wire u1_row_adr_12__FF_INPUT;
  wire u1_row_adr_1__FF_INPUT;
  wire u1_row_adr_2__FF_INPUT;
  wire u1_row_adr_3__FF_INPUT;
  wire u1_row_adr_4__FF_INPUT;
  wire u1_row_adr_5__FF_INPUT;
  wire u1_row_adr_6__FF_INPUT;
  wire u1_row_adr_7__FF_INPUT;
  wire u1_row_adr_8__FF_INPUT;
  wire u1_row_adr_9__FF_INPUT;
  wire u1_sram_addr_0_;
  wire u1_sram_addr_0__FF_INPUT;
  wire u1_sram_addr_10_;
  wire u1_sram_addr_10__FF_INPUT;
  wire u1_sram_addr_11_;
  wire u1_sram_addr_11__FF_INPUT;
  wire u1_sram_addr_12_;
  wire u1_sram_addr_12__FF_INPUT;
  wire u1_sram_addr_13_;
  wire u1_sram_addr_13__FF_INPUT;
  wire u1_sram_addr_14_;
  wire u1_sram_addr_14__FF_INPUT;
  wire u1_sram_addr_15_;
  wire u1_sram_addr_15__FF_INPUT;
  wire u1_sram_addr_16_;
  wire u1_sram_addr_16__FF_INPUT;
  wire u1_sram_addr_17_;
  wire u1_sram_addr_17__FF_INPUT;
  wire u1_sram_addr_18_;
  wire u1_sram_addr_18__FF_INPUT;
  wire u1_sram_addr_19_;
  wire u1_sram_addr_19__FF_INPUT;
  wire u1_sram_addr_1_;
  wire u1_sram_addr_1__FF_INPUT;
  wire u1_sram_addr_20_;
  wire u1_sram_addr_20__FF_INPUT;
  wire u1_sram_addr_21_;
  wire u1_sram_addr_21__FF_INPUT;
  wire u1_sram_addr_22_;
  wire u1_sram_addr_22__FF_INPUT;
  wire u1_sram_addr_23_;
  wire u1_sram_addr_23__FF_INPUT;
  wire u1_sram_addr_2_;
  wire u1_sram_addr_2__FF_INPUT;
  wire u1_sram_addr_3_;
  wire u1_sram_addr_3__FF_INPUT;
  wire u1_sram_addr_4_;
  wire u1_sram_addr_4__FF_INPUT;
  wire u1_sram_addr_5_;
  wire u1_sram_addr_5__FF_INPUT;
  wire u1_sram_addr_6_;
  wire u1_sram_addr_6__FF_INPUT;
  wire u1_sram_addr_7_;
  wire u1_sram_addr_7__FF_INPUT;
  wire u1_sram_addr_8_;
  wire u1_sram_addr_8__FF_INPUT;
  wire u1_sram_addr_9_;
  wire u1_sram_addr_9__FF_INPUT;
  wire u1_u0__abc_45749_n101;
  wire u1_u0__abc_45749_n102;
  wire u1_u0__abc_45749_n104;
  wire u1_u0__abc_45749_n105;
  wire u1_u0__abc_45749_n106;
  wire u1_u0__abc_45749_n108;
  wire u1_u0__abc_45749_n109;
  wire u1_u0__abc_45749_n110;
  wire u1_u0__abc_45749_n112;
  wire u1_u0__abc_45749_n113;
  wire u1_u0__abc_45749_n114;
  wire u1_u0__abc_45749_n116;
  wire u1_u0__abc_45749_n117;
  wire u1_u0__abc_45749_n118;
  wire u1_u0__abc_45749_n120;
  wire u1_u0__abc_45749_n121;
  wire u1_u0__abc_45749_n122;
  wire u1_u0__abc_45749_n123;
  wire u1_u0__abc_45749_n125;
  wire u1_u0__abc_45749_n126;
  wire u1_u0__abc_45749_n127;
  wire u1_u0__abc_45749_n129;
  wire u1_u0__abc_45749_n130;
  wire u1_u0__abc_45749_n131;
  wire u1_u0__abc_45749_n132;
  wire u1_u0__abc_45749_n133;
  wire u1_u0__abc_45749_n135;
  wire u1_u0__abc_45749_n136;
  wire u1_u0__abc_45749_n137;
  wire u1_u0__abc_45749_n139;
  wire u1_u0__abc_45749_n140;
  wire u1_u0__abc_45749_n141;
  wire u1_u0__abc_45749_n142;
  wire u1_u0__abc_45749_n144;
  wire u1_u0__abc_45749_n145;
  wire u1_u0__abc_45749_n146;
  wire u1_u0__abc_45749_n149;
  wire u1_u0__abc_45749_n150;
  wire u1_u0__abc_45749_n51;
  wire u1_u0__abc_45749_n52_1;
  wire u1_u0__abc_45749_n53_1;
  wire u1_u0__abc_45749_n54;
  wire u1_u0__abc_45749_n56_1;
  wire u1_u0__abc_45749_n57;
  wire u1_u0__abc_45749_n58;
  wire u1_u0__abc_45749_n60_1;
  wire u1_u0__abc_45749_n61;
  wire u1_u0__abc_45749_n62_1;
  wire u1_u0__abc_45749_n63_1;
  wire u1_u0__abc_45749_n65;
  wire u1_u0__abc_45749_n66;
  wire u1_u0__abc_45749_n67_1;
  wire u1_u0__abc_45749_n69;
  wire u1_u0__abc_45749_n70_1;
  wire u1_u0__abc_45749_n71_1;
  wire u1_u0__abc_45749_n72;
  wire u1_u0__abc_45749_n74_1;
  wire u1_u0__abc_45749_n75_1;
  wire u1_u0__abc_45749_n76;
  wire u1_u0__abc_45749_n78_1;
  wire u1_u0__abc_45749_n79_1;
  wire u1_u0__abc_45749_n80;
  wire u1_u0__abc_45749_n81;
  wire u1_u0__abc_45749_n82_1;
  wire u1_u0__abc_45749_n84;
  wire u1_u0__abc_45749_n85;
  wire u1_u0__abc_45749_n86;
  wire u1_u0__abc_45749_n88;
  wire u1_u0__abc_45749_n89;
  wire u1_u0__abc_45749_n90;
  wire u1_u0__abc_45749_n91;
  wire u1_u0__abc_45749_n93;
  wire u1_u0__abc_45749_n94;
  wire u1_u0__abc_45749_n95;
  wire u1_u0__abc_45749_n97;
  wire u1_u0__abc_45749_n98;
  wire u1_u0__abc_45749_n99;
  wire u1_u0_inc_next;
  wire u1_u0_out_r_0__FF_INPUT;
  wire u1_u0_out_r_10__FF_INPUT;
  wire u1_u0_out_r_11__FF_INPUT;
  wire u1_u0_out_r_12__FF_INPUT;
  wire u1_u0_out_r_1__FF_INPUT;
  wire u1_u0_out_r_2__FF_INPUT;
  wire u1_u0_out_r_3__FF_INPUT;
  wire u1_u0_out_r_4__FF_INPUT;
  wire u1_u0_out_r_5__FF_INPUT;
  wire u1_u0_out_r_6__FF_INPUT;
  wire u1_u0_out_r_7__FF_INPUT;
  wire u1_u0_out_r_8__FF_INPUT;
  wire u1_u0_out_r_9__FF_INPUT;
  wire u1_wb_write_go;
  wire u1_wr_cycle;
  wire u1_wr_hold;
  wire u2__abc_48153_n100;
  wire u2__abc_48153_n101;
  wire u2__abc_48153_n102;
  wire u2__abc_48153_n103;
  wire u2__abc_48153_n104;
  wire u2__abc_48153_n105;
  wire u2__abc_48153_n106;
  wire u2__abc_48153_n107;
  wire u2__abc_48153_n108;
  wire u2__abc_48153_n109;
  wire u2__abc_48153_n111;
  wire u2__abc_48153_n112;
  wire u2__abc_48153_n113;
  wire u2__abc_48153_n114;
  wire u2__abc_48153_n115;
  wire u2__abc_48153_n116;
  wire u2__abc_48153_n117;
  wire u2__abc_48153_n118;
  wire u2__abc_48153_n119;
  wire u2__abc_48153_n120;
  wire u2__abc_48153_n121;
  wire u2__abc_48153_n122;
  wire u2__abc_48153_n123;
  wire u2__abc_48153_n124;
  wire u2__abc_48153_n80;
  wire u2__abc_48153_n82_1;
  wire u2__abc_48153_n84_1;
  wire u2__abc_48153_n86;
  wire u2__abc_48153_n88_1;
  wire u2__abc_48153_n90;
  wire u2__abc_48153_n96;
  wire u2__abc_48153_n97;
  wire u2__abc_48153_n98;
  wire u2__abc_48153_n99;
  wire u2_bank_clr_0;
  wire u2_bank_clr_1;
  wire u2_bank_clr_2;
  wire u2_bank_clr_3;
  wire u2_bank_clr_4;
  wire u2_bank_clr_5;
  wire u2_bank_clr_all_0;
  wire u2_bank_clr_all_1;
  wire u2_bank_clr_all_2;
  wire u2_bank_clr_all_3;
  wire u2_bank_clr_all_4;
  wire u2_bank_clr_all_5;
  wire u2_bank_open_0;
  wire u2_bank_open_1;
  wire u2_bank_open_2;
  wire u2_bank_open_3;
  wire u2_bank_open_4;
  wire u2_bank_open_5;
  wire u2_bank_open_FF_INPUT;
  wire u2_bank_set_0;
  wire u2_bank_set_1;
  wire u2_bank_set_2;
  wire u2_bank_set_3;
  wire u2_bank_set_4;
  wire u2_bank_set_5;
  wire u2_row_same_0;
  wire u2_row_same_1;
  wire u2_row_same_2;
  wire u2_row_same_3;
  wire u2_row_same_4;
  wire u2_row_same_5;
  wire u2_row_same_FF_INPUT;
  wire u2_u0__abc_47660_n136;
  wire u2_u0__abc_47660_n137;
  wire u2_u0__abc_47660_n137_bF_buf0;
  wire u2_u0__abc_47660_n137_bF_buf1;
  wire u2_u0__abc_47660_n137_bF_buf2;
  wire u2_u0__abc_47660_n137_bF_buf3;
  wire u2_u0__abc_47660_n137_bF_buf4;
  wire u2_u0__abc_47660_n138;
  wire u2_u0__abc_47660_n139;
  wire u2_u0__abc_47660_n140;
  wire u2_u0__abc_47660_n141;
  wire u2_u0__abc_47660_n143;
  wire u2_u0__abc_47660_n144;
  wire u2_u0__abc_47660_n145;
  wire u2_u0__abc_47660_n146;
  wire u2_u0__abc_47660_n148;
  wire u2_u0__abc_47660_n149;
  wire u2_u0__abc_47660_n150;
  wire u2_u0__abc_47660_n151;
  wire u2_u0__abc_47660_n153;
  wire u2_u0__abc_47660_n154;
  wire u2_u0__abc_47660_n155;
  wire u2_u0__abc_47660_n156;
  wire u2_u0__abc_47660_n158;
  wire u2_u0__abc_47660_n159;
  wire u2_u0__abc_47660_n160;
  wire u2_u0__abc_47660_n161;
  wire u2_u0__abc_47660_n163;
  wire u2_u0__abc_47660_n164;
  wire u2_u0__abc_47660_n165;
  wire u2_u0__abc_47660_n166;
  wire u2_u0__abc_47660_n168;
  wire u2_u0__abc_47660_n169;
  wire u2_u0__abc_47660_n170;
  wire u2_u0__abc_47660_n171;
  wire u2_u0__abc_47660_n173;
  wire u2_u0__abc_47660_n174;
  wire u2_u0__abc_47660_n175;
  wire u2_u0__abc_47660_n176;
  wire u2_u0__abc_47660_n178;
  wire u2_u0__abc_47660_n179;
  wire u2_u0__abc_47660_n180;
  wire u2_u0__abc_47660_n181;
  wire u2_u0__abc_47660_n183;
  wire u2_u0__abc_47660_n184;
  wire u2_u0__abc_47660_n185;
  wire u2_u0__abc_47660_n186;
  wire u2_u0__abc_47660_n188;
  wire u2_u0__abc_47660_n189;
  wire u2_u0__abc_47660_n190;
  wire u2_u0__abc_47660_n191;
  wire u2_u0__abc_47660_n193;
  wire u2_u0__abc_47660_n194;
  wire u2_u0__abc_47660_n195;
  wire u2_u0__abc_47660_n196;
  wire u2_u0__abc_47660_n198;
  wire u2_u0__abc_47660_n199;
  wire u2_u0__abc_47660_n200;
  wire u2_u0__abc_47660_n201;
  wire u2_u0__abc_47660_n203;
  wire u2_u0__abc_47660_n204;
  wire u2_u0__abc_47660_n205;
  wire u2_u0__abc_47660_n206;
  wire u2_u0__abc_47660_n207;
  wire u2_u0__abc_47660_n208;
  wire u2_u0__abc_47660_n210;
  wire u2_u0__abc_47660_n211;
  wire u2_u0__abc_47660_n213;
  wire u2_u0__abc_47660_n214;
  wire u2_u0__abc_47660_n216;
  wire u2_u0__abc_47660_n217;
  wire u2_u0__abc_47660_n219;
  wire u2_u0__abc_47660_n220;
  wire u2_u0__abc_47660_n222;
  wire u2_u0__abc_47660_n223;
  wire u2_u0__abc_47660_n225;
  wire u2_u0__abc_47660_n226;
  wire u2_u0__abc_47660_n228;
  wire u2_u0__abc_47660_n229;
  wire u2_u0__abc_47660_n231;
  wire u2_u0__abc_47660_n232;
  wire u2_u0__abc_47660_n234;
  wire u2_u0__abc_47660_n235;
  wire u2_u0__abc_47660_n237;
  wire u2_u0__abc_47660_n238;
  wire u2_u0__abc_47660_n240;
  wire u2_u0__abc_47660_n241;
  wire u2_u0__abc_47660_n243;
  wire u2_u0__abc_47660_n244;
  wire u2_u0__abc_47660_n246;
  wire u2_u0__abc_47660_n247;
  wire u2_u0__abc_47660_n248;
  wire u2_u0__abc_47660_n249;
  wire u2_u0__abc_47660_n250;
  wire u2_u0__abc_47660_n251;
  wire u2_u0__abc_47660_n253;
  wire u2_u0__abc_47660_n254;
  wire u2_u0__abc_47660_n256;
  wire u2_u0__abc_47660_n257;
  wire u2_u0__abc_47660_n259;
  wire u2_u0__abc_47660_n260;
  wire u2_u0__abc_47660_n262;
  wire u2_u0__abc_47660_n263;
  wire u2_u0__abc_47660_n265;
  wire u2_u0__abc_47660_n266;
  wire u2_u0__abc_47660_n268;
  wire u2_u0__abc_47660_n269;
  wire u2_u0__abc_47660_n271;
  wire u2_u0__abc_47660_n272;
  wire u2_u0__abc_47660_n274;
  wire u2_u0__abc_47660_n275_1;
  wire u2_u0__abc_47660_n277;
  wire u2_u0__abc_47660_n278_1;
  wire u2_u0__abc_47660_n280;
  wire u2_u0__abc_47660_n281;
  wire u2_u0__abc_47660_n283_1;
  wire u2_u0__abc_47660_n284;
  wire u2_u0__abc_47660_n286_1;
  wire u2_u0__abc_47660_n287_1;
  wire u2_u0__abc_47660_n289;
  wire u2_u0__abc_47660_n290_1;
  wire u2_u0__abc_47660_n291;
  wire u2_u0__abc_47660_n292_1;
  wire u2_u0__abc_47660_n293;
  wire u2_u0__abc_47660_n295;
  wire u2_u0__abc_47660_n296_1;
  wire u2_u0__abc_47660_n298;
  wire u2_u0__abc_47660_n299;
  wire u2_u0__abc_47660_n301;
  wire u2_u0__abc_47660_n302;
  wire u2_u0__abc_47660_n304_1;
  wire u2_u0__abc_47660_n305;
  wire u2_u0__abc_47660_n305_1;
  wire u2_u0__abc_47660_n307;
  wire u2_u0__abc_47660_n308;
  wire u2_u0__abc_47660_n310;
  wire u2_u0__abc_47660_n311;
  wire u2_u0__abc_47660_n313;
  wire u2_u0__abc_47660_n314;
  wire u2_u0__abc_47660_n316;
  wire u2_u0__abc_47660_n317;
  wire u2_u0__abc_47660_n319;
  wire u2_u0__abc_47660_n320;
  wire u2_u0__abc_47660_n322;
  wire u2_u0__abc_47660_n323;
  wire u2_u0__abc_47660_n325;
  wire u2_u0__abc_47660_n326;
  wire u2_u0__abc_47660_n328;
  wire u2_u0__abc_47660_n329;
  wire u2_u0__abc_47660_n331;
  wire u2_u0__abc_47660_n332;
  wire u2_u0__abc_47660_n333;
  wire u2_u0__abc_47660_n334;
  wire u2_u0__abc_47660_n335;
  wire u2_u0__abc_47660_n336;
  wire u2_u0__abc_47660_n337;
  wire u2_u0__abc_47660_n338;
  wire u2_u0__abc_47660_n339;
  wire u2_u0__abc_47660_n340;
  wire u2_u0__abc_47660_n341;
  wire u2_u0__abc_47660_n342;
  wire u2_u0__abc_47660_n343;
  wire u2_u0__abc_47660_n344;
  wire u2_u0__abc_47660_n345;
  wire u2_u0__abc_47660_n346;
  wire u2_u0__abc_47660_n347;
  wire u2_u0__abc_47660_n348;
  wire u2_u0__abc_47660_n349;
  wire u2_u0__abc_47660_n350;
  wire u2_u0__abc_47660_n351;
  wire u2_u0__abc_47660_n352;
  wire u2_u0__abc_47660_n353;
  wire u2_u0__abc_47660_n354;
  wire u2_u0__abc_47660_n355;
  wire u2_u0__abc_47660_n356;
  wire u2_u0__abc_47660_n357;
  wire u2_u0__abc_47660_n358;
  wire u2_u0__abc_47660_n359;
  wire u2_u0__abc_47660_n360;
  wire u2_u0__abc_47660_n361;
  wire u2_u0__abc_47660_n362;
  wire u2_u0__abc_47660_n363;
  wire u2_u0__abc_47660_n364;
  wire u2_u0__abc_47660_n365;
  wire u2_u0__abc_47660_n366;
  wire u2_u0__abc_47660_n367;
  wire u2_u0__abc_47660_n368;
  wire u2_u0__abc_47660_n369;
  wire u2_u0__abc_47660_n370;
  wire u2_u0__abc_47660_n371;
  wire u2_u0__abc_47660_n372;
  wire u2_u0__abc_47660_n373;
  wire u2_u0__abc_47660_n374;
  wire u2_u0__abc_47660_n375;
  wire u2_u0__abc_47660_n376;
  wire u2_u0__abc_47660_n377;
  wire u2_u0__abc_47660_n378;
  wire u2_u0__abc_47660_n379;
  wire u2_u0__abc_47660_n380;
  wire u2_u0__abc_47660_n381;
  wire u2_u0__abc_47660_n382;
  wire u2_u0__abc_47660_n383;
  wire u2_u0__abc_47660_n384;
  wire u2_u0__abc_47660_n385;
  wire u2_u0__abc_47660_n386;
  wire u2_u0__abc_47660_n387;
  wire u2_u0__abc_47660_n388;
  wire u2_u0__abc_47660_n389;
  wire u2_u0__abc_47660_n390;
  wire u2_u0__abc_47660_n391;
  wire u2_u0__abc_47660_n392;
  wire u2_u0__abc_47660_n393;
  wire u2_u0__abc_47660_n394;
  wire u2_u0__abc_47660_n395;
  wire u2_u0__abc_47660_n396;
  wire u2_u0__abc_47660_n397;
  wire u2_u0__abc_47660_n398;
  wire u2_u0__abc_47660_n399;
  wire u2_u0__abc_47660_n400;
  wire u2_u0__abc_47660_n401;
  wire u2_u0__abc_47660_n402;
  wire u2_u0__abc_47660_n403;
  wire u2_u0__abc_47660_n404;
  wire u2_u0__abc_47660_n405;
  wire u2_u0__abc_47660_n406;
  wire u2_u0__abc_47660_n407;
  wire u2_u0__abc_47660_n408;
  wire u2_u0__abc_47660_n409;
  wire u2_u0__abc_47660_n410;
  wire u2_u0__abc_47660_n411;
  wire u2_u0__abc_47660_n412;
  wire u2_u0__abc_47660_n413;
  wire u2_u0__abc_47660_n414;
  wire u2_u0__abc_47660_n415;
  wire u2_u0__abc_47660_n416;
  wire u2_u0__abc_47660_n417;
  wire u2_u0__abc_47660_n418;
  wire u2_u0__abc_47660_n419;
  wire u2_u0__abc_47660_n420;
  wire u2_u0__abc_47660_n421;
  wire u2_u0__abc_47660_n422;
  wire u2_u0__abc_47660_n423;
  wire u2_u0__abc_47660_n424;
  wire u2_u0__abc_47660_n425;
  wire u2_u0__abc_47660_n426;
  wire u2_u0__abc_47660_n427;
  wire u2_u0__abc_47660_n428;
  wire u2_u0__abc_47660_n429;
  wire u2_u0__abc_47660_n430;
  wire u2_u0__abc_47660_n431;
  wire u2_u0__abc_47660_n432;
  wire u2_u0__abc_47660_n433;
  wire u2_u0__abc_47660_n434;
  wire u2_u0__abc_47660_n435;
  wire u2_u0__abc_47660_n436;
  wire u2_u0__abc_47660_n437;
  wire u2_u0__abc_47660_n438;
  wire u2_u0__abc_47660_n439;
  wire u2_u0__abc_47660_n440;
  wire u2_u0__abc_47660_n441;
  wire u2_u0__abc_47660_n442;
  wire u2_u0__abc_47660_n443;
  wire u2_u0__abc_47660_n444;
  wire u2_u0__abc_47660_n445;
  wire u2_u0__abc_47660_n446;
  wire u2_u0__abc_47660_n447;
  wire u2_u0__abc_47660_n448;
  wire u2_u0__abc_47660_n449;
  wire u2_u0__abc_47660_n450;
  wire u2_u0__abc_47660_n451;
  wire u2_u0__abc_47660_n452;
  wire u2_u0__abc_47660_n453;
  wire u2_u0__abc_47660_n454;
  wire u2_u0__abc_47660_n455;
  wire u2_u0__abc_47660_n456;
  wire u2_u0__abc_47660_n457;
  wire u2_u0__abc_47660_n458;
  wire u2_u0__abc_47660_n459;
  wire u2_u0__abc_47660_n460;
  wire u2_u0__abc_47660_n461;
  wire u2_u0__abc_47660_n462;
  wire u2_u0__abc_47660_n463;
  wire u2_u0__abc_47660_n464;
  wire u2_u0__abc_47660_n465;
  wire u2_u0__abc_47660_n466;
  wire u2_u0__abc_47660_n467;
  wire u2_u0__abc_47660_n468;
  wire u2_u0__abc_47660_n469;
  wire u2_u0__abc_47660_n470;
  wire u2_u0__abc_47660_n471;
  wire u2_u0__abc_47660_n472;
  wire u2_u0__abc_47660_n473;
  wire u2_u0__abc_47660_n474;
  wire u2_u0__abc_47660_n475;
  wire u2_u0__abc_47660_n476;
  wire u2_u0__abc_47660_n477;
  wire u2_u0__abc_47660_n478;
  wire u2_u0__abc_47660_n479;
  wire u2_u0__abc_47660_n480;
  wire u2_u0__abc_47660_n481;
  wire u2_u0__abc_47660_n482;
  wire u2_u0__abc_47660_n483;
  wire u2_u0__abc_47660_n484;
  wire u2_u0__abc_47660_n485;
  wire u2_u0__abc_47660_n486;
  wire u2_u0__abc_47660_n487;
  wire u2_u0__abc_47660_n488;
  wire u2_u0__abc_47660_n489;
  wire u2_u0__abc_47660_n490;
  wire u2_u0__abc_47660_n491;
  wire u2_u0__abc_47660_n492;
  wire u2_u0__abc_47660_n493;
  wire u2_u0__abc_47660_n494;
  wire u2_u0__abc_47660_n495;
  wire u2_u0__abc_47660_n496;
  wire u2_u0__abc_47660_n497;
  wire u2_u0__abc_47660_n498;
  wire u2_u0__abc_47660_n499;
  wire u2_u0__abc_47660_n500;
  wire u2_u0__abc_47660_n501;
  wire u2_u0__abc_47660_n502;
  wire u2_u0__abc_47660_n503;
  wire u2_u0__abc_47660_n504;
  wire u2_u0__abc_47660_n505;
  wire u2_u0__abc_47660_n506;
  wire u2_u0__abc_47660_n507;
  wire u2_u0__abc_47660_n508;
  wire u2_u0__abc_47660_n509;
  wire u2_u0__abc_47660_n510;
  wire u2_u0__abc_47660_n511;
  wire u2_u0__abc_47660_n512;
  wire u2_u0__abc_47660_n513;
  wire u2_u0__abc_47660_n514;
  wire u2_u0__abc_47660_n515;
  wire u2_u0__abc_47660_n516;
  wire u2_u0__abc_47660_n517;
  wire u2_u0__abc_47660_n518;
  wire u2_u0__abc_47660_n519;
  wire u2_u0__abc_47660_n520;
  wire u2_u0__abc_47660_n521;
  wire u2_u0__abc_47660_n522;
  wire u2_u0__abc_47660_n523;
  wire u2_u0__abc_47660_n524;
  wire u2_u0__abc_47660_n525;
  wire u2_u0__abc_47660_n526;
  wire u2_u0__abc_47660_n527;
  wire u2_u0__abc_47660_n528;
  wire u2_u0__abc_47660_n529;
  wire u2_u0__abc_47660_n530;
  wire u2_u0__abc_47660_n531;
  wire u2_u0__abc_47660_n532;
  wire u2_u0__abc_47660_n533;
  wire u2_u0__abc_47660_n534;
  wire u2_u0__abc_47660_n535;
  wire u2_u0__abc_47660_n536;
  wire u2_u0__abc_47660_n537;
  wire u2_u0__abc_47660_n538;
  wire u2_u0__abc_47660_n539;
  wire u2_u0__abc_47660_n540;
  wire u2_u0__abc_47660_n541;
  wire u2_u0__abc_47660_n542;
  wire u2_u0__abc_47660_n543;
  wire u2_u0__abc_47660_n544;
  wire u2_u0__abc_47660_n545;
  wire u2_u0__abc_47660_n546;
  wire u2_u0__abc_47660_n547;
  wire u2_u0__abc_47660_n548;
  wire u2_u0__abc_47660_n549;
  wire u2_u0__abc_47660_n550;
  wire u2_u0__abc_47660_n551;
  wire u2_u0__abc_47660_n552;
  wire u2_u0__abc_47660_n553;
  wire u2_u0__abc_47660_n554;
  wire u2_u0__abc_47660_n555;
  wire u2_u0__abc_47660_n556;
  wire u2_u0__abc_47660_n557;
  wire u2_u0__abc_47660_n558;
  wire u2_u0__abc_47660_n559;
  wire u2_u0__abc_47660_n560;
  wire u2_u0__abc_47660_n561;
  wire u2_u0__abc_47660_n562;
  wire u2_u0__abc_47660_n563;
  wire u2_u0__abc_47660_n564;
  wire u2_u0__abc_47660_n565;
  wire u2_u0__abc_47660_n566;
  wire u2_u0__abc_47660_n567;
  wire u2_u0__abc_47660_n568;
  wire u2_u0__abc_47660_n569;
  wire u2_u0__abc_47660_n570;
  wire u2_u0__abc_47660_n571;
  wire u2_u0__abc_47660_n572;
  wire u2_u0__abc_47660_n573;
  wire u2_u0__abc_47660_n574;
  wire u2_u0__abc_47660_n575;
  wire u2_u0__abc_47660_n576;
  wire u2_u0__abc_47660_n577;
  wire u2_u0__abc_47660_n578;
  wire u2_u0__abc_47660_n579;
  wire u2_u0__abc_47660_n580;
  wire u2_u0__abc_47660_n581;
  wire u2_u0__abc_47660_n582;
  wire u2_u0__abc_47660_n583;
  wire u2_u0__abc_47660_n584;
  wire u2_u0__abc_47660_n585;
  wire u2_u0__abc_47660_n586;
  wire u2_u0__abc_47660_n587;
  wire u2_u0__abc_47660_n588;
  wire u2_u0__abc_47660_n589;
  wire u2_u0__abc_47660_n590;
  wire u2_u0__abc_47660_n591;
  wire u2_u0__abc_47660_n592;
  wire u2_u0__abc_47660_n594;
  wire u2_u0__abc_47660_n595;
  wire u2_u0__abc_47660_n596;
  wire u2_u0__abc_47660_n597;
  wire u2_u0__abc_47660_n598;
  wire u2_u0__abc_47660_n599;
  wire u2_u0__abc_47660_n604;
  wire u2_u0__abc_47660_n605;
  wire u2_u0__abc_47660_n606;
  wire u2_u0__abc_47660_n607;
  wire u2_u0__abc_47660_n608;
  wire u2_u0__abc_47660_n610;
  wire u2_u0__abc_47660_n611;
  wire u2_u0__abc_47660_n612;
  wire u2_u0__abc_47660_n613;
  wire u2_u0__abc_47660_n614;
  wire u2_u0__abc_47660_n616;
  wire u2_u0__abc_47660_n617;
  wire u2_u0__abc_47660_n618;
  wire u2_u0__abc_47660_n619;
  wire u2_u0__abc_47660_n621;
  wire u2_u0__abc_47660_n622;
  wire u2_u0__abc_47660_n623;
  wire u2_u0__abc_47660_n624;
  wire u2_u0_b0_last_row_0_;
  wire u2_u0_b0_last_row_0__FF_INPUT;
  wire u2_u0_b0_last_row_10_;
  wire u2_u0_b0_last_row_10__FF_INPUT;
  wire u2_u0_b0_last_row_11_;
  wire u2_u0_b0_last_row_11__FF_INPUT;
  wire u2_u0_b0_last_row_12_;
  wire u2_u0_b0_last_row_12__FF_INPUT;
  wire u2_u0_b0_last_row_1_;
  wire u2_u0_b0_last_row_1__FF_INPUT;
  wire u2_u0_b0_last_row_2_;
  wire u2_u0_b0_last_row_2__FF_INPUT;
  wire u2_u0_b0_last_row_3_;
  wire u2_u0_b0_last_row_3__FF_INPUT;
  wire u2_u0_b0_last_row_4_;
  wire u2_u0_b0_last_row_4__FF_INPUT;
  wire u2_u0_b0_last_row_5_;
  wire u2_u0_b0_last_row_5__FF_INPUT;
  wire u2_u0_b0_last_row_6_;
  wire u2_u0_b0_last_row_6__FF_INPUT;
  wire u2_u0_b0_last_row_7_;
  wire u2_u0_b0_last_row_7__FF_INPUT;
  wire u2_u0_b0_last_row_8_;
  wire u2_u0_b0_last_row_8__FF_INPUT;
  wire u2_u0_b0_last_row_9_;
  wire u2_u0_b0_last_row_9__FF_INPUT;
  wire u2_u0_b1_last_row_0_;
  wire u2_u0_b1_last_row_0__FF_INPUT;
  wire u2_u0_b1_last_row_10_;
  wire u2_u0_b1_last_row_10__FF_INPUT;
  wire u2_u0_b1_last_row_11_;
  wire u2_u0_b1_last_row_11__FF_INPUT;
  wire u2_u0_b1_last_row_12_;
  wire u2_u0_b1_last_row_12__FF_INPUT;
  wire u2_u0_b1_last_row_1_;
  wire u2_u0_b1_last_row_1__FF_INPUT;
  wire u2_u0_b1_last_row_2_;
  wire u2_u0_b1_last_row_2__FF_INPUT;
  wire u2_u0_b1_last_row_3_;
  wire u2_u0_b1_last_row_3__FF_INPUT;
  wire u2_u0_b1_last_row_4_;
  wire u2_u0_b1_last_row_4__FF_INPUT;
  wire u2_u0_b1_last_row_5_;
  wire u2_u0_b1_last_row_5__FF_INPUT;
  wire u2_u0_b1_last_row_6_;
  wire u2_u0_b1_last_row_6__FF_INPUT;
  wire u2_u0_b1_last_row_7_;
  wire u2_u0_b1_last_row_7__FF_INPUT;
  wire u2_u0_b1_last_row_8_;
  wire u2_u0_b1_last_row_8__FF_INPUT;
  wire u2_u0_b1_last_row_9_;
  wire u2_u0_b1_last_row_9__FF_INPUT;
  wire u2_u0_b2_last_row_0_;
  wire u2_u0_b2_last_row_0__FF_INPUT;
  wire u2_u0_b2_last_row_10_;
  wire u2_u0_b2_last_row_10__FF_INPUT;
  wire u2_u0_b2_last_row_11_;
  wire u2_u0_b2_last_row_11__FF_INPUT;
  wire u2_u0_b2_last_row_12_;
  wire u2_u0_b2_last_row_12__FF_INPUT;
  wire u2_u0_b2_last_row_1_;
  wire u2_u0_b2_last_row_1__FF_INPUT;
  wire u2_u0_b2_last_row_2_;
  wire u2_u0_b2_last_row_2__FF_INPUT;
  wire u2_u0_b2_last_row_3_;
  wire u2_u0_b2_last_row_3__FF_INPUT;
  wire u2_u0_b2_last_row_4_;
  wire u2_u0_b2_last_row_4__FF_INPUT;
  wire u2_u0_b2_last_row_5_;
  wire u2_u0_b2_last_row_5__FF_INPUT;
  wire u2_u0_b2_last_row_6_;
  wire u2_u0_b2_last_row_6__FF_INPUT;
  wire u2_u0_b2_last_row_7_;
  wire u2_u0_b2_last_row_7__FF_INPUT;
  wire u2_u0_b2_last_row_8_;
  wire u2_u0_b2_last_row_8__FF_INPUT;
  wire u2_u0_b2_last_row_9_;
  wire u2_u0_b2_last_row_9__FF_INPUT;
  wire u2_u0_b3_last_row_0_;
  wire u2_u0_b3_last_row_0__FF_INPUT;
  wire u2_u0_b3_last_row_10_;
  wire u2_u0_b3_last_row_10__FF_INPUT;
  wire u2_u0_b3_last_row_11_;
  wire u2_u0_b3_last_row_11__FF_INPUT;
  wire u2_u0_b3_last_row_12_;
  wire u2_u0_b3_last_row_12__FF_INPUT;
  wire u2_u0_b3_last_row_1_;
  wire u2_u0_b3_last_row_1__FF_INPUT;
  wire u2_u0_b3_last_row_2_;
  wire u2_u0_b3_last_row_2__FF_INPUT;
  wire u2_u0_b3_last_row_3_;
  wire u2_u0_b3_last_row_3__FF_INPUT;
  wire u2_u0_b3_last_row_4_;
  wire u2_u0_b3_last_row_4__FF_INPUT;
  wire u2_u0_b3_last_row_5_;
  wire u2_u0_b3_last_row_5__FF_INPUT;
  wire u2_u0_b3_last_row_6_;
  wire u2_u0_b3_last_row_6__FF_INPUT;
  wire u2_u0_b3_last_row_7_;
  wire u2_u0_b3_last_row_7__FF_INPUT;
  wire u2_u0_b3_last_row_8_;
  wire u2_u0_b3_last_row_8__FF_INPUT;
  wire u2_u0_b3_last_row_9_;
  wire u2_u0_b3_last_row_9__FF_INPUT;
  wire u2_u0_bank0_open;
  wire u2_u0_bank0_open_FF_INPUT;
  wire u2_u0_bank1_open;
  wire u2_u0_bank1_open_FF_INPUT;
  wire u2_u0_bank2_open;
  wire u2_u0_bank2_open_FF_INPUT;
  wire u2_u0_bank3_open;
  wire u2_u0_bank3_open_FF_INPUT;
  wire u2_u1__abc_47660_n136;
  wire u2_u1__abc_47660_n137;
  wire u2_u1__abc_47660_n137_bF_buf0;
  wire u2_u1__abc_47660_n137_bF_buf1;
  wire u2_u1__abc_47660_n137_bF_buf2;
  wire u2_u1__abc_47660_n137_bF_buf3;
  wire u2_u1__abc_47660_n137_bF_buf4;
  wire u2_u1__abc_47660_n138;
  wire u2_u1__abc_47660_n139;
  wire u2_u1__abc_47660_n140;
  wire u2_u1__abc_47660_n141;
  wire u2_u1__abc_47660_n143;
  wire u2_u1__abc_47660_n144;
  wire u2_u1__abc_47660_n145;
  wire u2_u1__abc_47660_n146;
  wire u2_u1__abc_47660_n148;
  wire u2_u1__abc_47660_n149;
  wire u2_u1__abc_47660_n150;
  wire u2_u1__abc_47660_n151;
  wire u2_u1__abc_47660_n153;
  wire u2_u1__abc_47660_n154;
  wire u2_u1__abc_47660_n155;
  wire u2_u1__abc_47660_n156;
  wire u2_u1__abc_47660_n158;
  wire u2_u1__abc_47660_n159;
  wire u2_u1__abc_47660_n160;
  wire u2_u1__abc_47660_n161;
  wire u2_u1__abc_47660_n163;
  wire u2_u1__abc_47660_n164;
  wire u2_u1__abc_47660_n165;
  wire u2_u1__abc_47660_n166;
  wire u2_u1__abc_47660_n168;
  wire u2_u1__abc_47660_n169;
  wire u2_u1__abc_47660_n170;
  wire u2_u1__abc_47660_n171;
  wire u2_u1__abc_47660_n173;
  wire u2_u1__abc_47660_n174;
  wire u2_u1__abc_47660_n175;
  wire u2_u1__abc_47660_n176;
  wire u2_u1__abc_47660_n178;
  wire u2_u1__abc_47660_n179;
  wire u2_u1__abc_47660_n180;
  wire u2_u1__abc_47660_n181;
  wire u2_u1__abc_47660_n183;
  wire u2_u1__abc_47660_n184;
  wire u2_u1__abc_47660_n185;
  wire u2_u1__abc_47660_n186;
  wire u2_u1__abc_47660_n188;
  wire u2_u1__abc_47660_n189;
  wire u2_u1__abc_47660_n190;
  wire u2_u1__abc_47660_n191;
  wire u2_u1__abc_47660_n193;
  wire u2_u1__abc_47660_n194;
  wire u2_u1__abc_47660_n195;
  wire u2_u1__abc_47660_n196;
  wire u2_u1__abc_47660_n198;
  wire u2_u1__abc_47660_n199;
  wire u2_u1__abc_47660_n200;
  wire u2_u1__abc_47660_n201;
  wire u2_u1__abc_47660_n203;
  wire u2_u1__abc_47660_n204;
  wire u2_u1__abc_47660_n205;
  wire u2_u1__abc_47660_n206;
  wire u2_u1__abc_47660_n207;
  wire u2_u1__abc_47660_n208;
  wire u2_u1__abc_47660_n210;
  wire u2_u1__abc_47660_n211;
  wire u2_u1__abc_47660_n213;
  wire u2_u1__abc_47660_n214;
  wire u2_u1__abc_47660_n216;
  wire u2_u1__abc_47660_n217;
  wire u2_u1__abc_47660_n219;
  wire u2_u1__abc_47660_n220;
  wire u2_u1__abc_47660_n222;
  wire u2_u1__abc_47660_n223;
  wire u2_u1__abc_47660_n225;
  wire u2_u1__abc_47660_n226;
  wire u2_u1__abc_47660_n228;
  wire u2_u1__abc_47660_n229;
  wire u2_u1__abc_47660_n231;
  wire u2_u1__abc_47660_n232;
  wire u2_u1__abc_47660_n234;
  wire u2_u1__abc_47660_n235;
  wire u2_u1__abc_47660_n237;
  wire u2_u1__abc_47660_n238;
  wire u2_u1__abc_47660_n240;
  wire u2_u1__abc_47660_n241;
  wire u2_u1__abc_47660_n243;
  wire u2_u1__abc_47660_n244;
  wire u2_u1__abc_47660_n246;
  wire u2_u1__abc_47660_n247;
  wire u2_u1__abc_47660_n248;
  wire u2_u1__abc_47660_n249;
  wire u2_u1__abc_47660_n250;
  wire u2_u1__abc_47660_n251;
  wire u2_u1__abc_47660_n253;
  wire u2_u1__abc_47660_n254;
  wire u2_u1__abc_47660_n256;
  wire u2_u1__abc_47660_n257;
  wire u2_u1__abc_47660_n259;
  wire u2_u1__abc_47660_n260;
  wire u2_u1__abc_47660_n262;
  wire u2_u1__abc_47660_n263;
  wire u2_u1__abc_47660_n265;
  wire u2_u1__abc_47660_n266;
  wire u2_u1__abc_47660_n268;
  wire u2_u1__abc_47660_n269;
  wire u2_u1__abc_47660_n271;
  wire u2_u1__abc_47660_n272;
  wire u2_u1__abc_47660_n274;
  wire u2_u1__abc_47660_n275_1;
  wire u2_u1__abc_47660_n277;
  wire u2_u1__abc_47660_n278_1;
  wire u2_u1__abc_47660_n280;
  wire u2_u1__abc_47660_n281;
  wire u2_u1__abc_47660_n283_1;
  wire u2_u1__abc_47660_n284;
  wire u2_u1__abc_47660_n286_1;
  wire u2_u1__abc_47660_n287_1;
  wire u2_u1__abc_47660_n289;
  wire u2_u1__abc_47660_n290_1;
  wire u2_u1__abc_47660_n291;
  wire u2_u1__abc_47660_n292_1;
  wire u2_u1__abc_47660_n293;
  wire u2_u1__abc_47660_n295;
  wire u2_u1__abc_47660_n296_1;
  wire u2_u1__abc_47660_n298;
  wire u2_u1__abc_47660_n299;
  wire u2_u1__abc_47660_n301;
  wire u2_u1__abc_47660_n302;
  wire u2_u1__abc_47660_n304_1;
  wire u2_u1__abc_47660_n305;
  wire u2_u1__abc_47660_n305_1;
  wire u2_u1__abc_47660_n307;
  wire u2_u1__abc_47660_n308;
  wire u2_u1__abc_47660_n310;
  wire u2_u1__abc_47660_n311;
  wire u2_u1__abc_47660_n313;
  wire u2_u1__abc_47660_n314;
  wire u2_u1__abc_47660_n316;
  wire u2_u1__abc_47660_n317;
  wire u2_u1__abc_47660_n319;
  wire u2_u1__abc_47660_n320;
  wire u2_u1__abc_47660_n322;
  wire u2_u1__abc_47660_n323;
  wire u2_u1__abc_47660_n325;
  wire u2_u1__abc_47660_n326;
  wire u2_u1__abc_47660_n328;
  wire u2_u1__abc_47660_n329;
  wire u2_u1__abc_47660_n331;
  wire u2_u1__abc_47660_n332;
  wire u2_u1__abc_47660_n333;
  wire u2_u1__abc_47660_n334;
  wire u2_u1__abc_47660_n335;
  wire u2_u1__abc_47660_n336;
  wire u2_u1__abc_47660_n337;
  wire u2_u1__abc_47660_n338;
  wire u2_u1__abc_47660_n339;
  wire u2_u1__abc_47660_n340;
  wire u2_u1__abc_47660_n341;
  wire u2_u1__abc_47660_n342;
  wire u2_u1__abc_47660_n343;
  wire u2_u1__abc_47660_n344;
  wire u2_u1__abc_47660_n345;
  wire u2_u1__abc_47660_n346;
  wire u2_u1__abc_47660_n347;
  wire u2_u1__abc_47660_n348;
  wire u2_u1__abc_47660_n349;
  wire u2_u1__abc_47660_n350;
  wire u2_u1__abc_47660_n351;
  wire u2_u1__abc_47660_n352;
  wire u2_u1__abc_47660_n353;
  wire u2_u1__abc_47660_n354;
  wire u2_u1__abc_47660_n355;
  wire u2_u1__abc_47660_n356;
  wire u2_u1__abc_47660_n357;
  wire u2_u1__abc_47660_n358;
  wire u2_u1__abc_47660_n359;
  wire u2_u1__abc_47660_n360;
  wire u2_u1__abc_47660_n361;
  wire u2_u1__abc_47660_n362;
  wire u2_u1__abc_47660_n363;
  wire u2_u1__abc_47660_n364;
  wire u2_u1__abc_47660_n365;
  wire u2_u1__abc_47660_n366;
  wire u2_u1__abc_47660_n367;
  wire u2_u1__abc_47660_n368;
  wire u2_u1__abc_47660_n369;
  wire u2_u1__abc_47660_n370;
  wire u2_u1__abc_47660_n371;
  wire u2_u1__abc_47660_n372;
  wire u2_u1__abc_47660_n373;
  wire u2_u1__abc_47660_n374;
  wire u2_u1__abc_47660_n375;
  wire u2_u1__abc_47660_n376;
  wire u2_u1__abc_47660_n377;
  wire u2_u1__abc_47660_n378;
  wire u2_u1__abc_47660_n379;
  wire u2_u1__abc_47660_n380;
  wire u2_u1__abc_47660_n381;
  wire u2_u1__abc_47660_n382;
  wire u2_u1__abc_47660_n383;
  wire u2_u1__abc_47660_n384;
  wire u2_u1__abc_47660_n385;
  wire u2_u1__abc_47660_n386;
  wire u2_u1__abc_47660_n387;
  wire u2_u1__abc_47660_n388;
  wire u2_u1__abc_47660_n389;
  wire u2_u1__abc_47660_n390;
  wire u2_u1__abc_47660_n391;
  wire u2_u1__abc_47660_n392;
  wire u2_u1__abc_47660_n393;
  wire u2_u1__abc_47660_n394;
  wire u2_u1__abc_47660_n395;
  wire u2_u1__abc_47660_n396;
  wire u2_u1__abc_47660_n397;
  wire u2_u1__abc_47660_n398;
  wire u2_u1__abc_47660_n399;
  wire u2_u1__abc_47660_n400;
  wire u2_u1__abc_47660_n401;
  wire u2_u1__abc_47660_n402;
  wire u2_u1__abc_47660_n403;
  wire u2_u1__abc_47660_n404;
  wire u2_u1__abc_47660_n405;
  wire u2_u1__abc_47660_n406;
  wire u2_u1__abc_47660_n407;
  wire u2_u1__abc_47660_n408;
  wire u2_u1__abc_47660_n409;
  wire u2_u1__abc_47660_n410;
  wire u2_u1__abc_47660_n411;
  wire u2_u1__abc_47660_n412;
  wire u2_u1__abc_47660_n413;
  wire u2_u1__abc_47660_n414;
  wire u2_u1__abc_47660_n415;
  wire u2_u1__abc_47660_n416;
  wire u2_u1__abc_47660_n417;
  wire u2_u1__abc_47660_n418;
  wire u2_u1__abc_47660_n419;
  wire u2_u1__abc_47660_n420;
  wire u2_u1__abc_47660_n421;
  wire u2_u1__abc_47660_n422;
  wire u2_u1__abc_47660_n423;
  wire u2_u1__abc_47660_n424;
  wire u2_u1__abc_47660_n425;
  wire u2_u1__abc_47660_n426;
  wire u2_u1__abc_47660_n427;
  wire u2_u1__abc_47660_n428;
  wire u2_u1__abc_47660_n429;
  wire u2_u1__abc_47660_n430;
  wire u2_u1__abc_47660_n431;
  wire u2_u1__abc_47660_n432;
  wire u2_u1__abc_47660_n433;
  wire u2_u1__abc_47660_n434;
  wire u2_u1__abc_47660_n435;
  wire u2_u1__abc_47660_n436;
  wire u2_u1__abc_47660_n437;
  wire u2_u1__abc_47660_n438;
  wire u2_u1__abc_47660_n439;
  wire u2_u1__abc_47660_n440;
  wire u2_u1__abc_47660_n441;
  wire u2_u1__abc_47660_n442;
  wire u2_u1__abc_47660_n443;
  wire u2_u1__abc_47660_n444;
  wire u2_u1__abc_47660_n445;
  wire u2_u1__abc_47660_n446;
  wire u2_u1__abc_47660_n447;
  wire u2_u1__abc_47660_n448;
  wire u2_u1__abc_47660_n449;
  wire u2_u1__abc_47660_n450;
  wire u2_u1__abc_47660_n451;
  wire u2_u1__abc_47660_n452;
  wire u2_u1__abc_47660_n453;
  wire u2_u1__abc_47660_n454;
  wire u2_u1__abc_47660_n455;
  wire u2_u1__abc_47660_n456;
  wire u2_u1__abc_47660_n457;
  wire u2_u1__abc_47660_n458;
  wire u2_u1__abc_47660_n459;
  wire u2_u1__abc_47660_n460;
  wire u2_u1__abc_47660_n461;
  wire u2_u1__abc_47660_n462;
  wire u2_u1__abc_47660_n463;
  wire u2_u1__abc_47660_n464;
  wire u2_u1__abc_47660_n465;
  wire u2_u1__abc_47660_n466;
  wire u2_u1__abc_47660_n467;
  wire u2_u1__abc_47660_n468;
  wire u2_u1__abc_47660_n469;
  wire u2_u1__abc_47660_n470;
  wire u2_u1__abc_47660_n471;
  wire u2_u1__abc_47660_n472;
  wire u2_u1__abc_47660_n473;
  wire u2_u1__abc_47660_n474;
  wire u2_u1__abc_47660_n475;
  wire u2_u1__abc_47660_n476;
  wire u2_u1__abc_47660_n477;
  wire u2_u1__abc_47660_n478;
  wire u2_u1__abc_47660_n479;
  wire u2_u1__abc_47660_n480;
  wire u2_u1__abc_47660_n481;
  wire u2_u1__abc_47660_n482;
  wire u2_u1__abc_47660_n483;
  wire u2_u1__abc_47660_n484;
  wire u2_u1__abc_47660_n485;
  wire u2_u1__abc_47660_n486;
  wire u2_u1__abc_47660_n487;
  wire u2_u1__abc_47660_n488;
  wire u2_u1__abc_47660_n489;
  wire u2_u1__abc_47660_n490;
  wire u2_u1__abc_47660_n491;
  wire u2_u1__abc_47660_n492;
  wire u2_u1__abc_47660_n493;
  wire u2_u1__abc_47660_n494;
  wire u2_u1__abc_47660_n495;
  wire u2_u1__abc_47660_n496;
  wire u2_u1__abc_47660_n497;
  wire u2_u1__abc_47660_n498;
  wire u2_u1__abc_47660_n499;
  wire u2_u1__abc_47660_n500;
  wire u2_u1__abc_47660_n501;
  wire u2_u1__abc_47660_n502;
  wire u2_u1__abc_47660_n503;
  wire u2_u1__abc_47660_n504;
  wire u2_u1__abc_47660_n505;
  wire u2_u1__abc_47660_n506;
  wire u2_u1__abc_47660_n507;
  wire u2_u1__abc_47660_n508;
  wire u2_u1__abc_47660_n509;
  wire u2_u1__abc_47660_n510;
  wire u2_u1__abc_47660_n511;
  wire u2_u1__abc_47660_n512;
  wire u2_u1__abc_47660_n513;
  wire u2_u1__abc_47660_n514;
  wire u2_u1__abc_47660_n515;
  wire u2_u1__abc_47660_n516;
  wire u2_u1__abc_47660_n517;
  wire u2_u1__abc_47660_n518;
  wire u2_u1__abc_47660_n519;
  wire u2_u1__abc_47660_n520;
  wire u2_u1__abc_47660_n521;
  wire u2_u1__abc_47660_n522;
  wire u2_u1__abc_47660_n523;
  wire u2_u1__abc_47660_n524;
  wire u2_u1__abc_47660_n525;
  wire u2_u1__abc_47660_n526;
  wire u2_u1__abc_47660_n527;
  wire u2_u1__abc_47660_n528;
  wire u2_u1__abc_47660_n529;
  wire u2_u1__abc_47660_n530;
  wire u2_u1__abc_47660_n531;
  wire u2_u1__abc_47660_n532;
  wire u2_u1__abc_47660_n533;
  wire u2_u1__abc_47660_n534;
  wire u2_u1__abc_47660_n535;
  wire u2_u1__abc_47660_n536;
  wire u2_u1__abc_47660_n537;
  wire u2_u1__abc_47660_n538;
  wire u2_u1__abc_47660_n539;
  wire u2_u1__abc_47660_n540;
  wire u2_u1__abc_47660_n541;
  wire u2_u1__abc_47660_n542;
  wire u2_u1__abc_47660_n543;
  wire u2_u1__abc_47660_n544;
  wire u2_u1__abc_47660_n545;
  wire u2_u1__abc_47660_n546;
  wire u2_u1__abc_47660_n547;
  wire u2_u1__abc_47660_n548;
  wire u2_u1__abc_47660_n549;
  wire u2_u1__abc_47660_n550;
  wire u2_u1__abc_47660_n551;
  wire u2_u1__abc_47660_n552;
  wire u2_u1__abc_47660_n553;
  wire u2_u1__abc_47660_n554;
  wire u2_u1__abc_47660_n555;
  wire u2_u1__abc_47660_n556;
  wire u2_u1__abc_47660_n557;
  wire u2_u1__abc_47660_n558;
  wire u2_u1__abc_47660_n559;
  wire u2_u1__abc_47660_n560;
  wire u2_u1__abc_47660_n561;
  wire u2_u1__abc_47660_n562;
  wire u2_u1__abc_47660_n563;
  wire u2_u1__abc_47660_n564;
  wire u2_u1__abc_47660_n565;
  wire u2_u1__abc_47660_n566;
  wire u2_u1__abc_47660_n567;
  wire u2_u1__abc_47660_n568;
  wire u2_u1__abc_47660_n569;
  wire u2_u1__abc_47660_n570;
  wire u2_u1__abc_47660_n571;
  wire u2_u1__abc_47660_n572;
  wire u2_u1__abc_47660_n573;
  wire u2_u1__abc_47660_n574;
  wire u2_u1__abc_47660_n575;
  wire u2_u1__abc_47660_n576;
  wire u2_u1__abc_47660_n577;
  wire u2_u1__abc_47660_n578;
  wire u2_u1__abc_47660_n579;
  wire u2_u1__abc_47660_n580;
  wire u2_u1__abc_47660_n581;
  wire u2_u1__abc_47660_n582;
  wire u2_u1__abc_47660_n583;
  wire u2_u1__abc_47660_n584;
  wire u2_u1__abc_47660_n585;
  wire u2_u1__abc_47660_n586;
  wire u2_u1__abc_47660_n587;
  wire u2_u1__abc_47660_n588;
  wire u2_u1__abc_47660_n589;
  wire u2_u1__abc_47660_n590;
  wire u2_u1__abc_47660_n591;
  wire u2_u1__abc_47660_n592;
  wire u2_u1__abc_47660_n594;
  wire u2_u1__abc_47660_n595;
  wire u2_u1__abc_47660_n596;
  wire u2_u1__abc_47660_n597;
  wire u2_u1__abc_47660_n598;
  wire u2_u1__abc_47660_n599;
  wire u2_u1__abc_47660_n604;
  wire u2_u1__abc_47660_n605;
  wire u2_u1__abc_47660_n606;
  wire u2_u1__abc_47660_n607;
  wire u2_u1__abc_47660_n608;
  wire u2_u1__abc_47660_n610;
  wire u2_u1__abc_47660_n611;
  wire u2_u1__abc_47660_n612;
  wire u2_u1__abc_47660_n613;
  wire u2_u1__abc_47660_n614;
  wire u2_u1__abc_47660_n616;
  wire u2_u1__abc_47660_n617;
  wire u2_u1__abc_47660_n618;
  wire u2_u1__abc_47660_n619;
  wire u2_u1__abc_47660_n621;
  wire u2_u1__abc_47660_n622;
  wire u2_u1__abc_47660_n623;
  wire u2_u1__abc_47660_n624;
  wire u2_u1_b0_last_row_0_;
  wire u2_u1_b0_last_row_0__FF_INPUT;
  wire u2_u1_b0_last_row_10_;
  wire u2_u1_b0_last_row_10__FF_INPUT;
  wire u2_u1_b0_last_row_11_;
  wire u2_u1_b0_last_row_11__FF_INPUT;
  wire u2_u1_b0_last_row_12_;
  wire u2_u1_b0_last_row_12__FF_INPUT;
  wire u2_u1_b0_last_row_1_;
  wire u2_u1_b0_last_row_1__FF_INPUT;
  wire u2_u1_b0_last_row_2_;
  wire u2_u1_b0_last_row_2__FF_INPUT;
  wire u2_u1_b0_last_row_3_;
  wire u2_u1_b0_last_row_3__FF_INPUT;
  wire u2_u1_b0_last_row_4_;
  wire u2_u1_b0_last_row_4__FF_INPUT;
  wire u2_u1_b0_last_row_5_;
  wire u2_u1_b0_last_row_5__FF_INPUT;
  wire u2_u1_b0_last_row_6_;
  wire u2_u1_b0_last_row_6__FF_INPUT;
  wire u2_u1_b0_last_row_7_;
  wire u2_u1_b0_last_row_7__FF_INPUT;
  wire u2_u1_b0_last_row_8_;
  wire u2_u1_b0_last_row_8__FF_INPUT;
  wire u2_u1_b0_last_row_9_;
  wire u2_u1_b0_last_row_9__FF_INPUT;
  wire u2_u1_b1_last_row_0_;
  wire u2_u1_b1_last_row_0__FF_INPUT;
  wire u2_u1_b1_last_row_10_;
  wire u2_u1_b1_last_row_10__FF_INPUT;
  wire u2_u1_b1_last_row_11_;
  wire u2_u1_b1_last_row_11__FF_INPUT;
  wire u2_u1_b1_last_row_12_;
  wire u2_u1_b1_last_row_12__FF_INPUT;
  wire u2_u1_b1_last_row_1_;
  wire u2_u1_b1_last_row_1__FF_INPUT;
  wire u2_u1_b1_last_row_2_;
  wire u2_u1_b1_last_row_2__FF_INPUT;
  wire u2_u1_b1_last_row_3_;
  wire u2_u1_b1_last_row_3__FF_INPUT;
  wire u2_u1_b1_last_row_4_;
  wire u2_u1_b1_last_row_4__FF_INPUT;
  wire u2_u1_b1_last_row_5_;
  wire u2_u1_b1_last_row_5__FF_INPUT;
  wire u2_u1_b1_last_row_6_;
  wire u2_u1_b1_last_row_6__FF_INPUT;
  wire u2_u1_b1_last_row_7_;
  wire u2_u1_b1_last_row_7__FF_INPUT;
  wire u2_u1_b1_last_row_8_;
  wire u2_u1_b1_last_row_8__FF_INPUT;
  wire u2_u1_b1_last_row_9_;
  wire u2_u1_b1_last_row_9__FF_INPUT;
  wire u2_u1_b2_last_row_0_;
  wire u2_u1_b2_last_row_0__FF_INPUT;
  wire u2_u1_b2_last_row_10_;
  wire u2_u1_b2_last_row_10__FF_INPUT;
  wire u2_u1_b2_last_row_11_;
  wire u2_u1_b2_last_row_11__FF_INPUT;
  wire u2_u1_b2_last_row_12_;
  wire u2_u1_b2_last_row_12__FF_INPUT;
  wire u2_u1_b2_last_row_1_;
  wire u2_u1_b2_last_row_1__FF_INPUT;
  wire u2_u1_b2_last_row_2_;
  wire u2_u1_b2_last_row_2__FF_INPUT;
  wire u2_u1_b2_last_row_3_;
  wire u2_u1_b2_last_row_3__FF_INPUT;
  wire u2_u1_b2_last_row_4_;
  wire u2_u1_b2_last_row_4__FF_INPUT;
  wire u2_u1_b2_last_row_5_;
  wire u2_u1_b2_last_row_5__FF_INPUT;
  wire u2_u1_b2_last_row_6_;
  wire u2_u1_b2_last_row_6__FF_INPUT;
  wire u2_u1_b2_last_row_7_;
  wire u2_u1_b2_last_row_7__FF_INPUT;
  wire u2_u1_b2_last_row_8_;
  wire u2_u1_b2_last_row_8__FF_INPUT;
  wire u2_u1_b2_last_row_9_;
  wire u2_u1_b2_last_row_9__FF_INPUT;
  wire u2_u1_b3_last_row_0_;
  wire u2_u1_b3_last_row_0__FF_INPUT;
  wire u2_u1_b3_last_row_10_;
  wire u2_u1_b3_last_row_10__FF_INPUT;
  wire u2_u1_b3_last_row_11_;
  wire u2_u1_b3_last_row_11__FF_INPUT;
  wire u2_u1_b3_last_row_12_;
  wire u2_u1_b3_last_row_12__FF_INPUT;
  wire u2_u1_b3_last_row_1_;
  wire u2_u1_b3_last_row_1__FF_INPUT;
  wire u2_u1_b3_last_row_2_;
  wire u2_u1_b3_last_row_2__FF_INPUT;
  wire u2_u1_b3_last_row_3_;
  wire u2_u1_b3_last_row_3__FF_INPUT;
  wire u2_u1_b3_last_row_4_;
  wire u2_u1_b3_last_row_4__FF_INPUT;
  wire u2_u1_b3_last_row_5_;
  wire u2_u1_b3_last_row_5__FF_INPUT;
  wire u2_u1_b3_last_row_6_;
  wire u2_u1_b3_last_row_6__FF_INPUT;
  wire u2_u1_b3_last_row_7_;
  wire u2_u1_b3_last_row_7__FF_INPUT;
  wire u2_u1_b3_last_row_8_;
  wire u2_u1_b3_last_row_8__FF_INPUT;
  wire u2_u1_b3_last_row_9_;
  wire u2_u1_b3_last_row_9__FF_INPUT;
  wire u2_u1_bank0_open;
  wire u2_u1_bank0_open_FF_INPUT;
  wire u2_u1_bank1_open;
  wire u2_u1_bank1_open_FF_INPUT;
  wire u2_u1_bank2_open;
  wire u2_u1_bank2_open_FF_INPUT;
  wire u2_u1_bank3_open;
  wire u2_u1_bank3_open_FF_INPUT;
  wire u2_u2__abc_47660_n136;
  wire u2_u2__abc_47660_n137;
  wire u2_u2__abc_47660_n137_bF_buf0;
  wire u2_u2__abc_47660_n137_bF_buf1;
  wire u2_u2__abc_47660_n137_bF_buf2;
  wire u2_u2__abc_47660_n137_bF_buf3;
  wire u2_u2__abc_47660_n137_bF_buf4;
  wire u2_u2__abc_47660_n138;
  wire u2_u2__abc_47660_n139;
  wire u2_u2__abc_47660_n140;
  wire u2_u2__abc_47660_n141;
  wire u2_u2__abc_47660_n143;
  wire u2_u2__abc_47660_n144;
  wire u2_u2__abc_47660_n145;
  wire u2_u2__abc_47660_n146;
  wire u2_u2__abc_47660_n148;
  wire u2_u2__abc_47660_n149;
  wire u2_u2__abc_47660_n150;
  wire u2_u2__abc_47660_n151;
  wire u2_u2__abc_47660_n153;
  wire u2_u2__abc_47660_n154;
  wire u2_u2__abc_47660_n155;
  wire u2_u2__abc_47660_n156;
  wire u2_u2__abc_47660_n158;
  wire u2_u2__abc_47660_n159;
  wire u2_u2__abc_47660_n160;
  wire u2_u2__abc_47660_n161;
  wire u2_u2__abc_47660_n163;
  wire u2_u2__abc_47660_n164;
  wire u2_u2__abc_47660_n165;
  wire u2_u2__abc_47660_n166;
  wire u2_u2__abc_47660_n168;
  wire u2_u2__abc_47660_n169;
  wire u2_u2__abc_47660_n170;
  wire u2_u2__abc_47660_n171;
  wire u2_u2__abc_47660_n173;
  wire u2_u2__abc_47660_n174;
  wire u2_u2__abc_47660_n175;
  wire u2_u2__abc_47660_n176;
  wire u2_u2__abc_47660_n178;
  wire u2_u2__abc_47660_n179;
  wire u2_u2__abc_47660_n180;
  wire u2_u2__abc_47660_n181;
  wire u2_u2__abc_47660_n183;
  wire u2_u2__abc_47660_n184;
  wire u2_u2__abc_47660_n185;
  wire u2_u2__abc_47660_n186;
  wire u2_u2__abc_47660_n188;
  wire u2_u2__abc_47660_n189;
  wire u2_u2__abc_47660_n190;
  wire u2_u2__abc_47660_n191;
  wire u2_u2__abc_47660_n193;
  wire u2_u2__abc_47660_n194;
  wire u2_u2__abc_47660_n195;
  wire u2_u2__abc_47660_n196;
  wire u2_u2__abc_47660_n198;
  wire u2_u2__abc_47660_n199;
  wire u2_u2__abc_47660_n200;
  wire u2_u2__abc_47660_n201;
  wire u2_u2__abc_47660_n203;
  wire u2_u2__abc_47660_n204;
  wire u2_u2__abc_47660_n205;
  wire u2_u2__abc_47660_n206;
  wire u2_u2__abc_47660_n207;
  wire u2_u2__abc_47660_n208;
  wire u2_u2__abc_47660_n210;
  wire u2_u2__abc_47660_n211;
  wire u2_u2__abc_47660_n213;
  wire u2_u2__abc_47660_n214;
  wire u2_u2__abc_47660_n216;
  wire u2_u2__abc_47660_n217;
  wire u2_u2__abc_47660_n219;
  wire u2_u2__abc_47660_n220;
  wire u2_u2__abc_47660_n222;
  wire u2_u2__abc_47660_n223;
  wire u2_u2__abc_47660_n225;
  wire u2_u2__abc_47660_n226;
  wire u2_u2__abc_47660_n228;
  wire u2_u2__abc_47660_n229;
  wire u2_u2__abc_47660_n231;
  wire u2_u2__abc_47660_n232;
  wire u2_u2__abc_47660_n234;
  wire u2_u2__abc_47660_n235;
  wire u2_u2__abc_47660_n237;
  wire u2_u2__abc_47660_n238;
  wire u2_u2__abc_47660_n240;
  wire u2_u2__abc_47660_n241;
  wire u2_u2__abc_47660_n243;
  wire u2_u2__abc_47660_n244;
  wire u2_u2__abc_47660_n246;
  wire u2_u2__abc_47660_n247;
  wire u2_u2__abc_47660_n248;
  wire u2_u2__abc_47660_n249;
  wire u2_u2__abc_47660_n250;
  wire u2_u2__abc_47660_n251;
  wire u2_u2__abc_47660_n253;
  wire u2_u2__abc_47660_n254;
  wire u2_u2__abc_47660_n256;
  wire u2_u2__abc_47660_n257;
  wire u2_u2__abc_47660_n259;
  wire u2_u2__abc_47660_n260;
  wire u2_u2__abc_47660_n262;
  wire u2_u2__abc_47660_n263;
  wire u2_u2__abc_47660_n265;
  wire u2_u2__abc_47660_n266;
  wire u2_u2__abc_47660_n268;
  wire u2_u2__abc_47660_n269;
  wire u2_u2__abc_47660_n271;
  wire u2_u2__abc_47660_n272;
  wire u2_u2__abc_47660_n274;
  wire u2_u2__abc_47660_n275_1;
  wire u2_u2__abc_47660_n277;
  wire u2_u2__abc_47660_n278_1;
  wire u2_u2__abc_47660_n280;
  wire u2_u2__abc_47660_n281;
  wire u2_u2__abc_47660_n283_1;
  wire u2_u2__abc_47660_n284;
  wire u2_u2__abc_47660_n286_1;
  wire u2_u2__abc_47660_n287_1;
  wire u2_u2__abc_47660_n289;
  wire u2_u2__abc_47660_n290_1;
  wire u2_u2__abc_47660_n291;
  wire u2_u2__abc_47660_n292_1;
  wire u2_u2__abc_47660_n293;
  wire u2_u2__abc_47660_n295;
  wire u2_u2__abc_47660_n296_1;
  wire u2_u2__abc_47660_n298;
  wire u2_u2__abc_47660_n299;
  wire u2_u2__abc_47660_n301;
  wire u2_u2__abc_47660_n302;
  wire u2_u2__abc_47660_n304_1;
  wire u2_u2__abc_47660_n305;
  wire u2_u2__abc_47660_n305_1;
  wire u2_u2__abc_47660_n307;
  wire u2_u2__abc_47660_n308;
  wire u2_u2__abc_47660_n310;
  wire u2_u2__abc_47660_n311;
  wire u2_u2__abc_47660_n313;
  wire u2_u2__abc_47660_n314;
  wire u2_u2__abc_47660_n316;
  wire u2_u2__abc_47660_n317;
  wire u2_u2__abc_47660_n319;
  wire u2_u2__abc_47660_n320;
  wire u2_u2__abc_47660_n322;
  wire u2_u2__abc_47660_n323;
  wire u2_u2__abc_47660_n325;
  wire u2_u2__abc_47660_n326;
  wire u2_u2__abc_47660_n328;
  wire u2_u2__abc_47660_n329;
  wire u2_u2__abc_47660_n331;
  wire u2_u2__abc_47660_n332;
  wire u2_u2__abc_47660_n333;
  wire u2_u2__abc_47660_n334;
  wire u2_u2__abc_47660_n335;
  wire u2_u2__abc_47660_n336;
  wire u2_u2__abc_47660_n337;
  wire u2_u2__abc_47660_n338;
  wire u2_u2__abc_47660_n339;
  wire u2_u2__abc_47660_n340;
  wire u2_u2__abc_47660_n341;
  wire u2_u2__abc_47660_n342;
  wire u2_u2__abc_47660_n343;
  wire u2_u2__abc_47660_n344;
  wire u2_u2__abc_47660_n345;
  wire u2_u2__abc_47660_n346;
  wire u2_u2__abc_47660_n347;
  wire u2_u2__abc_47660_n348;
  wire u2_u2__abc_47660_n349;
  wire u2_u2__abc_47660_n350;
  wire u2_u2__abc_47660_n351;
  wire u2_u2__abc_47660_n352;
  wire u2_u2__abc_47660_n353;
  wire u2_u2__abc_47660_n354;
  wire u2_u2__abc_47660_n355;
  wire u2_u2__abc_47660_n356;
  wire u2_u2__abc_47660_n357;
  wire u2_u2__abc_47660_n358;
  wire u2_u2__abc_47660_n359;
  wire u2_u2__abc_47660_n360;
  wire u2_u2__abc_47660_n361;
  wire u2_u2__abc_47660_n362;
  wire u2_u2__abc_47660_n363;
  wire u2_u2__abc_47660_n364;
  wire u2_u2__abc_47660_n365;
  wire u2_u2__abc_47660_n366;
  wire u2_u2__abc_47660_n367;
  wire u2_u2__abc_47660_n368;
  wire u2_u2__abc_47660_n369;
  wire u2_u2__abc_47660_n370;
  wire u2_u2__abc_47660_n371;
  wire u2_u2__abc_47660_n372;
  wire u2_u2__abc_47660_n373;
  wire u2_u2__abc_47660_n374;
  wire u2_u2__abc_47660_n375;
  wire u2_u2__abc_47660_n376;
  wire u2_u2__abc_47660_n377;
  wire u2_u2__abc_47660_n378;
  wire u2_u2__abc_47660_n379;
  wire u2_u2__abc_47660_n380;
  wire u2_u2__abc_47660_n381;
  wire u2_u2__abc_47660_n382;
  wire u2_u2__abc_47660_n383;
  wire u2_u2__abc_47660_n384;
  wire u2_u2__abc_47660_n385;
  wire u2_u2__abc_47660_n386;
  wire u2_u2__abc_47660_n387;
  wire u2_u2__abc_47660_n388;
  wire u2_u2__abc_47660_n389;
  wire u2_u2__abc_47660_n390;
  wire u2_u2__abc_47660_n391;
  wire u2_u2__abc_47660_n392;
  wire u2_u2__abc_47660_n393;
  wire u2_u2__abc_47660_n394;
  wire u2_u2__abc_47660_n395;
  wire u2_u2__abc_47660_n396;
  wire u2_u2__abc_47660_n397;
  wire u2_u2__abc_47660_n398;
  wire u2_u2__abc_47660_n399;
  wire u2_u2__abc_47660_n400;
  wire u2_u2__abc_47660_n401;
  wire u2_u2__abc_47660_n402;
  wire u2_u2__abc_47660_n403;
  wire u2_u2__abc_47660_n404;
  wire u2_u2__abc_47660_n405;
  wire u2_u2__abc_47660_n406;
  wire u2_u2__abc_47660_n407;
  wire u2_u2__abc_47660_n408;
  wire u2_u2__abc_47660_n409;
  wire u2_u2__abc_47660_n410;
  wire u2_u2__abc_47660_n411;
  wire u2_u2__abc_47660_n412;
  wire u2_u2__abc_47660_n413;
  wire u2_u2__abc_47660_n414;
  wire u2_u2__abc_47660_n415;
  wire u2_u2__abc_47660_n416;
  wire u2_u2__abc_47660_n417;
  wire u2_u2__abc_47660_n418;
  wire u2_u2__abc_47660_n419;
  wire u2_u2__abc_47660_n420;
  wire u2_u2__abc_47660_n421;
  wire u2_u2__abc_47660_n422;
  wire u2_u2__abc_47660_n423;
  wire u2_u2__abc_47660_n424;
  wire u2_u2__abc_47660_n425;
  wire u2_u2__abc_47660_n426;
  wire u2_u2__abc_47660_n427;
  wire u2_u2__abc_47660_n428;
  wire u2_u2__abc_47660_n429;
  wire u2_u2__abc_47660_n430;
  wire u2_u2__abc_47660_n431;
  wire u2_u2__abc_47660_n432;
  wire u2_u2__abc_47660_n433;
  wire u2_u2__abc_47660_n434;
  wire u2_u2__abc_47660_n435;
  wire u2_u2__abc_47660_n436;
  wire u2_u2__abc_47660_n437;
  wire u2_u2__abc_47660_n438;
  wire u2_u2__abc_47660_n439;
  wire u2_u2__abc_47660_n440;
  wire u2_u2__abc_47660_n441;
  wire u2_u2__abc_47660_n442;
  wire u2_u2__abc_47660_n443;
  wire u2_u2__abc_47660_n444;
  wire u2_u2__abc_47660_n445;
  wire u2_u2__abc_47660_n446;
  wire u2_u2__abc_47660_n447;
  wire u2_u2__abc_47660_n448;
  wire u2_u2__abc_47660_n449;
  wire u2_u2__abc_47660_n450;
  wire u2_u2__abc_47660_n451;
  wire u2_u2__abc_47660_n452;
  wire u2_u2__abc_47660_n453;
  wire u2_u2__abc_47660_n454;
  wire u2_u2__abc_47660_n455;
  wire u2_u2__abc_47660_n456;
  wire u2_u2__abc_47660_n457;
  wire u2_u2__abc_47660_n458;
  wire u2_u2__abc_47660_n459;
  wire u2_u2__abc_47660_n460;
  wire u2_u2__abc_47660_n461;
  wire u2_u2__abc_47660_n462;
  wire u2_u2__abc_47660_n463;
  wire u2_u2__abc_47660_n464;
  wire u2_u2__abc_47660_n465;
  wire u2_u2__abc_47660_n466;
  wire u2_u2__abc_47660_n467;
  wire u2_u2__abc_47660_n468;
  wire u2_u2__abc_47660_n469;
  wire u2_u2__abc_47660_n470;
  wire u2_u2__abc_47660_n471;
  wire u2_u2__abc_47660_n472;
  wire u2_u2__abc_47660_n473;
  wire u2_u2__abc_47660_n474;
  wire u2_u2__abc_47660_n475;
  wire u2_u2__abc_47660_n476;
  wire u2_u2__abc_47660_n477;
  wire u2_u2__abc_47660_n478;
  wire u2_u2__abc_47660_n479;
  wire u2_u2__abc_47660_n480;
  wire u2_u2__abc_47660_n481;
  wire u2_u2__abc_47660_n482;
  wire u2_u2__abc_47660_n483;
  wire u2_u2__abc_47660_n484;
  wire u2_u2__abc_47660_n485;
  wire u2_u2__abc_47660_n486;
  wire u2_u2__abc_47660_n487;
  wire u2_u2__abc_47660_n488;
  wire u2_u2__abc_47660_n489;
  wire u2_u2__abc_47660_n490;
  wire u2_u2__abc_47660_n491;
  wire u2_u2__abc_47660_n492;
  wire u2_u2__abc_47660_n493;
  wire u2_u2__abc_47660_n494;
  wire u2_u2__abc_47660_n495;
  wire u2_u2__abc_47660_n496;
  wire u2_u2__abc_47660_n497;
  wire u2_u2__abc_47660_n498;
  wire u2_u2__abc_47660_n499;
  wire u2_u2__abc_47660_n500;
  wire u2_u2__abc_47660_n501;
  wire u2_u2__abc_47660_n502;
  wire u2_u2__abc_47660_n503;
  wire u2_u2__abc_47660_n504;
  wire u2_u2__abc_47660_n505;
  wire u2_u2__abc_47660_n506;
  wire u2_u2__abc_47660_n507;
  wire u2_u2__abc_47660_n508;
  wire u2_u2__abc_47660_n509;
  wire u2_u2__abc_47660_n510;
  wire u2_u2__abc_47660_n511;
  wire u2_u2__abc_47660_n512;
  wire u2_u2__abc_47660_n513;
  wire u2_u2__abc_47660_n514;
  wire u2_u2__abc_47660_n515;
  wire u2_u2__abc_47660_n516;
  wire u2_u2__abc_47660_n517;
  wire u2_u2__abc_47660_n518;
  wire u2_u2__abc_47660_n519;
  wire u2_u2__abc_47660_n520;
  wire u2_u2__abc_47660_n521;
  wire u2_u2__abc_47660_n522;
  wire u2_u2__abc_47660_n523;
  wire u2_u2__abc_47660_n524;
  wire u2_u2__abc_47660_n525;
  wire u2_u2__abc_47660_n526;
  wire u2_u2__abc_47660_n527;
  wire u2_u2__abc_47660_n528;
  wire u2_u2__abc_47660_n529;
  wire u2_u2__abc_47660_n530;
  wire u2_u2__abc_47660_n531;
  wire u2_u2__abc_47660_n532;
  wire u2_u2__abc_47660_n533;
  wire u2_u2__abc_47660_n534;
  wire u2_u2__abc_47660_n535;
  wire u2_u2__abc_47660_n536;
  wire u2_u2__abc_47660_n537;
  wire u2_u2__abc_47660_n538;
  wire u2_u2__abc_47660_n539;
  wire u2_u2__abc_47660_n540;
  wire u2_u2__abc_47660_n541;
  wire u2_u2__abc_47660_n542;
  wire u2_u2__abc_47660_n543;
  wire u2_u2__abc_47660_n544;
  wire u2_u2__abc_47660_n545;
  wire u2_u2__abc_47660_n546;
  wire u2_u2__abc_47660_n547;
  wire u2_u2__abc_47660_n548;
  wire u2_u2__abc_47660_n549;
  wire u2_u2__abc_47660_n550;
  wire u2_u2__abc_47660_n551;
  wire u2_u2__abc_47660_n552;
  wire u2_u2__abc_47660_n553;
  wire u2_u2__abc_47660_n554;
  wire u2_u2__abc_47660_n555;
  wire u2_u2__abc_47660_n556;
  wire u2_u2__abc_47660_n557;
  wire u2_u2__abc_47660_n558;
  wire u2_u2__abc_47660_n559;
  wire u2_u2__abc_47660_n560;
  wire u2_u2__abc_47660_n561;
  wire u2_u2__abc_47660_n562;
  wire u2_u2__abc_47660_n563;
  wire u2_u2__abc_47660_n564;
  wire u2_u2__abc_47660_n565;
  wire u2_u2__abc_47660_n566;
  wire u2_u2__abc_47660_n567;
  wire u2_u2__abc_47660_n568;
  wire u2_u2__abc_47660_n569;
  wire u2_u2__abc_47660_n570;
  wire u2_u2__abc_47660_n571;
  wire u2_u2__abc_47660_n572;
  wire u2_u2__abc_47660_n573;
  wire u2_u2__abc_47660_n574;
  wire u2_u2__abc_47660_n575;
  wire u2_u2__abc_47660_n576;
  wire u2_u2__abc_47660_n577;
  wire u2_u2__abc_47660_n578;
  wire u2_u2__abc_47660_n579;
  wire u2_u2__abc_47660_n580;
  wire u2_u2__abc_47660_n581;
  wire u2_u2__abc_47660_n582;
  wire u2_u2__abc_47660_n583;
  wire u2_u2__abc_47660_n584;
  wire u2_u2__abc_47660_n585;
  wire u2_u2__abc_47660_n586;
  wire u2_u2__abc_47660_n587;
  wire u2_u2__abc_47660_n588;
  wire u2_u2__abc_47660_n589;
  wire u2_u2__abc_47660_n590;
  wire u2_u2__abc_47660_n591;
  wire u2_u2__abc_47660_n592;
  wire u2_u2__abc_47660_n594;
  wire u2_u2__abc_47660_n595;
  wire u2_u2__abc_47660_n596;
  wire u2_u2__abc_47660_n597;
  wire u2_u2__abc_47660_n598;
  wire u2_u2__abc_47660_n599;
  wire u2_u2__abc_47660_n604;
  wire u2_u2__abc_47660_n605;
  wire u2_u2__abc_47660_n606;
  wire u2_u2__abc_47660_n607;
  wire u2_u2__abc_47660_n608;
  wire u2_u2__abc_47660_n610;
  wire u2_u2__abc_47660_n611;
  wire u2_u2__abc_47660_n612;
  wire u2_u2__abc_47660_n613;
  wire u2_u2__abc_47660_n614;
  wire u2_u2__abc_47660_n616;
  wire u2_u2__abc_47660_n617;
  wire u2_u2__abc_47660_n618;
  wire u2_u2__abc_47660_n619;
  wire u2_u2__abc_47660_n621;
  wire u2_u2__abc_47660_n622;
  wire u2_u2__abc_47660_n623;
  wire u2_u2__abc_47660_n624;
  wire u2_u2_b0_last_row_0_;
  wire u2_u2_b0_last_row_0__FF_INPUT;
  wire u2_u2_b0_last_row_10_;
  wire u2_u2_b0_last_row_10__FF_INPUT;
  wire u2_u2_b0_last_row_11_;
  wire u2_u2_b0_last_row_11__FF_INPUT;
  wire u2_u2_b0_last_row_12_;
  wire u2_u2_b0_last_row_12__FF_INPUT;
  wire u2_u2_b0_last_row_1_;
  wire u2_u2_b0_last_row_1__FF_INPUT;
  wire u2_u2_b0_last_row_2_;
  wire u2_u2_b0_last_row_2__FF_INPUT;
  wire u2_u2_b0_last_row_3_;
  wire u2_u2_b0_last_row_3__FF_INPUT;
  wire u2_u2_b0_last_row_4_;
  wire u2_u2_b0_last_row_4__FF_INPUT;
  wire u2_u2_b0_last_row_5_;
  wire u2_u2_b0_last_row_5__FF_INPUT;
  wire u2_u2_b0_last_row_6_;
  wire u2_u2_b0_last_row_6__FF_INPUT;
  wire u2_u2_b0_last_row_7_;
  wire u2_u2_b0_last_row_7__FF_INPUT;
  wire u2_u2_b0_last_row_8_;
  wire u2_u2_b0_last_row_8__FF_INPUT;
  wire u2_u2_b0_last_row_9_;
  wire u2_u2_b0_last_row_9__FF_INPUT;
  wire u2_u2_b1_last_row_0_;
  wire u2_u2_b1_last_row_0__FF_INPUT;
  wire u2_u2_b1_last_row_10_;
  wire u2_u2_b1_last_row_10__FF_INPUT;
  wire u2_u2_b1_last_row_11_;
  wire u2_u2_b1_last_row_11__FF_INPUT;
  wire u2_u2_b1_last_row_12_;
  wire u2_u2_b1_last_row_12__FF_INPUT;
  wire u2_u2_b1_last_row_1_;
  wire u2_u2_b1_last_row_1__FF_INPUT;
  wire u2_u2_b1_last_row_2_;
  wire u2_u2_b1_last_row_2__FF_INPUT;
  wire u2_u2_b1_last_row_3_;
  wire u2_u2_b1_last_row_3__FF_INPUT;
  wire u2_u2_b1_last_row_4_;
  wire u2_u2_b1_last_row_4__FF_INPUT;
  wire u2_u2_b1_last_row_5_;
  wire u2_u2_b1_last_row_5__FF_INPUT;
  wire u2_u2_b1_last_row_6_;
  wire u2_u2_b1_last_row_6__FF_INPUT;
  wire u2_u2_b1_last_row_7_;
  wire u2_u2_b1_last_row_7__FF_INPUT;
  wire u2_u2_b1_last_row_8_;
  wire u2_u2_b1_last_row_8__FF_INPUT;
  wire u2_u2_b1_last_row_9_;
  wire u2_u2_b1_last_row_9__FF_INPUT;
  wire u2_u2_b2_last_row_0_;
  wire u2_u2_b2_last_row_0__FF_INPUT;
  wire u2_u2_b2_last_row_10_;
  wire u2_u2_b2_last_row_10__FF_INPUT;
  wire u2_u2_b2_last_row_11_;
  wire u2_u2_b2_last_row_11__FF_INPUT;
  wire u2_u2_b2_last_row_12_;
  wire u2_u2_b2_last_row_12__FF_INPUT;
  wire u2_u2_b2_last_row_1_;
  wire u2_u2_b2_last_row_1__FF_INPUT;
  wire u2_u2_b2_last_row_2_;
  wire u2_u2_b2_last_row_2__FF_INPUT;
  wire u2_u2_b2_last_row_3_;
  wire u2_u2_b2_last_row_3__FF_INPUT;
  wire u2_u2_b2_last_row_4_;
  wire u2_u2_b2_last_row_4__FF_INPUT;
  wire u2_u2_b2_last_row_5_;
  wire u2_u2_b2_last_row_5__FF_INPUT;
  wire u2_u2_b2_last_row_6_;
  wire u2_u2_b2_last_row_6__FF_INPUT;
  wire u2_u2_b2_last_row_7_;
  wire u2_u2_b2_last_row_7__FF_INPUT;
  wire u2_u2_b2_last_row_8_;
  wire u2_u2_b2_last_row_8__FF_INPUT;
  wire u2_u2_b2_last_row_9_;
  wire u2_u2_b2_last_row_9__FF_INPUT;
  wire u2_u2_b3_last_row_0_;
  wire u2_u2_b3_last_row_0__FF_INPUT;
  wire u2_u2_b3_last_row_10_;
  wire u2_u2_b3_last_row_10__FF_INPUT;
  wire u2_u2_b3_last_row_11_;
  wire u2_u2_b3_last_row_11__FF_INPUT;
  wire u2_u2_b3_last_row_12_;
  wire u2_u2_b3_last_row_12__FF_INPUT;
  wire u2_u2_b3_last_row_1_;
  wire u2_u2_b3_last_row_1__FF_INPUT;
  wire u2_u2_b3_last_row_2_;
  wire u2_u2_b3_last_row_2__FF_INPUT;
  wire u2_u2_b3_last_row_3_;
  wire u2_u2_b3_last_row_3__FF_INPUT;
  wire u2_u2_b3_last_row_4_;
  wire u2_u2_b3_last_row_4__FF_INPUT;
  wire u2_u2_b3_last_row_5_;
  wire u2_u2_b3_last_row_5__FF_INPUT;
  wire u2_u2_b3_last_row_6_;
  wire u2_u2_b3_last_row_6__FF_INPUT;
  wire u2_u2_b3_last_row_7_;
  wire u2_u2_b3_last_row_7__FF_INPUT;
  wire u2_u2_b3_last_row_8_;
  wire u2_u2_b3_last_row_8__FF_INPUT;
  wire u2_u2_b3_last_row_9_;
  wire u2_u2_b3_last_row_9__FF_INPUT;
  wire u2_u2_bank0_open;
  wire u2_u2_bank0_open_FF_INPUT;
  wire u2_u2_bank1_open;
  wire u2_u2_bank1_open_FF_INPUT;
  wire u2_u2_bank2_open;
  wire u2_u2_bank2_open_FF_INPUT;
  wire u2_u2_bank3_open;
  wire u2_u2_bank3_open_FF_INPUT;
  wire u2_u3__abc_47660_n136;
  wire u2_u3__abc_47660_n137;
  wire u2_u3__abc_47660_n137_bF_buf0;
  wire u2_u3__abc_47660_n137_bF_buf1;
  wire u2_u3__abc_47660_n137_bF_buf2;
  wire u2_u3__abc_47660_n137_bF_buf3;
  wire u2_u3__abc_47660_n137_bF_buf4;
  wire u2_u3__abc_47660_n138;
  wire u2_u3__abc_47660_n139;
  wire u2_u3__abc_47660_n140;
  wire u2_u3__abc_47660_n141;
  wire u2_u3__abc_47660_n143;
  wire u2_u3__abc_47660_n144;
  wire u2_u3__abc_47660_n145;
  wire u2_u3__abc_47660_n146;
  wire u2_u3__abc_47660_n148;
  wire u2_u3__abc_47660_n149;
  wire u2_u3__abc_47660_n150;
  wire u2_u3__abc_47660_n151;
  wire u2_u3__abc_47660_n153;
  wire u2_u3__abc_47660_n154;
  wire u2_u3__abc_47660_n155;
  wire u2_u3__abc_47660_n156;
  wire u2_u3__abc_47660_n158;
  wire u2_u3__abc_47660_n159;
  wire u2_u3__abc_47660_n160;
  wire u2_u3__abc_47660_n161;
  wire u2_u3__abc_47660_n163;
  wire u2_u3__abc_47660_n164;
  wire u2_u3__abc_47660_n165;
  wire u2_u3__abc_47660_n166;
  wire u2_u3__abc_47660_n168;
  wire u2_u3__abc_47660_n169;
  wire u2_u3__abc_47660_n170;
  wire u2_u3__abc_47660_n171;
  wire u2_u3__abc_47660_n173;
  wire u2_u3__abc_47660_n174;
  wire u2_u3__abc_47660_n175;
  wire u2_u3__abc_47660_n176;
  wire u2_u3__abc_47660_n178;
  wire u2_u3__abc_47660_n179;
  wire u2_u3__abc_47660_n180;
  wire u2_u3__abc_47660_n181;
  wire u2_u3__abc_47660_n183;
  wire u2_u3__abc_47660_n184;
  wire u2_u3__abc_47660_n185;
  wire u2_u3__abc_47660_n186;
  wire u2_u3__abc_47660_n188;
  wire u2_u3__abc_47660_n189;
  wire u2_u3__abc_47660_n190;
  wire u2_u3__abc_47660_n191;
  wire u2_u3__abc_47660_n193;
  wire u2_u3__abc_47660_n194;
  wire u2_u3__abc_47660_n195;
  wire u2_u3__abc_47660_n196;
  wire u2_u3__abc_47660_n198;
  wire u2_u3__abc_47660_n199;
  wire u2_u3__abc_47660_n200;
  wire u2_u3__abc_47660_n201;
  wire u2_u3__abc_47660_n203;
  wire u2_u3__abc_47660_n204;
  wire u2_u3__abc_47660_n205;
  wire u2_u3__abc_47660_n206;
  wire u2_u3__abc_47660_n207;
  wire u2_u3__abc_47660_n208;
  wire u2_u3__abc_47660_n210;
  wire u2_u3__abc_47660_n211;
  wire u2_u3__abc_47660_n213;
  wire u2_u3__abc_47660_n214;
  wire u2_u3__abc_47660_n216;
  wire u2_u3__abc_47660_n217;
  wire u2_u3__abc_47660_n219;
  wire u2_u3__abc_47660_n220;
  wire u2_u3__abc_47660_n222;
  wire u2_u3__abc_47660_n223;
  wire u2_u3__abc_47660_n225;
  wire u2_u3__abc_47660_n226;
  wire u2_u3__abc_47660_n228;
  wire u2_u3__abc_47660_n229;
  wire u2_u3__abc_47660_n231;
  wire u2_u3__abc_47660_n232;
  wire u2_u3__abc_47660_n234;
  wire u2_u3__abc_47660_n235;
  wire u2_u3__abc_47660_n237;
  wire u2_u3__abc_47660_n238;
  wire u2_u3__abc_47660_n240;
  wire u2_u3__abc_47660_n241;
  wire u2_u3__abc_47660_n243;
  wire u2_u3__abc_47660_n244;
  wire u2_u3__abc_47660_n246;
  wire u2_u3__abc_47660_n247;
  wire u2_u3__abc_47660_n248;
  wire u2_u3__abc_47660_n249;
  wire u2_u3__abc_47660_n250;
  wire u2_u3__abc_47660_n251;
  wire u2_u3__abc_47660_n253;
  wire u2_u3__abc_47660_n254;
  wire u2_u3__abc_47660_n256;
  wire u2_u3__abc_47660_n257;
  wire u2_u3__abc_47660_n259;
  wire u2_u3__abc_47660_n260;
  wire u2_u3__abc_47660_n262;
  wire u2_u3__abc_47660_n263;
  wire u2_u3__abc_47660_n265;
  wire u2_u3__abc_47660_n266;
  wire u2_u3__abc_47660_n268;
  wire u2_u3__abc_47660_n269;
  wire u2_u3__abc_47660_n271;
  wire u2_u3__abc_47660_n272;
  wire u2_u3__abc_47660_n274;
  wire u2_u3__abc_47660_n275_1;
  wire u2_u3__abc_47660_n277;
  wire u2_u3__abc_47660_n278_1;
  wire u2_u3__abc_47660_n280;
  wire u2_u3__abc_47660_n281;
  wire u2_u3__abc_47660_n283_1;
  wire u2_u3__abc_47660_n284;
  wire u2_u3__abc_47660_n286_1;
  wire u2_u3__abc_47660_n287_1;
  wire u2_u3__abc_47660_n289;
  wire u2_u3__abc_47660_n290_1;
  wire u2_u3__abc_47660_n291;
  wire u2_u3__abc_47660_n292_1;
  wire u2_u3__abc_47660_n293;
  wire u2_u3__abc_47660_n295;
  wire u2_u3__abc_47660_n296_1;
  wire u2_u3__abc_47660_n298;
  wire u2_u3__abc_47660_n299;
  wire u2_u3__abc_47660_n301;
  wire u2_u3__abc_47660_n302;
  wire u2_u3__abc_47660_n304_1;
  wire u2_u3__abc_47660_n305;
  wire u2_u3__abc_47660_n305_1;
  wire u2_u3__abc_47660_n307;
  wire u2_u3__abc_47660_n308;
  wire u2_u3__abc_47660_n310;
  wire u2_u3__abc_47660_n311;
  wire u2_u3__abc_47660_n313;
  wire u2_u3__abc_47660_n314;
  wire u2_u3__abc_47660_n316;
  wire u2_u3__abc_47660_n317;
  wire u2_u3__abc_47660_n319;
  wire u2_u3__abc_47660_n320;
  wire u2_u3__abc_47660_n322;
  wire u2_u3__abc_47660_n323;
  wire u2_u3__abc_47660_n325;
  wire u2_u3__abc_47660_n326;
  wire u2_u3__abc_47660_n328;
  wire u2_u3__abc_47660_n329;
  wire u2_u3__abc_47660_n331;
  wire u2_u3__abc_47660_n332;
  wire u2_u3__abc_47660_n333;
  wire u2_u3__abc_47660_n334;
  wire u2_u3__abc_47660_n335;
  wire u2_u3__abc_47660_n336;
  wire u2_u3__abc_47660_n337;
  wire u2_u3__abc_47660_n338;
  wire u2_u3__abc_47660_n339;
  wire u2_u3__abc_47660_n340;
  wire u2_u3__abc_47660_n341;
  wire u2_u3__abc_47660_n342;
  wire u2_u3__abc_47660_n343;
  wire u2_u3__abc_47660_n344;
  wire u2_u3__abc_47660_n345;
  wire u2_u3__abc_47660_n346;
  wire u2_u3__abc_47660_n347;
  wire u2_u3__abc_47660_n348;
  wire u2_u3__abc_47660_n349;
  wire u2_u3__abc_47660_n350;
  wire u2_u3__abc_47660_n351;
  wire u2_u3__abc_47660_n352;
  wire u2_u3__abc_47660_n353;
  wire u2_u3__abc_47660_n354;
  wire u2_u3__abc_47660_n355;
  wire u2_u3__abc_47660_n356;
  wire u2_u3__abc_47660_n357;
  wire u2_u3__abc_47660_n358;
  wire u2_u3__abc_47660_n359;
  wire u2_u3__abc_47660_n360;
  wire u2_u3__abc_47660_n361;
  wire u2_u3__abc_47660_n362;
  wire u2_u3__abc_47660_n363;
  wire u2_u3__abc_47660_n364;
  wire u2_u3__abc_47660_n365;
  wire u2_u3__abc_47660_n366;
  wire u2_u3__abc_47660_n367;
  wire u2_u3__abc_47660_n368;
  wire u2_u3__abc_47660_n369;
  wire u2_u3__abc_47660_n370;
  wire u2_u3__abc_47660_n371;
  wire u2_u3__abc_47660_n372;
  wire u2_u3__abc_47660_n373;
  wire u2_u3__abc_47660_n374;
  wire u2_u3__abc_47660_n375;
  wire u2_u3__abc_47660_n376;
  wire u2_u3__abc_47660_n377;
  wire u2_u3__abc_47660_n378;
  wire u2_u3__abc_47660_n379;
  wire u2_u3__abc_47660_n380;
  wire u2_u3__abc_47660_n381;
  wire u2_u3__abc_47660_n382;
  wire u2_u3__abc_47660_n383;
  wire u2_u3__abc_47660_n384;
  wire u2_u3__abc_47660_n385;
  wire u2_u3__abc_47660_n386;
  wire u2_u3__abc_47660_n387;
  wire u2_u3__abc_47660_n388;
  wire u2_u3__abc_47660_n389;
  wire u2_u3__abc_47660_n390;
  wire u2_u3__abc_47660_n391;
  wire u2_u3__abc_47660_n392;
  wire u2_u3__abc_47660_n393;
  wire u2_u3__abc_47660_n394;
  wire u2_u3__abc_47660_n395;
  wire u2_u3__abc_47660_n396;
  wire u2_u3__abc_47660_n397;
  wire u2_u3__abc_47660_n398;
  wire u2_u3__abc_47660_n399;
  wire u2_u3__abc_47660_n400;
  wire u2_u3__abc_47660_n401;
  wire u2_u3__abc_47660_n402;
  wire u2_u3__abc_47660_n403;
  wire u2_u3__abc_47660_n404;
  wire u2_u3__abc_47660_n405;
  wire u2_u3__abc_47660_n406;
  wire u2_u3__abc_47660_n407;
  wire u2_u3__abc_47660_n408;
  wire u2_u3__abc_47660_n409;
  wire u2_u3__abc_47660_n410;
  wire u2_u3__abc_47660_n411;
  wire u2_u3__abc_47660_n412;
  wire u2_u3__abc_47660_n413;
  wire u2_u3__abc_47660_n414;
  wire u2_u3__abc_47660_n415;
  wire u2_u3__abc_47660_n416;
  wire u2_u3__abc_47660_n417;
  wire u2_u3__abc_47660_n418;
  wire u2_u3__abc_47660_n419;
  wire u2_u3__abc_47660_n420;
  wire u2_u3__abc_47660_n421;
  wire u2_u3__abc_47660_n422;
  wire u2_u3__abc_47660_n423;
  wire u2_u3__abc_47660_n424;
  wire u2_u3__abc_47660_n425;
  wire u2_u3__abc_47660_n426;
  wire u2_u3__abc_47660_n427;
  wire u2_u3__abc_47660_n428;
  wire u2_u3__abc_47660_n429;
  wire u2_u3__abc_47660_n430;
  wire u2_u3__abc_47660_n431;
  wire u2_u3__abc_47660_n432;
  wire u2_u3__abc_47660_n433;
  wire u2_u3__abc_47660_n434;
  wire u2_u3__abc_47660_n435;
  wire u2_u3__abc_47660_n436;
  wire u2_u3__abc_47660_n437;
  wire u2_u3__abc_47660_n438;
  wire u2_u3__abc_47660_n439;
  wire u2_u3__abc_47660_n440;
  wire u2_u3__abc_47660_n441;
  wire u2_u3__abc_47660_n442;
  wire u2_u3__abc_47660_n443;
  wire u2_u3__abc_47660_n444;
  wire u2_u3__abc_47660_n445;
  wire u2_u3__abc_47660_n446;
  wire u2_u3__abc_47660_n447;
  wire u2_u3__abc_47660_n448;
  wire u2_u3__abc_47660_n449;
  wire u2_u3__abc_47660_n450;
  wire u2_u3__abc_47660_n451;
  wire u2_u3__abc_47660_n452;
  wire u2_u3__abc_47660_n453;
  wire u2_u3__abc_47660_n454;
  wire u2_u3__abc_47660_n455;
  wire u2_u3__abc_47660_n456;
  wire u2_u3__abc_47660_n457;
  wire u2_u3__abc_47660_n458;
  wire u2_u3__abc_47660_n459;
  wire u2_u3__abc_47660_n460;
  wire u2_u3__abc_47660_n461;
  wire u2_u3__abc_47660_n462;
  wire u2_u3__abc_47660_n463;
  wire u2_u3__abc_47660_n464;
  wire u2_u3__abc_47660_n465;
  wire u2_u3__abc_47660_n466;
  wire u2_u3__abc_47660_n467;
  wire u2_u3__abc_47660_n468;
  wire u2_u3__abc_47660_n469;
  wire u2_u3__abc_47660_n470;
  wire u2_u3__abc_47660_n471;
  wire u2_u3__abc_47660_n472;
  wire u2_u3__abc_47660_n473;
  wire u2_u3__abc_47660_n474;
  wire u2_u3__abc_47660_n475;
  wire u2_u3__abc_47660_n476;
  wire u2_u3__abc_47660_n477;
  wire u2_u3__abc_47660_n478;
  wire u2_u3__abc_47660_n479;
  wire u2_u3__abc_47660_n480;
  wire u2_u3__abc_47660_n481;
  wire u2_u3__abc_47660_n482;
  wire u2_u3__abc_47660_n483;
  wire u2_u3__abc_47660_n484;
  wire u2_u3__abc_47660_n485;
  wire u2_u3__abc_47660_n486;
  wire u2_u3__abc_47660_n487;
  wire u2_u3__abc_47660_n488;
  wire u2_u3__abc_47660_n489;
  wire u2_u3__abc_47660_n490;
  wire u2_u3__abc_47660_n491;
  wire u2_u3__abc_47660_n492;
  wire u2_u3__abc_47660_n493;
  wire u2_u3__abc_47660_n494;
  wire u2_u3__abc_47660_n495;
  wire u2_u3__abc_47660_n496;
  wire u2_u3__abc_47660_n497;
  wire u2_u3__abc_47660_n498;
  wire u2_u3__abc_47660_n499;
  wire u2_u3__abc_47660_n500;
  wire u2_u3__abc_47660_n501;
  wire u2_u3__abc_47660_n502;
  wire u2_u3__abc_47660_n503;
  wire u2_u3__abc_47660_n504;
  wire u2_u3__abc_47660_n505;
  wire u2_u3__abc_47660_n506;
  wire u2_u3__abc_47660_n507;
  wire u2_u3__abc_47660_n508;
  wire u2_u3__abc_47660_n509;
  wire u2_u3__abc_47660_n510;
  wire u2_u3__abc_47660_n511;
  wire u2_u3__abc_47660_n512;
  wire u2_u3__abc_47660_n513;
  wire u2_u3__abc_47660_n514;
  wire u2_u3__abc_47660_n515;
  wire u2_u3__abc_47660_n516;
  wire u2_u3__abc_47660_n517;
  wire u2_u3__abc_47660_n518;
  wire u2_u3__abc_47660_n519;
  wire u2_u3__abc_47660_n520;
  wire u2_u3__abc_47660_n521;
  wire u2_u3__abc_47660_n522;
  wire u2_u3__abc_47660_n523;
  wire u2_u3__abc_47660_n524;
  wire u2_u3__abc_47660_n525;
  wire u2_u3__abc_47660_n526;
  wire u2_u3__abc_47660_n527;
  wire u2_u3__abc_47660_n528;
  wire u2_u3__abc_47660_n529;
  wire u2_u3__abc_47660_n530;
  wire u2_u3__abc_47660_n531;
  wire u2_u3__abc_47660_n532;
  wire u2_u3__abc_47660_n533;
  wire u2_u3__abc_47660_n534;
  wire u2_u3__abc_47660_n535;
  wire u2_u3__abc_47660_n536;
  wire u2_u3__abc_47660_n537;
  wire u2_u3__abc_47660_n538;
  wire u2_u3__abc_47660_n539;
  wire u2_u3__abc_47660_n540;
  wire u2_u3__abc_47660_n541;
  wire u2_u3__abc_47660_n542;
  wire u2_u3__abc_47660_n543;
  wire u2_u3__abc_47660_n544;
  wire u2_u3__abc_47660_n545;
  wire u2_u3__abc_47660_n546;
  wire u2_u3__abc_47660_n547;
  wire u2_u3__abc_47660_n548;
  wire u2_u3__abc_47660_n549;
  wire u2_u3__abc_47660_n550;
  wire u2_u3__abc_47660_n551;
  wire u2_u3__abc_47660_n552;
  wire u2_u3__abc_47660_n553;
  wire u2_u3__abc_47660_n554;
  wire u2_u3__abc_47660_n555;
  wire u2_u3__abc_47660_n556;
  wire u2_u3__abc_47660_n557;
  wire u2_u3__abc_47660_n558;
  wire u2_u3__abc_47660_n559;
  wire u2_u3__abc_47660_n560;
  wire u2_u3__abc_47660_n561;
  wire u2_u3__abc_47660_n562;
  wire u2_u3__abc_47660_n563;
  wire u2_u3__abc_47660_n564;
  wire u2_u3__abc_47660_n565;
  wire u2_u3__abc_47660_n566;
  wire u2_u3__abc_47660_n567;
  wire u2_u3__abc_47660_n568;
  wire u2_u3__abc_47660_n569;
  wire u2_u3__abc_47660_n570;
  wire u2_u3__abc_47660_n571;
  wire u2_u3__abc_47660_n572;
  wire u2_u3__abc_47660_n573;
  wire u2_u3__abc_47660_n574;
  wire u2_u3__abc_47660_n575;
  wire u2_u3__abc_47660_n576;
  wire u2_u3__abc_47660_n577;
  wire u2_u3__abc_47660_n578;
  wire u2_u3__abc_47660_n579;
  wire u2_u3__abc_47660_n580;
  wire u2_u3__abc_47660_n581;
  wire u2_u3__abc_47660_n582;
  wire u2_u3__abc_47660_n583;
  wire u2_u3__abc_47660_n584;
  wire u2_u3__abc_47660_n585;
  wire u2_u3__abc_47660_n586;
  wire u2_u3__abc_47660_n587;
  wire u2_u3__abc_47660_n588;
  wire u2_u3__abc_47660_n589;
  wire u2_u3__abc_47660_n590;
  wire u2_u3__abc_47660_n591;
  wire u2_u3__abc_47660_n592;
  wire u2_u3__abc_47660_n594;
  wire u2_u3__abc_47660_n595;
  wire u2_u3__abc_47660_n596;
  wire u2_u3__abc_47660_n597;
  wire u2_u3__abc_47660_n598;
  wire u2_u3__abc_47660_n599;
  wire u2_u3__abc_47660_n604;
  wire u2_u3__abc_47660_n605;
  wire u2_u3__abc_47660_n606;
  wire u2_u3__abc_47660_n607;
  wire u2_u3__abc_47660_n608;
  wire u2_u3__abc_47660_n610;
  wire u2_u3__abc_47660_n611;
  wire u2_u3__abc_47660_n612;
  wire u2_u3__abc_47660_n613;
  wire u2_u3__abc_47660_n614;
  wire u2_u3__abc_47660_n616;
  wire u2_u3__abc_47660_n617;
  wire u2_u3__abc_47660_n618;
  wire u2_u3__abc_47660_n619;
  wire u2_u3__abc_47660_n621;
  wire u2_u3__abc_47660_n622;
  wire u2_u3__abc_47660_n623;
  wire u2_u3__abc_47660_n624;
  wire u2_u3_b0_last_row_0_;
  wire u2_u3_b0_last_row_0__FF_INPUT;
  wire u2_u3_b0_last_row_10_;
  wire u2_u3_b0_last_row_10__FF_INPUT;
  wire u2_u3_b0_last_row_11_;
  wire u2_u3_b0_last_row_11__FF_INPUT;
  wire u2_u3_b0_last_row_12_;
  wire u2_u3_b0_last_row_12__FF_INPUT;
  wire u2_u3_b0_last_row_1_;
  wire u2_u3_b0_last_row_1__FF_INPUT;
  wire u2_u3_b0_last_row_2_;
  wire u2_u3_b0_last_row_2__FF_INPUT;
  wire u2_u3_b0_last_row_3_;
  wire u2_u3_b0_last_row_3__FF_INPUT;
  wire u2_u3_b0_last_row_4_;
  wire u2_u3_b0_last_row_4__FF_INPUT;
  wire u2_u3_b0_last_row_5_;
  wire u2_u3_b0_last_row_5__FF_INPUT;
  wire u2_u3_b0_last_row_6_;
  wire u2_u3_b0_last_row_6__FF_INPUT;
  wire u2_u3_b0_last_row_7_;
  wire u2_u3_b0_last_row_7__FF_INPUT;
  wire u2_u3_b0_last_row_8_;
  wire u2_u3_b0_last_row_8__FF_INPUT;
  wire u2_u3_b0_last_row_9_;
  wire u2_u3_b0_last_row_9__FF_INPUT;
  wire u2_u3_b1_last_row_0_;
  wire u2_u3_b1_last_row_0__FF_INPUT;
  wire u2_u3_b1_last_row_10_;
  wire u2_u3_b1_last_row_10__FF_INPUT;
  wire u2_u3_b1_last_row_11_;
  wire u2_u3_b1_last_row_11__FF_INPUT;
  wire u2_u3_b1_last_row_12_;
  wire u2_u3_b1_last_row_12__FF_INPUT;
  wire u2_u3_b1_last_row_1_;
  wire u2_u3_b1_last_row_1__FF_INPUT;
  wire u2_u3_b1_last_row_2_;
  wire u2_u3_b1_last_row_2__FF_INPUT;
  wire u2_u3_b1_last_row_3_;
  wire u2_u3_b1_last_row_3__FF_INPUT;
  wire u2_u3_b1_last_row_4_;
  wire u2_u3_b1_last_row_4__FF_INPUT;
  wire u2_u3_b1_last_row_5_;
  wire u2_u3_b1_last_row_5__FF_INPUT;
  wire u2_u3_b1_last_row_6_;
  wire u2_u3_b1_last_row_6__FF_INPUT;
  wire u2_u3_b1_last_row_7_;
  wire u2_u3_b1_last_row_7__FF_INPUT;
  wire u2_u3_b1_last_row_8_;
  wire u2_u3_b1_last_row_8__FF_INPUT;
  wire u2_u3_b1_last_row_9_;
  wire u2_u3_b1_last_row_9__FF_INPUT;
  wire u2_u3_b2_last_row_0_;
  wire u2_u3_b2_last_row_0__FF_INPUT;
  wire u2_u3_b2_last_row_10_;
  wire u2_u3_b2_last_row_10__FF_INPUT;
  wire u2_u3_b2_last_row_11_;
  wire u2_u3_b2_last_row_11__FF_INPUT;
  wire u2_u3_b2_last_row_12_;
  wire u2_u3_b2_last_row_12__FF_INPUT;
  wire u2_u3_b2_last_row_1_;
  wire u2_u3_b2_last_row_1__FF_INPUT;
  wire u2_u3_b2_last_row_2_;
  wire u2_u3_b2_last_row_2__FF_INPUT;
  wire u2_u3_b2_last_row_3_;
  wire u2_u3_b2_last_row_3__FF_INPUT;
  wire u2_u3_b2_last_row_4_;
  wire u2_u3_b2_last_row_4__FF_INPUT;
  wire u2_u3_b2_last_row_5_;
  wire u2_u3_b2_last_row_5__FF_INPUT;
  wire u2_u3_b2_last_row_6_;
  wire u2_u3_b2_last_row_6__FF_INPUT;
  wire u2_u3_b2_last_row_7_;
  wire u2_u3_b2_last_row_7__FF_INPUT;
  wire u2_u3_b2_last_row_8_;
  wire u2_u3_b2_last_row_8__FF_INPUT;
  wire u2_u3_b2_last_row_9_;
  wire u2_u3_b2_last_row_9__FF_INPUT;
  wire u2_u3_b3_last_row_0_;
  wire u2_u3_b3_last_row_0__FF_INPUT;
  wire u2_u3_b3_last_row_10_;
  wire u2_u3_b3_last_row_10__FF_INPUT;
  wire u2_u3_b3_last_row_11_;
  wire u2_u3_b3_last_row_11__FF_INPUT;
  wire u2_u3_b3_last_row_12_;
  wire u2_u3_b3_last_row_12__FF_INPUT;
  wire u2_u3_b3_last_row_1_;
  wire u2_u3_b3_last_row_1__FF_INPUT;
  wire u2_u3_b3_last_row_2_;
  wire u2_u3_b3_last_row_2__FF_INPUT;
  wire u2_u3_b3_last_row_3_;
  wire u2_u3_b3_last_row_3__FF_INPUT;
  wire u2_u3_b3_last_row_4_;
  wire u2_u3_b3_last_row_4__FF_INPUT;
  wire u2_u3_b3_last_row_5_;
  wire u2_u3_b3_last_row_5__FF_INPUT;
  wire u2_u3_b3_last_row_6_;
  wire u2_u3_b3_last_row_6__FF_INPUT;
  wire u2_u3_b3_last_row_7_;
  wire u2_u3_b3_last_row_7__FF_INPUT;
  wire u2_u3_b3_last_row_8_;
  wire u2_u3_b3_last_row_8__FF_INPUT;
  wire u2_u3_b3_last_row_9_;
  wire u2_u3_b3_last_row_9__FF_INPUT;
  wire u2_u3_bank0_open;
  wire u2_u3_bank0_open_FF_INPUT;
  wire u2_u3_bank1_open;
  wire u2_u3_bank1_open_FF_INPUT;
  wire u2_u3_bank2_open;
  wire u2_u3_bank2_open_FF_INPUT;
  wire u2_u3_bank3_open;
  wire u2_u3_bank3_open_FF_INPUT;
  wire u2_u4__abc_47660_n136;
  wire u2_u4__abc_47660_n137;
  wire u2_u4__abc_47660_n137_bF_buf0;
  wire u2_u4__abc_47660_n137_bF_buf1;
  wire u2_u4__abc_47660_n137_bF_buf2;
  wire u2_u4__abc_47660_n137_bF_buf3;
  wire u2_u4__abc_47660_n137_bF_buf4;
  wire u2_u4__abc_47660_n138;
  wire u2_u4__abc_47660_n139;
  wire u2_u4__abc_47660_n140;
  wire u2_u4__abc_47660_n141;
  wire u2_u4__abc_47660_n143;
  wire u2_u4__abc_47660_n144;
  wire u2_u4__abc_47660_n145;
  wire u2_u4__abc_47660_n146;
  wire u2_u4__abc_47660_n148;
  wire u2_u4__abc_47660_n149;
  wire u2_u4__abc_47660_n150;
  wire u2_u4__abc_47660_n151;
  wire u2_u4__abc_47660_n153;
  wire u2_u4__abc_47660_n154;
  wire u2_u4__abc_47660_n155;
  wire u2_u4__abc_47660_n156;
  wire u2_u4__abc_47660_n158;
  wire u2_u4__abc_47660_n159;
  wire u2_u4__abc_47660_n160;
  wire u2_u4__abc_47660_n161;
  wire u2_u4__abc_47660_n163;
  wire u2_u4__abc_47660_n164;
  wire u2_u4__abc_47660_n165;
  wire u2_u4__abc_47660_n166;
  wire u2_u4__abc_47660_n168;
  wire u2_u4__abc_47660_n169;
  wire u2_u4__abc_47660_n170;
  wire u2_u4__abc_47660_n171;
  wire u2_u4__abc_47660_n173;
  wire u2_u4__abc_47660_n174;
  wire u2_u4__abc_47660_n175;
  wire u2_u4__abc_47660_n176;
  wire u2_u4__abc_47660_n178;
  wire u2_u4__abc_47660_n179;
  wire u2_u4__abc_47660_n180;
  wire u2_u4__abc_47660_n181;
  wire u2_u4__abc_47660_n183;
  wire u2_u4__abc_47660_n184;
  wire u2_u4__abc_47660_n185;
  wire u2_u4__abc_47660_n186;
  wire u2_u4__abc_47660_n188;
  wire u2_u4__abc_47660_n189;
  wire u2_u4__abc_47660_n190;
  wire u2_u4__abc_47660_n191;
  wire u2_u4__abc_47660_n193;
  wire u2_u4__abc_47660_n194;
  wire u2_u4__abc_47660_n195;
  wire u2_u4__abc_47660_n196;
  wire u2_u4__abc_47660_n198;
  wire u2_u4__abc_47660_n199;
  wire u2_u4__abc_47660_n200;
  wire u2_u4__abc_47660_n201;
  wire u2_u4__abc_47660_n203;
  wire u2_u4__abc_47660_n204;
  wire u2_u4__abc_47660_n205;
  wire u2_u4__abc_47660_n206;
  wire u2_u4__abc_47660_n207;
  wire u2_u4__abc_47660_n208;
  wire u2_u4__abc_47660_n210;
  wire u2_u4__abc_47660_n211;
  wire u2_u4__abc_47660_n213;
  wire u2_u4__abc_47660_n214;
  wire u2_u4__abc_47660_n216;
  wire u2_u4__abc_47660_n217;
  wire u2_u4__abc_47660_n219;
  wire u2_u4__abc_47660_n220;
  wire u2_u4__abc_47660_n222;
  wire u2_u4__abc_47660_n223;
  wire u2_u4__abc_47660_n225;
  wire u2_u4__abc_47660_n226;
  wire u2_u4__abc_47660_n228;
  wire u2_u4__abc_47660_n229;
  wire u2_u4__abc_47660_n231;
  wire u2_u4__abc_47660_n232;
  wire u2_u4__abc_47660_n234;
  wire u2_u4__abc_47660_n235;
  wire u2_u4__abc_47660_n237;
  wire u2_u4__abc_47660_n238;
  wire u2_u4__abc_47660_n240;
  wire u2_u4__abc_47660_n241;
  wire u2_u4__abc_47660_n243;
  wire u2_u4__abc_47660_n244;
  wire u2_u4__abc_47660_n246;
  wire u2_u4__abc_47660_n247;
  wire u2_u4__abc_47660_n248;
  wire u2_u4__abc_47660_n249;
  wire u2_u4__abc_47660_n250;
  wire u2_u4__abc_47660_n251;
  wire u2_u4__abc_47660_n253;
  wire u2_u4__abc_47660_n254;
  wire u2_u4__abc_47660_n256;
  wire u2_u4__abc_47660_n257;
  wire u2_u4__abc_47660_n259;
  wire u2_u4__abc_47660_n260;
  wire u2_u4__abc_47660_n262;
  wire u2_u4__abc_47660_n263;
  wire u2_u4__abc_47660_n265;
  wire u2_u4__abc_47660_n266;
  wire u2_u4__abc_47660_n268;
  wire u2_u4__abc_47660_n269;
  wire u2_u4__abc_47660_n271;
  wire u2_u4__abc_47660_n272;
  wire u2_u4__abc_47660_n274;
  wire u2_u4__abc_47660_n275_1;
  wire u2_u4__abc_47660_n277;
  wire u2_u4__abc_47660_n278_1;
  wire u2_u4__abc_47660_n280;
  wire u2_u4__abc_47660_n281;
  wire u2_u4__abc_47660_n283_1;
  wire u2_u4__abc_47660_n284;
  wire u2_u4__abc_47660_n286_1;
  wire u2_u4__abc_47660_n287_1;
  wire u2_u4__abc_47660_n289;
  wire u2_u4__abc_47660_n290_1;
  wire u2_u4__abc_47660_n291;
  wire u2_u4__abc_47660_n292_1;
  wire u2_u4__abc_47660_n293;
  wire u2_u4__abc_47660_n295;
  wire u2_u4__abc_47660_n296_1;
  wire u2_u4__abc_47660_n298;
  wire u2_u4__abc_47660_n299;
  wire u2_u4__abc_47660_n301;
  wire u2_u4__abc_47660_n302;
  wire u2_u4__abc_47660_n304_1;
  wire u2_u4__abc_47660_n305;
  wire u2_u4__abc_47660_n305_1;
  wire u2_u4__abc_47660_n307;
  wire u2_u4__abc_47660_n308;
  wire u2_u4__abc_47660_n310;
  wire u2_u4__abc_47660_n311;
  wire u2_u4__abc_47660_n313;
  wire u2_u4__abc_47660_n314;
  wire u2_u4__abc_47660_n316;
  wire u2_u4__abc_47660_n317;
  wire u2_u4__abc_47660_n319;
  wire u2_u4__abc_47660_n320;
  wire u2_u4__abc_47660_n322;
  wire u2_u4__abc_47660_n323;
  wire u2_u4__abc_47660_n325;
  wire u2_u4__abc_47660_n326;
  wire u2_u4__abc_47660_n328;
  wire u2_u4__abc_47660_n329;
  wire u2_u4__abc_47660_n331;
  wire u2_u4__abc_47660_n332;
  wire u2_u4__abc_47660_n333;
  wire u2_u4__abc_47660_n334;
  wire u2_u4__abc_47660_n335;
  wire u2_u4__abc_47660_n336;
  wire u2_u4__abc_47660_n337;
  wire u2_u4__abc_47660_n338;
  wire u2_u4__abc_47660_n339;
  wire u2_u4__abc_47660_n340;
  wire u2_u4__abc_47660_n341;
  wire u2_u4__abc_47660_n342;
  wire u2_u4__abc_47660_n343;
  wire u2_u4__abc_47660_n344;
  wire u2_u4__abc_47660_n345;
  wire u2_u4__abc_47660_n346;
  wire u2_u4__abc_47660_n347;
  wire u2_u4__abc_47660_n348;
  wire u2_u4__abc_47660_n349;
  wire u2_u4__abc_47660_n350;
  wire u2_u4__abc_47660_n351;
  wire u2_u4__abc_47660_n352;
  wire u2_u4__abc_47660_n353;
  wire u2_u4__abc_47660_n354;
  wire u2_u4__abc_47660_n355;
  wire u2_u4__abc_47660_n356;
  wire u2_u4__abc_47660_n357;
  wire u2_u4__abc_47660_n358;
  wire u2_u4__abc_47660_n359;
  wire u2_u4__abc_47660_n360;
  wire u2_u4__abc_47660_n361;
  wire u2_u4__abc_47660_n362;
  wire u2_u4__abc_47660_n363;
  wire u2_u4__abc_47660_n364;
  wire u2_u4__abc_47660_n365;
  wire u2_u4__abc_47660_n366;
  wire u2_u4__abc_47660_n367;
  wire u2_u4__abc_47660_n368;
  wire u2_u4__abc_47660_n369;
  wire u2_u4__abc_47660_n370;
  wire u2_u4__abc_47660_n371;
  wire u2_u4__abc_47660_n372;
  wire u2_u4__abc_47660_n373;
  wire u2_u4__abc_47660_n374;
  wire u2_u4__abc_47660_n375;
  wire u2_u4__abc_47660_n376;
  wire u2_u4__abc_47660_n377;
  wire u2_u4__abc_47660_n378;
  wire u2_u4__abc_47660_n379;
  wire u2_u4__abc_47660_n380;
  wire u2_u4__abc_47660_n381;
  wire u2_u4__abc_47660_n382;
  wire u2_u4__abc_47660_n383;
  wire u2_u4__abc_47660_n384;
  wire u2_u4__abc_47660_n385;
  wire u2_u4__abc_47660_n386;
  wire u2_u4__abc_47660_n387;
  wire u2_u4__abc_47660_n388;
  wire u2_u4__abc_47660_n389;
  wire u2_u4__abc_47660_n390;
  wire u2_u4__abc_47660_n391;
  wire u2_u4__abc_47660_n392;
  wire u2_u4__abc_47660_n393;
  wire u2_u4__abc_47660_n394;
  wire u2_u4__abc_47660_n395;
  wire u2_u4__abc_47660_n396;
  wire u2_u4__abc_47660_n397;
  wire u2_u4__abc_47660_n398;
  wire u2_u4__abc_47660_n399;
  wire u2_u4__abc_47660_n400;
  wire u2_u4__abc_47660_n401;
  wire u2_u4__abc_47660_n402;
  wire u2_u4__abc_47660_n403;
  wire u2_u4__abc_47660_n404;
  wire u2_u4__abc_47660_n405;
  wire u2_u4__abc_47660_n406;
  wire u2_u4__abc_47660_n407;
  wire u2_u4__abc_47660_n408;
  wire u2_u4__abc_47660_n409;
  wire u2_u4__abc_47660_n410;
  wire u2_u4__abc_47660_n411;
  wire u2_u4__abc_47660_n412;
  wire u2_u4__abc_47660_n413;
  wire u2_u4__abc_47660_n414;
  wire u2_u4__abc_47660_n415;
  wire u2_u4__abc_47660_n416;
  wire u2_u4__abc_47660_n417;
  wire u2_u4__abc_47660_n418;
  wire u2_u4__abc_47660_n419;
  wire u2_u4__abc_47660_n420;
  wire u2_u4__abc_47660_n421;
  wire u2_u4__abc_47660_n422;
  wire u2_u4__abc_47660_n423;
  wire u2_u4__abc_47660_n424;
  wire u2_u4__abc_47660_n425;
  wire u2_u4__abc_47660_n426;
  wire u2_u4__abc_47660_n427;
  wire u2_u4__abc_47660_n428;
  wire u2_u4__abc_47660_n429;
  wire u2_u4__abc_47660_n430;
  wire u2_u4__abc_47660_n431;
  wire u2_u4__abc_47660_n432;
  wire u2_u4__abc_47660_n433;
  wire u2_u4__abc_47660_n434;
  wire u2_u4__abc_47660_n435;
  wire u2_u4__abc_47660_n436;
  wire u2_u4__abc_47660_n437;
  wire u2_u4__abc_47660_n438;
  wire u2_u4__abc_47660_n439;
  wire u2_u4__abc_47660_n440;
  wire u2_u4__abc_47660_n441;
  wire u2_u4__abc_47660_n442;
  wire u2_u4__abc_47660_n443;
  wire u2_u4__abc_47660_n444;
  wire u2_u4__abc_47660_n445;
  wire u2_u4__abc_47660_n446;
  wire u2_u4__abc_47660_n447;
  wire u2_u4__abc_47660_n448;
  wire u2_u4__abc_47660_n449;
  wire u2_u4__abc_47660_n450;
  wire u2_u4__abc_47660_n451;
  wire u2_u4__abc_47660_n452;
  wire u2_u4__abc_47660_n453;
  wire u2_u4__abc_47660_n454;
  wire u2_u4__abc_47660_n455;
  wire u2_u4__abc_47660_n456;
  wire u2_u4__abc_47660_n457;
  wire u2_u4__abc_47660_n458;
  wire u2_u4__abc_47660_n459;
  wire u2_u4__abc_47660_n460;
  wire u2_u4__abc_47660_n461;
  wire u2_u4__abc_47660_n462;
  wire u2_u4__abc_47660_n463;
  wire u2_u4__abc_47660_n464;
  wire u2_u4__abc_47660_n465;
  wire u2_u4__abc_47660_n466;
  wire u2_u4__abc_47660_n467;
  wire u2_u4__abc_47660_n468;
  wire u2_u4__abc_47660_n469;
  wire u2_u4__abc_47660_n470;
  wire u2_u4__abc_47660_n471;
  wire u2_u4__abc_47660_n472;
  wire u2_u4__abc_47660_n473;
  wire u2_u4__abc_47660_n474;
  wire u2_u4__abc_47660_n475;
  wire u2_u4__abc_47660_n476;
  wire u2_u4__abc_47660_n477;
  wire u2_u4__abc_47660_n478;
  wire u2_u4__abc_47660_n479;
  wire u2_u4__abc_47660_n480;
  wire u2_u4__abc_47660_n481;
  wire u2_u4__abc_47660_n482;
  wire u2_u4__abc_47660_n483;
  wire u2_u4__abc_47660_n484;
  wire u2_u4__abc_47660_n485;
  wire u2_u4__abc_47660_n486;
  wire u2_u4__abc_47660_n487;
  wire u2_u4__abc_47660_n488;
  wire u2_u4__abc_47660_n489;
  wire u2_u4__abc_47660_n490;
  wire u2_u4__abc_47660_n491;
  wire u2_u4__abc_47660_n492;
  wire u2_u4__abc_47660_n493;
  wire u2_u4__abc_47660_n494;
  wire u2_u4__abc_47660_n495;
  wire u2_u4__abc_47660_n496;
  wire u2_u4__abc_47660_n497;
  wire u2_u4__abc_47660_n498;
  wire u2_u4__abc_47660_n499;
  wire u2_u4__abc_47660_n500;
  wire u2_u4__abc_47660_n501;
  wire u2_u4__abc_47660_n502;
  wire u2_u4__abc_47660_n503;
  wire u2_u4__abc_47660_n504;
  wire u2_u4__abc_47660_n505;
  wire u2_u4__abc_47660_n506;
  wire u2_u4__abc_47660_n507;
  wire u2_u4__abc_47660_n508;
  wire u2_u4__abc_47660_n509;
  wire u2_u4__abc_47660_n510;
  wire u2_u4__abc_47660_n511;
  wire u2_u4__abc_47660_n512;
  wire u2_u4__abc_47660_n513;
  wire u2_u4__abc_47660_n514;
  wire u2_u4__abc_47660_n515;
  wire u2_u4__abc_47660_n516;
  wire u2_u4__abc_47660_n517;
  wire u2_u4__abc_47660_n518;
  wire u2_u4__abc_47660_n519;
  wire u2_u4__abc_47660_n520;
  wire u2_u4__abc_47660_n521;
  wire u2_u4__abc_47660_n522;
  wire u2_u4__abc_47660_n523;
  wire u2_u4__abc_47660_n524;
  wire u2_u4__abc_47660_n525;
  wire u2_u4__abc_47660_n526;
  wire u2_u4__abc_47660_n527;
  wire u2_u4__abc_47660_n528;
  wire u2_u4__abc_47660_n529;
  wire u2_u4__abc_47660_n530;
  wire u2_u4__abc_47660_n531;
  wire u2_u4__abc_47660_n532;
  wire u2_u4__abc_47660_n533;
  wire u2_u4__abc_47660_n534;
  wire u2_u4__abc_47660_n535;
  wire u2_u4__abc_47660_n536;
  wire u2_u4__abc_47660_n537;
  wire u2_u4__abc_47660_n538;
  wire u2_u4__abc_47660_n539;
  wire u2_u4__abc_47660_n540;
  wire u2_u4__abc_47660_n541;
  wire u2_u4__abc_47660_n542;
  wire u2_u4__abc_47660_n543;
  wire u2_u4__abc_47660_n544;
  wire u2_u4__abc_47660_n545;
  wire u2_u4__abc_47660_n546;
  wire u2_u4__abc_47660_n547;
  wire u2_u4__abc_47660_n548;
  wire u2_u4__abc_47660_n549;
  wire u2_u4__abc_47660_n550;
  wire u2_u4__abc_47660_n551;
  wire u2_u4__abc_47660_n552;
  wire u2_u4__abc_47660_n553;
  wire u2_u4__abc_47660_n554;
  wire u2_u4__abc_47660_n555;
  wire u2_u4__abc_47660_n556;
  wire u2_u4__abc_47660_n557;
  wire u2_u4__abc_47660_n558;
  wire u2_u4__abc_47660_n559;
  wire u2_u4__abc_47660_n560;
  wire u2_u4__abc_47660_n561;
  wire u2_u4__abc_47660_n562;
  wire u2_u4__abc_47660_n563;
  wire u2_u4__abc_47660_n564;
  wire u2_u4__abc_47660_n565;
  wire u2_u4__abc_47660_n566;
  wire u2_u4__abc_47660_n567;
  wire u2_u4__abc_47660_n568;
  wire u2_u4__abc_47660_n569;
  wire u2_u4__abc_47660_n570;
  wire u2_u4__abc_47660_n571;
  wire u2_u4__abc_47660_n572;
  wire u2_u4__abc_47660_n573;
  wire u2_u4__abc_47660_n574;
  wire u2_u4__abc_47660_n575;
  wire u2_u4__abc_47660_n576;
  wire u2_u4__abc_47660_n577;
  wire u2_u4__abc_47660_n578;
  wire u2_u4__abc_47660_n579;
  wire u2_u4__abc_47660_n580;
  wire u2_u4__abc_47660_n581;
  wire u2_u4__abc_47660_n582;
  wire u2_u4__abc_47660_n583;
  wire u2_u4__abc_47660_n584;
  wire u2_u4__abc_47660_n585;
  wire u2_u4__abc_47660_n586;
  wire u2_u4__abc_47660_n587;
  wire u2_u4__abc_47660_n588;
  wire u2_u4__abc_47660_n589;
  wire u2_u4__abc_47660_n590;
  wire u2_u4__abc_47660_n591;
  wire u2_u4__abc_47660_n592;
  wire u2_u4__abc_47660_n594;
  wire u2_u4__abc_47660_n595;
  wire u2_u4__abc_47660_n596;
  wire u2_u4__abc_47660_n597;
  wire u2_u4__abc_47660_n598;
  wire u2_u4__abc_47660_n599;
  wire u2_u4__abc_47660_n604;
  wire u2_u4__abc_47660_n605;
  wire u2_u4__abc_47660_n606;
  wire u2_u4__abc_47660_n607;
  wire u2_u4__abc_47660_n608;
  wire u2_u4__abc_47660_n610;
  wire u2_u4__abc_47660_n611;
  wire u2_u4__abc_47660_n612;
  wire u2_u4__abc_47660_n613;
  wire u2_u4__abc_47660_n614;
  wire u2_u4__abc_47660_n616;
  wire u2_u4__abc_47660_n617;
  wire u2_u4__abc_47660_n618;
  wire u2_u4__abc_47660_n619;
  wire u2_u4__abc_47660_n621;
  wire u2_u4__abc_47660_n622;
  wire u2_u4__abc_47660_n623;
  wire u2_u4__abc_47660_n624;
  wire u2_u4_b0_last_row_0_;
  wire u2_u4_b0_last_row_0__FF_INPUT;
  wire u2_u4_b0_last_row_10_;
  wire u2_u4_b0_last_row_10__FF_INPUT;
  wire u2_u4_b0_last_row_11_;
  wire u2_u4_b0_last_row_11__FF_INPUT;
  wire u2_u4_b0_last_row_12_;
  wire u2_u4_b0_last_row_12__FF_INPUT;
  wire u2_u4_b0_last_row_1_;
  wire u2_u4_b0_last_row_1__FF_INPUT;
  wire u2_u4_b0_last_row_2_;
  wire u2_u4_b0_last_row_2__FF_INPUT;
  wire u2_u4_b0_last_row_3_;
  wire u2_u4_b0_last_row_3__FF_INPUT;
  wire u2_u4_b0_last_row_4_;
  wire u2_u4_b0_last_row_4__FF_INPUT;
  wire u2_u4_b0_last_row_5_;
  wire u2_u4_b0_last_row_5__FF_INPUT;
  wire u2_u4_b0_last_row_6_;
  wire u2_u4_b0_last_row_6__FF_INPUT;
  wire u2_u4_b0_last_row_7_;
  wire u2_u4_b0_last_row_7__FF_INPUT;
  wire u2_u4_b0_last_row_8_;
  wire u2_u4_b0_last_row_8__FF_INPUT;
  wire u2_u4_b0_last_row_9_;
  wire u2_u4_b0_last_row_9__FF_INPUT;
  wire u2_u4_b1_last_row_0_;
  wire u2_u4_b1_last_row_0__FF_INPUT;
  wire u2_u4_b1_last_row_10_;
  wire u2_u4_b1_last_row_10__FF_INPUT;
  wire u2_u4_b1_last_row_11_;
  wire u2_u4_b1_last_row_11__FF_INPUT;
  wire u2_u4_b1_last_row_12_;
  wire u2_u4_b1_last_row_12__FF_INPUT;
  wire u2_u4_b1_last_row_1_;
  wire u2_u4_b1_last_row_1__FF_INPUT;
  wire u2_u4_b1_last_row_2_;
  wire u2_u4_b1_last_row_2__FF_INPUT;
  wire u2_u4_b1_last_row_3_;
  wire u2_u4_b1_last_row_3__FF_INPUT;
  wire u2_u4_b1_last_row_4_;
  wire u2_u4_b1_last_row_4__FF_INPUT;
  wire u2_u4_b1_last_row_5_;
  wire u2_u4_b1_last_row_5__FF_INPUT;
  wire u2_u4_b1_last_row_6_;
  wire u2_u4_b1_last_row_6__FF_INPUT;
  wire u2_u4_b1_last_row_7_;
  wire u2_u4_b1_last_row_7__FF_INPUT;
  wire u2_u4_b1_last_row_8_;
  wire u2_u4_b1_last_row_8__FF_INPUT;
  wire u2_u4_b1_last_row_9_;
  wire u2_u4_b1_last_row_9__FF_INPUT;
  wire u2_u4_b2_last_row_0_;
  wire u2_u4_b2_last_row_0__FF_INPUT;
  wire u2_u4_b2_last_row_10_;
  wire u2_u4_b2_last_row_10__FF_INPUT;
  wire u2_u4_b2_last_row_11_;
  wire u2_u4_b2_last_row_11__FF_INPUT;
  wire u2_u4_b2_last_row_12_;
  wire u2_u4_b2_last_row_12__FF_INPUT;
  wire u2_u4_b2_last_row_1_;
  wire u2_u4_b2_last_row_1__FF_INPUT;
  wire u2_u4_b2_last_row_2_;
  wire u2_u4_b2_last_row_2__FF_INPUT;
  wire u2_u4_b2_last_row_3_;
  wire u2_u4_b2_last_row_3__FF_INPUT;
  wire u2_u4_b2_last_row_4_;
  wire u2_u4_b2_last_row_4__FF_INPUT;
  wire u2_u4_b2_last_row_5_;
  wire u2_u4_b2_last_row_5__FF_INPUT;
  wire u2_u4_b2_last_row_6_;
  wire u2_u4_b2_last_row_6__FF_INPUT;
  wire u2_u4_b2_last_row_7_;
  wire u2_u4_b2_last_row_7__FF_INPUT;
  wire u2_u4_b2_last_row_8_;
  wire u2_u4_b2_last_row_8__FF_INPUT;
  wire u2_u4_b2_last_row_9_;
  wire u2_u4_b2_last_row_9__FF_INPUT;
  wire u2_u4_b3_last_row_0_;
  wire u2_u4_b3_last_row_0__FF_INPUT;
  wire u2_u4_b3_last_row_10_;
  wire u2_u4_b3_last_row_10__FF_INPUT;
  wire u2_u4_b3_last_row_11_;
  wire u2_u4_b3_last_row_11__FF_INPUT;
  wire u2_u4_b3_last_row_12_;
  wire u2_u4_b3_last_row_12__FF_INPUT;
  wire u2_u4_b3_last_row_1_;
  wire u2_u4_b3_last_row_1__FF_INPUT;
  wire u2_u4_b3_last_row_2_;
  wire u2_u4_b3_last_row_2__FF_INPUT;
  wire u2_u4_b3_last_row_3_;
  wire u2_u4_b3_last_row_3__FF_INPUT;
  wire u2_u4_b3_last_row_4_;
  wire u2_u4_b3_last_row_4__FF_INPUT;
  wire u2_u4_b3_last_row_5_;
  wire u2_u4_b3_last_row_5__FF_INPUT;
  wire u2_u4_b3_last_row_6_;
  wire u2_u4_b3_last_row_6__FF_INPUT;
  wire u2_u4_b3_last_row_7_;
  wire u2_u4_b3_last_row_7__FF_INPUT;
  wire u2_u4_b3_last_row_8_;
  wire u2_u4_b3_last_row_8__FF_INPUT;
  wire u2_u4_b3_last_row_9_;
  wire u2_u4_b3_last_row_9__FF_INPUT;
  wire u2_u4_bank0_open;
  wire u2_u4_bank0_open_FF_INPUT;
  wire u2_u4_bank1_open;
  wire u2_u4_bank1_open_FF_INPUT;
  wire u2_u4_bank2_open;
  wire u2_u4_bank2_open_FF_INPUT;
  wire u2_u4_bank3_open;
  wire u2_u4_bank3_open_FF_INPUT;
  wire u2_u5__abc_47660_n136;
  wire u2_u5__abc_47660_n137;
  wire u2_u5__abc_47660_n137_bF_buf0;
  wire u2_u5__abc_47660_n137_bF_buf1;
  wire u2_u5__abc_47660_n137_bF_buf2;
  wire u2_u5__abc_47660_n137_bF_buf3;
  wire u2_u5__abc_47660_n137_bF_buf4;
  wire u2_u5__abc_47660_n138;
  wire u2_u5__abc_47660_n139;
  wire u2_u5__abc_47660_n140;
  wire u2_u5__abc_47660_n141;
  wire u2_u5__abc_47660_n143;
  wire u2_u5__abc_47660_n144;
  wire u2_u5__abc_47660_n145;
  wire u2_u5__abc_47660_n146;
  wire u2_u5__abc_47660_n148;
  wire u2_u5__abc_47660_n149;
  wire u2_u5__abc_47660_n150;
  wire u2_u5__abc_47660_n151;
  wire u2_u5__abc_47660_n153;
  wire u2_u5__abc_47660_n154;
  wire u2_u5__abc_47660_n155;
  wire u2_u5__abc_47660_n156;
  wire u2_u5__abc_47660_n158;
  wire u2_u5__abc_47660_n159;
  wire u2_u5__abc_47660_n160;
  wire u2_u5__abc_47660_n161;
  wire u2_u5__abc_47660_n163;
  wire u2_u5__abc_47660_n164;
  wire u2_u5__abc_47660_n165;
  wire u2_u5__abc_47660_n166;
  wire u2_u5__abc_47660_n168;
  wire u2_u5__abc_47660_n169;
  wire u2_u5__abc_47660_n170;
  wire u2_u5__abc_47660_n171;
  wire u2_u5__abc_47660_n173;
  wire u2_u5__abc_47660_n174;
  wire u2_u5__abc_47660_n175;
  wire u2_u5__abc_47660_n176;
  wire u2_u5__abc_47660_n178;
  wire u2_u5__abc_47660_n179;
  wire u2_u5__abc_47660_n180;
  wire u2_u5__abc_47660_n181;
  wire u2_u5__abc_47660_n183;
  wire u2_u5__abc_47660_n184;
  wire u2_u5__abc_47660_n185;
  wire u2_u5__abc_47660_n186;
  wire u2_u5__abc_47660_n188;
  wire u2_u5__abc_47660_n189;
  wire u2_u5__abc_47660_n190;
  wire u2_u5__abc_47660_n191;
  wire u2_u5__abc_47660_n193;
  wire u2_u5__abc_47660_n194;
  wire u2_u5__abc_47660_n195;
  wire u2_u5__abc_47660_n196;
  wire u2_u5__abc_47660_n198;
  wire u2_u5__abc_47660_n199;
  wire u2_u5__abc_47660_n200;
  wire u2_u5__abc_47660_n201;
  wire u2_u5__abc_47660_n203;
  wire u2_u5__abc_47660_n204;
  wire u2_u5__abc_47660_n205;
  wire u2_u5__abc_47660_n206;
  wire u2_u5__abc_47660_n207;
  wire u2_u5__abc_47660_n208;
  wire u2_u5__abc_47660_n210;
  wire u2_u5__abc_47660_n211;
  wire u2_u5__abc_47660_n213;
  wire u2_u5__abc_47660_n214;
  wire u2_u5__abc_47660_n216;
  wire u2_u5__abc_47660_n217;
  wire u2_u5__abc_47660_n219;
  wire u2_u5__abc_47660_n220;
  wire u2_u5__abc_47660_n222;
  wire u2_u5__abc_47660_n223;
  wire u2_u5__abc_47660_n225;
  wire u2_u5__abc_47660_n226;
  wire u2_u5__abc_47660_n228;
  wire u2_u5__abc_47660_n229;
  wire u2_u5__abc_47660_n231;
  wire u2_u5__abc_47660_n232;
  wire u2_u5__abc_47660_n234;
  wire u2_u5__abc_47660_n235;
  wire u2_u5__abc_47660_n237;
  wire u2_u5__abc_47660_n238;
  wire u2_u5__abc_47660_n240;
  wire u2_u5__abc_47660_n241;
  wire u2_u5__abc_47660_n243;
  wire u2_u5__abc_47660_n244;
  wire u2_u5__abc_47660_n246;
  wire u2_u5__abc_47660_n247;
  wire u2_u5__abc_47660_n248;
  wire u2_u5__abc_47660_n249;
  wire u2_u5__abc_47660_n250;
  wire u2_u5__abc_47660_n251;
  wire u2_u5__abc_47660_n253;
  wire u2_u5__abc_47660_n254;
  wire u2_u5__abc_47660_n256;
  wire u2_u5__abc_47660_n257;
  wire u2_u5__abc_47660_n259;
  wire u2_u5__abc_47660_n260;
  wire u2_u5__abc_47660_n262;
  wire u2_u5__abc_47660_n263;
  wire u2_u5__abc_47660_n265;
  wire u2_u5__abc_47660_n266;
  wire u2_u5__abc_47660_n268;
  wire u2_u5__abc_47660_n269;
  wire u2_u5__abc_47660_n271;
  wire u2_u5__abc_47660_n272;
  wire u2_u5__abc_47660_n274;
  wire u2_u5__abc_47660_n275_1;
  wire u2_u5__abc_47660_n277;
  wire u2_u5__abc_47660_n278_1;
  wire u2_u5__abc_47660_n280;
  wire u2_u5__abc_47660_n281;
  wire u2_u5__abc_47660_n283_1;
  wire u2_u5__abc_47660_n284;
  wire u2_u5__abc_47660_n286_1;
  wire u2_u5__abc_47660_n287_1;
  wire u2_u5__abc_47660_n289;
  wire u2_u5__abc_47660_n290_1;
  wire u2_u5__abc_47660_n291;
  wire u2_u5__abc_47660_n292_1;
  wire u2_u5__abc_47660_n293;
  wire u2_u5__abc_47660_n295;
  wire u2_u5__abc_47660_n296_1;
  wire u2_u5__abc_47660_n298;
  wire u2_u5__abc_47660_n299;
  wire u2_u5__abc_47660_n301;
  wire u2_u5__abc_47660_n302;
  wire u2_u5__abc_47660_n304_1;
  wire u2_u5__abc_47660_n305;
  wire u2_u5__abc_47660_n305_1;
  wire u2_u5__abc_47660_n307;
  wire u2_u5__abc_47660_n308;
  wire u2_u5__abc_47660_n310;
  wire u2_u5__abc_47660_n311;
  wire u2_u5__abc_47660_n313;
  wire u2_u5__abc_47660_n314;
  wire u2_u5__abc_47660_n316;
  wire u2_u5__abc_47660_n317;
  wire u2_u5__abc_47660_n319;
  wire u2_u5__abc_47660_n320;
  wire u2_u5__abc_47660_n322;
  wire u2_u5__abc_47660_n323;
  wire u2_u5__abc_47660_n325;
  wire u2_u5__abc_47660_n326;
  wire u2_u5__abc_47660_n328;
  wire u2_u5__abc_47660_n329;
  wire u2_u5__abc_47660_n331;
  wire u2_u5__abc_47660_n332;
  wire u2_u5__abc_47660_n333;
  wire u2_u5__abc_47660_n334;
  wire u2_u5__abc_47660_n335;
  wire u2_u5__abc_47660_n336;
  wire u2_u5__abc_47660_n337;
  wire u2_u5__abc_47660_n338;
  wire u2_u5__abc_47660_n339;
  wire u2_u5__abc_47660_n340;
  wire u2_u5__abc_47660_n341;
  wire u2_u5__abc_47660_n342;
  wire u2_u5__abc_47660_n343;
  wire u2_u5__abc_47660_n344;
  wire u2_u5__abc_47660_n345;
  wire u2_u5__abc_47660_n346;
  wire u2_u5__abc_47660_n347;
  wire u2_u5__abc_47660_n348;
  wire u2_u5__abc_47660_n349;
  wire u2_u5__abc_47660_n350;
  wire u2_u5__abc_47660_n351;
  wire u2_u5__abc_47660_n352;
  wire u2_u5__abc_47660_n353;
  wire u2_u5__abc_47660_n354;
  wire u2_u5__abc_47660_n355;
  wire u2_u5__abc_47660_n356;
  wire u2_u5__abc_47660_n357;
  wire u2_u5__abc_47660_n358;
  wire u2_u5__abc_47660_n359;
  wire u2_u5__abc_47660_n360;
  wire u2_u5__abc_47660_n361;
  wire u2_u5__abc_47660_n362;
  wire u2_u5__abc_47660_n363;
  wire u2_u5__abc_47660_n364;
  wire u2_u5__abc_47660_n365;
  wire u2_u5__abc_47660_n366;
  wire u2_u5__abc_47660_n367;
  wire u2_u5__abc_47660_n368;
  wire u2_u5__abc_47660_n369;
  wire u2_u5__abc_47660_n370;
  wire u2_u5__abc_47660_n371;
  wire u2_u5__abc_47660_n372;
  wire u2_u5__abc_47660_n373;
  wire u2_u5__abc_47660_n374;
  wire u2_u5__abc_47660_n375;
  wire u2_u5__abc_47660_n376;
  wire u2_u5__abc_47660_n377;
  wire u2_u5__abc_47660_n378;
  wire u2_u5__abc_47660_n379;
  wire u2_u5__abc_47660_n380;
  wire u2_u5__abc_47660_n381;
  wire u2_u5__abc_47660_n382;
  wire u2_u5__abc_47660_n383;
  wire u2_u5__abc_47660_n384;
  wire u2_u5__abc_47660_n385;
  wire u2_u5__abc_47660_n386;
  wire u2_u5__abc_47660_n387;
  wire u2_u5__abc_47660_n388;
  wire u2_u5__abc_47660_n389;
  wire u2_u5__abc_47660_n390;
  wire u2_u5__abc_47660_n391;
  wire u2_u5__abc_47660_n392;
  wire u2_u5__abc_47660_n393;
  wire u2_u5__abc_47660_n394;
  wire u2_u5__abc_47660_n395;
  wire u2_u5__abc_47660_n396;
  wire u2_u5__abc_47660_n397;
  wire u2_u5__abc_47660_n398;
  wire u2_u5__abc_47660_n399;
  wire u2_u5__abc_47660_n400;
  wire u2_u5__abc_47660_n401;
  wire u2_u5__abc_47660_n402;
  wire u2_u5__abc_47660_n403;
  wire u2_u5__abc_47660_n404;
  wire u2_u5__abc_47660_n405;
  wire u2_u5__abc_47660_n406;
  wire u2_u5__abc_47660_n407;
  wire u2_u5__abc_47660_n408;
  wire u2_u5__abc_47660_n409;
  wire u2_u5__abc_47660_n410;
  wire u2_u5__abc_47660_n411;
  wire u2_u5__abc_47660_n412;
  wire u2_u5__abc_47660_n413;
  wire u2_u5__abc_47660_n414;
  wire u2_u5__abc_47660_n415;
  wire u2_u5__abc_47660_n416;
  wire u2_u5__abc_47660_n417;
  wire u2_u5__abc_47660_n418;
  wire u2_u5__abc_47660_n419;
  wire u2_u5__abc_47660_n420;
  wire u2_u5__abc_47660_n421;
  wire u2_u5__abc_47660_n422;
  wire u2_u5__abc_47660_n423;
  wire u2_u5__abc_47660_n424;
  wire u2_u5__abc_47660_n425;
  wire u2_u5__abc_47660_n426;
  wire u2_u5__abc_47660_n427;
  wire u2_u5__abc_47660_n428;
  wire u2_u5__abc_47660_n429;
  wire u2_u5__abc_47660_n430;
  wire u2_u5__abc_47660_n431;
  wire u2_u5__abc_47660_n432;
  wire u2_u5__abc_47660_n433;
  wire u2_u5__abc_47660_n434;
  wire u2_u5__abc_47660_n435;
  wire u2_u5__abc_47660_n436;
  wire u2_u5__abc_47660_n437;
  wire u2_u5__abc_47660_n438;
  wire u2_u5__abc_47660_n439;
  wire u2_u5__abc_47660_n440;
  wire u2_u5__abc_47660_n441;
  wire u2_u5__abc_47660_n442;
  wire u2_u5__abc_47660_n443;
  wire u2_u5__abc_47660_n444;
  wire u2_u5__abc_47660_n445;
  wire u2_u5__abc_47660_n446;
  wire u2_u5__abc_47660_n447;
  wire u2_u5__abc_47660_n448;
  wire u2_u5__abc_47660_n449;
  wire u2_u5__abc_47660_n450;
  wire u2_u5__abc_47660_n451;
  wire u2_u5__abc_47660_n452;
  wire u2_u5__abc_47660_n453;
  wire u2_u5__abc_47660_n454;
  wire u2_u5__abc_47660_n455;
  wire u2_u5__abc_47660_n456;
  wire u2_u5__abc_47660_n457;
  wire u2_u5__abc_47660_n458;
  wire u2_u5__abc_47660_n459;
  wire u2_u5__abc_47660_n460;
  wire u2_u5__abc_47660_n461;
  wire u2_u5__abc_47660_n462;
  wire u2_u5__abc_47660_n463;
  wire u2_u5__abc_47660_n464;
  wire u2_u5__abc_47660_n465;
  wire u2_u5__abc_47660_n466;
  wire u2_u5__abc_47660_n467;
  wire u2_u5__abc_47660_n468;
  wire u2_u5__abc_47660_n469;
  wire u2_u5__abc_47660_n470;
  wire u2_u5__abc_47660_n471;
  wire u2_u5__abc_47660_n472;
  wire u2_u5__abc_47660_n473;
  wire u2_u5__abc_47660_n474;
  wire u2_u5__abc_47660_n475;
  wire u2_u5__abc_47660_n476;
  wire u2_u5__abc_47660_n477;
  wire u2_u5__abc_47660_n478;
  wire u2_u5__abc_47660_n479;
  wire u2_u5__abc_47660_n480;
  wire u2_u5__abc_47660_n481;
  wire u2_u5__abc_47660_n482;
  wire u2_u5__abc_47660_n483;
  wire u2_u5__abc_47660_n484;
  wire u2_u5__abc_47660_n485;
  wire u2_u5__abc_47660_n486;
  wire u2_u5__abc_47660_n487;
  wire u2_u5__abc_47660_n488;
  wire u2_u5__abc_47660_n489;
  wire u2_u5__abc_47660_n490;
  wire u2_u5__abc_47660_n491;
  wire u2_u5__abc_47660_n492;
  wire u2_u5__abc_47660_n493;
  wire u2_u5__abc_47660_n494;
  wire u2_u5__abc_47660_n495;
  wire u2_u5__abc_47660_n496;
  wire u2_u5__abc_47660_n497;
  wire u2_u5__abc_47660_n498;
  wire u2_u5__abc_47660_n499;
  wire u2_u5__abc_47660_n500;
  wire u2_u5__abc_47660_n501;
  wire u2_u5__abc_47660_n502;
  wire u2_u5__abc_47660_n503;
  wire u2_u5__abc_47660_n504;
  wire u2_u5__abc_47660_n505;
  wire u2_u5__abc_47660_n506;
  wire u2_u5__abc_47660_n507;
  wire u2_u5__abc_47660_n508;
  wire u2_u5__abc_47660_n509;
  wire u2_u5__abc_47660_n510;
  wire u2_u5__abc_47660_n511;
  wire u2_u5__abc_47660_n512;
  wire u2_u5__abc_47660_n513;
  wire u2_u5__abc_47660_n514;
  wire u2_u5__abc_47660_n515;
  wire u2_u5__abc_47660_n516;
  wire u2_u5__abc_47660_n517;
  wire u2_u5__abc_47660_n518;
  wire u2_u5__abc_47660_n519;
  wire u2_u5__abc_47660_n520;
  wire u2_u5__abc_47660_n521;
  wire u2_u5__abc_47660_n522;
  wire u2_u5__abc_47660_n523;
  wire u2_u5__abc_47660_n524;
  wire u2_u5__abc_47660_n525;
  wire u2_u5__abc_47660_n526;
  wire u2_u5__abc_47660_n527;
  wire u2_u5__abc_47660_n528;
  wire u2_u5__abc_47660_n529;
  wire u2_u5__abc_47660_n530;
  wire u2_u5__abc_47660_n531;
  wire u2_u5__abc_47660_n532;
  wire u2_u5__abc_47660_n533;
  wire u2_u5__abc_47660_n534;
  wire u2_u5__abc_47660_n535;
  wire u2_u5__abc_47660_n536;
  wire u2_u5__abc_47660_n537;
  wire u2_u5__abc_47660_n538;
  wire u2_u5__abc_47660_n539;
  wire u2_u5__abc_47660_n540;
  wire u2_u5__abc_47660_n541;
  wire u2_u5__abc_47660_n542;
  wire u2_u5__abc_47660_n543;
  wire u2_u5__abc_47660_n544;
  wire u2_u5__abc_47660_n545;
  wire u2_u5__abc_47660_n546;
  wire u2_u5__abc_47660_n547;
  wire u2_u5__abc_47660_n548;
  wire u2_u5__abc_47660_n549;
  wire u2_u5__abc_47660_n550;
  wire u2_u5__abc_47660_n551;
  wire u2_u5__abc_47660_n552;
  wire u2_u5__abc_47660_n553;
  wire u2_u5__abc_47660_n554;
  wire u2_u5__abc_47660_n555;
  wire u2_u5__abc_47660_n556;
  wire u2_u5__abc_47660_n557;
  wire u2_u5__abc_47660_n558;
  wire u2_u5__abc_47660_n559;
  wire u2_u5__abc_47660_n560;
  wire u2_u5__abc_47660_n561;
  wire u2_u5__abc_47660_n562;
  wire u2_u5__abc_47660_n563;
  wire u2_u5__abc_47660_n564;
  wire u2_u5__abc_47660_n565;
  wire u2_u5__abc_47660_n566;
  wire u2_u5__abc_47660_n567;
  wire u2_u5__abc_47660_n568;
  wire u2_u5__abc_47660_n569;
  wire u2_u5__abc_47660_n570;
  wire u2_u5__abc_47660_n571;
  wire u2_u5__abc_47660_n572;
  wire u2_u5__abc_47660_n573;
  wire u2_u5__abc_47660_n574;
  wire u2_u5__abc_47660_n575;
  wire u2_u5__abc_47660_n576;
  wire u2_u5__abc_47660_n577;
  wire u2_u5__abc_47660_n578;
  wire u2_u5__abc_47660_n579;
  wire u2_u5__abc_47660_n580;
  wire u2_u5__abc_47660_n581;
  wire u2_u5__abc_47660_n582;
  wire u2_u5__abc_47660_n583;
  wire u2_u5__abc_47660_n584;
  wire u2_u5__abc_47660_n585;
  wire u2_u5__abc_47660_n586;
  wire u2_u5__abc_47660_n587;
  wire u2_u5__abc_47660_n588;
  wire u2_u5__abc_47660_n589;
  wire u2_u5__abc_47660_n590;
  wire u2_u5__abc_47660_n591;
  wire u2_u5__abc_47660_n592;
  wire u2_u5__abc_47660_n594;
  wire u2_u5__abc_47660_n595;
  wire u2_u5__abc_47660_n596;
  wire u2_u5__abc_47660_n597;
  wire u2_u5__abc_47660_n598;
  wire u2_u5__abc_47660_n599;
  wire u2_u5__abc_47660_n604;
  wire u2_u5__abc_47660_n605;
  wire u2_u5__abc_47660_n606;
  wire u2_u5__abc_47660_n607;
  wire u2_u5__abc_47660_n608;
  wire u2_u5__abc_47660_n610;
  wire u2_u5__abc_47660_n611;
  wire u2_u5__abc_47660_n612;
  wire u2_u5__abc_47660_n613;
  wire u2_u5__abc_47660_n614;
  wire u2_u5__abc_47660_n616;
  wire u2_u5__abc_47660_n617;
  wire u2_u5__abc_47660_n618;
  wire u2_u5__abc_47660_n619;
  wire u2_u5__abc_47660_n621;
  wire u2_u5__abc_47660_n622;
  wire u2_u5__abc_47660_n623;
  wire u2_u5__abc_47660_n624;
  wire u2_u5_b0_last_row_0_;
  wire u2_u5_b0_last_row_0__FF_INPUT;
  wire u2_u5_b0_last_row_10_;
  wire u2_u5_b0_last_row_10__FF_INPUT;
  wire u2_u5_b0_last_row_11_;
  wire u2_u5_b0_last_row_11__FF_INPUT;
  wire u2_u5_b0_last_row_12_;
  wire u2_u5_b0_last_row_12__FF_INPUT;
  wire u2_u5_b0_last_row_1_;
  wire u2_u5_b0_last_row_1__FF_INPUT;
  wire u2_u5_b0_last_row_2_;
  wire u2_u5_b0_last_row_2__FF_INPUT;
  wire u2_u5_b0_last_row_3_;
  wire u2_u5_b0_last_row_3__FF_INPUT;
  wire u2_u5_b0_last_row_4_;
  wire u2_u5_b0_last_row_4__FF_INPUT;
  wire u2_u5_b0_last_row_5_;
  wire u2_u5_b0_last_row_5__FF_INPUT;
  wire u2_u5_b0_last_row_6_;
  wire u2_u5_b0_last_row_6__FF_INPUT;
  wire u2_u5_b0_last_row_7_;
  wire u2_u5_b0_last_row_7__FF_INPUT;
  wire u2_u5_b0_last_row_8_;
  wire u2_u5_b0_last_row_8__FF_INPUT;
  wire u2_u5_b0_last_row_9_;
  wire u2_u5_b0_last_row_9__FF_INPUT;
  wire u2_u5_b1_last_row_0_;
  wire u2_u5_b1_last_row_0__FF_INPUT;
  wire u2_u5_b1_last_row_10_;
  wire u2_u5_b1_last_row_10__FF_INPUT;
  wire u2_u5_b1_last_row_11_;
  wire u2_u5_b1_last_row_11__FF_INPUT;
  wire u2_u5_b1_last_row_12_;
  wire u2_u5_b1_last_row_12__FF_INPUT;
  wire u2_u5_b1_last_row_1_;
  wire u2_u5_b1_last_row_1__FF_INPUT;
  wire u2_u5_b1_last_row_2_;
  wire u2_u5_b1_last_row_2__FF_INPUT;
  wire u2_u5_b1_last_row_3_;
  wire u2_u5_b1_last_row_3__FF_INPUT;
  wire u2_u5_b1_last_row_4_;
  wire u2_u5_b1_last_row_4__FF_INPUT;
  wire u2_u5_b1_last_row_5_;
  wire u2_u5_b1_last_row_5__FF_INPUT;
  wire u2_u5_b1_last_row_6_;
  wire u2_u5_b1_last_row_6__FF_INPUT;
  wire u2_u5_b1_last_row_7_;
  wire u2_u5_b1_last_row_7__FF_INPUT;
  wire u2_u5_b1_last_row_8_;
  wire u2_u5_b1_last_row_8__FF_INPUT;
  wire u2_u5_b1_last_row_9_;
  wire u2_u5_b1_last_row_9__FF_INPUT;
  wire u2_u5_b2_last_row_0_;
  wire u2_u5_b2_last_row_0__FF_INPUT;
  wire u2_u5_b2_last_row_10_;
  wire u2_u5_b2_last_row_10__FF_INPUT;
  wire u2_u5_b2_last_row_11_;
  wire u2_u5_b2_last_row_11__FF_INPUT;
  wire u2_u5_b2_last_row_12_;
  wire u2_u5_b2_last_row_12__FF_INPUT;
  wire u2_u5_b2_last_row_1_;
  wire u2_u5_b2_last_row_1__FF_INPUT;
  wire u2_u5_b2_last_row_2_;
  wire u2_u5_b2_last_row_2__FF_INPUT;
  wire u2_u5_b2_last_row_3_;
  wire u2_u5_b2_last_row_3__FF_INPUT;
  wire u2_u5_b2_last_row_4_;
  wire u2_u5_b2_last_row_4__FF_INPUT;
  wire u2_u5_b2_last_row_5_;
  wire u2_u5_b2_last_row_5__FF_INPUT;
  wire u2_u5_b2_last_row_6_;
  wire u2_u5_b2_last_row_6__FF_INPUT;
  wire u2_u5_b2_last_row_7_;
  wire u2_u5_b2_last_row_7__FF_INPUT;
  wire u2_u5_b2_last_row_8_;
  wire u2_u5_b2_last_row_8__FF_INPUT;
  wire u2_u5_b2_last_row_9_;
  wire u2_u5_b2_last_row_9__FF_INPUT;
  wire u2_u5_b3_last_row_0_;
  wire u2_u5_b3_last_row_0__FF_INPUT;
  wire u2_u5_b3_last_row_10_;
  wire u2_u5_b3_last_row_10__FF_INPUT;
  wire u2_u5_b3_last_row_11_;
  wire u2_u5_b3_last_row_11__FF_INPUT;
  wire u2_u5_b3_last_row_12_;
  wire u2_u5_b3_last_row_12__FF_INPUT;
  wire u2_u5_b3_last_row_1_;
  wire u2_u5_b3_last_row_1__FF_INPUT;
  wire u2_u5_b3_last_row_2_;
  wire u2_u5_b3_last_row_2__FF_INPUT;
  wire u2_u5_b3_last_row_3_;
  wire u2_u5_b3_last_row_3__FF_INPUT;
  wire u2_u5_b3_last_row_4_;
  wire u2_u5_b3_last_row_4__FF_INPUT;
  wire u2_u5_b3_last_row_5_;
  wire u2_u5_b3_last_row_5__FF_INPUT;
  wire u2_u5_b3_last_row_6_;
  wire u2_u5_b3_last_row_6__FF_INPUT;
  wire u2_u5_b3_last_row_7_;
  wire u2_u5_b3_last_row_7__FF_INPUT;
  wire u2_u5_b3_last_row_8_;
  wire u2_u5_b3_last_row_8__FF_INPUT;
  wire u2_u5_b3_last_row_9_;
  wire u2_u5_b3_last_row_9__FF_INPUT;
  wire u2_u5_bank0_open;
  wire u2_u5_bank0_open_FF_INPUT;
  wire u2_u5_bank1_open;
  wire u2_u5_bank1_open_FF_INPUT;
  wire u2_u5_bank2_open;
  wire u2_u5_bank2_open_FF_INPUT;
  wire u2_u5_bank3_open;
  wire u2_u5_bank3_open_FF_INPUT;
  wire u3__abc_46775_n1000;
  wire u3__abc_46775_n1001;
  wire u3__abc_46775_n1002;
  wire u3__abc_46775_n1003;
  wire u3__abc_46775_n1004;
  wire u3__abc_46775_n1005;
  wire u3__abc_46775_n1006;
  wire u3__abc_46775_n1007;
  wire u3__abc_46775_n1008;
  wire u3__abc_46775_n1009;
  wire u3__abc_46775_n1010;
  wire u3__abc_46775_n1011;
  wire u3__abc_46775_n1012;
  wire u3__abc_46775_n1013;
  wire u3__abc_46775_n1014;
  wire u3__abc_46775_n1015;
  wire u3__abc_46775_n1016;
  wire u3__abc_46775_n1017;
  wire u3__abc_46775_n1018;
  wire u3__abc_46775_n1019;
  wire u3__abc_46775_n1020;
  wire u3__abc_46775_n1021;
  wire u3__abc_46775_n1022;
  wire u3__abc_46775_n1023;
  wire u3__abc_46775_n1024;
  wire u3__abc_46775_n1025;
  wire u3__abc_46775_n1026;
  wire u3__abc_46775_n1027;
  wire u3__abc_46775_n1028;
  wire u3__abc_46775_n1029;
  wire u3__abc_46775_n1030;
  wire u3__abc_46775_n1031;
  wire u3__abc_46775_n1032;
  wire u3__abc_46775_n275;
  wire u3__abc_46775_n275_bF_buf0;
  wire u3__abc_46775_n275_bF_buf1;
  wire u3__abc_46775_n275_bF_buf2;
  wire u3__abc_46775_n275_bF_buf3;
  wire u3__abc_46775_n275_bF_buf4;
  wire u3__abc_46775_n276;
  wire u3__abc_46775_n277_1;
  wire u3__abc_46775_n277_1_bF_buf0;
  wire u3__abc_46775_n277_1_bF_buf1;
  wire u3__abc_46775_n277_1_bF_buf2;
  wire u3__abc_46775_n277_1_bF_buf3;
  wire u3__abc_46775_n277_1_bF_buf4;
  wire u3__abc_46775_n277_1_bF_buf5;
  wire u3__abc_46775_n278_1;
  wire u3__abc_46775_n279;
  wire u3__abc_46775_n279_bF_buf0;
  wire u3__abc_46775_n279_bF_buf1;
  wire u3__abc_46775_n279_bF_buf2;
  wire u3__abc_46775_n279_bF_buf3;
  wire u3__abc_46775_n279_bF_buf4;
  wire u3__abc_46775_n279_bF_buf5;
  wire u3__abc_46775_n280;
  wire u3__abc_46775_n281_1;
  wire u3__abc_46775_n282_1;
  wire u3__abc_46775_n283;
  wire u3__abc_46775_n284;
  wire u3__abc_46775_n285_1;
  wire u3__abc_46775_n286_1;
  wire u3__abc_46775_n287_1;
  wire u3__abc_46775_n288;
  wire u3__abc_46775_n289;
  wire u3__abc_46775_n290_1;
  wire u3__abc_46775_n291_1;
  wire u3__abc_46775_n292_1;
  wire u3__abc_46775_n293;
  wire u3__abc_46775_n294;
  wire u3__abc_46775_n295_1;
  wire u3__abc_46775_n296_1;
  wire u3__abc_46775_n297_1;
  wire u3__abc_46775_n298;
  wire u3__abc_46775_n299;
  wire u3__abc_46775_n300_1;
  wire u3__abc_46775_n301_1;
  wire u3__abc_46775_n302_1;
  wire u3__abc_46775_n303;
  wire u3__abc_46775_n304;
  wire u3__abc_46775_n305_1;
  wire u3__abc_46775_n306_1;
  wire u3__abc_46775_n307_1;
  wire u3__abc_46775_n308;
  wire u3__abc_46775_n309;
  wire u3__abc_46775_n310_1;
  wire u3__abc_46775_n311_1;
  wire u3__abc_46775_n312_1;
  wire u3__abc_46775_n313;
  wire u3__abc_46775_n315_1;
  wire u3__abc_46775_n316_1;
  wire u3__abc_46775_n317_1;
  wire u3__abc_46775_n318;
  wire u3__abc_46775_n319;
  wire u3__abc_46775_n320_1;
  wire u3__abc_46775_n321_1;
  wire u3__abc_46775_n322_1;
  wire u3__abc_46775_n323;
  wire u3__abc_46775_n324;
  wire u3__abc_46775_n325_1;
  wire u3__abc_46775_n326_1;
  wire u3__abc_46775_n327_1;
  wire u3__abc_46775_n328;
  wire u3__abc_46775_n329;
  wire u3__abc_46775_n330_1;
  wire u3__abc_46775_n331_1;
  wire u3__abc_46775_n332_1;
  wire u3__abc_46775_n333;
  wire u3__abc_46775_n334;
  wire u3__abc_46775_n335_1;
  wire u3__abc_46775_n336_1;
  wire u3__abc_46775_n337_1;
  wire u3__abc_46775_n338;
  wire u3__abc_46775_n339;
  wire u3__abc_46775_n340_1;
  wire u3__abc_46775_n341_1;
  wire u3__abc_46775_n342_1;
  wire u3__abc_46775_n343;
  wire u3__abc_46775_n344;
  wire u3__abc_46775_n345_1;
  wire u3__abc_46775_n346_1;
  wire u3__abc_46775_n347_1;
  wire u3__abc_46775_n348;
  wire u3__abc_46775_n349;
  wire u3__abc_46775_n351_1;
  wire u3__abc_46775_n352_1;
  wire u3__abc_46775_n353;
  wire u3__abc_46775_n354;
  wire u3__abc_46775_n355_1;
  wire u3__abc_46775_n356_1;
  wire u3__abc_46775_n357_1;
  wire u3__abc_46775_n358;
  wire u3__abc_46775_n359;
  wire u3__abc_46775_n360_1;
  wire u3__abc_46775_n361_1;
  wire u3__abc_46775_n362_1;
  wire u3__abc_46775_n363;
  wire u3__abc_46775_n364;
  wire u3__abc_46775_n365_1;
  wire u3__abc_46775_n366_1;
  wire u3__abc_46775_n367_1;
  wire u3__abc_46775_n368_1;
  wire u3__abc_46775_n369;
  wire u3__abc_46775_n370_1;
  wire u3__abc_46775_n371_1;
  wire u3__abc_46775_n372_1;
  wire u3__abc_46775_n373_1;
  wire u3__abc_46775_n374;
  wire u3__abc_46775_n375;
  wire u3__abc_46775_n376;
  wire u3__abc_46775_n377;
  wire u3__abc_46775_n378;
  wire u3__abc_46775_n379;
  wire u3__abc_46775_n380;
  wire u3__abc_46775_n381_1;
  wire u3__abc_46775_n382;
  wire u3__abc_46775_n383;
  wire u3__abc_46775_n384;
  wire u3__abc_46775_n385;
  wire u3__abc_46775_n387;
  wire u3__abc_46775_n388;
  wire u3__abc_46775_n389;
  wire u3__abc_46775_n390_1;
  wire u3__abc_46775_n391;
  wire u3__abc_46775_n392_1;
  wire u3__abc_46775_n393_1;
  wire u3__abc_46775_n394;
  wire u3__abc_46775_n395;
  wire u3__abc_46775_n396;
  wire u3__abc_46775_n397;
  wire u3__abc_46775_n398;
  wire u3__abc_46775_n399;
  wire u3__abc_46775_n400;
  wire u3__abc_46775_n401;
  wire u3__abc_46775_n402_1;
  wire u3__abc_46775_n403;
  wire u3__abc_46775_n404;
  wire u3__abc_46775_n405;
  wire u3__abc_46775_n406;
  wire u3__abc_46775_n407;
  wire u3__abc_46775_n408;
  wire u3__abc_46775_n409;
  wire u3__abc_46775_n410;
  wire u3__abc_46775_n411_1;
  wire u3__abc_46775_n412;
  wire u3__abc_46775_n413_1;
  wire u3__abc_46775_n414_1;
  wire u3__abc_46775_n415;
  wire u3__abc_46775_n416_1;
  wire u3__abc_46775_n417;
  wire u3__abc_46775_n418;
  wire u3__abc_46775_n419_1;
  wire u3__abc_46775_n420;
  wire u3__abc_46775_n421_1;
  wire u3__abc_46775_n423;
  wire u3__abc_46775_n424;
  wire u3__abc_46775_n425;
  wire u3__abc_46775_n427;
  wire u3__abc_46775_n428;
  wire u3__abc_46775_n430;
  wire u3__abc_46775_n431;
  wire u3__abc_46775_n433;
  wire u3__abc_46775_n434;
  wire u3__abc_46775_n436;
  wire u3__abc_46775_n437;
  wire u3__abc_46775_n439;
  wire u3__abc_46775_n440;
  wire u3__abc_46775_n442;
  wire u3__abc_46775_n443;
  wire u3__abc_46775_n445;
  wire u3__abc_46775_n446;
  wire u3__abc_46775_n448;
  wire u3__abc_46775_n448_bF_buf0;
  wire u3__abc_46775_n448_bF_buf1;
  wire u3__abc_46775_n448_bF_buf2;
  wire u3__abc_46775_n448_bF_buf3;
  wire u3__abc_46775_n449;
  wire u3__abc_46775_n450;
  wire u3__abc_46775_n450_bF_buf0;
  wire u3__abc_46775_n450_bF_buf1;
  wire u3__abc_46775_n450_bF_buf2;
  wire u3__abc_46775_n450_bF_buf3;
  wire u3__abc_46775_n451;
  wire u3__abc_46775_n452;
  wire u3__abc_46775_n452_bF_buf0;
  wire u3__abc_46775_n452_bF_buf1;
  wire u3__abc_46775_n452_bF_buf2;
  wire u3__abc_46775_n452_bF_buf3;
  wire u3__abc_46775_n453;
  wire u3__abc_46775_n454;
  wire u3__abc_46775_n455;
  wire u3__abc_46775_n456;
  wire u3__abc_46775_n457;
  wire u3__abc_46775_n458;
  wire u3__abc_46775_n459;
  wire u3__abc_46775_n460;
  wire u3__abc_46775_n462;
  wire u3__abc_46775_n463;
  wire u3__abc_46775_n464;
  wire u3__abc_46775_n465;
  wire u3__abc_46775_n466;
  wire u3__abc_46775_n468;
  wire u3__abc_46775_n469;
  wire u3__abc_46775_n470;
  wire u3__abc_46775_n471;
  wire u3__abc_46775_n472;
  wire u3__abc_46775_n474;
  wire u3__abc_46775_n475;
  wire u3__abc_46775_n476;
  wire u3__abc_46775_n477;
  wire u3__abc_46775_n478;
  wire u3__abc_46775_n480;
  wire u3__abc_46775_n481;
  wire u3__abc_46775_n482;
  wire u3__abc_46775_n483;
  wire u3__abc_46775_n484;
  wire u3__abc_46775_n486;
  wire u3__abc_46775_n487;
  wire u3__abc_46775_n488;
  wire u3__abc_46775_n489;
  wire u3__abc_46775_n490;
  wire u3__abc_46775_n492;
  wire u3__abc_46775_n493;
  wire u3__abc_46775_n494;
  wire u3__abc_46775_n495;
  wire u3__abc_46775_n496;
  wire u3__abc_46775_n498;
  wire u3__abc_46775_n499;
  wire u3__abc_46775_n500;
  wire u3__abc_46775_n501;
  wire u3__abc_46775_n502;
  wire u3__abc_46775_n504;
  wire u3__abc_46775_n505;
  wire u3__abc_46775_n506;
  wire u3__abc_46775_n508;
  wire u3__abc_46775_n509;
  wire u3__abc_46775_n511;
  wire u3__abc_46775_n512;
  wire u3__abc_46775_n514;
  wire u3__abc_46775_n515;
  wire u3__abc_46775_n517;
  wire u3__abc_46775_n518;
  wire u3__abc_46775_n520;
  wire u3__abc_46775_n521;
  wire u3__abc_46775_n523;
  wire u3__abc_46775_n524;
  wire u3__abc_46775_n526;
  wire u3__abc_46775_n527;
  wire u3__abc_46775_n529;
  wire u3__abc_46775_n530;
  wire u3__abc_46775_n532;
  wire u3__abc_46775_n533;
  wire u3__abc_46775_n535;
  wire u3__abc_46775_n536;
  wire u3__abc_46775_n538;
  wire u3__abc_46775_n539;
  wire u3__abc_46775_n541;
  wire u3__abc_46775_n542;
  wire u3__abc_46775_n544;
  wire u3__abc_46775_n545;
  wire u3__abc_46775_n547;
  wire u3__abc_46775_n548;
  wire u3__abc_46775_n550;
  wire u3__abc_46775_n551;
  wire u3__abc_46775_n553;
  wire u3__abc_46775_n554;
  wire u3__abc_46775_n556;
  wire u3__abc_46775_n557;
  wire u3__abc_46775_n559;
  wire u3__abc_46775_n560;
  wire u3__abc_46775_n562;
  wire u3__abc_46775_n563;
  wire u3__abc_46775_n565;
  wire u3__abc_46775_n566;
  wire u3__abc_46775_n568;
  wire u3__abc_46775_n569;
  wire u3__abc_46775_n571;
  wire u3__abc_46775_n572;
  wire u3__abc_46775_n574;
  wire u3__abc_46775_n575;
  wire u3__abc_46775_n577;
  wire u3__abc_46775_n578;
  wire u3__abc_46775_n580;
  wire u3__abc_46775_n581;
  wire u3__abc_46775_n583;
  wire u3__abc_46775_n584;
  wire u3__abc_46775_n586;
  wire u3__abc_46775_n587;
  wire u3__abc_46775_n589;
  wire u3__abc_46775_n590;
  wire u3__abc_46775_n592;
  wire u3__abc_46775_n593;
  wire u3__abc_46775_n595;
  wire u3__abc_46775_n596;
  wire u3__abc_46775_n598;
  wire u3__abc_46775_n599;
  wire u3__abc_46775_n601;
  wire u3__abc_46775_n602;
  wire u3__abc_46775_n604;
  wire u3__abc_46775_n605;
  wire u3__abc_46775_n607;
  wire u3__abc_46775_n608;
  wire u3__abc_46775_n610;
  wire u3__abc_46775_n611;
  wire u3__abc_46775_n613;
  wire u3__abc_46775_n614;
  wire u3__abc_46775_n616;
  wire u3__abc_46775_n617;
  wire u3__abc_46775_n619;
  wire u3__abc_46775_n620;
  wire u3__abc_46775_n622;
  wire u3__abc_46775_n623;
  wire u3__abc_46775_n625;
  wire u3__abc_46775_n625_bF_buf0;
  wire u3__abc_46775_n625_bF_buf1;
  wire u3__abc_46775_n625_bF_buf2;
  wire u3__abc_46775_n625_bF_buf3;
  wire u3__abc_46775_n625_bF_buf4;
  wire u3__abc_46775_n626;
  wire u3__abc_46775_n627;
  wire u3__abc_46775_n628;
  wire u3__abc_46775_n629;
  wire u3__abc_46775_n630;
  wire u3__abc_46775_n632;
  wire u3__abc_46775_n633;
  wire u3__abc_46775_n634;
  wire u3__abc_46775_n635;
  wire u3__abc_46775_n636;
  wire u3__abc_46775_n638;
  wire u3__abc_46775_n639;
  wire u3__abc_46775_n640;
  wire u3__abc_46775_n641;
  wire u3__abc_46775_n642;
  wire u3__abc_46775_n644;
  wire u3__abc_46775_n645;
  wire u3__abc_46775_n646;
  wire u3__abc_46775_n647;
  wire u3__abc_46775_n648;
  wire u3__abc_46775_n650;
  wire u3__abc_46775_n651;
  wire u3__abc_46775_n652;
  wire u3__abc_46775_n653;
  wire u3__abc_46775_n654;
  wire u3__abc_46775_n656;
  wire u3__abc_46775_n657;
  wire u3__abc_46775_n658;
  wire u3__abc_46775_n659;
  wire u3__abc_46775_n660;
  wire u3__abc_46775_n662;
  wire u3__abc_46775_n663;
  wire u3__abc_46775_n664;
  wire u3__abc_46775_n665;
  wire u3__abc_46775_n666;
  wire u3__abc_46775_n668;
  wire u3__abc_46775_n669;
  wire u3__abc_46775_n670;
  wire u3__abc_46775_n671;
  wire u3__abc_46775_n672;
  wire u3__abc_46775_n674;
  wire u3__abc_46775_n675;
  wire u3__abc_46775_n676;
  wire u3__abc_46775_n677;
  wire u3__abc_46775_n678;
  wire u3__abc_46775_n680;
  wire u3__abc_46775_n681;
  wire u3__abc_46775_n682;
  wire u3__abc_46775_n683;
  wire u3__abc_46775_n684;
  wire u3__abc_46775_n686;
  wire u3__abc_46775_n687;
  wire u3__abc_46775_n688;
  wire u3__abc_46775_n689;
  wire u3__abc_46775_n690;
  wire u3__abc_46775_n692;
  wire u3__abc_46775_n693;
  wire u3__abc_46775_n694;
  wire u3__abc_46775_n695;
  wire u3__abc_46775_n696;
  wire u3__abc_46775_n698;
  wire u3__abc_46775_n699;
  wire u3__abc_46775_n700;
  wire u3__abc_46775_n701;
  wire u3__abc_46775_n702;
  wire u3__abc_46775_n704;
  wire u3__abc_46775_n705;
  wire u3__abc_46775_n706;
  wire u3__abc_46775_n707;
  wire u3__abc_46775_n708;
  wire u3__abc_46775_n710;
  wire u3__abc_46775_n711;
  wire u3__abc_46775_n712;
  wire u3__abc_46775_n713;
  wire u3__abc_46775_n714;
  wire u3__abc_46775_n716;
  wire u3__abc_46775_n717;
  wire u3__abc_46775_n718;
  wire u3__abc_46775_n719;
  wire u3__abc_46775_n720;
  wire u3__abc_46775_n722;
  wire u3__abc_46775_n723;
  wire u3__abc_46775_n724;
  wire u3__abc_46775_n725;
  wire u3__abc_46775_n726;
  wire u3__abc_46775_n727;
  wire u3__abc_46775_n728;
  wire u3__abc_46775_n730;
  wire u3__abc_46775_n731;
  wire u3__abc_46775_n732;
  wire u3__abc_46775_n733;
  wire u3__abc_46775_n734;
  wire u3__abc_46775_n735;
  wire u3__abc_46775_n736;
  wire u3__abc_46775_n738;
  wire u3__abc_46775_n739;
  wire u3__abc_46775_n740;
  wire u3__abc_46775_n741;
  wire u3__abc_46775_n742;
  wire u3__abc_46775_n743;
  wire u3__abc_46775_n744;
  wire u3__abc_46775_n746;
  wire u3__abc_46775_n747;
  wire u3__abc_46775_n748;
  wire u3__abc_46775_n749;
  wire u3__abc_46775_n750;
  wire u3__abc_46775_n751;
  wire u3__abc_46775_n752;
  wire u3__abc_46775_n754;
  wire u3__abc_46775_n755;
  wire u3__abc_46775_n756;
  wire u3__abc_46775_n757;
  wire u3__abc_46775_n758;
  wire u3__abc_46775_n759;
  wire u3__abc_46775_n760;
  wire u3__abc_46775_n762;
  wire u3__abc_46775_n763;
  wire u3__abc_46775_n764;
  wire u3__abc_46775_n765;
  wire u3__abc_46775_n766;
  wire u3__abc_46775_n767;
  wire u3__abc_46775_n768;
  wire u3__abc_46775_n770;
  wire u3__abc_46775_n771;
  wire u3__abc_46775_n772;
  wire u3__abc_46775_n773;
  wire u3__abc_46775_n774;
  wire u3__abc_46775_n775;
  wire u3__abc_46775_n776;
  wire u3__abc_46775_n778;
  wire u3__abc_46775_n779;
  wire u3__abc_46775_n780;
  wire u3__abc_46775_n781;
  wire u3__abc_46775_n782;
  wire u3__abc_46775_n783;
  wire u3__abc_46775_n784;
  wire u3__abc_46775_n786;
  wire u3__abc_46775_n787;
  wire u3__abc_46775_n788;
  wire u3__abc_46775_n789;
  wire u3__abc_46775_n790;
  wire u3__abc_46775_n791;
  wire u3__abc_46775_n792;
  wire u3__abc_46775_n794;
  wire u3__abc_46775_n795;
  wire u3__abc_46775_n796;
  wire u3__abc_46775_n797;
  wire u3__abc_46775_n798;
  wire u3__abc_46775_n799;
  wire u3__abc_46775_n800;
  wire u3__abc_46775_n802;
  wire u3__abc_46775_n803;
  wire u3__abc_46775_n804;
  wire u3__abc_46775_n805;
  wire u3__abc_46775_n806;
  wire u3__abc_46775_n807;
  wire u3__abc_46775_n808;
  wire u3__abc_46775_n810;
  wire u3__abc_46775_n811;
  wire u3__abc_46775_n812;
  wire u3__abc_46775_n813;
  wire u3__abc_46775_n814;
  wire u3__abc_46775_n815;
  wire u3__abc_46775_n816;
  wire u3__abc_46775_n818;
  wire u3__abc_46775_n819;
  wire u3__abc_46775_n820;
  wire u3__abc_46775_n821;
  wire u3__abc_46775_n822;
  wire u3__abc_46775_n823;
  wire u3__abc_46775_n824;
  wire u3__abc_46775_n826;
  wire u3__abc_46775_n827;
  wire u3__abc_46775_n828;
  wire u3__abc_46775_n829;
  wire u3__abc_46775_n830;
  wire u3__abc_46775_n831;
  wire u3__abc_46775_n832;
  wire u3__abc_46775_n834;
  wire u3__abc_46775_n835;
  wire u3__abc_46775_n836;
  wire u3__abc_46775_n837;
  wire u3__abc_46775_n838;
  wire u3__abc_46775_n839;
  wire u3__abc_46775_n840;
  wire u3__abc_46775_n842;
  wire u3__abc_46775_n843;
  wire u3__abc_46775_n844;
  wire u3__abc_46775_n845;
  wire u3__abc_46775_n846;
  wire u3__abc_46775_n847;
  wire u3__abc_46775_n848;
  wire u3__abc_46775_n850;
  wire u3__abc_46775_n851;
  wire u3__abc_46775_n854;
  wire u3__abc_46775_n855;
  wire u3__abc_46775_n856;
  wire u3__abc_46775_n857;
  wire u3__abc_46775_n858;
  wire u3__abc_46775_n859;
  wire u3__abc_46775_n860;
  wire u3__abc_46775_n861;
  wire u3__abc_46775_n862;
  wire u3__abc_46775_n863;
  wire u3__abc_46775_n864;
  wire u3__abc_46775_n865;
  wire u3__abc_46775_n866;
  wire u3__abc_46775_n867;
  wire u3__abc_46775_n868;
  wire u3__abc_46775_n869;
  wire u3__abc_46775_n870;
  wire u3__abc_46775_n871;
  wire u3__abc_46775_n872;
  wire u3__abc_46775_n873;
  wire u3__abc_46775_n874;
  wire u3__abc_46775_n875;
  wire u3__abc_46775_n876;
  wire u3__abc_46775_n877;
  wire u3__abc_46775_n878;
  wire u3__abc_46775_n879;
  wire u3__abc_46775_n880;
  wire u3__abc_46775_n881;
  wire u3__abc_46775_n882;
  wire u3__abc_46775_n883;
  wire u3__abc_46775_n884;
  wire u3__abc_46775_n885;
  wire u3__abc_46775_n886;
  wire u3__abc_46775_n887;
  wire u3__abc_46775_n888;
  wire u3__abc_46775_n889;
  wire u3__abc_46775_n890;
  wire u3__abc_46775_n891;
  wire u3__abc_46775_n892;
  wire u3__abc_46775_n893;
  wire u3__abc_46775_n894;
  wire u3__abc_46775_n895;
  wire u3__abc_46775_n896;
  wire u3__abc_46775_n897;
  wire u3__abc_46775_n898;
  wire u3__abc_46775_n899;
  wire u3__abc_46775_n900;
  wire u3__abc_46775_n901;
  wire u3__abc_46775_n902;
  wire u3__abc_46775_n903;
  wire u3__abc_46775_n904;
  wire u3__abc_46775_n905;
  wire u3__abc_46775_n906;
  wire u3__abc_46775_n907;
  wire u3__abc_46775_n908;
  wire u3__abc_46775_n909;
  wire u3__abc_46775_n910;
  wire u3__abc_46775_n911;
  wire u3__abc_46775_n912;
  wire u3__abc_46775_n913;
  wire u3__abc_46775_n914;
  wire u3__abc_46775_n915;
  wire u3__abc_46775_n916;
  wire u3__abc_46775_n917;
  wire u3__abc_46775_n918;
  wire u3__abc_46775_n919;
  wire u3__abc_46775_n920;
  wire u3__abc_46775_n921;
  wire u3__abc_46775_n922;
  wire u3__abc_46775_n923;
  wire u3__abc_46775_n924;
  wire u3__abc_46775_n925;
  wire u3__abc_46775_n926;
  wire u3__abc_46775_n927;
  wire u3__abc_46775_n928;
  wire u3__abc_46775_n929;
  wire u3__abc_46775_n930;
  wire u3__abc_46775_n931;
  wire u3__abc_46775_n932;
  wire u3__abc_46775_n933;
  wire u3__abc_46775_n934;
  wire u3__abc_46775_n935;
  wire u3__abc_46775_n936;
  wire u3__abc_46775_n937;
  wire u3__abc_46775_n938;
  wire u3__abc_46775_n939;
  wire u3__abc_46775_n940;
  wire u3__abc_46775_n941;
  wire u3__abc_46775_n942;
  wire u3__abc_46775_n943;
  wire u3__abc_46775_n944;
  wire u3__abc_46775_n945;
  wire u3__abc_46775_n946;
  wire u3__abc_46775_n947;
  wire u3__abc_46775_n948;
  wire u3__abc_46775_n949;
  wire u3__abc_46775_n950;
  wire u3__abc_46775_n951;
  wire u3__abc_46775_n952;
  wire u3__abc_46775_n953;
  wire u3__abc_46775_n954;
  wire u3__abc_46775_n955;
  wire u3__abc_46775_n956;
  wire u3__abc_46775_n957;
  wire u3__abc_46775_n958;
  wire u3__abc_46775_n959;
  wire u3__abc_46775_n960;
  wire u3__abc_46775_n961;
  wire u3__abc_46775_n962;
  wire u3__abc_46775_n963;
  wire u3__abc_46775_n964;
  wire u3__abc_46775_n965;
  wire u3__abc_46775_n966;
  wire u3__abc_46775_n967;
  wire u3__abc_46775_n968;
  wire u3__abc_46775_n969;
  wire u3__abc_46775_n970;
  wire u3__abc_46775_n971;
  wire u3__abc_46775_n972;
  wire u3__abc_46775_n973;
  wire u3__abc_46775_n974;
  wire u3__abc_46775_n975;
  wire u3__abc_46775_n976;
  wire u3__abc_46775_n977;
  wire u3__abc_46775_n978;
  wire u3__abc_46775_n979;
  wire u3__abc_46775_n980;
  wire u3__abc_46775_n981;
  wire u3__abc_46775_n982;
  wire u3__abc_46775_n983;
  wire u3__abc_46775_n984;
  wire u3__abc_46775_n985;
  wire u3__abc_46775_n986;
  wire u3__abc_46775_n987;
  wire u3__abc_46775_n988;
  wire u3__abc_46775_n989;
  wire u3__abc_46775_n990;
  wire u3__abc_46775_n991;
  wire u3__abc_46775_n992;
  wire u3__abc_46775_n993;
  wire u3__abc_46775_n994;
  wire u3__abc_46775_n995;
  wire u3__abc_46775_n996;
  wire u3__abc_46775_n997;
  wire u3__abc_46775_n998;
  wire u3__abc_46775_n999;
  wire u3_byte0_0_;
  wire u3_byte0_0__FF_INPUT;
  wire u3_byte0_1_;
  wire u3_byte0_1__FF_INPUT;
  wire u3_byte0_2_;
  wire u3_byte0_2__FF_INPUT;
  wire u3_byte0_3_;
  wire u3_byte0_3__FF_INPUT;
  wire u3_byte0_4_;
  wire u3_byte0_4__FF_INPUT;
  wire u3_byte0_5_;
  wire u3_byte0_5__FF_INPUT;
  wire u3_byte0_6_;
  wire u3_byte0_6__FF_INPUT;
  wire u3_byte0_7_;
  wire u3_byte0_7__FF_INPUT;
  wire u3_byte1_0_;
  wire u3_byte1_0__FF_INPUT;
  wire u3_byte1_1_;
  wire u3_byte1_1__FF_INPUT;
  wire u3_byte1_2_;
  wire u3_byte1_2__FF_INPUT;
  wire u3_byte1_3_;
  wire u3_byte1_3__FF_INPUT;
  wire u3_byte1_4_;
  wire u3_byte1_4__FF_INPUT;
  wire u3_byte1_5_;
  wire u3_byte1_5__FF_INPUT;
  wire u3_byte1_6_;
  wire u3_byte1_6__FF_INPUT;
  wire u3_byte1_7_;
  wire u3_byte1_7__FF_INPUT;
  wire u3_byte2_0_;
  wire u3_byte2_0__FF_INPUT;
  wire u3_byte2_1_;
  wire u3_byte2_1__FF_INPUT;
  wire u3_byte2_2_;
  wire u3_byte2_2__FF_INPUT;
  wire u3_byte2_3_;
  wire u3_byte2_3__FF_INPUT;
  wire u3_byte2_4_;
  wire u3_byte2_4__FF_INPUT;
  wire u3_byte2_5_;
  wire u3_byte2_5__FF_INPUT;
  wire u3_byte2_6_;
  wire u3_byte2_6__FF_INPUT;
  wire u3_byte2_7_;
  wire u3_byte2_7__FF_INPUT;
  wire u3_mc_data_o_0__FF_INPUT;
  wire u3_mc_data_o_10__FF_INPUT;
  wire u3_mc_data_o_11__FF_INPUT;
  wire u3_mc_data_o_12__FF_INPUT;
  wire u3_mc_data_o_13__FF_INPUT;
  wire u3_mc_data_o_14__FF_INPUT;
  wire u3_mc_data_o_15__FF_INPUT;
  wire u3_mc_data_o_16__FF_INPUT;
  wire u3_mc_data_o_17__FF_INPUT;
  wire u3_mc_data_o_18__FF_INPUT;
  wire u3_mc_data_o_19__FF_INPUT;
  wire u3_mc_data_o_1__FF_INPUT;
  wire u3_mc_data_o_20__FF_INPUT;
  wire u3_mc_data_o_21__FF_INPUT;
  wire u3_mc_data_o_22__FF_INPUT;
  wire u3_mc_data_o_23__FF_INPUT;
  wire u3_mc_data_o_24__FF_INPUT;
  wire u3_mc_data_o_25__FF_INPUT;
  wire u3_mc_data_o_26__FF_INPUT;
  wire u3_mc_data_o_27__FF_INPUT;
  wire u3_mc_data_o_28__FF_INPUT;
  wire u3_mc_data_o_29__FF_INPUT;
  wire u3_mc_data_o_2__FF_INPUT;
  wire u3_mc_data_o_30__FF_INPUT;
  wire u3_mc_data_o_31__FF_INPUT;
  wire u3_mc_data_o_3__FF_INPUT;
  wire u3_mc_data_o_4__FF_INPUT;
  wire u3_mc_data_o_5__FF_INPUT;
  wire u3_mc_data_o_6__FF_INPUT;
  wire u3_mc_data_o_7__FF_INPUT;
  wire u3_mc_data_o_8__FF_INPUT;
  wire u3_mc_data_o_9__FF_INPUT;
  wire u3_mc_dp_o_0__FF_INPUT;
  wire u3_mc_dp_o_1__FF_INPUT;
  wire u3_mc_dp_o_2__FF_INPUT;
  wire u3_mc_dp_o_3__FF_INPUT;
  wire u3_pen;
  wire u3_rd_fifo_clr;
  wire u3_rd_fifo_out_0_;
  wire u3_rd_fifo_out_10_;
  wire u3_rd_fifo_out_11_;
  wire u3_rd_fifo_out_12_;
  wire u3_rd_fifo_out_13_;
  wire u3_rd_fifo_out_14_;
  wire u3_rd_fifo_out_15_;
  wire u3_rd_fifo_out_16_;
  wire u3_rd_fifo_out_17_;
  wire u3_rd_fifo_out_18_;
  wire u3_rd_fifo_out_19_;
  wire u3_rd_fifo_out_1_;
  wire u3_rd_fifo_out_20_;
  wire u3_rd_fifo_out_21_;
  wire u3_rd_fifo_out_22_;
  wire u3_rd_fifo_out_23_;
  wire u3_rd_fifo_out_24_;
  wire u3_rd_fifo_out_25_;
  wire u3_rd_fifo_out_26_;
  wire u3_rd_fifo_out_27_;
  wire u3_rd_fifo_out_28_;
  wire u3_rd_fifo_out_29_;
  wire u3_rd_fifo_out_2_;
  wire u3_rd_fifo_out_30_;
  wire u3_rd_fifo_out_31_;
  wire u3_rd_fifo_out_32_;
  wire u3_rd_fifo_out_33_;
  wire u3_rd_fifo_out_34_;
  wire u3_rd_fifo_out_35_;
  wire u3_rd_fifo_out_3_;
  wire u3_rd_fifo_out_4_;
  wire u3_rd_fifo_out_5_;
  wire u3_rd_fifo_out_6_;
  wire u3_rd_fifo_out_7_;
  wire u3_rd_fifo_out_8_;
  wire u3_rd_fifo_out_9_;
  wire u3_re;
  wire u3_u0__abc_48231_n1000;
  wire u3_u0__abc_48231_n1002;
  wire u3_u0__abc_48231_n1003;
  wire u3_u0__abc_48231_n1004;
  wire u3_u0__abc_48231_n1006;
  wire u3_u0__abc_48231_n1007;
  wire u3_u0__abc_48231_n1009;
  wire u3_u0__abc_48231_n1010;
  wire u3_u0__abc_48231_n1012;
  wire u3_u0__abc_48231_n1013;
  wire u3_u0__abc_48231_n1014;
  wire u3_u0__abc_48231_n1015;
  wire u3_u0__abc_48231_n1017;
  wire u3_u0__abc_48231_n1018;
  wire u3_u0__abc_48231_n1019;
  wire u3_u0__abc_48231_n1021;
  wire u3_u0__abc_48231_n1022;
  wire u3_u0__abc_48231_n1023;
  wire u3_u0__abc_48231_n1025;
  wire u3_u0__abc_48231_n1026;
  wire u3_u0__abc_48231_n1027;
  wire u3_u0__abc_48231_n1029;
  wire u3_u0__abc_48231_n1030;
  wire u3_u0__abc_48231_n1031;
  wire u3_u0__abc_48231_n1032;
  wire u3_u0__abc_48231_n1033;
  wire u3_u0__abc_48231_n1034;
  wire u3_u0__abc_48231_n1034_bF_buf0;
  wire u3_u0__abc_48231_n1034_bF_buf1;
  wire u3_u0__abc_48231_n1034_bF_buf2;
  wire u3_u0__abc_48231_n1034_bF_buf3;
  wire u3_u0__abc_48231_n1034_bF_buf4;
  wire u3_u0__abc_48231_n1034_bF_buf5;
  wire u3_u0__abc_48231_n1035;
  wire u3_u0__abc_48231_n1036;
  wire u3_u0__abc_48231_n1037;
  wire u3_u0__abc_48231_n1038;
  wire u3_u0__abc_48231_n1039;
  wire u3_u0__abc_48231_n1040;
  wire u3_u0__abc_48231_n1041;
  wire u3_u0__abc_48231_n1042;
  wire u3_u0__abc_48231_n1042_bF_buf0;
  wire u3_u0__abc_48231_n1042_bF_buf1;
  wire u3_u0__abc_48231_n1042_bF_buf2;
  wire u3_u0__abc_48231_n1042_bF_buf3;
  wire u3_u0__abc_48231_n1042_bF_buf4;
  wire u3_u0__abc_48231_n1042_bF_buf5;
  wire u3_u0__abc_48231_n1043;
  wire u3_u0__abc_48231_n1044;
  wire u3_u0__abc_48231_n1045;
  wire u3_u0__abc_48231_n1046;
  wire u3_u0__abc_48231_n1047;
  wire u3_u0__abc_48231_n1047_bF_buf0;
  wire u3_u0__abc_48231_n1047_bF_buf1;
  wire u3_u0__abc_48231_n1047_bF_buf2;
  wire u3_u0__abc_48231_n1047_bF_buf3;
  wire u3_u0__abc_48231_n1047_bF_buf4;
  wire u3_u0__abc_48231_n1047_bF_buf5;
  wire u3_u0__abc_48231_n1048;
  wire u3_u0__abc_48231_n1049;
  wire u3_u0__abc_48231_n1050;
  wire u3_u0__abc_48231_n1050_bF_buf0;
  wire u3_u0__abc_48231_n1050_bF_buf1;
  wire u3_u0__abc_48231_n1050_bF_buf2;
  wire u3_u0__abc_48231_n1050_bF_buf3;
  wire u3_u0__abc_48231_n1050_bF_buf4;
  wire u3_u0__abc_48231_n1050_bF_buf5;
  wire u3_u0__abc_48231_n1051;
  wire u3_u0__abc_48231_n1052;
  wire u3_u0__abc_48231_n1053;
  wire u3_u0__abc_48231_n1054;
  wire u3_u0__abc_48231_n1056;
  wire u3_u0__abc_48231_n1057;
  wire u3_u0__abc_48231_n1058;
  wire u3_u0__abc_48231_n1059;
  wire u3_u0__abc_48231_n1060;
  wire u3_u0__abc_48231_n1061;
  wire u3_u0__abc_48231_n1063;
  wire u3_u0__abc_48231_n1064;
  wire u3_u0__abc_48231_n1065;
  wire u3_u0__abc_48231_n1066;
  wire u3_u0__abc_48231_n1067;
  wire u3_u0__abc_48231_n1068;
  wire u3_u0__abc_48231_n1070;
  wire u3_u0__abc_48231_n1071;
  wire u3_u0__abc_48231_n1072;
  wire u3_u0__abc_48231_n1073;
  wire u3_u0__abc_48231_n1074;
  wire u3_u0__abc_48231_n1075;
  wire u3_u0__abc_48231_n1077;
  wire u3_u0__abc_48231_n1078;
  wire u3_u0__abc_48231_n1079;
  wire u3_u0__abc_48231_n1080;
  wire u3_u0__abc_48231_n1081;
  wire u3_u0__abc_48231_n1082;
  wire u3_u0__abc_48231_n1084;
  wire u3_u0__abc_48231_n1085;
  wire u3_u0__abc_48231_n1086;
  wire u3_u0__abc_48231_n1087;
  wire u3_u0__abc_48231_n1088;
  wire u3_u0__abc_48231_n1089;
  wire u3_u0__abc_48231_n1091;
  wire u3_u0__abc_48231_n1092;
  wire u3_u0__abc_48231_n1093;
  wire u3_u0__abc_48231_n1094;
  wire u3_u0__abc_48231_n1095;
  wire u3_u0__abc_48231_n1096;
  wire u3_u0__abc_48231_n1098;
  wire u3_u0__abc_48231_n1099;
  wire u3_u0__abc_48231_n1100;
  wire u3_u0__abc_48231_n1101;
  wire u3_u0__abc_48231_n1102;
  wire u3_u0__abc_48231_n1103;
  wire u3_u0__abc_48231_n1105;
  wire u3_u0__abc_48231_n1106;
  wire u3_u0__abc_48231_n1107;
  wire u3_u0__abc_48231_n1108;
  wire u3_u0__abc_48231_n1109;
  wire u3_u0__abc_48231_n1110;
  wire u3_u0__abc_48231_n1112;
  wire u3_u0__abc_48231_n1113;
  wire u3_u0__abc_48231_n1114;
  wire u3_u0__abc_48231_n1115;
  wire u3_u0__abc_48231_n1116;
  wire u3_u0__abc_48231_n1117;
  wire u3_u0__abc_48231_n1119;
  wire u3_u0__abc_48231_n1120;
  wire u3_u0__abc_48231_n1121;
  wire u3_u0__abc_48231_n1122;
  wire u3_u0__abc_48231_n1123;
  wire u3_u0__abc_48231_n1124;
  wire u3_u0__abc_48231_n1126;
  wire u3_u0__abc_48231_n1127;
  wire u3_u0__abc_48231_n1128;
  wire u3_u0__abc_48231_n1129;
  wire u3_u0__abc_48231_n1130;
  wire u3_u0__abc_48231_n1131;
  wire u3_u0__abc_48231_n1133;
  wire u3_u0__abc_48231_n1134;
  wire u3_u0__abc_48231_n1135;
  wire u3_u0__abc_48231_n1136;
  wire u3_u0__abc_48231_n1137;
  wire u3_u0__abc_48231_n1138;
  wire u3_u0__abc_48231_n1140;
  wire u3_u0__abc_48231_n1141;
  wire u3_u0__abc_48231_n1142;
  wire u3_u0__abc_48231_n1143;
  wire u3_u0__abc_48231_n1144;
  wire u3_u0__abc_48231_n1145;
  wire u3_u0__abc_48231_n1147;
  wire u3_u0__abc_48231_n1148;
  wire u3_u0__abc_48231_n1149;
  wire u3_u0__abc_48231_n1150;
  wire u3_u0__abc_48231_n1151;
  wire u3_u0__abc_48231_n1152;
  wire u3_u0__abc_48231_n1154;
  wire u3_u0__abc_48231_n1155;
  wire u3_u0__abc_48231_n1156;
  wire u3_u0__abc_48231_n1157;
  wire u3_u0__abc_48231_n1158;
  wire u3_u0__abc_48231_n1159;
  wire u3_u0__abc_48231_n1161;
  wire u3_u0__abc_48231_n1162;
  wire u3_u0__abc_48231_n1163;
  wire u3_u0__abc_48231_n1164;
  wire u3_u0__abc_48231_n1165;
  wire u3_u0__abc_48231_n1166;
  wire u3_u0__abc_48231_n1168;
  wire u3_u0__abc_48231_n1169;
  wire u3_u0__abc_48231_n1170;
  wire u3_u0__abc_48231_n1171;
  wire u3_u0__abc_48231_n1172;
  wire u3_u0__abc_48231_n1173;
  wire u3_u0__abc_48231_n1175;
  wire u3_u0__abc_48231_n1176;
  wire u3_u0__abc_48231_n1177;
  wire u3_u0__abc_48231_n1178;
  wire u3_u0__abc_48231_n1179;
  wire u3_u0__abc_48231_n1180;
  wire u3_u0__abc_48231_n1182;
  wire u3_u0__abc_48231_n1183;
  wire u3_u0__abc_48231_n1184;
  wire u3_u0__abc_48231_n1185;
  wire u3_u0__abc_48231_n1186;
  wire u3_u0__abc_48231_n1187;
  wire u3_u0__abc_48231_n1189;
  wire u3_u0__abc_48231_n1190;
  wire u3_u0__abc_48231_n1191;
  wire u3_u0__abc_48231_n1192;
  wire u3_u0__abc_48231_n1193;
  wire u3_u0__abc_48231_n1194;
  wire u3_u0__abc_48231_n1196;
  wire u3_u0__abc_48231_n1197;
  wire u3_u0__abc_48231_n1198;
  wire u3_u0__abc_48231_n1199;
  wire u3_u0__abc_48231_n1200;
  wire u3_u0__abc_48231_n1201;
  wire u3_u0__abc_48231_n1203;
  wire u3_u0__abc_48231_n1204;
  wire u3_u0__abc_48231_n1205;
  wire u3_u0__abc_48231_n1206;
  wire u3_u0__abc_48231_n1207;
  wire u3_u0__abc_48231_n1208;
  wire u3_u0__abc_48231_n1210;
  wire u3_u0__abc_48231_n1211;
  wire u3_u0__abc_48231_n1212;
  wire u3_u0__abc_48231_n1213;
  wire u3_u0__abc_48231_n1214;
  wire u3_u0__abc_48231_n1215;
  wire u3_u0__abc_48231_n1217;
  wire u3_u0__abc_48231_n1218;
  wire u3_u0__abc_48231_n1219;
  wire u3_u0__abc_48231_n1220;
  wire u3_u0__abc_48231_n1221;
  wire u3_u0__abc_48231_n1222;
  wire u3_u0__abc_48231_n1224;
  wire u3_u0__abc_48231_n1225;
  wire u3_u0__abc_48231_n1226;
  wire u3_u0__abc_48231_n1227;
  wire u3_u0__abc_48231_n1228;
  wire u3_u0__abc_48231_n1229;
  wire u3_u0__abc_48231_n1231;
  wire u3_u0__abc_48231_n1232;
  wire u3_u0__abc_48231_n1233;
  wire u3_u0__abc_48231_n1234;
  wire u3_u0__abc_48231_n1235;
  wire u3_u0__abc_48231_n1236;
  wire u3_u0__abc_48231_n1238;
  wire u3_u0__abc_48231_n1239;
  wire u3_u0__abc_48231_n1240;
  wire u3_u0__abc_48231_n1241;
  wire u3_u0__abc_48231_n1242;
  wire u3_u0__abc_48231_n1243;
  wire u3_u0__abc_48231_n1245;
  wire u3_u0__abc_48231_n1246;
  wire u3_u0__abc_48231_n1247;
  wire u3_u0__abc_48231_n1248;
  wire u3_u0__abc_48231_n1249;
  wire u3_u0__abc_48231_n1250;
  wire u3_u0__abc_48231_n1252;
  wire u3_u0__abc_48231_n1253;
  wire u3_u0__abc_48231_n1254;
  wire u3_u0__abc_48231_n1255;
  wire u3_u0__abc_48231_n1256;
  wire u3_u0__abc_48231_n1257;
  wire u3_u0__abc_48231_n1259;
  wire u3_u0__abc_48231_n1260;
  wire u3_u0__abc_48231_n1261;
  wire u3_u0__abc_48231_n1262;
  wire u3_u0__abc_48231_n1263;
  wire u3_u0__abc_48231_n1264;
  wire u3_u0__abc_48231_n1266;
  wire u3_u0__abc_48231_n1267;
  wire u3_u0__abc_48231_n1268;
  wire u3_u0__abc_48231_n1269;
  wire u3_u0__abc_48231_n1270;
  wire u3_u0__abc_48231_n1271;
  wire u3_u0__abc_48231_n1273;
  wire u3_u0__abc_48231_n1274;
  wire u3_u0__abc_48231_n1275;
  wire u3_u0__abc_48231_n1276;
  wire u3_u0__abc_48231_n1277;
  wire u3_u0__abc_48231_n1278;
  wire u3_u0__abc_48231_n1280;
  wire u3_u0__abc_48231_n1281;
  wire u3_u0__abc_48231_n1282;
  wire u3_u0__abc_48231_n1283;
  wire u3_u0__abc_48231_n1284;
  wire u3_u0__abc_48231_n1285;
  wire u3_u0__abc_48231_n1287;
  wire u3_u0__abc_48231_n1288;
  wire u3_u0__abc_48231_n1289;
  wire u3_u0__abc_48231_n1290;
  wire u3_u0__abc_48231_n1291;
  wire u3_u0__abc_48231_n1292;
  wire u3_u0__abc_48231_n1294;
  wire u3_u0__abc_48231_n1295;
  wire u3_u0__abc_48231_n1296;
  wire u3_u0__abc_48231_n1297;
  wire u3_u0__abc_48231_n1298;
  wire u3_u0__abc_48231_n1299;
  wire u3_u0__abc_48231_n382;
  wire u3_u0__abc_48231_n382_bF_buf0;
  wire u3_u0__abc_48231_n382_bF_buf1;
  wire u3_u0__abc_48231_n382_bF_buf2;
  wire u3_u0__abc_48231_n382_bF_buf3;
  wire u3_u0__abc_48231_n382_bF_buf4;
  wire u3_u0__abc_48231_n382_bF_buf5;
  wire u3_u0__abc_48231_n382_bF_buf6;
  wire u3_u0__abc_48231_n382_bF_buf7;
  wire u3_u0__abc_48231_n383;
  wire u3_u0__abc_48231_n384_1;
  wire u3_u0__abc_48231_n385;
  wire u3_u0__abc_48231_n386;
  wire u3_u0__abc_48231_n388_1;
  wire u3_u0__abc_48231_n389;
  wire u3_u0__abc_48231_n390;
  wire u3_u0__abc_48231_n391;
  wire u3_u0__abc_48231_n393;
  wire u3_u0__abc_48231_n394;
  wire u3_u0__abc_48231_n395;
  wire u3_u0__abc_48231_n396_1;
  wire u3_u0__abc_48231_n398;
  wire u3_u0__abc_48231_n399;
  wire u3_u0__abc_48231_n400_1;
  wire u3_u0__abc_48231_n401;
  wire u3_u0__abc_48231_n403;
  wire u3_u0__abc_48231_n404_1;
  wire u3_u0__abc_48231_n405;
  wire u3_u0__abc_48231_n406;
  wire u3_u0__abc_48231_n408_1;
  wire u3_u0__abc_48231_n409;
  wire u3_u0__abc_48231_n410;
  wire u3_u0__abc_48231_n411;
  wire u3_u0__abc_48231_n413;
  wire u3_u0__abc_48231_n414;
  wire u3_u0__abc_48231_n415;
  wire u3_u0__abc_48231_n416_1;
  wire u3_u0__abc_48231_n418;
  wire u3_u0__abc_48231_n419;
  wire u3_u0__abc_48231_n420_1;
  wire u3_u0__abc_48231_n421;
  wire u3_u0__abc_48231_n423;
  wire u3_u0__abc_48231_n424_1;
  wire u3_u0__abc_48231_n425;
  wire u3_u0__abc_48231_n426;
  wire u3_u0__abc_48231_n428_1;
  wire u3_u0__abc_48231_n429;
  wire u3_u0__abc_48231_n430;
  wire u3_u0__abc_48231_n431;
  wire u3_u0__abc_48231_n433;
  wire u3_u0__abc_48231_n434;
  wire u3_u0__abc_48231_n435;
  wire u3_u0__abc_48231_n436_1;
  wire u3_u0__abc_48231_n438;
  wire u3_u0__abc_48231_n439;
  wire u3_u0__abc_48231_n440_1;
  wire u3_u0__abc_48231_n441;
  wire u3_u0__abc_48231_n443;
  wire u3_u0__abc_48231_n444_1;
  wire u3_u0__abc_48231_n445;
  wire u3_u0__abc_48231_n446;
  wire u3_u0__abc_48231_n448_1;
  wire u3_u0__abc_48231_n449;
  wire u3_u0__abc_48231_n450;
  wire u3_u0__abc_48231_n451;
  wire u3_u0__abc_48231_n453;
  wire u3_u0__abc_48231_n454;
  wire u3_u0__abc_48231_n455;
  wire u3_u0__abc_48231_n456_1;
  wire u3_u0__abc_48231_n458;
  wire u3_u0__abc_48231_n459;
  wire u3_u0__abc_48231_n460_1;
  wire u3_u0__abc_48231_n461;
  wire u3_u0__abc_48231_n463;
  wire u3_u0__abc_48231_n464_1;
  wire u3_u0__abc_48231_n465;
  wire u3_u0__abc_48231_n466;
  wire u3_u0__abc_48231_n468_1;
  wire u3_u0__abc_48231_n469;
  wire u3_u0__abc_48231_n470;
  wire u3_u0__abc_48231_n471;
  wire u3_u0__abc_48231_n473;
  wire u3_u0__abc_48231_n474;
  wire u3_u0__abc_48231_n475;
  wire u3_u0__abc_48231_n476_1;
  wire u3_u0__abc_48231_n478;
  wire u3_u0__abc_48231_n479;
  wire u3_u0__abc_48231_n480_1;
  wire u3_u0__abc_48231_n481;
  wire u3_u0__abc_48231_n483;
  wire u3_u0__abc_48231_n484_1;
  wire u3_u0__abc_48231_n485;
  wire u3_u0__abc_48231_n486;
  wire u3_u0__abc_48231_n488_1;
  wire u3_u0__abc_48231_n489;
  wire u3_u0__abc_48231_n490;
  wire u3_u0__abc_48231_n491;
  wire u3_u0__abc_48231_n493;
  wire u3_u0__abc_48231_n494;
  wire u3_u0__abc_48231_n495;
  wire u3_u0__abc_48231_n496_1;
  wire u3_u0__abc_48231_n498;
  wire u3_u0__abc_48231_n499;
  wire u3_u0__abc_48231_n500_1;
  wire u3_u0__abc_48231_n501;
  wire u3_u0__abc_48231_n503;
  wire u3_u0__abc_48231_n504_1;
  wire u3_u0__abc_48231_n505;
  wire u3_u0__abc_48231_n506;
  wire u3_u0__abc_48231_n508_1;
  wire u3_u0__abc_48231_n509;
  wire u3_u0__abc_48231_n510;
  wire u3_u0__abc_48231_n511;
  wire u3_u0__abc_48231_n513_1;
  wire u3_u0__abc_48231_n514;
  wire u3_u0__abc_48231_n514_1;
  wire u3_u0__abc_48231_n515;
  wire u3_u0__abc_48231_n516;
  wire u3_u0__abc_48231_n518;
  wire u3_u0__abc_48231_n519;
  wire u3_u0__abc_48231_n520;
  wire u3_u0__abc_48231_n521;
  wire u3_u0__abc_48231_n523;
  wire u3_u0__abc_48231_n524;
  wire u3_u0__abc_48231_n525;
  wire u3_u0__abc_48231_n526;
  wire u3_u0__abc_48231_n528;
  wire u3_u0__abc_48231_n529;
  wire u3_u0__abc_48231_n530;
  wire u3_u0__abc_48231_n531;
  wire u3_u0__abc_48231_n533;
  wire u3_u0__abc_48231_n534;
  wire u3_u0__abc_48231_n535;
  wire u3_u0__abc_48231_n536;
  wire u3_u0__abc_48231_n538;
  wire u3_u0__abc_48231_n539;
  wire u3_u0__abc_48231_n540;
  wire u3_u0__abc_48231_n541;
  wire u3_u0__abc_48231_n543;
  wire u3_u0__abc_48231_n544;
  wire u3_u0__abc_48231_n545;
  wire u3_u0__abc_48231_n546;
  wire u3_u0__abc_48231_n548;
  wire u3_u0__abc_48231_n549;
  wire u3_u0__abc_48231_n550;
  wire u3_u0__abc_48231_n551;
  wire u3_u0__abc_48231_n553;
  wire u3_u0__abc_48231_n554;
  wire u3_u0__abc_48231_n555;
  wire u3_u0__abc_48231_n556;
  wire u3_u0__abc_48231_n558;
  wire u3_u0__abc_48231_n559;
  wire u3_u0__abc_48231_n560;
  wire u3_u0__abc_48231_n561;
  wire u3_u0__abc_48231_n563;
  wire u3_u0__abc_48231_n563_bF_buf0;
  wire u3_u0__abc_48231_n563_bF_buf1;
  wire u3_u0__abc_48231_n563_bF_buf2;
  wire u3_u0__abc_48231_n563_bF_buf3;
  wire u3_u0__abc_48231_n563_bF_buf4;
  wire u3_u0__abc_48231_n563_bF_buf5;
  wire u3_u0__abc_48231_n563_bF_buf6;
  wire u3_u0__abc_48231_n563_bF_buf7;
  wire u3_u0__abc_48231_n564;
  wire u3_u0__abc_48231_n565;
  wire u3_u0__abc_48231_n566;
  wire u3_u0__abc_48231_n568;
  wire u3_u0__abc_48231_n569;
  wire u3_u0__abc_48231_n570;
  wire u3_u0__abc_48231_n572;
  wire u3_u0__abc_48231_n573;
  wire u3_u0__abc_48231_n574;
  wire u3_u0__abc_48231_n576;
  wire u3_u0__abc_48231_n577;
  wire u3_u0__abc_48231_n578;
  wire u3_u0__abc_48231_n580;
  wire u3_u0__abc_48231_n581;
  wire u3_u0__abc_48231_n582;
  wire u3_u0__abc_48231_n584;
  wire u3_u0__abc_48231_n585;
  wire u3_u0__abc_48231_n586;
  wire u3_u0__abc_48231_n588;
  wire u3_u0__abc_48231_n589;
  wire u3_u0__abc_48231_n590;
  wire u3_u0__abc_48231_n592;
  wire u3_u0__abc_48231_n593;
  wire u3_u0__abc_48231_n594;
  wire u3_u0__abc_48231_n596;
  wire u3_u0__abc_48231_n597;
  wire u3_u0__abc_48231_n598;
  wire u3_u0__abc_48231_n600;
  wire u3_u0__abc_48231_n601;
  wire u3_u0__abc_48231_n602;
  wire u3_u0__abc_48231_n604;
  wire u3_u0__abc_48231_n605;
  wire u3_u0__abc_48231_n606;
  wire u3_u0__abc_48231_n608;
  wire u3_u0__abc_48231_n609;
  wire u3_u0__abc_48231_n610;
  wire u3_u0__abc_48231_n612;
  wire u3_u0__abc_48231_n613;
  wire u3_u0__abc_48231_n614;
  wire u3_u0__abc_48231_n616;
  wire u3_u0__abc_48231_n617;
  wire u3_u0__abc_48231_n618;
  wire u3_u0__abc_48231_n620;
  wire u3_u0__abc_48231_n621;
  wire u3_u0__abc_48231_n622;
  wire u3_u0__abc_48231_n624;
  wire u3_u0__abc_48231_n625;
  wire u3_u0__abc_48231_n626;
  wire u3_u0__abc_48231_n628;
  wire u3_u0__abc_48231_n629;
  wire u3_u0__abc_48231_n630;
  wire u3_u0__abc_48231_n632;
  wire u3_u0__abc_48231_n633;
  wire u3_u0__abc_48231_n634;
  wire u3_u0__abc_48231_n636;
  wire u3_u0__abc_48231_n637;
  wire u3_u0__abc_48231_n638;
  wire u3_u0__abc_48231_n640;
  wire u3_u0__abc_48231_n641;
  wire u3_u0__abc_48231_n642;
  wire u3_u0__abc_48231_n644;
  wire u3_u0__abc_48231_n645;
  wire u3_u0__abc_48231_n646;
  wire u3_u0__abc_48231_n648;
  wire u3_u0__abc_48231_n649;
  wire u3_u0__abc_48231_n650;
  wire u3_u0__abc_48231_n652;
  wire u3_u0__abc_48231_n653;
  wire u3_u0__abc_48231_n654;
  wire u3_u0__abc_48231_n656;
  wire u3_u0__abc_48231_n657;
  wire u3_u0__abc_48231_n658;
  wire u3_u0__abc_48231_n660;
  wire u3_u0__abc_48231_n661;
  wire u3_u0__abc_48231_n662;
  wire u3_u0__abc_48231_n664;
  wire u3_u0__abc_48231_n665;
  wire u3_u0__abc_48231_n666;
  wire u3_u0__abc_48231_n668;
  wire u3_u0__abc_48231_n669;
  wire u3_u0__abc_48231_n670;
  wire u3_u0__abc_48231_n672;
  wire u3_u0__abc_48231_n673;
  wire u3_u0__abc_48231_n674;
  wire u3_u0__abc_48231_n676;
  wire u3_u0__abc_48231_n677;
  wire u3_u0__abc_48231_n678;
  wire u3_u0__abc_48231_n680;
  wire u3_u0__abc_48231_n681;
  wire u3_u0__abc_48231_n682;
  wire u3_u0__abc_48231_n684;
  wire u3_u0__abc_48231_n685;
  wire u3_u0__abc_48231_n686;
  wire u3_u0__abc_48231_n688;
  wire u3_u0__abc_48231_n689;
  wire u3_u0__abc_48231_n690;
  wire u3_u0__abc_48231_n692;
  wire u3_u0__abc_48231_n693;
  wire u3_u0__abc_48231_n694;
  wire u3_u0__abc_48231_n696;
  wire u3_u0__abc_48231_n697;
  wire u3_u0__abc_48231_n698;
  wire u3_u0__abc_48231_n700;
  wire u3_u0__abc_48231_n701;
  wire u3_u0__abc_48231_n702;
  wire u3_u0__abc_48231_n704;
  wire u3_u0__abc_48231_n705;
  wire u3_u0__abc_48231_n706;
  wire u3_u0__abc_48231_n708;
  wire u3_u0__abc_48231_n708_bF_buf0;
  wire u3_u0__abc_48231_n708_bF_buf1;
  wire u3_u0__abc_48231_n708_bF_buf2;
  wire u3_u0__abc_48231_n708_bF_buf3;
  wire u3_u0__abc_48231_n708_bF_buf4;
  wire u3_u0__abc_48231_n708_bF_buf5;
  wire u3_u0__abc_48231_n708_bF_buf6;
  wire u3_u0__abc_48231_n708_bF_buf7;
  wire u3_u0__abc_48231_n709;
  wire u3_u0__abc_48231_n710;
  wire u3_u0__abc_48231_n711;
  wire u3_u0__abc_48231_n713;
  wire u3_u0__abc_48231_n714;
  wire u3_u0__abc_48231_n715;
  wire u3_u0__abc_48231_n717;
  wire u3_u0__abc_48231_n718;
  wire u3_u0__abc_48231_n719;
  wire u3_u0__abc_48231_n721;
  wire u3_u0__abc_48231_n722;
  wire u3_u0__abc_48231_n723;
  wire u3_u0__abc_48231_n725;
  wire u3_u0__abc_48231_n726;
  wire u3_u0__abc_48231_n727;
  wire u3_u0__abc_48231_n729;
  wire u3_u0__abc_48231_n730;
  wire u3_u0__abc_48231_n731;
  wire u3_u0__abc_48231_n733;
  wire u3_u0__abc_48231_n734;
  wire u3_u0__abc_48231_n735;
  wire u3_u0__abc_48231_n737;
  wire u3_u0__abc_48231_n738;
  wire u3_u0__abc_48231_n739;
  wire u3_u0__abc_48231_n741;
  wire u3_u0__abc_48231_n742;
  wire u3_u0__abc_48231_n743;
  wire u3_u0__abc_48231_n745;
  wire u3_u0__abc_48231_n746;
  wire u3_u0__abc_48231_n747;
  wire u3_u0__abc_48231_n749;
  wire u3_u0__abc_48231_n750;
  wire u3_u0__abc_48231_n751;
  wire u3_u0__abc_48231_n753;
  wire u3_u0__abc_48231_n754;
  wire u3_u0__abc_48231_n755;
  wire u3_u0__abc_48231_n757;
  wire u3_u0__abc_48231_n758;
  wire u3_u0__abc_48231_n759;
  wire u3_u0__abc_48231_n761;
  wire u3_u0__abc_48231_n762;
  wire u3_u0__abc_48231_n763;
  wire u3_u0__abc_48231_n765;
  wire u3_u0__abc_48231_n766;
  wire u3_u0__abc_48231_n767;
  wire u3_u0__abc_48231_n769;
  wire u3_u0__abc_48231_n770;
  wire u3_u0__abc_48231_n771;
  wire u3_u0__abc_48231_n773;
  wire u3_u0__abc_48231_n774;
  wire u3_u0__abc_48231_n775;
  wire u3_u0__abc_48231_n777;
  wire u3_u0__abc_48231_n778;
  wire u3_u0__abc_48231_n779;
  wire u3_u0__abc_48231_n781;
  wire u3_u0__abc_48231_n782;
  wire u3_u0__abc_48231_n783;
  wire u3_u0__abc_48231_n785;
  wire u3_u0__abc_48231_n786;
  wire u3_u0__abc_48231_n787;
  wire u3_u0__abc_48231_n789;
  wire u3_u0__abc_48231_n790;
  wire u3_u0__abc_48231_n791;
  wire u3_u0__abc_48231_n793;
  wire u3_u0__abc_48231_n794;
  wire u3_u0__abc_48231_n795;
  wire u3_u0__abc_48231_n797;
  wire u3_u0__abc_48231_n798;
  wire u3_u0__abc_48231_n799;
  wire u3_u0__abc_48231_n801;
  wire u3_u0__abc_48231_n802;
  wire u3_u0__abc_48231_n803;
  wire u3_u0__abc_48231_n805;
  wire u3_u0__abc_48231_n806;
  wire u3_u0__abc_48231_n807;
  wire u3_u0__abc_48231_n809;
  wire u3_u0__abc_48231_n810;
  wire u3_u0__abc_48231_n811;
  wire u3_u0__abc_48231_n813;
  wire u3_u0__abc_48231_n814;
  wire u3_u0__abc_48231_n815;
  wire u3_u0__abc_48231_n817;
  wire u3_u0__abc_48231_n818;
  wire u3_u0__abc_48231_n819;
  wire u3_u0__abc_48231_n821;
  wire u3_u0__abc_48231_n822;
  wire u3_u0__abc_48231_n823;
  wire u3_u0__abc_48231_n825;
  wire u3_u0__abc_48231_n826;
  wire u3_u0__abc_48231_n827;
  wire u3_u0__abc_48231_n829;
  wire u3_u0__abc_48231_n830;
  wire u3_u0__abc_48231_n831;
  wire u3_u0__abc_48231_n833;
  wire u3_u0__abc_48231_n834;
  wire u3_u0__abc_48231_n835;
  wire u3_u0__abc_48231_n837;
  wire u3_u0__abc_48231_n838;
  wire u3_u0__abc_48231_n839;
  wire u3_u0__abc_48231_n841;
  wire u3_u0__abc_48231_n842;
  wire u3_u0__abc_48231_n843;
  wire u3_u0__abc_48231_n845;
  wire u3_u0__abc_48231_n846;
  wire u3_u0__abc_48231_n847;
  wire u3_u0__abc_48231_n849;
  wire u3_u0__abc_48231_n850;
  wire u3_u0__abc_48231_n851;
  wire u3_u0__abc_48231_n853;
  wire u3_u0__abc_48231_n853_bF_buf0;
  wire u3_u0__abc_48231_n853_bF_buf1;
  wire u3_u0__abc_48231_n853_bF_buf2;
  wire u3_u0__abc_48231_n853_bF_buf3;
  wire u3_u0__abc_48231_n853_bF_buf4;
  wire u3_u0__abc_48231_n853_bF_buf5;
  wire u3_u0__abc_48231_n853_bF_buf6;
  wire u3_u0__abc_48231_n853_bF_buf7;
  wire u3_u0__abc_48231_n854;
  wire u3_u0__abc_48231_n855;
  wire u3_u0__abc_48231_n856;
  wire u3_u0__abc_48231_n858;
  wire u3_u0__abc_48231_n859;
  wire u3_u0__abc_48231_n860;
  wire u3_u0__abc_48231_n862;
  wire u3_u0__abc_48231_n863;
  wire u3_u0__abc_48231_n864;
  wire u3_u0__abc_48231_n866;
  wire u3_u0__abc_48231_n867;
  wire u3_u0__abc_48231_n868;
  wire u3_u0__abc_48231_n870;
  wire u3_u0__abc_48231_n871;
  wire u3_u0__abc_48231_n872;
  wire u3_u0__abc_48231_n874;
  wire u3_u0__abc_48231_n875;
  wire u3_u0__abc_48231_n876;
  wire u3_u0__abc_48231_n878;
  wire u3_u0__abc_48231_n879;
  wire u3_u0__abc_48231_n880;
  wire u3_u0__abc_48231_n882;
  wire u3_u0__abc_48231_n883;
  wire u3_u0__abc_48231_n884;
  wire u3_u0__abc_48231_n886;
  wire u3_u0__abc_48231_n887;
  wire u3_u0__abc_48231_n888;
  wire u3_u0__abc_48231_n890;
  wire u3_u0__abc_48231_n891;
  wire u3_u0__abc_48231_n892;
  wire u3_u0__abc_48231_n894;
  wire u3_u0__abc_48231_n895;
  wire u3_u0__abc_48231_n896;
  wire u3_u0__abc_48231_n898;
  wire u3_u0__abc_48231_n899;
  wire u3_u0__abc_48231_n900;
  wire u3_u0__abc_48231_n902;
  wire u3_u0__abc_48231_n903;
  wire u3_u0__abc_48231_n904;
  wire u3_u0__abc_48231_n906;
  wire u3_u0__abc_48231_n907;
  wire u3_u0__abc_48231_n908;
  wire u3_u0__abc_48231_n910;
  wire u3_u0__abc_48231_n911;
  wire u3_u0__abc_48231_n912;
  wire u3_u0__abc_48231_n914;
  wire u3_u0__abc_48231_n915;
  wire u3_u0__abc_48231_n916;
  wire u3_u0__abc_48231_n918;
  wire u3_u0__abc_48231_n919;
  wire u3_u0__abc_48231_n920;
  wire u3_u0__abc_48231_n922;
  wire u3_u0__abc_48231_n923;
  wire u3_u0__abc_48231_n924;
  wire u3_u0__abc_48231_n926;
  wire u3_u0__abc_48231_n927;
  wire u3_u0__abc_48231_n928;
  wire u3_u0__abc_48231_n930;
  wire u3_u0__abc_48231_n931;
  wire u3_u0__abc_48231_n932;
  wire u3_u0__abc_48231_n934;
  wire u3_u0__abc_48231_n935;
  wire u3_u0__abc_48231_n936;
  wire u3_u0__abc_48231_n938;
  wire u3_u0__abc_48231_n939;
  wire u3_u0__abc_48231_n940;
  wire u3_u0__abc_48231_n942;
  wire u3_u0__abc_48231_n943;
  wire u3_u0__abc_48231_n944;
  wire u3_u0__abc_48231_n946;
  wire u3_u0__abc_48231_n947;
  wire u3_u0__abc_48231_n948;
  wire u3_u0__abc_48231_n950;
  wire u3_u0__abc_48231_n951;
  wire u3_u0__abc_48231_n952;
  wire u3_u0__abc_48231_n954;
  wire u3_u0__abc_48231_n955;
  wire u3_u0__abc_48231_n956;
  wire u3_u0__abc_48231_n958;
  wire u3_u0__abc_48231_n959;
  wire u3_u0__abc_48231_n960;
  wire u3_u0__abc_48231_n962;
  wire u3_u0__abc_48231_n963;
  wire u3_u0__abc_48231_n964;
  wire u3_u0__abc_48231_n966;
  wire u3_u0__abc_48231_n967;
  wire u3_u0__abc_48231_n968;
  wire u3_u0__abc_48231_n970;
  wire u3_u0__abc_48231_n971;
  wire u3_u0__abc_48231_n972;
  wire u3_u0__abc_48231_n974;
  wire u3_u0__abc_48231_n975;
  wire u3_u0__abc_48231_n976;
  wire u3_u0__abc_48231_n978;
  wire u3_u0__abc_48231_n979;
  wire u3_u0__abc_48231_n980;
  wire u3_u0__abc_48231_n982;
  wire u3_u0__abc_48231_n983;
  wire u3_u0__abc_48231_n984;
  wire u3_u0__abc_48231_n986;
  wire u3_u0__abc_48231_n987;
  wire u3_u0__abc_48231_n988;
  wire u3_u0__abc_48231_n990;
  wire u3_u0__abc_48231_n991;
  wire u3_u0__abc_48231_n992;
  wire u3_u0__abc_48231_n994;
  wire u3_u0__abc_48231_n995;
  wire u3_u0__abc_48231_n996;
  wire u3_u0__abc_48231_n998;
  wire u3_u0__abc_48231_n999;
  wire u3_u0_r0_0_;
  wire u3_u0_r0_0__FF_INPUT;
  wire u3_u0_r0_10_;
  wire u3_u0_r0_10__FF_INPUT;
  wire u3_u0_r0_11_;
  wire u3_u0_r0_11__FF_INPUT;
  wire u3_u0_r0_12_;
  wire u3_u0_r0_12__FF_INPUT;
  wire u3_u0_r0_13_;
  wire u3_u0_r0_13__FF_INPUT;
  wire u3_u0_r0_14_;
  wire u3_u0_r0_14__FF_INPUT;
  wire u3_u0_r0_15_;
  wire u3_u0_r0_15__FF_INPUT;
  wire u3_u0_r0_16_;
  wire u3_u0_r0_16__FF_INPUT;
  wire u3_u0_r0_17_;
  wire u3_u0_r0_17__FF_INPUT;
  wire u3_u0_r0_18_;
  wire u3_u0_r0_18__FF_INPUT;
  wire u3_u0_r0_19_;
  wire u3_u0_r0_19__FF_INPUT;
  wire u3_u0_r0_1_;
  wire u3_u0_r0_1__FF_INPUT;
  wire u3_u0_r0_20_;
  wire u3_u0_r0_20__FF_INPUT;
  wire u3_u0_r0_21_;
  wire u3_u0_r0_21__FF_INPUT;
  wire u3_u0_r0_22_;
  wire u3_u0_r0_22__FF_INPUT;
  wire u3_u0_r0_23_;
  wire u3_u0_r0_23__FF_INPUT;
  wire u3_u0_r0_24_;
  wire u3_u0_r0_24__FF_INPUT;
  wire u3_u0_r0_25_;
  wire u3_u0_r0_25__FF_INPUT;
  wire u3_u0_r0_26_;
  wire u3_u0_r0_26__FF_INPUT;
  wire u3_u0_r0_27_;
  wire u3_u0_r0_27__FF_INPUT;
  wire u3_u0_r0_28_;
  wire u3_u0_r0_28__FF_INPUT;
  wire u3_u0_r0_29_;
  wire u3_u0_r0_29__FF_INPUT;
  wire u3_u0_r0_2_;
  wire u3_u0_r0_2__FF_INPUT;
  wire u3_u0_r0_30_;
  wire u3_u0_r0_30__FF_INPUT;
  wire u3_u0_r0_31_;
  wire u3_u0_r0_31__FF_INPUT;
  wire u3_u0_r0_32_;
  wire u3_u0_r0_32__FF_INPUT;
  wire u3_u0_r0_33_;
  wire u3_u0_r0_33__FF_INPUT;
  wire u3_u0_r0_34_;
  wire u3_u0_r0_34__FF_INPUT;
  wire u3_u0_r0_35_;
  wire u3_u0_r0_35__FF_INPUT;
  wire u3_u0_r0_3_;
  wire u3_u0_r0_3__FF_INPUT;
  wire u3_u0_r0_4_;
  wire u3_u0_r0_4__FF_INPUT;
  wire u3_u0_r0_5_;
  wire u3_u0_r0_5__FF_INPUT;
  wire u3_u0_r0_6_;
  wire u3_u0_r0_6__FF_INPUT;
  wire u3_u0_r0_7_;
  wire u3_u0_r0_7__FF_INPUT;
  wire u3_u0_r0_8_;
  wire u3_u0_r0_8__FF_INPUT;
  wire u3_u0_r0_9_;
  wire u3_u0_r0_9__FF_INPUT;
  wire u3_u0_r1_0_;
  wire u3_u0_r1_0__FF_INPUT;
  wire u3_u0_r1_10_;
  wire u3_u0_r1_10__FF_INPUT;
  wire u3_u0_r1_11_;
  wire u3_u0_r1_11__FF_INPUT;
  wire u3_u0_r1_12_;
  wire u3_u0_r1_12__FF_INPUT;
  wire u3_u0_r1_13_;
  wire u3_u0_r1_13__FF_INPUT;
  wire u3_u0_r1_14_;
  wire u3_u0_r1_14__FF_INPUT;
  wire u3_u0_r1_15_;
  wire u3_u0_r1_15__FF_INPUT;
  wire u3_u0_r1_16_;
  wire u3_u0_r1_16__FF_INPUT;
  wire u3_u0_r1_17_;
  wire u3_u0_r1_17__FF_INPUT;
  wire u3_u0_r1_18_;
  wire u3_u0_r1_18__FF_INPUT;
  wire u3_u0_r1_19_;
  wire u3_u0_r1_19__FF_INPUT;
  wire u3_u0_r1_1_;
  wire u3_u0_r1_1__FF_INPUT;
  wire u3_u0_r1_20_;
  wire u3_u0_r1_20__FF_INPUT;
  wire u3_u0_r1_21_;
  wire u3_u0_r1_21__FF_INPUT;
  wire u3_u0_r1_22_;
  wire u3_u0_r1_22__FF_INPUT;
  wire u3_u0_r1_23_;
  wire u3_u0_r1_23__FF_INPUT;
  wire u3_u0_r1_24_;
  wire u3_u0_r1_24__FF_INPUT;
  wire u3_u0_r1_25_;
  wire u3_u0_r1_25__FF_INPUT;
  wire u3_u0_r1_26_;
  wire u3_u0_r1_26__FF_INPUT;
  wire u3_u0_r1_27_;
  wire u3_u0_r1_27__FF_INPUT;
  wire u3_u0_r1_28_;
  wire u3_u0_r1_28__FF_INPUT;
  wire u3_u0_r1_29_;
  wire u3_u0_r1_29__FF_INPUT;
  wire u3_u0_r1_2_;
  wire u3_u0_r1_2__FF_INPUT;
  wire u3_u0_r1_30_;
  wire u3_u0_r1_30__FF_INPUT;
  wire u3_u0_r1_31_;
  wire u3_u0_r1_31__FF_INPUT;
  wire u3_u0_r1_32_;
  wire u3_u0_r1_32__FF_INPUT;
  wire u3_u0_r1_33_;
  wire u3_u0_r1_33__FF_INPUT;
  wire u3_u0_r1_34_;
  wire u3_u0_r1_34__FF_INPUT;
  wire u3_u0_r1_35_;
  wire u3_u0_r1_35__FF_INPUT;
  wire u3_u0_r1_3_;
  wire u3_u0_r1_3__FF_INPUT;
  wire u3_u0_r1_4_;
  wire u3_u0_r1_4__FF_INPUT;
  wire u3_u0_r1_5_;
  wire u3_u0_r1_5__FF_INPUT;
  wire u3_u0_r1_6_;
  wire u3_u0_r1_6__FF_INPUT;
  wire u3_u0_r1_7_;
  wire u3_u0_r1_7__FF_INPUT;
  wire u3_u0_r1_8_;
  wire u3_u0_r1_8__FF_INPUT;
  wire u3_u0_r1_9_;
  wire u3_u0_r1_9__FF_INPUT;
  wire u3_u0_r2_0_;
  wire u3_u0_r2_0__FF_INPUT;
  wire u3_u0_r2_10_;
  wire u3_u0_r2_10__FF_INPUT;
  wire u3_u0_r2_11_;
  wire u3_u0_r2_11__FF_INPUT;
  wire u3_u0_r2_12_;
  wire u3_u0_r2_12__FF_INPUT;
  wire u3_u0_r2_13_;
  wire u3_u0_r2_13__FF_INPUT;
  wire u3_u0_r2_14_;
  wire u3_u0_r2_14__FF_INPUT;
  wire u3_u0_r2_15_;
  wire u3_u0_r2_15__FF_INPUT;
  wire u3_u0_r2_16_;
  wire u3_u0_r2_16__FF_INPUT;
  wire u3_u0_r2_17_;
  wire u3_u0_r2_17__FF_INPUT;
  wire u3_u0_r2_18_;
  wire u3_u0_r2_18__FF_INPUT;
  wire u3_u0_r2_19_;
  wire u3_u0_r2_19__FF_INPUT;
  wire u3_u0_r2_1_;
  wire u3_u0_r2_1__FF_INPUT;
  wire u3_u0_r2_20_;
  wire u3_u0_r2_20__FF_INPUT;
  wire u3_u0_r2_21_;
  wire u3_u0_r2_21__FF_INPUT;
  wire u3_u0_r2_22_;
  wire u3_u0_r2_22__FF_INPUT;
  wire u3_u0_r2_23_;
  wire u3_u0_r2_23__FF_INPUT;
  wire u3_u0_r2_24_;
  wire u3_u0_r2_24__FF_INPUT;
  wire u3_u0_r2_25_;
  wire u3_u0_r2_25__FF_INPUT;
  wire u3_u0_r2_26_;
  wire u3_u0_r2_26__FF_INPUT;
  wire u3_u0_r2_27_;
  wire u3_u0_r2_27__FF_INPUT;
  wire u3_u0_r2_28_;
  wire u3_u0_r2_28__FF_INPUT;
  wire u3_u0_r2_29_;
  wire u3_u0_r2_29__FF_INPUT;
  wire u3_u0_r2_2_;
  wire u3_u0_r2_2__FF_INPUT;
  wire u3_u0_r2_30_;
  wire u3_u0_r2_30__FF_INPUT;
  wire u3_u0_r2_31_;
  wire u3_u0_r2_31__FF_INPUT;
  wire u3_u0_r2_32_;
  wire u3_u0_r2_32__FF_INPUT;
  wire u3_u0_r2_33_;
  wire u3_u0_r2_33__FF_INPUT;
  wire u3_u0_r2_34_;
  wire u3_u0_r2_34__FF_INPUT;
  wire u3_u0_r2_35_;
  wire u3_u0_r2_35__FF_INPUT;
  wire u3_u0_r2_3_;
  wire u3_u0_r2_3__FF_INPUT;
  wire u3_u0_r2_4_;
  wire u3_u0_r2_4__FF_INPUT;
  wire u3_u0_r2_5_;
  wire u3_u0_r2_5__FF_INPUT;
  wire u3_u0_r2_6_;
  wire u3_u0_r2_6__FF_INPUT;
  wire u3_u0_r2_7_;
  wire u3_u0_r2_7__FF_INPUT;
  wire u3_u0_r2_8_;
  wire u3_u0_r2_8__FF_INPUT;
  wire u3_u0_r2_9_;
  wire u3_u0_r2_9__FF_INPUT;
  wire u3_u0_r3_0_;
  wire u3_u0_r3_0__FF_INPUT;
  wire u3_u0_r3_10_;
  wire u3_u0_r3_10__FF_INPUT;
  wire u3_u0_r3_11_;
  wire u3_u0_r3_11__FF_INPUT;
  wire u3_u0_r3_12_;
  wire u3_u0_r3_12__FF_INPUT;
  wire u3_u0_r3_13_;
  wire u3_u0_r3_13__FF_INPUT;
  wire u3_u0_r3_14_;
  wire u3_u0_r3_14__FF_INPUT;
  wire u3_u0_r3_15_;
  wire u3_u0_r3_15__FF_INPUT;
  wire u3_u0_r3_16_;
  wire u3_u0_r3_16__FF_INPUT;
  wire u3_u0_r3_17_;
  wire u3_u0_r3_17__FF_INPUT;
  wire u3_u0_r3_18_;
  wire u3_u0_r3_18__FF_INPUT;
  wire u3_u0_r3_19_;
  wire u3_u0_r3_19__FF_INPUT;
  wire u3_u0_r3_1_;
  wire u3_u0_r3_1__FF_INPUT;
  wire u3_u0_r3_20_;
  wire u3_u0_r3_20__FF_INPUT;
  wire u3_u0_r3_21_;
  wire u3_u0_r3_21__FF_INPUT;
  wire u3_u0_r3_22_;
  wire u3_u0_r3_22__FF_INPUT;
  wire u3_u0_r3_23_;
  wire u3_u0_r3_23__FF_INPUT;
  wire u3_u0_r3_24_;
  wire u3_u0_r3_24__FF_INPUT;
  wire u3_u0_r3_25_;
  wire u3_u0_r3_25__FF_INPUT;
  wire u3_u0_r3_26_;
  wire u3_u0_r3_26__FF_INPUT;
  wire u3_u0_r3_27_;
  wire u3_u0_r3_27__FF_INPUT;
  wire u3_u0_r3_28_;
  wire u3_u0_r3_28__FF_INPUT;
  wire u3_u0_r3_29_;
  wire u3_u0_r3_29__FF_INPUT;
  wire u3_u0_r3_2_;
  wire u3_u0_r3_2__FF_INPUT;
  wire u3_u0_r3_30_;
  wire u3_u0_r3_30__FF_INPUT;
  wire u3_u0_r3_31_;
  wire u3_u0_r3_31__FF_INPUT;
  wire u3_u0_r3_32_;
  wire u3_u0_r3_32__FF_INPUT;
  wire u3_u0_r3_33_;
  wire u3_u0_r3_33__FF_INPUT;
  wire u3_u0_r3_34_;
  wire u3_u0_r3_34__FF_INPUT;
  wire u3_u0_r3_35_;
  wire u3_u0_r3_35__FF_INPUT;
  wire u3_u0_r3_3_;
  wire u3_u0_r3_3__FF_INPUT;
  wire u3_u0_r3_4_;
  wire u3_u0_r3_4__FF_INPUT;
  wire u3_u0_r3_5_;
  wire u3_u0_r3_5__FF_INPUT;
  wire u3_u0_r3_6_;
  wire u3_u0_r3_6__FF_INPUT;
  wire u3_u0_r3_7_;
  wire u3_u0_r3_7__FF_INPUT;
  wire u3_u0_r3_8_;
  wire u3_u0_r3_8__FF_INPUT;
  wire u3_u0_r3_9_;
  wire u3_u0_r3_9__FF_INPUT;
  wire u3_u0_rd_adr_0_;
  wire u3_u0_rd_adr_0__FF_INPUT;
  wire u3_u0_rd_adr_1_;
  wire u3_u0_rd_adr_1__FF_INPUT;
  wire u3_u0_rd_adr_2_;
  wire u3_u0_rd_adr_2__FF_INPUT;
  wire u3_u0_rd_adr_3_;
  wire u3_u0_rd_adr_3__FF_INPUT;
  wire u3_u0_wr_adr_0_;
  wire u3_u0_wr_adr_0__FF_INPUT;
  wire u3_u0_wr_adr_1_;
  wire u3_u0_wr_adr_1__FF_INPUT;
  wire u3_u0_wr_adr_2_;
  wire u3_u0_wr_adr_2__FF_INPUT;
  wire u3_u0_wr_adr_3_;
  wire u3_u0_wr_adr_3__FF_INPUT;
  wire u3_wb_read_go;
  wire u4__abc_49152_n100;
  wire u4__abc_49152_n101_1;
  wire u4__abc_49152_n102_1;
  wire u4__abc_49152_n103;
  wire u4__abc_49152_n104_1;
  wire u4__abc_49152_n105;
  wire u4__abc_49152_n106;
  wire u4__abc_49152_n107;
  wire u4__abc_49152_n108_1;
  wire u4__abc_49152_n109;
  wire u4__abc_49152_n110;
  wire u4__abc_49152_n111;
  wire u4__abc_49152_n112;
  wire u4__abc_49152_n113_1;
  wire u4__abc_49152_n114;
  wire u4__abc_49152_n115;
  wire u4__abc_49152_n116;
  wire u4__abc_49152_n117;
  wire u4__abc_49152_n119;
  wire u4__abc_49152_n120;
  wire u4__abc_49152_n122;
  wire u4__abc_49152_n123;
  wire u4__abc_49152_n124_1;
  wire u4__abc_49152_n125;
  wire u4__abc_49152_n127;
  wire u4__abc_49152_n128;
  wire u4__abc_49152_n129_1;
  wire u4__abc_49152_n130;
  wire u4__abc_49152_n131;
  wire u4__abc_49152_n133;
  wire u4__abc_49152_n134_1;
  wire u4__abc_49152_n135;
  wire u4__abc_49152_n136;
  wire u4__abc_49152_n137;
  wire u4__abc_49152_n139_1;
  wire u4__abc_49152_n140;
  wire u4__abc_49152_n141_1;
  wire u4__abc_49152_n142;
  wire u4__abc_49152_n143_1;
  wire u4__abc_49152_n145;
  wire u4__abc_49152_n146;
  wire u4__abc_49152_n147;
  wire u4__abc_49152_n148;
  wire u4__abc_49152_n150;
  wire u4__abc_49152_n151;
  wire u4__abc_49152_n152;
  wire u4__abc_49152_n153;
  wire u4__abc_49152_n154;
  wire u4__abc_49152_n156;
  wire u4__abc_49152_n157;
  wire u4__abc_49152_n158;
  wire u4__abc_49152_n159_1;
  wire u4__abc_49152_n161;
  wire u4__abc_49152_n162;
  wire u4__abc_49152_n163;
  wire u4__abc_49152_n164;
  wire u4__abc_49152_n165;
  wire u4__abc_49152_n167;
  wire u4__abc_49152_n168;
  wire u4__abc_49152_n169;
  wire u4__abc_49152_n170;
  wire u4__abc_49152_n171;
  wire u4__abc_49152_n172;
  wire u4__abc_49152_n173;
  wire u4__abc_49152_n174;
  wire u4__abc_49152_n175;
  wire u4__abc_49152_n177;
  wire u4__abc_49152_n178;
  wire u4__abc_49152_n179;
  wire u4__abc_49152_n180;
  wire u4__abc_49152_n182;
  wire u4__abc_49152_n183;
  wire u4__abc_49152_n184;
  wire u4__abc_49152_n185;
  wire u4__abc_49152_n187;
  wire u4__abc_49152_n188;
  wire u4__abc_49152_n189_1;
  wire u4__abc_49152_n191;
  wire u4__abc_49152_n191_1;
  wire u4__abc_49152_n191_bF_buf0;
  wire u4__abc_49152_n191_bF_buf1;
  wire u4__abc_49152_n191_bF_buf2;
  wire u4__abc_49152_n191_bF_buf3;
  wire u4__abc_49152_n192;
  wire u4__abc_49152_n193;
  wire u4__abc_49152_n194;
  wire u4__abc_49152_n195;
  wire u4__abc_49152_n196;
  wire u4__abc_49152_n198;
  wire u4__abc_49152_n199;
  wire u4__abc_49152_n200;
  wire u4__abc_49152_n201;
  wire u4__abc_49152_n202;
  wire u4__abc_49152_n204;
  wire u4__abc_49152_n205;
  wire u4__abc_49152_n206;
  wire u4__abc_49152_n207;
  wire u4__abc_49152_n209;
  wire u4__abc_49152_n210;
  wire u4__abc_49152_n211;
  wire u4__abc_49152_n212;
  wire u4__abc_49152_n213;
  wire u4__abc_49152_n214;
  wire u4__abc_49152_n215;
  wire u4__abc_49152_n216;
  wire u4__abc_49152_n217;
  wire u4__abc_49152_n219;
  wire u4__abc_49152_n220;
  wire u4__abc_49152_n221;
  wire u4__abc_49152_n222;
  wire u4__abc_49152_n224;
  wire u4__abc_49152_n225;
  wire u4__abc_49152_n226;
  wire u4__abc_49152_n227;
  wire u4__abc_49152_n228;
  wire u4__abc_49152_n229;
  wire u4__abc_49152_n230;
  wire u4__abc_49152_n231;
  wire u4__abc_49152_n232;
  wire u4__abc_49152_n233;
  wire u4__abc_49152_n234;
  wire u4__abc_49152_n235;
  wire u4__abc_49152_n236;
  wire u4__abc_49152_n237;
  wire u4__abc_49152_n238;
  wire u4__abc_49152_n239;
  wire u4__abc_49152_n240;
  wire u4__abc_49152_n241;
  wire u4__abc_49152_n242;
  wire u4__abc_49152_n243;
  wire u4__abc_49152_n244;
  wire u4__abc_49152_n245;
  wire u4__abc_49152_n246;
  wire u4__abc_49152_n247;
  wire u4__abc_49152_n248;
  wire u4__abc_49152_n249;
  wire u4__abc_49152_n250;
  wire u4__abc_49152_n251;
  wire u4__abc_49152_n252;
  wire u4__abc_49152_n253;
  wire u4__abc_49152_n254;
  wire u4__abc_49152_n255;
  wire u4__abc_49152_n256;
  wire u4__abc_49152_n65;
  wire u4__abc_49152_n66_1;
  wire u4__abc_49152_n67;
  wire u4__abc_49152_n68;
  wire u4__abc_49152_n69_1;
  wire u4__abc_49152_n70;
  wire u4__abc_49152_n72;
  wire u4__abc_49152_n73_1;
  wire u4__abc_49152_n74;
  wire u4__abc_49152_n75;
  wire u4__abc_49152_n76_1;
  wire u4__abc_49152_n77;
  wire u4__abc_49152_n78;
  wire u4__abc_49152_n79_1;
  wire u4__abc_49152_n80;
  wire u4__abc_49152_n81;
  wire u4__abc_49152_n82_1;
  wire u4__abc_49152_n83;
  wire u4__abc_49152_n84;
  wire u4__abc_49152_n85_1;
  wire u4__abc_49152_n86;
  wire u4__abc_49152_n87;
  wire u4__abc_49152_n88_1;
  wire u4__abc_49152_n89;
  wire u4__abc_49152_n90_1;
  wire u4__abc_49152_n91;
  wire u4__abc_49152_n92;
  wire u4__abc_49152_n93_1;
  wire u4__abc_49152_n94;
  wire u4__abc_49152_n95;
  wire u4__abc_49152_n96;
  wire u4__abc_49152_n97;
  wire u4__abc_49152_n98;
  wire u4__abc_49152_n99;
  wire u4_ps_cnt_0_;
  wire u4_ps_cnt_0__FF_INPUT;
  wire u4_ps_cnt_1_;
  wire u4_ps_cnt_1__FF_INPUT;
  wire u4_ps_cnt_2_;
  wire u4_ps_cnt_2__FF_INPUT;
  wire u4_ps_cnt_3_;
  wire u4_ps_cnt_3__FF_INPUT;
  wire u4_ps_cnt_4_;
  wire u4_ps_cnt_4__FF_INPUT;
  wire u4_ps_cnt_5_;
  wire u4_ps_cnt_5__FF_INPUT;
  wire u4_ps_cnt_6_;
  wire u4_ps_cnt_6__FF_INPUT;
  wire u4_ps_cnt_7_;
  wire u4_ps_cnt_7__FF_INPUT;
  wire u4_ps_cnt_clr;
  wire u4_rfr_ce;
  wire u4_rfr_clr;
  wire u4_rfr_clr_FF_INPUT;
  wire u4_rfr_cnt_0_;
  wire u4_rfr_cnt_0__FF_INPUT;
  wire u4_rfr_cnt_1_;
  wire u4_rfr_cnt_1__FF_INPUT;
  wire u4_rfr_cnt_2_;
  wire u4_rfr_cnt_2__FF_INPUT;
  wire u4_rfr_cnt_3_;
  wire u4_rfr_cnt_3__FF_INPUT;
  wire u4_rfr_cnt_4_;
  wire u4_rfr_cnt_4__FF_INPUT;
  wire u4_rfr_cnt_5_;
  wire u4_rfr_cnt_5__FF_INPUT;
  wire u4_rfr_cnt_6_;
  wire u4_rfr_cnt_6__FF_INPUT;
  wire u4_rfr_cnt_7_;
  wire u4_rfr_cnt_7__FF_INPUT;
  wire u4_rfr_early;
  wire u4_rfr_early_FF_INPUT;
  wire u4_rfr_en;
  wire u4_rfr_en_FF_INPUT;
  wire u4_rfr_req_FF_INPUT;
  wire u5__abc_41027_n1845;
  wire u5__abc_41027_n1846;
  wire u5__abc_41027_n1847;
  wire u5__abc_41027_n1848;
  wire u5__abc_41027_n1849;
  wire u5__abc_41027_n1850;
  wire u5__abc_41027_n1851;
  wire u5__abc_54027_n1000_1;
  wire u5__abc_54027_n1001;
  wire u5__abc_54027_n1002;
  wire u5__abc_54027_n1003;
  wire u5__abc_54027_n1004;
  wire u5__abc_54027_n1005;
  wire u5__abc_54027_n1007;
  wire u5__abc_54027_n1008;
  wire u5__abc_54027_n1009;
  wire u5__abc_54027_n1010;
  wire u5__abc_54027_n1011;
  wire u5__abc_54027_n1012;
  wire u5__abc_54027_n1013;
  wire u5__abc_54027_n1014;
  wire u5__abc_54027_n1015;
  wire u5__abc_54027_n1016;
  wire u5__abc_54027_n1017;
  wire u5__abc_54027_n1018;
  wire u5__abc_54027_n1019;
  wire u5__abc_54027_n1020;
  wire u5__abc_54027_n1021;
  wire u5__abc_54027_n1022;
  wire u5__abc_54027_n1023;
  wire u5__abc_54027_n1024;
  wire u5__abc_54027_n1025;
  wire u5__abc_54027_n1026;
  wire u5__abc_54027_n1027;
  wire u5__abc_54027_n1028;
  wire u5__abc_54027_n1029;
  wire u5__abc_54027_n1030;
  wire u5__abc_54027_n1031;
  wire u5__abc_54027_n1032;
  wire u5__abc_54027_n1033;
  wire u5__abc_54027_n1034;
  wire u5__abc_54027_n1035;
  wire u5__abc_54027_n1036;
  wire u5__abc_54027_n1037;
  wire u5__abc_54027_n1038;
  wire u5__abc_54027_n1040;
  wire u5__abc_54027_n1041;
  wire u5__abc_54027_n1042;
  wire u5__abc_54027_n1043;
  wire u5__abc_54027_n1044;
  wire u5__abc_54027_n1045;
  wire u5__abc_54027_n1046;
  wire u5__abc_54027_n1047;
  wire u5__abc_54027_n1048;
  wire u5__abc_54027_n1049;
  wire u5__abc_54027_n1050;
  wire u5__abc_54027_n1051;
  wire u5__abc_54027_n1052_1;
  wire u5__abc_54027_n1053_1;
  wire u5__abc_54027_n1054;
  wire u5__abc_54027_n1055;
  wire u5__abc_54027_n1057;
  wire u5__abc_54027_n1058_1;
  wire u5__abc_54027_n1059;
  wire u5__abc_54027_n1060;
  wire u5__abc_54027_n1061;
  wire u5__abc_54027_n1062;
  wire u5__abc_54027_n1063;
  wire u5__abc_54027_n1065;
  wire u5__abc_54027_n1066;
  wire u5__abc_54027_n1067;
  wire u5__abc_54027_n1068;
  wire u5__abc_54027_n1069;
  wire u5__abc_54027_n1070;
  wire u5__abc_54027_n1071;
  wire u5__abc_54027_n1072;
  wire u5__abc_54027_n1073;
  wire u5__abc_54027_n1074;
  wire u5__abc_54027_n1075;
  wire u5__abc_54027_n1077;
  wire u5__abc_54027_n1078;
  wire u5__abc_54027_n1079;
  wire u5__abc_54027_n1080;
  wire u5__abc_54027_n1081;
  wire u5__abc_54027_n1082;
  wire u5__abc_54027_n1084;
  wire u5__abc_54027_n1085;
  wire u5__abc_54027_n1086;
  wire u5__abc_54027_n1087;
  wire u5__abc_54027_n1088;
  wire u5__abc_54027_n1089;
  wire u5__abc_54027_n1090;
  wire u5__abc_54027_n1091;
  wire u5__abc_54027_n1092;
  wire u5__abc_54027_n1093;
  wire u5__abc_54027_n1094;
  wire u5__abc_54027_n1095;
  wire u5__abc_54027_n1096;
  wire u5__abc_54027_n1097;
  wire u5__abc_54027_n1098;
  wire u5__abc_54027_n1099;
  wire u5__abc_54027_n1100;
  wire u5__abc_54027_n1101;
  wire u5__abc_54027_n1102;
  wire u5__abc_54027_n1103;
  wire u5__abc_54027_n1104;
  wire u5__abc_54027_n1105;
  wire u5__abc_54027_n1106;
  wire u5__abc_54027_n1107;
  wire u5__abc_54027_n1108;
  wire u5__abc_54027_n1109;
  wire u5__abc_54027_n1110;
  wire u5__abc_54027_n1111;
  wire u5__abc_54027_n1112;
  wire u5__abc_54027_n1113;
  wire u5__abc_54027_n1114;
  wire u5__abc_54027_n1115;
  wire u5__abc_54027_n1116;
  wire u5__abc_54027_n1117;
  wire u5__abc_54027_n1119;
  wire u5__abc_54027_n1120;
  wire u5__abc_54027_n1121;
  wire u5__abc_54027_n1122;
  wire u5__abc_54027_n1123;
  wire u5__abc_54027_n1124;
  wire u5__abc_54027_n1125;
  wire u5__abc_54027_n1126;
  wire u5__abc_54027_n1127;
  wire u5__abc_54027_n1128;
  wire u5__abc_54027_n1129;
  wire u5__abc_54027_n1130;
  wire u5__abc_54027_n1131;
  wire u5__abc_54027_n1132;
  wire u5__abc_54027_n1133;
  wire u5__abc_54027_n1134;
  wire u5__abc_54027_n1135;
  wire u5__abc_54027_n1136;
  wire u5__abc_54027_n1137;
  wire u5__abc_54027_n1138;
  wire u5__abc_54027_n1139;
  wire u5__abc_54027_n1140;
  wire u5__abc_54027_n1142;
  wire u5__abc_54027_n1143;
  wire u5__abc_54027_n1144;
  wire u5__abc_54027_n1145;
  wire u5__abc_54027_n1146;
  wire u5__abc_54027_n1147;
  wire u5__abc_54027_n1148;
  wire u5__abc_54027_n1149;
  wire u5__abc_54027_n1150;
  wire u5__abc_54027_n1151;
  wire u5__abc_54027_n1152;
  wire u5__abc_54027_n1153;
  wire u5__abc_54027_n1154;
  wire u5__abc_54027_n1155;
  wire u5__abc_54027_n1156;
  wire u5__abc_54027_n1157;
  wire u5__abc_54027_n1158;
  wire u5__abc_54027_n1159;
  wire u5__abc_54027_n1160;
  wire u5__abc_54027_n1161;
  wire u5__abc_54027_n1162;
  wire u5__abc_54027_n1163;
  wire u5__abc_54027_n1165;
  wire u5__abc_54027_n1166;
  wire u5__abc_54027_n1167;
  wire u5__abc_54027_n1168;
  wire u5__abc_54027_n1169;
  wire u5__abc_54027_n1170;
  wire u5__abc_54027_n1171;
  wire u5__abc_54027_n1172;
  wire u5__abc_54027_n1173;
  wire u5__abc_54027_n1174;
  wire u5__abc_54027_n1175;
  wire u5__abc_54027_n1176;
  wire u5__abc_54027_n1177;
  wire u5__abc_54027_n1178;
  wire u5__abc_54027_n1179;
  wire u5__abc_54027_n1180;
  wire u5__abc_54027_n1181;
  wire u5__abc_54027_n1182;
  wire u5__abc_54027_n1183;
  wire u5__abc_54027_n1184;
  wire u5__abc_54027_n1185;
  wire u5__abc_54027_n1187;
  wire u5__abc_54027_n1188;
  wire u5__abc_54027_n1189;
  wire u5__abc_54027_n1190;
  wire u5__abc_54027_n1191;
  wire u5__abc_54027_n1192;
  wire u5__abc_54027_n1193;
  wire u5__abc_54027_n1194;
  wire u5__abc_54027_n1195;
  wire u5__abc_54027_n1196;
  wire u5__abc_54027_n1197;
  wire u5__abc_54027_n1198;
  wire u5__abc_54027_n1199;
  wire u5__abc_54027_n1200;
  wire u5__abc_54027_n1201;
  wire u5__abc_54027_n1202;
  wire u5__abc_54027_n1203;
  wire u5__abc_54027_n1204;
  wire u5__abc_54027_n1205_1;
  wire u5__abc_54027_n1207;
  wire u5__abc_54027_n1208;
  wire u5__abc_54027_n1209;
  wire u5__abc_54027_n1210;
  wire u5__abc_54027_n1211;
  wire u5__abc_54027_n1212;
  wire u5__abc_54027_n1213;
  wire u5__abc_54027_n1214;
  wire u5__abc_54027_n1215;
  wire u5__abc_54027_n1216;
  wire u5__abc_54027_n1217;
  wire u5__abc_54027_n1218;
  wire u5__abc_54027_n1219;
  wire u5__abc_54027_n1221;
  wire u5__abc_54027_n1222;
  wire u5__abc_54027_n1223;
  wire u5__abc_54027_n1224;
  wire u5__abc_54027_n1225;
  wire u5__abc_54027_n1226;
  wire u5__abc_54027_n1227;
  wire u5__abc_54027_n1228;
  wire u5__abc_54027_n1229;
  wire u5__abc_54027_n1230;
  wire u5__abc_54027_n1232;
  wire u5__abc_54027_n1233_1;
  wire u5__abc_54027_n1234;
  wire u5__abc_54027_n1235_1;
  wire u5__abc_54027_n1236;
  wire u5__abc_54027_n1237;
  wire u5__abc_54027_n1238;
  wire u5__abc_54027_n1239;
  wire u5__abc_54027_n1240;
  wire u5__abc_54027_n1242;
  wire u5__abc_54027_n1243;
  wire u5__abc_54027_n1244;
  wire u5__abc_54027_n1245;
  wire u5__abc_54027_n1246;
  wire u5__abc_54027_n1247;
  wire u5__abc_54027_n1249;
  wire u5__abc_54027_n1250;
  wire u5__abc_54027_n1251;
  wire u5__abc_54027_n1252;
  wire u5__abc_54027_n1253;
  wire u5__abc_54027_n1254;
  wire u5__abc_54027_n1255;
  wire u5__abc_54027_n1256;
  wire u5__abc_54027_n1257;
  wire u5__abc_54027_n1259;
  wire u5__abc_54027_n1260;
  wire u5__abc_54027_n1261;
  wire u5__abc_54027_n1262;
  wire u5__abc_54027_n1263;
  wire u5__abc_54027_n1264;
  wire u5__abc_54027_n1265;
  wire u5__abc_54027_n1267;
  wire u5__abc_54027_n1268;
  wire u5__abc_54027_n1269;
  wire u5__abc_54027_n1270;
  wire u5__abc_54027_n1271;
  wire u5__abc_54027_n1272;
  wire u5__abc_54027_n1273;
  wire u5__abc_54027_n1274;
  wire u5__abc_54027_n1276;
  wire u5__abc_54027_n1277;
  wire u5__abc_54027_n1278;
  wire u5__abc_54027_n1279;
  wire u5__abc_54027_n1280;
  wire u5__abc_54027_n1281;
  wire u5__abc_54027_n1282;
  wire u5__abc_54027_n1283;
  wire u5__abc_54027_n1285;
  wire u5__abc_54027_n1286;
  wire u5__abc_54027_n1288;
  wire u5__abc_54027_n1289;
  wire u5__abc_54027_n1291;
  wire u5__abc_54027_n1292;
  wire u5__abc_54027_n1294;
  wire u5__abc_54027_n1295;
  wire u5__abc_54027_n1296;
  wire u5__abc_54027_n1297;
  wire u5__abc_54027_n1298;
  wire u5__abc_54027_n1299;
  wire u5__abc_54027_n1300;
  wire u5__abc_54027_n1301;
  wire u5__abc_54027_n1303;
  wire u5__abc_54027_n1304;
  wire u5__abc_54027_n1306;
  wire u5__abc_54027_n1307;
  wire u5__abc_54027_n1308;
  wire u5__abc_54027_n1309;
  wire u5__abc_54027_n1310;
  wire u5__abc_54027_n1311;
  wire u5__abc_54027_n1312_1;
  wire u5__abc_54027_n1313;
  wire u5__abc_54027_n1314;
  wire u5__abc_54027_n1315;
  wire u5__abc_54027_n1316;
  wire u5__abc_54027_n1317;
  wire u5__abc_54027_n1318;
  wire u5__abc_54027_n1319;
  wire u5__abc_54027_n1320;
  wire u5__abc_54027_n1321;
  wire u5__abc_54027_n1322;
  wire u5__abc_54027_n1323;
  wire u5__abc_54027_n1324;
  wire u5__abc_54027_n1325;
  wire u5__abc_54027_n1326;
  wire u5__abc_54027_n1327;
  wire u5__abc_54027_n1328;
  wire u5__abc_54027_n1329;
  wire u5__abc_54027_n1330;
  wire u5__abc_54027_n1331;
  wire u5__abc_54027_n1332;
  wire u5__abc_54027_n1333;
  wire u5__abc_54027_n1334;
  wire u5__abc_54027_n1335;
  wire u5__abc_54027_n1336;
  wire u5__abc_54027_n1337;
  wire u5__abc_54027_n1338;
  wire u5__abc_54027_n1339;
  wire u5__abc_54027_n1340;
  wire u5__abc_54027_n1341_1;
  wire u5__abc_54027_n1342;
  wire u5__abc_54027_n1343;
  wire u5__abc_54027_n1344;
  wire u5__abc_54027_n1345;
  wire u5__abc_54027_n1346;
  wire u5__abc_54027_n1347;
  wire u5__abc_54027_n1348;
  wire u5__abc_54027_n1349;
  wire u5__abc_54027_n1350;
  wire u5__abc_54027_n1351;
  wire u5__abc_54027_n1352;
  wire u5__abc_54027_n1353;
  wire u5__abc_54027_n1354;
  wire u5__abc_54027_n1355;
  wire u5__abc_54027_n1356;
  wire u5__abc_54027_n1357;
  wire u5__abc_54027_n1358;
  wire u5__abc_54027_n1359;
  wire u5__abc_54027_n1360;
  wire u5__abc_54027_n1361;
  wire u5__abc_54027_n1362;
  wire u5__abc_54027_n1363;
  wire u5__abc_54027_n1364_1;
  wire u5__abc_54027_n1365;
  wire u5__abc_54027_n1366;
  wire u5__abc_54027_n1367;
  wire u5__abc_54027_n1368;
  wire u5__abc_54027_n1369;
  wire u5__abc_54027_n1370;
  wire u5__abc_54027_n1371;
  wire u5__abc_54027_n1372;
  wire u5__abc_54027_n1373_1;
  wire u5__abc_54027_n1374;
  wire u5__abc_54027_n1375;
  wire u5__abc_54027_n1376;
  wire u5__abc_54027_n1377;
  wire u5__abc_54027_n1378_1;
  wire u5__abc_54027_n1379;
  wire u5__abc_54027_n1380_1;
  wire u5__abc_54027_n1381_1;
  wire u5__abc_54027_n1382;
  wire u5__abc_54027_n1383_1;
  wire u5__abc_54027_n1384;
  wire u5__abc_54027_n1385;
  wire u5__abc_54027_n1386;
  wire u5__abc_54027_n1387;
  wire u5__abc_54027_n1388;
  wire u5__abc_54027_n1389;
  wire u5__abc_54027_n1390;
  wire u5__abc_54027_n1391_1;
  wire u5__abc_54027_n1392;
  wire u5__abc_54027_n1393;
  wire u5__abc_54027_n1394;
  wire u5__abc_54027_n1395;
  wire u5__abc_54027_n1396_1;
  wire u5__abc_54027_n1397;
  wire u5__abc_54027_n1398;
  wire u5__abc_54027_n1399;
  wire u5__abc_54027_n1400;
  wire u5__abc_54027_n1401;
  wire u5__abc_54027_n1402;
  wire u5__abc_54027_n1403;
  wire u5__abc_54027_n1404;
  wire u5__abc_54027_n1405;
  wire u5__abc_54027_n1406;
  wire u5__abc_54027_n1407_1;
  wire u5__abc_54027_n1408;
  wire u5__abc_54027_n1409;
  wire u5__abc_54027_n1410;
  wire u5__abc_54027_n1411;
  wire u5__abc_54027_n1412_1;
  wire u5__abc_54027_n1413;
  wire u5__abc_54027_n1414;
  wire u5__abc_54027_n1415;
  wire u5__abc_54027_n1416;
  wire u5__abc_54027_n1417;
  wire u5__abc_54027_n1418;
  wire u5__abc_54027_n1419;
  wire u5__abc_54027_n1420;
  wire u5__abc_54027_n1421;
  wire u5__abc_54027_n1422;
  wire u5__abc_54027_n1423;
  wire u5__abc_54027_n1424;
  wire u5__abc_54027_n1425;
  wire u5__abc_54027_n1426;
  wire u5__abc_54027_n1427;
  wire u5__abc_54027_n1428;
  wire u5__abc_54027_n1429;
  wire u5__abc_54027_n1430;
  wire u5__abc_54027_n1431;
  wire u5__abc_54027_n1432;
  wire u5__abc_54027_n1433;
  wire u5__abc_54027_n1434;
  wire u5__abc_54027_n1435;
  wire u5__abc_54027_n1436;
  wire u5__abc_54027_n1437;
  wire u5__abc_54027_n1438_1;
  wire u5__abc_54027_n1439;
  wire u5__abc_54027_n1440;
  wire u5__abc_54027_n1441;
  wire u5__abc_54027_n1442;
  wire u5__abc_54027_n1443;
  wire u5__abc_54027_n1444;
  wire u5__abc_54027_n1445_1;
  wire u5__abc_54027_n1446;
  wire u5__abc_54027_n1447;
  wire u5__abc_54027_n1448_1;
  wire u5__abc_54027_n1449;
  wire u5__abc_54027_n1450_1;
  wire u5__abc_54027_n1451;
  wire u5__abc_54027_n1452;
  wire u5__abc_54027_n1453;
  wire u5__abc_54027_n1454_1;
  wire u5__abc_54027_n1455_1;
  wire u5__abc_54027_n1456;
  wire u5__abc_54027_n1457;
  wire u5__abc_54027_n1458;
  wire u5__abc_54027_n1459;
  wire u5__abc_54027_n1460;
  wire u5__abc_54027_n1461;
  wire u5__abc_54027_n1462;
  wire u5__abc_54027_n1463;
  wire u5__abc_54027_n1464;
  wire u5__abc_54027_n1465;
  wire u5__abc_54027_n1466;
  wire u5__abc_54027_n1467_1;
  wire u5__abc_54027_n1468;
  wire u5__abc_54027_n1469;
  wire u5__abc_54027_n1470;
  wire u5__abc_54027_n1471;
  wire u5__abc_54027_n1472;
  wire u5__abc_54027_n1473;
  wire u5__abc_54027_n1474;
  wire u5__abc_54027_n1475;
  wire u5__abc_54027_n1476_1;
  wire u5__abc_54027_n1477;
  wire u5__abc_54027_n1478;
  wire u5__abc_54027_n1479;
  wire u5__abc_54027_n1480;
  wire u5__abc_54027_n1481;
  wire u5__abc_54027_n1482;
  wire u5__abc_54027_n1483;
  wire u5__abc_54027_n1484;
  wire u5__abc_54027_n1485;
  wire u5__abc_54027_n1486;
  wire u5__abc_54027_n1487;
  wire u5__abc_54027_n1488;
  wire u5__abc_54027_n1489;
  wire u5__abc_54027_n1490;
  wire u5__abc_54027_n1491_1;
  wire u5__abc_54027_n1492;
  wire u5__abc_54027_n1493;
  wire u5__abc_54027_n1494;
  wire u5__abc_54027_n1495;
  wire u5__abc_54027_n1496;
  wire u5__abc_54027_n1497;
  wire u5__abc_54027_n1498;
  wire u5__abc_54027_n1499;
  wire u5__abc_54027_n1500;
  wire u5__abc_54027_n1501;
  wire u5__abc_54027_n1502;
  wire u5__abc_54027_n1503;
  wire u5__abc_54027_n1504;
  wire u5__abc_54027_n1505;
  wire u5__abc_54027_n1506;
  wire u5__abc_54027_n1507;
  wire u5__abc_54027_n1508;
  wire u5__abc_54027_n1509;
  wire u5__abc_54027_n1510;
  wire u5__abc_54027_n1511;
  wire u5__abc_54027_n1512;
  wire u5__abc_54027_n1513;
  wire u5__abc_54027_n1514;
  wire u5__abc_54027_n1515;
  wire u5__abc_54027_n1516;
  wire u5__abc_54027_n1517;
  wire u5__abc_54027_n1518;
  wire u5__abc_54027_n1519;
  wire u5__abc_54027_n1520;
  wire u5__abc_54027_n1521;
  wire u5__abc_54027_n1522;
  wire u5__abc_54027_n1523;
  wire u5__abc_54027_n1524;
  wire u5__abc_54027_n1525;
  wire u5__abc_54027_n1526;
  wire u5__abc_54027_n1527;
  wire u5__abc_54027_n1528;
  wire u5__abc_54027_n1529;
  wire u5__abc_54027_n1530;
  wire u5__abc_54027_n1531;
  wire u5__abc_54027_n1532;
  wire u5__abc_54027_n1533_1;
  wire u5__abc_54027_n1534;
  wire u5__abc_54027_n1535;
  wire u5__abc_54027_n1536;
  wire u5__abc_54027_n1537_1;
  wire u5__abc_54027_n1538;
  wire u5__abc_54027_n1539;
  wire u5__abc_54027_n1540_1;
  wire u5__abc_54027_n1541_1;
  wire u5__abc_54027_n1542_1;
  wire u5__abc_54027_n1543;
  wire u5__abc_54027_n1544_1;
  wire u5__abc_54027_n1545;
  wire u5__abc_54027_n1547_1;
  wire u5__abc_54027_n1548;
  wire u5__abc_54027_n1549;
  wire u5__abc_54027_n1550;
  wire u5__abc_54027_n1551_1;
  wire u5__abc_54027_n1552_1;
  wire u5__abc_54027_n1553;
  wire u5__abc_54027_n1554_1;
  wire u5__abc_54027_n1555_1;
  wire u5__abc_54027_n1556;
  wire u5__abc_54027_n1557;
  wire u5__abc_54027_n1558_1;
  wire u5__abc_54027_n1559;
  wire u5__abc_54027_n1560;
  wire u5__abc_54027_n1561_1;
  wire u5__abc_54027_n1562_1;
  wire u5__abc_54027_n1563;
  wire u5__abc_54027_n1564;
  wire u5__abc_54027_n1565;
  wire u5__abc_54027_n1566;
  wire u5__abc_54027_n1567;
  wire u5__abc_54027_n1568;
  wire u5__abc_54027_n1569;
  wire u5__abc_54027_n1570;
  wire u5__abc_54027_n1571_1;
  wire u5__abc_54027_n1572_1;
  wire u5__abc_54027_n1573;
  wire u5__abc_54027_n1573_1;
  wire u5__abc_54027_n1574_1;
  wire u5__abc_54027_n1575;
  wire u5__abc_54027_n1575_1;
  wire u5__abc_54027_n1575_bF_buf0;
  wire u5__abc_54027_n1575_bF_buf1;
  wire u5__abc_54027_n1575_bF_buf2;
  wire u5__abc_54027_n1575_bF_buf3;
  wire u5__abc_54027_n1575_bF_buf4;
  wire u5__abc_54027_n1575_bF_buf5;
  wire u5__abc_54027_n1575_bF_buf6;
  wire u5__abc_54027_n1576;
  wire u5__abc_54027_n1577;
  wire u5__abc_54027_n1578;
  wire u5__abc_54027_n1579;
  wire u5__abc_54027_n1580;
  wire u5__abc_54027_n1581;
  wire u5__abc_54027_n1582;
  wire u5__abc_54027_n1583;
  wire u5__abc_54027_n1584;
  wire u5__abc_54027_n1585;
  wire u5__abc_54027_n1586;
  wire u5__abc_54027_n1587;
  wire u5__abc_54027_n1588;
  wire u5__abc_54027_n1589;
  wire u5__abc_54027_n1590;
  wire u5__abc_54027_n1591;
  wire u5__abc_54027_n1592;
  wire u5__abc_54027_n1593;
  wire u5__abc_54027_n1594;
  wire u5__abc_54027_n1595;
  wire u5__abc_54027_n1596;
  wire u5__abc_54027_n1597;
  wire u5__abc_54027_n1598;
  wire u5__abc_54027_n1599;
  wire u5__abc_54027_n1600;
  wire u5__abc_54027_n1601;
  wire u5__abc_54027_n1602;
  wire u5__abc_54027_n1603;
  wire u5__abc_54027_n1604;
  wire u5__abc_54027_n1605;
  wire u5__abc_54027_n1606;
  wire u5__abc_54027_n1607;
  wire u5__abc_54027_n1608;
  wire u5__abc_54027_n1609;
  wire u5__abc_54027_n1610;
  wire u5__abc_54027_n1611;
  wire u5__abc_54027_n1612;
  wire u5__abc_54027_n1613;
  wire u5__abc_54027_n1614;
  wire u5__abc_54027_n1615;
  wire u5__abc_54027_n1616;
  wire u5__abc_54027_n1617;
  wire u5__abc_54027_n1618;
  wire u5__abc_54027_n1619;
  wire u5__abc_54027_n1620;
  wire u5__abc_54027_n1621;
  wire u5__abc_54027_n1622;
  wire u5__abc_54027_n1623;
  wire u5__abc_54027_n1624;
  wire u5__abc_54027_n1625;
  wire u5__abc_54027_n1626;
  wire u5__abc_54027_n1627;
  wire u5__abc_54027_n1628;
  wire u5__abc_54027_n1629;
  wire u5__abc_54027_n1630;
  wire u5__abc_54027_n1631;
  wire u5__abc_54027_n1632;
  wire u5__abc_54027_n1633;
  wire u5__abc_54027_n1634;
  wire u5__abc_54027_n1635;
  wire u5__abc_54027_n1636;
  wire u5__abc_54027_n1637;
  wire u5__abc_54027_n1638;
  wire u5__abc_54027_n1639;
  wire u5__abc_54027_n1640;
  wire u5__abc_54027_n1641;
  wire u5__abc_54027_n1642;
  wire u5__abc_54027_n1643;
  wire u5__abc_54027_n1644;
  wire u5__abc_54027_n1645;
  wire u5__abc_54027_n1646;
  wire u5__abc_54027_n1647;
  wire u5__abc_54027_n1648;
  wire u5__abc_54027_n1649;
  wire u5__abc_54027_n1650;
  wire u5__abc_54027_n1651;
  wire u5__abc_54027_n1652;
  wire u5__abc_54027_n1653;
  wire u5__abc_54027_n1654;
  wire u5__abc_54027_n1655;
  wire u5__abc_54027_n1656;
  wire u5__abc_54027_n1657;
  wire u5__abc_54027_n1658;
  wire u5__abc_54027_n1659;
  wire u5__abc_54027_n1660;
  wire u5__abc_54027_n1661;
  wire u5__abc_54027_n1662;
  wire u5__abc_54027_n1663;
  wire u5__abc_54027_n1664;
  wire u5__abc_54027_n1665;
  wire u5__abc_54027_n1666;
  wire u5__abc_54027_n1667;
  wire u5__abc_54027_n1668;
  wire u5__abc_54027_n1669;
  wire u5__abc_54027_n1670;
  wire u5__abc_54027_n1672;
  wire u5__abc_54027_n1673;
  wire u5__abc_54027_n1674;
  wire u5__abc_54027_n1675;
  wire u5__abc_54027_n1676;
  wire u5__abc_54027_n1677;
  wire u5__abc_54027_n1678;
  wire u5__abc_54027_n1679;
  wire u5__abc_54027_n1680;
  wire u5__abc_54027_n1681;
  wire u5__abc_54027_n1682;
  wire u5__abc_54027_n1683;
  wire u5__abc_54027_n1684;
  wire u5__abc_54027_n1685;
  wire u5__abc_54027_n1686;
  wire u5__abc_54027_n1687;
  wire u5__abc_54027_n1688;
  wire u5__abc_54027_n1689;
  wire u5__abc_54027_n1690;
  wire u5__abc_54027_n1691;
  wire u5__abc_54027_n1692;
  wire u5__abc_54027_n1693;
  wire u5__abc_54027_n1694;
  wire u5__abc_54027_n1695;
  wire u5__abc_54027_n1696;
  wire u5__abc_54027_n1697;
  wire u5__abc_54027_n1698;
  wire u5__abc_54027_n1699;
  wire u5__abc_54027_n1700;
  wire u5__abc_54027_n1701;
  wire u5__abc_54027_n1702;
  wire u5__abc_54027_n1703;
  wire u5__abc_54027_n1704;
  wire u5__abc_54027_n1705;
  wire u5__abc_54027_n1706;
  wire u5__abc_54027_n1707;
  wire u5__abc_54027_n1708;
  wire u5__abc_54027_n1709;
  wire u5__abc_54027_n1710;
  wire u5__abc_54027_n1711;
  wire u5__abc_54027_n1712;
  wire u5__abc_54027_n1713;
  wire u5__abc_54027_n1714;
  wire u5__abc_54027_n1715;
  wire u5__abc_54027_n1716;
  wire u5__abc_54027_n1717;
  wire u5__abc_54027_n1718;
  wire u5__abc_54027_n1719;
  wire u5__abc_54027_n1720;
  wire u5__abc_54027_n1721;
  wire u5__abc_54027_n1722;
  wire u5__abc_54027_n1723;
  wire u5__abc_54027_n1724;
  wire u5__abc_54027_n1725;
  wire u5__abc_54027_n1726;
  wire u5__abc_54027_n1727;
  wire u5__abc_54027_n1728;
  wire u5__abc_54027_n1729;
  wire u5__abc_54027_n1730;
  wire u5__abc_54027_n1731;
  wire u5__abc_54027_n1732;
  wire u5__abc_54027_n1733;
  wire u5__abc_54027_n1734;
  wire u5__abc_54027_n1735;
  wire u5__abc_54027_n1736;
  wire u5__abc_54027_n1737;
  wire u5__abc_54027_n1738;
  wire u5__abc_54027_n1739;
  wire u5__abc_54027_n1740;
  wire u5__abc_54027_n1741;
  wire u5__abc_54027_n1742;
  wire u5__abc_54027_n1743;
  wire u5__abc_54027_n1744;
  wire u5__abc_54027_n1745;
  wire u5__abc_54027_n1747;
  wire u5__abc_54027_n1748;
  wire u5__abc_54027_n1749;
  wire u5__abc_54027_n1750;
  wire u5__abc_54027_n1751;
  wire u5__abc_54027_n1752;
  wire u5__abc_54027_n1753;
  wire u5__abc_54027_n1754;
  wire u5__abc_54027_n1755;
  wire u5__abc_54027_n1756;
  wire u5__abc_54027_n1757;
  wire u5__abc_54027_n1758;
  wire u5__abc_54027_n1759;
  wire u5__abc_54027_n1760;
  wire u5__abc_54027_n1761;
  wire u5__abc_54027_n1762;
  wire u5__abc_54027_n1763;
  wire u5__abc_54027_n1764;
  wire u5__abc_54027_n1765;
  wire u5__abc_54027_n1766;
  wire u5__abc_54027_n1767;
  wire u5__abc_54027_n1768;
  wire u5__abc_54027_n1769;
  wire u5__abc_54027_n1770;
  wire u5__abc_54027_n1771;
  wire u5__abc_54027_n1772;
  wire u5__abc_54027_n1773;
  wire u5__abc_54027_n1774;
  wire u5__abc_54027_n1775;
  wire u5__abc_54027_n1776;
  wire u5__abc_54027_n1777;
  wire u5__abc_54027_n1778;
  wire u5__abc_54027_n1779;
  wire u5__abc_54027_n1780;
  wire u5__abc_54027_n1781;
  wire u5__abc_54027_n1782;
  wire u5__abc_54027_n1783;
  wire u5__abc_54027_n1784;
  wire u5__abc_54027_n1786;
  wire u5__abc_54027_n1787;
  wire u5__abc_54027_n1788;
  wire u5__abc_54027_n1789;
  wire u5__abc_54027_n1790;
  wire u5__abc_54027_n1791;
  wire u5__abc_54027_n1792;
  wire u5__abc_54027_n1793;
  wire u5__abc_54027_n1794;
  wire u5__abc_54027_n1795;
  wire u5__abc_54027_n1796;
  wire u5__abc_54027_n1797;
  wire u5__abc_54027_n1798;
  wire u5__abc_54027_n1799;
  wire u5__abc_54027_n1800;
  wire u5__abc_54027_n1801;
  wire u5__abc_54027_n1802;
  wire u5__abc_54027_n1803;
  wire u5__abc_54027_n1804;
  wire u5__abc_54027_n1805;
  wire u5__abc_54027_n1806;
  wire u5__abc_54027_n1807;
  wire u5__abc_54027_n1809;
  wire u5__abc_54027_n1810;
  wire u5__abc_54027_n1811;
  wire u5__abc_54027_n1812;
  wire u5__abc_54027_n1813;
  wire u5__abc_54027_n1814;
  wire u5__abc_54027_n1815;
  wire u5__abc_54027_n1816;
  wire u5__abc_54027_n1817;
  wire u5__abc_54027_n1818;
  wire u5__abc_54027_n1819;
  wire u5__abc_54027_n1820;
  wire u5__abc_54027_n1821;
  wire u5__abc_54027_n1823;
  wire u5__abc_54027_n1824;
  wire u5__abc_54027_n1825;
  wire u5__abc_54027_n1826;
  wire u5__abc_54027_n1827;
  wire u5__abc_54027_n1828;
  wire u5__abc_54027_n1829;
  wire u5__abc_54027_n1830;
  wire u5__abc_54027_n1831;
  wire u5__abc_54027_n1832;
  wire u5__abc_54027_n1833;
  wire u5__abc_54027_n1834;
  wire u5__abc_54027_n1835;
  wire u5__abc_54027_n1836;
  wire u5__abc_54027_n1837;
  wire u5__abc_54027_n1838;
  wire u5__abc_54027_n1839;
  wire u5__abc_54027_n1840;
  wire u5__abc_54027_n1841;
  wire u5__abc_54027_n1842;
  wire u5__abc_54027_n1843;
  wire u5__abc_54027_n1844;
  wire u5__abc_54027_n1845;
  wire u5__abc_54027_n1846;
  wire u5__abc_54027_n1847;
  wire u5__abc_54027_n1848;
  wire u5__abc_54027_n1849;
  wire u5__abc_54027_n1850;
  wire u5__abc_54027_n1851;
  wire u5__abc_54027_n1853;
  wire u5__abc_54027_n1855;
  wire u5__abc_54027_n1856;
  wire u5__abc_54027_n1857;
  wire u5__abc_54027_n1858;
  wire u5__abc_54027_n1859;
  wire u5__abc_54027_n1860;
  wire u5__abc_54027_n1861;
  wire u5__abc_54027_n1862;
  wire u5__abc_54027_n1863;
  wire u5__abc_54027_n1865;
  wire u5__abc_54027_n1866;
  wire u5__abc_54027_n1868;
  wire u5__abc_54027_n1869;
  wire u5__abc_54027_n1870;
  wire u5__abc_54027_n1871;
  wire u5__abc_54027_n1872;
  wire u5__abc_54027_n1873;
  wire u5__abc_54027_n1875;
  wire u5__abc_54027_n1876;
  wire u5__abc_54027_n1877;
  wire u5__abc_54027_n1878;
  wire u5__abc_54027_n1879;
  wire u5__abc_54027_n1880;
  wire u5__abc_54027_n1881;
  wire u5__abc_54027_n1883;
  wire u5__abc_54027_n1884;
  wire u5__abc_54027_n1885;
  wire u5__abc_54027_n1886;
  wire u5__abc_54027_n1887;
  wire u5__abc_54027_n1888;
  wire u5__abc_54027_n1889;
  wire u5__abc_54027_n1890;
  wire u5__abc_54027_n1891;
  wire u5__abc_54027_n1892;
  wire u5__abc_54027_n1893;
  wire u5__abc_54027_n1894;
  wire u5__abc_54027_n1895;
  wire u5__abc_54027_n1896;
  wire u5__abc_54027_n1897;
  wire u5__abc_54027_n1898;
  wire u5__abc_54027_n1899;
  wire u5__abc_54027_n1900;
  wire u5__abc_54027_n1901;
  wire u5__abc_54027_n1902;
  wire u5__abc_54027_n1904;
  wire u5__abc_54027_n1905;
  wire u5__abc_54027_n1906;
  wire u5__abc_54027_n1908;
  wire u5__abc_54027_n1909;
  wire u5__abc_54027_n1911;
  wire u5__abc_54027_n1913;
  wire u5__abc_54027_n1914;
  wire u5__abc_54027_n1915;
  wire u5__abc_54027_n1918;
  wire u5__abc_54027_n1919;
  wire u5__abc_54027_n1920;
  wire u5__abc_54027_n1921;
  wire u5__abc_54027_n1922;
  wire u5__abc_54027_n1923;
  wire u5__abc_54027_n1924;
  wire u5__abc_54027_n1925;
  wire u5__abc_54027_n1926;
  wire u5__abc_54027_n1927;
  wire u5__abc_54027_n1928;
  wire u5__abc_54027_n1929;
  wire u5__abc_54027_n1930;
  wire u5__abc_54027_n1931;
  wire u5__abc_54027_n1933;
  wire u5__abc_54027_n1934;
  wire u5__abc_54027_n1935;
  wire u5__abc_54027_n1936;
  wire u5__abc_54027_n1937;
  wire u5__abc_54027_n1938;
  wire u5__abc_54027_n1939;
  wire u5__abc_54027_n1941;
  wire u5__abc_54027_n1942;
  wire u5__abc_54027_n1943;
  wire u5__abc_54027_n1944;
  wire u5__abc_54027_n1945;
  wire u5__abc_54027_n1946;
  wire u5__abc_54027_n1947;
  wire u5__abc_54027_n1948;
  wire u5__abc_54027_n1949;
  wire u5__abc_54027_n1950;
  wire u5__abc_54027_n1951;
  wire u5__abc_54027_n1952;
  wire u5__abc_54027_n1953;
  wire u5__abc_54027_n1954;
  wire u5__abc_54027_n1955;
  wire u5__abc_54027_n1956;
  wire u5__abc_54027_n1957;
  wire u5__abc_54027_n1958;
  wire u5__abc_54027_n1959;
  wire u5__abc_54027_n1960;
  wire u5__abc_54027_n1961;
  wire u5__abc_54027_n1962;
  wire u5__abc_54027_n1963;
  wire u5__abc_54027_n1964;
  wire u5__abc_54027_n1965;
  wire u5__abc_54027_n1966;
  wire u5__abc_54027_n1967;
  wire u5__abc_54027_n1968;
  wire u5__abc_54027_n1969;
  wire u5__abc_54027_n1970;
  wire u5__abc_54027_n1971;
  wire u5__abc_54027_n1972;
  wire u5__abc_54027_n1973;
  wire u5__abc_54027_n1974;
  wire u5__abc_54027_n1975;
  wire u5__abc_54027_n1976;
  wire u5__abc_54027_n1977;
  wire u5__abc_54027_n1978;
  wire u5__abc_54027_n1979;
  wire u5__abc_54027_n1980;
  wire u5__abc_54027_n1981;
  wire u5__abc_54027_n1982;
  wire u5__abc_54027_n1983;
  wire u5__abc_54027_n1984;
  wire u5__abc_54027_n1985;
  wire u5__abc_54027_n1986;
  wire u5__abc_54027_n1988;
  wire u5__abc_54027_n1989;
  wire u5__abc_54027_n1990;
  wire u5__abc_54027_n1991;
  wire u5__abc_54027_n1992;
  wire u5__abc_54027_n1993;
  wire u5__abc_54027_n1994;
  wire u5__abc_54027_n1995;
  wire u5__abc_54027_n1997;
  wire u5__abc_54027_n2000;
  wire u5__abc_54027_n2001;
  wire u5__abc_54027_n2002;
  wire u5__abc_54027_n2004;
  wire u5__abc_54027_n2006;
  wire u5__abc_54027_n2009;
  wire u5__abc_54027_n2010;
  wire u5__abc_54027_n2012;
  wire u5__abc_54027_n2013;
  wire u5__abc_54027_n2014;
  wire u5__abc_54027_n2016;
  wire u5__abc_54027_n2017;
  wire u5__abc_54027_n2018;
  wire u5__abc_54027_n2019;
  wire u5__abc_54027_n2020;
  wire u5__abc_54027_n2021;
  wire u5__abc_54027_n248_1;
  wire u5__abc_54027_n249_1;
  wire u5__abc_54027_n250;
  wire u5__abc_54027_n251;
  wire u5__abc_54027_n252_1;
  wire u5__abc_54027_n253_1;
  wire u5__abc_54027_n254;
  wire u5__abc_54027_n255_1;
  wire u5__abc_54027_n256_1;
  wire u5__abc_54027_n257;
  wire u5__abc_54027_n258;
  wire u5__abc_54027_n259_1;
  wire u5__abc_54027_n260_1;
  wire u5__abc_54027_n261;
  wire u5__abc_54027_n262;
  wire u5__abc_54027_n263;
  wire u5__abc_54027_n264_1;
  wire u5__abc_54027_n265;
  wire u5__abc_54027_n267;
  wire u5__abc_54027_n268_1;
  wire u5__abc_54027_n269;
  wire u5__abc_54027_n270;
  wire u5__abc_54027_n271;
  wire u5__abc_54027_n272;
  wire u5__abc_54027_n273;
  wire u5__abc_54027_n274;
  wire u5__abc_54027_n276;
  wire u5__abc_54027_n277;
  wire u5__abc_54027_n278;
  wire u5__abc_54027_n279;
  wire u5__abc_54027_n280;
  wire u5__abc_54027_n281;
  wire u5__abc_54027_n282;
  wire u5__abc_54027_n283;
  wire u5__abc_54027_n285_1;
  wire u5__abc_54027_n286;
  wire u5__abc_54027_n287;
  wire u5__abc_54027_n288_1;
  wire u5__abc_54027_n289;
  wire u5__abc_54027_n290_1;
  wire u5__abc_54027_n291;
  wire u5__abc_54027_n292;
  wire u5__abc_54027_n293;
  wire u5__abc_54027_n294;
  wire u5__abc_54027_n295;
  wire u5__abc_54027_n296;
  wire u5__abc_54027_n297;
  wire u5__abc_54027_n298_1;
  wire u5__abc_54027_n299_1;
  wire u5__abc_54027_n300_1;
  wire u5__abc_54027_n301_1;
  wire u5__abc_54027_n302;
  wire u5__abc_54027_n303;
  wire u5__abc_54027_n304;
  wire u5__abc_54027_n305;
  wire u5__abc_54027_n306;
  wire u5__abc_54027_n307;
  wire u5__abc_54027_n308;
  wire u5__abc_54027_n309;
  wire u5__abc_54027_n311_1;
  wire u5__abc_54027_n312_1;
  wire u5__abc_54027_n313_1;
  wire u5__abc_54027_n314;
  wire u5__abc_54027_n315;
  wire u5__abc_54027_n316_1;
  wire u5__abc_54027_n317;
  wire u5__abc_54027_n318;
  wire u5__abc_54027_n319;
  wire u5__abc_54027_n320;
  wire u5__abc_54027_n321_1;
  wire u5__abc_54027_n322_1;
  wire u5__abc_54027_n325;
  wire u5__abc_54027_n326;
  wire u5__abc_54027_n327;
  wire u5__abc_54027_n328_1;
  wire u5__abc_54027_n329;
  wire u5__abc_54027_n330_1;
  wire u5__abc_54027_n331;
  wire u5__abc_54027_n332;
  wire u5__abc_54027_n333_1;
  wire u5__abc_54027_n334;
  wire u5__abc_54027_n336;
  wire u5__abc_54027_n337;
  wire u5__abc_54027_n338;
  wire u5__abc_54027_n339;
  wire u5__abc_54027_n340;
  wire u5__abc_54027_n341;
  wire u5__abc_54027_n343;
  wire u5__abc_54027_n344_1;
  wire u5__abc_54027_n345;
  wire u5__abc_54027_n346;
  wire u5__abc_54027_n347;
  wire u5__abc_54027_n348;
  wire u5__abc_54027_n349;
  wire u5__abc_54027_n350;
  wire u5__abc_54027_n351;
  wire u5__abc_54027_n351_bF_buf0;
  wire u5__abc_54027_n351_bF_buf1;
  wire u5__abc_54027_n351_bF_buf2;
  wire u5__abc_54027_n351_bF_buf3;
  wire u5__abc_54027_n352;
  wire u5__abc_54027_n353;
  wire u5__abc_54027_n354;
  wire u5__abc_54027_n355;
  wire u5__abc_54027_n356;
  wire u5__abc_54027_n357;
  wire u5__abc_54027_n359;
  wire u5__abc_54027_n360;
  wire u5__abc_54027_n361;
  wire u5__abc_54027_n362;
  wire u5__abc_54027_n363;
  wire u5__abc_54027_n364;
  wire u5__abc_54027_n365_1;
  wire u5__abc_54027_n366_1;
  wire u5__abc_54027_n367_1;
  wire u5__abc_54027_n368;
  wire u5__abc_54027_n369;
  wire u5__abc_54027_n370;
  wire u5__abc_54027_n371;
  wire u5__abc_54027_n372;
  wire u5__abc_54027_n373;
  wire u5__abc_54027_n374;
  wire u5__abc_54027_n375;
  wire u5__abc_54027_n376;
  wire u5__abc_54027_n377;
  wire u5__abc_54027_n378;
  wire u5__abc_54027_n379;
  wire u5__abc_54027_n380;
  wire u5__abc_54027_n381;
  wire u5__abc_54027_n382;
  wire u5__abc_54027_n383;
  wire u5__abc_54027_n384;
  wire u5__abc_54027_n385;
  wire u5__abc_54027_n386_1;
  wire u5__abc_54027_n387_1;
  wire u5__abc_54027_n388_1;
  wire u5__abc_54027_n389_1;
  wire u5__abc_54027_n390_1;
  wire u5__abc_54027_n391;
  wire u5__abc_54027_n392;
  wire u5__abc_54027_n393;
  wire u5__abc_54027_n394_1;
  wire u5__abc_54027_n395;
  wire u5__abc_54027_n396;
  wire u5__abc_54027_n397;
  wire u5__abc_54027_n398;
  wire u5__abc_54027_n399;
  wire u5__abc_54027_n400;
  wire u5__abc_54027_n401;
  wire u5__abc_54027_n402;
  wire u5__abc_54027_n403;
  wire u5__abc_54027_n404;
  wire u5__abc_54027_n405;
  wire u5__abc_54027_n406;
  wire u5__abc_54027_n407;
  wire u5__abc_54027_n408;
  wire u5__abc_54027_n409;
  wire u5__abc_54027_n410;
  wire u5__abc_54027_n411;
  wire u5__abc_54027_n412;
  wire u5__abc_54027_n413;
  wire u5__abc_54027_n414;
  wire u5__abc_54027_n415;
  wire u5__abc_54027_n416;
  wire u5__abc_54027_n417;
  wire u5__abc_54027_n418;
  wire u5__abc_54027_n419;
  wire u5__abc_54027_n420;
  wire u5__abc_54027_n421;
  wire u5__abc_54027_n422;
  wire u5__abc_54027_n423;
  wire u5__abc_54027_n424;
  wire u5__abc_54027_n425;
  wire u5__abc_54027_n426;
  wire u5__abc_54027_n427;
  wire u5__abc_54027_n428;
  wire u5__abc_54027_n429_1;
  wire u5__abc_54027_n430_1;
  wire u5__abc_54027_n431;
  wire u5__abc_54027_n432_1;
  wire u5__abc_54027_n433_1;
  wire u5__abc_54027_n434;
  wire u5__abc_54027_n435;
  wire u5__abc_54027_n436;
  wire u5__abc_54027_n437_1;
  wire u5__abc_54027_n438_1;
  wire u5__abc_54027_n439;
  wire u5__abc_54027_n440;
  wire u5__abc_54027_n441;
  wire u5__abc_54027_n442;
  wire u5__abc_54027_n443;
  wire u5__abc_54027_n444;
  wire u5__abc_54027_n445;
  wire u5__abc_54027_n446_1;
  wire u5__abc_54027_n447_1;
  wire u5__abc_54027_n448;
  wire u5__abc_54027_n449_1;
  wire u5__abc_54027_n450;
  wire u5__abc_54027_n451_1;
  wire u5__abc_54027_n452_1;
  wire u5__abc_54027_n453;
  wire u5__abc_54027_n454;
  wire u5__abc_54027_n455;
  wire u5__abc_54027_n456;
  wire u5__abc_54027_n457;
  wire u5__abc_54027_n458;
  wire u5__abc_54027_n459;
  wire u5__abc_54027_n460;
  wire u5__abc_54027_n461_1;
  wire u5__abc_54027_n462;
  wire u5__abc_54027_n463_1;
  wire u5__abc_54027_n464;
  wire u5__abc_54027_n465;
  wire u5__abc_54027_n466;
  wire u5__abc_54027_n467;
  wire u5__abc_54027_n468_1;
  wire u5__abc_54027_n469;
  wire u5__abc_54027_n470_1;
  wire u5__abc_54027_n471;
  wire u5__abc_54027_n472;
  wire u5__abc_54027_n473;
  wire u5__abc_54027_n474;
  wire u5__abc_54027_n475_1;
  wire u5__abc_54027_n476;
  wire u5__abc_54027_n477;
  wire u5__abc_54027_n478_1;
  wire u5__abc_54027_n479;
  wire u5__abc_54027_n480;
  wire u5__abc_54027_n481;
  wire u5__abc_54027_n482;
  wire u5__abc_54027_n483;
  wire u5__abc_54027_n484_1;
  wire u5__abc_54027_n485;
  wire u5__abc_54027_n486_1;
  wire u5__abc_54027_n487;
  wire u5__abc_54027_n488;
  wire u5__abc_54027_n489;
  wire u5__abc_54027_n490;
  wire u5__abc_54027_n491;
  wire u5__abc_54027_n492;
  wire u5__abc_54027_n493_1;
  wire u5__abc_54027_n494;
  wire u5__abc_54027_n495_1;
  wire u5__abc_54027_n496;
  wire u5__abc_54027_n497;
  wire u5__abc_54027_n498;
  wire u5__abc_54027_n499;
  wire u5__abc_54027_n500;
  wire u5__abc_54027_n501;
  wire u5__abc_54027_n503;
  wire u5__abc_54027_n504_1;
  wire u5__abc_54027_n505_1;
  wire u5__abc_54027_n506;
  wire u5__abc_54027_n507;
  wire u5__abc_54027_n508;
  wire u5__abc_54027_n509;
  wire u5__abc_54027_n510;
  wire u5__abc_54027_n511;
  wire u5__abc_54027_n512_1;
  wire u5__abc_54027_n513_1;
  wire u5__abc_54027_n514;
  wire u5__abc_54027_n515;
  wire u5__abc_54027_n516;
  wire u5__abc_54027_n517;
  wire u5__abc_54027_n518;
  wire u5__abc_54027_n519;
  wire u5__abc_54027_n520;
  wire u5__abc_54027_n521;
  wire u5__abc_54027_n522;
  wire u5__abc_54027_n523_1;
  wire u5__abc_54027_n524_1;
  wire u5__abc_54027_n525;
  wire u5__abc_54027_n526;
  wire u5__abc_54027_n527;
  wire u5__abc_54027_n528;
  wire u5__abc_54027_n529;
  wire u5__abc_54027_n530;
  wire u5__abc_54027_n532_1;
  wire u5__abc_54027_n533;
  wire u5__abc_54027_n534;
  wire u5__abc_54027_n536;
  wire u5__abc_54027_n537;
  wire u5__abc_54027_n538;
  wire u5__abc_54027_n539;
  wire u5__abc_54027_n541;
  wire u5__abc_54027_n542;
  wire u5__abc_54027_n544_1;
  wire u5__abc_54027_n545_1;
  wire u5__abc_54027_n546;
  wire u5__abc_54027_n547;
  wire u5__abc_54027_n548;
  wire u5__abc_54027_n549;
  wire u5__abc_54027_n550;
  wire u5__abc_54027_n551;
  wire u5__abc_54027_n553_1;
  wire u5__abc_54027_n554;
  wire u5__abc_54027_n556;
  wire u5__abc_54027_n557;
  wire u5__abc_54027_n558;
  wire u5__abc_54027_n559;
  wire u5__abc_54027_n560;
  wire u5__abc_54027_n561;
  wire u5__abc_54027_n562;
  wire u5__abc_54027_n563_1;
  wire u5__abc_54027_n564;
  wire u5__abc_54027_n565;
  wire u5__abc_54027_n565_bF_buf0;
  wire u5__abc_54027_n565_bF_buf1;
  wire u5__abc_54027_n565_bF_buf2;
  wire u5__abc_54027_n565_bF_buf3;
  wire u5__abc_54027_n565_bF_buf4;
  wire u5__abc_54027_n566_1;
  wire u5__abc_54027_n567;
  wire u5__abc_54027_n568;
  wire u5__abc_54027_n569_1;
  wire u5__abc_54027_n570;
  wire u5__abc_54027_n571;
  wire u5__abc_54027_n572_1;
  wire u5__abc_54027_n573;
  wire u5__abc_54027_n574;
  wire u5__abc_54027_n575;
  wire u5__abc_54027_n576;
  wire u5__abc_54027_n577_1;
  wire u5__abc_54027_n578;
  wire u5__abc_54027_n579_1;
  wire u5__abc_54027_n580;
  wire u5__abc_54027_n581;
  wire u5__abc_54027_n582;
  wire u5__abc_54027_n583;
  wire u5__abc_54027_n584;
  wire u5__abc_54027_n585;
  wire u5__abc_54027_n586;
  wire u5__abc_54027_n587;
  wire u5__abc_54027_n588;
  wire u5__abc_54027_n589;
  wire u5__abc_54027_n590;
  wire u5__abc_54027_n591;
  wire u5__abc_54027_n592_1;
  wire u5__abc_54027_n593;
  wire u5__abc_54027_n594;
  wire u5__abc_54027_n595;
  wire u5__abc_54027_n596;
  wire u5__abc_54027_n597;
  wire u5__abc_54027_n598;
  wire u5__abc_54027_n599;
  wire u5__abc_54027_n600;
  wire u5__abc_54027_n601_1;
  wire u5__abc_54027_n602;
  wire u5__abc_54027_n603;
  wire u5__abc_54027_n604;
  wire u5__abc_54027_n605_1;
  wire u5__abc_54027_n606;
  wire u5__abc_54027_n607;
  wire u5__abc_54027_n609;
  wire u5__abc_54027_n610;
  wire u5__abc_54027_n612;
  wire u5__abc_54027_n613;
  wire u5__abc_54027_n614;
  wire u5__abc_54027_n615;
  wire u5__abc_54027_n616;
  wire u5__abc_54027_n617;
  wire u5__abc_54027_n618;
  wire u5__abc_54027_n619;
  wire u5__abc_54027_n620_1;
  wire u5__abc_54027_n621;
  wire u5__abc_54027_n622;
  wire u5__abc_54027_n623;
  wire u5__abc_54027_n624;
  wire u5__abc_54027_n626;
  wire u5__abc_54027_n627;
  wire u5__abc_54027_n629;
  wire u5__abc_54027_n630_1;
  wire u5__abc_54027_n631;
  wire u5__abc_54027_n632_1;
  wire u5__abc_54027_n633;
  wire u5__abc_54027_n634;
  wire u5__abc_54027_n635;
  wire u5__abc_54027_n636;
  wire u5__abc_54027_n637;
  wire u5__abc_54027_n638_1;
  wire u5__abc_54027_n639;
  wire u5__abc_54027_n640;
  wire u5__abc_54027_n641;
  wire u5__abc_54027_n642;
  wire u5__abc_54027_n643_1;
  wire u5__abc_54027_n644;
  wire u5__abc_54027_n645;
  wire u5__abc_54027_n646;
  wire u5__abc_54027_n647;
  wire u5__abc_54027_n648;
  wire u5__abc_54027_n649;
  wire u5__abc_54027_n650;
  wire u5__abc_54027_n651;
  wire u5__abc_54027_n652;
  wire u5__abc_54027_n653;
  wire u5__abc_54027_n654_1;
  wire u5__abc_54027_n655;
  wire u5__abc_54027_n656;
  wire u5__abc_54027_n657_1;
  wire u5__abc_54027_n658;
  wire u5__abc_54027_n659;
  wire u5__abc_54027_n660;
  wire u5__abc_54027_n661;
  wire u5__abc_54027_n662;
  wire u5__abc_54027_n663;
  wire u5__abc_54027_n664;
  wire u5__abc_54027_n665;
  wire u5__abc_54027_n666_1;
  wire u5__abc_54027_n667;
  wire u5__abc_54027_n668;
  wire u5__abc_54027_n669;
  wire u5__abc_54027_n670;
  wire u5__abc_54027_n671;
  wire u5__abc_54027_n672_1;
  wire u5__abc_54027_n673;
  wire u5__abc_54027_n674;
  wire u5__abc_54027_n675;
  wire u5__abc_54027_n676;
  wire u5__abc_54027_n677;
  wire u5__abc_54027_n678;
  wire u5__abc_54027_n679;
  wire u5__abc_54027_n680;
  wire u5__abc_54027_n681_1;
  wire u5__abc_54027_n682;
  wire u5__abc_54027_n683;
  wire u5__abc_54027_n684;
  wire u5__abc_54027_n685_1;
  wire u5__abc_54027_n686;
  wire u5__abc_54027_n687_1;
  wire u5__abc_54027_n688;
  wire u5__abc_54027_n689;
  wire u5__abc_54027_n691;
  wire u5__abc_54027_n692;
  wire u5__abc_54027_n694_1;
  wire u5__abc_54027_n695;
  wire u5__abc_54027_n696;
  wire u5__abc_54027_n698;
  wire u5__abc_54027_n699_1;
  wire u5__abc_54027_n700;
  wire u5__abc_54027_n701;
  wire u5__abc_54027_n702;
  wire u5__abc_54027_n703;
  wire u5__abc_54027_n704;
  wire u5__abc_54027_n705_1;
  wire u5__abc_54027_n706;
  wire u5__abc_54027_n707;
  wire u5__abc_54027_n708;
  wire u5__abc_54027_n709_1;
  wire u5__abc_54027_n710;
  wire u5__abc_54027_n711;
  wire u5__abc_54027_n712;
  wire u5__abc_54027_n713_1;
  wire u5__abc_54027_n715;
  wire u5__abc_54027_n716;
  wire u5__abc_54027_n717;
  wire u5__abc_54027_n718;
  wire u5__abc_54027_n719;
  wire u5__abc_54027_n720;
  wire u5__abc_54027_n721;
  wire u5__abc_54027_n722;
  wire u5__abc_54027_n723;
  wire u5__abc_54027_n724;
  wire u5__abc_54027_n725;
  wire u5__abc_54027_n726;
  wire u5__abc_54027_n728;
  wire u5__abc_54027_n729_1;
  wire u5__abc_54027_n730;
  wire u5__abc_54027_n731;
  wire u5__abc_54027_n732;
  wire u5__abc_54027_n733;
  wire u5__abc_54027_n734;
  wire u5__abc_54027_n735;
  wire u5__abc_54027_n736;
  wire u5__abc_54027_n737_1;
  wire u5__abc_54027_n738;
  wire u5__abc_54027_n739;
  wire u5__abc_54027_n741;
  wire u5__abc_54027_n742;
  wire u5__abc_54027_n743;
  wire u5__abc_54027_n744_1;
  wire u5__abc_54027_n745;
  wire u5__abc_54027_n746;
  wire u5__abc_54027_n747_1;
  wire u5__abc_54027_n748;
  wire u5__abc_54027_n749;
  wire u5__abc_54027_n750;
  wire u5__abc_54027_n752_1;
  wire u5__abc_54027_n753;
  wire u5__abc_54027_n754;
  wire u5__abc_54027_n755_1;
  wire u5__abc_54027_n756;
  wire u5__abc_54027_n757;
  wire u5__abc_54027_n758;
  wire u5__abc_54027_n759_1;
  wire u5__abc_54027_n761;
  wire u5__abc_54027_n762_1;
  wire u5__abc_54027_n763_1;
  wire u5__abc_54027_n764;
  wire u5__abc_54027_n765;
  wire u5__abc_54027_n766_1;
  wire u5__abc_54027_n767_1;
  wire u5__abc_54027_n768;
  wire u5__abc_54027_n770;
  wire u5__abc_54027_n771_1;
  wire u5__abc_54027_n772_1;
  wire u5__abc_54027_n773;
  wire u5__abc_54027_n774;
  wire u5__abc_54027_n775;
  wire u5__abc_54027_n776;
  wire u5__abc_54027_n777;
  wire u5__abc_54027_n779;
  wire u5__abc_54027_n780;
  wire u5__abc_54027_n781;
  wire u5__abc_54027_n782;
  wire u5__abc_54027_n783;
  wire u5__abc_54027_n784;
  wire u5__abc_54027_n785;
  wire u5__abc_54027_n786;
  wire u5__abc_54027_n788;
  wire u5__abc_54027_n789;
  wire u5__abc_54027_n790;
  wire u5__abc_54027_n791_1;
  wire u5__abc_54027_n792;
  wire u5__abc_54027_n793;
  wire u5__abc_54027_n794;
  wire u5__abc_54027_n795;
  wire u5__abc_54027_n796;
  wire u5__abc_54027_n797;
  wire u5__abc_54027_n799;
  wire u5__abc_54027_n800;
  wire u5__abc_54027_n801_1;
  wire u5__abc_54027_n802;
  wire u5__abc_54027_n803;
  wire u5__abc_54027_n804;
  wire u5__abc_54027_n805;
  wire u5__abc_54027_n806;
  wire u5__abc_54027_n807;
  wire u5__abc_54027_n808;
  wire u5__abc_54027_n809;
  wire u5__abc_54027_n810_1;
  wire u5__abc_54027_n812;
  wire u5__abc_54027_n813;
  wire u5__abc_54027_n814;
  wire u5__abc_54027_n815;
  wire u5__abc_54027_n816;
  wire u5__abc_54027_n817;
  wire u5__abc_54027_n818;
  wire u5__abc_54027_n819;
  wire u5__abc_54027_n820;
  wire u5__abc_54027_n821_1;
  wire u5__abc_54027_n822;
  wire u5__abc_54027_n823;
  wire u5__abc_54027_n825;
  wire u5__abc_54027_n826;
  wire u5__abc_54027_n827;
  wire u5__abc_54027_n828;
  wire u5__abc_54027_n829;
  wire u5__abc_54027_n831;
  wire u5__abc_54027_n832;
  wire u5__abc_54027_n833_1;
  wire u5__abc_54027_n834;
  wire u5__abc_54027_n836;
  wire u5__abc_54027_n837;
  wire u5__abc_54027_n838;
  wire u5__abc_54027_n839;
  wire u5__abc_54027_n841;
  wire u5__abc_54027_n842;
  wire u5__abc_54027_n843_1;
  wire u5__abc_54027_n844;
  wire u5__abc_54027_n846;
  wire u5__abc_54027_n847;
  wire u5__abc_54027_n848;
  wire u5__abc_54027_n849;
  wire u5__abc_54027_n850;
  wire u5__abc_54027_n851;
  wire u5__abc_54027_n852;
  wire u5__abc_54027_n853;
  wire u5__abc_54027_n854;
  wire u5__abc_54027_n855_1;
  wire u5__abc_54027_n856;
  wire u5__abc_54027_n857;
  wire u5__abc_54027_n858;
  wire u5__abc_54027_n859;
  wire u5__abc_54027_n860;
  wire u5__abc_54027_n861_1;
  wire u5__abc_54027_n862;
  wire u5__abc_54027_n863;
  wire u5__abc_54027_n864;
  wire u5__abc_54027_n865;
  wire u5__abc_54027_n866;
  wire u5__abc_54027_n867;
  wire u5__abc_54027_n868_1;
  wire u5__abc_54027_n869_1;
  wire u5__abc_54027_n870;
  wire u5__abc_54027_n871;
  wire u5__abc_54027_n872;
  wire u5__abc_54027_n873;
  wire u5__abc_54027_n874;
  wire u5__abc_54027_n875;
  wire u5__abc_54027_n876_1;
  wire u5__abc_54027_n877;
  wire u5__abc_54027_n878;
  wire u5__abc_54027_n879;
  wire u5__abc_54027_n880;
  wire u5__abc_54027_n881;
  wire u5__abc_54027_n882_1;
  wire u5__abc_54027_n883;
  wire u5__abc_54027_n884;
  wire u5__abc_54027_n885;
  wire u5__abc_54027_n886;
  wire u5__abc_54027_n887_1;
  wire u5__abc_54027_n888;
  wire u5__abc_54027_n889;
  wire u5__abc_54027_n890;
  wire u5__abc_54027_n891;
  wire u5__abc_54027_n892;
  wire u5__abc_54027_n893;
  wire u5__abc_54027_n894;
  wire u5__abc_54027_n895_1;
  wire u5__abc_54027_n896_1;
  wire u5__abc_54027_n897_1;
  wire u5__abc_54027_n898_1;
  wire u5__abc_54027_n899_1;
  wire u5__abc_54027_n900_1;
  wire u5__abc_54027_n901;
  wire u5__abc_54027_n902;
  wire u5__abc_54027_n903;
  wire u5__abc_54027_n904;
  wire u5__abc_54027_n905_1;
  wire u5__abc_54027_n906_1;
  wire u5__abc_54027_n907;
  wire u5__abc_54027_n908;
  wire u5__abc_54027_n909;
  wire u5__abc_54027_n910;
  wire u5__abc_54027_n911;
  wire u5__abc_54027_n912;
  wire u5__abc_54027_n913;
  wire u5__abc_54027_n915;
  wire u5__abc_54027_n916;
  wire u5__abc_54027_n917;
  wire u5__abc_54027_n918;
  wire u5__abc_54027_n919;
  wire u5__abc_54027_n920;
  wire u5__abc_54027_n921;
  wire u5__abc_54027_n922;
  wire u5__abc_54027_n923;
  wire u5__abc_54027_n924;
  wire u5__abc_54027_n925;
  wire u5__abc_54027_n926;
  wire u5__abc_54027_n927;
  wire u5__abc_54027_n928;
  wire u5__abc_54027_n929;
  wire u5__abc_54027_n930;
  wire u5__abc_54027_n931;
  wire u5__abc_54027_n932;
  wire u5__abc_54027_n933;
  wire u5__abc_54027_n934;
  wire u5__abc_54027_n935;
  wire u5__abc_54027_n936;
  wire u5__abc_54027_n937;
  wire u5__abc_54027_n938;
  wire u5__abc_54027_n939;
  wire u5__abc_54027_n940;
  wire u5__abc_54027_n941;
  wire u5__abc_54027_n942_1;
  wire u5__abc_54027_n943;
  wire u5__abc_54027_n944;
  wire u5__abc_54027_n945;
  wire u5__abc_54027_n946;
  wire u5__abc_54027_n947;
  wire u5__abc_54027_n948;
  wire u5__abc_54027_n949;
  wire u5__abc_54027_n950;
  wire u5__abc_54027_n951;
  wire u5__abc_54027_n952;
  wire u5__abc_54027_n953_1;
  wire u5__abc_54027_n954;
  wire u5__abc_54027_n955;
  wire u5__abc_54027_n956;
  wire u5__abc_54027_n957;
  wire u5__abc_54027_n958;
  wire u5__abc_54027_n959;
  wire u5__abc_54027_n960;
  wire u5__abc_54027_n961;
  wire u5__abc_54027_n962;
  wire u5__abc_54027_n963;
  wire u5__abc_54027_n964;
  wire u5__abc_54027_n966;
  wire u5__abc_54027_n967;
  wire u5__abc_54027_n968;
  wire u5__abc_54027_n969;
  wire u5__abc_54027_n970;
  wire u5__abc_54027_n971;
  wire u5__abc_54027_n972;
  wire u5__abc_54027_n973;
  wire u5__abc_54027_n974;
  wire u5__abc_54027_n975;
  wire u5__abc_54027_n976;
  wire u5__abc_54027_n977;
  wire u5__abc_54027_n978;
  wire u5__abc_54027_n979;
  wire u5__abc_54027_n980;
  wire u5__abc_54027_n981;
  wire u5__abc_54027_n982;
  wire u5__abc_54027_n983;
  wire u5__abc_54027_n984;
  wire u5__abc_54027_n985;
  wire u5__abc_54027_n986;
  wire u5__abc_54027_n987;
  wire u5__abc_54027_n988;
  wire u5__abc_54027_n989;
  wire u5__abc_54027_n990;
  wire u5__abc_54027_n991;
  wire u5__abc_54027_n992;
  wire u5__abc_54027_n993;
  wire u5__abc_54027_n994;
  wire u5__abc_54027_n995;
  wire u5__abc_54027_n996;
  wire u5__abc_54027_n997;
  wire u5__abc_54027_n998;
  wire u5__abc_54027_n999;
  wire u5_ack_cnt_0_;
  wire u5_ack_cnt_0__FF_INPUT;
  wire u5_ack_cnt_1_;
  wire u5_ack_cnt_1__FF_INPUT;
  wire u5_ack_cnt_2_;
  wire u5_ack_cnt_2__FF_INPUT;
  wire u5_ack_cnt_3_;
  wire u5_ack_cnt_3__FF_INPUT;
  wire u5_ap_en;
  wire u5_ap_en_FF_INPUT;
  wire u5_burst_act_rd;
  wire u5_burst_act_rd_FF_INPUT;
  wire u5_burst_cnt_0_;
  wire u5_burst_cnt_0__FF_INPUT;
  wire u5_burst_cnt_10_;
  wire u5_burst_cnt_10__FF_INPUT;
  wire u5_burst_cnt_1_;
  wire u5_burst_cnt_1__FF_INPUT;
  wire u5_burst_cnt_2_;
  wire u5_burst_cnt_2__FF_INPUT;
  wire u5_burst_cnt_3_;
  wire u5_burst_cnt_3__FF_INPUT;
  wire u5_burst_cnt_4_;
  wire u5_burst_cnt_4__FF_INPUT;
  wire u5_burst_cnt_5_;
  wire u5_burst_cnt_5__FF_INPUT;
  wire u5_burst_cnt_6_;
  wire u5_burst_cnt_6__FF_INPUT;
  wire u5_burst_cnt_7_;
  wire u5_burst_cnt_7__FF_INPUT;
  wire u5_burst_cnt_8_;
  wire u5_burst_cnt_8__FF_INPUT;
  wire u5_burst_cnt_9_;
  wire u5_burst_cnt_9__FF_INPUT;
  wire u5_cke__FF_INPUT;
  wire u5_cke_d;
  wire u5_cke_o_del;
  wire u5_cke_o_r1;
  wire u5_cke_o_r2;
  wire u5_cke_r;
  wire u5_cmd_0_;
  wire u5_cmd_1_;
  wire u5_cmd_2_;
  wire u5_cmd_3_;
  wire u5_cmd_a10_r;
  wire u5_cmd_asserted;
  wire u5_cmd_asserted2;
  wire u5_cmd_asserted2_FF_INPUT;
  wire u5_cmd_asserted_FF_INPUT;
  wire u5_cmd_asserted_bF_buf0;
  wire u5_cmd_asserted_bF_buf1;
  wire u5_cmd_asserted_bF_buf2;
  wire u5_cmd_asserted_bF_buf3;
  wire u5_cmd_del_0_;
  wire u5_cmd_del_1_;
  wire u5_cmd_del_2_;
  wire u5_cmd_del_3_;
  wire u5_cmd_r_0_;
  wire u5_cmd_r_1_;
  wire u5_cmd_r_2_;
  wire u5_cmd_r_3_;
  wire u5_cnt;
  wire u5_cnt_next;
  wire u5_cs_le_r;
  wire u5_cs_le_r1;
  wire u5_data_oe_FF_INPUT;
  wire u5_data_oe_d;
  wire u5_data_oe_r;
  wire u5_data_oe_r2;
  wire u5_dv_r;
  wire u5_ir_cnt_0_;
  wire u5_ir_cnt_0__FF_INPUT;
  wire u5_ir_cnt_1_;
  wire u5_ir_cnt_1__FF_INPUT;
  wire u5_ir_cnt_2_;
  wire u5_ir_cnt_2__FF_INPUT;
  wire u5_ir_cnt_3_;
  wire u5_ir_cnt_3__FF_INPUT;
  wire u5_ir_cnt_done;
  wire u5_ir_cnt_done_FF_INPUT;
  wire u5_kro;
  wire u5_lmr_ack_d;
  wire u5_lookup_ready1;
  wire u5_lookup_ready1_FF_INPUT;
  wire u5_lookup_ready2;
  wire u5_lookup_ready2_FF_INPUT;
  wire u5_mc_adv_r;
  wire u5_mc_adv_r1;
  wire u5_mc_adv_r1_FF_INPUT;
  wire u5_mc_adv_r_FF_INPUT;
  wire u5_mc_c_oe_d;
  wire u5_mc_le;
  wire u5_mc_le_FF_INPUT;
  wire u5_mem_ack_r;
  wire u5_no_wb_cycle;
  wire u5_no_wb_cycle_FF_INPUT;
  wire u5_oe__FF_INPUT;
  wire u5_pack_le0_d;
  wire u5_pack_le1_d;
  wire u5_pack_le2_d;
  wire u5_resume_req_r;
  wire u5_rfr_ack_d;
  wire u5_rsts;
  wire u5_rsts1;
  wire u5_state_0_;
  wire u5_state_1_;
  wire u5_state_2_;
  wire u5_state_3_;
  wire u5_state_4_;
  wire u5_state_5_;
  wire u5_state_6_;
  wire u5_susp_req_r;
  wire u5_susp_sel_r_FF_INPUT;
  wire u5_suspended_d;
  wire u5_timer2_0_;
  wire u5_timer2_0__FF_INPUT;
  wire u5_timer2_1_;
  wire u5_timer2_1__FF_INPUT;
  wire u5_timer2_2_;
  wire u5_timer2_2__FF_INPUT;
  wire u5_timer2_3_;
  wire u5_timer2_3__FF_INPUT;
  wire u5_timer2_4_;
  wire u5_timer2_4__FF_INPUT;
  wire u5_timer2_5_;
  wire u5_timer2_5__FF_INPUT;
  wire u5_timer2_6_;
  wire u5_timer2_6__FF_INPUT;
  wire u5_timer2_7_;
  wire u5_timer2_7__FF_INPUT;
  wire u5_timer2_8_;
  wire u5_timer2_8__FF_INPUT;
  wire u5_timer_0_;
  wire u5_timer_0__FF_INPUT;
  wire u5_timer_1_;
  wire u5_timer_1__FF_INPUT;
  wire u5_timer_2_;
  wire u5_timer_2__FF_INPUT;
  wire u5_timer_3_;
  wire u5_timer_3__FF_INPUT;
  wire u5_timer_4_;
  wire u5_timer_4__FF_INPUT;
  wire u5_timer_5_;
  wire u5_timer_5__FF_INPUT;
  wire u5_timer_6_;
  wire u5_timer_6__FF_INPUT;
  wire u5_timer_7_;
  wire u5_timer_7__FF_INPUT;
  wire u5_timer_is_zero;
  wire u5_tmr2_done;
  wire u5_tmr2_done_FF_INPUT;
  wire u5_tmr_done;
  wire u5_wb_cycle;
  wire u5_wb_cycle_FF_INPUT;
  wire u5_wb_first;
  wire u5_wb_stb_first;
  wire u5_wb_stb_first_FF_INPUT;
  wire u5_wb_wait;
  wire u5_wb_wait_r;
  wire u5_wb_wait_r2;
  wire u5_wb_write_go_r;
  wire u5_we_;
  wire u5_wr_cycle_FF_INPUT;
  wire u6__abc_56056_n132;
  wire u6__abc_56056_n133;
  wire u6__abc_56056_n134;
  wire u6__abc_56056_n135_1;
  wire u6__abc_56056_n136;
  wire u6__abc_56056_n137;
  wire u6__abc_56056_n138_1;
  wire u6__abc_56056_n139_1;
  wire u6__abc_56056_n140_1;
  wire u6__abc_56056_n141_1;
  wire u6__abc_56056_n142_1;
  wire u6__abc_56056_n143;
  wire u6__abc_56056_n144;
  wire u6__abc_56056_n144_bF_buf0;
  wire u6__abc_56056_n144_bF_buf1;
  wire u6__abc_56056_n144_bF_buf2;
  wire u6__abc_56056_n144_bF_buf3;
  wire u6__abc_56056_n144_bF_buf4;
  wire u6__abc_56056_n144_bF_buf5;
  wire u6__abc_56056_n145_1;
  wire u6__abc_56056_n146_1;
  wire u6__abc_56056_n147;
  wire u6__abc_56056_n148_1;
  wire u6__abc_56056_n149_1;
  wire u6__abc_56056_n150_1;
  wire u6__abc_56056_n151;
  wire u6__abc_56056_n153;
  wire u6__abc_56056_n154;
  wire u6__abc_56056_n154_bF_buf0;
  wire u6__abc_56056_n154_bF_buf1;
  wire u6__abc_56056_n154_bF_buf2;
  wire u6__abc_56056_n154_bF_buf3;
  wire u6__abc_56056_n154_bF_buf4;
  wire u6__abc_56056_n155_1;
  wire u6__abc_56056_n157_1;
  wire u6__abc_56056_n158;
  wire u6__abc_56056_n160;
  wire u6__abc_56056_n161;
  wire u6__abc_56056_n163_1;
  wire u6__abc_56056_n164;
  wire u6__abc_56056_n166_1;
  wire u6__abc_56056_n167;
  wire u6__abc_56056_n167_1;
  wire u6__abc_56056_n169;
  wire u6__abc_56056_n170;
  wire u6__abc_56056_n172;
  wire u6__abc_56056_n173;
  wire u6__abc_56056_n175;
  wire u6__abc_56056_n176;
  wire u6__abc_56056_n178;
  wire u6__abc_56056_n179;
  wire u6__abc_56056_n181;
  wire u6__abc_56056_n182;
  wire u6__abc_56056_n184;
  wire u6__abc_56056_n185;
  wire u6__abc_56056_n187;
  wire u6__abc_56056_n188;
  wire u6__abc_56056_n190;
  wire u6__abc_56056_n191;
  wire u6__abc_56056_n193;
  wire u6__abc_56056_n194;
  wire u6__abc_56056_n196;
  wire u6__abc_56056_n197;
  wire u6__abc_56056_n199;
  wire u6__abc_56056_n200;
  wire u6__abc_56056_n202;
  wire u6__abc_56056_n203;
  wire u6__abc_56056_n205;
  wire u6__abc_56056_n206;
  wire u6__abc_56056_n208;
  wire u6__abc_56056_n209;
  wire u6__abc_56056_n211;
  wire u6__abc_56056_n212;
  wire u6__abc_56056_n214;
  wire u6__abc_56056_n215;
  wire u6__abc_56056_n217;
  wire u6__abc_56056_n218;
  wire u6__abc_56056_n220;
  wire u6__abc_56056_n221;
  wire u6__abc_56056_n223;
  wire u6__abc_56056_n224;
  wire u6__abc_56056_n226;
  wire u6__abc_56056_n227;
  wire u6__abc_56056_n229;
  wire u6__abc_56056_n230;
  wire u6__abc_56056_n232;
  wire u6__abc_56056_n233;
  wire u6__abc_56056_n235;
  wire u6__abc_56056_n236;
  wire u6__abc_56056_n238;
  wire u6__abc_56056_n239;
  wire u6__abc_56056_n241;
  wire u6__abc_56056_n242;
  wire u6__abc_56056_n244;
  wire u6__abc_56056_n245;
  wire u6__abc_56056_n247;
  wire u6__abc_56056_n248;
  wire u6__abc_56056_n250;
  wire u6__abc_56056_n251;
  wire u6__abc_56056_n253;
  wire u6__abc_56056_n254;
  wire u6__abc_56056_n256;
  wire u6__abc_56056_n257;
  wire u6__abc_56056_n258;
  wire u6__abc_56056_n259;
  wire u6__abc_56056_n260;
  wire u6__abc_56056_n261;
  wire u6__abc_56056_n262;
  wire u6__abc_56056_n263;
  wire u6__abc_56056_n267;
  wire u6__abc_56056_n268;
  wire u6__abc_56056_n270;
  wire u6__abc_56056_n271;
  wire u6__abc_56056_n272;
  wire u6__abc_56056_n275;
  wire u6__abc_56056_n276;
  wire u6__abc_56056_n277;
  wire u6__abc_56056_n278;
  wire u6__abc_56056_n279;
  wire u6__abc_56056_n280;
  wire u6__abc_56056_n281;
  wire u6__abc_56056_n282;
  wire u6__abc_56056_n284;
  wire u6__abc_56056_n285;
  wire u6__abc_56056_n287;
  wire u6__abc_56056_n288;
  wire u6__abc_56056_n290;
  wire u6_read_go_r;
  wire u6_read_go_r1;
  wire u6_read_go_r1_FF_INPUT;
  wire u6_read_go_r_FF_INPUT;
  wire u6_rmw_en;
  wire u6_rmw_en_FF_INPUT;
  wire u6_rmw_r;
  wire u6_rmw_r_FF_INPUT;
  wire u6_wb_ack_o_FF_INPUT;
  wire u6_wb_data_o_0__FF_INPUT;
  wire u6_wb_data_o_10__FF_INPUT;
  wire u6_wb_data_o_11__FF_INPUT;
  wire u6_wb_data_o_12__FF_INPUT;
  wire u6_wb_data_o_13__FF_INPUT;
  wire u6_wb_data_o_14__FF_INPUT;
  wire u6_wb_data_o_15__FF_INPUT;
  wire u6_wb_data_o_16__FF_INPUT;
  wire u6_wb_data_o_17__FF_INPUT;
  wire u6_wb_data_o_18__FF_INPUT;
  wire u6_wb_data_o_19__FF_INPUT;
  wire u6_wb_data_o_1__FF_INPUT;
  wire u6_wb_data_o_20__FF_INPUT;
  wire u6_wb_data_o_21__FF_INPUT;
  wire u6_wb_data_o_22__FF_INPUT;
  wire u6_wb_data_o_23__FF_INPUT;
  wire u6_wb_data_o_24__FF_INPUT;
  wire u6_wb_data_o_25__FF_INPUT;
  wire u6_wb_data_o_26__FF_INPUT;
  wire u6_wb_data_o_27__FF_INPUT;
  wire u6_wb_data_o_28__FF_INPUT;
  wire u6_wb_data_o_29__FF_INPUT;
  wire u6_wb_data_o_2__FF_INPUT;
  wire u6_wb_data_o_30__FF_INPUT;
  wire u6_wb_data_o_31__FF_INPUT;
  wire u6_wb_data_o_3__FF_INPUT;
  wire u6_wb_data_o_4__FF_INPUT;
  wire u6_wb_data_o_5__FF_INPUT;
  wire u6_wb_data_o_6__FF_INPUT;
  wire u6_wb_data_o_7__FF_INPUT;
  wire u6_wb_data_o_8__FF_INPUT;
  wire u6_wb_data_o_9__FF_INPUT;
  wire u6_wb_err_FF_INPUT;
  wire u6_wb_first_r;
  wire u6_wr_hold_FF_INPUT;
  wire u6_write_go_r;
  wire u6_write_go_r1;
  wire u6_write_go_r1_FF_INPUT;
  wire u6_write_go_r_FF_INPUT;
  wire u7__abc_47535_n100;
  wire u7__abc_47535_n101;
  wire u7__abc_47535_n103;
  wire u7__abc_47535_n104;
  wire u7__abc_47535_n106;
  wire u7__abc_47535_n107;
  wire u7__abc_47535_n108;
  wire u7__abc_47535_n109;
  wire u7__abc_47535_n110;
  wire u7__abc_47535_n111;
  wire u7__abc_47535_n112;
  wire u7__abc_47535_n113;
  wire u7__abc_47535_n114;
  wire u7__abc_47535_n115;
  wire u7__abc_47535_n116;
  wire u7__abc_47535_n117;
  wire u7__abc_47535_n119;
  wire u7__abc_47535_n120;
  wire u7__abc_47535_n121;
  wire u7__abc_47535_n122;
  wire u7__abc_47535_n123;
  wire u7__abc_47535_n124;
  wire u7__abc_47535_n125;
  wire u7__abc_47535_n126;
  wire u7__abc_47535_n127;
  wire u7__abc_47535_n129;
  wire u7__abc_47535_n130;
  wire u7__abc_47535_n131;
  wire u7__abc_47535_n132;
  wire u7__abc_47535_n133;
  wire u7__abc_47535_n134;
  wire u7__abc_47535_n135;
  wire u7__abc_47535_n136;
  wire u7__abc_47535_n137;
  wire u7__abc_47535_n139;
  wire u7__abc_47535_n140;
  wire u7__abc_47535_n141;
  wire u7__abc_47535_n142;
  wire u7__abc_47535_n143;
  wire u7__abc_47535_n144;
  wire u7__abc_47535_n145;
  wire u7__abc_47535_n146;
  wire u7__abc_47535_n147;
  wire u7__abc_47535_n149;
  wire u7__abc_47535_n150;
  wire u7__abc_47535_n151;
  wire u7__abc_47535_n152;
  wire u7__abc_47535_n153;
  wire u7__abc_47535_n154;
  wire u7__abc_47535_n155;
  wire u7__abc_47535_n156;
  wire u7__abc_47535_n157;
  wire u7__abc_47535_n159;
  wire u7__abc_47535_n160;
  wire u7__abc_47535_n161;
  wire u7__abc_47535_n162;
  wire u7__abc_47535_n163;
  wire u7__abc_47535_n164;
  wire u7__abc_47535_n165;
  wire u7__abc_47535_n166;
  wire u7__abc_47535_n167;
  wire u7__abc_47535_n169;
  wire u7__abc_47535_n170;
  wire u7__abc_47535_n171;
  wire u7__abc_47535_n172;
  wire u7__abc_47535_n173;
  wire u7__abc_47535_n174;
  wire u7__abc_47535_n175;
  wire u7__abc_47535_n176;
  wire u7__abc_47535_n177;
  wire u7__abc_47535_n179;
  wire u7__abc_47535_n180;
  wire u7__abc_47535_n181;
  wire u7__abc_47535_n182;
  wire u7__abc_47535_n183;
  wire u7__abc_47535_n184;
  wire u7__abc_47535_n185;
  wire u7__abc_47535_n186;
  wire u7__abc_47535_n187;
  wire u7__abc_47535_n191;
  wire u7__abc_47535_n192;
  wire u7__abc_47535_n194;
  wire u7__abc_47535_n195;
  wire u7__abc_47535_n75_1;
  wire u7__abc_47535_n76;
  wire u7__abc_47535_n77_1;
  wire u7__abc_47535_n78;
  wire u7__abc_47535_n79_1;
  wire u7__abc_47535_n80_1;
  wire u7__abc_47535_n81_1;
  wire u7__abc_47535_n83_1;
  wire u7__abc_47535_n84;
  wire u7__abc_47535_n86_1;
  wire u7__abc_47535_n87_1;
  wire u7__abc_47535_n89_1;
  wire u7__abc_47535_n90_1;
  wire u7__abc_47535_n92_1;
  wire u7__abc_47535_n93;
  wire u7__abc_47535_n94_1;
  wire u7__abc_47535_n95_1;
  wire u7__abc_47535_n97_1;
  wire u7__abc_47535_n98_1;
  wire u7__abc_47535_n99;
  wire u7_mc_adsc__FF_INPUT;
  wire u7_mc_adv__FF_INPUT;
  wire u7_mc_cs__FF_INPUT;
  wire u7_mc_data_oe_FF_INPUT;
  wire u7_mc_dqm_0__FF_INPUT;
  wire u7_mc_dqm_1__FF_INPUT;
  wire u7_mc_dqm_2__FF_INPUT;
  wire u7_mc_dqm_3__FF_INPUT;
  wire u7_mc_dqm_r2_0_;
  wire u7_mc_dqm_r2_1_;
  wire u7_mc_dqm_r2_2_;
  wire u7_mc_dqm_r2_3_;
  wire u7_mc_dqm_r_0_;
  wire u7_mc_dqm_r_0__FF_INPUT;
  wire u7_mc_dqm_r_1_;
  wire u7_mc_dqm_r_1__FF_INPUT;
  wire u7_mc_dqm_r_2_;
  wire u7_mc_dqm_r_2__FF_INPUT;
  wire u7_mc_dqm_r_3_;
  wire u7_mc_dqm_r_3__FF_INPUT;
  wire u7_mc_oe__FF_INPUT;
  wire u7_mc_rp_FF_INPUT;
  output wb_ack_o;
  input \wb_addr_i[0] ;
  input \wb_addr_i[10] ;
  input \wb_addr_i[11] ;
  input \wb_addr_i[12] ;
  input \wb_addr_i[13] ;
  input \wb_addr_i[14] ;
  input \wb_addr_i[15] ;
  input \wb_addr_i[16] ;
  input \wb_addr_i[17] ;
  input \wb_addr_i[18] ;
  input \wb_addr_i[19] ;
  input \wb_addr_i[1] ;
  input \wb_addr_i[20] ;
  input \wb_addr_i[21] ;
  input \wb_addr_i[22] ;
  input \wb_addr_i[23] ;
  input \wb_addr_i[24] ;
  input \wb_addr_i[25] ;
  input \wb_addr_i[26] ;
  input \wb_addr_i[27] ;
  input \wb_addr_i[28] ;
  input \wb_addr_i[29] ;
  input \wb_addr_i[2] ;
  input \wb_addr_i[30] ;
  input \wb_addr_i[31] ;
  input \wb_addr_i[3] ;
  input \wb_addr_i[4] ;
  input \wb_addr_i[5] ;
  input \wb_addr_i[6] ;
  input \wb_addr_i[7] ;
  input \wb_addr_i[8] ;
  input \wb_addr_i[9] ;
  wire wb_addr_i_23_bF_buf0;
  wire wb_addr_i_23_bF_buf1;
  wire wb_addr_i_23_bF_buf2;
  wire wb_addr_i_23_bF_buf3;
  wire wb_addr_i_25_bF_buf0;
  wire wb_addr_i_25_bF_buf1;
  wire wb_addr_i_25_bF_buf2;
  wire wb_addr_i_25_bF_buf3;
  input wb_cyc_i;
  input \wb_data_i[0] ;
  input \wb_data_i[10] ;
  input \wb_data_i[11] ;
  input \wb_data_i[12] ;
  input \wb_data_i[13] ;
  input \wb_data_i[14] ;
  input \wb_data_i[15] ;
  input \wb_data_i[16] ;
  input \wb_data_i[17] ;
  input \wb_data_i[18] ;
  input \wb_data_i[19] ;
  input \wb_data_i[1] ;
  input \wb_data_i[20] ;
  input \wb_data_i[21] ;
  input \wb_data_i[22] ;
  input \wb_data_i[23] ;
  input \wb_data_i[24] ;
  input \wb_data_i[25] ;
  input \wb_data_i[26] ;
  input \wb_data_i[27] ;
  input \wb_data_i[28] ;
  input \wb_data_i[29] ;
  input \wb_data_i[2] ;
  input \wb_data_i[30] ;
  input \wb_data_i[31] ;
  input \wb_data_i[3] ;
  input \wb_data_i[4] ;
  input \wb_data_i[5] ;
  input \wb_data_i[6] ;
  input \wb_data_i[7] ;
  input \wb_data_i[8] ;
  input \wb_data_i[9] ;
  output \wb_data_o[0] ;
  output \wb_data_o[10] ;
  output \wb_data_o[11] ;
  output \wb_data_o[12] ;
  output \wb_data_o[13] ;
  output \wb_data_o[14] ;
  output \wb_data_o[15] ;
  output \wb_data_o[16] ;
  output \wb_data_o[17] ;
  output \wb_data_o[18] ;
  output \wb_data_o[19] ;
  output \wb_data_o[1] ;
  output \wb_data_o[20] ;
  output \wb_data_o[21] ;
  output \wb_data_o[22] ;
  output \wb_data_o[23] ;
  output \wb_data_o[24] ;
  output \wb_data_o[25] ;
  output \wb_data_o[26] ;
  output \wb_data_o[27] ;
  output \wb_data_o[28] ;
  output \wb_data_o[29] ;
  output \wb_data_o[2] ;
  output \wb_data_o[30] ;
  output \wb_data_o[31] ;
  output \wb_data_o[3] ;
  output \wb_data_o[4] ;
  output \wb_data_o[5] ;
  output \wb_data_o[6] ;
  output \wb_data_o[7] ;
  output \wb_data_o[8] ;
  output \wb_data_o[9] ;
  output wb_err_o;
  input \wb_sel_i[0] ;
  input \wb_sel_i[1] ;
  input \wb_sel_i[2] ;
  input \wb_sel_i[3] ;
  input wb_stb_i;
  wire wb_stb_i_bF_buf0;
  wire wb_stb_i_bF_buf1;
  wire wb_stb_i_bF_buf2;
  wire wb_stb_i_bF_buf3;
  wire wb_stb_i_bF_buf4;
  wire wb_stb_i_bF_buf5;
  input wb_we_i;
  AND2X2 AND2X2_1 ( .A(_abc_55805_n238_1), .B(_abc_55805_n239_1), .Y(_abc_55805_n240) );
  AND2X2 AND2X2_10 ( .A(_abc_55805_n266), .B(_abc_55805_n267), .Y(_abc_55805_n268) );
  AND2X2 AND2X2_100 ( .A(u0__abc_49347_n1168_1), .B(u0__abc_49347_n1154_1), .Y(u0__abc_49347_n1169) );
  AND2X2 AND2X2_1000 ( .A(u0__abc_49347_n1175_bF_buf0), .B(u0__abc_49347_n3373), .Y(u0__abc_49347_n3374) );
  AND2X2 AND2X2_1001 ( .A(u0__abc_49347_n3372), .B(u0__abc_49347_n3374), .Y(u0__abc_49347_n3375) );
  AND2X2 AND2X2_1002 ( .A(u0__abc_49347_n1176_1_bF_buf0), .B(tms_27_), .Y(u0__abc_49347_n3377) );
  AND2X2 AND2X2_1003 ( .A(u0_tms5_27_), .B(u0_cs5_bF_buf1), .Y(u0__abc_49347_n3378) );
  AND2X2 AND2X2_1004 ( .A(u0__abc_49347_n3380), .B(u0__abc_49347_n2730_bF_buf2), .Y(u0__abc_49347_n3381) );
  AND2X2 AND2X2_1005 ( .A(u0__abc_49347_n3381), .B(u0__abc_49347_n3379), .Y(u0__abc_49347_n3382) );
  AND2X2 AND2X2_1006 ( .A(u0__abc_49347_n3383), .B(u0__abc_49347_n2726_bF_buf2), .Y(u0__abc_49347_n3384) );
  AND2X2 AND2X2_1007 ( .A(u0_tms4_27_), .B(u0_cs4_bF_buf1), .Y(u0__abc_49347_n3385) );
  AND2X2 AND2X2_1008 ( .A(u0__abc_49347_n3386), .B(u0__abc_49347_n2725_bF_buf2), .Y(u0__abc_49347_n3387) );
  AND2X2 AND2X2_1009 ( .A(u0_tms3_27_), .B(u0_cs3_bF_buf1), .Y(u0__abc_49347_n3388) );
  AND2X2 AND2X2_101 ( .A(u0__abc_49347_n1169), .B(u0__abc_49347_n1149_1), .Y(u0__abc_49347_n1170_1) );
  AND2X2 AND2X2_1010 ( .A(u0__abc_49347_n3389), .B(u0__abc_49347_n2724_bF_buf2), .Y(u0__abc_49347_n3390) );
  AND2X2 AND2X2_1011 ( .A(u0_tms2_27_), .B(u0_cs2_bF_buf1), .Y(u0__abc_49347_n3391) );
  AND2X2 AND2X2_1012 ( .A(u0__abc_49347_n3392), .B(u0__abc_49347_n2723_bF_buf2), .Y(u0__abc_49347_n3393) );
  AND2X2 AND2X2_1013 ( .A(u0_tms1_27_), .B(u0_cs1_bF_buf1), .Y(u0__abc_49347_n3394) );
  AND2X2 AND2X2_1014 ( .A(u0__abc_49347_n1175_bF_buf6), .B(u0__abc_49347_n3397), .Y(u0__abc_49347_n3398) );
  AND2X2 AND2X2_1015 ( .A(u0__abc_49347_n3396), .B(u0__abc_49347_n3398), .Y(u0__abc_49347_n3399) );
  AND2X2 AND2X2_1016 ( .A(u0__abc_49347_n1953_1_bF_buf2), .B(csc_1_), .Y(u0__abc_49347_n3521) );
  AND2X2 AND2X2_1017 ( .A(u0_csc5_1_), .B(u0_cs5_bF_buf0), .Y(u0__abc_49347_n3522) );
  AND2X2 AND2X2_1018 ( .A(u0__abc_49347_n3524), .B(u0__abc_49347_n2730_bF_buf1), .Y(u0__abc_49347_n3525) );
  AND2X2 AND2X2_1019 ( .A(u0__abc_49347_n3525), .B(u0__abc_49347_n3523), .Y(u0__abc_49347_n3526) );
  AND2X2 AND2X2_102 ( .A(u0__abc_49347_n1170_1), .B(u0__abc_49347_n1135_1), .Y(u0__abc_49347_n1171) );
  AND2X2 AND2X2_1020 ( .A(u0__abc_49347_n3527), .B(u0__abc_49347_n2726_bF_buf1), .Y(u0__abc_49347_n3528) );
  AND2X2 AND2X2_1021 ( .A(u0_csc4_1_), .B(u0_cs4_bF_buf0), .Y(u0__abc_49347_n3529) );
  AND2X2 AND2X2_1022 ( .A(u0__abc_49347_n3530), .B(u0__abc_49347_n2725_bF_buf1), .Y(u0__abc_49347_n3531) );
  AND2X2 AND2X2_1023 ( .A(u0_csc3_1_), .B(u0_cs3_bF_buf0), .Y(u0__abc_49347_n3532) );
  AND2X2 AND2X2_1024 ( .A(u0__abc_49347_n3533), .B(u0__abc_49347_n2724_bF_buf1), .Y(u0__abc_49347_n3534) );
  AND2X2 AND2X2_1025 ( .A(u0_csc2_1_), .B(u0_cs2_bF_buf0), .Y(u0__abc_49347_n3535) );
  AND2X2 AND2X2_1026 ( .A(u0__abc_49347_n3536), .B(u0__abc_49347_n2723_bF_buf1), .Y(u0__abc_49347_n3537) );
  AND2X2 AND2X2_1027 ( .A(u0_csc1_1_), .B(u0_cs1_bF_buf0), .Y(u0__abc_49347_n3538) );
  AND2X2 AND2X2_1028 ( .A(u0__abc_49347_n1952_1_bF_buf1), .B(u0__abc_49347_n3541), .Y(u0__abc_49347_n3542) );
  AND2X2 AND2X2_1029 ( .A(u0__abc_49347_n3540), .B(u0__abc_49347_n3542), .Y(u0__abc_49347_n3543) );
  AND2X2 AND2X2_103 ( .A(wb_stb_i_bF_buf4), .B(wb_cyc_i), .Y(u0__abc_49347_n1173) );
  AND2X2 AND2X2_1030 ( .A(u0__abc_49347_n1953_1_bF_buf1), .B(csc_2_), .Y(u0__abc_49347_n3545) );
  AND2X2 AND2X2_1031 ( .A(u0_csc5_2_), .B(u0_cs5_bF_buf5), .Y(u0__abc_49347_n3546) );
  AND2X2 AND2X2_1032 ( .A(u0__abc_49347_n3548), .B(u0__abc_49347_n2730_bF_buf0), .Y(u0__abc_49347_n3549) );
  AND2X2 AND2X2_1033 ( .A(u0__abc_49347_n3549), .B(u0__abc_49347_n3547), .Y(u0__abc_49347_n3550) );
  AND2X2 AND2X2_1034 ( .A(u0__abc_49347_n3551), .B(u0__abc_49347_n2726_bF_buf0), .Y(u0__abc_49347_n3552) );
  AND2X2 AND2X2_1035 ( .A(u0_csc4_2_), .B(u0_cs4_bF_buf5), .Y(u0__abc_49347_n3553) );
  AND2X2 AND2X2_1036 ( .A(u0__abc_49347_n3554), .B(u0__abc_49347_n2725_bF_buf0), .Y(u0__abc_49347_n3555) );
  AND2X2 AND2X2_1037 ( .A(u0_csc3_2_), .B(u0_cs3_bF_buf5), .Y(u0__abc_49347_n3556) );
  AND2X2 AND2X2_1038 ( .A(u0__abc_49347_n3557), .B(u0__abc_49347_n2724_bF_buf0), .Y(u0__abc_49347_n3558) );
  AND2X2 AND2X2_1039 ( .A(u0_csc2_2_), .B(u0_cs2_bF_buf5), .Y(u0__abc_49347_n3559) );
  AND2X2 AND2X2_104 ( .A(u0__abc_49347_n1174_1), .B(u0__abc_49347_n1173), .Y(u0__abc_49347_n1175) );
  AND2X2 AND2X2_1040 ( .A(u0__abc_49347_n3560), .B(u0__abc_49347_n2723_bF_buf0), .Y(u0__abc_49347_n3561) );
  AND2X2 AND2X2_1041 ( .A(u0_csc1_2_), .B(u0_cs1_bF_buf5), .Y(u0__abc_49347_n3562) );
  AND2X2 AND2X2_1042 ( .A(u0__abc_49347_n1952_1_bF_buf0), .B(u0__abc_49347_n3565), .Y(u0__abc_49347_n3566) );
  AND2X2 AND2X2_1043 ( .A(u0__abc_49347_n3564), .B(u0__abc_49347_n3566), .Y(u0__abc_49347_n3567) );
  AND2X2 AND2X2_1044 ( .A(u0__abc_49347_n1953_1_bF_buf0), .B(csc_3_), .Y(u0__abc_49347_n3569) );
  AND2X2 AND2X2_1045 ( .A(u0_csc5_3_), .B(u0_cs5_bF_buf4), .Y(u0__abc_49347_n3570) );
  AND2X2 AND2X2_1046 ( .A(u0__abc_49347_n3572), .B(u0__abc_49347_n2730_bF_buf5), .Y(u0__abc_49347_n3573) );
  AND2X2 AND2X2_1047 ( .A(u0__abc_49347_n3573), .B(u0__abc_49347_n3571), .Y(u0__abc_49347_n3574) );
  AND2X2 AND2X2_1048 ( .A(u0__abc_49347_n3575), .B(u0__abc_49347_n2726_bF_buf5), .Y(u0__abc_49347_n3576) );
  AND2X2 AND2X2_1049 ( .A(u0_csc4_3_), .B(u0_cs4_bF_buf4), .Y(u0__abc_49347_n3577) );
  AND2X2 AND2X2_105 ( .A(u0__abc_49347_n1176_1_bF_buf6), .B(sp_tms_0_), .Y(u0__abc_49347_n1177) );
  AND2X2 AND2X2_1050 ( .A(u0__abc_49347_n3578), .B(u0__abc_49347_n2725_bF_buf5), .Y(u0__abc_49347_n3579) );
  AND2X2 AND2X2_1051 ( .A(u0_csc3_3_), .B(u0_cs3_bF_buf4), .Y(u0__abc_49347_n3580) );
  AND2X2 AND2X2_1052 ( .A(u0__abc_49347_n3581), .B(u0__abc_49347_n2724_bF_buf5), .Y(u0__abc_49347_n3582) );
  AND2X2 AND2X2_1053 ( .A(u0_csc2_3_), .B(u0_cs2_bF_buf4), .Y(u0__abc_49347_n3583) );
  AND2X2 AND2X2_1054 ( .A(u0__abc_49347_n3584), .B(u0__abc_49347_n2723_bF_buf5), .Y(u0__abc_49347_n3585) );
  AND2X2 AND2X2_1055 ( .A(u0_csc1_3_), .B(u0_cs1_bF_buf4), .Y(u0__abc_49347_n3586) );
  AND2X2 AND2X2_1056 ( .A(u0__abc_49347_n1952_1_bF_buf3), .B(u0__abc_49347_n3589), .Y(u0__abc_49347_n3590) );
  AND2X2 AND2X2_1057 ( .A(u0__abc_49347_n3588), .B(u0__abc_49347_n3590), .Y(u0__abc_49347_n3591) );
  AND2X2 AND2X2_1058 ( .A(u0__abc_49347_n1953_1_bF_buf3), .B(csc_4_), .Y(u0__abc_49347_n3593) );
  AND2X2 AND2X2_1059 ( .A(u0_csc5_4_), .B(u0_cs5_bF_buf3), .Y(u0__abc_49347_n3594) );
  AND2X2 AND2X2_106 ( .A(spec_req_cs_5_bF_buf3), .B(u0_tms5_0_), .Y(u0__abc_49347_n1182_1) );
  AND2X2 AND2X2_1060 ( .A(u0__abc_49347_n3596), .B(u0__abc_49347_n2730_bF_buf4), .Y(u0__abc_49347_n3597) );
  AND2X2 AND2X2_1061 ( .A(u0__abc_49347_n3597), .B(u0__abc_49347_n3595), .Y(u0__abc_49347_n3598) );
  AND2X2 AND2X2_1062 ( .A(u0__abc_49347_n3599), .B(u0__abc_49347_n2726_bF_buf4), .Y(u0__abc_49347_n3600) );
  AND2X2 AND2X2_1063 ( .A(u0_csc4_4_), .B(u0_cs4_bF_buf3), .Y(u0__abc_49347_n3601) );
  AND2X2 AND2X2_1064 ( .A(u0__abc_49347_n3602), .B(u0__abc_49347_n2725_bF_buf4), .Y(u0__abc_49347_n3603) );
  AND2X2 AND2X2_1065 ( .A(u0_csc3_4_), .B(u0_cs3_bF_buf3), .Y(u0__abc_49347_n3604) );
  AND2X2 AND2X2_1066 ( .A(u0__abc_49347_n3605), .B(u0__abc_49347_n2724_bF_buf4), .Y(u0__abc_49347_n3606) );
  AND2X2 AND2X2_1067 ( .A(u0_csc2_4_), .B(u0_cs2_bF_buf3), .Y(u0__abc_49347_n3607) );
  AND2X2 AND2X2_1068 ( .A(u0__abc_49347_n3608), .B(u0__abc_49347_n2723_bF_buf4), .Y(u0__abc_49347_n3609) );
  AND2X2 AND2X2_1069 ( .A(u0_csc1_4_), .B(u0_cs1_bF_buf3), .Y(u0__abc_49347_n3610) );
  AND2X2 AND2X2_107 ( .A(u0__abc_49347_n1186), .B(u0__abc_49347_n1185_bF_buf5), .Y(u0__abc_49347_n1187) );
  AND2X2 AND2X2_1070 ( .A(u0__abc_49347_n1952_1_bF_buf2), .B(u0__abc_49347_n3613), .Y(u0__abc_49347_n3614) );
  AND2X2 AND2X2_1071 ( .A(u0__abc_49347_n3612), .B(u0__abc_49347_n3614), .Y(u0__abc_49347_n3615) );
  AND2X2 AND2X2_1072 ( .A(u0__abc_49347_n1953_1_bF_buf2), .B(csc_5_bF_buf3), .Y(u0__abc_49347_n3617) );
  AND2X2 AND2X2_1073 ( .A(u0_csc5_5_), .B(u0_cs5_bF_buf2), .Y(u0__abc_49347_n3618) );
  AND2X2 AND2X2_1074 ( .A(u0__abc_49347_n3620), .B(u0__abc_49347_n2730_bF_buf3), .Y(u0__abc_49347_n3621) );
  AND2X2 AND2X2_1075 ( .A(u0__abc_49347_n3621), .B(u0__abc_49347_n3619), .Y(u0__abc_49347_n3622) );
  AND2X2 AND2X2_1076 ( .A(u0__abc_49347_n3623), .B(u0__abc_49347_n2726_bF_buf3), .Y(u0__abc_49347_n3624) );
  AND2X2 AND2X2_1077 ( .A(u0_csc4_5_), .B(u0_cs4_bF_buf2), .Y(u0__abc_49347_n3625) );
  AND2X2 AND2X2_1078 ( .A(u0__abc_49347_n3626), .B(u0__abc_49347_n2725_bF_buf3), .Y(u0__abc_49347_n3627) );
  AND2X2 AND2X2_1079 ( .A(u0_csc3_5_), .B(u0_cs3_bF_buf2), .Y(u0__abc_49347_n3628) );
  AND2X2 AND2X2_108 ( .A(u0__abc_49347_n1187), .B(u0__abc_49347_n1184), .Y(u0__abc_49347_n1188) );
  AND2X2 AND2X2_1080 ( .A(u0__abc_49347_n3629), .B(u0__abc_49347_n2724_bF_buf3), .Y(u0__abc_49347_n3630) );
  AND2X2 AND2X2_1081 ( .A(u0_csc2_5_), .B(u0_cs2_bF_buf2), .Y(u0__abc_49347_n3631) );
  AND2X2 AND2X2_1082 ( .A(u0__abc_49347_n3632), .B(u0__abc_49347_n2723_bF_buf3), .Y(u0__abc_49347_n3633) );
  AND2X2 AND2X2_1083 ( .A(u0_csc1_5_), .B(u0_cs1_bF_buf2), .Y(u0__abc_49347_n3634) );
  AND2X2 AND2X2_1084 ( .A(u0__abc_49347_n1952_1_bF_buf1), .B(u0__abc_49347_n3637), .Y(u0__abc_49347_n3638) );
  AND2X2 AND2X2_1085 ( .A(u0__abc_49347_n3636), .B(u0__abc_49347_n3638), .Y(u0__abc_49347_n3639) );
  AND2X2 AND2X2_1086 ( .A(u0__abc_49347_n1953_1_bF_buf1), .B(csc_6_), .Y(u0__abc_49347_n3641) );
  AND2X2 AND2X2_1087 ( .A(u0_csc5_6_), .B(u0_cs5_bF_buf1), .Y(u0__abc_49347_n3642) );
  AND2X2 AND2X2_1088 ( .A(u0__abc_49347_n3644), .B(u0__abc_49347_n2730_bF_buf2), .Y(u0__abc_49347_n3645) );
  AND2X2 AND2X2_1089 ( .A(u0__abc_49347_n3645), .B(u0__abc_49347_n3643), .Y(u0__abc_49347_n3646) );
  AND2X2 AND2X2_109 ( .A(u0__abc_49347_n1189), .B(u0__abc_49347_n1181_bF_buf5), .Y(u0__abc_49347_n1190) );
  AND2X2 AND2X2_1090 ( .A(u0__abc_49347_n3647), .B(u0__abc_49347_n2726_bF_buf2), .Y(u0__abc_49347_n3648) );
  AND2X2 AND2X2_1091 ( .A(u0_csc4_6_), .B(u0_cs4_bF_buf1), .Y(u0__abc_49347_n3649) );
  AND2X2 AND2X2_1092 ( .A(u0__abc_49347_n3650), .B(u0__abc_49347_n2725_bF_buf2), .Y(u0__abc_49347_n3651) );
  AND2X2 AND2X2_1093 ( .A(u0_csc3_6_), .B(u0_cs3_bF_buf1), .Y(u0__abc_49347_n3652) );
  AND2X2 AND2X2_1094 ( .A(u0__abc_49347_n3653), .B(u0__abc_49347_n2724_bF_buf2), .Y(u0__abc_49347_n3654) );
  AND2X2 AND2X2_1095 ( .A(u0_csc2_6_), .B(u0_cs2_bF_buf1), .Y(u0__abc_49347_n3655) );
  AND2X2 AND2X2_1096 ( .A(u0__abc_49347_n3656), .B(u0__abc_49347_n2723_bF_buf2), .Y(u0__abc_49347_n3657) );
  AND2X2 AND2X2_1097 ( .A(u0_csc1_6_), .B(u0_cs1_bF_buf1), .Y(u0__abc_49347_n3658) );
  AND2X2 AND2X2_1098 ( .A(u0__abc_49347_n1952_1_bF_buf0), .B(u0__abc_49347_n3661), .Y(u0__abc_49347_n3662) );
  AND2X2 AND2X2_1099 ( .A(u0__abc_49347_n3660), .B(u0__abc_49347_n3662), .Y(u0__abc_49347_n3663) );
  AND2X2 AND2X2_11 ( .A(_abc_55805_n269), .B(_abc_55805_n270), .Y(obct_cs_4_) );
  AND2X2 AND2X2_110 ( .A(spec_req_cs_4_bF_buf2), .B(u0_tms4_0_), .Y(u0__abc_49347_n1191_1) );
  AND2X2 AND2X2_1100 ( .A(u0__abc_49347_n1953_1_bF_buf0), .B(csc_7_), .Y(u0__abc_49347_n3665) );
  AND2X2 AND2X2_1101 ( .A(u0_csc5_7_), .B(u0_cs5_bF_buf0), .Y(u0__abc_49347_n3666) );
  AND2X2 AND2X2_1102 ( .A(u0__abc_49347_n3668), .B(u0__abc_49347_n2730_bF_buf1), .Y(u0__abc_49347_n3669) );
  AND2X2 AND2X2_1103 ( .A(u0__abc_49347_n3669), .B(u0__abc_49347_n3667), .Y(u0__abc_49347_n3670) );
  AND2X2 AND2X2_1104 ( .A(u0__abc_49347_n3671), .B(u0__abc_49347_n2726_bF_buf1), .Y(u0__abc_49347_n3672) );
  AND2X2 AND2X2_1105 ( .A(u0_csc4_7_), .B(u0_cs4_bF_buf0), .Y(u0__abc_49347_n3673) );
  AND2X2 AND2X2_1106 ( .A(u0__abc_49347_n3674), .B(u0__abc_49347_n2725_bF_buf1), .Y(u0__abc_49347_n3675) );
  AND2X2 AND2X2_1107 ( .A(u0_csc3_7_), .B(u0_cs3_bF_buf0), .Y(u0__abc_49347_n3676) );
  AND2X2 AND2X2_1108 ( .A(u0__abc_49347_n3677), .B(u0__abc_49347_n2724_bF_buf1), .Y(u0__abc_49347_n3678) );
  AND2X2 AND2X2_1109 ( .A(u0_csc2_7_), .B(u0_cs2_bF_buf0), .Y(u0__abc_49347_n3679) );
  AND2X2 AND2X2_111 ( .A(u0__abc_49347_n1192_1), .B(u0__abc_49347_n1180_1_bF_buf5), .Y(u0__abc_49347_n1193) );
  AND2X2 AND2X2_1110 ( .A(u0__abc_49347_n3680), .B(u0__abc_49347_n2723_bF_buf1), .Y(u0__abc_49347_n3681) );
  AND2X2 AND2X2_1111 ( .A(u0_csc1_7_), .B(u0_cs1_bF_buf0), .Y(u0__abc_49347_n3682) );
  AND2X2 AND2X2_1112 ( .A(u0__abc_49347_n1952_1_bF_buf3), .B(u0__abc_49347_n3685), .Y(u0__abc_49347_n3686) );
  AND2X2 AND2X2_1113 ( .A(u0__abc_49347_n3684), .B(u0__abc_49347_n3686), .Y(u0__abc_49347_n3687) );
  AND2X2 AND2X2_1114 ( .A(u0__abc_49347_n1953_1_bF_buf3), .B(csc_9_), .Y(u0__abc_49347_n3713) );
  AND2X2 AND2X2_1115 ( .A(u0_csc5_9_), .B(u0_cs5_bF_buf5), .Y(u0__abc_49347_n3714) );
  AND2X2 AND2X2_1116 ( .A(u0__abc_49347_n3716), .B(u0__abc_49347_n2730_bF_buf0), .Y(u0__abc_49347_n3717) );
  AND2X2 AND2X2_1117 ( .A(u0__abc_49347_n3717), .B(u0__abc_49347_n3715), .Y(u0__abc_49347_n3718) );
  AND2X2 AND2X2_1118 ( .A(u0__abc_49347_n3719), .B(u0__abc_49347_n2726_bF_buf0), .Y(u0__abc_49347_n3720) );
  AND2X2 AND2X2_1119 ( .A(u0_csc4_9_), .B(u0_cs4_bF_buf5), .Y(u0__abc_49347_n3721) );
  AND2X2 AND2X2_112 ( .A(spec_req_cs_3_bF_buf2), .B(u0_tms3_0_), .Y(u0__abc_49347_n1194) );
  AND2X2 AND2X2_1120 ( .A(u0__abc_49347_n3722), .B(u0__abc_49347_n2725_bF_buf0), .Y(u0__abc_49347_n3723) );
  AND2X2 AND2X2_1121 ( .A(u0_csc3_9_), .B(u0_cs3_bF_buf5), .Y(u0__abc_49347_n3724) );
  AND2X2 AND2X2_1122 ( .A(u0__abc_49347_n3725), .B(u0__abc_49347_n2724_bF_buf0), .Y(u0__abc_49347_n3726) );
  AND2X2 AND2X2_1123 ( .A(u0_csc2_9_), .B(u0_cs2_bF_buf5), .Y(u0__abc_49347_n3727) );
  AND2X2 AND2X2_1124 ( .A(u0__abc_49347_n3728), .B(u0__abc_49347_n2723_bF_buf0), .Y(u0__abc_49347_n3729) );
  AND2X2 AND2X2_1125 ( .A(u0_csc1_9_), .B(u0_cs1_bF_buf5), .Y(u0__abc_49347_n3730) );
  AND2X2 AND2X2_1126 ( .A(u0__abc_49347_n1952_1_bF_buf2), .B(u0__abc_49347_n3733), .Y(u0__abc_49347_n3734) );
  AND2X2 AND2X2_1127 ( .A(u0__abc_49347_n3732), .B(u0__abc_49347_n3734), .Y(u0__abc_49347_n3735) );
  AND2X2 AND2X2_1128 ( .A(u0__abc_49347_n1953_1_bF_buf2), .B(csc_10_), .Y(u0__abc_49347_n3737) );
  AND2X2 AND2X2_1129 ( .A(u0_csc5_10_), .B(u0_cs5_bF_buf4), .Y(u0__abc_49347_n3738) );
  AND2X2 AND2X2_113 ( .A(u0__abc_49347_n1195), .B(u0__abc_49347_n1179_bF_buf5), .Y(u0__abc_49347_n1196) );
  AND2X2 AND2X2_1130 ( .A(u0__abc_49347_n3740), .B(u0__abc_49347_n2730_bF_buf5), .Y(u0__abc_49347_n3741) );
  AND2X2 AND2X2_1131 ( .A(u0__abc_49347_n3741), .B(u0__abc_49347_n3739), .Y(u0__abc_49347_n3742) );
  AND2X2 AND2X2_1132 ( .A(u0__abc_49347_n3743), .B(u0__abc_49347_n2726_bF_buf5), .Y(u0__abc_49347_n3744) );
  AND2X2 AND2X2_1133 ( .A(u0_csc4_10_), .B(u0_cs4_bF_buf4), .Y(u0__abc_49347_n3745) );
  AND2X2 AND2X2_1134 ( .A(u0__abc_49347_n3746), .B(u0__abc_49347_n2725_bF_buf5), .Y(u0__abc_49347_n3747) );
  AND2X2 AND2X2_1135 ( .A(u0_csc3_10_), .B(u0_cs3_bF_buf4), .Y(u0__abc_49347_n3748) );
  AND2X2 AND2X2_1136 ( .A(u0__abc_49347_n3749), .B(u0__abc_49347_n2724_bF_buf5), .Y(u0__abc_49347_n3750) );
  AND2X2 AND2X2_1137 ( .A(u0_csc2_10_), .B(u0_cs2_bF_buf4), .Y(u0__abc_49347_n3751) );
  AND2X2 AND2X2_1138 ( .A(u0__abc_49347_n3752), .B(u0__abc_49347_n2723_bF_buf5), .Y(u0__abc_49347_n3753) );
  AND2X2 AND2X2_1139 ( .A(u0_csc1_10_), .B(u0_cs1_bF_buf4), .Y(u0__abc_49347_n3754) );
  AND2X2 AND2X2_114 ( .A(spec_req_cs_2_bF_buf2), .B(u0_tms2_0_), .Y(u0__abc_49347_n1197) );
  AND2X2 AND2X2_1140 ( .A(u0__abc_49347_n1952_1_bF_buf1), .B(u0__abc_49347_n3757), .Y(u0__abc_49347_n3758) );
  AND2X2 AND2X2_1141 ( .A(u0__abc_49347_n3756), .B(u0__abc_49347_n3758), .Y(u0__abc_49347_n3759) );
  AND2X2 AND2X2_1142 ( .A(u0__abc_49347_n1953_1_bF_buf1), .B(u3_pen), .Y(u0__abc_49347_n3761) );
  AND2X2 AND2X2_1143 ( .A(u0_csc5_11_), .B(u0_cs5_bF_buf3), .Y(u0__abc_49347_n3762) );
  AND2X2 AND2X2_1144 ( .A(u0__abc_49347_n3764), .B(u0__abc_49347_n2730_bF_buf4), .Y(u0__abc_49347_n3765) );
  AND2X2 AND2X2_1145 ( .A(u0__abc_49347_n3765), .B(u0__abc_49347_n3763), .Y(u0__abc_49347_n3766) );
  AND2X2 AND2X2_1146 ( .A(u0__abc_49347_n3767), .B(u0__abc_49347_n2726_bF_buf4), .Y(u0__abc_49347_n3768) );
  AND2X2 AND2X2_1147 ( .A(u0_csc4_11_), .B(u0_cs4_bF_buf3), .Y(u0__abc_49347_n3769) );
  AND2X2 AND2X2_1148 ( .A(u0__abc_49347_n3770), .B(u0__abc_49347_n2725_bF_buf4), .Y(u0__abc_49347_n3771) );
  AND2X2 AND2X2_1149 ( .A(u0_csc3_11_), .B(u0_cs3_bF_buf3), .Y(u0__abc_49347_n3772) );
  AND2X2 AND2X2_115 ( .A(u0__abc_49347_n1198), .B(u0__abc_49347_n1178_1_bF_buf5), .Y(u0__abc_49347_n1199) );
  AND2X2 AND2X2_1150 ( .A(u0__abc_49347_n3773), .B(u0__abc_49347_n2724_bF_buf4), .Y(u0__abc_49347_n3774) );
  AND2X2 AND2X2_1151 ( .A(u0_csc2_11_), .B(u0_cs2_bF_buf3), .Y(u0__abc_49347_n3775) );
  AND2X2 AND2X2_1152 ( .A(u0__abc_49347_n3776), .B(u0__abc_49347_n2723_bF_buf4), .Y(u0__abc_49347_n3777) );
  AND2X2 AND2X2_1153 ( .A(u0_csc1_11_), .B(u0_cs1_bF_buf3), .Y(u0__abc_49347_n3778) );
  AND2X2 AND2X2_1154 ( .A(u0__abc_49347_n1952_1_bF_buf0), .B(u0__abc_49347_n3781), .Y(u0__abc_49347_n3782) );
  AND2X2 AND2X2_1155 ( .A(u0__abc_49347_n3780), .B(u0__abc_49347_n3782), .Y(u0__abc_49347_n3783) );
  AND2X2 AND2X2_1156 ( .A(u0__abc_49347_n1173), .B(cs_le_bF_buf4), .Y(u0__abc_49347_n4265) );
  AND2X2 AND2X2_1157 ( .A(u0__abc_49347_n4272), .B(u0__abc_49347_n4265), .Y(u0__abc_49347_n4273) );
  AND2X2 AND2X2_1158 ( .A(wb_cyc_i), .B(u0_wp_err), .Y(u0__abc_49347_n4275) );
  AND2X2 AND2X2_1159 ( .A(u0__abc_49347_n4274), .B(u0__abc_49347_n4275), .Y(u0__abc_49347_n4276) );
  AND2X2 AND2X2_116 ( .A(spec_req_cs_1_bF_buf2), .B(u0_tms1_0_), .Y(u0__abc_49347_n1200_1) );
  AND2X2 AND2X2_1160 ( .A(u0__abc_49347_n4280), .B(u0__abc_49347_n4278), .Y(u0_cs_0__FF_INPUT) );
  AND2X2 AND2X2_1161 ( .A(u0__abc_49347_n4283), .B(u0__abc_49347_n4282), .Y(u0_cs_1__FF_INPUT) );
  AND2X2 AND2X2_1162 ( .A(u0__abc_49347_n4286), .B(u0__abc_49347_n4285), .Y(u0_cs_2__FF_INPUT) );
  AND2X2 AND2X2_1163 ( .A(u0__abc_49347_n4289), .B(u0__abc_49347_n4288), .Y(u0_cs_3__FF_INPUT) );
  AND2X2 AND2X2_1164 ( .A(u0__abc_49347_n4292), .B(u0__abc_49347_n4291), .Y(u0_cs_4__FF_INPUT) );
  AND2X2 AND2X2_1165 ( .A(u0__abc_49347_n4295), .B(u0__abc_49347_n4294), .Y(u0_cs_5__FF_INPUT) );
  AND2X2 AND2X2_1166 ( .A(u0__abc_49347_n4298), .B(u0__abc_49347_n4297), .Y(u0_cs_6__FF_INPUT) );
  AND2X2 AND2X2_1167 ( .A(u0__abc_49347_n4301), .B(u0__abc_49347_n4300), .Y(u0_cs_7__FF_INPUT) );
  AND2X2 AND2X2_1168 ( .A(u0__abc_49347_n4305), .B(u0__abc_49347_n4303), .Y(u0_poc_0__FF_INPUT) );
  AND2X2 AND2X2_1169 ( .A(u0__abc_49347_n4308), .B(u0__abc_49347_n4307), .Y(u0_poc_1__FF_INPUT) );
  AND2X2 AND2X2_117 ( .A(u0__abc_49347_n1175_bF_buf5), .B(u0__abc_49347_n1204), .Y(u0__abc_49347_n1205) );
  AND2X2 AND2X2_1170 ( .A(u0__abc_49347_n4311), .B(u0__abc_49347_n4310), .Y(u0_poc_2__FF_INPUT) );
  AND2X2 AND2X2_1171 ( .A(u0__abc_49347_n4314), .B(u0__abc_49347_n4313), .Y(u0_poc_3__FF_INPUT) );
  AND2X2 AND2X2_1172 ( .A(u0__abc_49347_n4317), .B(u0__abc_49347_n4316), .Y(u0_poc_4__FF_INPUT) );
  AND2X2 AND2X2_1173 ( .A(u0__abc_49347_n4320), .B(u0__abc_49347_n4319), .Y(u0_poc_5__FF_INPUT) );
  AND2X2 AND2X2_1174 ( .A(u0__abc_49347_n4323), .B(u0__abc_49347_n4322), .Y(u0_poc_6__FF_INPUT) );
  AND2X2 AND2X2_1175 ( .A(u0__abc_49347_n4326), .B(u0__abc_49347_n4325), .Y(u0_poc_7__FF_INPUT) );
  AND2X2 AND2X2_1176 ( .A(u0__abc_49347_n4329), .B(u0__abc_49347_n4328), .Y(u0_poc_8__FF_INPUT) );
  AND2X2 AND2X2_1177 ( .A(u0__abc_49347_n4332), .B(u0__abc_49347_n4331), .Y(u0_poc_9__FF_INPUT) );
  AND2X2 AND2X2_1178 ( .A(u0__abc_49347_n4335), .B(u0__abc_49347_n4334), .Y(u0_poc_10__FF_INPUT) );
  AND2X2 AND2X2_1179 ( .A(u0__abc_49347_n4338), .B(u0__abc_49347_n4337), .Y(u0_poc_11__FF_INPUT) );
  AND2X2 AND2X2_118 ( .A(u0__abc_49347_n1202), .B(u0__abc_49347_n1205), .Y(u0__abc_49347_n1206) );
  AND2X2 AND2X2_1180 ( .A(u0__abc_49347_n4341), .B(u0__abc_49347_n4340), .Y(u0_poc_12__FF_INPUT) );
  AND2X2 AND2X2_1181 ( .A(u0__abc_49347_n4344), .B(u0__abc_49347_n4343), .Y(u0_poc_13__FF_INPUT) );
  AND2X2 AND2X2_1182 ( .A(u0__abc_49347_n4347), .B(u0__abc_49347_n4346), .Y(u0_poc_14__FF_INPUT) );
  AND2X2 AND2X2_1183 ( .A(u0__abc_49347_n4350), .B(u0__abc_49347_n4349), .Y(u0_poc_15__FF_INPUT) );
  AND2X2 AND2X2_1184 ( .A(u0__abc_49347_n4353), .B(u0__abc_49347_n4352), .Y(u0_poc_16__FF_INPUT) );
  AND2X2 AND2X2_1185 ( .A(u0__abc_49347_n4356), .B(u0__abc_49347_n4355), .Y(u0_poc_17__FF_INPUT) );
  AND2X2 AND2X2_1186 ( .A(u0__abc_49347_n4359), .B(u0__abc_49347_n4358), .Y(u0_poc_18__FF_INPUT) );
  AND2X2 AND2X2_1187 ( .A(u0__abc_49347_n4362), .B(u0__abc_49347_n4361), .Y(u0_poc_19__FF_INPUT) );
  AND2X2 AND2X2_1188 ( .A(u0__abc_49347_n4365), .B(u0__abc_49347_n4364), .Y(u0_poc_20__FF_INPUT) );
  AND2X2 AND2X2_1189 ( .A(u0__abc_49347_n4368), .B(u0__abc_49347_n4367), .Y(u0_poc_21__FF_INPUT) );
  AND2X2 AND2X2_119 ( .A(u0__abc_49347_n1176_1_bF_buf5), .B(sp_tms_1_), .Y(u0__abc_49347_n1208) );
  AND2X2 AND2X2_1190 ( .A(u0__abc_49347_n4371), .B(u0__abc_49347_n4370), .Y(u0_poc_22__FF_INPUT) );
  AND2X2 AND2X2_1191 ( .A(u0__abc_49347_n4374), .B(u0__abc_49347_n4373), .Y(u0_poc_23__FF_INPUT) );
  AND2X2 AND2X2_1192 ( .A(u0__abc_49347_n4377), .B(u0__abc_49347_n4376), .Y(u0_poc_24__FF_INPUT) );
  AND2X2 AND2X2_1193 ( .A(u0__abc_49347_n4380), .B(u0__abc_49347_n4379), .Y(u0_poc_25__FF_INPUT) );
  AND2X2 AND2X2_1194 ( .A(u0__abc_49347_n4383), .B(u0__abc_49347_n4382), .Y(u0_poc_26__FF_INPUT) );
  AND2X2 AND2X2_1195 ( .A(u0__abc_49347_n4386), .B(u0__abc_49347_n4385), .Y(u0_poc_27__FF_INPUT) );
  AND2X2 AND2X2_1196 ( .A(u0__abc_49347_n4389), .B(u0__abc_49347_n4388), .Y(u0_poc_28__FF_INPUT) );
  AND2X2 AND2X2_1197 ( .A(u0__abc_49347_n4392), .B(u0__abc_49347_n4391), .Y(u0_poc_29__FF_INPUT) );
  AND2X2 AND2X2_1198 ( .A(u0__abc_49347_n4395), .B(u0__abc_49347_n4394), .Y(u0_poc_30__FF_INPUT) );
  AND2X2 AND2X2_1199 ( .A(u0__abc_49347_n4398), .B(u0__abc_49347_n4397), .Y(u0_poc_31__FF_INPUT) );
  AND2X2 AND2X2_12 ( .A(_abc_55805_n272), .B(_abc_55805_n273), .Y(_abc_55805_n274) );
  AND2X2 AND2X2_120 ( .A(spec_req_cs_5_bF_buf1), .B(u0_tms5_1_), .Y(u0__abc_49347_n1209_1) );
  AND2X2 AND2X2_1200 ( .A(u0__abc_49347_n4405), .B(u0_wb_addr_r_3_), .Y(u0__abc_49347_n4406) );
  AND2X2 AND2X2_1201 ( .A(u0__abc_49347_n4403), .B(u0__abc_49347_n4406), .Y(u0__abc_49347_n4407) );
  AND2X2 AND2X2_1202 ( .A(u0__abc_49347_n4410), .B(u0__abc_49347_n4408), .Y(u0_csc_mask_r_0__FF_INPUT) );
  AND2X2 AND2X2_1203 ( .A(u0__abc_49347_n4413), .B(u0__abc_49347_n4412), .Y(u0_csc_mask_r_1__FF_INPUT) );
  AND2X2 AND2X2_1204 ( .A(u0__abc_49347_n4416), .B(u0__abc_49347_n4415), .Y(u0_csc_mask_r_2__FF_INPUT) );
  AND2X2 AND2X2_1205 ( .A(u0__abc_49347_n4419), .B(u0__abc_49347_n4418), .Y(u0_csc_mask_r_3__FF_INPUT) );
  AND2X2 AND2X2_1206 ( .A(u0__abc_49347_n4422), .B(u0__abc_49347_n4421), .Y(u0_csc_mask_r_4__FF_INPUT) );
  AND2X2 AND2X2_1207 ( .A(u0__abc_49347_n4425), .B(u0__abc_49347_n4424), .Y(u0_csc_mask_r_5__FF_INPUT) );
  AND2X2 AND2X2_1208 ( .A(u0__abc_49347_n4428), .B(u0__abc_49347_n4427), .Y(u0_csc_mask_r_6__FF_INPUT) );
  AND2X2 AND2X2_1209 ( .A(u0__abc_49347_n4431), .B(u0__abc_49347_n4430), .Y(u0_csc_mask_r_7__FF_INPUT) );
  AND2X2 AND2X2_121 ( .A(u0__abc_49347_n1211), .B(u0__abc_49347_n1185_bF_buf4), .Y(u0__abc_49347_n1212) );
  AND2X2 AND2X2_1210 ( .A(u0__abc_49347_n4434), .B(u0__abc_49347_n4433), .Y(u0_csc_mask_r_8__FF_INPUT) );
  AND2X2 AND2X2_1211 ( .A(u0__abc_49347_n4437), .B(u0__abc_49347_n4436), .Y(u0_csc_mask_r_9__FF_INPUT) );
  AND2X2 AND2X2_1212 ( .A(u0__abc_49347_n4440), .B(u0__abc_49347_n4439), .Y(u0_csc_mask_r_10__FF_INPUT) );
  AND2X2 AND2X2_1213 ( .A(u0__abc_49347_n4445), .B(u0__abc_49347_n4446), .Y(u0_csr_r_0__FF_INPUT) );
  AND2X2 AND2X2_1214 ( .A(u0__abc_49347_n4448), .B(u0__abc_49347_n4449), .Y(u0_csr_r_1__FF_INPUT) );
  AND2X2 AND2X2_1215 ( .A(u0__abc_49347_n4451), .B(u0__abc_49347_n4452), .Y(u0_csr_r_2__FF_INPUT) );
  AND2X2 AND2X2_1216 ( .A(u0__abc_49347_n4454), .B(u0__abc_49347_n4455), .Y(u0_csr_r_3__FF_INPUT) );
  AND2X2 AND2X2_1217 ( .A(u0__abc_49347_n4457), .B(u0__abc_49347_n4458), .Y(u0_csr_r_4__FF_INPUT) );
  AND2X2 AND2X2_1218 ( .A(u0__abc_49347_n4460), .B(u0__abc_49347_n4461), .Y(u0_csr_r_5__FF_INPUT) );
  AND2X2 AND2X2_1219 ( .A(u0__abc_49347_n4463), .B(u0__abc_49347_n4464), .Y(u0_csr_r_6__FF_INPUT) );
  AND2X2 AND2X2_122 ( .A(u0__abc_49347_n1212), .B(u0__abc_49347_n1210_1), .Y(u0__abc_49347_n1213) );
  AND2X2 AND2X2_1220 ( .A(u0__abc_49347_n4466), .B(u0__abc_49347_n4467), .Y(u0_csr_r_7__FF_INPUT) );
  AND2X2 AND2X2_1221 ( .A(u0__abc_49347_n4469), .B(u0__abc_49347_n4470), .Y(u0_csr_r_8__FF_INPUT) );
  AND2X2 AND2X2_1222 ( .A(u0__abc_49347_n4472), .B(u0__abc_49347_n4473), .Y(u0_csr_r_9__FF_INPUT) );
  AND2X2 AND2X2_1223 ( .A(u0__abc_49347_n4475), .B(u0__abc_49347_n4476), .Y(u0_csr_r2_0__FF_INPUT) );
  AND2X2 AND2X2_1224 ( .A(u0__abc_49347_n4478), .B(u0__abc_49347_n4479), .Y(u0_csr_r2_1__FF_INPUT) );
  AND2X2 AND2X2_1225 ( .A(u0__abc_49347_n4481), .B(u0__abc_49347_n4482), .Y(u0_csr_r2_2__FF_INPUT) );
  AND2X2 AND2X2_1226 ( .A(u0__abc_49347_n4484), .B(u0__abc_49347_n4485), .Y(u0_csr_r2_3__FF_INPUT) );
  AND2X2 AND2X2_1227 ( .A(u0__abc_49347_n4487), .B(u0__abc_49347_n4488), .Y(u0_csr_r2_4__FF_INPUT) );
  AND2X2 AND2X2_1228 ( .A(u0__abc_49347_n4490), .B(u0__abc_49347_n4491), .Y(u0_csr_r2_5__FF_INPUT) );
  AND2X2 AND2X2_1229 ( .A(u0__abc_49347_n4493), .B(u0__abc_49347_n4494), .Y(u0_csr_r2_6__FF_INPUT) );
  AND2X2 AND2X2_123 ( .A(u0__abc_49347_n1214), .B(u0__abc_49347_n1181_bF_buf4), .Y(u0__abc_49347_n1215) );
  AND2X2 AND2X2_1230 ( .A(u0__abc_49347_n4496), .B(u0__abc_49347_n4497), .Y(u0_csr_r2_7__FF_INPUT) );
  AND2X2 AND2X2_1231 ( .A(u0__abc_49347_n4499), .B(u0__abc_49347_n4500), .Y(u0__abc_49347_n4501) );
  AND2X2 AND2X2_1232 ( .A(u0__abc_49347_n4503), .B(u0__abc_49347_n4504), .Y(u0__abc_49347_n4505) );
  AND2X2 AND2X2_1233 ( .A(u0__abc_49347_n4505), .B(u0__abc_49347_n4502), .Y(u0__abc_49347_n4506) );
  AND2X2 AND2X2_1234 ( .A(u0__abc_49347_n4506), .B(u0__abc_49347_n4501), .Y(u0__abc_49347_n4507) );
  AND2X2 AND2X2_1235 ( .A(u0__abc_49347_n4507_bF_buf3), .B(u0_csr_0_), .Y(u0__abc_49347_n4508) );
  AND2X2 AND2X2_1236 ( .A(u0__abc_49347_n4503), .B(\wb_addr_i[2] ), .Y(u0__abc_49347_n4509) );
  AND2X2 AND2X2_1237 ( .A(u0__abc_49347_n4509), .B(u0__abc_49347_n4502), .Y(u0__abc_49347_n4510) );
  AND2X2 AND2X2_1238 ( .A(u0__abc_49347_n4510), .B(u0__abc_49347_n4501), .Y(u0__abc_49347_n4511) );
  AND2X2 AND2X2_1239 ( .A(u0__abc_49347_n4511_bF_buf4), .B(_auto_iopadmap_cc_313_execute_56321_0_), .Y(u0__abc_49347_n4512) );
  AND2X2 AND2X2_124 ( .A(spec_req_cs_4_bF_buf1), .B(u0_tms4_1_), .Y(u0__abc_49347_n1216) );
  AND2X2 AND2X2_1240 ( .A(u0__abc_49347_n4499), .B(\wb_addr_i[4] ), .Y(u0__abc_49347_n4513) );
  AND2X2 AND2X2_1241 ( .A(\wb_addr_i[3] ), .B(\wb_addr_i[2] ), .Y(u0__abc_49347_n4514) );
  AND2X2 AND2X2_1242 ( .A(u0__abc_49347_n4514), .B(u0__abc_49347_n4502), .Y(u0__abc_49347_n4515) );
  AND2X2 AND2X2_1243 ( .A(u0__abc_49347_n4515), .B(u0__abc_49347_n4513), .Y(u0__abc_49347_n4516) );
  AND2X2 AND2X2_1244 ( .A(u0__abc_49347_n4516_bF_buf4), .B(u0_tms1_0_), .Y(u0__abc_49347_n4517) );
  AND2X2 AND2X2_1245 ( .A(u0__abc_49347_n4500), .B(\wb_addr_i[5] ), .Y(u0__abc_49347_n4518) );
  AND2X2 AND2X2_1246 ( .A(u0__abc_49347_n4506), .B(u0__abc_49347_n4518), .Y(u0__abc_49347_n4519) );
  AND2X2 AND2X2_1247 ( .A(u0__abc_49347_n4519_bF_buf4), .B(u0_csc2_0_), .Y(u0__abc_49347_n4520) );
  AND2X2 AND2X2_1248 ( .A(u0__abc_49347_n4504), .B(\wb_addr_i[3] ), .Y(u0__abc_49347_n4524) );
  AND2X2 AND2X2_1249 ( .A(u0__abc_49347_n4524), .B(u0__abc_49347_n4502), .Y(u0__abc_49347_n4525) );
  AND2X2 AND2X2_125 ( .A(u0__abc_49347_n1217), .B(u0__abc_49347_n1180_1_bF_buf4), .Y(u0__abc_49347_n1218_1) );
  AND2X2 AND2X2_1250 ( .A(u0__abc_49347_n4525), .B(u0__abc_49347_n4513), .Y(u0__abc_49347_n4526) );
  AND2X2 AND2X2_1251 ( .A(u0__abc_49347_n4526_bF_buf4), .B(u0_csc1_0_), .Y(u0__abc_49347_n4527) );
  AND2X2 AND2X2_1252 ( .A(u0__abc_49347_n4515), .B(u0__abc_49347_n4518), .Y(u0__abc_49347_n4528) );
  AND2X2 AND2X2_1253 ( .A(u0__abc_49347_n4528_bF_buf4), .B(u0_tms3_0_), .Y(u0__abc_49347_n4529) );
  AND2X2 AND2X2_1254 ( .A(\wb_addr_i[5] ), .B(\wb_addr_i[4] ), .Y(u0__abc_49347_n4530) );
  AND2X2 AND2X2_1255 ( .A(u0__abc_49347_n4506), .B(u0__abc_49347_n4530), .Y(u0__abc_49347_n4531) );
  AND2X2 AND2X2_1256 ( .A(u0__abc_49347_n4531_bF_buf4), .B(u0_csc4_0_), .Y(u0__abc_49347_n4532) );
  AND2X2 AND2X2_1257 ( .A(u0__abc_49347_n4510), .B(u0__abc_49347_n4513), .Y(u0__abc_49347_n4535) );
  AND2X2 AND2X2_1258 ( .A(u0__abc_49347_n4535_bF_buf4), .B(u0_tms0_0_), .Y(u0__abc_49347_n4536) );
  AND2X2 AND2X2_1259 ( .A(u0__abc_49347_n4510), .B(u0__abc_49347_n4518), .Y(u0__abc_49347_n4537) );
  AND2X2 AND2X2_126 ( .A(spec_req_cs_3_bF_buf1), .B(u0_tms3_1_), .Y(u0__abc_49347_n1219_1) );
  AND2X2 AND2X2_1260 ( .A(u0__abc_49347_n4537_bF_buf4), .B(u0_tms2_0_), .Y(u0__abc_49347_n4538) );
  AND2X2 AND2X2_1261 ( .A(u0__abc_49347_n4525), .B(u0__abc_49347_n4518), .Y(u0__abc_49347_n4539) );
  AND2X2 AND2X2_1262 ( .A(u0__abc_49347_n4539_bF_buf4), .B(u0_csc3_0_), .Y(u0__abc_49347_n4540) );
  AND2X2 AND2X2_1263 ( .A(u0__abc_49347_n4545), .B(u0__abc_49347_n4546), .Y(u0__abc_49347_n4547) );
  AND2X2 AND2X2_1264 ( .A(u0__abc_49347_n4549), .B(u0__abc_49347_n4548), .Y(u0__abc_49347_n4550) );
  AND2X2 AND2X2_1265 ( .A(u0__abc_49347_n4547), .B(u0__abc_49347_n4550), .Y(u0__abc_49347_n4551) );
  AND2X2 AND2X2_1266 ( .A(u0__abc_49347_n4552), .B(u0__abc_49347_n4553), .Y(u0__abc_49347_n4554) );
  AND2X2 AND2X2_1267 ( .A(u0__abc_49347_n4555), .B(u0__abc_49347_n4556), .Y(u0__abc_49347_n4557) );
  AND2X2 AND2X2_1268 ( .A(u0__abc_49347_n4557), .B(u0__abc_49347_n4554), .Y(u0__abc_49347_n4558) );
  AND2X2 AND2X2_1269 ( .A(u0__abc_49347_n4558), .B(u0__abc_49347_n4551), .Y(u0__abc_49347_n4559) );
  AND2X2 AND2X2_127 ( .A(u0__abc_49347_n1220), .B(u0__abc_49347_n1179_bF_buf4), .Y(u0__abc_49347_n1221) );
  AND2X2 AND2X2_1270 ( .A(u0__abc_49347_n4506), .B(u0__abc_49347_n4513), .Y(u0__abc_49347_n4560) );
  AND2X2 AND2X2_1271 ( .A(u0__abc_49347_n4525), .B(u0__abc_49347_n4530), .Y(u0__abc_49347_n4562) );
  AND2X2 AND2X2_1272 ( .A(u0__abc_49347_n4561), .B(u0__abc_49347_n4563), .Y(u0__abc_49347_n4564) );
  AND2X2 AND2X2_1273 ( .A(u0__abc_49347_n4525), .B(u0__abc_49347_n4501), .Y(u0__abc_49347_n4565) );
  AND2X2 AND2X2_1274 ( .A(u0__abc_49347_n4510), .B(u0__abc_49347_n4530), .Y(u0__abc_49347_n4567) );
  AND2X2 AND2X2_1275 ( .A(u0__abc_49347_n4566), .B(u0__abc_49347_n4568), .Y(u0__abc_49347_n4569) );
  AND2X2 AND2X2_1276 ( .A(u0__abc_49347_n4569), .B(u0__abc_49347_n4564), .Y(u0__abc_49347_n4570) );
  AND2X2 AND2X2_1277 ( .A(u0__abc_49347_n4515), .B(u0__abc_49347_n4530), .Y(u0__abc_49347_n4571) );
  AND2X2 AND2X2_1278 ( .A(u0__abc_49347_n4501), .B(\wb_addr_i[6] ), .Y(u0__abc_49347_n4573) );
  AND2X2 AND2X2_1279 ( .A(u0__abc_49347_n4575), .B(u0__abc_49347_n4572), .Y(u0__abc_49347_n4576) );
  AND2X2 AND2X2_128 ( .A(spec_req_cs_2_bF_buf1), .B(u0_tms2_1_), .Y(u0__abc_49347_n1222) );
  AND2X2 AND2X2_1280 ( .A(u0__abc_49347_n4577), .B(u0__abc_49347_n4578), .Y(u0__abc_49347_n4579) );
  AND2X2 AND2X2_1281 ( .A(u0__abc_49347_n4576), .B(u0__abc_49347_n4579), .Y(u0__abc_49347_n4580) );
  AND2X2 AND2X2_1282 ( .A(u0__abc_49347_n4580), .B(u0__abc_49347_n4570), .Y(u0__abc_49347_n4581) );
  AND2X2 AND2X2_1283 ( .A(u0__abc_49347_n4581), .B(u0__abc_49347_n4559), .Y(u0__abc_49347_n4582) );
  AND2X2 AND2X2_1284 ( .A(u0__abc_49347_n4582_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n4583) );
  AND2X2 AND2X2_1285 ( .A(u0__abc_49347_n4573), .B(u0__abc_49347_n4524), .Y(u0__abc_49347_n4584) );
  AND2X2 AND2X2_1286 ( .A(u0__abc_49347_n4584_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n4585) );
  AND2X2 AND2X2_1287 ( .A(u0__abc_49347_n4573), .B(u0__abc_49347_n4509), .Y(u0__abc_49347_n4586) );
  AND2X2 AND2X2_1288 ( .A(u0__abc_49347_n4586_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n4587) );
  AND2X2 AND2X2_1289 ( .A(u0__abc_49347_n4571_bF_buf3), .B(u0_tms5_0_), .Y(u0__abc_49347_n4588) );
  AND2X2 AND2X2_129 ( .A(u0__abc_49347_n1223), .B(u0__abc_49347_n1178_1_bF_buf4), .Y(u0__abc_49347_n1224) );
  AND2X2 AND2X2_1290 ( .A(u0__abc_49347_n4573), .B(u0__abc_49347_n4505), .Y(u0__abc_49347_n4589) );
  AND2X2 AND2X2_1291 ( .A(u0__abc_49347_n4589_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n4590) );
  AND2X2 AND2X2_1292 ( .A(u0__abc_49347_n4565), .B(u0_csc_mask_0_), .Y(u0__abc_49347_n4594) );
  AND2X2 AND2X2_1293 ( .A(u0__abc_49347_n4560_bF_buf3), .B(u0_csc0_0_), .Y(u0__abc_49347_n4595) );
  AND2X2 AND2X2_1294 ( .A(u0__abc_49347_n4562_bF_buf3), .B(u0_csc5_0_), .Y(u0__abc_49347_n4597) );
  AND2X2 AND2X2_1295 ( .A(u0__abc_49347_n4567_bF_buf3), .B(u0_tms4_0_), .Y(u0__abc_49347_n4598) );
  AND2X2 AND2X2_1296 ( .A(u0__abc_49347_n4526_bF_buf2), .B(u0_csc1_1_), .Y(u0__abc_49347_n4604) );
  AND2X2 AND2X2_1297 ( .A(u0__abc_49347_n4531_bF_buf2), .B(u0_csc4_1_), .Y(u0__abc_49347_n4605) );
  AND2X2 AND2X2_1298 ( .A(u0__abc_49347_n4528_bF_buf2), .B(u0_tms3_1_), .Y(u0__abc_49347_n4606) );
  AND2X2 AND2X2_1299 ( .A(u0__abc_49347_n4535_bF_buf2), .B(u0_tms0_1_), .Y(u0__abc_49347_n4609) );
  AND2X2 AND2X2_13 ( .A(_abc_55805_n275), .B(_abc_55805_n276), .Y(obct_cs_5_) );
  AND2X2 AND2X2_130 ( .A(spec_req_cs_1_bF_buf1), .B(u0_tms1_1_), .Y(u0__abc_49347_n1225) );
  AND2X2 AND2X2_1300 ( .A(u0__abc_49347_n4539_bF_buf2), .B(u0_csc3_1_), .Y(u0__abc_49347_n4610) );
  AND2X2 AND2X2_1301 ( .A(u0__abc_49347_n4537_bF_buf2), .B(u0_tms2_1_), .Y(u0__abc_49347_n4611) );
  AND2X2 AND2X2_1302 ( .A(u0__abc_49347_n4562_bF_buf2), .B(u0_csc5_1_), .Y(u0__abc_49347_n4615) );
  AND2X2 AND2X2_1303 ( .A(u0__abc_49347_n4560_bF_buf2), .B(u0_csc0_1_), .Y(u0__abc_49347_n4616) );
  AND2X2 AND2X2_1304 ( .A(u0__abc_49347_n4565), .B(u0_csc_mask_1_), .Y(u0__abc_49347_n4617) );
  AND2X2 AND2X2_1305 ( .A(u0__abc_49347_n4582_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n4621) );
  AND2X2 AND2X2_1306 ( .A(u0__abc_49347_n4586_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n4622) );
  AND2X2 AND2X2_1307 ( .A(u0__abc_49347_n4584_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n4623) );
  AND2X2 AND2X2_1308 ( .A(u0__abc_49347_n4571_bF_buf2), .B(u0_tms5_1_), .Y(u0__abc_49347_n4624) );
  AND2X2 AND2X2_1309 ( .A(u0__abc_49347_n4589_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n4625) );
  AND2X2 AND2X2_131 ( .A(u0__abc_49347_n1175_bF_buf4), .B(u0__abc_49347_n1228_1), .Y(u0__abc_49347_n1229) );
  AND2X2 AND2X2_1310 ( .A(u0__abc_49347_n4507_bF_buf1), .B(_auto_iopadmap_cc_313_execute_56315), .Y(u0__abc_49347_n4629) );
  AND2X2 AND2X2_1311 ( .A(u0__abc_49347_n4519_bF_buf2), .B(u0_csc2_1_), .Y(u0__abc_49347_n4630) );
  AND2X2 AND2X2_1312 ( .A(u0__abc_49347_n4516_bF_buf2), .B(u0_tms1_1_), .Y(u0__abc_49347_n4631) );
  AND2X2 AND2X2_1313 ( .A(u0__abc_49347_n4511_bF_buf2), .B(_auto_iopadmap_cc_313_execute_56321_1_), .Y(u0__abc_49347_n4634) );
  AND2X2 AND2X2_1314 ( .A(u0__abc_49347_n4567_bF_buf2), .B(u0_tms4_1_), .Y(u0__abc_49347_n4635) );
  AND2X2 AND2X2_1315 ( .A(u0__abc_49347_n4507_bF_buf0), .B(fs), .Y(u0__abc_49347_n4641) );
  AND2X2 AND2X2_1316 ( .A(u0__abc_49347_n4511_bF_buf1), .B(_auto_iopadmap_cc_313_execute_56321_2_), .Y(u0__abc_49347_n4642) );
  AND2X2 AND2X2_1317 ( .A(u0__abc_49347_n4516_bF_buf1), .B(u0_tms1_2_), .Y(u0__abc_49347_n4643) );
  AND2X2 AND2X2_1318 ( .A(u0__abc_49347_n4519_bF_buf1), .B(u0_csc2_2_), .Y(u0__abc_49347_n4644) );
  AND2X2 AND2X2_1319 ( .A(u0__abc_49347_n4535_bF_buf1), .B(u0_tms0_2_), .Y(u0__abc_49347_n4648) );
  AND2X2 AND2X2_132 ( .A(u0__abc_49347_n1227_1), .B(u0__abc_49347_n1229), .Y(u0__abc_49347_n1230) );
  AND2X2 AND2X2_1320 ( .A(u0__abc_49347_n4528_bF_buf1), .B(u0_tms3_2_), .Y(u0__abc_49347_n4649) );
  AND2X2 AND2X2_1321 ( .A(u0__abc_49347_n4531_bF_buf1), .B(u0_csc4_2_), .Y(u0__abc_49347_n4650) );
  AND2X2 AND2X2_1322 ( .A(u0__abc_49347_n4526_bF_buf1), .B(u0_csc1_2_), .Y(u0__abc_49347_n4653) );
  AND2X2 AND2X2_1323 ( .A(u0__abc_49347_n4539_bF_buf1), .B(u0_csc3_2_), .Y(u0__abc_49347_n4654) );
  AND2X2 AND2X2_1324 ( .A(u0__abc_49347_n4537_bF_buf1), .B(u0_tms2_2_), .Y(u0__abc_49347_n4655) );
  AND2X2 AND2X2_1325 ( .A(u0__abc_49347_n4582_bF_buf2), .B(1'b0), .Y(u0__abc_49347_n4660) );
  AND2X2 AND2X2_1326 ( .A(u0__abc_49347_n4586_bF_buf2), .B(1'b0), .Y(u0__abc_49347_n4661) );
  AND2X2 AND2X2_1327 ( .A(u0__abc_49347_n4584_bF_buf2), .B(1'b0), .Y(u0__abc_49347_n4662) );
  AND2X2 AND2X2_1328 ( .A(u0__abc_49347_n4571_bF_buf1), .B(u0_tms5_2_), .Y(u0__abc_49347_n4663) );
  AND2X2 AND2X2_1329 ( .A(u0__abc_49347_n4589_bF_buf2), .B(1'b0), .Y(u0__abc_49347_n4664) );
  AND2X2 AND2X2_133 ( .A(u0__abc_49347_n1176_1_bF_buf4), .B(sp_tms_2_), .Y(u0__abc_49347_n1232) );
  AND2X2 AND2X2_1330 ( .A(u0__abc_49347_n4565), .B(u0_csc_mask_2_), .Y(u0__abc_49347_n4668) );
  AND2X2 AND2X2_1331 ( .A(u0__abc_49347_n4560_bF_buf1), .B(u0_csc0_2_), .Y(u0__abc_49347_n4669) );
  AND2X2 AND2X2_1332 ( .A(u0__abc_49347_n4567_bF_buf1), .B(u0_tms4_2_), .Y(u0__abc_49347_n4671) );
  AND2X2 AND2X2_1333 ( .A(u0__abc_49347_n4562_bF_buf1), .B(u0_csc5_2_), .Y(u0__abc_49347_n4672) );
  AND2X2 AND2X2_1334 ( .A(u0__abc_49347_n4511_bF_buf0), .B(_auto_iopadmap_cc_313_execute_56321_3_), .Y(u0__abc_49347_n4678) );
  AND2X2 AND2X2_1335 ( .A(u0__abc_49347_n4507_bF_buf3), .B(u0_csr_3_), .Y(u0__abc_49347_n4679) );
  AND2X2 AND2X2_1336 ( .A(u0__abc_49347_n4516_bF_buf0), .B(u0_tms1_3_), .Y(u0__abc_49347_n4680) );
  AND2X2 AND2X2_1337 ( .A(u0__abc_49347_n4519_bF_buf0), .B(u0_csc2_3_), .Y(u0__abc_49347_n4681) );
  AND2X2 AND2X2_1338 ( .A(u0__abc_49347_n4535_bF_buf0), .B(u0_tms0_3_), .Y(u0__abc_49347_n4685) );
  AND2X2 AND2X2_1339 ( .A(u0__abc_49347_n4528_bF_buf0), .B(u0_tms3_3_), .Y(u0__abc_49347_n4686) );
  AND2X2 AND2X2_134 ( .A(spec_req_cs_5_bF_buf0), .B(u0_tms5_2_), .Y(u0__abc_49347_n1233) );
  AND2X2 AND2X2_1340 ( .A(u0__abc_49347_n4531_bF_buf0), .B(u0_csc4_3_), .Y(u0__abc_49347_n4687) );
  AND2X2 AND2X2_1341 ( .A(u0__abc_49347_n4526_bF_buf0), .B(u0_csc1_3_), .Y(u0__abc_49347_n4690) );
  AND2X2 AND2X2_1342 ( .A(u0__abc_49347_n4539_bF_buf0), .B(u0_csc3_3_), .Y(u0__abc_49347_n4691) );
  AND2X2 AND2X2_1343 ( .A(u0__abc_49347_n4537_bF_buf0), .B(u0_tms2_3_), .Y(u0__abc_49347_n4692) );
  AND2X2 AND2X2_1344 ( .A(u0__abc_49347_n4582_bF_buf1), .B(1'b0), .Y(u0__abc_49347_n4697) );
  AND2X2 AND2X2_1345 ( .A(u0__abc_49347_n4586_bF_buf1), .B(1'b0), .Y(u0__abc_49347_n4698) );
  AND2X2 AND2X2_1346 ( .A(u0__abc_49347_n4584_bF_buf1), .B(1'b0), .Y(u0__abc_49347_n4699) );
  AND2X2 AND2X2_1347 ( .A(u0__abc_49347_n4571_bF_buf0), .B(u0_tms5_3_), .Y(u0__abc_49347_n4700) );
  AND2X2 AND2X2_1348 ( .A(u0__abc_49347_n4589_bF_buf1), .B(1'b0), .Y(u0__abc_49347_n4701) );
  AND2X2 AND2X2_1349 ( .A(u0__abc_49347_n4560_bF_buf0), .B(u0_csc0_3_), .Y(u0__abc_49347_n4705) );
  AND2X2 AND2X2_135 ( .A(u0__abc_49347_n1235), .B(u0__abc_49347_n1185_bF_buf3), .Y(u0__abc_49347_n1236_1) );
  AND2X2 AND2X2_1350 ( .A(u0__abc_49347_n4565), .B(u0_csc_mask_3_), .Y(u0__abc_49347_n4706) );
  AND2X2 AND2X2_1351 ( .A(u0__abc_49347_n4562_bF_buf0), .B(u0_csc5_3_), .Y(u0__abc_49347_n4708) );
  AND2X2 AND2X2_1352 ( .A(u0__abc_49347_n4567_bF_buf0), .B(u0_tms4_3_), .Y(u0__abc_49347_n4709) );
  AND2X2 AND2X2_1353 ( .A(u0__abc_49347_n4526_bF_buf4), .B(u0_csc1_4_), .Y(u0__abc_49347_n4715) );
  AND2X2 AND2X2_1354 ( .A(u0__abc_49347_n4531_bF_buf4), .B(u0_csc4_4_), .Y(u0__abc_49347_n4716) );
  AND2X2 AND2X2_1355 ( .A(u0__abc_49347_n4528_bF_buf4), .B(u0_tms3_4_), .Y(u0__abc_49347_n4717) );
  AND2X2 AND2X2_1356 ( .A(u0__abc_49347_n4535_bF_buf4), .B(u0_tms0_4_), .Y(u0__abc_49347_n4720) );
  AND2X2 AND2X2_1357 ( .A(u0__abc_49347_n4537_bF_buf4), .B(u0_tms2_4_), .Y(u0__abc_49347_n4721) );
  AND2X2 AND2X2_1358 ( .A(u0__abc_49347_n4539_bF_buf4), .B(u0_csc3_4_), .Y(u0__abc_49347_n4722) );
  AND2X2 AND2X2_1359 ( .A(u0__abc_49347_n4567_bF_buf4), .B(u0_tms4_4_), .Y(u0__abc_49347_n4726) );
  AND2X2 AND2X2_136 ( .A(u0__abc_49347_n1236_1), .B(u0__abc_49347_n1234), .Y(u0__abc_49347_n1237_1) );
  AND2X2 AND2X2_1360 ( .A(u0__abc_49347_n4560_bF_buf4), .B(u0_csc0_4_), .Y(u0__abc_49347_n4727) );
  AND2X2 AND2X2_1361 ( .A(u0__abc_49347_n4565), .B(u0_csc_mask_4_), .Y(u0__abc_49347_n4728) );
  AND2X2 AND2X2_1362 ( .A(u0__abc_49347_n4582_bF_buf0), .B(1'b0), .Y(u0__abc_49347_n4732) );
  AND2X2 AND2X2_1363 ( .A(u0__abc_49347_n4586_bF_buf0), .B(1'b0), .Y(u0__abc_49347_n4733) );
  AND2X2 AND2X2_1364 ( .A(u0__abc_49347_n4584_bF_buf0), .B(1'b0), .Y(u0__abc_49347_n4734) );
  AND2X2 AND2X2_1365 ( .A(u0__abc_49347_n4571_bF_buf4), .B(u0_tms5_4_), .Y(u0__abc_49347_n4735) );
  AND2X2 AND2X2_1366 ( .A(u0__abc_49347_n4589_bF_buf0), .B(1'b0), .Y(u0__abc_49347_n4736) );
  AND2X2 AND2X2_1367 ( .A(u0__abc_49347_n4511_bF_buf4), .B(_auto_iopadmap_cc_313_execute_56321_4_), .Y(u0__abc_49347_n4740) );
  AND2X2 AND2X2_1368 ( .A(u0__abc_49347_n4516_bF_buf4), .B(u0_tms1_4_), .Y(u0__abc_49347_n4741) );
  AND2X2 AND2X2_1369 ( .A(u0__abc_49347_n4519_bF_buf4), .B(u0_csc2_4_), .Y(u0__abc_49347_n4742) );
  AND2X2 AND2X2_137 ( .A(u0__abc_49347_n1238), .B(u0__abc_49347_n1181_bF_buf3), .Y(u0__abc_49347_n1239) );
  AND2X2 AND2X2_1370 ( .A(u0__abc_49347_n4507_bF_buf2), .B(u0_csr_4_), .Y(u0__abc_49347_n4745) );
  AND2X2 AND2X2_1371 ( .A(u0__abc_49347_n4562_bF_buf4), .B(u0_csc5_4_), .Y(u0__abc_49347_n4746) );
  AND2X2 AND2X2_1372 ( .A(u0__abc_49347_n4526_bF_buf3), .B(u0_csc1_5_), .Y(u0__abc_49347_n4752) );
  AND2X2 AND2X2_1373 ( .A(u0__abc_49347_n4531_bF_buf3), .B(u0_csc4_5_), .Y(u0__abc_49347_n4753) );
  AND2X2 AND2X2_1374 ( .A(u0__abc_49347_n4528_bF_buf3), .B(u0_tms3_5_), .Y(u0__abc_49347_n4754) );
  AND2X2 AND2X2_1375 ( .A(u0__abc_49347_n4535_bF_buf3), .B(u0_tms0_5_), .Y(u0__abc_49347_n4757) );
  AND2X2 AND2X2_1376 ( .A(u0__abc_49347_n4539_bF_buf3), .B(u0_csc3_5_), .Y(u0__abc_49347_n4758) );
  AND2X2 AND2X2_1377 ( .A(u0__abc_49347_n4537_bF_buf3), .B(u0_tms2_5_), .Y(u0__abc_49347_n4759) );
  AND2X2 AND2X2_1378 ( .A(u0__abc_49347_n4562_bF_buf3), .B(u0_csc5_5_), .Y(u0__abc_49347_n4763) );
  AND2X2 AND2X2_1379 ( .A(u0__abc_49347_n4560_bF_buf3), .B(u0_csc0_5_), .Y(u0__abc_49347_n4764) );
  AND2X2 AND2X2_138 ( .A(spec_req_cs_4_bF_buf0), .B(u0_tms4_2_), .Y(u0__abc_49347_n1240) );
  AND2X2 AND2X2_1380 ( .A(u0__abc_49347_n4565), .B(u0_csc_mask_5_), .Y(u0__abc_49347_n4765) );
  AND2X2 AND2X2_1381 ( .A(u0__abc_49347_n4582_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n4769) );
  AND2X2 AND2X2_1382 ( .A(u0__abc_49347_n4584_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n4770) );
  AND2X2 AND2X2_1383 ( .A(u0__abc_49347_n4586_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n4771) );
  AND2X2 AND2X2_1384 ( .A(u0__abc_49347_n4571_bF_buf3), .B(u0_tms5_5_), .Y(u0__abc_49347_n4772) );
  AND2X2 AND2X2_1385 ( .A(u0__abc_49347_n4589_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n4773) );
  AND2X2 AND2X2_1386 ( .A(u0__abc_49347_n4507_bF_buf1), .B(u0_csr_5_), .Y(u0__abc_49347_n4777) );
  AND2X2 AND2X2_1387 ( .A(u0__abc_49347_n4519_bF_buf3), .B(u0_csc2_5_), .Y(u0__abc_49347_n4778) );
  AND2X2 AND2X2_1388 ( .A(u0__abc_49347_n4516_bF_buf3), .B(u0_tms1_5_), .Y(u0__abc_49347_n4779) );
  AND2X2 AND2X2_1389 ( .A(u0__abc_49347_n4567_bF_buf3), .B(u0_tms4_5_), .Y(u0__abc_49347_n4782) );
  AND2X2 AND2X2_139 ( .A(u0__abc_49347_n1241), .B(u0__abc_49347_n1180_1_bF_buf3), .Y(u0__abc_49347_n1242) );
  AND2X2 AND2X2_1390 ( .A(u0__abc_49347_n4511_bF_buf3), .B(_auto_iopadmap_cc_313_execute_56321_5_), .Y(u0__abc_49347_n4783) );
  AND2X2 AND2X2_1391 ( .A(u0__abc_49347_n4535_bF_buf2), .B(u0_tms0_6_), .Y(u0__abc_49347_n4789) );
  AND2X2 AND2X2_1392 ( .A(u0__abc_49347_n4531_bF_buf2), .B(u0_csc4_6_), .Y(u0__abc_49347_n4790) );
  AND2X2 AND2X2_1393 ( .A(u0__abc_49347_n4528_bF_buf2), .B(u0_tms3_6_), .Y(u0__abc_49347_n4791) );
  AND2X2 AND2X2_1394 ( .A(u0__abc_49347_n4526_bF_buf2), .B(u0_csc1_6_), .Y(u0__abc_49347_n4794) );
  AND2X2 AND2X2_1395 ( .A(u0__abc_49347_n4537_bF_buf2), .B(u0_tms2_6_), .Y(u0__abc_49347_n4795) );
  AND2X2 AND2X2_1396 ( .A(u0__abc_49347_n4539_bF_buf2), .B(u0_csc3_6_), .Y(u0__abc_49347_n4796) );
  AND2X2 AND2X2_1397 ( .A(u0__abc_49347_n4567_bF_buf2), .B(u0_tms4_6_), .Y(u0__abc_49347_n4800) );
  AND2X2 AND2X2_1398 ( .A(u0__abc_49347_n4560_bF_buf2), .B(u0_csc0_6_), .Y(u0__abc_49347_n4801) );
  AND2X2 AND2X2_1399 ( .A(u0__abc_49347_n4565), .B(u0_csc_mask_6_), .Y(u0__abc_49347_n4802) );
  AND2X2 AND2X2_14 ( .A(_abc_55805_n278), .B(_abc_55805_n279), .Y(_abc_55805_n280) );
  AND2X2 AND2X2_140 ( .A(spec_req_cs_3_bF_buf0), .B(u0_tms3_2_), .Y(u0__abc_49347_n1243) );
  AND2X2 AND2X2_1400 ( .A(u0__abc_49347_n4582_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n4806) );
  AND2X2 AND2X2_1401 ( .A(u0__abc_49347_n4586_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n4807) );
  AND2X2 AND2X2_1402 ( .A(u0__abc_49347_n4584_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n4808) );
  AND2X2 AND2X2_1403 ( .A(u0__abc_49347_n4571_bF_buf2), .B(u0_tms5_6_), .Y(u0__abc_49347_n4809) );
  AND2X2 AND2X2_1404 ( .A(u0__abc_49347_n4589_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n4810) );
  AND2X2 AND2X2_1405 ( .A(u0__abc_49347_n4511_bF_buf2), .B(_auto_iopadmap_cc_313_execute_56321_6_), .Y(u0__abc_49347_n4814) );
  AND2X2 AND2X2_1406 ( .A(u0__abc_49347_n4516_bF_buf2), .B(u0_tms1_6_), .Y(u0__abc_49347_n4815) );
  AND2X2 AND2X2_1407 ( .A(u0__abc_49347_n4519_bF_buf2), .B(u0_csc2_6_), .Y(u0__abc_49347_n4816) );
  AND2X2 AND2X2_1408 ( .A(u0__abc_49347_n4562_bF_buf2), .B(u0_csc5_6_), .Y(u0__abc_49347_n4819) );
  AND2X2 AND2X2_1409 ( .A(u0__abc_49347_n4507_bF_buf0), .B(u0_csr_6_), .Y(u0__abc_49347_n4820) );
  AND2X2 AND2X2_141 ( .A(u0__abc_49347_n1244), .B(u0__abc_49347_n1179_bF_buf3), .Y(u0__abc_49347_n1245_1) );
  AND2X2 AND2X2_1410 ( .A(u0__abc_49347_n4526_bF_buf1), .B(u0_csc1_7_), .Y(u0__abc_49347_n4826) );
  AND2X2 AND2X2_1411 ( .A(u0__abc_49347_n4531_bF_buf1), .B(u0_csc4_7_), .Y(u0__abc_49347_n4827) );
  AND2X2 AND2X2_1412 ( .A(u0__abc_49347_n4528_bF_buf1), .B(u0_tms3_7_), .Y(u0__abc_49347_n4828) );
  AND2X2 AND2X2_1413 ( .A(u0__abc_49347_n4535_bF_buf1), .B(u0_tms0_7_), .Y(u0__abc_49347_n4831) );
  AND2X2 AND2X2_1414 ( .A(u0__abc_49347_n4539_bF_buf1), .B(u0_csc3_7_), .Y(u0__abc_49347_n4832) );
  AND2X2 AND2X2_1415 ( .A(u0__abc_49347_n4537_bF_buf1), .B(u0_tms2_7_), .Y(u0__abc_49347_n4833) );
  AND2X2 AND2X2_1416 ( .A(u0__abc_49347_n4562_bF_buf1), .B(u0_csc5_7_), .Y(u0__abc_49347_n4837) );
  AND2X2 AND2X2_1417 ( .A(u0__abc_49347_n4560_bF_buf1), .B(u0_csc0_7_), .Y(u0__abc_49347_n4838) );
  AND2X2 AND2X2_1418 ( .A(u0__abc_49347_n4565), .B(u0_csc_mask_7_), .Y(u0__abc_49347_n4839) );
  AND2X2 AND2X2_1419 ( .A(u0__abc_49347_n4582_bF_buf2), .B(1'b0), .Y(u0__abc_49347_n4843) );
  AND2X2 AND2X2_142 ( .A(spec_req_cs_2_bF_buf0), .B(u0_tms2_2_), .Y(u0__abc_49347_n1246_1) );
  AND2X2 AND2X2_1420 ( .A(u0__abc_49347_n4584_bF_buf2), .B(1'b0), .Y(u0__abc_49347_n4844) );
  AND2X2 AND2X2_1421 ( .A(u0__abc_49347_n4586_bF_buf2), .B(1'b0), .Y(u0__abc_49347_n4845) );
  AND2X2 AND2X2_1422 ( .A(u0__abc_49347_n4571_bF_buf1), .B(u0_tms5_7_), .Y(u0__abc_49347_n4846) );
  AND2X2 AND2X2_1423 ( .A(u0__abc_49347_n4589_bF_buf2), .B(1'b0), .Y(u0__abc_49347_n4847) );
  AND2X2 AND2X2_1424 ( .A(u0__abc_49347_n4511_bF_buf1), .B(_auto_iopadmap_cc_313_execute_56321_7_), .Y(u0__abc_49347_n4851) );
  AND2X2 AND2X2_1425 ( .A(u0__abc_49347_n4519_bF_buf1), .B(u0_csc2_7_), .Y(u0__abc_49347_n4852) );
  AND2X2 AND2X2_1426 ( .A(u0__abc_49347_n4516_bF_buf1), .B(u0_tms1_7_), .Y(u0__abc_49347_n4853) );
  AND2X2 AND2X2_1427 ( .A(u0__abc_49347_n4567_bF_buf1), .B(u0_tms4_7_), .Y(u0__abc_49347_n4856) );
  AND2X2 AND2X2_1428 ( .A(u0__abc_49347_n4507_bF_buf3), .B(u0_csr_7_), .Y(u0__abc_49347_n4857) );
  AND2X2 AND2X2_1429 ( .A(u0__abc_49347_n4535_bF_buf0), .B(u0_tms0_8_), .Y(u0__abc_49347_n4863) );
  AND2X2 AND2X2_143 ( .A(u0__abc_49347_n1247), .B(u0__abc_49347_n1178_1_bF_buf3), .Y(u0__abc_49347_n1248) );
  AND2X2 AND2X2_1430 ( .A(u0__abc_49347_n4531_bF_buf0), .B(u0_csc4_8_), .Y(u0__abc_49347_n4864) );
  AND2X2 AND2X2_1431 ( .A(u0__abc_49347_n4528_bF_buf0), .B(u0_tms3_8_), .Y(u0__abc_49347_n4865) );
  AND2X2 AND2X2_1432 ( .A(u0__abc_49347_n4526_bF_buf0), .B(u0_csc1_8_), .Y(u0__abc_49347_n4868) );
  AND2X2 AND2X2_1433 ( .A(u0__abc_49347_n4537_bF_buf0), .B(u0_tms2_8_), .Y(u0__abc_49347_n4869) );
  AND2X2 AND2X2_1434 ( .A(u0__abc_49347_n4539_bF_buf0), .B(u0_csc3_8_), .Y(u0__abc_49347_n4870) );
  AND2X2 AND2X2_1435 ( .A(u0__abc_49347_n4562_bF_buf0), .B(u0_csc5_8_), .Y(u0__abc_49347_n4874) );
  AND2X2 AND2X2_1436 ( .A(u0__abc_49347_n4560_bF_buf0), .B(u0_csc0_8_), .Y(u0__abc_49347_n4875) );
  AND2X2 AND2X2_1437 ( .A(u0__abc_49347_n4565), .B(u0_csc_mask_8_), .Y(u0__abc_49347_n4876) );
  AND2X2 AND2X2_1438 ( .A(u0__abc_49347_n4582_bF_buf1), .B(1'b0), .Y(u0__abc_49347_n4880) );
  AND2X2 AND2X2_1439 ( .A(u0__abc_49347_n4586_bF_buf1), .B(1'b0), .Y(u0__abc_49347_n4881) );
  AND2X2 AND2X2_144 ( .A(spec_req_cs_1_bF_buf0), .B(u0_tms1_2_), .Y(u0__abc_49347_n1249) );
  AND2X2 AND2X2_1440 ( .A(u0__abc_49347_n4584_bF_buf1), .B(1'b0), .Y(u0__abc_49347_n4882) );
  AND2X2 AND2X2_1441 ( .A(u0__abc_49347_n4571_bF_buf0), .B(u0_tms5_8_), .Y(u0__abc_49347_n4883) );
  AND2X2 AND2X2_1442 ( .A(u0__abc_49347_n4589_bF_buf1), .B(1'b0), .Y(u0__abc_49347_n4884) );
  AND2X2 AND2X2_1443 ( .A(u0__abc_49347_n4507_bF_buf2), .B(ref_int_0_), .Y(u0__abc_49347_n4888) );
  AND2X2 AND2X2_1444 ( .A(u0__abc_49347_n4519_bF_buf0), .B(u0_csc2_8_), .Y(u0__abc_49347_n4889) );
  AND2X2 AND2X2_1445 ( .A(u0__abc_49347_n4516_bF_buf0), .B(u0_tms1_8_), .Y(u0__abc_49347_n4890) );
  AND2X2 AND2X2_1446 ( .A(u0__abc_49347_n4511_bF_buf0), .B(_auto_iopadmap_cc_313_execute_56321_8_), .Y(u0__abc_49347_n4893) );
  AND2X2 AND2X2_1447 ( .A(u0__abc_49347_n4567_bF_buf0), .B(u0_tms4_8_), .Y(u0__abc_49347_n4894) );
  AND2X2 AND2X2_1448 ( .A(u0__abc_49347_n4535_bF_buf4), .B(u0_tms0_9_), .Y(u0__abc_49347_n4900) );
  AND2X2 AND2X2_1449 ( .A(u0__abc_49347_n4531_bF_buf4), .B(u0_csc4_9_), .Y(u0__abc_49347_n4901) );
  AND2X2 AND2X2_145 ( .A(u0__abc_49347_n1175_bF_buf3), .B(u0__abc_49347_n1252), .Y(u0__abc_49347_n1253) );
  AND2X2 AND2X2_1450 ( .A(u0__abc_49347_n4528_bF_buf4), .B(u0_tms3_9_), .Y(u0__abc_49347_n4902) );
  AND2X2 AND2X2_1451 ( .A(u0__abc_49347_n4526_bF_buf4), .B(u0_csc1_9_), .Y(u0__abc_49347_n4905) );
  AND2X2 AND2X2_1452 ( .A(u0__abc_49347_n4539_bF_buf4), .B(u0_csc3_9_), .Y(u0__abc_49347_n4906) );
  AND2X2 AND2X2_1453 ( .A(u0__abc_49347_n4537_bF_buf4), .B(u0_tms2_9_), .Y(u0__abc_49347_n4907) );
  AND2X2 AND2X2_1454 ( .A(u0__abc_49347_n4562_bF_buf4), .B(u0_csc5_9_), .Y(u0__abc_49347_n4911) );
  AND2X2 AND2X2_1455 ( .A(u0__abc_49347_n4565), .B(u0_csc_mask_9_), .Y(u0__abc_49347_n4912) );
  AND2X2 AND2X2_1456 ( .A(u0__abc_49347_n4560_bF_buf4), .B(u0_csc0_9_), .Y(u0__abc_49347_n4913) );
  AND2X2 AND2X2_1457 ( .A(u0__abc_49347_n4582_bF_buf0), .B(1'b0), .Y(u0__abc_49347_n4917) );
  AND2X2 AND2X2_1458 ( .A(u0__abc_49347_n4586_bF_buf0), .B(1'b0), .Y(u0__abc_49347_n4918) );
  AND2X2 AND2X2_1459 ( .A(u0__abc_49347_n4584_bF_buf0), .B(1'b0), .Y(u0__abc_49347_n4919) );
  AND2X2 AND2X2_146 ( .A(u0__abc_49347_n1251), .B(u0__abc_49347_n1253), .Y(u0__abc_49347_n1254_1) );
  AND2X2 AND2X2_1460 ( .A(u0__abc_49347_n4571_bF_buf4), .B(u0_tms5_9_), .Y(u0__abc_49347_n4920) );
  AND2X2 AND2X2_1461 ( .A(u0__abc_49347_n4589_bF_buf0), .B(1'b0), .Y(u0__abc_49347_n4921) );
  AND2X2 AND2X2_1462 ( .A(u0__abc_49347_n4511_bF_buf4), .B(_auto_iopadmap_cc_313_execute_56321_9_), .Y(u0__abc_49347_n4925) );
  AND2X2 AND2X2_1463 ( .A(u0__abc_49347_n4516_bF_buf4), .B(u0_tms1_9_), .Y(u0__abc_49347_n4926) );
  AND2X2 AND2X2_1464 ( .A(u0__abc_49347_n4519_bF_buf4), .B(u0_csc2_9_), .Y(u0__abc_49347_n4927) );
  AND2X2 AND2X2_1465 ( .A(u0__abc_49347_n4507_bF_buf1), .B(ref_int_1_), .Y(u0__abc_49347_n4930) );
  AND2X2 AND2X2_1466 ( .A(u0__abc_49347_n4567_bF_buf4), .B(u0_tms4_9_), .Y(u0__abc_49347_n4931) );
  AND2X2 AND2X2_1467 ( .A(u0__abc_49347_n4511_bF_buf3), .B(_auto_iopadmap_cc_313_execute_56321_10_), .Y(u0__abc_49347_n4937) );
  AND2X2 AND2X2_1468 ( .A(u0__abc_49347_n4507_bF_buf0), .B(ref_int_2_), .Y(u0__abc_49347_n4938) );
  AND2X2 AND2X2_1469 ( .A(u0__abc_49347_n4516_bF_buf3), .B(u0_tms1_10_), .Y(u0__abc_49347_n4939) );
  AND2X2 AND2X2_147 ( .A(u0__abc_49347_n1176_1_bF_buf3), .B(sp_tms_3_), .Y(u0__abc_49347_n1256) );
  AND2X2 AND2X2_1470 ( .A(u0__abc_49347_n4519_bF_buf3), .B(u0_csc2_10_), .Y(u0__abc_49347_n4940) );
  AND2X2 AND2X2_1471 ( .A(u0__abc_49347_n4526_bF_buf3), .B(u0_csc1_10_), .Y(u0__abc_49347_n4944) );
  AND2X2 AND2X2_1472 ( .A(u0__abc_49347_n4528_bF_buf3), .B(u0_tms3_10_), .Y(u0__abc_49347_n4945) );
  AND2X2 AND2X2_1473 ( .A(u0__abc_49347_n4531_bF_buf3), .B(u0_csc4_10_), .Y(u0__abc_49347_n4946) );
  AND2X2 AND2X2_1474 ( .A(u0__abc_49347_n4535_bF_buf3), .B(u0_tms0_10_), .Y(u0__abc_49347_n4949) );
  AND2X2 AND2X2_1475 ( .A(u0__abc_49347_n4537_bF_buf3), .B(u0_tms2_10_), .Y(u0__abc_49347_n4950) );
  AND2X2 AND2X2_1476 ( .A(u0__abc_49347_n4539_bF_buf3), .B(u0_csc3_10_), .Y(u0__abc_49347_n4951) );
  AND2X2 AND2X2_1477 ( .A(u0__abc_49347_n4582_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n4956) );
  AND2X2 AND2X2_1478 ( .A(u0__abc_49347_n4586_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n4957) );
  AND2X2 AND2X2_1479 ( .A(u0__abc_49347_n4584_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n4958) );
  AND2X2 AND2X2_148 ( .A(spec_req_cs_5_bF_buf5), .B(u0_tms5_3_), .Y(u0__abc_49347_n1257) );
  AND2X2 AND2X2_1480 ( .A(u0__abc_49347_n4571_bF_buf3), .B(u0_tms5_10_), .Y(u0__abc_49347_n4959) );
  AND2X2 AND2X2_1481 ( .A(u0__abc_49347_n4589_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n4960) );
  AND2X2 AND2X2_1482 ( .A(u0__abc_49347_n4565), .B(u0_csc_mask_10_), .Y(u0__abc_49347_n4964) );
  AND2X2 AND2X2_1483 ( .A(u0__abc_49347_n4560_bF_buf3), .B(u0_csc0_10_), .Y(u0__abc_49347_n4965) );
  AND2X2 AND2X2_1484 ( .A(u0__abc_49347_n4562_bF_buf3), .B(u0_csc5_10_), .Y(u0__abc_49347_n4967) );
  AND2X2 AND2X2_1485 ( .A(u0__abc_49347_n4567_bF_buf3), .B(u0_tms4_10_), .Y(u0__abc_49347_n4968) );
  AND2X2 AND2X2_1486 ( .A(u0__abc_49347_n4582_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n4974) );
  AND2X2 AND2X2_1487 ( .A(u0__abc_49347_n4539_bF_buf2), .B(u0_csc3_11_), .Y(u0__abc_49347_n4975) );
  AND2X2 AND2X2_1488 ( .A(u0__abc_49347_n4562_bF_buf2), .B(u0_csc5_11_), .Y(u0__abc_49347_n4976) );
  AND2X2 AND2X2_1489 ( .A(u0__abc_49347_n4511_bF_buf2), .B(_auto_iopadmap_cc_313_execute_56321_11_), .Y(u0__abc_49347_n4978) );
  AND2X2 AND2X2_149 ( .A(u0__abc_49347_n1259), .B(u0__abc_49347_n1185_bF_buf2), .Y(u0__abc_49347_n1260) );
  AND2X2 AND2X2_1490 ( .A(u0__abc_49347_n4528_bF_buf2), .B(u0_tms3_11_), .Y(u0__abc_49347_n4979) );
  AND2X2 AND2X2_1491 ( .A(u0__abc_49347_n4560_bF_buf2), .B(u0_csc0_11_), .Y(u0__abc_49347_n4982) );
  AND2X2 AND2X2_1492 ( .A(u0__abc_49347_n4526_bF_buf2), .B(u0_csc1_11_), .Y(u0__abc_49347_n4983) );
  AND2X2 AND2X2_1493 ( .A(u0__abc_49347_n4535_bF_buf2), .B(u0_tms0_11_), .Y(u0__abc_49347_n4985) );
  AND2X2 AND2X2_1494 ( .A(u0__abc_49347_n4531_bF_buf2), .B(u0_csc4_11_), .Y(u0__abc_49347_n4986) );
  AND2X2 AND2X2_1495 ( .A(u0__abc_49347_n4537_bF_buf2), .B(u0_tms2_11_), .Y(u0__abc_49347_n4990) );
  AND2X2 AND2X2_1496 ( .A(u0__abc_49347_n4567_bF_buf2), .B(u0_tms4_11_), .Y(u0__abc_49347_n4991) );
  AND2X2 AND2X2_1497 ( .A(u0__abc_49347_n4571_bF_buf2), .B(u0_tms5_11_), .Y(u0__abc_49347_n4993) );
  AND2X2 AND2X2_1498 ( .A(u0__abc_49347_n4584_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n4994) );
  AND2X2 AND2X2_1499 ( .A(u0__abc_49347_n4516_bF_buf2), .B(u0_tms1_11_), .Y(u0__abc_49347_n4997) );
  AND2X2 AND2X2_15 ( .A(_abc_55805_n281), .B(_abc_55805_n282), .Y(obct_cs_6_) );
  AND2X2 AND2X2_150 ( .A(u0__abc_49347_n1260), .B(u0__abc_49347_n1258), .Y(u0__abc_49347_n1261) );
  AND2X2 AND2X2_1500 ( .A(u0__abc_49347_n4519_bF_buf2), .B(u0_csc2_11_), .Y(u0__abc_49347_n4998) );
  AND2X2 AND2X2_1501 ( .A(u0__abc_49347_n4589_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n5000) );
  AND2X2 AND2X2_1502 ( .A(u0__abc_49347_n4586_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n5001) );
  AND2X2 AND2X2_1503 ( .A(u0__abc_49347_n4582_bF_buf2), .B(1'b0), .Y(u0__abc_49347_n5007) );
  AND2X2 AND2X2_1504 ( .A(u0__abc_49347_n4511_bF_buf1), .B(_auto_iopadmap_cc_313_execute_56321_12_), .Y(u0__abc_49347_n5008) );
  AND2X2 AND2X2_1505 ( .A(u0__abc_49347_n4560_bF_buf1), .B(u0_csc0_12_), .Y(u0__abc_49347_n5009) );
  AND2X2 AND2X2_1506 ( .A(u0__abc_49347_n4526_bF_buf1), .B(u0_csc1_12_), .Y(u0__abc_49347_n5011) );
  AND2X2 AND2X2_1507 ( .A(u0__abc_49347_n4535_bF_buf1), .B(u0_tms0_12_), .Y(u0__abc_49347_n5012) );
  AND2X2 AND2X2_1508 ( .A(u0__abc_49347_n4519_bF_buf1), .B(u0_csc2_12_), .Y(u0__abc_49347_n5015) );
  AND2X2 AND2X2_1509 ( .A(u0__abc_49347_n4516_bF_buf1), .B(u0_tms1_12_), .Y(u0__abc_49347_n5016) );
  AND2X2 AND2X2_151 ( .A(u0__abc_49347_n1262), .B(u0__abc_49347_n1181_bF_buf2), .Y(u0__abc_49347_n1263_1) );
  AND2X2 AND2X2_1510 ( .A(u0__abc_49347_n4537_bF_buf1), .B(u0_tms2_12_), .Y(u0__abc_49347_n5018) );
  AND2X2 AND2X2_1511 ( .A(u0__abc_49347_n4539_bF_buf1), .B(u0_csc3_12_), .Y(u0__abc_49347_n5019) );
  AND2X2 AND2X2_1512 ( .A(u0__abc_49347_n4589_bF_buf2), .B(1'b0), .Y(u0__abc_49347_n5023) );
  AND2X2 AND2X2_1513 ( .A(u0__abc_49347_n4571_bF_buf1), .B(u0_tms5_12_), .Y(u0__abc_49347_n5024) );
  AND2X2 AND2X2_1514 ( .A(u0__abc_49347_n4584_bF_buf2), .B(1'b0), .Y(u0__abc_49347_n5026) );
  AND2X2 AND2X2_1515 ( .A(u0__abc_49347_n4586_bF_buf2), .B(1'b0), .Y(u0__abc_49347_n5027) );
  AND2X2 AND2X2_1516 ( .A(u0__abc_49347_n4531_bF_buf1), .B(u0_csc4_12_), .Y(u0__abc_49347_n5030) );
  AND2X2 AND2X2_1517 ( .A(u0__abc_49347_n4528_bF_buf1), .B(u0_tms3_12_), .Y(u0__abc_49347_n5031) );
  AND2X2 AND2X2_1518 ( .A(u0__abc_49347_n4567_bF_buf1), .B(u0_tms4_12_), .Y(u0__abc_49347_n5033) );
  AND2X2 AND2X2_1519 ( .A(u0__abc_49347_n4562_bF_buf1), .B(u0_csc5_12_), .Y(u0__abc_49347_n5034) );
  AND2X2 AND2X2_152 ( .A(spec_req_cs_4_bF_buf5), .B(u0_tms4_3_), .Y(u0__abc_49347_n1264_1) );
  AND2X2 AND2X2_1520 ( .A(u0__abc_49347_n4582_bF_buf1), .B(1'b0), .Y(u0__abc_49347_n5040) );
  AND2X2 AND2X2_1521 ( .A(u0__abc_49347_n4589_bF_buf1), .B(1'b0), .Y(u0__abc_49347_n5041) );
  AND2X2 AND2X2_1522 ( .A(u0__abc_49347_n4586_bF_buf1), .B(1'b0), .Y(u0__abc_49347_n5042) );
  AND2X2 AND2X2_1523 ( .A(u0__abc_49347_n4562_bF_buf0), .B(u0_csc5_13_), .Y(u0__abc_49347_n5044) );
  AND2X2 AND2X2_1524 ( .A(u0__abc_49347_n4584_bF_buf1), .B(1'b0), .Y(u0__abc_49347_n5045) );
  AND2X2 AND2X2_1525 ( .A(u0__abc_49347_n4531_bF_buf0), .B(u0_csc4_13_), .Y(u0__abc_49347_n5048) );
  AND2X2 AND2X2_1526 ( .A(u0__abc_49347_n4567_bF_buf0), .B(u0_tms4_13_), .Y(u0__abc_49347_n5049) );
  AND2X2 AND2X2_1527 ( .A(u0__abc_49347_n4528_bF_buf0), .B(u0_tms3_13_), .Y(u0__abc_49347_n5051) );
  AND2X2 AND2X2_1528 ( .A(u0__abc_49347_n4571_bF_buf0), .B(u0_tms5_13_), .Y(u0__abc_49347_n5052) );
  AND2X2 AND2X2_1529 ( .A(u0__abc_49347_n4560_bF_buf0), .B(u0_csc0_13_), .Y(u0__abc_49347_n5056) );
  AND2X2 AND2X2_153 ( .A(u0__abc_49347_n1265), .B(u0__abc_49347_n1180_1_bF_buf2), .Y(u0__abc_49347_n1266) );
  AND2X2 AND2X2_1530 ( .A(u0__abc_49347_n4511_bF_buf0), .B(_auto_iopadmap_cc_313_execute_56321_13_), .Y(u0__abc_49347_n5057) );
  AND2X2 AND2X2_1531 ( .A(u0__abc_49347_n4516_bF_buf0), .B(u0_tms1_13_), .Y(u0__abc_49347_n5059) );
  AND2X2 AND2X2_1532 ( .A(u0__abc_49347_n4537_bF_buf0), .B(u0_tms2_13_), .Y(u0__abc_49347_n5060) );
  AND2X2 AND2X2_1533 ( .A(u0__abc_49347_n4535_bF_buf0), .B(u0_tms0_13_), .Y(u0__abc_49347_n5063) );
  AND2X2 AND2X2_1534 ( .A(u0__abc_49347_n4526_bF_buf0), .B(u0_csc1_13_), .Y(u0__abc_49347_n5064) );
  AND2X2 AND2X2_1535 ( .A(u0__abc_49347_n4519_bF_buf0), .B(u0_csc2_13_), .Y(u0__abc_49347_n5066) );
  AND2X2 AND2X2_1536 ( .A(u0__abc_49347_n4539_bF_buf0), .B(u0_csc3_13_), .Y(u0__abc_49347_n5067) );
  AND2X2 AND2X2_1537 ( .A(u0__abc_49347_n4582_bF_buf0), .B(1'b0), .Y(u0__abc_49347_n5073) );
  AND2X2 AND2X2_1538 ( .A(u0__abc_49347_n4516_bF_buf4), .B(u0_tms1_14_), .Y(u0__abc_49347_n5074) );
  AND2X2 AND2X2_1539 ( .A(u0__abc_49347_n4539_bF_buf4), .B(u0_csc3_14_), .Y(u0__abc_49347_n5075) );
  AND2X2 AND2X2_154 ( .A(spec_req_cs_3_bF_buf5), .B(u0_tms3_3_), .Y(u0__abc_49347_n1267) );
  AND2X2 AND2X2_1540 ( .A(u0__abc_49347_n4511_bF_buf4), .B(_auto_iopadmap_cc_313_execute_56321_14_), .Y(u0__abc_49347_n5077) );
  AND2X2 AND2X2_1541 ( .A(u0__abc_49347_n4571_bF_buf4), .B(u0_tms5_14_), .Y(u0__abc_49347_n5078) );
  AND2X2 AND2X2_1542 ( .A(u0__abc_49347_n4519_bF_buf4), .B(u0_csc2_14_), .Y(u0__abc_49347_n5081) );
  AND2X2 AND2X2_1543 ( .A(u0__abc_49347_n4531_bF_buf4), .B(u0_csc4_14_), .Y(u0__abc_49347_n5082) );
  AND2X2 AND2X2_1544 ( .A(u0__abc_49347_n4535_bF_buf4), .B(u0_tms0_14_), .Y(u0__abc_49347_n5084) );
  AND2X2 AND2X2_1545 ( .A(u0__abc_49347_n4567_bF_buf4), .B(u0_tms4_14_), .Y(u0__abc_49347_n5085) );
  AND2X2 AND2X2_1546 ( .A(u0__abc_49347_n4537_bF_buf4), .B(u0_tms2_14_), .Y(u0__abc_49347_n5089) );
  AND2X2 AND2X2_1547 ( .A(u0__abc_49347_n4562_bF_buf4), .B(u0_csc5_14_), .Y(u0__abc_49347_n5090) );
  AND2X2 AND2X2_1548 ( .A(u0__abc_49347_n4560_bF_buf4), .B(u0_csc0_14_), .Y(u0__abc_49347_n5092) );
  AND2X2 AND2X2_1549 ( .A(u0__abc_49347_n4528_bF_buf4), .B(u0_tms3_14_), .Y(u0__abc_49347_n5093) );
  AND2X2 AND2X2_155 ( .A(u0__abc_49347_n1268), .B(u0__abc_49347_n1179_bF_buf2), .Y(u0__abc_49347_n1269) );
  AND2X2 AND2X2_1550 ( .A(u0__abc_49347_n4589_bF_buf0), .B(1'b0), .Y(u0__abc_49347_n5096) );
  AND2X2 AND2X2_1551 ( .A(u0__abc_49347_n4584_bF_buf0), .B(1'b0), .Y(u0__abc_49347_n5097) );
  AND2X2 AND2X2_1552 ( .A(u0__abc_49347_n4526_bF_buf4), .B(u0_csc1_14_), .Y(u0__abc_49347_n5099) );
  AND2X2 AND2X2_1553 ( .A(u0__abc_49347_n4586_bF_buf0), .B(1'b0), .Y(u0__abc_49347_n5100) );
  AND2X2 AND2X2_1554 ( .A(u0__abc_49347_n4582_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n5106) );
  AND2X2 AND2X2_1555 ( .A(u0__abc_49347_n4586_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n5107) );
  AND2X2 AND2X2_1556 ( .A(u0__abc_49347_n4584_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n5108) );
  AND2X2 AND2X2_1557 ( .A(u0__abc_49347_n4562_bF_buf3), .B(u0_csc5_15_), .Y(u0__abc_49347_n5110) );
  AND2X2 AND2X2_1558 ( .A(u0__abc_49347_n4589_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n5111) );
  AND2X2 AND2X2_1559 ( .A(u0__abc_49347_n4531_bF_buf3), .B(u0_csc4_15_), .Y(u0__abc_49347_n5114) );
  AND2X2 AND2X2_156 ( .A(spec_req_cs_2_bF_buf5), .B(u0_tms2_3_), .Y(u0__abc_49347_n1270) );
  AND2X2 AND2X2_1560 ( .A(u0__abc_49347_n4567_bF_buf3), .B(u0_tms4_15_), .Y(u0__abc_49347_n5115) );
  AND2X2 AND2X2_1561 ( .A(u0__abc_49347_n4528_bF_buf3), .B(u0_tms3_15_), .Y(u0__abc_49347_n5117) );
  AND2X2 AND2X2_1562 ( .A(u0__abc_49347_n4571_bF_buf3), .B(u0_tms5_15_), .Y(u0__abc_49347_n5118) );
  AND2X2 AND2X2_1563 ( .A(u0__abc_49347_n4560_bF_buf3), .B(u0_csc0_15_), .Y(u0__abc_49347_n5122) );
  AND2X2 AND2X2_1564 ( .A(u0__abc_49347_n4511_bF_buf3), .B(_auto_iopadmap_cc_313_execute_56321_15_), .Y(u0__abc_49347_n5123) );
  AND2X2 AND2X2_1565 ( .A(u0__abc_49347_n4516_bF_buf3), .B(u0_tms1_15_), .Y(u0__abc_49347_n5125) );
  AND2X2 AND2X2_1566 ( .A(u0__abc_49347_n4537_bF_buf3), .B(u0_tms2_15_), .Y(u0__abc_49347_n5126) );
  AND2X2 AND2X2_1567 ( .A(u0__abc_49347_n4535_bF_buf3), .B(u0_tms0_15_), .Y(u0__abc_49347_n5129) );
  AND2X2 AND2X2_1568 ( .A(u0__abc_49347_n4526_bF_buf3), .B(u0_csc1_15_), .Y(u0__abc_49347_n5130) );
  AND2X2 AND2X2_1569 ( .A(u0__abc_49347_n4519_bF_buf3), .B(u0_csc2_15_), .Y(u0__abc_49347_n5132) );
  AND2X2 AND2X2_157 ( .A(u0__abc_49347_n1271), .B(u0__abc_49347_n1178_1_bF_buf2), .Y(u0__abc_49347_n1272_1) );
  AND2X2 AND2X2_1570 ( .A(u0__abc_49347_n4539_bF_buf3), .B(u0_csc3_15_), .Y(u0__abc_49347_n5133) );
  AND2X2 AND2X2_1571 ( .A(u0__abc_49347_n4582_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n5139) );
  AND2X2 AND2X2_1572 ( .A(u0__abc_49347_n4511_bF_buf2), .B(_auto_iopadmap_cc_313_execute_56321_16_), .Y(u0__abc_49347_n5140) );
  AND2X2 AND2X2_1573 ( .A(u0__abc_49347_n4560_bF_buf2), .B(u0_csc0_16_), .Y(u0__abc_49347_n5141) );
  AND2X2 AND2X2_1574 ( .A(u0__abc_49347_n4526_bF_buf2), .B(u0_csc1_16_), .Y(u0__abc_49347_n5143) );
  AND2X2 AND2X2_1575 ( .A(u0__abc_49347_n4535_bF_buf2), .B(u0_tms0_16_), .Y(u0__abc_49347_n5144) );
  AND2X2 AND2X2_1576 ( .A(u0__abc_49347_n4519_bF_buf2), .B(u0_csc2_16_), .Y(u0__abc_49347_n5147) );
  AND2X2 AND2X2_1577 ( .A(u0__abc_49347_n4516_bF_buf2), .B(u0_tms1_16_), .Y(u0__abc_49347_n5148) );
  AND2X2 AND2X2_1578 ( .A(u0__abc_49347_n4537_bF_buf2), .B(u0_tms2_16_), .Y(u0__abc_49347_n5150) );
  AND2X2 AND2X2_1579 ( .A(u0__abc_49347_n4539_bF_buf2), .B(u0_csc3_16_), .Y(u0__abc_49347_n5151) );
  AND2X2 AND2X2_158 ( .A(spec_req_cs_1_bF_buf5), .B(u0_tms1_3_), .Y(u0__abc_49347_n1273_1) );
  AND2X2 AND2X2_1580 ( .A(u0__abc_49347_n4571_bF_buf2), .B(u0_tms5_16_), .Y(u0__abc_49347_n5155) );
  AND2X2 AND2X2_1581 ( .A(u0__abc_49347_n4589_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n5156) );
  AND2X2 AND2X2_1582 ( .A(u0__abc_49347_n4584_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n5158) );
  AND2X2 AND2X2_1583 ( .A(u0__abc_49347_n4528_bF_buf2), .B(u0_tms3_16_), .Y(u0__abc_49347_n5159) );
  AND2X2 AND2X2_1584 ( .A(u0__abc_49347_n4586_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n5162) );
  AND2X2 AND2X2_1585 ( .A(u0__abc_49347_n4562_bF_buf2), .B(u0_csc5_16_), .Y(u0__abc_49347_n5163) );
  AND2X2 AND2X2_1586 ( .A(u0__abc_49347_n4531_bF_buf2), .B(u0_csc4_16_), .Y(u0__abc_49347_n5165) );
  AND2X2 AND2X2_1587 ( .A(u0__abc_49347_n4567_bF_buf2), .B(u0_tms4_16_), .Y(u0__abc_49347_n5166) );
  AND2X2 AND2X2_1588 ( .A(u0__abc_49347_n4582_bF_buf2), .B(1'b0), .Y(u0__abc_49347_n5172) );
  AND2X2 AND2X2_1589 ( .A(u0__abc_49347_n4528_bF_buf1), .B(u0_tms3_17_), .Y(u0__abc_49347_n5173) );
  AND2X2 AND2X2_159 ( .A(u0__abc_49347_n1175_bF_buf2), .B(u0__abc_49347_n1276), .Y(u0__abc_49347_n1277) );
  AND2X2 AND2X2_1590 ( .A(u0__abc_49347_n4531_bF_buf1), .B(u0_csc4_17_), .Y(u0__abc_49347_n5174) );
  AND2X2 AND2X2_1591 ( .A(u0__abc_49347_n4567_bF_buf1), .B(u0_tms4_17_), .Y(u0__abc_49347_n5176) );
  AND2X2 AND2X2_1592 ( .A(u0__abc_49347_n4562_bF_buf1), .B(u0_csc5_17_), .Y(u0__abc_49347_n5177) );
  AND2X2 AND2X2_1593 ( .A(u0__abc_49347_n4589_bF_buf2), .B(1'b0), .Y(u0__abc_49347_n5180) );
  AND2X2 AND2X2_1594 ( .A(u0__abc_49347_n4571_bF_buf1), .B(u0_tms5_17_), .Y(u0__abc_49347_n5181) );
  AND2X2 AND2X2_1595 ( .A(u0__abc_49347_n4584_bF_buf2), .B(1'b0), .Y(u0__abc_49347_n5183) );
  AND2X2 AND2X2_1596 ( .A(u0__abc_49347_n4586_bF_buf2), .B(1'b0), .Y(u0__abc_49347_n5184) );
  AND2X2 AND2X2_1597 ( .A(u0__abc_49347_n4516_bF_buf1), .B(u0_tms1_17_), .Y(u0__abc_49347_n5188) );
  AND2X2 AND2X2_1598 ( .A(u0__abc_49347_n4539_bF_buf1), .B(u0_csc3_17_), .Y(u0__abc_49347_n5189) );
  AND2X2 AND2X2_1599 ( .A(u0__abc_49347_n4519_bF_buf1), .B(u0_csc2_17_), .Y(u0__abc_49347_n5191) );
  AND2X2 AND2X2_16 ( .A(_abc_55805_n284), .B(_abc_55805_n285), .Y(_abc_55805_n286) );
  AND2X2 AND2X2_160 ( .A(u0__abc_49347_n1275), .B(u0__abc_49347_n1277), .Y(u0__abc_49347_n1278) );
  AND2X2 AND2X2_1600 ( .A(u0__abc_49347_n4526_bF_buf1), .B(u0_csc1_17_), .Y(u0__abc_49347_n5192) );
  AND2X2 AND2X2_1601 ( .A(u0__abc_49347_n4511_bF_buf1), .B(_auto_iopadmap_cc_313_execute_56321_17_), .Y(u0__abc_49347_n5195) );
  AND2X2 AND2X2_1602 ( .A(u0__abc_49347_n4535_bF_buf1), .B(u0_tms0_17_), .Y(u0__abc_49347_n5196) );
  AND2X2 AND2X2_1603 ( .A(u0__abc_49347_n4537_bF_buf1), .B(u0_tms2_17_), .Y(u0__abc_49347_n5198) );
  AND2X2 AND2X2_1604 ( .A(u0__abc_49347_n4560_bF_buf1), .B(u0_csc0_17_), .Y(u0__abc_49347_n5199) );
  AND2X2 AND2X2_1605 ( .A(u0__abc_49347_n4582_bF_buf1), .B(1'b0), .Y(u0__abc_49347_n5205) );
  AND2X2 AND2X2_1606 ( .A(u0__abc_49347_n4560_bF_buf0), .B(u0_csc0_18_), .Y(u0__abc_49347_n5206) );
  AND2X2 AND2X2_1607 ( .A(u0__abc_49347_n4511_bF_buf0), .B(_auto_iopadmap_cc_313_execute_56321_18_), .Y(u0__abc_49347_n5207) );
  AND2X2 AND2X2_1608 ( .A(u0__abc_49347_n4516_bF_buf0), .B(u0_tms1_18_), .Y(u0__abc_49347_n5209) );
  AND2X2 AND2X2_1609 ( .A(u0__abc_49347_n4537_bF_buf0), .B(u0_tms2_18_), .Y(u0__abc_49347_n5210) );
  AND2X2 AND2X2_161 ( .A(u0__abc_49347_n1176_1_bF_buf2), .B(sp_tms_4_), .Y(u0__abc_49347_n1280) );
  AND2X2 AND2X2_1610 ( .A(u0__abc_49347_n4535_bF_buf0), .B(u0_tms0_18_), .Y(u0__abc_49347_n5213) );
  AND2X2 AND2X2_1611 ( .A(u0__abc_49347_n4526_bF_buf0), .B(u0_csc1_18_), .Y(u0__abc_49347_n5214) );
  AND2X2 AND2X2_1612 ( .A(u0__abc_49347_n4519_bF_buf0), .B(u0_csc2_18_), .Y(u0__abc_49347_n5216) );
  AND2X2 AND2X2_1613 ( .A(u0__abc_49347_n4539_bF_buf0), .B(u0_csc3_18_), .Y(u0__abc_49347_n5217) );
  AND2X2 AND2X2_1614 ( .A(u0__abc_49347_n4589_bF_buf1), .B(1'b0), .Y(u0__abc_49347_n5221) );
  AND2X2 AND2X2_1615 ( .A(u0__abc_49347_n4571_bF_buf0), .B(u0_tms5_18_), .Y(u0__abc_49347_n5222) );
  AND2X2 AND2X2_1616 ( .A(u0__abc_49347_n4584_bF_buf1), .B(1'b0), .Y(u0__abc_49347_n5224) );
  AND2X2 AND2X2_1617 ( .A(u0__abc_49347_n4586_bF_buf1), .B(1'b0), .Y(u0__abc_49347_n5225) );
  AND2X2 AND2X2_1618 ( .A(u0__abc_49347_n4531_bF_buf0), .B(u0_csc4_18_), .Y(u0__abc_49347_n5228) );
  AND2X2 AND2X2_1619 ( .A(u0__abc_49347_n4528_bF_buf0), .B(u0_tms3_18_), .Y(u0__abc_49347_n5229) );
  AND2X2 AND2X2_162 ( .A(spec_req_cs_5_bF_buf4), .B(u0_tms5_4_), .Y(u0__abc_49347_n1281_1) );
  AND2X2 AND2X2_1620 ( .A(u0__abc_49347_n4562_bF_buf0), .B(u0_csc5_18_), .Y(u0__abc_49347_n5231) );
  AND2X2 AND2X2_1621 ( .A(u0__abc_49347_n4567_bF_buf0), .B(u0_tms4_18_), .Y(u0__abc_49347_n5232) );
  AND2X2 AND2X2_1622 ( .A(u0__abc_49347_n4582_bF_buf0), .B(1'b0), .Y(u0__abc_49347_n5238) );
  AND2X2 AND2X2_1623 ( .A(u0__abc_49347_n4537_bF_buf4), .B(u0_tms2_19_), .Y(u0__abc_49347_n5239) );
  AND2X2 AND2X2_1624 ( .A(u0__abc_49347_n4528_bF_buf4), .B(u0_tms3_19_), .Y(u0__abc_49347_n5240) );
  AND2X2 AND2X2_1625 ( .A(u0__abc_49347_n4511_bF_buf4), .B(_auto_iopadmap_cc_313_execute_56321_19_), .Y(u0__abc_49347_n5242) );
  AND2X2 AND2X2_1626 ( .A(u0__abc_49347_n4562_bF_buf4), .B(u0_csc5_19_), .Y(u0__abc_49347_n5243) );
  AND2X2 AND2X2_1627 ( .A(u0__abc_49347_n4560_bF_buf4), .B(u0_csc0_19_), .Y(u0__abc_49347_n5246) );
  AND2X2 AND2X2_1628 ( .A(u0__abc_49347_n4526_bF_buf4), .B(u0_csc1_19_), .Y(u0__abc_49347_n5247) );
  AND2X2 AND2X2_1629 ( .A(u0__abc_49347_n4535_bF_buf4), .B(u0_tms0_19_), .Y(u0__abc_49347_n5249) );
  AND2X2 AND2X2_163 ( .A(u0__abc_49347_n1283), .B(u0__abc_49347_n1185_bF_buf1), .Y(u0__abc_49347_n1284) );
  AND2X2 AND2X2_1630 ( .A(u0__abc_49347_n4531_bF_buf4), .B(u0_csc4_19_), .Y(u0__abc_49347_n5250) );
  AND2X2 AND2X2_1631 ( .A(u0__abc_49347_n4589_bF_buf0), .B(1'b0), .Y(u0__abc_49347_n5254) );
  AND2X2 AND2X2_1632 ( .A(u0__abc_49347_n4571_bF_buf4), .B(u0_tms5_19_), .Y(u0__abc_49347_n5255) );
  AND2X2 AND2X2_1633 ( .A(u0__abc_49347_n4516_bF_buf4), .B(u0_tms1_19_), .Y(u0__abc_49347_n5257) );
  AND2X2 AND2X2_1634 ( .A(u0__abc_49347_n4567_bF_buf4), .B(u0_tms4_19_), .Y(u0__abc_49347_n5258) );
  AND2X2 AND2X2_1635 ( .A(u0__abc_49347_n4519_bF_buf4), .B(u0_csc2_19_), .Y(u0__abc_49347_n5261) );
  AND2X2 AND2X2_1636 ( .A(u0__abc_49347_n4586_bF_buf0), .B(1'b0), .Y(u0__abc_49347_n5262) );
  AND2X2 AND2X2_1637 ( .A(u0__abc_49347_n4539_bF_buf4), .B(u0_csc3_19_), .Y(u0__abc_49347_n5264) );
  AND2X2 AND2X2_1638 ( .A(u0__abc_49347_n4584_bF_buf0), .B(1'b0), .Y(u0__abc_49347_n5265) );
  AND2X2 AND2X2_1639 ( .A(u0__abc_49347_n4582_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n5271) );
  AND2X2 AND2X2_164 ( .A(u0__abc_49347_n1284), .B(u0__abc_49347_n1282_1), .Y(u0__abc_49347_n1285) );
  AND2X2 AND2X2_1640 ( .A(u0__abc_49347_n4511_bF_buf3), .B(_auto_iopadmap_cc_313_execute_56321_20_), .Y(u0__abc_49347_n5272) );
  AND2X2 AND2X2_1641 ( .A(u0__abc_49347_n4560_bF_buf3), .B(u0_csc0_20_), .Y(u0__abc_49347_n5273) );
  AND2X2 AND2X2_1642 ( .A(u0__abc_49347_n4526_bF_buf3), .B(u0_csc1_20_), .Y(u0__abc_49347_n5275) );
  AND2X2 AND2X2_1643 ( .A(u0__abc_49347_n4535_bF_buf3), .B(u0_tms0_20_), .Y(u0__abc_49347_n5276) );
  AND2X2 AND2X2_1644 ( .A(u0__abc_49347_n4537_bF_buf3), .B(u0_tms2_20_), .Y(u0__abc_49347_n5279) );
  AND2X2 AND2X2_1645 ( .A(u0__abc_49347_n4539_bF_buf3), .B(u0_csc3_20_), .Y(u0__abc_49347_n5280) );
  AND2X2 AND2X2_1646 ( .A(u0__abc_49347_n4519_bF_buf3), .B(u0_csc2_20_), .Y(u0__abc_49347_n5282) );
  AND2X2 AND2X2_1647 ( .A(u0__abc_49347_n4516_bF_buf3), .B(u0_tms1_20_), .Y(u0__abc_49347_n5283) );
  AND2X2 AND2X2_1648 ( .A(u0__abc_49347_n4589_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n5287) );
  AND2X2 AND2X2_1649 ( .A(u0__abc_49347_n4571_bF_buf3), .B(u0_tms5_20_), .Y(u0__abc_49347_n5288) );
  AND2X2 AND2X2_165 ( .A(u0__abc_49347_n1286), .B(u0__abc_49347_n1181_bF_buf1), .Y(u0__abc_49347_n1287) );
  AND2X2 AND2X2_1650 ( .A(u0__abc_49347_n4586_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n5290) );
  AND2X2 AND2X2_1651 ( .A(u0__abc_49347_n4584_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n5291) );
  AND2X2 AND2X2_1652 ( .A(u0__abc_49347_n4528_bF_buf3), .B(u0_tms3_20_), .Y(u0__abc_49347_n5294) );
  AND2X2 AND2X2_1653 ( .A(u0__abc_49347_n4531_bF_buf3), .B(u0_csc4_20_), .Y(u0__abc_49347_n5295) );
  AND2X2 AND2X2_1654 ( .A(u0__abc_49347_n4567_bF_buf3), .B(u0_tms4_20_), .Y(u0__abc_49347_n5297) );
  AND2X2 AND2X2_1655 ( .A(u0__abc_49347_n4562_bF_buf3), .B(u0_csc5_20_), .Y(u0__abc_49347_n5298) );
  AND2X2 AND2X2_1656 ( .A(u0__abc_49347_n4582_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n5304) );
  AND2X2 AND2X2_1657 ( .A(u0__abc_49347_n4560_bF_buf2), .B(u0_csc0_21_), .Y(u0__abc_49347_n5305) );
  AND2X2 AND2X2_1658 ( .A(u0__abc_49347_n4511_bF_buf2), .B(_auto_iopadmap_cc_313_execute_56321_21_), .Y(u0__abc_49347_n5306) );
  AND2X2 AND2X2_1659 ( .A(u0__abc_49347_n4535_bF_buf2), .B(u0_tms0_21_), .Y(u0__abc_49347_n5308) );
  AND2X2 AND2X2_166 ( .A(spec_req_cs_4_bF_buf4), .B(u0_tms4_4_), .Y(u0__abc_49347_n1288) );
  AND2X2 AND2X2_1660 ( .A(u0__abc_49347_n4526_bF_buf2), .B(u0_csc1_21_), .Y(u0__abc_49347_n5309) );
  AND2X2 AND2X2_1661 ( .A(u0__abc_49347_n4516_bF_buf2), .B(u0_tms1_21_), .Y(u0__abc_49347_n5312) );
  AND2X2 AND2X2_1662 ( .A(u0__abc_49347_n4519_bF_buf2), .B(u0_csc2_21_), .Y(u0__abc_49347_n5313) );
  AND2X2 AND2X2_1663 ( .A(u0__abc_49347_n4537_bF_buf2), .B(u0_tms2_21_), .Y(u0__abc_49347_n5315) );
  AND2X2 AND2X2_1664 ( .A(u0__abc_49347_n4539_bF_buf2), .B(u0_csc3_21_), .Y(u0__abc_49347_n5316) );
  AND2X2 AND2X2_1665 ( .A(u0__abc_49347_n4589_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n5320) );
  AND2X2 AND2X2_1666 ( .A(u0__abc_49347_n4571_bF_buf2), .B(u0_tms5_21_), .Y(u0__abc_49347_n5321) );
  AND2X2 AND2X2_1667 ( .A(u0__abc_49347_n4586_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n5323) );
  AND2X2 AND2X2_1668 ( .A(u0__abc_49347_n4584_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n5324) );
  AND2X2 AND2X2_1669 ( .A(u0__abc_49347_n4528_bF_buf2), .B(u0_tms3_21_), .Y(u0__abc_49347_n5327) );
  AND2X2 AND2X2_167 ( .A(u0__abc_49347_n1289), .B(u0__abc_49347_n1180_1_bF_buf1), .Y(u0__abc_49347_n1290_1) );
  AND2X2 AND2X2_1670 ( .A(u0__abc_49347_n4531_bF_buf2), .B(u0_csc4_21_), .Y(u0__abc_49347_n5328) );
  AND2X2 AND2X2_1671 ( .A(u0__abc_49347_n4562_bF_buf2), .B(u0_csc5_21_), .Y(u0__abc_49347_n5330) );
  AND2X2 AND2X2_1672 ( .A(u0__abc_49347_n4567_bF_buf2), .B(u0_tms4_21_), .Y(u0__abc_49347_n5331) );
  AND2X2 AND2X2_1673 ( .A(u0__abc_49347_n4582_bF_buf2), .B(1'b0), .Y(u0__abc_49347_n5337) );
  AND2X2 AND2X2_1674 ( .A(u0__abc_49347_n4560_bF_buf1), .B(u0_csc0_22_), .Y(u0__abc_49347_n5338) );
  AND2X2 AND2X2_1675 ( .A(u0__abc_49347_n4535_bF_buf1), .B(u0_tms0_22_), .Y(u0__abc_49347_n5339) );
  AND2X2 AND2X2_1676 ( .A(u0__abc_49347_n4516_bF_buf1), .B(u0_tms1_22_), .Y(u0__abc_49347_n5341) );
  AND2X2 AND2X2_1677 ( .A(u0__abc_49347_n4539_bF_buf1), .B(u0_csc3_22_), .Y(u0__abc_49347_n5342) );
  AND2X2 AND2X2_1678 ( .A(u0__abc_49347_n4526_bF_buf1), .B(u0_csc1_22_), .Y(u0__abc_49347_n5345) );
  AND2X2 AND2X2_1679 ( .A(u0__abc_49347_n4519_bF_buf1), .B(u0_csc2_22_), .Y(u0__abc_49347_n5346) );
  AND2X2 AND2X2_168 ( .A(spec_req_cs_3_bF_buf4), .B(u0_tms3_4_), .Y(u0__abc_49347_n1291_1) );
  AND2X2 AND2X2_1680 ( .A(u0__abc_49347_n4511_bF_buf1), .B(_auto_iopadmap_cc_313_execute_56321_22_), .Y(u0__abc_49347_n5348) );
  AND2X2 AND2X2_1681 ( .A(u0__abc_49347_n4537_bF_buf1), .B(u0_tms2_22_), .Y(u0__abc_49347_n5349) );
  AND2X2 AND2X2_1682 ( .A(u0__abc_49347_n4589_bF_buf2), .B(1'b0), .Y(u0__abc_49347_n5353) );
  AND2X2 AND2X2_1683 ( .A(u0__abc_49347_n4571_bF_buf1), .B(u0_tms5_22_), .Y(u0__abc_49347_n5354) );
  AND2X2 AND2X2_1684 ( .A(u0__abc_49347_n4586_bF_buf2), .B(1'b0), .Y(u0__abc_49347_n5356) );
  AND2X2 AND2X2_1685 ( .A(u0__abc_49347_n4584_bF_buf2), .B(1'b0), .Y(u0__abc_49347_n5357) );
  AND2X2 AND2X2_1686 ( .A(u0__abc_49347_n4531_bF_buf1), .B(u0_csc4_22_), .Y(u0__abc_49347_n5360) );
  AND2X2 AND2X2_1687 ( .A(u0__abc_49347_n4528_bF_buf1), .B(u0_tms3_22_), .Y(u0__abc_49347_n5361) );
  AND2X2 AND2X2_1688 ( .A(u0__abc_49347_n4562_bF_buf1), .B(u0_csc5_22_), .Y(u0__abc_49347_n5363) );
  AND2X2 AND2X2_1689 ( .A(u0__abc_49347_n4567_bF_buf1), .B(u0_tms4_22_), .Y(u0__abc_49347_n5364) );
  AND2X2 AND2X2_169 ( .A(u0__abc_49347_n1292), .B(u0__abc_49347_n1179_bF_buf1), .Y(u0__abc_49347_n1293) );
  AND2X2 AND2X2_1690 ( .A(u0__abc_49347_n4582_bF_buf1), .B(1'b0), .Y(u0__abc_49347_n5370) );
  AND2X2 AND2X2_1691 ( .A(u0__abc_49347_n4516_bF_buf0), .B(u0_tms1_23_), .Y(u0__abc_49347_n5371) );
  AND2X2 AND2X2_1692 ( .A(u0__abc_49347_n4539_bF_buf0), .B(u0_csc3_23_), .Y(u0__abc_49347_n5372) );
  AND2X2 AND2X2_1693 ( .A(u0__abc_49347_n4571_bF_buf0), .B(u0_tms5_23_), .Y(u0__abc_49347_n5374) );
  AND2X2 AND2X2_1694 ( .A(u0__abc_49347_n4586_bF_buf1), .B(1'b0), .Y(u0__abc_49347_n5375) );
  AND2X2 AND2X2_1695 ( .A(u0__abc_49347_n4537_bF_buf0), .B(u0_tms2_23_), .Y(u0__abc_49347_n5378) );
  AND2X2 AND2X2_1696 ( .A(u0__abc_49347_n4560_bF_buf0), .B(u0_csc0_23_), .Y(u0__abc_49347_n5379) );
  AND2X2 AND2X2_1697 ( .A(u0__abc_49347_n4526_bF_buf0), .B(u0_csc1_23_), .Y(u0__abc_49347_n5381) );
  AND2X2 AND2X2_1698 ( .A(u0__abc_49347_n4562_bF_buf0), .B(u0_csc5_23_), .Y(u0__abc_49347_n5382) );
  AND2X2 AND2X2_1699 ( .A(u0__abc_49347_n4511_bF_buf0), .B(_auto_iopadmap_cc_313_execute_56321_23_), .Y(u0__abc_49347_n5386) );
  AND2X2 AND2X2_17 ( .A(_abc_55805_n287), .B(_abc_55805_n288), .Y(obct_cs_7_) );
  AND2X2 AND2X2_170 ( .A(spec_req_cs_2_bF_buf4), .B(u0_tms2_4_), .Y(u0__abc_49347_n1294) );
  AND2X2 AND2X2_1700 ( .A(u0__abc_49347_n4567_bF_buf0), .B(u0_tms4_23_), .Y(u0__abc_49347_n5387) );
  AND2X2 AND2X2_1701 ( .A(u0__abc_49347_n4535_bF_buf0), .B(u0_tms0_23_), .Y(u0__abc_49347_n5389) );
  AND2X2 AND2X2_1702 ( .A(u0__abc_49347_n4584_bF_buf1), .B(1'b0), .Y(u0__abc_49347_n5390) );
  AND2X2 AND2X2_1703 ( .A(u0__abc_49347_n4528_bF_buf0), .B(u0_tms3_23_), .Y(u0__abc_49347_n5393) );
  AND2X2 AND2X2_1704 ( .A(u0__abc_49347_n4531_bF_buf0), .B(u0_csc4_23_), .Y(u0__abc_49347_n5394) );
  AND2X2 AND2X2_1705 ( .A(u0__abc_49347_n4519_bF_buf0), .B(u0_csc2_23_), .Y(u0__abc_49347_n5396) );
  AND2X2 AND2X2_1706 ( .A(u0__abc_49347_n4589_bF_buf1), .B(1'b0), .Y(u0__abc_49347_n5397) );
  AND2X2 AND2X2_1707 ( .A(u0__abc_49347_n4560_bF_buf4), .B(u0_csc0_24_), .Y(u0__abc_49347_n5403) );
  AND2X2 AND2X2_1708 ( .A(u0__abc_49347_n4511_bF_buf4), .B(_auto_iopadmap_cc_313_execute_56321_24_), .Y(u0__abc_49347_n5404) );
  AND2X2 AND2X2_1709 ( .A(u0__abc_49347_n4516_bF_buf4), .B(u0_tms1_24_), .Y(u0__abc_49347_n5405) );
  AND2X2 AND2X2_171 ( .A(u0__abc_49347_n1295), .B(u0__abc_49347_n1178_1_bF_buf1), .Y(u0__abc_49347_n1296) );
  AND2X2 AND2X2_1710 ( .A(u0__abc_49347_n4519_bF_buf4), .B(u0_csc2_24_), .Y(u0__abc_49347_n5406) );
  AND2X2 AND2X2_1711 ( .A(u0__abc_49347_n4526_bF_buf4), .B(u0_csc1_24_), .Y(u0__abc_49347_n5410) );
  AND2X2 AND2X2_1712 ( .A(u0__abc_49347_n4528_bF_buf4), .B(u0_tms3_24_), .Y(u0__abc_49347_n5411) );
  AND2X2 AND2X2_1713 ( .A(u0__abc_49347_n4531_bF_buf4), .B(u0_csc4_24_), .Y(u0__abc_49347_n5412) );
  AND2X2 AND2X2_1714 ( .A(u0__abc_49347_n4535_bF_buf4), .B(u0_tms0_24_), .Y(u0__abc_49347_n5415) );
  AND2X2 AND2X2_1715 ( .A(u0__abc_49347_n4537_bF_buf4), .B(u0_tms2_24_), .Y(u0__abc_49347_n5416) );
  AND2X2 AND2X2_1716 ( .A(u0__abc_49347_n4539_bF_buf4), .B(u0_csc3_24_), .Y(u0__abc_49347_n5417) );
  AND2X2 AND2X2_1717 ( .A(u0__abc_49347_n4582_bF_buf0), .B(1'b0), .Y(u0__abc_49347_n5422) );
  AND2X2 AND2X2_1718 ( .A(u0__abc_49347_n4589_bF_buf0), .B(1'b0), .Y(u0__abc_49347_n5423) );
  AND2X2 AND2X2_1719 ( .A(u0__abc_49347_n4584_bF_buf0), .B(1'b0), .Y(u0__abc_49347_n5424) );
  AND2X2 AND2X2_172 ( .A(spec_req_cs_1_bF_buf4), .B(u0_tms1_4_), .Y(u0__abc_49347_n1297) );
  AND2X2 AND2X2_1720 ( .A(u0__abc_49347_n4586_bF_buf0), .B(1'b0), .Y(u0__abc_49347_n5426) );
  AND2X2 AND2X2_1721 ( .A(u0__abc_49347_n4507_bF_buf3), .B(rfr_ps_val_0_), .Y(u0__abc_49347_n5428) );
  AND2X2 AND2X2_1722 ( .A(u0__abc_49347_n4567_bF_buf4), .B(u0_tms4_24_), .Y(u0__abc_49347_n5429) );
  AND2X2 AND2X2_1723 ( .A(u0__abc_49347_n4562_bF_buf4), .B(u0_csc5_24_), .Y(u0__abc_49347_n5431) );
  AND2X2 AND2X2_1724 ( .A(u0__abc_49347_n4571_bF_buf4), .B(u0_tms5_24_), .Y(u0__abc_49347_n5432) );
  AND2X2 AND2X2_1725 ( .A(u0__abc_49347_n4582_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n5438) );
  AND2X2 AND2X2_1726 ( .A(u0__abc_49347_n4535_bF_buf3), .B(u0_tms0_25_), .Y(u0__abc_49347_n5439) );
  AND2X2 AND2X2_1727 ( .A(u0__abc_49347_n4531_bF_buf3), .B(u0_csc4_25_), .Y(u0__abc_49347_n5440) );
  AND2X2 AND2X2_1728 ( .A(u0__abc_49347_n4528_bF_buf3), .B(u0_tms3_25_), .Y(u0__abc_49347_n5441) );
  AND2X2 AND2X2_1729 ( .A(u0__abc_49347_n4526_bF_buf3), .B(u0_csc1_25_), .Y(u0__abc_49347_n5444) );
  AND2X2 AND2X2_173 ( .A(u0__abc_49347_n1175_bF_buf1), .B(u0__abc_49347_n1300_1), .Y(u0__abc_49347_n1301) );
  AND2X2 AND2X2_1730 ( .A(u0__abc_49347_n4537_bF_buf3), .B(u0_tms2_25_), .Y(u0__abc_49347_n5445) );
  AND2X2 AND2X2_1731 ( .A(u0__abc_49347_n4539_bF_buf3), .B(u0_csc3_25_), .Y(u0__abc_49347_n5446) );
  AND2X2 AND2X2_1732 ( .A(u0__abc_49347_n4560_bF_buf3), .B(u0_csc0_25_), .Y(u0__abc_49347_n5450) );
  AND2X2 AND2X2_1733 ( .A(u0__abc_49347_n4511_bF_buf3), .B(_auto_iopadmap_cc_313_execute_56321_25_), .Y(u0__abc_49347_n5451) );
  AND2X2 AND2X2_1734 ( .A(u0__abc_49347_n4516_bF_buf3), .B(u0_tms1_25_), .Y(u0__abc_49347_n5452) );
  AND2X2 AND2X2_1735 ( .A(u0__abc_49347_n4519_bF_buf3), .B(u0_csc2_25_), .Y(u0__abc_49347_n5453) );
  AND2X2 AND2X2_1736 ( .A(u0__abc_49347_n4586_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n5457) );
  AND2X2 AND2X2_1737 ( .A(u0__abc_49347_n4584_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n5458) );
  AND2X2 AND2X2_1738 ( .A(u0__abc_49347_n4589_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n5459) );
  AND2X2 AND2X2_1739 ( .A(u0__abc_49347_n4562_bF_buf3), .B(u0_csc5_25_), .Y(u0__abc_49347_n5462) );
  AND2X2 AND2X2_174 ( .A(u0__abc_49347_n1299_1), .B(u0__abc_49347_n1301), .Y(u0__abc_49347_n1302) );
  AND2X2 AND2X2_1740 ( .A(u0__abc_49347_n4571_bF_buf3), .B(u0_tms5_25_), .Y(u0__abc_49347_n5463) );
  AND2X2 AND2X2_1741 ( .A(u0__abc_49347_n4567_bF_buf3), .B(u0_tms4_25_), .Y(u0__abc_49347_n5465) );
  AND2X2 AND2X2_1742 ( .A(u0__abc_49347_n4507_bF_buf2), .B(rfr_ps_val_1_), .Y(u0__abc_49347_n5466) );
  AND2X2 AND2X2_1743 ( .A(u0__abc_49347_n4582_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n5473) );
  AND2X2 AND2X2_1744 ( .A(u0__abc_49347_n4531_bF_buf2), .B(u0_csc4_26_), .Y(u0__abc_49347_n5474) );
  AND2X2 AND2X2_1745 ( .A(u0__abc_49347_n4535_bF_buf2), .B(u0_tms0_26_), .Y(u0__abc_49347_n5475) );
  AND2X2 AND2X2_1746 ( .A(u0__abc_49347_n4537_bF_buf2), .B(u0_tms2_26_), .Y(u0__abc_49347_n5477) );
  AND2X2 AND2X2_1747 ( .A(u0__abc_49347_n4526_bF_buf2), .B(u0_csc1_26_), .Y(u0__abc_49347_n5478) );
  AND2X2 AND2X2_1748 ( .A(u0__abc_49347_n4528_bF_buf2), .B(u0_tms3_26_), .Y(u0__abc_49347_n5480) );
  AND2X2 AND2X2_1749 ( .A(u0__abc_49347_n4560_bF_buf2), .B(u0_csc0_26_), .Y(u0__abc_49347_n5481) );
  AND2X2 AND2X2_175 ( .A(u0__abc_49347_n1176_1_bF_buf1), .B(sp_tms_5_), .Y(u0__abc_49347_n1304) );
  AND2X2 AND2X2_1750 ( .A(u0__abc_49347_n4507_bF_buf1), .B(rfr_ps_val_2_), .Y(u0__abc_49347_n5485) );
  AND2X2 AND2X2_1751 ( .A(u0__abc_49347_n4589_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n5486) );
  AND2X2 AND2X2_1752 ( .A(u0__abc_49347_n4571_bF_buf2), .B(u0_tms5_26_), .Y(u0__abc_49347_n5487) );
  AND2X2 AND2X2_1753 ( .A(u0__abc_49347_n4584_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n5490) );
  AND2X2 AND2X2_1754 ( .A(u0__abc_49347_n4586_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n5491) );
  AND2X2 AND2X2_1755 ( .A(u0__abc_49347_n4567_bF_buf2), .B(u0_tms4_26_), .Y(u0__abc_49347_n5493) );
  AND2X2 AND2X2_1756 ( .A(u0__abc_49347_n4562_bF_buf2), .B(u0_csc5_26_), .Y(u0__abc_49347_n5494) );
  AND2X2 AND2X2_1757 ( .A(u0__abc_49347_n4539_bF_buf2), .B(u0_csc3_26_), .Y(u0__abc_49347_n5497) );
  AND2X2 AND2X2_1758 ( .A(u0__abc_49347_n4516_bF_buf2), .B(u0_tms1_26_), .Y(u0__abc_49347_n5498) );
  AND2X2 AND2X2_1759 ( .A(u0__abc_49347_n4519_bF_buf2), .B(u0_csc2_26_), .Y(u0__abc_49347_n5500) );
  AND2X2 AND2X2_176 ( .A(spec_req_cs_5_bF_buf3), .B(u0_tms5_5_), .Y(u0__abc_49347_n1305) );
  AND2X2 AND2X2_1760 ( .A(u0__abc_49347_n4511_bF_buf2), .B(_auto_iopadmap_cc_313_execute_56321_26_), .Y(u0__abc_49347_n5501) );
  AND2X2 AND2X2_1761 ( .A(u0__abc_49347_n4582_bF_buf2), .B(1'b0), .Y(u0__abc_49347_n5508) );
  AND2X2 AND2X2_1762 ( .A(u0__abc_49347_n4586_bF_buf2), .B(1'b0), .Y(u0__abc_49347_n5509) );
  AND2X2 AND2X2_1763 ( .A(u0__abc_49347_n4584_bF_buf2), .B(1'b0), .Y(u0__abc_49347_n5510) );
  AND2X2 AND2X2_1764 ( .A(u0__abc_49347_n4589_bF_buf2), .B(1'b0), .Y(u0__abc_49347_n5511) );
  AND2X2 AND2X2_1765 ( .A(u0__abc_49347_n4571_bF_buf1), .B(u0_tms5_27_), .Y(u0__abc_49347_n5514) );
  AND2X2 AND2X2_1766 ( .A(u0__abc_49347_n4567_bF_buf1), .B(u0_tms4_27_), .Y(u0__abc_49347_n5515) );
  AND2X2 AND2X2_1767 ( .A(u0__abc_49347_n4507_bF_buf0), .B(rfr_ps_val_3_), .Y(u0__abc_49347_n5516) );
  AND2X2 AND2X2_1768 ( .A(u0__abc_49347_n4526_bF_buf1), .B(u0_csc1_27_), .Y(u0__abc_49347_n5520) );
  AND2X2 AND2X2_1769 ( .A(u0__abc_49347_n4528_bF_buf1), .B(u0_tms3_27_), .Y(u0__abc_49347_n5521) );
  AND2X2 AND2X2_177 ( .A(u0__abc_49347_n1307), .B(u0__abc_49347_n1185_bF_buf0), .Y(u0__abc_49347_n1308_1) );
  AND2X2 AND2X2_1770 ( .A(u0__abc_49347_n4531_bF_buf1), .B(u0_csc4_27_), .Y(u0__abc_49347_n5522) );
  AND2X2 AND2X2_1771 ( .A(u0__abc_49347_n4535_bF_buf1), .B(u0_tms0_27_), .Y(u0__abc_49347_n5525) );
  AND2X2 AND2X2_1772 ( .A(u0__abc_49347_n4539_bF_buf1), .B(u0_csc3_27_), .Y(u0__abc_49347_n5526) );
  AND2X2 AND2X2_1773 ( .A(u0__abc_49347_n4537_bF_buf1), .B(u0_tms2_27_), .Y(u0__abc_49347_n5527) );
  AND2X2 AND2X2_1774 ( .A(u0__abc_49347_n4560_bF_buf1), .B(u0_csc0_27_), .Y(u0__abc_49347_n5531) );
  AND2X2 AND2X2_1775 ( .A(u0__abc_49347_n4516_bF_buf1), .B(u0_tms1_27_), .Y(u0__abc_49347_n5532) );
  AND2X2 AND2X2_1776 ( .A(u0__abc_49347_n4519_bF_buf1), .B(u0_csc2_27_), .Y(u0__abc_49347_n5533) );
  AND2X2 AND2X2_1777 ( .A(u0__abc_49347_n4562_bF_buf1), .B(u0_csc5_27_), .Y(u0__abc_49347_n5536) );
  AND2X2 AND2X2_1778 ( .A(u0__abc_49347_n4511_bF_buf1), .B(_auto_iopadmap_cc_313_execute_56321_27_), .Y(u0__abc_49347_n5537) );
  AND2X2 AND2X2_1779 ( .A(u0__abc_49347_n4582_bF_buf1), .B(1'b0), .Y(u0__abc_49347_n5543) );
  AND2X2 AND2X2_178 ( .A(u0__abc_49347_n1308_1), .B(u0__abc_49347_n1306), .Y(u0__abc_49347_n1309_1) );
  AND2X2 AND2X2_1780 ( .A(u0__abc_49347_n4535_bF_buf0), .B(u0_tms0_28_), .Y(u0__abc_49347_n5544) );
  AND2X2 AND2X2_1781 ( .A(u0__abc_49347_n4531_bF_buf0), .B(u0_csc4_28_), .Y(u0__abc_49347_n5545) );
  AND2X2 AND2X2_1782 ( .A(u0__abc_49347_n4528_bF_buf0), .B(u0_tms3_28_), .Y(u0__abc_49347_n5546) );
  AND2X2 AND2X2_1783 ( .A(u0__abc_49347_n4526_bF_buf0), .B(u0_csc1_28_), .Y(u0__abc_49347_n5549) );
  AND2X2 AND2X2_1784 ( .A(u0__abc_49347_n4537_bF_buf0), .B(u0_tms2_28_), .Y(u0__abc_49347_n5550) );
  AND2X2 AND2X2_1785 ( .A(u0__abc_49347_n4539_bF_buf0), .B(u0_csc3_28_), .Y(u0__abc_49347_n5551) );
  AND2X2 AND2X2_1786 ( .A(u0__abc_49347_n4511_bF_buf0), .B(_auto_iopadmap_cc_313_execute_56321_28_), .Y(u0__abc_49347_n5555) );
  AND2X2 AND2X2_1787 ( .A(u0__abc_49347_n4560_bF_buf0), .B(u0_csc0_28_), .Y(u0__abc_49347_n5556) );
  AND2X2 AND2X2_1788 ( .A(u0__abc_49347_n4516_bF_buf0), .B(u0_tms1_28_), .Y(u0__abc_49347_n5557) );
  AND2X2 AND2X2_1789 ( .A(u0__abc_49347_n4519_bF_buf0), .B(u0_csc2_28_), .Y(u0__abc_49347_n5558) );
  AND2X2 AND2X2_179 ( .A(u0__abc_49347_n1310), .B(u0__abc_49347_n1181_bF_buf0), .Y(u0__abc_49347_n1311) );
  AND2X2 AND2X2_1790 ( .A(u0__abc_49347_n4586_bF_buf1), .B(1'b0), .Y(u0__abc_49347_n5562) );
  AND2X2 AND2X2_1791 ( .A(u0__abc_49347_n4584_bF_buf1), .B(1'b0), .Y(u0__abc_49347_n5563) );
  AND2X2 AND2X2_1792 ( .A(u0__abc_49347_n4589_bF_buf1), .B(1'b0), .Y(u0__abc_49347_n5564) );
  AND2X2 AND2X2_1793 ( .A(u0__abc_49347_n4562_bF_buf0), .B(u0_csc5_28_), .Y(u0__abc_49347_n5567) );
  AND2X2 AND2X2_1794 ( .A(u0__abc_49347_n4571_bF_buf0), .B(u0_tms5_28_), .Y(u0__abc_49347_n5568) );
  AND2X2 AND2X2_1795 ( .A(u0__abc_49347_n4567_bF_buf0), .B(u0_tms4_28_), .Y(u0__abc_49347_n5570) );
  AND2X2 AND2X2_1796 ( .A(u0__abc_49347_n4507_bF_buf3), .B(rfr_ps_val_4_), .Y(u0__abc_49347_n5571) );
  AND2X2 AND2X2_1797 ( .A(u0__abc_49347_n4526_bF_buf4), .B(u0_csc1_29_), .Y(u0__abc_49347_n5578) );
  AND2X2 AND2X2_1798 ( .A(u0__abc_49347_n4531_bF_buf4), .B(u0_csc4_29_), .Y(u0__abc_49347_n5579) );
  AND2X2 AND2X2_1799 ( .A(u0__abc_49347_n4528_bF_buf4), .B(u0_tms3_29_), .Y(u0__abc_49347_n5581) );
  AND2X2 AND2X2_18 ( .A(_abc_55805_n290), .B(_abc_55805_n291), .Y(tms_s_0_) );
  AND2X2 AND2X2_180 ( .A(spec_req_cs_4_bF_buf3), .B(u0_tms4_5_), .Y(u0__abc_49347_n1312) );
  AND2X2 AND2X2_1800 ( .A(u0__abc_49347_n4539_bF_buf4), .B(u0_csc3_29_), .Y(u0__abc_49347_n5582) );
  AND2X2 AND2X2_1801 ( .A(u0__abc_49347_n4535_bF_buf4), .B(u0_tms0_29_), .Y(u0__abc_49347_n5584) );
  AND2X2 AND2X2_1802 ( .A(u0__abc_49347_n4537_bF_buf4), .B(u0_tms2_29_), .Y(u0__abc_49347_n5585) );
  AND2X2 AND2X2_1803 ( .A(u0__abc_49347_n4586_bF_buf0), .B(1'b0), .Y(u0__abc_49347_n5589) );
  AND2X2 AND2X2_1804 ( .A(u0__abc_49347_n4589_bF_buf0), .B(1'b0), .Y(u0__abc_49347_n5590) );
  AND2X2 AND2X2_1805 ( .A(u0__abc_49347_n4584_bF_buf0), .B(1'b0), .Y(u0__abc_49347_n5591) );
  AND2X2 AND2X2_1806 ( .A(u0__abc_49347_n4571_bF_buf4), .B(u0_tms5_29_), .Y(u0__abc_49347_n5594) );
  AND2X2 AND2X2_1807 ( .A(u0__abc_49347_n4507_bF_buf2), .B(rfr_ps_val_5_), .Y(u0__abc_49347_n5595) );
  AND2X2 AND2X2_1808 ( .A(u0__abc_49347_n4567_bF_buf4), .B(u0_tms4_29_), .Y(u0__abc_49347_n5596) );
  AND2X2 AND2X2_1809 ( .A(u0__abc_49347_n4582_bF_buf0), .B(1'b0), .Y(u0__abc_49347_n5601) );
  AND2X2 AND2X2_181 ( .A(u0__abc_49347_n1313), .B(u0__abc_49347_n1180_1_bF_buf0), .Y(u0__abc_49347_n1314) );
  AND2X2 AND2X2_1810 ( .A(u0__abc_49347_n4560_bF_buf4), .B(u0_csc0_29_), .Y(u0__abc_49347_n5602) );
  AND2X2 AND2X2_1811 ( .A(u0__abc_49347_n4516_bF_buf4), .B(u0_tms1_29_), .Y(u0__abc_49347_n5603) );
  AND2X2 AND2X2_1812 ( .A(u0__abc_49347_n4519_bF_buf4), .B(u0_csc2_29_), .Y(u0__abc_49347_n5604) );
  AND2X2 AND2X2_1813 ( .A(u0__abc_49347_n4511_bF_buf4), .B(_auto_iopadmap_cc_313_execute_56321_29_), .Y(u0__abc_49347_n5607) );
  AND2X2 AND2X2_1814 ( .A(u0__abc_49347_n4562_bF_buf4), .B(u0_csc5_29_), .Y(u0__abc_49347_n5608) );
  AND2X2 AND2X2_1815 ( .A(u0__abc_49347_n4582_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n5613) );
  AND2X2 AND2X2_1816 ( .A(u0__abc_49347_n4586_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n5614) );
  AND2X2 AND2X2_1817 ( .A(u0__abc_49347_n4584_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n5615) );
  AND2X2 AND2X2_1818 ( .A(u0__abc_49347_n4567_bF_buf3), .B(u0_tms4_30_), .Y(u0__abc_49347_n5617) );
  AND2X2 AND2X2_1819 ( .A(u0__abc_49347_n4589_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n5618) );
  AND2X2 AND2X2_182 ( .A(spec_req_cs_3_bF_buf3), .B(u0_tms3_5_), .Y(u0__abc_49347_n1315) );
  AND2X2 AND2X2_1820 ( .A(u0__abc_49347_n4507_bF_buf1), .B(rfr_ps_val_6_), .Y(u0__abc_49347_n5620) );
  AND2X2 AND2X2_1821 ( .A(u0__abc_49347_n4571_bF_buf3), .B(u0_tms5_30_), .Y(u0__abc_49347_n5621) );
  AND2X2 AND2X2_1822 ( .A(u0__abc_49347_n4535_bF_buf3), .B(u0_tms0_30_), .Y(u0__abc_49347_n5625) );
  AND2X2 AND2X2_1823 ( .A(u0__abc_49347_n4531_bF_buf3), .B(u0_csc4_30_), .Y(u0__abc_49347_n5626) );
  AND2X2 AND2X2_1824 ( .A(u0__abc_49347_n4528_bF_buf3), .B(u0_tms3_30_), .Y(u0__abc_49347_n5627) );
  AND2X2 AND2X2_1825 ( .A(u0__abc_49347_n4526_bF_buf3), .B(u0_csc1_30_), .Y(u0__abc_49347_n5630) );
  AND2X2 AND2X2_1826 ( .A(u0__abc_49347_n4537_bF_buf3), .B(u0_tms2_30_), .Y(u0__abc_49347_n5631) );
  AND2X2 AND2X2_1827 ( .A(u0__abc_49347_n4539_bF_buf3), .B(u0_csc3_30_), .Y(u0__abc_49347_n5632) );
  AND2X2 AND2X2_1828 ( .A(u0__abc_49347_n4560_bF_buf3), .B(u0_csc0_30_), .Y(u0__abc_49347_n5636) );
  AND2X2 AND2X2_1829 ( .A(u0__abc_49347_n4516_bF_buf3), .B(u0_tms1_30_), .Y(u0__abc_49347_n5637) );
  AND2X2 AND2X2_183 ( .A(u0__abc_49347_n1316), .B(u0__abc_49347_n1179_bF_buf0), .Y(u0__abc_49347_n1317_1) );
  AND2X2 AND2X2_1830 ( .A(u0__abc_49347_n4519_bF_buf3), .B(u0_csc2_30_), .Y(u0__abc_49347_n5638) );
  AND2X2 AND2X2_1831 ( .A(u0__abc_49347_n4511_bF_buf3), .B(_auto_iopadmap_cc_313_execute_56321_30_), .Y(u0__abc_49347_n5641) );
  AND2X2 AND2X2_1832 ( .A(u0__abc_49347_n4562_bF_buf3), .B(u0_csc5_30_), .Y(u0__abc_49347_n5642) );
  AND2X2 AND2X2_1833 ( .A(u0__abc_49347_n4582_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n5648) );
  AND2X2 AND2X2_1834 ( .A(u0__abc_49347_n4531_bF_buf2), .B(u0_csc4_31_), .Y(u0__abc_49347_n5649) );
  AND2X2 AND2X2_1835 ( .A(u0__abc_49347_n4526_bF_buf2), .B(u0_csc1_31_), .Y(u0__abc_49347_n5650) );
  AND2X2 AND2X2_1836 ( .A(u0__abc_49347_n4528_bF_buf2), .B(u0_tms3_31_), .Y(u0__abc_49347_n5652) );
  AND2X2 AND2X2_1837 ( .A(u0__abc_49347_n4537_bF_buf2), .B(u0_tms2_31_), .Y(u0__abc_49347_n5653) );
  AND2X2 AND2X2_1838 ( .A(u0__abc_49347_n4539_bF_buf2), .B(u0_csc3_31_), .Y(u0__abc_49347_n5655) );
  AND2X2 AND2X2_1839 ( .A(u0__abc_49347_n4535_bF_buf2), .B(u0_tms0_31_), .Y(u0__abc_49347_n5656) );
  AND2X2 AND2X2_184 ( .A(spec_req_cs_2_bF_buf3), .B(u0_tms2_5_), .Y(u0__abc_49347_n1318_1) );
  AND2X2 AND2X2_1840 ( .A(u0__abc_49347_n4511_bF_buf2), .B(_auto_iopadmap_cc_313_execute_56321_31_), .Y(u0__abc_49347_n5660) );
  AND2X2 AND2X2_1841 ( .A(u0__abc_49347_n4560_bF_buf2), .B(u0_csc0_31_), .Y(u0__abc_49347_n5661) );
  AND2X2 AND2X2_1842 ( .A(u0__abc_49347_n4516_bF_buf2), .B(u0_tms1_31_), .Y(u0__abc_49347_n5662) );
  AND2X2 AND2X2_1843 ( .A(u0__abc_49347_n4519_bF_buf2), .B(u0_csc2_31_), .Y(u0__abc_49347_n5663) );
  AND2X2 AND2X2_1844 ( .A(u0__abc_49347_n4589_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n5667) );
  AND2X2 AND2X2_1845 ( .A(u0__abc_49347_n4584_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n5668) );
  AND2X2 AND2X2_1846 ( .A(u0__abc_49347_n4586_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n5670) );
  AND2X2 AND2X2_1847 ( .A(u0__abc_49347_n4507_bF_buf0), .B(rfr_ps_val_7_), .Y(u0__abc_49347_n5672) );
  AND2X2 AND2X2_1848 ( .A(u0__abc_49347_n4567_bF_buf2), .B(u0_tms4_31_), .Y(u0__abc_49347_n5673) );
  AND2X2 AND2X2_1849 ( .A(u0__abc_49347_n4562_bF_buf2), .B(u0_csc5_31_), .Y(u0__abc_49347_n5675) );
  AND2X2 AND2X2_185 ( .A(u0__abc_49347_n1319), .B(u0__abc_49347_n1178_1_bF_buf0), .Y(u0__abc_49347_n1320) );
  AND2X2 AND2X2_1850 ( .A(u0__abc_49347_n4571_bF_buf2), .B(u0_tms5_31_), .Y(u0__abc_49347_n5676) );
  AND2X2 AND2X2_1851 ( .A(\wb_addr_i[29] ), .B(\wb_addr_i[30] ), .Y(u0__abc_49347_n5684) );
  AND2X2 AND2X2_1852 ( .A(u0__abc_49347_n5684), .B(u0__abc_49347_n5683), .Y(u0__abc_49347_n5685) );
  AND2X2 AND2X2_1853 ( .A(u0__abc_49347_n4400), .B(wb_we_i), .Y(u0__abc_49347_n5686) );
  AND2X2 AND2X2_1854 ( .A(u0__abc_49347_n5686), .B(u0__abc_49347_n1173), .Y(u0__abc_49347_n5687) );
  AND2X2 AND2X2_1855 ( .A(u0__abc_49347_n5687), .B(u0__abc_49347_n5685), .Y(u0_rf_we_FF_INPUT) );
  AND2X2 AND2X2_1856 ( .A(u0__abc_49347_n5692), .B(u0_csc0_0_), .Y(u0__abc_49347_n5693) );
  AND2X2 AND2X2_1857 ( .A(u0__abc_49347_n5694), .B(u0__abc_49347_n5695), .Y(u0__abc_49347_n5696) );
  AND2X2 AND2X2_1858 ( .A(u0__abc_49347_n5696), .B(u0__abc_49347_n5693), .Y(cs_need_rfr_0_) );
  AND2X2 AND2X2_1859 ( .A(u0__abc_49347_n5698), .B(u0_csc1_0_), .Y(u0__abc_49347_n5699) );
  AND2X2 AND2X2_186 ( .A(spec_req_cs_1_bF_buf3), .B(u0_tms1_5_), .Y(u0__abc_49347_n1321) );
  AND2X2 AND2X2_1860 ( .A(u0__abc_49347_n5700), .B(u0__abc_49347_n5701), .Y(u0__abc_49347_n5702) );
  AND2X2 AND2X2_1861 ( .A(u0__abc_49347_n5702), .B(u0__abc_49347_n5699), .Y(cs_need_rfr_1_) );
  AND2X2 AND2X2_1862 ( .A(u0__abc_49347_n5704), .B(u0_csc2_0_), .Y(u0__abc_49347_n5705) );
  AND2X2 AND2X2_1863 ( .A(u0__abc_49347_n5706), .B(u0__abc_49347_n5707), .Y(u0__abc_49347_n5708) );
  AND2X2 AND2X2_1864 ( .A(u0__abc_49347_n5708), .B(u0__abc_49347_n5705), .Y(cs_need_rfr_2_) );
  AND2X2 AND2X2_1865 ( .A(u0__abc_49347_n5710), .B(u0_csc3_0_), .Y(u0__abc_49347_n5711) );
  AND2X2 AND2X2_1866 ( .A(u0__abc_49347_n5712), .B(u0__abc_49347_n5713), .Y(u0__abc_49347_n5714) );
  AND2X2 AND2X2_1867 ( .A(u0__abc_49347_n5714), .B(u0__abc_49347_n5711), .Y(cs_need_rfr_3_) );
  AND2X2 AND2X2_1868 ( .A(u0__abc_49347_n5716), .B(u0_csc4_0_), .Y(u0__abc_49347_n5717) );
  AND2X2 AND2X2_1869 ( .A(u0__abc_49347_n5718), .B(u0__abc_49347_n5719), .Y(u0__abc_49347_n5720) );
  AND2X2 AND2X2_187 ( .A(u0__abc_49347_n1175_bF_buf0), .B(u0__abc_49347_n1324), .Y(u0__abc_49347_n1325) );
  AND2X2 AND2X2_1870 ( .A(u0__abc_49347_n5720), .B(u0__abc_49347_n5717), .Y(cs_need_rfr_4_) );
  AND2X2 AND2X2_1871 ( .A(u0__abc_49347_n5722), .B(u0_csc5_0_), .Y(u0__abc_49347_n5723) );
  AND2X2 AND2X2_1872 ( .A(u0__abc_49347_n5724), .B(u0__abc_49347_n5725), .Y(u0__abc_49347_n5726) );
  AND2X2 AND2X2_1873 ( .A(u0__abc_49347_n5726), .B(u0__abc_49347_n5723), .Y(cs_need_rfr_5_) );
  AND2X2 AND2X2_1874 ( .A(u0__abc_49347_n5728), .B(1'b0), .Y(u0__abc_49347_n5729) );
  AND2X2 AND2X2_1875 ( .A(u0__abc_49347_n5730), .B(u0__abc_49347_n5731), .Y(u0__abc_49347_n5732) );
  AND2X2 AND2X2_1876 ( .A(u0__abc_49347_n5732), .B(u0__abc_49347_n5729), .Y(cs_need_rfr_6_) );
  AND2X2 AND2X2_1877 ( .A(u0__abc_49347_n5734), .B(1'b0), .Y(u0__abc_49347_n5735) );
  AND2X2 AND2X2_1878 ( .A(u0__abc_49347_n5736), .B(u0__abc_49347_n5737), .Y(u0__abc_49347_n5738) );
  AND2X2 AND2X2_1879 ( .A(u0__abc_49347_n5738), .B(u0__abc_49347_n5735), .Y(cs_need_rfr_7_) );
  AND2X2 AND2X2_188 ( .A(u0__abc_49347_n1323), .B(u0__abc_49347_n1325), .Y(u0__abc_49347_n1326_1) );
  AND2X2 AND2X2_1880 ( .A(u0__abc_49347_n1100_1), .B(u0__abc_49347_n5740), .Y(u0__abc_49347_n5741) );
  AND2X2 AND2X2_1881 ( .A(u0__abc_49347_n5742), .B(u0_init_ack_r), .Y(u0__abc_49347_n5743) );
  AND2X2 AND2X2_1882 ( .A(u0__abc_49347_n5744), .B(u0_lmr_ack_r), .Y(u0__abc_49347_n5745) );
  AND2X2 AND2X2_1883 ( .A(u0__abc_49347_n5745), .B(spec_req_cs_0_bF_buf1), .Y(u0_lmr_ack0) );
  AND2X2 AND2X2_1884 ( .A(u0__abc_49347_n5745), .B(spec_req_cs_1_bF_buf1), .Y(u0_lmr_ack1) );
  AND2X2 AND2X2_1885 ( .A(u0__abc_49347_n5745), .B(spec_req_cs_2_bF_buf1), .Y(u0_lmr_ack2) );
  AND2X2 AND2X2_1886 ( .A(u0__abc_49347_n5745), .B(spec_req_cs_3_bF_buf1), .Y(u0_lmr_ack3) );
  AND2X2 AND2X2_1887 ( .A(u0__abc_49347_n5745), .B(spec_req_cs_4_bF_buf1), .Y(u0_lmr_ack4) );
  AND2X2 AND2X2_1888 ( .A(u0__abc_49347_n5745), .B(spec_req_cs_5_bF_buf1), .Y(u0_lmr_ack5) );
  AND2X2 AND2X2_1889 ( .A(u0__abc_49347_n5743), .B(spec_req_cs_0_bF_buf0), .Y(u0_init_ack0) );
  AND2X2 AND2X2_189 ( .A(u0__abc_49347_n1176_1_bF_buf0), .B(sp_tms_6_), .Y(u0__abc_49347_n1328) );
  AND2X2 AND2X2_1890 ( .A(u0__abc_49347_n5743), .B(spec_req_cs_1_bF_buf0), .Y(u0_init_ack1) );
  AND2X2 AND2X2_1891 ( .A(u0__abc_49347_n5743), .B(spec_req_cs_2_bF_buf0), .Y(u0_init_ack2) );
  AND2X2 AND2X2_1892 ( .A(u0__abc_49347_n5743), .B(spec_req_cs_3_bF_buf0), .Y(u0_init_ack3) );
  AND2X2 AND2X2_1893 ( .A(u0__abc_49347_n5743), .B(spec_req_cs_4_bF_buf0), .Y(u0_init_ack4) );
  AND2X2 AND2X2_1894 ( .A(u0__abc_49347_n5743), .B(spec_req_cs_5_bF_buf0), .Y(u0_init_ack5) );
  AND2X2 AND2X2_1895 ( .A(u0_u0__abc_43300_n203), .B(u0_u0_lmr_req_we), .Y(u0_u0__abc_43300_n204_1) );
  AND2X2 AND2X2_1896 ( .A(u0_u0__abc_43300_n204_1), .B(u0_u0_inited), .Y(u0_u0__abc_43300_n205_1) );
  AND2X2 AND2X2_1897 ( .A(u0_u0__abc_43300_n207_1), .B(u0_lmr_req0), .Y(u0_u0__abc_43300_n208_1) );
  AND2X2 AND2X2_1898 ( .A(u0_u0__abc_43300_n206), .B(u0_u0__abc_43300_n208_1), .Y(u0_u0__abc_43300_n209) );
  AND2X2 AND2X2_1899 ( .A(u0_u0_addr_r_4_), .B(u0_rf_we), .Y(u0_u0__abc_43300_n211_1) );
  AND2X2 AND2X2_19 ( .A(_abc_55805_n293), .B(_abc_55805_n294), .Y(tms_s_1_) );
  AND2X2 AND2X2_190 ( .A(spec_req_cs_5_bF_buf2), .B(u0_tms5_6_), .Y(u0__abc_49347_n1329) );
  AND2X2 AND2X2_1900 ( .A(u0_u0__abc_43300_n214_1), .B(u0_u0__abc_43300_n211_1), .Y(u0_u0__abc_43300_n215) );
  AND2X2 AND2X2_1901 ( .A(u0_u0__abc_43300_n215), .B(u0_u0_addr_r_2_), .Y(u0_u0_lmr_req_we_FF_INPUT) );
  AND2X2 AND2X2_1902 ( .A(u0_u0__abc_43300_n220_1), .B(u0_u0__abc_43300_n218_bF_buf7), .Y(u0_u0__abc_43300_n221) );
  AND2X2 AND2X2_1903 ( .A(u0_u0__abc_43300_n221), .B(u0_u0__abc_43300_n217_1), .Y(u0_u0_tms_0__FF_INPUT) );
  AND2X2 AND2X2_1904 ( .A(u0_u0__abc_43300_n224), .B(u0_u0__abc_43300_n218_bF_buf6), .Y(u0_u0__abc_43300_n225_1) );
  AND2X2 AND2X2_1905 ( .A(u0_u0__abc_43300_n225_1), .B(u0_u0__abc_43300_n223_1), .Y(u0_u0_tms_1__FF_INPUT) );
  AND2X2 AND2X2_1906 ( .A(u0_u0__abc_43300_n228_1), .B(u0_u0__abc_43300_n218_bF_buf5), .Y(u0_u0__abc_43300_n229_1) );
  AND2X2 AND2X2_1907 ( .A(u0_u0__abc_43300_n229_1), .B(u0_u0__abc_43300_n227), .Y(u0_u0_tms_2__FF_INPUT) );
  AND2X2 AND2X2_1908 ( .A(u0_u0__abc_43300_n232_1), .B(u0_u0__abc_43300_n218_bF_buf4), .Y(u0_u0__abc_43300_n233) );
  AND2X2 AND2X2_1909 ( .A(u0_u0__abc_43300_n233), .B(u0_u0__abc_43300_n231_1), .Y(u0_u0_tms_3__FF_INPUT) );
  AND2X2 AND2X2_191 ( .A(u0__abc_49347_n1331), .B(u0__abc_49347_n1185_bF_buf5), .Y(u0__abc_49347_n1332) );
  AND2X2 AND2X2_1910 ( .A(u0_u0__abc_43300_n236), .B(u0_u0__abc_43300_n218_bF_buf3), .Y(u0_u0__abc_43300_n237_1) );
  AND2X2 AND2X2_1911 ( .A(u0_u0__abc_43300_n237_1), .B(u0_u0__abc_43300_n235_1), .Y(u0_u0_tms_4__FF_INPUT) );
  AND2X2 AND2X2_1912 ( .A(u0_u0__abc_43300_n240_1), .B(u0_u0__abc_43300_n218_bF_buf2), .Y(u0_u0__abc_43300_n241_1) );
  AND2X2 AND2X2_1913 ( .A(u0_u0__abc_43300_n241_1), .B(u0_u0__abc_43300_n239), .Y(u0_u0_tms_5__FF_INPUT) );
  AND2X2 AND2X2_1914 ( .A(u0_u0__abc_43300_n244_1), .B(u0_u0__abc_43300_n218_bF_buf1), .Y(u0_u0__abc_43300_n245) );
  AND2X2 AND2X2_1915 ( .A(u0_u0__abc_43300_n245), .B(u0_u0__abc_43300_n243_1), .Y(u0_u0_tms_6__FF_INPUT) );
  AND2X2 AND2X2_1916 ( .A(u0_u0__abc_43300_n248), .B(u0_u0__abc_43300_n218_bF_buf0), .Y(u0_u0__abc_43300_n249_1) );
  AND2X2 AND2X2_1917 ( .A(u0_u0__abc_43300_n249_1), .B(u0_u0__abc_43300_n247_1), .Y(u0_u0_tms_7__FF_INPUT) );
  AND2X2 AND2X2_1918 ( .A(u0_u0__abc_43300_n252_1), .B(u0_u0__abc_43300_n218_bF_buf7), .Y(u0_u0__abc_43300_n253_1) );
  AND2X2 AND2X2_1919 ( .A(u0_u0__abc_43300_n253_1), .B(u0_u0__abc_43300_n251), .Y(u0_u0_tms_8__FF_INPUT) );
  AND2X2 AND2X2_192 ( .A(u0__abc_49347_n1332), .B(u0__abc_49347_n1330), .Y(u0__abc_49347_n1333) );
  AND2X2 AND2X2_1920 ( .A(u0_u0__abc_43300_n256), .B(u0_u0__abc_43300_n218_bF_buf6), .Y(u0_u0__abc_43300_n257) );
  AND2X2 AND2X2_1921 ( .A(u0_u0__abc_43300_n257), .B(u0_u0__abc_43300_n255_1), .Y(u0_u0_tms_9__FF_INPUT) );
  AND2X2 AND2X2_1922 ( .A(u0_u0__abc_43300_n260_1), .B(u0_u0__abc_43300_n218_bF_buf5), .Y(u0_u0__abc_43300_n261) );
  AND2X2 AND2X2_1923 ( .A(u0_u0__abc_43300_n261), .B(u0_u0__abc_43300_n259), .Y(u0_u0_tms_10__FF_INPUT) );
  AND2X2 AND2X2_1924 ( .A(u0_u0__abc_43300_n264), .B(u0_u0__abc_43300_n218_bF_buf4), .Y(u0_u0__abc_43300_n265) );
  AND2X2 AND2X2_1925 ( .A(u0_u0__abc_43300_n265), .B(u0_u0__abc_43300_n263), .Y(u0_u0_tms_11__FF_INPUT) );
  AND2X2 AND2X2_1926 ( .A(u0_u0__abc_43300_n268_1), .B(u0_u0__abc_43300_n218_bF_buf3), .Y(u0_u0__abc_43300_n269) );
  AND2X2 AND2X2_1927 ( .A(u0_u0__abc_43300_n269), .B(u0_u0__abc_43300_n267), .Y(u0_u0_tms_12__FF_INPUT) );
  AND2X2 AND2X2_1928 ( .A(u0_u0__abc_43300_n272), .B(u0_u0__abc_43300_n218_bF_buf2), .Y(u0_u0__abc_43300_n273_1) );
  AND2X2 AND2X2_1929 ( .A(u0_u0__abc_43300_n273_1), .B(u0_u0__abc_43300_n271), .Y(u0_u0_tms_13__FF_INPUT) );
  AND2X2 AND2X2_193 ( .A(u0__abc_49347_n1334), .B(u0__abc_49347_n1181_bF_buf5), .Y(u0__abc_49347_n1335_1) );
  AND2X2 AND2X2_1930 ( .A(u0_u0__abc_43300_n276), .B(u0_u0__abc_43300_n218_bF_buf1), .Y(u0_u0__abc_43300_n277_1) );
  AND2X2 AND2X2_1931 ( .A(u0_u0__abc_43300_n277_1), .B(u0_u0__abc_43300_n275_1), .Y(u0_u0_tms_14__FF_INPUT) );
  AND2X2 AND2X2_1932 ( .A(u0_u0__abc_43300_n280), .B(u0_u0__abc_43300_n218_bF_buf0), .Y(u0_u0__abc_43300_n281) );
  AND2X2 AND2X2_1933 ( .A(u0_u0__abc_43300_n281), .B(u0_u0__abc_43300_n279_1), .Y(u0_u0_tms_15__FF_INPUT) );
  AND2X2 AND2X2_1934 ( .A(u0_u0__abc_43300_n284), .B(u0_u0__abc_43300_n218_bF_buf7), .Y(u0_u0__abc_43300_n285_1) );
  AND2X2 AND2X2_1935 ( .A(u0_u0__abc_43300_n285_1), .B(u0_u0__abc_43300_n283_1), .Y(u0_u0_tms_16__FF_INPUT) );
  AND2X2 AND2X2_1936 ( .A(u0_u0__abc_43300_n288), .B(u0_u0__abc_43300_n218_bF_buf6), .Y(u0_u0__abc_43300_n289_1) );
  AND2X2 AND2X2_1937 ( .A(u0_u0__abc_43300_n289_1), .B(u0_u0__abc_43300_n287_1), .Y(u0_u0_tms_17__FF_INPUT) );
  AND2X2 AND2X2_1938 ( .A(u0_u0__abc_43300_n292), .B(u0_u0__abc_43300_n218_bF_buf5), .Y(u0_u0__abc_43300_n293) );
  AND2X2 AND2X2_1939 ( .A(u0_u0__abc_43300_n293), .B(u0_u0__abc_43300_n291), .Y(u0_u0_tms_18__FF_INPUT) );
  AND2X2 AND2X2_194 ( .A(spec_req_cs_4_bF_buf2), .B(u0_tms4_6_), .Y(u0__abc_49347_n1336_1) );
  AND2X2 AND2X2_1940 ( .A(u0_u0__abc_43300_n296_1), .B(u0_u0__abc_43300_n218_bF_buf4), .Y(u0_u0__abc_43300_n297) );
  AND2X2 AND2X2_1941 ( .A(u0_u0__abc_43300_n297), .B(u0_u0__abc_43300_n295), .Y(u0_u0_tms_19__FF_INPUT) );
  AND2X2 AND2X2_1942 ( .A(u0_u0__abc_43300_n300), .B(u0_u0__abc_43300_n218_bF_buf3), .Y(u0_u0__abc_43300_n301) );
  AND2X2 AND2X2_1943 ( .A(u0_u0__abc_43300_n301), .B(u0_u0__abc_43300_n299), .Y(u0_u0_tms_20__FF_INPUT) );
  AND2X2 AND2X2_1944 ( .A(u0_u0__abc_43300_n304), .B(u0_u0__abc_43300_n218_bF_buf2), .Y(u0_u0__abc_43300_n305) );
  AND2X2 AND2X2_1945 ( .A(u0_u0__abc_43300_n305), .B(u0_u0__abc_43300_n303), .Y(u0_u0_tms_21__FF_INPUT) );
  AND2X2 AND2X2_1946 ( .A(u0_u0__abc_43300_n308), .B(u0_u0__abc_43300_n218_bF_buf1), .Y(u0_u0__abc_43300_n309) );
  AND2X2 AND2X2_1947 ( .A(u0_u0__abc_43300_n309), .B(u0_u0__abc_43300_n307), .Y(u0_u0_tms_22__FF_INPUT) );
  AND2X2 AND2X2_1948 ( .A(u0_u0__abc_43300_n312_1), .B(u0_u0__abc_43300_n218_bF_buf0), .Y(u0_u0__abc_43300_n313) );
  AND2X2 AND2X2_1949 ( .A(u0_u0__abc_43300_n313), .B(u0_u0__abc_43300_n311), .Y(u0_u0_tms_23__FF_INPUT) );
  AND2X2 AND2X2_195 ( .A(u0__abc_49347_n1337), .B(u0__abc_49347_n1180_1_bF_buf5), .Y(u0__abc_49347_n1338) );
  AND2X2 AND2X2_1950 ( .A(u0_u0__abc_43300_n316_1), .B(u0_u0__abc_43300_n218_bF_buf7), .Y(u0_u0__abc_43300_n317_1) );
  AND2X2 AND2X2_1951 ( .A(u0_u0__abc_43300_n317_1), .B(u0_u0__abc_43300_n315_1), .Y(u0_u0_tms_24__FF_INPUT) );
  AND2X2 AND2X2_1952 ( .A(u0_u0__abc_43300_n320), .B(u0_u0__abc_43300_n218_bF_buf6), .Y(u0_u0__abc_43300_n321_1) );
  AND2X2 AND2X2_1953 ( .A(u0_u0__abc_43300_n321_1), .B(u0_u0__abc_43300_n319), .Y(u0_u0_tms_25__FF_INPUT) );
  AND2X2 AND2X2_1954 ( .A(u0_u0__abc_43300_n324_1), .B(u0_u0__abc_43300_n218_bF_buf5), .Y(u0_u0__abc_43300_n325_1) );
  AND2X2 AND2X2_1955 ( .A(u0_u0__abc_43300_n325_1), .B(u0_u0__abc_43300_n323_1), .Y(u0_u0_tms_26__FF_INPUT) );
  AND2X2 AND2X2_1956 ( .A(u0_u0__abc_43300_n328), .B(u0_u0__abc_43300_n218_bF_buf4), .Y(u0_u0__abc_43300_n329) );
  AND2X2 AND2X2_1957 ( .A(u0_u0__abc_43300_n329), .B(u0_u0__abc_43300_n327), .Y(u0_u0_tms_27__FF_INPUT) );
  AND2X2 AND2X2_1958 ( .A(u0_u0__abc_43300_n332), .B(u0_u0__abc_43300_n218_bF_buf3), .Y(u0_u0__abc_43300_n333) );
  AND2X2 AND2X2_1959 ( .A(u0_u0__abc_43300_n333), .B(u0_u0__abc_43300_n331), .Y(u0_u0_tms_28__FF_INPUT) );
  AND2X2 AND2X2_196 ( .A(spec_req_cs_3_bF_buf2), .B(u0_tms3_6_), .Y(u0__abc_49347_n1339) );
  AND2X2 AND2X2_1960 ( .A(u0_u0__abc_43300_n336), .B(u0_u0__abc_43300_n218_bF_buf2), .Y(u0_u0__abc_43300_n337) );
  AND2X2 AND2X2_1961 ( .A(u0_u0__abc_43300_n337), .B(u0_u0__abc_43300_n335), .Y(u0_u0_tms_29__FF_INPUT) );
  AND2X2 AND2X2_1962 ( .A(u0_u0__abc_43300_n340), .B(u0_u0__abc_43300_n218_bF_buf1), .Y(u0_u0__abc_43300_n341) );
  AND2X2 AND2X2_1963 ( .A(u0_u0__abc_43300_n341), .B(u0_u0__abc_43300_n339), .Y(u0_u0_tms_30__FF_INPUT) );
  AND2X2 AND2X2_1964 ( .A(u0_u0__abc_43300_n344), .B(u0_u0__abc_43300_n218_bF_buf0), .Y(u0_u0__abc_43300_n345) );
  AND2X2 AND2X2_1965 ( .A(u0_u0__abc_43300_n345), .B(u0_u0__abc_43300_n343), .Y(u0_u0_tms_31__FF_INPUT) );
  AND2X2 AND2X2_1966 ( .A(u0_u0__abc_43300_n215), .B(u0_u0__abc_43300_n347), .Y(u0_u0_init_req_we_FF_INPUT) );
  AND2X2 AND2X2_1967 ( .A(u0_u0__abc_43300_n351), .B(u0_u0__abc_43300_n218_bF_buf7), .Y(u0_u0__abc_43300_n352) );
  AND2X2 AND2X2_1968 ( .A(u0_u0__abc_43300_n352), .B(u0_u0__abc_43300_n349), .Y(u0_u0_csc_0__FF_INPUT) );
  AND2X2 AND2X2_1969 ( .A(u0_u0__abc_43300_n355), .B(u0_u0__abc_43300_n218_bF_buf6), .Y(u0_u0__abc_43300_n356) );
  AND2X2 AND2X2_197 ( .A(u0__abc_49347_n1340), .B(u0__abc_49347_n1179_bF_buf5), .Y(u0__abc_49347_n1341) );
  AND2X2 AND2X2_1970 ( .A(u0_u0__abc_43300_n356), .B(u0_u0__abc_43300_n354), .Y(u0_u0_csc_1__FF_INPUT) );
  AND2X2 AND2X2_1971 ( .A(u0_u0__abc_43300_n359), .B(u0_u0__abc_43300_n218_bF_buf5), .Y(u0_u0__abc_43300_n360) );
  AND2X2 AND2X2_1972 ( .A(u0_u0__abc_43300_n360), .B(u0_u0__abc_43300_n358), .Y(u0_u0_csc_2__FF_INPUT) );
  AND2X2 AND2X2_1973 ( .A(u0_u0__abc_43300_n363), .B(u0_u0__abc_43300_n218_bF_buf4), .Y(u0_u0__abc_43300_n364) );
  AND2X2 AND2X2_1974 ( .A(u0_u0__abc_43300_n364), .B(u0_u0__abc_43300_n362), .Y(u0_u0_csc_3__FF_INPUT) );
  AND2X2 AND2X2_1975 ( .A(u0_u0__abc_43300_n367), .B(u0_u0__abc_43300_n218_bF_buf3), .Y(u0_u0__abc_43300_n368) );
  AND2X2 AND2X2_1976 ( .A(u0_u0__abc_43300_n368), .B(u0_u0__abc_43300_n366), .Y(u0_u0_csc_4__FF_INPUT) );
  AND2X2 AND2X2_1977 ( .A(u0_u0__abc_43300_n371), .B(u0_u0__abc_43300_n218_bF_buf2), .Y(u0_u0__abc_43300_n372) );
  AND2X2 AND2X2_1978 ( .A(u0_u0__abc_43300_n372), .B(u0_u0__abc_43300_n370), .Y(u0_u0_csc_5__FF_INPUT) );
  AND2X2 AND2X2_1979 ( .A(u0_u0__abc_43300_n375), .B(u0_u0__abc_43300_n218_bF_buf1), .Y(u0_u0__abc_43300_n376) );
  AND2X2 AND2X2_198 ( .A(spec_req_cs_2_bF_buf2), .B(u0_tms2_6_), .Y(u0__abc_49347_n1342) );
  AND2X2 AND2X2_1980 ( .A(u0_u0__abc_43300_n376), .B(u0_u0__abc_43300_n374), .Y(u0_u0_csc_6__FF_INPUT) );
  AND2X2 AND2X2_1981 ( .A(u0_u0__abc_43300_n379), .B(u0_u0__abc_43300_n218_bF_buf0), .Y(u0_u0__abc_43300_n380) );
  AND2X2 AND2X2_1982 ( .A(u0_u0__abc_43300_n380), .B(u0_u0__abc_43300_n378), .Y(u0_u0_csc_7__FF_INPUT) );
  AND2X2 AND2X2_1983 ( .A(u0_u0__abc_43300_n383), .B(u0_u0__abc_43300_n218_bF_buf7), .Y(u0_u0__abc_43300_n384) );
  AND2X2 AND2X2_1984 ( .A(u0_u0__abc_43300_n384), .B(u0_u0__abc_43300_n382), .Y(u0_u0_csc_8__FF_INPUT) );
  AND2X2 AND2X2_1985 ( .A(u0_u0__abc_43300_n387), .B(u0_u0__abc_43300_n218_bF_buf6), .Y(u0_u0__abc_43300_n388) );
  AND2X2 AND2X2_1986 ( .A(u0_u0__abc_43300_n388), .B(u0_u0__abc_43300_n386), .Y(u0_u0_csc_9__FF_INPUT) );
  AND2X2 AND2X2_1987 ( .A(u0_u0__abc_43300_n391), .B(u0_u0__abc_43300_n218_bF_buf5), .Y(u0_u0__abc_43300_n392) );
  AND2X2 AND2X2_1988 ( .A(u0_u0__abc_43300_n392), .B(u0_u0__abc_43300_n390), .Y(u0_u0_csc_10__FF_INPUT) );
  AND2X2 AND2X2_1989 ( .A(u0_u0__abc_43300_n395), .B(u0_u0__abc_43300_n218_bF_buf4), .Y(u0_u0__abc_43300_n396) );
  AND2X2 AND2X2_199 ( .A(u0__abc_49347_n1343), .B(u0__abc_49347_n1178_1_bF_buf5), .Y(u0__abc_49347_n1344_1) );
  AND2X2 AND2X2_1990 ( .A(u0_u0__abc_43300_n396), .B(u0_u0__abc_43300_n394), .Y(u0_u0_csc_11__FF_INPUT) );
  AND2X2 AND2X2_1991 ( .A(u0_u0__abc_43300_n399), .B(u0_u0__abc_43300_n218_bF_buf3), .Y(u0_u0__abc_43300_n400) );
  AND2X2 AND2X2_1992 ( .A(u0_u0__abc_43300_n400), .B(u0_u0__abc_43300_n398), .Y(u0_u0_csc_12__FF_INPUT) );
  AND2X2 AND2X2_1993 ( .A(u0_u0__abc_43300_n403), .B(u0_u0__abc_43300_n218_bF_buf2), .Y(u0_u0__abc_43300_n404) );
  AND2X2 AND2X2_1994 ( .A(u0_u0__abc_43300_n404), .B(u0_u0__abc_43300_n402), .Y(u0_u0_csc_13__FF_INPUT) );
  AND2X2 AND2X2_1995 ( .A(u0_u0__abc_43300_n407), .B(u0_u0__abc_43300_n218_bF_buf1), .Y(u0_u0__abc_43300_n408) );
  AND2X2 AND2X2_1996 ( .A(u0_u0__abc_43300_n408), .B(u0_u0__abc_43300_n406), .Y(u0_u0_csc_14__FF_INPUT) );
  AND2X2 AND2X2_1997 ( .A(u0_u0__abc_43300_n411), .B(u0_u0__abc_43300_n218_bF_buf0), .Y(u0_u0__abc_43300_n412) );
  AND2X2 AND2X2_1998 ( .A(u0_u0__abc_43300_n412), .B(u0_u0__abc_43300_n410), .Y(u0_u0_csc_15__FF_INPUT) );
  AND2X2 AND2X2_1999 ( .A(u0_u0__abc_43300_n415), .B(u0_u0__abc_43300_n218_bF_buf7), .Y(u0_u0__abc_43300_n416) );
  AND2X2 AND2X2_2 ( .A(_abc_55805_n241_1), .B(_abc_55805_n242_1), .Y(_abc_55805_n243) );
  AND2X2 AND2X2_20 ( .A(_abc_55805_n296), .B(_abc_55805_n297), .Y(tms_s_2_) );
  AND2X2 AND2X2_200 ( .A(spec_req_cs_1_bF_buf2), .B(u0_tms1_6_), .Y(u0__abc_49347_n1345_1) );
  AND2X2 AND2X2_2000 ( .A(u0_u0__abc_43300_n416), .B(u0_u0__abc_43300_n414), .Y(u0_u0_csc_16__FF_INPUT) );
  AND2X2 AND2X2_2001 ( .A(u0_u0__abc_43300_n419), .B(u0_u0__abc_43300_n218_bF_buf6), .Y(u0_u0__abc_43300_n420) );
  AND2X2 AND2X2_2002 ( .A(u0_u0__abc_43300_n420), .B(u0_u0__abc_43300_n418), .Y(u0_u0_csc_17__FF_INPUT) );
  AND2X2 AND2X2_2003 ( .A(u0_u0__abc_43300_n423), .B(u0_u0__abc_43300_n218_bF_buf5), .Y(u0_u0__abc_43300_n424) );
  AND2X2 AND2X2_2004 ( .A(u0_u0__abc_43300_n424), .B(u0_u0__abc_43300_n422), .Y(u0_u0_csc_18__FF_INPUT) );
  AND2X2 AND2X2_2005 ( .A(u0_u0__abc_43300_n427), .B(u0_u0__abc_43300_n218_bF_buf4), .Y(u0_u0__abc_43300_n428) );
  AND2X2 AND2X2_2006 ( .A(u0_u0__abc_43300_n428), .B(u0_u0__abc_43300_n426), .Y(u0_u0_csc_19__FF_INPUT) );
  AND2X2 AND2X2_2007 ( .A(u0_u0__abc_43300_n431), .B(u0_u0__abc_43300_n218_bF_buf3), .Y(u0_u0__abc_43300_n432) );
  AND2X2 AND2X2_2008 ( .A(u0_u0__abc_43300_n432), .B(u0_u0__abc_43300_n430), .Y(u0_u0_csc_20__FF_INPUT) );
  AND2X2 AND2X2_2009 ( .A(u0_u0__abc_43300_n435), .B(u0_u0__abc_43300_n218_bF_buf2), .Y(u0_u0__abc_43300_n436) );
  AND2X2 AND2X2_201 ( .A(u0__abc_49347_n1175_bF_buf6), .B(u0__abc_49347_n1348), .Y(u0__abc_49347_n1349) );
  AND2X2 AND2X2_2010 ( .A(u0_u0__abc_43300_n436), .B(u0_u0__abc_43300_n434), .Y(u0_u0_csc_21__FF_INPUT) );
  AND2X2 AND2X2_2011 ( .A(u0_u0__abc_43300_n439), .B(u0_u0__abc_43300_n218_bF_buf1), .Y(u0_u0__abc_43300_n440) );
  AND2X2 AND2X2_2012 ( .A(u0_u0__abc_43300_n440), .B(u0_u0__abc_43300_n438), .Y(u0_u0_csc_22__FF_INPUT) );
  AND2X2 AND2X2_2013 ( .A(u0_u0__abc_43300_n443), .B(u0_u0__abc_43300_n218_bF_buf0), .Y(u0_u0__abc_43300_n444) );
  AND2X2 AND2X2_2014 ( .A(u0_u0__abc_43300_n444), .B(u0_u0__abc_43300_n442), .Y(u0_u0_csc_23__FF_INPUT) );
  AND2X2 AND2X2_2015 ( .A(u0_u0__abc_43300_n447), .B(u0_u0__abc_43300_n218_bF_buf7), .Y(u0_u0__abc_43300_n448) );
  AND2X2 AND2X2_2016 ( .A(u0_u0__abc_43300_n448), .B(u0_u0__abc_43300_n446), .Y(u0_u0_csc_24__FF_INPUT) );
  AND2X2 AND2X2_2017 ( .A(u0_u0__abc_43300_n451), .B(u0_u0__abc_43300_n218_bF_buf6), .Y(u0_u0__abc_43300_n452) );
  AND2X2 AND2X2_2018 ( .A(u0_u0__abc_43300_n452), .B(u0_u0__abc_43300_n450), .Y(u0_u0_csc_25__FF_INPUT) );
  AND2X2 AND2X2_2019 ( .A(u0_u0__abc_43300_n455), .B(u0_u0__abc_43300_n218_bF_buf5), .Y(u0_u0__abc_43300_n456) );
  AND2X2 AND2X2_202 ( .A(u0__abc_49347_n1347), .B(u0__abc_49347_n1349), .Y(u0__abc_49347_n1350) );
  AND2X2 AND2X2_2020 ( .A(u0_u0__abc_43300_n456), .B(u0_u0__abc_43300_n454), .Y(u0_u0_csc_26__FF_INPUT) );
  AND2X2 AND2X2_2021 ( .A(u0_u0__abc_43300_n459), .B(u0_u0__abc_43300_n218_bF_buf4), .Y(u0_u0__abc_43300_n460) );
  AND2X2 AND2X2_2022 ( .A(u0_u0__abc_43300_n460), .B(u0_u0__abc_43300_n458), .Y(u0_u0_csc_27__FF_INPUT) );
  AND2X2 AND2X2_2023 ( .A(u0_u0__abc_43300_n463), .B(u0_u0__abc_43300_n218_bF_buf3), .Y(u0_u0__abc_43300_n464) );
  AND2X2 AND2X2_2024 ( .A(u0_u0__abc_43300_n464), .B(u0_u0__abc_43300_n462), .Y(u0_u0_csc_28__FF_INPUT) );
  AND2X2 AND2X2_2025 ( .A(u0_u0__abc_43300_n467), .B(u0_u0__abc_43300_n218_bF_buf2), .Y(u0_u0__abc_43300_n468) );
  AND2X2 AND2X2_2026 ( .A(u0_u0__abc_43300_n468), .B(u0_u0__abc_43300_n466), .Y(u0_u0_csc_29__FF_INPUT) );
  AND2X2 AND2X2_2027 ( .A(u0_u0__abc_43300_n471), .B(u0_u0__abc_43300_n218_bF_buf1), .Y(u0_u0__abc_43300_n472) );
  AND2X2 AND2X2_2028 ( .A(u0_u0__abc_43300_n472), .B(u0_u0__abc_43300_n470), .Y(u0_u0_csc_30__FF_INPUT) );
  AND2X2 AND2X2_2029 ( .A(u0_u0__abc_43300_n475), .B(u0_u0__abc_43300_n218_bF_buf0), .Y(u0_u0__abc_43300_n476) );
  AND2X2 AND2X2_203 ( .A(u0__abc_49347_n1176_1_bF_buf6), .B(sp_tms_7_), .Y(u0__abc_49347_n1352) );
  AND2X2 AND2X2_2030 ( .A(u0_u0__abc_43300_n476), .B(u0_u0__abc_43300_n474), .Y(u0_u0_csc_31__FF_INPUT) );
  AND2X2 AND2X2_2031 ( .A(u0_csc0_8_), .B(wb_we_i), .Y(u0_u0__abc_43300_n478) );
  AND2X2 AND2X2_2032 ( .A(u0_csc0_20_), .B(u0_csc_mask_4_), .Y(u0_u0__abc_43300_n479) );
  AND2X2 AND2X2_2033 ( .A(u0_csc_mask_4_), .B(wb_addr_i_25_bF_buf3), .Y(u0_u0__abc_43300_n480) );
  AND2X2 AND2X2_2034 ( .A(u0_csc_mask_3_), .B(\wb_addr_i[24] ), .Y(u0_u0__abc_43300_n483) );
  AND2X2 AND2X2_2035 ( .A(u0_csc0_19_), .B(u0_csc_mask_3_), .Y(u0_u0__abc_43300_n484) );
  AND2X2 AND2X2_2036 ( .A(u0_u0__abc_43300_n482), .B(u0_u0__abc_43300_n486), .Y(u0_u0__abc_43300_n487) );
  AND2X2 AND2X2_2037 ( .A(u0_csc0_18_), .B(u0_csc_mask_2_), .Y(u0_u0__abc_43300_n489) );
  AND2X2 AND2X2_2038 ( .A(u0_u0__abc_43300_n489), .B(u0_u0__abc_43300_n488), .Y(u0_u0__abc_43300_n490) );
  AND2X2 AND2X2_2039 ( .A(u0_u0__abc_43300_n493), .B(u0_u0__abc_43300_n491), .Y(u0_u0__abc_43300_n494) );
  AND2X2 AND2X2_204 ( .A(spec_req_cs_5_bF_buf1), .B(u0_tms5_7_), .Y(u0__abc_49347_n1353_1) );
  AND2X2 AND2X2_2040 ( .A(u0_u0__abc_43300_n487), .B(u0_u0__abc_43300_n494), .Y(u0_u0__abc_43300_n495) );
  AND2X2 AND2X2_2041 ( .A(u0_csc0_22_), .B(u0_csc_mask_6_), .Y(u0_u0__abc_43300_n496) );
  AND2X2 AND2X2_2042 ( .A(u0_csc_mask_6_), .B(\wb_addr_i[27] ), .Y(u0_u0__abc_43300_n497) );
  AND2X2 AND2X2_2043 ( .A(u0_csc_mask_5_), .B(\wb_addr_i[26] ), .Y(u0_u0__abc_43300_n500) );
  AND2X2 AND2X2_2044 ( .A(u0_csc0_21_), .B(u0_csc_mask_5_), .Y(u0_u0__abc_43300_n501) );
  AND2X2 AND2X2_2045 ( .A(u0_u0__abc_43300_n499), .B(u0_u0__abc_43300_n503), .Y(u0_u0__abc_43300_n504) );
  AND2X2 AND2X2_2046 ( .A(u0_u0__abc_43300_n479), .B(u0_u0__abc_43300_n505), .Y(u0_u0__abc_43300_n506) );
  AND2X2 AND2X2_2047 ( .A(u0_u0__abc_43300_n509), .B(u0_u0__abc_43300_n507), .Y(u0_u0__abc_43300_n510) );
  AND2X2 AND2X2_2048 ( .A(u0_u0__abc_43300_n504), .B(u0_u0__abc_43300_n510), .Y(u0_u0__abc_43300_n511) );
  AND2X2 AND2X2_2049 ( .A(u0_u0__abc_43300_n495), .B(u0_u0__abc_43300_n511), .Y(u0_u0__abc_43300_n512) );
  AND2X2 AND2X2_205 ( .A(u0__abc_49347_n1355), .B(u0__abc_49347_n1185_bF_buf4), .Y(u0__abc_49347_n1356) );
  AND2X2 AND2X2_2050 ( .A(u0_u0__abc_43300_n498), .B(u0_u0__abc_43300_n496), .Y(u0_u0__abc_43300_n513) );
  AND2X2 AND2X2_2051 ( .A(u0_csc_mask_7_), .B(\wb_addr_i[28] ), .Y(u0_u0__abc_43300_n515) );
  AND2X2 AND2X2_2052 ( .A(u0_csc0_23_), .B(u0_csc_mask_7_), .Y(u0_u0__abc_43300_n517) );
  AND2X2 AND2X2_2053 ( .A(u0_u0__abc_43300_n514), .B(u0_u0__abc_43300_n518), .Y(u0_u0__abc_43300_n519) );
  AND2X2 AND2X2_2054 ( .A(u0_u0__abc_43300_n519), .B(u0_u0__abc_43300_n521), .Y(u0_u0__abc_43300_n522) );
  AND2X2 AND2X2_2055 ( .A(u0_u0__abc_43300_n512), .B(u0_u0__abc_43300_n522), .Y(u0_u0__abc_43300_n523) );
  AND2X2 AND2X2_2056 ( .A(u0_csc_mask_2_), .B(wb_addr_i_23_bF_buf2), .Y(u0_u0__abc_43300_n524) );
  AND2X2 AND2X2_2057 ( .A(u0_csc_mask_1_), .B(\wb_addr_i[22] ), .Y(u0_u0__abc_43300_n527) );
  AND2X2 AND2X2_2058 ( .A(u0_csc0_17_), .B(u0_csc_mask_1_), .Y(u0_u0__abc_43300_n528) );
  AND2X2 AND2X2_2059 ( .A(u0_u0__abc_43300_n526), .B(u0_u0__abc_43300_n530), .Y(u0_u0__abc_43300_n531) );
  AND2X2 AND2X2_206 ( .A(u0__abc_49347_n1356), .B(u0__abc_49347_n1354_1), .Y(u0__abc_49347_n1357) );
  AND2X2 AND2X2_2060 ( .A(u0_csc_mask_0_), .B(\wb_addr_i[21] ), .Y(u0_u0__abc_43300_n532) );
  AND2X2 AND2X2_2061 ( .A(u0_csc0_16_), .B(u0_csc_mask_0_), .Y(u0_u0__abc_43300_n533) );
  AND2X2 AND2X2_2062 ( .A(u0_u0__abc_43300_n535), .B(u0_u0__abc_43300_n537), .Y(u0_u0__abc_43300_n538) );
  AND2X2 AND2X2_2063 ( .A(u0_u0__abc_43300_n531), .B(u0_u0__abc_43300_n538), .Y(u0_u0__abc_43300_n539) );
  AND2X2 AND2X2_2064 ( .A(u0_u0__abc_43300_n541), .B(u0_csc0_0_), .Y(u0_u0__abc_43300_n542) );
  AND2X2 AND2X2_2065 ( .A(u0_u0__abc_43300_n539), .B(u0_u0__abc_43300_n542), .Y(u0_u0__abc_43300_n543) );
  AND2X2 AND2X2_2066 ( .A(u0_u0__abc_43300_n523), .B(u0_u0__abc_43300_n543), .Y(u0_u0__abc_43300_n544) );
  AND2X2 AND2X2_2067 ( .A(u0_u0__abc_43300_n544), .B(u0_u0__abc_43300_n478), .Y(u0_u0_wp_err) );
  AND2X2 AND2X2_2068 ( .A(u0_u0__abc_43300_n544), .B(u0_u0__abc_43300_n546), .Y(u0_cs0) );
  AND2X2 AND2X2_2069 ( .A(u0_u0__abc_43300_n549), .B(u0_init_req0), .Y(u0_u0__abc_43300_n550) );
  AND2X2 AND2X2_207 ( .A(u0__abc_49347_n1358), .B(u0__abc_49347_n1181_bF_buf4), .Y(u0__abc_49347_n1359) );
  AND2X2 AND2X2_2070 ( .A(u0_u0__abc_43300_n551), .B(u0_csc0_0_), .Y(u0_u0__abc_43300_n552) );
  AND2X2 AND2X2_2071 ( .A(u0_u0__abc_43300_n552), .B(u0_u0_init_req_we), .Y(u0_u0__abc_43300_n553) );
  AND2X2 AND2X2_2072 ( .A(u0_u0__abc_43300_n203), .B(u0_u0__abc_43300_n553), .Y(u0_u0__abc_43300_n554) );
  AND2X2 AND2X2_2073 ( .A(u0_u1__abc_43657_n203_1), .B(u0_u1_lmr_req_we), .Y(u0_u1__abc_43657_n204_1) );
  AND2X2 AND2X2_2074 ( .A(u0_u1__abc_43657_n204_1), .B(u0_u1_inited), .Y(u0_u1__abc_43657_n205) );
  AND2X2 AND2X2_2075 ( .A(u0_u1__abc_43657_n207_1), .B(u0_lmr_req1), .Y(u0_u1__abc_43657_n208) );
  AND2X2 AND2X2_2076 ( .A(u0_u1__abc_43657_n206_1), .B(u0_u1__abc_43657_n208), .Y(u0_u1__abc_43657_n209_1) );
  AND2X2 AND2X2_2077 ( .A(u0_u1__abc_43657_n211), .B(u0_u1__abc_43657_n212_1), .Y(u0_u1__abc_43657_n213_1) );
  AND2X2 AND2X2_2078 ( .A(u0_u1_addr_r_4_), .B(u0_u1_addr_r_3_), .Y(u0_u1__abc_43657_n214) );
  AND2X2 AND2X2_2079 ( .A(u0_u1__abc_43657_n214), .B(u0_rf_we), .Y(u0_u1__abc_43657_n215_1) );
  AND2X2 AND2X2_208 ( .A(spec_req_cs_4_bF_buf1), .B(u0_tms4_7_), .Y(u0__abc_49347_n1360) );
  AND2X2 AND2X2_2080 ( .A(u0_u1__abc_43657_n215_1), .B(u0_u1__abc_43657_n213_1), .Y(u0_u1__abc_43657_n216_1) );
  AND2X2 AND2X2_2081 ( .A(u0_u1__abc_43657_n216_1), .B(u0_u1_addr_r_2_), .Y(u0_u1_lmr_req_we_FF_INPUT) );
  AND2X2 AND2X2_2082 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf6), .B(u0_u1__abc_43657_n220), .Y(u0_u1__abc_43657_n221_1) );
  AND2X2 AND2X2_2083 ( .A(u0_u1__abc_43657_n222_1), .B(u0_u1__abc_43657_n219_1_bF_buf7), .Y(u0_u1__abc_43657_n223) );
  AND2X2 AND2X2_2084 ( .A(u0_u1__abc_43657_n223), .B(u0_u1__abc_43657_n218_1), .Y(u0_u1_tms_0__FF_INPUT) );
  AND2X2 AND2X2_2085 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf4), .B(u0_u1__abc_43657_n226), .Y(u0_u1__abc_43657_n227_1) );
  AND2X2 AND2X2_2086 ( .A(u0_u1__abc_43657_n228_1), .B(u0_u1__abc_43657_n219_1_bF_buf6), .Y(u0_u1__abc_43657_n229) );
  AND2X2 AND2X2_2087 ( .A(u0_u1__abc_43657_n229), .B(u0_u1__abc_43657_n225_1), .Y(u0_u1_tms_1__FF_INPUT) );
  AND2X2 AND2X2_2088 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf2), .B(u0_u1__abc_43657_n232), .Y(u0_u1__abc_43657_n233_1) );
  AND2X2 AND2X2_2089 ( .A(u0_u1__abc_43657_n234_1), .B(u0_u1__abc_43657_n219_1_bF_buf5), .Y(u0_u1__abc_43657_n235) );
  AND2X2 AND2X2_209 ( .A(u0__abc_49347_n1361), .B(u0__abc_49347_n1180_1_bF_buf4), .Y(u0__abc_49347_n1362_1) );
  AND2X2 AND2X2_2090 ( .A(u0_u1__abc_43657_n235), .B(u0_u1__abc_43657_n231_1), .Y(u0_u1_tms_2__FF_INPUT) );
  AND2X2 AND2X2_2091 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf0), .B(u0_u1__abc_43657_n238), .Y(u0_u1__abc_43657_n239_1) );
  AND2X2 AND2X2_2092 ( .A(u0_u1__abc_43657_n240_1), .B(u0_u1__abc_43657_n219_1_bF_buf4), .Y(u0_u1__abc_43657_n241) );
  AND2X2 AND2X2_2093 ( .A(u0_u1__abc_43657_n241), .B(u0_u1__abc_43657_n237_1), .Y(u0_u1_tms_3__FF_INPUT) );
  AND2X2 AND2X2_2094 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf6), .B(u0_u1__abc_43657_n244), .Y(u0_u1__abc_43657_n245_1) );
  AND2X2 AND2X2_2095 ( .A(u0_u1__abc_43657_n246_1), .B(u0_u1__abc_43657_n219_1_bF_buf3), .Y(u0_u1__abc_43657_n247) );
  AND2X2 AND2X2_2096 ( .A(u0_u1__abc_43657_n247), .B(u0_u1__abc_43657_n243_1), .Y(u0_u1_tms_4__FF_INPUT) );
  AND2X2 AND2X2_2097 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf4), .B(u0_u1__abc_43657_n250), .Y(u0_u1__abc_43657_n251_1) );
  AND2X2 AND2X2_2098 ( .A(u0_u1__abc_43657_n252_1), .B(u0_u1__abc_43657_n219_1_bF_buf2), .Y(u0_u1__abc_43657_n253) );
  AND2X2 AND2X2_2099 ( .A(u0_u1__abc_43657_n253), .B(u0_u1__abc_43657_n249_1), .Y(u0_u1_tms_5__FF_INPUT) );
  AND2X2 AND2X2_21 ( .A(_abc_55805_n299), .B(_abc_55805_n300), .Y(tms_s_3_) );
  AND2X2 AND2X2_210 ( .A(spec_req_cs_3_bF_buf1), .B(u0_tms3_7_), .Y(u0__abc_49347_n1363_1) );
  AND2X2 AND2X2_2100 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf2), .B(u0_u1__abc_43657_n256), .Y(u0_u1__abc_43657_n257) );
  AND2X2 AND2X2_2101 ( .A(u0_u1__abc_43657_n258), .B(u0_u1__abc_43657_n219_1_bF_buf1), .Y(u0_u1__abc_43657_n259_1) );
  AND2X2 AND2X2_2102 ( .A(u0_u1__abc_43657_n259_1), .B(u0_u1__abc_43657_n255), .Y(u0_u1_tms_6__FF_INPUT) );
  AND2X2 AND2X2_2103 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf0), .B(u0_u1__abc_43657_n262), .Y(u0_u1__abc_43657_n263) );
  AND2X2 AND2X2_2104 ( .A(u0_u1__abc_43657_n264), .B(u0_u1__abc_43657_n219_1_bF_buf0), .Y(u0_u1__abc_43657_n265_1) );
  AND2X2 AND2X2_2105 ( .A(u0_u1__abc_43657_n265_1), .B(u0_u1__abc_43657_n261_1), .Y(u0_u1_tms_7__FF_INPUT) );
  AND2X2 AND2X2_2106 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf6), .B(u0_u1__abc_43657_n268), .Y(u0_u1__abc_43657_n269) );
  AND2X2 AND2X2_2107 ( .A(u0_u1__abc_43657_n270), .B(u0_u1__abc_43657_n219_1_bF_buf7), .Y(u0_u1__abc_43657_n271) );
  AND2X2 AND2X2_2108 ( .A(u0_u1__abc_43657_n271), .B(u0_u1__abc_43657_n267_1), .Y(u0_u1_tms_8__FF_INPUT) );
  AND2X2 AND2X2_2109 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf4), .B(u0_u1__abc_43657_n274_1), .Y(u0_u1__abc_43657_n275) );
  AND2X2 AND2X2_211 ( .A(u0__abc_49347_n1364), .B(u0__abc_49347_n1179_bF_buf4), .Y(u0__abc_49347_n1365) );
  AND2X2 AND2X2_2110 ( .A(u0_u1__abc_43657_n276_1), .B(u0_u1__abc_43657_n219_1_bF_buf6), .Y(u0_u1__abc_43657_n277) );
  AND2X2 AND2X2_2111 ( .A(u0_u1__abc_43657_n277), .B(u0_u1__abc_43657_n273), .Y(u0_u1_tms_9__FF_INPUT) );
  AND2X2 AND2X2_2112 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf2), .B(u0_u1__abc_43657_n280), .Y(u0_u1__abc_43657_n281) );
  AND2X2 AND2X2_2113 ( .A(u0_u1__abc_43657_n282_1), .B(u0_u1__abc_43657_n219_1_bF_buf5), .Y(u0_u1__abc_43657_n283) );
  AND2X2 AND2X2_2114 ( .A(u0_u1__abc_43657_n283), .B(u0_u1__abc_43657_n279), .Y(u0_u1_tms_10__FF_INPUT) );
  AND2X2 AND2X2_2115 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf0), .B(u0_u1__abc_43657_n286_1), .Y(u0_u1__abc_43657_n287) );
  AND2X2 AND2X2_2116 ( .A(u0_u1__abc_43657_n288_1), .B(u0_u1__abc_43657_n219_1_bF_buf4), .Y(u0_u1__abc_43657_n289) );
  AND2X2 AND2X2_2117 ( .A(u0_u1__abc_43657_n289), .B(u0_u1__abc_43657_n285), .Y(u0_u1_tms_11__FF_INPUT) );
  AND2X2 AND2X2_2118 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf6), .B(u0_u1__abc_43657_n292), .Y(u0_u1__abc_43657_n293) );
  AND2X2 AND2X2_2119 ( .A(u0_u1__abc_43657_n294), .B(u0_u1__abc_43657_n219_1_bF_buf3), .Y(u0_u1__abc_43657_n295_1) );
  AND2X2 AND2X2_212 ( .A(spec_req_cs_2_bF_buf1), .B(u0_tms2_7_), .Y(u0__abc_49347_n1366) );
  AND2X2 AND2X2_2120 ( .A(u0_u1__abc_43657_n295_1), .B(u0_u1__abc_43657_n291), .Y(u0_u1_tms_12__FF_INPUT) );
  AND2X2 AND2X2_2121 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf4), .B(u0_u1__abc_43657_n298), .Y(u0_u1__abc_43657_n299) );
  AND2X2 AND2X2_2122 ( .A(u0_u1__abc_43657_n300), .B(u0_u1__abc_43657_n219_1_bF_buf2), .Y(u0_u1__abc_43657_n301) );
  AND2X2 AND2X2_2123 ( .A(u0_u1__abc_43657_n301), .B(u0_u1__abc_43657_n297_1), .Y(u0_u1_tms_13__FF_INPUT) );
  AND2X2 AND2X2_2124 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf2), .B(u0_u1__abc_43657_n304), .Y(u0_u1__abc_43657_n305) );
  AND2X2 AND2X2_2125 ( .A(u0_u1__abc_43657_n306), .B(u0_u1__abc_43657_n219_1_bF_buf1), .Y(u0_u1__abc_43657_n307) );
  AND2X2 AND2X2_2126 ( .A(u0_u1__abc_43657_n307), .B(u0_u1__abc_43657_n303), .Y(u0_u1_tms_14__FF_INPUT) );
  AND2X2 AND2X2_2127 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf0), .B(u0_u1__abc_43657_n310), .Y(u0_u1__abc_43657_n311_1) );
  AND2X2 AND2X2_2128 ( .A(u0_u1__abc_43657_n312), .B(u0_u1__abc_43657_n219_1_bF_buf0), .Y(u0_u1__abc_43657_n313_1) );
  AND2X2 AND2X2_2129 ( .A(u0_u1__abc_43657_n313_1), .B(u0_u1__abc_43657_n309_1), .Y(u0_u1_tms_15__FF_INPUT) );
  AND2X2 AND2X2_213 ( .A(u0__abc_49347_n1367), .B(u0__abc_49347_n1178_1_bF_buf4), .Y(u0__abc_49347_n1368) );
  AND2X2 AND2X2_2130 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf6), .B(u0_u1__abc_43657_n316_1), .Y(u0_u1__abc_43657_n317) );
  AND2X2 AND2X2_2131 ( .A(u0_u1__abc_43657_n318), .B(u0_u1__abc_43657_n219_1_bF_buf7), .Y(u0_u1__abc_43657_n319) );
  AND2X2 AND2X2_2132 ( .A(u0_u1__abc_43657_n319), .B(u0_u1__abc_43657_n315_1), .Y(u0_u1_tms_16__FF_INPUT) );
  AND2X2 AND2X2_2133 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf4), .B(u0_u1__abc_43657_n322_1), .Y(u0_u1__abc_43657_n323_1) );
  AND2X2 AND2X2_2134 ( .A(u0_u1__abc_43657_n324_1), .B(u0_u1__abc_43657_n219_1_bF_buf6), .Y(u0_u1__abc_43657_n325) );
  AND2X2 AND2X2_2135 ( .A(u0_u1__abc_43657_n325), .B(u0_u1__abc_43657_n321), .Y(u0_u1_tms_17__FF_INPUT) );
  AND2X2 AND2X2_2136 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf2), .B(u0_u1__abc_43657_n328), .Y(u0_u1__abc_43657_n329) );
  AND2X2 AND2X2_2137 ( .A(u0_u1__abc_43657_n330), .B(u0_u1__abc_43657_n219_1_bF_buf5), .Y(u0_u1__abc_43657_n331) );
  AND2X2 AND2X2_2138 ( .A(u0_u1__abc_43657_n331), .B(u0_u1__abc_43657_n327), .Y(u0_u1_tms_18__FF_INPUT) );
  AND2X2 AND2X2_2139 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf0), .B(u0_u1__abc_43657_n334), .Y(u0_u1__abc_43657_n335) );
  AND2X2 AND2X2_214 ( .A(spec_req_cs_1_bF_buf1), .B(u0_tms1_7_), .Y(u0__abc_49347_n1369) );
  AND2X2 AND2X2_2140 ( .A(u0_u1__abc_43657_n336), .B(u0_u1__abc_43657_n219_1_bF_buf4), .Y(u0_u1__abc_43657_n337) );
  AND2X2 AND2X2_2141 ( .A(u0_u1__abc_43657_n337), .B(u0_u1__abc_43657_n333), .Y(u0_u1_tms_19__FF_INPUT) );
  AND2X2 AND2X2_2142 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf6), .B(u0_u1__abc_43657_n340), .Y(u0_u1__abc_43657_n341) );
  AND2X2 AND2X2_2143 ( .A(u0_u1__abc_43657_n342), .B(u0_u1__abc_43657_n219_1_bF_buf3), .Y(u0_u1__abc_43657_n343) );
  AND2X2 AND2X2_2144 ( .A(u0_u1__abc_43657_n343), .B(u0_u1__abc_43657_n339), .Y(u0_u1_tms_20__FF_INPUT) );
  AND2X2 AND2X2_2145 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf4), .B(u0_u1__abc_43657_n346), .Y(u0_u1__abc_43657_n347) );
  AND2X2 AND2X2_2146 ( .A(u0_u1__abc_43657_n348), .B(u0_u1__abc_43657_n219_1_bF_buf2), .Y(u0_u1__abc_43657_n349) );
  AND2X2 AND2X2_2147 ( .A(u0_u1__abc_43657_n349), .B(u0_u1__abc_43657_n345), .Y(u0_u1_tms_21__FF_INPUT) );
  AND2X2 AND2X2_2148 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf2), .B(u0_u1__abc_43657_n352), .Y(u0_u1__abc_43657_n353) );
  AND2X2 AND2X2_2149 ( .A(u0_u1__abc_43657_n354), .B(u0_u1__abc_43657_n219_1_bF_buf1), .Y(u0_u1__abc_43657_n355) );
  AND2X2 AND2X2_215 ( .A(u0__abc_49347_n1175_bF_buf5), .B(u0__abc_49347_n1372_1), .Y(u0__abc_49347_n1373) );
  AND2X2 AND2X2_2150 ( .A(u0_u1__abc_43657_n355), .B(u0_u1__abc_43657_n351), .Y(u0_u1_tms_22__FF_INPUT) );
  AND2X2 AND2X2_2151 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf0), .B(u0_u1__abc_43657_n358), .Y(u0_u1__abc_43657_n359) );
  AND2X2 AND2X2_2152 ( .A(u0_u1__abc_43657_n360), .B(u0_u1__abc_43657_n219_1_bF_buf0), .Y(u0_u1__abc_43657_n361) );
  AND2X2 AND2X2_2153 ( .A(u0_u1__abc_43657_n361), .B(u0_u1__abc_43657_n357), .Y(u0_u1_tms_23__FF_INPUT) );
  AND2X2 AND2X2_2154 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf6), .B(u0_u1__abc_43657_n364), .Y(u0_u1__abc_43657_n365) );
  AND2X2 AND2X2_2155 ( .A(u0_u1__abc_43657_n366), .B(u0_u1__abc_43657_n219_1_bF_buf7), .Y(u0_u1__abc_43657_n367) );
  AND2X2 AND2X2_2156 ( .A(u0_u1__abc_43657_n367), .B(u0_u1__abc_43657_n363), .Y(u0_u1_tms_24__FF_INPUT) );
  AND2X2 AND2X2_2157 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf4), .B(u0_u1__abc_43657_n370), .Y(u0_u1__abc_43657_n371) );
  AND2X2 AND2X2_2158 ( .A(u0_u1__abc_43657_n372), .B(u0_u1__abc_43657_n219_1_bF_buf6), .Y(u0_u1__abc_43657_n373) );
  AND2X2 AND2X2_2159 ( .A(u0_u1__abc_43657_n373), .B(u0_u1__abc_43657_n369), .Y(u0_u1_tms_25__FF_INPUT) );
  AND2X2 AND2X2_216 ( .A(u0__abc_49347_n1371_1), .B(u0__abc_49347_n1373), .Y(u0__abc_49347_n1374) );
  AND2X2 AND2X2_2160 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf2), .B(u0_u1__abc_43657_n376), .Y(u0_u1__abc_43657_n377) );
  AND2X2 AND2X2_2161 ( .A(u0_u1__abc_43657_n378), .B(u0_u1__abc_43657_n219_1_bF_buf5), .Y(u0_u1__abc_43657_n379) );
  AND2X2 AND2X2_2162 ( .A(u0_u1__abc_43657_n379), .B(u0_u1__abc_43657_n375), .Y(u0_u1_tms_26__FF_INPUT) );
  AND2X2 AND2X2_2163 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf0), .B(u0_u1__abc_43657_n382), .Y(u0_u1__abc_43657_n383) );
  AND2X2 AND2X2_2164 ( .A(u0_u1__abc_43657_n384), .B(u0_u1__abc_43657_n219_1_bF_buf4), .Y(u0_u1__abc_43657_n385) );
  AND2X2 AND2X2_2165 ( .A(u0_u1__abc_43657_n385), .B(u0_u1__abc_43657_n381), .Y(u0_u1_tms_27__FF_INPUT) );
  AND2X2 AND2X2_2166 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf6), .B(u0_u1__abc_43657_n388), .Y(u0_u1__abc_43657_n389) );
  AND2X2 AND2X2_2167 ( .A(u0_u1__abc_43657_n390), .B(u0_u1__abc_43657_n219_1_bF_buf3), .Y(u0_u1__abc_43657_n391) );
  AND2X2 AND2X2_2168 ( .A(u0_u1__abc_43657_n391), .B(u0_u1__abc_43657_n387), .Y(u0_u1_tms_28__FF_INPUT) );
  AND2X2 AND2X2_2169 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf4), .B(u0_u1__abc_43657_n394), .Y(u0_u1__abc_43657_n395) );
  AND2X2 AND2X2_217 ( .A(u0__abc_49347_n1176_1_bF_buf5), .B(sp_tms_8_), .Y(u0__abc_49347_n1376) );
  AND2X2 AND2X2_2170 ( .A(u0_u1__abc_43657_n396), .B(u0_u1__abc_43657_n219_1_bF_buf2), .Y(u0_u1__abc_43657_n397) );
  AND2X2 AND2X2_2171 ( .A(u0_u1__abc_43657_n397), .B(u0_u1__abc_43657_n393), .Y(u0_u1_tms_29__FF_INPUT) );
  AND2X2 AND2X2_2172 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf2), .B(u0_u1__abc_43657_n400), .Y(u0_u1__abc_43657_n401) );
  AND2X2 AND2X2_2173 ( .A(u0_u1__abc_43657_n402), .B(u0_u1__abc_43657_n219_1_bF_buf1), .Y(u0_u1__abc_43657_n403) );
  AND2X2 AND2X2_2174 ( .A(u0_u1__abc_43657_n403), .B(u0_u1__abc_43657_n399), .Y(u0_u1_tms_30__FF_INPUT) );
  AND2X2 AND2X2_2175 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf0), .B(u0_u1__abc_43657_n406), .Y(u0_u1__abc_43657_n407) );
  AND2X2 AND2X2_2176 ( .A(u0_u1__abc_43657_n408), .B(u0_u1__abc_43657_n219_1_bF_buf0), .Y(u0_u1__abc_43657_n409) );
  AND2X2 AND2X2_2177 ( .A(u0_u1__abc_43657_n409), .B(u0_u1__abc_43657_n405), .Y(u0_u1_tms_31__FF_INPUT) );
  AND2X2 AND2X2_2178 ( .A(u0_u1__abc_43657_n216_1), .B(u0_u1__abc_43657_n411), .Y(u0_u1_init_req_we_FF_INPUT) );
  AND2X2 AND2X2_2179 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf6), .B(u0_u1__abc_43657_n220), .Y(u0_u1__abc_43657_n414) );
  AND2X2 AND2X2_218 ( .A(spec_req_cs_5_bF_buf0), .B(u0_tms5_8_), .Y(u0__abc_49347_n1377) );
  AND2X2 AND2X2_2180 ( .A(u0_u1__abc_43657_n415), .B(u0_u1__abc_43657_n219_1_bF_buf7), .Y(u0_u1__abc_43657_n416) );
  AND2X2 AND2X2_2181 ( .A(u0_u1__abc_43657_n416), .B(u0_u1__abc_43657_n413), .Y(u0_u1_csc_0__FF_INPUT) );
  AND2X2 AND2X2_2182 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf4), .B(u0_u1__abc_43657_n226), .Y(u0_u1__abc_43657_n419) );
  AND2X2 AND2X2_2183 ( .A(u0_u1__abc_43657_n420), .B(u0_u1__abc_43657_n219_1_bF_buf6), .Y(u0_u1__abc_43657_n421) );
  AND2X2 AND2X2_2184 ( .A(u0_u1__abc_43657_n421), .B(u0_u1__abc_43657_n418), .Y(u0_u1_csc_1__FF_INPUT) );
  AND2X2 AND2X2_2185 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf2), .B(u0_u1__abc_43657_n232), .Y(u0_u1__abc_43657_n424) );
  AND2X2 AND2X2_2186 ( .A(u0_u1__abc_43657_n425), .B(u0_u1__abc_43657_n219_1_bF_buf5), .Y(u0_u1__abc_43657_n426) );
  AND2X2 AND2X2_2187 ( .A(u0_u1__abc_43657_n426), .B(u0_u1__abc_43657_n423), .Y(u0_u1_csc_2__FF_INPUT) );
  AND2X2 AND2X2_2188 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf0), .B(u0_u1__abc_43657_n238), .Y(u0_u1__abc_43657_n429) );
  AND2X2 AND2X2_2189 ( .A(u0_u1__abc_43657_n430), .B(u0_u1__abc_43657_n219_1_bF_buf4), .Y(u0_u1__abc_43657_n431) );
  AND2X2 AND2X2_219 ( .A(u0__abc_49347_n1379), .B(u0__abc_49347_n1185_bF_buf3), .Y(u0__abc_49347_n1380_1) );
  AND2X2 AND2X2_2190 ( .A(u0_u1__abc_43657_n431), .B(u0_u1__abc_43657_n428), .Y(u0_u1_csc_3__FF_INPUT) );
  AND2X2 AND2X2_2191 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf6), .B(u0_u1__abc_43657_n244), .Y(u0_u1__abc_43657_n434) );
  AND2X2 AND2X2_2192 ( .A(u0_u1__abc_43657_n435), .B(u0_u1__abc_43657_n219_1_bF_buf3), .Y(u0_u1__abc_43657_n436) );
  AND2X2 AND2X2_2193 ( .A(u0_u1__abc_43657_n436), .B(u0_u1__abc_43657_n433), .Y(u0_u1_csc_4__FF_INPUT) );
  AND2X2 AND2X2_2194 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf4), .B(u0_u1__abc_43657_n250), .Y(u0_u1__abc_43657_n439) );
  AND2X2 AND2X2_2195 ( .A(u0_u1__abc_43657_n440), .B(u0_u1__abc_43657_n219_1_bF_buf2), .Y(u0_u1__abc_43657_n441) );
  AND2X2 AND2X2_2196 ( .A(u0_u1__abc_43657_n441), .B(u0_u1__abc_43657_n438), .Y(u0_u1_csc_5__FF_INPUT) );
  AND2X2 AND2X2_2197 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf2), .B(u0_u1__abc_43657_n256), .Y(u0_u1__abc_43657_n444) );
  AND2X2 AND2X2_2198 ( .A(u0_u1__abc_43657_n445), .B(u0_u1__abc_43657_n219_1_bF_buf1), .Y(u0_u1__abc_43657_n446) );
  AND2X2 AND2X2_2199 ( .A(u0_u1__abc_43657_n446), .B(u0_u1__abc_43657_n443), .Y(u0_u1_csc_6__FF_INPUT) );
  AND2X2 AND2X2_22 ( .A(_abc_55805_n302), .B(_abc_55805_n303), .Y(tms_s_4_) );
  AND2X2 AND2X2_220 ( .A(u0__abc_49347_n1380_1), .B(u0__abc_49347_n1378), .Y(u0__abc_49347_n1381_1) );
  AND2X2 AND2X2_2200 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf0), .B(u0_u1__abc_43657_n262), .Y(u0_u1__abc_43657_n449) );
  AND2X2 AND2X2_2201 ( .A(u0_u1__abc_43657_n450), .B(u0_u1__abc_43657_n219_1_bF_buf0), .Y(u0_u1__abc_43657_n451) );
  AND2X2 AND2X2_2202 ( .A(u0_u1__abc_43657_n451), .B(u0_u1__abc_43657_n448), .Y(u0_u1_csc_7__FF_INPUT) );
  AND2X2 AND2X2_2203 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf6), .B(u0_u1__abc_43657_n268), .Y(u0_u1__abc_43657_n454) );
  AND2X2 AND2X2_2204 ( .A(u0_u1__abc_43657_n455), .B(u0_u1__abc_43657_n219_1_bF_buf7), .Y(u0_u1__abc_43657_n456) );
  AND2X2 AND2X2_2205 ( .A(u0_u1__abc_43657_n456), .B(u0_u1__abc_43657_n453), .Y(u0_u1_csc_8__FF_INPUT) );
  AND2X2 AND2X2_2206 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf4), .B(u0_u1__abc_43657_n274_1), .Y(u0_u1__abc_43657_n459) );
  AND2X2 AND2X2_2207 ( .A(u0_u1__abc_43657_n460), .B(u0_u1__abc_43657_n219_1_bF_buf6), .Y(u0_u1__abc_43657_n461) );
  AND2X2 AND2X2_2208 ( .A(u0_u1__abc_43657_n461), .B(u0_u1__abc_43657_n458), .Y(u0_u1_csc_9__FF_INPUT) );
  AND2X2 AND2X2_2209 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf2), .B(u0_u1__abc_43657_n280), .Y(u0_u1__abc_43657_n464) );
  AND2X2 AND2X2_221 ( .A(u0__abc_49347_n1382), .B(u0__abc_49347_n1181_bF_buf3), .Y(u0__abc_49347_n1383) );
  AND2X2 AND2X2_2210 ( .A(u0_u1__abc_43657_n465), .B(u0_u1__abc_43657_n219_1_bF_buf5), .Y(u0_u1__abc_43657_n466) );
  AND2X2 AND2X2_2211 ( .A(u0_u1__abc_43657_n466), .B(u0_u1__abc_43657_n463), .Y(u0_u1_csc_10__FF_INPUT) );
  AND2X2 AND2X2_2212 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf0), .B(u0_u1__abc_43657_n286_1), .Y(u0_u1__abc_43657_n469) );
  AND2X2 AND2X2_2213 ( .A(u0_u1__abc_43657_n470), .B(u0_u1__abc_43657_n219_1_bF_buf4), .Y(u0_u1__abc_43657_n471) );
  AND2X2 AND2X2_2214 ( .A(u0_u1__abc_43657_n471), .B(u0_u1__abc_43657_n468), .Y(u0_u1_csc_11__FF_INPUT) );
  AND2X2 AND2X2_2215 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf6), .B(u0_u1__abc_43657_n292), .Y(u0_u1__abc_43657_n474) );
  AND2X2 AND2X2_2216 ( .A(u0_u1__abc_43657_n475), .B(u0_u1__abc_43657_n219_1_bF_buf3), .Y(u0_u1__abc_43657_n476) );
  AND2X2 AND2X2_2217 ( .A(u0_u1__abc_43657_n476), .B(u0_u1__abc_43657_n473), .Y(u0_u1_csc_12__FF_INPUT) );
  AND2X2 AND2X2_2218 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf4), .B(u0_u1__abc_43657_n298), .Y(u0_u1__abc_43657_n479) );
  AND2X2 AND2X2_2219 ( .A(u0_u1__abc_43657_n480), .B(u0_u1__abc_43657_n219_1_bF_buf2), .Y(u0_u1__abc_43657_n481) );
  AND2X2 AND2X2_222 ( .A(spec_req_cs_4_bF_buf0), .B(u0_tms4_8_), .Y(u0__abc_49347_n1384) );
  AND2X2 AND2X2_2220 ( .A(u0_u1__abc_43657_n481), .B(u0_u1__abc_43657_n478), .Y(u0_u1_csc_13__FF_INPUT) );
  AND2X2 AND2X2_2221 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf2), .B(u0_u1__abc_43657_n304), .Y(u0_u1__abc_43657_n484) );
  AND2X2 AND2X2_2222 ( .A(u0_u1__abc_43657_n485), .B(u0_u1__abc_43657_n219_1_bF_buf1), .Y(u0_u1__abc_43657_n486) );
  AND2X2 AND2X2_2223 ( .A(u0_u1__abc_43657_n486), .B(u0_u1__abc_43657_n483), .Y(u0_u1_csc_14__FF_INPUT) );
  AND2X2 AND2X2_2224 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf0), .B(u0_u1__abc_43657_n310), .Y(u0_u1__abc_43657_n489) );
  AND2X2 AND2X2_2225 ( .A(u0_u1__abc_43657_n490), .B(u0_u1__abc_43657_n219_1_bF_buf0), .Y(u0_u1__abc_43657_n491) );
  AND2X2 AND2X2_2226 ( .A(u0_u1__abc_43657_n491), .B(u0_u1__abc_43657_n488), .Y(u0_u1_csc_15__FF_INPUT) );
  AND2X2 AND2X2_2227 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf6), .B(u0_u1__abc_43657_n316_1), .Y(u0_u1__abc_43657_n494) );
  AND2X2 AND2X2_2228 ( .A(u0_u1__abc_43657_n495), .B(u0_u1__abc_43657_n219_1_bF_buf7), .Y(u0_u1__abc_43657_n496) );
  AND2X2 AND2X2_2229 ( .A(u0_u1__abc_43657_n496), .B(u0_u1__abc_43657_n493), .Y(u0_u1_csc_16__FF_INPUT) );
  AND2X2 AND2X2_223 ( .A(u0__abc_49347_n1385), .B(u0__abc_49347_n1180_1_bF_buf3), .Y(u0__abc_49347_n1386) );
  AND2X2 AND2X2_2230 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf4), .B(u0_u1__abc_43657_n322_1), .Y(u0_u1__abc_43657_n499) );
  AND2X2 AND2X2_2231 ( .A(u0_u1__abc_43657_n500), .B(u0_u1__abc_43657_n219_1_bF_buf6), .Y(u0_u1__abc_43657_n501) );
  AND2X2 AND2X2_2232 ( .A(u0_u1__abc_43657_n501), .B(u0_u1__abc_43657_n498), .Y(u0_u1_csc_17__FF_INPUT) );
  AND2X2 AND2X2_2233 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf2), .B(u0_u1__abc_43657_n328), .Y(u0_u1__abc_43657_n504) );
  AND2X2 AND2X2_2234 ( .A(u0_u1__abc_43657_n505), .B(u0_u1__abc_43657_n219_1_bF_buf5), .Y(u0_u1__abc_43657_n506) );
  AND2X2 AND2X2_2235 ( .A(u0_u1__abc_43657_n506), .B(u0_u1__abc_43657_n503), .Y(u0_u1_csc_18__FF_INPUT) );
  AND2X2 AND2X2_2236 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf0), .B(u0_u1__abc_43657_n334), .Y(u0_u1__abc_43657_n509) );
  AND2X2 AND2X2_2237 ( .A(u0_u1__abc_43657_n510), .B(u0_u1__abc_43657_n219_1_bF_buf4), .Y(u0_u1__abc_43657_n511) );
  AND2X2 AND2X2_2238 ( .A(u0_u1__abc_43657_n511), .B(u0_u1__abc_43657_n508), .Y(u0_u1_csc_19__FF_INPUT) );
  AND2X2 AND2X2_2239 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf6), .B(u0_u1__abc_43657_n340), .Y(u0_u1__abc_43657_n514) );
  AND2X2 AND2X2_224 ( .A(spec_req_cs_3_bF_buf0), .B(u0_tms3_8_), .Y(u0__abc_49347_n1387) );
  AND2X2 AND2X2_2240 ( .A(u0_u1__abc_43657_n515), .B(u0_u1__abc_43657_n219_1_bF_buf3), .Y(u0_u1__abc_43657_n516) );
  AND2X2 AND2X2_2241 ( .A(u0_u1__abc_43657_n516), .B(u0_u1__abc_43657_n513), .Y(u0_u1_csc_20__FF_INPUT) );
  AND2X2 AND2X2_2242 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf4), .B(u0_u1__abc_43657_n346), .Y(u0_u1__abc_43657_n519) );
  AND2X2 AND2X2_2243 ( .A(u0_u1__abc_43657_n520), .B(u0_u1__abc_43657_n219_1_bF_buf2), .Y(u0_u1__abc_43657_n521) );
  AND2X2 AND2X2_2244 ( .A(u0_u1__abc_43657_n521), .B(u0_u1__abc_43657_n518), .Y(u0_u1_csc_21__FF_INPUT) );
  AND2X2 AND2X2_2245 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf2), .B(u0_u1__abc_43657_n352), .Y(u0_u1__abc_43657_n524) );
  AND2X2 AND2X2_2246 ( .A(u0_u1__abc_43657_n525), .B(u0_u1__abc_43657_n219_1_bF_buf1), .Y(u0_u1__abc_43657_n526) );
  AND2X2 AND2X2_2247 ( .A(u0_u1__abc_43657_n526), .B(u0_u1__abc_43657_n523), .Y(u0_u1_csc_22__FF_INPUT) );
  AND2X2 AND2X2_2248 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf0), .B(u0_u1__abc_43657_n358), .Y(u0_u1__abc_43657_n529) );
  AND2X2 AND2X2_2249 ( .A(u0_u1__abc_43657_n530), .B(u0_u1__abc_43657_n219_1_bF_buf0), .Y(u0_u1__abc_43657_n531) );
  AND2X2 AND2X2_225 ( .A(u0__abc_49347_n1388), .B(u0__abc_49347_n1179_bF_buf3), .Y(u0__abc_49347_n1389_1) );
  AND2X2 AND2X2_2250 ( .A(u0_u1__abc_43657_n531), .B(u0_u1__abc_43657_n528), .Y(u0_u1_csc_23__FF_INPUT) );
  AND2X2 AND2X2_2251 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf6), .B(u0_u1__abc_43657_n364), .Y(u0_u1__abc_43657_n534) );
  AND2X2 AND2X2_2252 ( .A(u0_u1__abc_43657_n535), .B(u0_u1__abc_43657_n219_1_bF_buf7), .Y(u0_u1__abc_43657_n536) );
  AND2X2 AND2X2_2253 ( .A(u0_u1__abc_43657_n536), .B(u0_u1__abc_43657_n533), .Y(u0_u1_csc_24__FF_INPUT) );
  AND2X2 AND2X2_2254 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf4), .B(u0_u1__abc_43657_n370), .Y(u0_u1__abc_43657_n539) );
  AND2X2 AND2X2_2255 ( .A(u0_u1__abc_43657_n540), .B(u0_u1__abc_43657_n219_1_bF_buf6), .Y(u0_u1__abc_43657_n541) );
  AND2X2 AND2X2_2256 ( .A(u0_u1__abc_43657_n541), .B(u0_u1__abc_43657_n538), .Y(u0_u1_csc_25__FF_INPUT) );
  AND2X2 AND2X2_2257 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf2), .B(u0_u1__abc_43657_n376), .Y(u0_u1__abc_43657_n544) );
  AND2X2 AND2X2_2258 ( .A(u0_u1__abc_43657_n545), .B(u0_u1__abc_43657_n219_1_bF_buf5), .Y(u0_u1__abc_43657_n546) );
  AND2X2 AND2X2_2259 ( .A(u0_u1__abc_43657_n546), .B(u0_u1__abc_43657_n543), .Y(u0_u1_csc_26__FF_INPUT) );
  AND2X2 AND2X2_226 ( .A(spec_req_cs_2_bF_buf0), .B(u0_tms2_8_), .Y(u0__abc_49347_n1390_1) );
  AND2X2 AND2X2_2260 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf0), .B(u0_u1__abc_43657_n382), .Y(u0_u1__abc_43657_n549) );
  AND2X2 AND2X2_2261 ( .A(u0_u1__abc_43657_n550), .B(u0_u1__abc_43657_n219_1_bF_buf4), .Y(u0_u1__abc_43657_n551) );
  AND2X2 AND2X2_2262 ( .A(u0_u1__abc_43657_n551), .B(u0_u1__abc_43657_n548), .Y(u0_u1_csc_27__FF_INPUT) );
  AND2X2 AND2X2_2263 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf6), .B(u0_u1__abc_43657_n388), .Y(u0_u1__abc_43657_n554) );
  AND2X2 AND2X2_2264 ( .A(u0_u1__abc_43657_n555), .B(u0_u1__abc_43657_n219_1_bF_buf3), .Y(u0_u1__abc_43657_n556) );
  AND2X2 AND2X2_2265 ( .A(u0_u1__abc_43657_n556), .B(u0_u1__abc_43657_n553), .Y(u0_u1_csc_28__FF_INPUT) );
  AND2X2 AND2X2_2266 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf4), .B(u0_u1__abc_43657_n394), .Y(u0_u1__abc_43657_n559) );
  AND2X2 AND2X2_2267 ( .A(u0_u1__abc_43657_n560), .B(u0_u1__abc_43657_n219_1_bF_buf2), .Y(u0_u1__abc_43657_n561) );
  AND2X2 AND2X2_2268 ( .A(u0_u1__abc_43657_n561), .B(u0_u1__abc_43657_n558), .Y(u0_u1_csc_29__FF_INPUT) );
  AND2X2 AND2X2_2269 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf2), .B(u0_u1__abc_43657_n400), .Y(u0_u1__abc_43657_n564) );
  AND2X2 AND2X2_227 ( .A(u0__abc_49347_n1391), .B(u0__abc_49347_n1178_1_bF_buf3), .Y(u0__abc_49347_n1392) );
  AND2X2 AND2X2_2270 ( .A(u0_u1__abc_43657_n565), .B(u0_u1__abc_43657_n219_1_bF_buf1), .Y(u0_u1__abc_43657_n566) );
  AND2X2 AND2X2_2271 ( .A(u0_u1__abc_43657_n566), .B(u0_u1__abc_43657_n563), .Y(u0_u1_csc_30__FF_INPUT) );
  AND2X2 AND2X2_2272 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf0), .B(u0_u1__abc_43657_n406), .Y(u0_u1__abc_43657_n569) );
  AND2X2 AND2X2_2273 ( .A(u0_u1__abc_43657_n570), .B(u0_u1__abc_43657_n219_1_bF_buf0), .Y(u0_u1__abc_43657_n571) );
  AND2X2 AND2X2_2274 ( .A(u0_u1__abc_43657_n571), .B(u0_u1__abc_43657_n568), .Y(u0_u1_csc_31__FF_INPUT) );
  AND2X2 AND2X2_2275 ( .A(u0_csc1_8_), .B(wb_we_i), .Y(u0_u1__abc_43657_n573) );
  AND2X2 AND2X2_2276 ( .A(u0_csc1_20_), .B(u0_csc_mask_4_), .Y(u0_u1__abc_43657_n574) );
  AND2X2 AND2X2_2277 ( .A(u0_csc_mask_4_), .B(wb_addr_i_25_bF_buf1), .Y(u0_u1__abc_43657_n575) );
  AND2X2 AND2X2_2278 ( .A(u0_csc_mask_3_), .B(\wb_addr_i[24] ), .Y(u0_u1__abc_43657_n578) );
  AND2X2 AND2X2_2279 ( .A(u0_csc1_19_), .B(u0_csc_mask_3_), .Y(u0_u1__abc_43657_n579) );
  AND2X2 AND2X2_228 ( .A(spec_req_cs_1_bF_buf0), .B(u0_tms1_8_), .Y(u0__abc_49347_n1393) );
  AND2X2 AND2X2_2280 ( .A(u0_u1__abc_43657_n577), .B(u0_u1__abc_43657_n581), .Y(u0_u1__abc_43657_n582) );
  AND2X2 AND2X2_2281 ( .A(u0_csc1_18_), .B(u0_csc_mask_2_), .Y(u0_u1__abc_43657_n584) );
  AND2X2 AND2X2_2282 ( .A(u0_u1__abc_43657_n584), .B(u0_u1__abc_43657_n583), .Y(u0_u1__abc_43657_n585) );
  AND2X2 AND2X2_2283 ( .A(u0_u1__abc_43657_n588), .B(u0_u1__abc_43657_n586), .Y(u0_u1__abc_43657_n589) );
  AND2X2 AND2X2_2284 ( .A(u0_u1__abc_43657_n582), .B(u0_u1__abc_43657_n589), .Y(u0_u1__abc_43657_n590) );
  AND2X2 AND2X2_2285 ( .A(u0_csc1_22_), .B(u0_csc_mask_6_), .Y(u0_u1__abc_43657_n591) );
  AND2X2 AND2X2_2286 ( .A(u0_csc_mask_6_), .B(\wb_addr_i[27] ), .Y(u0_u1__abc_43657_n592) );
  AND2X2 AND2X2_2287 ( .A(u0_csc_mask_5_), .B(\wb_addr_i[26] ), .Y(u0_u1__abc_43657_n595) );
  AND2X2 AND2X2_2288 ( .A(u0_csc1_21_), .B(u0_csc_mask_5_), .Y(u0_u1__abc_43657_n596) );
  AND2X2 AND2X2_2289 ( .A(u0_u1__abc_43657_n594), .B(u0_u1__abc_43657_n598), .Y(u0_u1__abc_43657_n599) );
  AND2X2 AND2X2_229 ( .A(u0__abc_49347_n1175_bF_buf4), .B(u0__abc_49347_n1396), .Y(u0__abc_49347_n1397) );
  AND2X2 AND2X2_2290 ( .A(u0_u1__abc_43657_n574), .B(u0_u1__abc_43657_n600), .Y(u0_u1__abc_43657_n601) );
  AND2X2 AND2X2_2291 ( .A(u0_u1__abc_43657_n604), .B(u0_u1__abc_43657_n602), .Y(u0_u1__abc_43657_n605) );
  AND2X2 AND2X2_2292 ( .A(u0_u1__abc_43657_n599), .B(u0_u1__abc_43657_n605), .Y(u0_u1__abc_43657_n606) );
  AND2X2 AND2X2_2293 ( .A(u0_u1__abc_43657_n590), .B(u0_u1__abc_43657_n606), .Y(u0_u1__abc_43657_n607) );
  AND2X2 AND2X2_2294 ( .A(u0_u1__abc_43657_n593), .B(u0_u1__abc_43657_n591), .Y(u0_u1__abc_43657_n608) );
  AND2X2 AND2X2_2295 ( .A(u0_csc_mask_7_), .B(\wb_addr_i[28] ), .Y(u0_u1__abc_43657_n610) );
  AND2X2 AND2X2_2296 ( .A(u0_csc1_23_), .B(u0_csc_mask_7_), .Y(u0_u1__abc_43657_n612) );
  AND2X2 AND2X2_2297 ( .A(u0_u1__abc_43657_n609), .B(u0_u1__abc_43657_n613), .Y(u0_u1__abc_43657_n614) );
  AND2X2 AND2X2_2298 ( .A(u0_u1__abc_43657_n614), .B(u0_u1__abc_43657_n616), .Y(u0_u1__abc_43657_n617) );
  AND2X2 AND2X2_2299 ( .A(u0_u1__abc_43657_n607), .B(u0_u1__abc_43657_n617), .Y(u0_u1__abc_43657_n618) );
  AND2X2 AND2X2_23 ( .A(_abc_55805_n305), .B(_abc_55805_n306), .Y(tms_s_5_) );
  AND2X2 AND2X2_230 ( .A(u0__abc_49347_n1395), .B(u0__abc_49347_n1397), .Y(u0__abc_49347_n1398_1) );
  AND2X2 AND2X2_2300 ( .A(u0_csc_mask_2_), .B(wb_addr_i_23_bF_buf0), .Y(u0_u1__abc_43657_n619) );
  AND2X2 AND2X2_2301 ( .A(u0_csc_mask_1_), .B(\wb_addr_i[22] ), .Y(u0_u1__abc_43657_n622) );
  AND2X2 AND2X2_2302 ( .A(u0_csc1_17_), .B(u0_csc_mask_1_), .Y(u0_u1__abc_43657_n623) );
  AND2X2 AND2X2_2303 ( .A(u0_u1__abc_43657_n621), .B(u0_u1__abc_43657_n625), .Y(u0_u1__abc_43657_n626) );
  AND2X2 AND2X2_2304 ( .A(u0_csc_mask_0_), .B(\wb_addr_i[21] ), .Y(u0_u1__abc_43657_n627) );
  AND2X2 AND2X2_2305 ( .A(u0_csc1_16_), .B(u0_csc_mask_0_), .Y(u0_u1__abc_43657_n628) );
  AND2X2 AND2X2_2306 ( .A(u0_u1__abc_43657_n630), .B(u0_u1__abc_43657_n632), .Y(u0_u1__abc_43657_n633) );
  AND2X2 AND2X2_2307 ( .A(u0_u1__abc_43657_n626), .B(u0_u1__abc_43657_n633), .Y(u0_u1__abc_43657_n634) );
  AND2X2 AND2X2_2308 ( .A(u0_u1__abc_43657_n636), .B(u0_csc1_0_), .Y(u0_u1__abc_43657_n637) );
  AND2X2 AND2X2_2309 ( .A(u0_u1__abc_43657_n634), .B(u0_u1__abc_43657_n637), .Y(u0_u1__abc_43657_n638) );
  AND2X2 AND2X2_231 ( .A(u0__abc_49347_n1176_1_bF_buf4), .B(sp_tms_9_), .Y(u0__abc_49347_n1400) );
  AND2X2 AND2X2_2310 ( .A(u0_u1__abc_43657_n618), .B(u0_u1__abc_43657_n638), .Y(u0_u1__abc_43657_n639) );
  AND2X2 AND2X2_2311 ( .A(u0_u1__abc_43657_n639), .B(u0_u1__abc_43657_n573), .Y(u0_u1_wp_err) );
  AND2X2 AND2X2_2312 ( .A(u0_u1__abc_43657_n639), .B(u0_u1__abc_43657_n641), .Y(u0_cs1) );
  AND2X2 AND2X2_2313 ( .A(u0_u1__abc_43657_n644), .B(u0_init_req1), .Y(u0_u1__abc_43657_n645) );
  AND2X2 AND2X2_2314 ( .A(u0_u1__abc_43657_n646), .B(u0_csc1_0_), .Y(u0_u1__abc_43657_n647) );
  AND2X2 AND2X2_2315 ( .A(u0_u1__abc_43657_n647), .B(u0_u1_init_req_we), .Y(u0_u1__abc_43657_n648) );
  AND2X2 AND2X2_2316 ( .A(u0_u1__abc_43657_n203_1), .B(u0_u1__abc_43657_n648), .Y(u0_u1__abc_43657_n649) );
  AND2X2 AND2X2_2317 ( .A(u0_u2_addr_r_5_), .B(u0_rf_we), .Y(u0_u2__abc_44109_n202_1) );
  AND2X2 AND2X2_2318 ( .A(u0_u2__abc_44109_n205_1), .B(u0_u2__abc_44109_n202_1), .Y(u0_u2__abc_44109_n206) );
  AND2X2 AND2X2_2319 ( .A(u0_u2__abc_44109_n206), .B(u0_u2__abc_44109_n201_1), .Y(u0_u2_init_req_we_FF_INPUT) );
  AND2X2 AND2X2_232 ( .A(spec_req_cs_5_bF_buf5), .B(u0_tms5_9_), .Y(u0__abc_49347_n1401) );
  AND2X2 AND2X2_2320 ( .A(u0_u2__abc_44109_n211_1), .B(u0_u2__abc_44109_n209_bF_buf7), .Y(u0_u2__abc_44109_n212) );
  AND2X2 AND2X2_2321 ( .A(u0_u2__abc_44109_n212), .B(u0_u2__abc_44109_n208_1), .Y(u0_u2_csc_0__FF_INPUT) );
  AND2X2 AND2X2_2322 ( .A(u0_u2__abc_44109_n215), .B(u0_u2__abc_44109_n209_bF_buf6), .Y(u0_u2__abc_44109_n216_1) );
  AND2X2 AND2X2_2323 ( .A(u0_u2__abc_44109_n216_1), .B(u0_u2__abc_44109_n214_1), .Y(u0_u2_csc_1__FF_INPUT) );
  AND2X2 AND2X2_2324 ( .A(u0_u2__abc_44109_n219_1), .B(u0_u2__abc_44109_n209_bF_buf5), .Y(u0_u2__abc_44109_n220_1) );
  AND2X2 AND2X2_2325 ( .A(u0_u2__abc_44109_n220_1), .B(u0_u2__abc_44109_n218), .Y(u0_u2_csc_2__FF_INPUT) );
  AND2X2 AND2X2_2326 ( .A(u0_u2__abc_44109_n223_1), .B(u0_u2__abc_44109_n209_bF_buf4), .Y(u0_u2__abc_44109_n224) );
  AND2X2 AND2X2_2327 ( .A(u0_u2__abc_44109_n224), .B(u0_u2__abc_44109_n222_1), .Y(u0_u2_csc_3__FF_INPUT) );
  AND2X2 AND2X2_2328 ( .A(u0_u2__abc_44109_n227), .B(u0_u2__abc_44109_n209_bF_buf3), .Y(u0_u2__abc_44109_n228_1) );
  AND2X2 AND2X2_2329 ( .A(u0_u2__abc_44109_n228_1), .B(u0_u2__abc_44109_n226_1), .Y(u0_u2_csc_4__FF_INPUT) );
  AND2X2 AND2X2_233 ( .A(u0__abc_49347_n1403), .B(u0__abc_49347_n1185_bF_buf2), .Y(u0__abc_49347_n1404) );
  AND2X2 AND2X2_2330 ( .A(u0_u2__abc_44109_n231_1), .B(u0_u2__abc_44109_n209_bF_buf2), .Y(u0_u2__abc_44109_n232_1) );
  AND2X2 AND2X2_2331 ( .A(u0_u2__abc_44109_n232_1), .B(u0_u2__abc_44109_n230), .Y(u0_u2_csc_5__FF_INPUT) );
  AND2X2 AND2X2_2332 ( .A(u0_u2__abc_44109_n235_1), .B(u0_u2__abc_44109_n209_bF_buf1), .Y(u0_u2__abc_44109_n236) );
  AND2X2 AND2X2_2333 ( .A(u0_u2__abc_44109_n236), .B(u0_u2__abc_44109_n234_1), .Y(u0_u2_csc_6__FF_INPUT) );
  AND2X2 AND2X2_2334 ( .A(u0_u2__abc_44109_n239), .B(u0_u2__abc_44109_n209_bF_buf0), .Y(u0_u2__abc_44109_n240_1) );
  AND2X2 AND2X2_2335 ( .A(u0_u2__abc_44109_n240_1), .B(u0_u2__abc_44109_n238_1), .Y(u0_u2_csc_7__FF_INPUT) );
  AND2X2 AND2X2_2336 ( .A(u0_u2__abc_44109_n243), .B(u0_u2__abc_44109_n209_bF_buf7), .Y(u0_u2__abc_44109_n244) );
  AND2X2 AND2X2_2337 ( .A(u0_u2__abc_44109_n244), .B(u0_u2__abc_44109_n242), .Y(u0_u2_csc_8__FF_INPUT) );
  AND2X2 AND2X2_2338 ( .A(u0_u2__abc_44109_n247), .B(u0_u2__abc_44109_n209_bF_buf6), .Y(u0_u2__abc_44109_n248_1) );
  AND2X2 AND2X2_2339 ( .A(u0_u2__abc_44109_n248_1), .B(u0_u2__abc_44109_n246_1), .Y(u0_u2_csc_9__FF_INPUT) );
  AND2X2 AND2X2_234 ( .A(u0__abc_49347_n1404), .B(u0__abc_49347_n1402), .Y(u0__abc_49347_n1405) );
  AND2X2 AND2X2_2340 ( .A(u0_u2__abc_44109_n251_1), .B(u0_u2__abc_44109_n209_bF_buf5), .Y(u0_u2__abc_44109_n252_1) );
  AND2X2 AND2X2_2341 ( .A(u0_u2__abc_44109_n252_1), .B(u0_u2__abc_44109_n250_1), .Y(u0_u2_csc_10__FF_INPUT) );
  AND2X2 AND2X2_2342 ( .A(u0_u2__abc_44109_n255), .B(u0_u2__abc_44109_n209_bF_buf4), .Y(u0_u2__abc_44109_n256_1) );
  AND2X2 AND2X2_2343 ( .A(u0_u2__abc_44109_n256_1), .B(u0_u2__abc_44109_n254), .Y(u0_u2_csc_11__FF_INPUT) );
  AND2X2 AND2X2_2344 ( .A(u0_u2__abc_44109_n259_1), .B(u0_u2__abc_44109_n209_bF_buf3), .Y(u0_u2__abc_44109_n260_1) );
  AND2X2 AND2X2_2345 ( .A(u0_u2__abc_44109_n260_1), .B(u0_u2__abc_44109_n258_1), .Y(u0_u2_csc_12__FF_INPUT) );
  AND2X2 AND2X2_2346 ( .A(u0_u2__abc_44109_n263_1), .B(u0_u2__abc_44109_n209_bF_buf2), .Y(u0_u2__abc_44109_n264) );
  AND2X2 AND2X2_2347 ( .A(u0_u2__abc_44109_n264), .B(u0_u2__abc_44109_n262), .Y(u0_u2_csc_13__FF_INPUT) );
  AND2X2 AND2X2_2348 ( .A(u0_u2__abc_44109_n267), .B(u0_u2__abc_44109_n209_bF_buf1), .Y(u0_u2__abc_44109_n268_1) );
  AND2X2 AND2X2_2349 ( .A(u0_u2__abc_44109_n268_1), .B(u0_u2__abc_44109_n266), .Y(u0_u2_csc_14__FF_INPUT) );
  AND2X2 AND2X2_235 ( .A(u0__abc_49347_n1406), .B(u0__abc_49347_n1181_bF_buf2), .Y(u0__abc_49347_n1407_1) );
  AND2X2 AND2X2_2350 ( .A(u0_u2__abc_44109_n271), .B(u0_u2__abc_44109_n209_bF_buf0), .Y(u0_u2__abc_44109_n272) );
  AND2X2 AND2X2_2351 ( .A(u0_u2__abc_44109_n272), .B(u0_u2__abc_44109_n270_1), .Y(u0_u2_csc_15__FF_INPUT) );
  AND2X2 AND2X2_2352 ( .A(u0_u2__abc_44109_n275), .B(u0_u2__abc_44109_n209_bF_buf7), .Y(u0_u2__abc_44109_n276_1) );
  AND2X2 AND2X2_2353 ( .A(u0_u2__abc_44109_n276_1), .B(u0_u2__abc_44109_n274_1), .Y(u0_u2_csc_16__FF_INPUT) );
  AND2X2 AND2X2_2354 ( .A(u0_u2__abc_44109_n279), .B(u0_u2__abc_44109_n209_bF_buf6), .Y(u0_u2__abc_44109_n280) );
  AND2X2 AND2X2_2355 ( .A(u0_u2__abc_44109_n280), .B(u0_u2__abc_44109_n278), .Y(u0_u2_csc_17__FF_INPUT) );
  AND2X2 AND2X2_2356 ( .A(u0_u2__abc_44109_n283_1), .B(u0_u2__abc_44109_n209_bF_buf5), .Y(u0_u2__abc_44109_n284) );
  AND2X2 AND2X2_2357 ( .A(u0_u2__abc_44109_n284), .B(u0_u2__abc_44109_n282), .Y(u0_u2_csc_18__FF_INPUT) );
  AND2X2 AND2X2_2358 ( .A(u0_u2__abc_44109_n287_1), .B(u0_u2__abc_44109_n209_bF_buf4), .Y(u0_u2__abc_44109_n288) );
  AND2X2 AND2X2_2359 ( .A(u0_u2__abc_44109_n288), .B(u0_u2__abc_44109_n286), .Y(u0_u2_csc_19__FF_INPUT) );
  AND2X2 AND2X2_236 ( .A(spec_req_cs_4_bF_buf5), .B(u0_tms4_9_), .Y(u0__abc_49347_n1408_1) );
  AND2X2 AND2X2_2360 ( .A(u0_u2__abc_44109_n291_1), .B(u0_u2__abc_44109_n209_bF_buf3), .Y(u0_u2__abc_44109_n292) );
  AND2X2 AND2X2_2361 ( .A(u0_u2__abc_44109_n292), .B(u0_u2__abc_44109_n290), .Y(u0_u2_csc_20__FF_INPUT) );
  AND2X2 AND2X2_2362 ( .A(u0_u2__abc_44109_n295_1), .B(u0_u2__abc_44109_n209_bF_buf2), .Y(u0_u2__abc_44109_n296) );
  AND2X2 AND2X2_2363 ( .A(u0_u2__abc_44109_n296), .B(u0_u2__abc_44109_n294), .Y(u0_u2_csc_21__FF_INPUT) );
  AND2X2 AND2X2_2364 ( .A(u0_u2__abc_44109_n299), .B(u0_u2__abc_44109_n209_bF_buf1), .Y(u0_u2__abc_44109_n300) );
  AND2X2 AND2X2_2365 ( .A(u0_u2__abc_44109_n300), .B(u0_u2__abc_44109_n298), .Y(u0_u2_csc_22__FF_INPUT) );
  AND2X2 AND2X2_2366 ( .A(u0_u2__abc_44109_n303), .B(u0_u2__abc_44109_n209_bF_buf0), .Y(u0_u2__abc_44109_n304_1) );
  AND2X2 AND2X2_2367 ( .A(u0_u2__abc_44109_n304_1), .B(u0_u2__abc_44109_n302), .Y(u0_u2_csc_23__FF_INPUT) );
  AND2X2 AND2X2_2368 ( .A(u0_u2__abc_44109_n307), .B(u0_u2__abc_44109_n209_bF_buf7), .Y(u0_u2__abc_44109_n308) );
  AND2X2 AND2X2_2369 ( .A(u0_u2__abc_44109_n308), .B(u0_u2__abc_44109_n306_1), .Y(u0_u2_csc_24__FF_INPUT) );
  AND2X2 AND2X2_237 ( .A(u0__abc_49347_n1409), .B(u0__abc_49347_n1180_1_bF_buf2), .Y(u0__abc_49347_n1410) );
  AND2X2 AND2X2_2370 ( .A(u0_u2__abc_44109_n311), .B(u0_u2__abc_44109_n209_bF_buf6), .Y(u0_u2__abc_44109_n312) );
  AND2X2 AND2X2_2371 ( .A(u0_u2__abc_44109_n312), .B(u0_u2__abc_44109_n310), .Y(u0_u2_csc_25__FF_INPUT) );
  AND2X2 AND2X2_2372 ( .A(u0_u2__abc_44109_n315), .B(u0_u2__abc_44109_n209_bF_buf5), .Y(u0_u2__abc_44109_n316) );
  AND2X2 AND2X2_2373 ( .A(u0_u2__abc_44109_n316), .B(u0_u2__abc_44109_n314), .Y(u0_u2_csc_26__FF_INPUT) );
  AND2X2 AND2X2_2374 ( .A(u0_u2__abc_44109_n319), .B(u0_u2__abc_44109_n209_bF_buf4), .Y(u0_u2__abc_44109_n320_1) );
  AND2X2 AND2X2_2375 ( .A(u0_u2__abc_44109_n320_1), .B(u0_u2__abc_44109_n318_1), .Y(u0_u2_csc_27__FF_INPUT) );
  AND2X2 AND2X2_2376 ( .A(u0_u2__abc_44109_n323_1), .B(u0_u2__abc_44109_n209_bF_buf3), .Y(u0_u2__abc_44109_n324_1) );
  AND2X2 AND2X2_2377 ( .A(u0_u2__abc_44109_n324_1), .B(u0_u2__abc_44109_n322_1), .Y(u0_u2_csc_28__FF_INPUT) );
  AND2X2 AND2X2_2378 ( .A(u0_u2__abc_44109_n327), .B(u0_u2__abc_44109_n209_bF_buf2), .Y(u0_u2__abc_44109_n328) );
  AND2X2 AND2X2_2379 ( .A(u0_u2__abc_44109_n328), .B(u0_u2__abc_44109_n326), .Y(u0_u2_csc_29__FF_INPUT) );
  AND2X2 AND2X2_238 ( .A(spec_req_cs_3_bF_buf5), .B(u0_tms3_9_), .Y(u0__abc_49347_n1411) );
  AND2X2 AND2X2_2380 ( .A(u0_u2__abc_44109_n331), .B(u0_u2__abc_44109_n209_bF_buf1), .Y(u0_u2__abc_44109_n332) );
  AND2X2 AND2X2_2381 ( .A(u0_u2__abc_44109_n332), .B(u0_u2__abc_44109_n330), .Y(u0_u2_csc_30__FF_INPUT) );
  AND2X2 AND2X2_2382 ( .A(u0_u2__abc_44109_n335), .B(u0_u2__abc_44109_n209_bF_buf0), .Y(u0_u2__abc_44109_n336) );
  AND2X2 AND2X2_2383 ( .A(u0_u2__abc_44109_n336), .B(u0_u2__abc_44109_n334), .Y(u0_u2_csc_31__FF_INPUT) );
  AND2X2 AND2X2_2384 ( .A(u0_u2__abc_44109_n206), .B(u0_u2_addr_r_2_), .Y(u0_u2_lmr_req_we_FF_INPUT) );
  AND2X2 AND2X2_2385 ( .A(u0_u2__abc_44109_n341), .B(u0_u2__abc_44109_n209_bF_buf7), .Y(u0_u2__abc_44109_n342) );
  AND2X2 AND2X2_2386 ( .A(u0_u2__abc_44109_n342), .B(u0_u2__abc_44109_n339), .Y(u0_u2_tms_0__FF_INPUT) );
  AND2X2 AND2X2_2387 ( .A(u0_u2__abc_44109_n345), .B(u0_u2__abc_44109_n209_bF_buf6), .Y(u0_u2__abc_44109_n346) );
  AND2X2 AND2X2_2388 ( .A(u0_u2__abc_44109_n346), .B(u0_u2__abc_44109_n344), .Y(u0_u2_tms_1__FF_INPUT) );
  AND2X2 AND2X2_2389 ( .A(u0_u2__abc_44109_n349), .B(u0_u2__abc_44109_n209_bF_buf5), .Y(u0_u2__abc_44109_n350) );
  AND2X2 AND2X2_239 ( .A(u0__abc_49347_n1412), .B(u0__abc_49347_n1179_bF_buf2), .Y(u0__abc_49347_n1413) );
  AND2X2 AND2X2_2390 ( .A(u0_u2__abc_44109_n350), .B(u0_u2__abc_44109_n348), .Y(u0_u2_tms_2__FF_INPUT) );
  AND2X2 AND2X2_2391 ( .A(u0_u2__abc_44109_n353), .B(u0_u2__abc_44109_n209_bF_buf4), .Y(u0_u2__abc_44109_n354) );
  AND2X2 AND2X2_2392 ( .A(u0_u2__abc_44109_n354), .B(u0_u2__abc_44109_n352), .Y(u0_u2_tms_3__FF_INPUT) );
  AND2X2 AND2X2_2393 ( .A(u0_u2__abc_44109_n357), .B(u0_u2__abc_44109_n209_bF_buf3), .Y(u0_u2__abc_44109_n358) );
  AND2X2 AND2X2_2394 ( .A(u0_u2__abc_44109_n358), .B(u0_u2__abc_44109_n356), .Y(u0_u2_tms_4__FF_INPUT) );
  AND2X2 AND2X2_2395 ( .A(u0_u2__abc_44109_n361), .B(u0_u2__abc_44109_n209_bF_buf2), .Y(u0_u2__abc_44109_n362) );
  AND2X2 AND2X2_2396 ( .A(u0_u2__abc_44109_n362), .B(u0_u2__abc_44109_n360), .Y(u0_u2_tms_5__FF_INPUT) );
  AND2X2 AND2X2_2397 ( .A(u0_u2__abc_44109_n365), .B(u0_u2__abc_44109_n209_bF_buf1), .Y(u0_u2__abc_44109_n366) );
  AND2X2 AND2X2_2398 ( .A(u0_u2__abc_44109_n366), .B(u0_u2__abc_44109_n364), .Y(u0_u2_tms_6__FF_INPUT) );
  AND2X2 AND2X2_2399 ( .A(u0_u2__abc_44109_n369), .B(u0_u2__abc_44109_n209_bF_buf0), .Y(u0_u2__abc_44109_n370) );
  AND2X2 AND2X2_24 ( .A(_abc_55805_n308), .B(_abc_55805_n309), .Y(tms_s_6_) );
  AND2X2 AND2X2_240 ( .A(spec_req_cs_2_bF_buf5), .B(u0_tms2_9_), .Y(u0__abc_49347_n1414) );
  AND2X2 AND2X2_2400 ( .A(u0_u2__abc_44109_n370), .B(u0_u2__abc_44109_n368), .Y(u0_u2_tms_7__FF_INPUT) );
  AND2X2 AND2X2_2401 ( .A(u0_u2__abc_44109_n373), .B(u0_u2__abc_44109_n209_bF_buf7), .Y(u0_u2__abc_44109_n374) );
  AND2X2 AND2X2_2402 ( .A(u0_u2__abc_44109_n374), .B(u0_u2__abc_44109_n372), .Y(u0_u2_tms_8__FF_INPUT) );
  AND2X2 AND2X2_2403 ( .A(u0_u2__abc_44109_n377), .B(u0_u2__abc_44109_n209_bF_buf6), .Y(u0_u2__abc_44109_n378) );
  AND2X2 AND2X2_2404 ( .A(u0_u2__abc_44109_n378), .B(u0_u2__abc_44109_n376), .Y(u0_u2_tms_9__FF_INPUT) );
  AND2X2 AND2X2_2405 ( .A(u0_u2__abc_44109_n381), .B(u0_u2__abc_44109_n209_bF_buf5), .Y(u0_u2__abc_44109_n382) );
  AND2X2 AND2X2_2406 ( .A(u0_u2__abc_44109_n382), .B(u0_u2__abc_44109_n380), .Y(u0_u2_tms_10__FF_INPUT) );
  AND2X2 AND2X2_2407 ( .A(u0_u2__abc_44109_n385), .B(u0_u2__abc_44109_n209_bF_buf4), .Y(u0_u2__abc_44109_n386) );
  AND2X2 AND2X2_2408 ( .A(u0_u2__abc_44109_n386), .B(u0_u2__abc_44109_n384), .Y(u0_u2_tms_11__FF_INPUT) );
  AND2X2 AND2X2_2409 ( .A(u0_u2__abc_44109_n389), .B(u0_u2__abc_44109_n209_bF_buf3), .Y(u0_u2__abc_44109_n390) );
  AND2X2 AND2X2_241 ( .A(u0__abc_49347_n1415), .B(u0__abc_49347_n1178_1_bF_buf2), .Y(u0__abc_49347_n1416_1) );
  AND2X2 AND2X2_2410 ( .A(u0_u2__abc_44109_n390), .B(u0_u2__abc_44109_n388), .Y(u0_u2_tms_12__FF_INPUT) );
  AND2X2 AND2X2_2411 ( .A(u0_u2__abc_44109_n393), .B(u0_u2__abc_44109_n209_bF_buf2), .Y(u0_u2__abc_44109_n394) );
  AND2X2 AND2X2_2412 ( .A(u0_u2__abc_44109_n394), .B(u0_u2__abc_44109_n392), .Y(u0_u2_tms_13__FF_INPUT) );
  AND2X2 AND2X2_2413 ( .A(u0_u2__abc_44109_n397), .B(u0_u2__abc_44109_n209_bF_buf1), .Y(u0_u2__abc_44109_n398) );
  AND2X2 AND2X2_2414 ( .A(u0_u2__abc_44109_n398), .B(u0_u2__abc_44109_n396), .Y(u0_u2_tms_14__FF_INPUT) );
  AND2X2 AND2X2_2415 ( .A(u0_u2__abc_44109_n401), .B(u0_u2__abc_44109_n209_bF_buf0), .Y(u0_u2__abc_44109_n402) );
  AND2X2 AND2X2_2416 ( .A(u0_u2__abc_44109_n402), .B(u0_u2__abc_44109_n400), .Y(u0_u2_tms_15__FF_INPUT) );
  AND2X2 AND2X2_2417 ( .A(u0_u2__abc_44109_n405), .B(u0_u2__abc_44109_n209_bF_buf7), .Y(u0_u2__abc_44109_n406) );
  AND2X2 AND2X2_2418 ( .A(u0_u2__abc_44109_n406), .B(u0_u2__abc_44109_n404), .Y(u0_u2_tms_16__FF_INPUT) );
  AND2X2 AND2X2_2419 ( .A(u0_u2__abc_44109_n409), .B(u0_u2__abc_44109_n209_bF_buf6), .Y(u0_u2__abc_44109_n410) );
  AND2X2 AND2X2_242 ( .A(spec_req_cs_1_bF_buf5), .B(u0_tms1_9_), .Y(u0__abc_49347_n1417_1) );
  AND2X2 AND2X2_2420 ( .A(u0_u2__abc_44109_n410), .B(u0_u2__abc_44109_n408), .Y(u0_u2_tms_17__FF_INPUT) );
  AND2X2 AND2X2_2421 ( .A(u0_u2__abc_44109_n413), .B(u0_u2__abc_44109_n209_bF_buf5), .Y(u0_u2__abc_44109_n414) );
  AND2X2 AND2X2_2422 ( .A(u0_u2__abc_44109_n414), .B(u0_u2__abc_44109_n412), .Y(u0_u2_tms_18__FF_INPUT) );
  AND2X2 AND2X2_2423 ( .A(u0_u2__abc_44109_n417), .B(u0_u2__abc_44109_n209_bF_buf4), .Y(u0_u2__abc_44109_n418) );
  AND2X2 AND2X2_2424 ( .A(u0_u2__abc_44109_n418), .B(u0_u2__abc_44109_n416), .Y(u0_u2_tms_19__FF_INPUT) );
  AND2X2 AND2X2_2425 ( .A(u0_u2__abc_44109_n421), .B(u0_u2__abc_44109_n209_bF_buf3), .Y(u0_u2__abc_44109_n422) );
  AND2X2 AND2X2_2426 ( .A(u0_u2__abc_44109_n422), .B(u0_u2__abc_44109_n420), .Y(u0_u2_tms_20__FF_INPUT) );
  AND2X2 AND2X2_2427 ( .A(u0_u2__abc_44109_n425), .B(u0_u2__abc_44109_n209_bF_buf2), .Y(u0_u2__abc_44109_n426) );
  AND2X2 AND2X2_2428 ( .A(u0_u2__abc_44109_n426), .B(u0_u2__abc_44109_n424), .Y(u0_u2_tms_21__FF_INPUT) );
  AND2X2 AND2X2_2429 ( .A(u0_u2__abc_44109_n429), .B(u0_u2__abc_44109_n209_bF_buf1), .Y(u0_u2__abc_44109_n430) );
  AND2X2 AND2X2_243 ( .A(u0__abc_49347_n1175_bF_buf3), .B(u0__abc_49347_n1420), .Y(u0__abc_49347_n1421) );
  AND2X2 AND2X2_2430 ( .A(u0_u2__abc_44109_n430), .B(u0_u2__abc_44109_n428), .Y(u0_u2_tms_22__FF_INPUT) );
  AND2X2 AND2X2_2431 ( .A(u0_u2__abc_44109_n433), .B(u0_u2__abc_44109_n209_bF_buf0), .Y(u0_u2__abc_44109_n434) );
  AND2X2 AND2X2_2432 ( .A(u0_u2__abc_44109_n434), .B(u0_u2__abc_44109_n432), .Y(u0_u2_tms_23__FF_INPUT) );
  AND2X2 AND2X2_2433 ( .A(u0_u2__abc_44109_n437), .B(u0_u2__abc_44109_n209_bF_buf7), .Y(u0_u2__abc_44109_n438) );
  AND2X2 AND2X2_2434 ( .A(u0_u2__abc_44109_n438), .B(u0_u2__abc_44109_n436), .Y(u0_u2_tms_24__FF_INPUT) );
  AND2X2 AND2X2_2435 ( .A(u0_u2__abc_44109_n441), .B(u0_u2__abc_44109_n209_bF_buf6), .Y(u0_u2__abc_44109_n442) );
  AND2X2 AND2X2_2436 ( .A(u0_u2__abc_44109_n442), .B(u0_u2__abc_44109_n440), .Y(u0_u2_tms_25__FF_INPUT) );
  AND2X2 AND2X2_2437 ( .A(u0_u2__abc_44109_n445), .B(u0_u2__abc_44109_n209_bF_buf5), .Y(u0_u2__abc_44109_n446) );
  AND2X2 AND2X2_2438 ( .A(u0_u2__abc_44109_n446), .B(u0_u2__abc_44109_n444), .Y(u0_u2_tms_26__FF_INPUT) );
  AND2X2 AND2X2_2439 ( .A(u0_u2__abc_44109_n449), .B(u0_u2__abc_44109_n209_bF_buf4), .Y(u0_u2__abc_44109_n450) );
  AND2X2 AND2X2_244 ( .A(u0__abc_49347_n1419), .B(u0__abc_49347_n1421), .Y(u0__abc_49347_n1422) );
  AND2X2 AND2X2_2440 ( .A(u0_u2__abc_44109_n450), .B(u0_u2__abc_44109_n448), .Y(u0_u2_tms_27__FF_INPUT) );
  AND2X2 AND2X2_2441 ( .A(u0_u2__abc_44109_n453), .B(u0_u2__abc_44109_n209_bF_buf3), .Y(u0_u2__abc_44109_n454) );
  AND2X2 AND2X2_2442 ( .A(u0_u2__abc_44109_n454), .B(u0_u2__abc_44109_n452), .Y(u0_u2_tms_28__FF_INPUT) );
  AND2X2 AND2X2_2443 ( .A(u0_u2__abc_44109_n457), .B(u0_u2__abc_44109_n209_bF_buf2), .Y(u0_u2__abc_44109_n458) );
  AND2X2 AND2X2_2444 ( .A(u0_u2__abc_44109_n458), .B(u0_u2__abc_44109_n456), .Y(u0_u2_tms_29__FF_INPUT) );
  AND2X2 AND2X2_2445 ( .A(u0_u2__abc_44109_n461), .B(u0_u2__abc_44109_n209_bF_buf1), .Y(u0_u2__abc_44109_n462) );
  AND2X2 AND2X2_2446 ( .A(u0_u2__abc_44109_n462), .B(u0_u2__abc_44109_n460), .Y(u0_u2_tms_30__FF_INPUT) );
  AND2X2 AND2X2_2447 ( .A(u0_u2__abc_44109_n465), .B(u0_u2__abc_44109_n209_bF_buf0), .Y(u0_u2__abc_44109_n466) );
  AND2X2 AND2X2_2448 ( .A(u0_u2__abc_44109_n466), .B(u0_u2__abc_44109_n464), .Y(u0_u2_tms_31__FF_INPUT) );
  AND2X2 AND2X2_2449 ( .A(u0_u2__abc_44109_n470), .B(u0_u2_lmr_req_we), .Y(u0_u2__abc_44109_n471) );
  AND2X2 AND2X2_245 ( .A(u0__abc_49347_n1176_1_bF_buf3), .B(sp_tms_10_), .Y(u0__abc_49347_n1424) );
  AND2X2 AND2X2_2450 ( .A(u0_u2__abc_44109_n471), .B(u0_u2_inited), .Y(u0_u2__abc_44109_n472) );
  AND2X2 AND2X2_2451 ( .A(u0_u2__abc_44109_n474), .B(u0_lmr_req2), .Y(u0_u2__abc_44109_n475) );
  AND2X2 AND2X2_2452 ( .A(u0_u2__abc_44109_n473), .B(u0_u2__abc_44109_n475), .Y(u0_u2__abc_44109_n476) );
  AND2X2 AND2X2_2453 ( .A(u0_u2__abc_44109_n478), .B(u0_init_req2), .Y(u0_u2__abc_44109_n479) );
  AND2X2 AND2X2_2454 ( .A(u0_u2__abc_44109_n480), .B(u0_csc2_0_), .Y(u0_u2__abc_44109_n481) );
  AND2X2 AND2X2_2455 ( .A(u0_u2__abc_44109_n481), .B(u0_u2_init_req_we), .Y(u0_u2__abc_44109_n482) );
  AND2X2 AND2X2_2456 ( .A(u0_u2__abc_44109_n470), .B(u0_u2__abc_44109_n482), .Y(u0_u2__abc_44109_n483) );
  AND2X2 AND2X2_2457 ( .A(u0_csc2_8_), .B(wb_we_i), .Y(u0_u2__abc_44109_n486) );
  AND2X2 AND2X2_2458 ( .A(u0_csc2_20_), .B(u0_csc_mask_4_), .Y(u0_u2__abc_44109_n487) );
  AND2X2 AND2X2_2459 ( .A(u0_csc_mask_4_), .B(wb_addr_i_25_bF_buf3), .Y(u0_u2__abc_44109_n488) );
  AND2X2 AND2X2_246 ( .A(spec_req_cs_5_bF_buf4), .B(u0_tms5_10_), .Y(u0__abc_49347_n1425_1) );
  AND2X2 AND2X2_2460 ( .A(u0_csc_mask_3_), .B(\wb_addr_i[24] ), .Y(u0_u2__abc_44109_n491) );
  AND2X2 AND2X2_2461 ( .A(u0_csc2_19_), .B(u0_csc_mask_3_), .Y(u0_u2__abc_44109_n492) );
  AND2X2 AND2X2_2462 ( .A(u0_u2__abc_44109_n490), .B(u0_u2__abc_44109_n494), .Y(u0_u2__abc_44109_n495) );
  AND2X2 AND2X2_2463 ( .A(u0_csc2_18_), .B(u0_csc_mask_2_), .Y(u0_u2__abc_44109_n497) );
  AND2X2 AND2X2_2464 ( .A(u0_u2__abc_44109_n497), .B(u0_u2__abc_44109_n496), .Y(u0_u2__abc_44109_n498) );
  AND2X2 AND2X2_2465 ( .A(u0_u2__abc_44109_n501), .B(u0_u2__abc_44109_n499), .Y(u0_u2__abc_44109_n502) );
  AND2X2 AND2X2_2466 ( .A(u0_u2__abc_44109_n495), .B(u0_u2__abc_44109_n502), .Y(u0_u2__abc_44109_n503) );
  AND2X2 AND2X2_2467 ( .A(u0_csc2_22_), .B(u0_csc_mask_6_), .Y(u0_u2__abc_44109_n504) );
  AND2X2 AND2X2_2468 ( .A(u0_csc_mask_6_), .B(\wb_addr_i[27] ), .Y(u0_u2__abc_44109_n505) );
  AND2X2 AND2X2_2469 ( .A(u0_csc_mask_5_), .B(\wb_addr_i[26] ), .Y(u0_u2__abc_44109_n508) );
  AND2X2 AND2X2_247 ( .A(u0__abc_49347_n1427), .B(u0__abc_49347_n1185_bF_buf1), .Y(u0__abc_49347_n1428) );
  AND2X2 AND2X2_2470 ( .A(u0_csc2_21_), .B(u0_csc_mask_5_), .Y(u0_u2__abc_44109_n509) );
  AND2X2 AND2X2_2471 ( .A(u0_u2__abc_44109_n507), .B(u0_u2__abc_44109_n511), .Y(u0_u2__abc_44109_n512) );
  AND2X2 AND2X2_2472 ( .A(u0_u2__abc_44109_n487), .B(u0_u2__abc_44109_n513), .Y(u0_u2__abc_44109_n514) );
  AND2X2 AND2X2_2473 ( .A(u0_u2__abc_44109_n517), .B(u0_u2__abc_44109_n515), .Y(u0_u2__abc_44109_n518) );
  AND2X2 AND2X2_2474 ( .A(u0_u2__abc_44109_n512), .B(u0_u2__abc_44109_n518), .Y(u0_u2__abc_44109_n519) );
  AND2X2 AND2X2_2475 ( .A(u0_u2__abc_44109_n503), .B(u0_u2__abc_44109_n519), .Y(u0_u2__abc_44109_n520) );
  AND2X2 AND2X2_2476 ( .A(u0_u2__abc_44109_n506), .B(u0_u2__abc_44109_n504), .Y(u0_u2__abc_44109_n521) );
  AND2X2 AND2X2_2477 ( .A(u0_csc_mask_7_), .B(\wb_addr_i[28] ), .Y(u0_u2__abc_44109_n523) );
  AND2X2 AND2X2_2478 ( .A(u0_csc2_23_), .B(u0_csc_mask_7_), .Y(u0_u2__abc_44109_n525) );
  AND2X2 AND2X2_2479 ( .A(u0_u2__abc_44109_n522), .B(u0_u2__abc_44109_n526), .Y(u0_u2__abc_44109_n527) );
  AND2X2 AND2X2_248 ( .A(u0__abc_49347_n1428), .B(u0__abc_49347_n1426_1), .Y(u0__abc_49347_n1429) );
  AND2X2 AND2X2_2480 ( .A(u0_u2__abc_44109_n527), .B(u0_u2__abc_44109_n529), .Y(u0_u2__abc_44109_n530) );
  AND2X2 AND2X2_2481 ( .A(u0_u2__abc_44109_n520), .B(u0_u2__abc_44109_n530), .Y(u0_u2__abc_44109_n531) );
  AND2X2 AND2X2_2482 ( .A(u0_csc_mask_2_), .B(wb_addr_i_23_bF_buf2), .Y(u0_u2__abc_44109_n532) );
  AND2X2 AND2X2_2483 ( .A(u0_csc_mask_1_), .B(\wb_addr_i[22] ), .Y(u0_u2__abc_44109_n535) );
  AND2X2 AND2X2_2484 ( .A(u0_csc2_17_), .B(u0_csc_mask_1_), .Y(u0_u2__abc_44109_n536) );
  AND2X2 AND2X2_2485 ( .A(u0_u2__abc_44109_n534), .B(u0_u2__abc_44109_n538), .Y(u0_u2__abc_44109_n539) );
  AND2X2 AND2X2_2486 ( .A(u0_csc_mask_0_), .B(\wb_addr_i[21] ), .Y(u0_u2__abc_44109_n540) );
  AND2X2 AND2X2_2487 ( .A(u0_csc2_16_), .B(u0_csc_mask_0_), .Y(u0_u2__abc_44109_n541) );
  AND2X2 AND2X2_2488 ( .A(u0_u2__abc_44109_n543), .B(u0_u2__abc_44109_n545), .Y(u0_u2__abc_44109_n546) );
  AND2X2 AND2X2_2489 ( .A(u0_u2__abc_44109_n539), .B(u0_u2__abc_44109_n546), .Y(u0_u2__abc_44109_n547) );
  AND2X2 AND2X2_249 ( .A(u0__abc_49347_n1430), .B(u0__abc_49347_n1181_bF_buf1), .Y(u0__abc_49347_n1431) );
  AND2X2 AND2X2_2490 ( .A(u0_u2__abc_44109_n549), .B(u0_csc2_0_), .Y(u0_u2__abc_44109_n550) );
  AND2X2 AND2X2_2491 ( .A(u0_u2__abc_44109_n547), .B(u0_u2__abc_44109_n550), .Y(u0_u2__abc_44109_n551) );
  AND2X2 AND2X2_2492 ( .A(u0_u2__abc_44109_n531), .B(u0_u2__abc_44109_n551), .Y(u0_u2__abc_44109_n552) );
  AND2X2 AND2X2_2493 ( .A(u0_u2__abc_44109_n552), .B(u0_u2__abc_44109_n486), .Y(u0_u2_wp_err) );
  AND2X2 AND2X2_2494 ( .A(u0_u2__abc_44109_n552), .B(u0_u2__abc_44109_n554), .Y(u0_cs2) );
  AND2X2 AND2X2_2495 ( .A(u0_u3__abc_44466_n207), .B(u0_u3__abc_44466_n208_1), .Y(u0_u3__abc_44466_n209_1) );
  AND2X2 AND2X2_2496 ( .A(u0_u3_addr_r_5_), .B(u0_u3_addr_r_3_), .Y(u0_u3__abc_44466_n210) );
  AND2X2 AND2X2_2497 ( .A(u0_u3__abc_44466_n210), .B(u0_rf_we), .Y(u0_u3__abc_44466_n211_1) );
  AND2X2 AND2X2_2498 ( .A(u0_u3__abc_44466_n211_1), .B(u0_u3__abc_44466_n209_1), .Y(u0_u3__abc_44466_n212_1) );
  AND2X2 AND2X2_2499 ( .A(u0_u3__abc_44466_n212_1), .B(u0_u3__abc_44466_n206_1), .Y(u0_u3_init_req_we_FF_INPUT) );
  AND2X2 AND2X2_25 ( .A(_abc_55805_n311), .B(_abc_55805_n312), .Y(tms_s_7_) );
  AND2X2 AND2X2_250 ( .A(spec_req_cs_4_bF_buf4), .B(u0_tms4_10_), .Y(u0__abc_49347_n1432) );
  AND2X2 AND2X2_2500 ( .A(u0_u3_init_req_we_FF_INPUT_bF_buf4), .B(u0_u3__abc_44466_n215_1), .Y(u0_u3__abc_44466_n216) );
  AND2X2 AND2X2_2501 ( .A(u0_u3__abc_44466_n217_1), .B(u0_u3__abc_44466_n214_1), .Y(u0_u3__abc_44466_n218_1) );
  AND2X2 AND2X2_2502 ( .A(u0_u3__abc_44466_n218_1), .B(u0_u3__abc_44466_n205_1_bF_buf4), .Y(u0_u3__abc_44466_n219) );
  AND2X2 AND2X2_2503 ( .A(u0_u3_rst_r2_bF_buf4), .B(_auto_iopadmap_cc_313_execute_56321_2_), .Y(u0_u3__abc_44466_n220_1) );
  AND2X2 AND2X2_2504 ( .A(u0_u3_rst_r2_bF_buf3), .B(_auto_iopadmap_cc_313_execute_56321_3_), .Y(u0_u3__abc_44466_n221_1) );
  AND2X2 AND2X2_2505 ( .A(u0_u3_init_req_we_FF_INPUT_bF_buf2), .B(u0_u3__abc_44466_n225), .Y(u0_u3__abc_44466_n226_1) );
  AND2X2 AND2X2_2506 ( .A(u0_u3__abc_44466_n227_1), .B(u0_u3__abc_44466_n205_1_bF_buf3), .Y(u0_u3__abc_44466_n228) );
  AND2X2 AND2X2_2507 ( .A(u0_u3__abc_44466_n228), .B(u0_u3__abc_44466_n224_1), .Y(u0_u3__abc_44466_n229_1) );
  AND2X2 AND2X2_2508 ( .A(u0_u3_init_req_we_FF_INPUT_bF_buf0), .B(u0_u3__abc_44466_n232_1), .Y(u0_u3__abc_44466_n233_1) );
  AND2X2 AND2X2_2509 ( .A(u0_u3__abc_44466_n234), .B(u0_u3__abc_44466_n205_1_bF_buf2), .Y(u0_u3__abc_44466_n235_1) );
  AND2X2 AND2X2_251 ( .A(u0__abc_49347_n1433), .B(u0__abc_49347_n1180_1_bF_buf1), .Y(u0__abc_49347_n1434_1) );
  AND2X2 AND2X2_2510 ( .A(u0_u3__abc_44466_n235_1), .B(u0_u3__abc_44466_n231), .Y(u0_u3__abc_44466_n236_1) );
  AND2X2 AND2X2_2511 ( .A(u0_u3_init_req_we_FF_INPUT_bF_buf5), .B(\wb_data_i[3] ), .Y(u0_u3__abc_44466_n238_1) );
  AND2X2 AND2X2_2512 ( .A(u0_u3__abc_44466_n239_1_bF_buf4), .B(u0_csc3_3_), .Y(u0_u3__abc_44466_n240) );
  AND2X2 AND2X2_2513 ( .A(u0_u3__abc_44466_n241_1), .B(u0_u3__abc_44466_n205_1_bF_buf1), .Y(u0_u3_csc_3__FF_INPUT) );
  AND2X2 AND2X2_2514 ( .A(u0_u3_init_req_we_FF_INPUT_bF_buf2), .B(u0_u3__abc_44466_n244_1), .Y(u0_u3__abc_44466_n245_1) );
  AND2X2 AND2X2_2515 ( .A(u0_u3__abc_44466_n246), .B(u0_u3__abc_44466_n243), .Y(u0_u3__abc_44466_n247) );
  AND2X2 AND2X2_2516 ( .A(u0_u3__abc_44466_n248), .B(u0_u3__abc_44466_n249), .Y(u0_u3_csc_4__FF_INPUT) );
  AND2X2 AND2X2_2517 ( .A(u0_u3_init_req_we_FF_INPUT_bF_buf0), .B(u0_u3__abc_44466_n252_1), .Y(u0_u3__abc_44466_n253) );
  AND2X2 AND2X2_2518 ( .A(u0_u3__abc_44466_n254_1), .B(u0_u3__abc_44466_n251), .Y(u0_u3__abc_44466_n255_1) );
  AND2X2 AND2X2_2519 ( .A(u0_u3__abc_44466_n256_1), .B(u0_u3__abc_44466_n257), .Y(u0_u3_csc_5__FF_INPUT) );
  AND2X2 AND2X2_252 ( .A(spec_req_cs_3_bF_buf4), .B(u0_tms3_10_), .Y(u0__abc_49347_n1435_1) );
  AND2X2 AND2X2_2520 ( .A(u0_u3_init_req_we_FF_INPUT_bF_buf5), .B(\wb_data_i[6] ), .Y(u0_u3__abc_44466_n259) );
  AND2X2 AND2X2_2521 ( .A(u0_u3__abc_44466_n239_1_bF_buf3), .B(u0_csc3_6_), .Y(u0_u3__abc_44466_n260_1) );
  AND2X2 AND2X2_2522 ( .A(u0_u3__abc_44466_n261), .B(u0_u3__abc_44466_n205_1_bF_buf3), .Y(u0_u3_csc_6__FF_INPUT) );
  AND2X2 AND2X2_2523 ( .A(u0_u3_init_req_we_FF_INPUT_bF_buf4), .B(\wb_data_i[7] ), .Y(u0_u3__abc_44466_n263_1) );
  AND2X2 AND2X2_2524 ( .A(u0_u3__abc_44466_n239_1_bF_buf2), .B(u0_csc3_7_), .Y(u0_u3__abc_44466_n264_1) );
  AND2X2 AND2X2_2525 ( .A(u0_u3__abc_44466_n265_1), .B(u0_u3__abc_44466_n205_1_bF_buf2), .Y(u0_u3_csc_7__FF_INPUT) );
  AND2X2 AND2X2_2526 ( .A(u0_u3_init_req_we_FF_INPUT_bF_buf3), .B(\wb_data_i[8] ), .Y(u0_u3__abc_44466_n267_1) );
  AND2X2 AND2X2_2527 ( .A(u0_u3__abc_44466_n239_1_bF_buf1), .B(u0_csc3_8_), .Y(u0_u3__abc_44466_n268) );
  AND2X2 AND2X2_2528 ( .A(u0_u3__abc_44466_n269), .B(u0_u3__abc_44466_n205_1_bF_buf1), .Y(u0_u3_csc_8__FF_INPUT) );
  AND2X2 AND2X2_2529 ( .A(u0_u3_init_req_we_FF_INPUT_bF_buf2), .B(\wb_data_i[9] ), .Y(u0_u3__abc_44466_n271) );
  AND2X2 AND2X2_253 ( .A(u0__abc_49347_n1436), .B(u0__abc_49347_n1179_bF_buf1), .Y(u0__abc_49347_n1437) );
  AND2X2 AND2X2_2530 ( .A(u0_u3__abc_44466_n239_1_bF_buf0), .B(u0_csc3_9_), .Y(u0_u3__abc_44466_n272_1) );
  AND2X2 AND2X2_2531 ( .A(u0_u3__abc_44466_n273), .B(u0_u3__abc_44466_n205_1_bF_buf0), .Y(u0_u3_csc_9__FF_INPUT) );
  AND2X2 AND2X2_2532 ( .A(u0_u3_init_req_we_FF_INPUT_bF_buf1), .B(\wb_data_i[10] ), .Y(u0_u3__abc_44466_n275) );
  AND2X2 AND2X2_2533 ( .A(u0_u3__abc_44466_n239_1_bF_buf4), .B(u0_csc3_10_), .Y(u0_u3__abc_44466_n276) );
  AND2X2 AND2X2_2534 ( .A(u0_u3__abc_44466_n277), .B(u0_u3__abc_44466_n205_1_bF_buf4), .Y(u0_u3_csc_10__FF_INPUT) );
  AND2X2 AND2X2_2535 ( .A(u0_u3_init_req_we_FF_INPUT_bF_buf0), .B(\wb_data_i[11] ), .Y(u0_u3__abc_44466_n279) );
  AND2X2 AND2X2_2536 ( .A(u0_u3__abc_44466_n239_1_bF_buf3), .B(u0_csc3_11_), .Y(u0_u3__abc_44466_n280_1) );
  AND2X2 AND2X2_2537 ( .A(u0_u3__abc_44466_n281), .B(u0_u3__abc_44466_n205_1_bF_buf3), .Y(u0_u3_csc_11__FF_INPUT) );
  AND2X2 AND2X2_2538 ( .A(u0_u3_init_req_we_FF_INPUT_bF_buf5), .B(\wb_data_i[12] ), .Y(u0_u3__abc_44466_n283) );
  AND2X2 AND2X2_2539 ( .A(u0_u3__abc_44466_n239_1_bF_buf2), .B(u0_csc3_12_), .Y(u0_u3__abc_44466_n284) );
  AND2X2 AND2X2_254 ( .A(spec_req_cs_2_bF_buf4), .B(u0_tms2_10_), .Y(u0__abc_49347_n1438) );
  AND2X2 AND2X2_2540 ( .A(u0_u3__abc_44466_n285_1), .B(u0_u3__abc_44466_n205_1_bF_buf2), .Y(u0_u3_csc_12__FF_INPUT) );
  AND2X2 AND2X2_2541 ( .A(u0_u3_init_req_we_FF_INPUT_bF_buf4), .B(\wb_data_i[13] ), .Y(u0_u3__abc_44466_n287_1) );
  AND2X2 AND2X2_2542 ( .A(u0_u3__abc_44466_n239_1_bF_buf1), .B(u0_csc3_13_), .Y(u0_u3__abc_44466_n288) );
  AND2X2 AND2X2_2543 ( .A(u0_u3__abc_44466_n289_1), .B(u0_u3__abc_44466_n205_1_bF_buf1), .Y(u0_u3_csc_13__FF_INPUT) );
  AND2X2 AND2X2_2544 ( .A(u0_u3_init_req_we_FF_INPUT_bF_buf3), .B(\wb_data_i[14] ), .Y(u0_u3__abc_44466_n291_1) );
  AND2X2 AND2X2_2545 ( .A(u0_u3__abc_44466_n239_1_bF_buf0), .B(u0_csc3_14_), .Y(u0_u3__abc_44466_n292) );
  AND2X2 AND2X2_2546 ( .A(u0_u3__abc_44466_n293), .B(u0_u3__abc_44466_n205_1_bF_buf0), .Y(u0_u3_csc_14__FF_INPUT) );
  AND2X2 AND2X2_2547 ( .A(u0_u3_init_req_we_FF_INPUT_bF_buf2), .B(\wb_data_i[15] ), .Y(u0_u3__abc_44466_n295_1) );
  AND2X2 AND2X2_2548 ( .A(u0_u3__abc_44466_n239_1_bF_buf4), .B(u0_csc3_15_), .Y(u0_u3__abc_44466_n296) );
  AND2X2 AND2X2_2549 ( .A(u0_u3__abc_44466_n297_1), .B(u0_u3__abc_44466_n205_1_bF_buf4), .Y(u0_u3_csc_15__FF_INPUT) );
  AND2X2 AND2X2_255 ( .A(u0__abc_49347_n1439), .B(u0__abc_49347_n1178_1_bF_buf1), .Y(u0__abc_49347_n1440) );
  AND2X2 AND2X2_2550 ( .A(u0_u3_init_req_we_FF_INPUT_bF_buf1), .B(\wb_data_i[16] ), .Y(u0_u3__abc_44466_n299_1) );
  AND2X2 AND2X2_2551 ( .A(u0_u3__abc_44466_n239_1_bF_buf3), .B(u0_csc3_16_), .Y(u0_u3__abc_44466_n300) );
  AND2X2 AND2X2_2552 ( .A(u0_u3__abc_44466_n301_1), .B(u0_u3__abc_44466_n205_1_bF_buf3), .Y(u0_u3_csc_16__FF_INPUT) );
  AND2X2 AND2X2_2553 ( .A(u0_u3_init_req_we_FF_INPUT_bF_buf0), .B(\wb_data_i[17] ), .Y(u0_u3__abc_44466_n303) );
  AND2X2 AND2X2_2554 ( .A(u0_u3__abc_44466_n239_1_bF_buf2), .B(u0_csc3_17_), .Y(u0_u3__abc_44466_n304) );
  AND2X2 AND2X2_2555 ( .A(u0_u3__abc_44466_n305), .B(u0_u3__abc_44466_n205_1_bF_buf2), .Y(u0_u3_csc_17__FF_INPUT) );
  AND2X2 AND2X2_2556 ( .A(u0_u3_init_req_we_FF_INPUT_bF_buf5), .B(\wb_data_i[18] ), .Y(u0_u3__abc_44466_n307) );
  AND2X2 AND2X2_2557 ( .A(u0_u3__abc_44466_n239_1_bF_buf1), .B(u0_csc3_18_), .Y(u0_u3__abc_44466_n308_1) );
  AND2X2 AND2X2_2558 ( .A(u0_u3__abc_44466_n309), .B(u0_u3__abc_44466_n205_1_bF_buf1), .Y(u0_u3_csc_18__FF_INPUT) );
  AND2X2 AND2X2_2559 ( .A(u0_u3_init_req_we_FF_INPUT_bF_buf4), .B(\wb_data_i[19] ), .Y(u0_u3__abc_44466_n311) );
  AND2X2 AND2X2_256 ( .A(spec_req_cs_1_bF_buf4), .B(u0_tms1_10_), .Y(u0__abc_49347_n1441) );
  AND2X2 AND2X2_2560 ( .A(u0_u3__abc_44466_n239_1_bF_buf0), .B(u0_csc3_19_), .Y(u0_u3__abc_44466_n312) );
  AND2X2 AND2X2_2561 ( .A(u0_u3__abc_44466_n313), .B(u0_u3__abc_44466_n205_1_bF_buf0), .Y(u0_u3_csc_19__FF_INPUT) );
  AND2X2 AND2X2_2562 ( .A(u0_u3_init_req_we_FF_INPUT_bF_buf3), .B(\wb_data_i[20] ), .Y(u0_u3__abc_44466_n315) );
  AND2X2 AND2X2_2563 ( .A(u0_u3__abc_44466_n239_1_bF_buf4), .B(u0_csc3_20_), .Y(u0_u3__abc_44466_n316) );
  AND2X2 AND2X2_2564 ( .A(u0_u3__abc_44466_n317), .B(u0_u3__abc_44466_n205_1_bF_buf4), .Y(u0_u3_csc_20__FF_INPUT) );
  AND2X2 AND2X2_2565 ( .A(u0_u3_init_req_we_FF_INPUT_bF_buf2), .B(\wb_data_i[21] ), .Y(u0_u3__abc_44466_n319) );
  AND2X2 AND2X2_2566 ( .A(u0_u3__abc_44466_n239_1_bF_buf3), .B(u0_csc3_21_), .Y(u0_u3__abc_44466_n320) );
  AND2X2 AND2X2_2567 ( .A(u0_u3__abc_44466_n321), .B(u0_u3__abc_44466_n205_1_bF_buf3), .Y(u0_u3_csc_21__FF_INPUT) );
  AND2X2 AND2X2_2568 ( .A(u0_u3_init_req_we_FF_INPUT_bF_buf1), .B(\wb_data_i[22] ), .Y(u0_u3__abc_44466_n323) );
  AND2X2 AND2X2_2569 ( .A(u0_u3__abc_44466_n239_1_bF_buf2), .B(u0_csc3_22_), .Y(u0_u3__abc_44466_n324_1) );
  AND2X2 AND2X2_257 ( .A(u0__abc_49347_n1175_bF_buf2), .B(u0__abc_49347_n1444_1), .Y(u0__abc_49347_n1445) );
  AND2X2 AND2X2_2570 ( .A(u0_u3__abc_44466_n325), .B(u0_u3__abc_44466_n205_1_bF_buf2), .Y(u0_u3_csc_22__FF_INPUT) );
  AND2X2 AND2X2_2571 ( .A(u0_u3_init_req_we_FF_INPUT_bF_buf0), .B(\wb_data_i[23] ), .Y(u0_u3__abc_44466_n327_1) );
  AND2X2 AND2X2_2572 ( .A(u0_u3__abc_44466_n239_1_bF_buf1), .B(u0_csc3_23_), .Y(u0_u3__abc_44466_n328_1) );
  AND2X2 AND2X2_2573 ( .A(u0_u3__abc_44466_n329), .B(u0_u3__abc_44466_n205_1_bF_buf1), .Y(u0_u3_csc_23__FF_INPUT) );
  AND2X2 AND2X2_2574 ( .A(u0_u3_init_req_we_FF_INPUT_bF_buf5), .B(\wb_data_i[24] ), .Y(u0_u3__abc_44466_n331) );
  AND2X2 AND2X2_2575 ( .A(u0_u3__abc_44466_n239_1_bF_buf0), .B(u0_csc3_24_), .Y(u0_u3__abc_44466_n332) );
  AND2X2 AND2X2_2576 ( .A(u0_u3__abc_44466_n333), .B(u0_u3__abc_44466_n205_1_bF_buf0), .Y(u0_u3_csc_24__FF_INPUT) );
  AND2X2 AND2X2_2577 ( .A(u0_u3_init_req_we_FF_INPUT_bF_buf4), .B(\wb_data_i[25] ), .Y(u0_u3__abc_44466_n335) );
  AND2X2 AND2X2_2578 ( .A(u0_u3__abc_44466_n239_1_bF_buf4), .B(u0_csc3_25_), .Y(u0_u3__abc_44466_n336) );
  AND2X2 AND2X2_2579 ( .A(u0_u3__abc_44466_n337), .B(u0_u3__abc_44466_n205_1_bF_buf4), .Y(u0_u3_csc_25__FF_INPUT) );
  AND2X2 AND2X2_258 ( .A(u0__abc_49347_n1443_1), .B(u0__abc_49347_n1445), .Y(u0__abc_49347_n1446) );
  AND2X2 AND2X2_2580 ( .A(u0_u3_init_req_we_FF_INPUT_bF_buf3), .B(\wb_data_i[26] ), .Y(u0_u3__abc_44466_n339) );
  AND2X2 AND2X2_2581 ( .A(u0_u3__abc_44466_n239_1_bF_buf3), .B(u0_csc3_26_), .Y(u0_u3__abc_44466_n340) );
  AND2X2 AND2X2_2582 ( .A(u0_u3__abc_44466_n341), .B(u0_u3__abc_44466_n205_1_bF_buf3), .Y(u0_u3_csc_26__FF_INPUT) );
  AND2X2 AND2X2_2583 ( .A(u0_u3_init_req_we_FF_INPUT_bF_buf2), .B(\wb_data_i[27] ), .Y(u0_u3__abc_44466_n343) );
  AND2X2 AND2X2_2584 ( .A(u0_u3__abc_44466_n239_1_bF_buf2), .B(u0_csc3_27_), .Y(u0_u3__abc_44466_n344) );
  AND2X2 AND2X2_2585 ( .A(u0_u3__abc_44466_n345), .B(u0_u3__abc_44466_n205_1_bF_buf2), .Y(u0_u3_csc_27__FF_INPUT) );
  AND2X2 AND2X2_2586 ( .A(u0_u3_init_req_we_FF_INPUT_bF_buf1), .B(\wb_data_i[28] ), .Y(u0_u3__abc_44466_n347) );
  AND2X2 AND2X2_2587 ( .A(u0_u3__abc_44466_n239_1_bF_buf1), .B(u0_csc3_28_), .Y(u0_u3__abc_44466_n348) );
  AND2X2 AND2X2_2588 ( .A(u0_u3__abc_44466_n349), .B(u0_u3__abc_44466_n205_1_bF_buf1), .Y(u0_u3_csc_28__FF_INPUT) );
  AND2X2 AND2X2_2589 ( .A(u0_u3_init_req_we_FF_INPUT_bF_buf0), .B(\wb_data_i[29] ), .Y(u0_u3__abc_44466_n351) );
  AND2X2 AND2X2_259 ( .A(u0__abc_49347_n1176_1_bF_buf2), .B(sp_tms_11_), .Y(u0__abc_49347_n1448) );
  AND2X2 AND2X2_2590 ( .A(u0_u3__abc_44466_n239_1_bF_buf0), .B(u0_csc3_29_), .Y(u0_u3__abc_44466_n352) );
  AND2X2 AND2X2_2591 ( .A(u0_u3__abc_44466_n353), .B(u0_u3__abc_44466_n205_1_bF_buf0), .Y(u0_u3_csc_29__FF_INPUT) );
  AND2X2 AND2X2_2592 ( .A(u0_u3_init_req_we_FF_INPUT_bF_buf5), .B(\wb_data_i[30] ), .Y(u0_u3__abc_44466_n355) );
  AND2X2 AND2X2_2593 ( .A(u0_u3__abc_44466_n239_1_bF_buf4), .B(u0_csc3_30_), .Y(u0_u3__abc_44466_n356) );
  AND2X2 AND2X2_2594 ( .A(u0_u3__abc_44466_n357), .B(u0_u3__abc_44466_n205_1_bF_buf4), .Y(u0_u3_csc_30__FF_INPUT) );
  AND2X2 AND2X2_2595 ( .A(u0_u3_init_req_we_FF_INPUT_bF_buf4), .B(\wb_data_i[31] ), .Y(u0_u3__abc_44466_n359) );
  AND2X2 AND2X2_2596 ( .A(u0_u3__abc_44466_n239_1_bF_buf3), .B(u0_csc3_31_), .Y(u0_u3__abc_44466_n360) );
  AND2X2 AND2X2_2597 ( .A(u0_u3__abc_44466_n361), .B(u0_u3__abc_44466_n205_1_bF_buf3), .Y(u0_u3_csc_31__FF_INPUT) );
  AND2X2 AND2X2_2598 ( .A(u0_u3__abc_44466_n212_1), .B(u0_u3_addr_r_2_), .Y(u0_u3_lmr_req_we_FF_INPUT) );
  AND2X2 AND2X2_2599 ( .A(u0_u3__abc_44466_n364_bF_buf4), .B(u0_tms3_0_), .Y(u0_u3__abc_44466_n365) );
  AND2X2 AND2X2_26 ( .A(_abc_55805_n314), .B(_abc_55805_n315), .Y(tms_s_8_) );
  AND2X2 AND2X2_260 ( .A(spec_req_cs_5_bF_buf3), .B(u0_tms5_11_), .Y(u0__abc_49347_n1449) );
  AND2X2 AND2X2_2600 ( .A(u0_u3_lmr_req_we_FF_INPUT_bF_buf3), .B(\wb_data_i[0] ), .Y(u0_u3__abc_44466_n366) );
  AND2X2 AND2X2_2601 ( .A(u0_u3__abc_44466_n364_bF_buf3), .B(u0_tms3_1_), .Y(u0_u3__abc_44466_n369) );
  AND2X2 AND2X2_2602 ( .A(u0_u3_lmr_req_we_FF_INPUT_bF_buf2), .B(\wb_data_i[1] ), .Y(u0_u3__abc_44466_n370) );
  AND2X2 AND2X2_2603 ( .A(u0_u3__abc_44466_n364_bF_buf2), .B(u0_tms3_2_), .Y(u0_u3__abc_44466_n373) );
  AND2X2 AND2X2_2604 ( .A(u0_u3_lmr_req_we_FF_INPUT_bF_buf1), .B(\wb_data_i[2] ), .Y(u0_u3__abc_44466_n374) );
  AND2X2 AND2X2_2605 ( .A(u0_u3__abc_44466_n364_bF_buf1), .B(u0_tms3_3_), .Y(u0_u3__abc_44466_n377) );
  AND2X2 AND2X2_2606 ( .A(u0_u3_lmr_req_we_FF_INPUT_bF_buf0), .B(\wb_data_i[3] ), .Y(u0_u3__abc_44466_n378) );
  AND2X2 AND2X2_2607 ( .A(u0_u3__abc_44466_n364_bF_buf0), .B(u0_tms3_4_), .Y(u0_u3__abc_44466_n381) );
  AND2X2 AND2X2_2608 ( .A(u0_u3_lmr_req_we_FF_INPUT_bF_buf4), .B(\wb_data_i[4] ), .Y(u0_u3__abc_44466_n382) );
  AND2X2 AND2X2_2609 ( .A(u0_u3__abc_44466_n364_bF_buf4), .B(u0_tms3_5_), .Y(u0_u3__abc_44466_n385) );
  AND2X2 AND2X2_261 ( .A(u0__abc_49347_n1451), .B(u0__abc_49347_n1185_bF_buf0), .Y(u0__abc_49347_n1452_1) );
  AND2X2 AND2X2_2610 ( .A(u0_u3_lmr_req_we_FF_INPUT_bF_buf3), .B(\wb_data_i[5] ), .Y(u0_u3__abc_44466_n386) );
  AND2X2 AND2X2_2611 ( .A(u0_u3__abc_44466_n364_bF_buf3), .B(u0_tms3_6_), .Y(u0_u3__abc_44466_n389) );
  AND2X2 AND2X2_2612 ( .A(u0_u3_lmr_req_we_FF_INPUT_bF_buf2), .B(\wb_data_i[6] ), .Y(u0_u3__abc_44466_n390) );
  AND2X2 AND2X2_2613 ( .A(u0_u3__abc_44466_n364_bF_buf2), .B(u0_tms3_7_), .Y(u0_u3__abc_44466_n393) );
  AND2X2 AND2X2_2614 ( .A(u0_u3_lmr_req_we_FF_INPUT_bF_buf1), .B(\wb_data_i[7] ), .Y(u0_u3__abc_44466_n394) );
  AND2X2 AND2X2_2615 ( .A(u0_u3__abc_44466_n364_bF_buf1), .B(u0_tms3_8_), .Y(u0_u3__abc_44466_n397) );
  AND2X2 AND2X2_2616 ( .A(u0_u3_lmr_req_we_FF_INPUT_bF_buf0), .B(\wb_data_i[8] ), .Y(u0_u3__abc_44466_n398) );
  AND2X2 AND2X2_2617 ( .A(u0_u3__abc_44466_n364_bF_buf0), .B(u0_tms3_9_), .Y(u0_u3__abc_44466_n401) );
  AND2X2 AND2X2_2618 ( .A(u0_u3_lmr_req_we_FF_INPUT_bF_buf4), .B(\wb_data_i[9] ), .Y(u0_u3__abc_44466_n402) );
  AND2X2 AND2X2_2619 ( .A(u0_u3__abc_44466_n364_bF_buf4), .B(u0_tms3_10_), .Y(u0_u3__abc_44466_n405) );
  AND2X2 AND2X2_262 ( .A(u0__abc_49347_n1452_1), .B(u0__abc_49347_n1450), .Y(u0__abc_49347_n1453_1) );
  AND2X2 AND2X2_2620 ( .A(u0_u3_lmr_req_we_FF_INPUT_bF_buf3), .B(\wb_data_i[10] ), .Y(u0_u3__abc_44466_n406) );
  AND2X2 AND2X2_2621 ( .A(u0_u3__abc_44466_n364_bF_buf3), .B(u0_tms3_11_), .Y(u0_u3__abc_44466_n409) );
  AND2X2 AND2X2_2622 ( .A(u0_u3_lmr_req_we_FF_INPUT_bF_buf2), .B(\wb_data_i[11] ), .Y(u0_u3__abc_44466_n410) );
  AND2X2 AND2X2_2623 ( .A(u0_u3__abc_44466_n364_bF_buf2), .B(u0_tms3_12_), .Y(u0_u3__abc_44466_n413) );
  AND2X2 AND2X2_2624 ( .A(u0_u3_lmr_req_we_FF_INPUT_bF_buf1), .B(\wb_data_i[12] ), .Y(u0_u3__abc_44466_n414) );
  AND2X2 AND2X2_2625 ( .A(u0_u3__abc_44466_n364_bF_buf1), .B(u0_tms3_13_), .Y(u0_u3__abc_44466_n417) );
  AND2X2 AND2X2_2626 ( .A(u0_u3_lmr_req_we_FF_INPUT_bF_buf0), .B(\wb_data_i[13] ), .Y(u0_u3__abc_44466_n418) );
  AND2X2 AND2X2_2627 ( .A(u0_u3__abc_44466_n364_bF_buf0), .B(u0_tms3_14_), .Y(u0_u3__abc_44466_n421) );
  AND2X2 AND2X2_2628 ( .A(u0_u3_lmr_req_we_FF_INPUT_bF_buf4), .B(\wb_data_i[14] ), .Y(u0_u3__abc_44466_n422) );
  AND2X2 AND2X2_2629 ( .A(u0_u3__abc_44466_n364_bF_buf4), .B(u0_tms3_15_), .Y(u0_u3__abc_44466_n425) );
  AND2X2 AND2X2_263 ( .A(u0__abc_49347_n1454), .B(u0__abc_49347_n1181_bF_buf0), .Y(u0__abc_49347_n1455) );
  AND2X2 AND2X2_2630 ( .A(u0_u3_lmr_req_we_FF_INPUT_bF_buf3), .B(\wb_data_i[15] ), .Y(u0_u3__abc_44466_n426) );
  AND2X2 AND2X2_2631 ( .A(u0_u3__abc_44466_n364_bF_buf3), .B(u0_tms3_16_), .Y(u0_u3__abc_44466_n429) );
  AND2X2 AND2X2_2632 ( .A(u0_u3_lmr_req_we_FF_INPUT_bF_buf2), .B(\wb_data_i[16] ), .Y(u0_u3__abc_44466_n430) );
  AND2X2 AND2X2_2633 ( .A(u0_u3__abc_44466_n364_bF_buf2), .B(u0_tms3_17_), .Y(u0_u3__abc_44466_n433) );
  AND2X2 AND2X2_2634 ( .A(u0_u3_lmr_req_we_FF_INPUT_bF_buf1), .B(\wb_data_i[17] ), .Y(u0_u3__abc_44466_n434) );
  AND2X2 AND2X2_2635 ( .A(u0_u3__abc_44466_n364_bF_buf1), .B(u0_tms3_18_), .Y(u0_u3__abc_44466_n437) );
  AND2X2 AND2X2_2636 ( .A(u0_u3_lmr_req_we_FF_INPUT_bF_buf0), .B(\wb_data_i[18] ), .Y(u0_u3__abc_44466_n438) );
  AND2X2 AND2X2_2637 ( .A(u0_u3__abc_44466_n364_bF_buf0), .B(u0_tms3_19_), .Y(u0_u3__abc_44466_n441) );
  AND2X2 AND2X2_2638 ( .A(u0_u3_lmr_req_we_FF_INPUT_bF_buf4), .B(\wb_data_i[19] ), .Y(u0_u3__abc_44466_n442) );
  AND2X2 AND2X2_2639 ( .A(u0_u3__abc_44466_n364_bF_buf4), .B(u0_tms3_20_), .Y(u0_u3__abc_44466_n445) );
  AND2X2 AND2X2_264 ( .A(spec_req_cs_4_bF_buf3), .B(u0_tms4_11_), .Y(u0__abc_49347_n1456) );
  AND2X2 AND2X2_2640 ( .A(u0_u3_lmr_req_we_FF_INPUT_bF_buf3), .B(\wb_data_i[20] ), .Y(u0_u3__abc_44466_n446) );
  AND2X2 AND2X2_2641 ( .A(u0_u3__abc_44466_n364_bF_buf3), .B(u0_tms3_21_), .Y(u0_u3__abc_44466_n449) );
  AND2X2 AND2X2_2642 ( .A(u0_u3_lmr_req_we_FF_INPUT_bF_buf2), .B(\wb_data_i[21] ), .Y(u0_u3__abc_44466_n450) );
  AND2X2 AND2X2_2643 ( .A(u0_u3__abc_44466_n364_bF_buf2), .B(u0_tms3_22_), .Y(u0_u3__abc_44466_n453) );
  AND2X2 AND2X2_2644 ( .A(u0_u3_lmr_req_we_FF_INPUT_bF_buf1), .B(\wb_data_i[22] ), .Y(u0_u3__abc_44466_n454) );
  AND2X2 AND2X2_2645 ( .A(u0_u3__abc_44466_n364_bF_buf1), .B(u0_tms3_23_), .Y(u0_u3__abc_44466_n457) );
  AND2X2 AND2X2_2646 ( .A(u0_u3_lmr_req_we_FF_INPUT_bF_buf0), .B(\wb_data_i[23] ), .Y(u0_u3__abc_44466_n458) );
  AND2X2 AND2X2_2647 ( .A(u0_u3__abc_44466_n364_bF_buf0), .B(u0_tms3_24_), .Y(u0_u3__abc_44466_n461) );
  AND2X2 AND2X2_2648 ( .A(u0_u3_lmr_req_we_FF_INPUT_bF_buf4), .B(\wb_data_i[24] ), .Y(u0_u3__abc_44466_n462) );
  AND2X2 AND2X2_2649 ( .A(u0_u3__abc_44466_n364_bF_buf4), .B(u0_tms3_25_), .Y(u0_u3__abc_44466_n465) );
  AND2X2 AND2X2_265 ( .A(u0__abc_49347_n1457), .B(u0__abc_49347_n1180_1_bF_buf0), .Y(u0__abc_49347_n1458) );
  AND2X2 AND2X2_2650 ( .A(u0_u3_lmr_req_we_FF_INPUT_bF_buf3), .B(\wb_data_i[25] ), .Y(u0_u3__abc_44466_n466) );
  AND2X2 AND2X2_2651 ( .A(u0_u3__abc_44466_n364_bF_buf3), .B(u0_tms3_26_), .Y(u0_u3__abc_44466_n469) );
  AND2X2 AND2X2_2652 ( .A(u0_u3_lmr_req_we_FF_INPUT_bF_buf2), .B(\wb_data_i[26] ), .Y(u0_u3__abc_44466_n470) );
  AND2X2 AND2X2_2653 ( .A(u0_u3__abc_44466_n364_bF_buf2), .B(u0_tms3_27_), .Y(u0_u3__abc_44466_n473) );
  AND2X2 AND2X2_2654 ( .A(u0_u3_lmr_req_we_FF_INPUT_bF_buf1), .B(\wb_data_i[27] ), .Y(u0_u3__abc_44466_n474) );
  AND2X2 AND2X2_2655 ( .A(u0_u3__abc_44466_n364_bF_buf1), .B(u0_tms3_28_), .Y(u0_u3__abc_44466_n477) );
  AND2X2 AND2X2_2656 ( .A(u0_u3_lmr_req_we_FF_INPUT_bF_buf0), .B(\wb_data_i[28] ), .Y(u0_u3__abc_44466_n478) );
  AND2X2 AND2X2_2657 ( .A(u0_u3__abc_44466_n364_bF_buf0), .B(u0_tms3_29_), .Y(u0_u3__abc_44466_n481) );
  AND2X2 AND2X2_2658 ( .A(u0_u3_lmr_req_we_FF_INPUT_bF_buf4), .B(\wb_data_i[29] ), .Y(u0_u3__abc_44466_n482) );
  AND2X2 AND2X2_2659 ( .A(u0_u3__abc_44466_n364_bF_buf4), .B(u0_tms3_30_), .Y(u0_u3__abc_44466_n485) );
  AND2X2 AND2X2_266 ( .A(spec_req_cs_3_bF_buf3), .B(u0_tms3_11_), .Y(u0__abc_49347_n1459) );
  AND2X2 AND2X2_2660 ( .A(u0_u3_lmr_req_we_FF_INPUT_bF_buf3), .B(\wb_data_i[30] ), .Y(u0_u3__abc_44466_n486) );
  AND2X2 AND2X2_2661 ( .A(u0_u3__abc_44466_n364_bF_buf3), .B(u0_tms3_31_), .Y(u0_u3__abc_44466_n489) );
  AND2X2 AND2X2_2662 ( .A(u0_u3_lmr_req_we_FF_INPUT_bF_buf2), .B(\wb_data_i[31] ), .Y(u0_u3__abc_44466_n490) );
  AND2X2 AND2X2_2663 ( .A(u0_u3__abc_44466_n495), .B(u0_u3_lmr_req_we), .Y(u0_u3__abc_44466_n496) );
  AND2X2 AND2X2_2664 ( .A(u0_u3__abc_44466_n496), .B(u0_u3_inited), .Y(u0_u3__abc_44466_n497) );
  AND2X2 AND2X2_2665 ( .A(u0_u3__abc_44466_n499), .B(u0_lmr_req3), .Y(u0_u3__abc_44466_n500) );
  AND2X2 AND2X2_2666 ( .A(u0_u3__abc_44466_n498), .B(u0_u3__abc_44466_n500), .Y(u0_u3__abc_44466_n501) );
  AND2X2 AND2X2_2667 ( .A(u0_u3__abc_44466_n503), .B(u0_init_req3), .Y(u0_u3__abc_44466_n504) );
  AND2X2 AND2X2_2668 ( .A(u0_u3__abc_44466_n505), .B(u0_csc3_0_), .Y(u0_u3__abc_44466_n506) );
  AND2X2 AND2X2_2669 ( .A(u0_u3__abc_44466_n506), .B(u0_u3_init_req_we), .Y(u0_u3__abc_44466_n507) );
  AND2X2 AND2X2_267 ( .A(u0__abc_49347_n1460), .B(u0__abc_49347_n1179_bF_buf0), .Y(u0__abc_49347_n1461_1) );
  AND2X2 AND2X2_2670 ( .A(u0_u3__abc_44466_n495), .B(u0_u3__abc_44466_n507), .Y(u0_u3__abc_44466_n508) );
  AND2X2 AND2X2_2671 ( .A(u0_csc3_8_), .B(wb_we_i), .Y(u0_u3__abc_44466_n511) );
  AND2X2 AND2X2_2672 ( .A(u0_csc3_20_), .B(u0_csc_mask_4_), .Y(u0_u3__abc_44466_n512) );
  AND2X2 AND2X2_2673 ( .A(u0_csc_mask_4_), .B(wb_addr_i_25_bF_buf1), .Y(u0_u3__abc_44466_n513) );
  AND2X2 AND2X2_2674 ( .A(u0_csc_mask_3_), .B(\wb_addr_i[24] ), .Y(u0_u3__abc_44466_n516) );
  AND2X2 AND2X2_2675 ( .A(u0_csc3_19_), .B(u0_csc_mask_3_), .Y(u0_u3__abc_44466_n517) );
  AND2X2 AND2X2_2676 ( .A(u0_u3__abc_44466_n515), .B(u0_u3__abc_44466_n519), .Y(u0_u3__abc_44466_n520) );
  AND2X2 AND2X2_2677 ( .A(u0_csc3_18_), .B(u0_csc_mask_2_), .Y(u0_u3__abc_44466_n522) );
  AND2X2 AND2X2_2678 ( .A(u0_u3__abc_44466_n522), .B(u0_u3__abc_44466_n521), .Y(u0_u3__abc_44466_n523) );
  AND2X2 AND2X2_2679 ( .A(u0_u3__abc_44466_n526), .B(u0_u3__abc_44466_n524), .Y(u0_u3__abc_44466_n527) );
  AND2X2 AND2X2_268 ( .A(spec_req_cs_2_bF_buf3), .B(u0_tms2_11_), .Y(u0__abc_49347_n1462_1) );
  AND2X2 AND2X2_2680 ( .A(u0_u3__abc_44466_n520), .B(u0_u3__abc_44466_n527), .Y(u0_u3__abc_44466_n528) );
  AND2X2 AND2X2_2681 ( .A(u0_csc3_22_), .B(u0_csc_mask_6_), .Y(u0_u3__abc_44466_n529) );
  AND2X2 AND2X2_2682 ( .A(u0_csc_mask_6_), .B(\wb_addr_i[27] ), .Y(u0_u3__abc_44466_n530) );
  AND2X2 AND2X2_2683 ( .A(u0_csc_mask_5_), .B(\wb_addr_i[26] ), .Y(u0_u3__abc_44466_n533) );
  AND2X2 AND2X2_2684 ( .A(u0_csc3_21_), .B(u0_csc_mask_5_), .Y(u0_u3__abc_44466_n534) );
  AND2X2 AND2X2_2685 ( .A(u0_u3__abc_44466_n532), .B(u0_u3__abc_44466_n536), .Y(u0_u3__abc_44466_n537) );
  AND2X2 AND2X2_2686 ( .A(u0_u3__abc_44466_n512), .B(u0_u3__abc_44466_n538), .Y(u0_u3__abc_44466_n539) );
  AND2X2 AND2X2_2687 ( .A(u0_u3__abc_44466_n542), .B(u0_u3__abc_44466_n540), .Y(u0_u3__abc_44466_n543) );
  AND2X2 AND2X2_2688 ( .A(u0_u3__abc_44466_n537), .B(u0_u3__abc_44466_n543), .Y(u0_u3__abc_44466_n544) );
  AND2X2 AND2X2_2689 ( .A(u0_u3__abc_44466_n528), .B(u0_u3__abc_44466_n544), .Y(u0_u3__abc_44466_n545) );
  AND2X2 AND2X2_269 ( .A(u0__abc_49347_n1463), .B(u0__abc_49347_n1178_1_bF_buf0), .Y(u0__abc_49347_n1464) );
  AND2X2 AND2X2_2690 ( .A(u0_u3__abc_44466_n531), .B(u0_u3__abc_44466_n529), .Y(u0_u3__abc_44466_n546) );
  AND2X2 AND2X2_2691 ( .A(u0_csc_mask_7_), .B(\wb_addr_i[28] ), .Y(u0_u3__abc_44466_n548) );
  AND2X2 AND2X2_2692 ( .A(u0_csc3_23_), .B(u0_csc_mask_7_), .Y(u0_u3__abc_44466_n550) );
  AND2X2 AND2X2_2693 ( .A(u0_u3__abc_44466_n547), .B(u0_u3__abc_44466_n551), .Y(u0_u3__abc_44466_n552) );
  AND2X2 AND2X2_2694 ( .A(u0_u3__abc_44466_n552), .B(u0_u3__abc_44466_n554), .Y(u0_u3__abc_44466_n555) );
  AND2X2 AND2X2_2695 ( .A(u0_u3__abc_44466_n545), .B(u0_u3__abc_44466_n555), .Y(u0_u3__abc_44466_n556) );
  AND2X2 AND2X2_2696 ( .A(u0_csc_mask_2_), .B(wb_addr_i_23_bF_buf0), .Y(u0_u3__abc_44466_n557) );
  AND2X2 AND2X2_2697 ( .A(u0_csc_mask_1_), .B(\wb_addr_i[22] ), .Y(u0_u3__abc_44466_n560) );
  AND2X2 AND2X2_2698 ( .A(u0_csc3_17_), .B(u0_csc_mask_1_), .Y(u0_u3__abc_44466_n561) );
  AND2X2 AND2X2_2699 ( .A(u0_u3__abc_44466_n559), .B(u0_u3__abc_44466_n563), .Y(u0_u3__abc_44466_n564) );
  AND2X2 AND2X2_27 ( .A(_abc_55805_n317), .B(_abc_55805_n318), .Y(tms_s_9_) );
  AND2X2 AND2X2_270 ( .A(spec_req_cs_1_bF_buf3), .B(u0_tms1_11_), .Y(u0__abc_49347_n1465) );
  AND2X2 AND2X2_2700 ( .A(u0_csc_mask_0_), .B(\wb_addr_i[21] ), .Y(u0_u3__abc_44466_n565) );
  AND2X2 AND2X2_2701 ( .A(u0_csc3_16_), .B(u0_csc_mask_0_), .Y(u0_u3__abc_44466_n566) );
  AND2X2 AND2X2_2702 ( .A(u0_u3__abc_44466_n568), .B(u0_u3__abc_44466_n570), .Y(u0_u3__abc_44466_n571) );
  AND2X2 AND2X2_2703 ( .A(u0_u3__abc_44466_n564), .B(u0_u3__abc_44466_n571), .Y(u0_u3__abc_44466_n572) );
  AND2X2 AND2X2_2704 ( .A(u0_u3__abc_44466_n574), .B(u0_csc3_0_), .Y(u0_u3__abc_44466_n575) );
  AND2X2 AND2X2_2705 ( .A(u0_u3__abc_44466_n572), .B(u0_u3__abc_44466_n575), .Y(u0_u3__abc_44466_n576) );
  AND2X2 AND2X2_2706 ( .A(u0_u3__abc_44466_n556), .B(u0_u3__abc_44466_n576), .Y(u0_u3__abc_44466_n577) );
  AND2X2 AND2X2_2707 ( .A(u0_u3__abc_44466_n577), .B(u0_u3__abc_44466_n511), .Y(u0_u3_wp_err) );
  AND2X2 AND2X2_2708 ( .A(u0_u3__abc_44466_n577), .B(u0_u3__abc_44466_n579), .Y(u0_cs3) );
  AND2X2 AND2X2_2709 ( .A(u0_u4__abc_44844_n201_1), .B(u0_u4__abc_44844_n202), .Y(u0_u4__abc_44844_n203_1) );
  AND2X2 AND2X2_271 ( .A(u0__abc_49347_n1175_bF_buf1), .B(u0__abc_49347_n1468), .Y(u0__abc_49347_n1469) );
  AND2X2 AND2X2_2710 ( .A(u0_u4_addr_r_5_), .B(u0_u4_addr_r_4_), .Y(u0_u4__abc_44844_n204_1) );
  AND2X2 AND2X2_2711 ( .A(u0_u4__abc_44844_n204_1), .B(u0_rf_we), .Y(u0_u4__abc_44844_n205) );
  AND2X2 AND2X2_2712 ( .A(u0_u4__abc_44844_n205), .B(u0_u4__abc_44844_n203_1), .Y(u0_u4__abc_44844_n206_1) );
  AND2X2 AND2X2_2713 ( .A(u0_u4__abc_44844_n206_1), .B(u0_u4_addr_r_2_), .Y(u0_u4_lmr_req_we_FF_INPUT) );
  AND2X2 AND2X2_2714 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf6), .B(u0_u4__abc_44844_n210_1), .Y(u0_u4__abc_44844_n211) );
  AND2X2 AND2X2_2715 ( .A(u0_u4__abc_44844_n212_1), .B(u0_u4__abc_44844_n209_1_bF_buf7), .Y(u0_u4__abc_44844_n213_1) );
  AND2X2 AND2X2_2716 ( .A(u0_u4__abc_44844_n213_1), .B(u0_u4__abc_44844_n208), .Y(u0_u4_tms_0__FF_INPUT) );
  AND2X2 AND2X2_2717 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf4), .B(u0_u4__abc_44844_n216_1), .Y(u0_u4__abc_44844_n217) );
  AND2X2 AND2X2_2718 ( .A(u0_u4__abc_44844_n218_1), .B(u0_u4__abc_44844_n209_1_bF_buf6), .Y(u0_u4__abc_44844_n219_1) );
  AND2X2 AND2X2_2719 ( .A(u0_u4__abc_44844_n219_1), .B(u0_u4__abc_44844_n215_1), .Y(u0_u4_tms_1__FF_INPUT) );
  AND2X2 AND2X2_272 ( .A(u0__abc_49347_n1467), .B(u0__abc_49347_n1469), .Y(u0__abc_49347_n1470_1) );
  AND2X2 AND2X2_2720 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf2), .B(u0_u4__abc_44844_n222_1), .Y(u0_u4__abc_44844_n223) );
  AND2X2 AND2X2_2721 ( .A(u0_u4__abc_44844_n224_1), .B(u0_u4__abc_44844_n209_1_bF_buf5), .Y(u0_u4__abc_44844_n225_1) );
  AND2X2 AND2X2_2722 ( .A(u0_u4__abc_44844_n225_1), .B(u0_u4__abc_44844_n221_1), .Y(u0_u4_tms_2__FF_INPUT) );
  AND2X2 AND2X2_2723 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf0), .B(u0_u4__abc_44844_n228_1), .Y(u0_u4__abc_44844_n229) );
  AND2X2 AND2X2_2724 ( .A(u0_u4__abc_44844_n230_1), .B(u0_u4__abc_44844_n209_1_bF_buf4), .Y(u0_u4__abc_44844_n231_1) );
  AND2X2 AND2X2_2725 ( .A(u0_u4__abc_44844_n231_1), .B(u0_u4__abc_44844_n227_1), .Y(u0_u4_tms_3__FF_INPUT) );
  AND2X2 AND2X2_2726 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf6), .B(u0_u4__abc_44844_n234_1), .Y(u0_u4__abc_44844_n235) );
  AND2X2 AND2X2_2727 ( .A(u0_u4__abc_44844_n236_1), .B(u0_u4__abc_44844_n209_1_bF_buf3), .Y(u0_u4__abc_44844_n237_1) );
  AND2X2 AND2X2_2728 ( .A(u0_u4__abc_44844_n237_1), .B(u0_u4__abc_44844_n233_1), .Y(u0_u4_tms_4__FF_INPUT) );
  AND2X2 AND2X2_2729 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf4), .B(u0_u4__abc_44844_n240_1), .Y(u0_u4__abc_44844_n241) );
  AND2X2 AND2X2_273 ( .A(u0__abc_49347_n1176_1_bF_buf1), .B(sp_tms_12_), .Y(u0__abc_49347_n1472) );
  AND2X2 AND2X2_2730 ( .A(u0_u4__abc_44844_n242_1), .B(u0_u4__abc_44844_n209_1_bF_buf2), .Y(u0_u4__abc_44844_n243_1) );
  AND2X2 AND2X2_2731 ( .A(u0_u4__abc_44844_n243_1), .B(u0_u4__abc_44844_n239_1), .Y(u0_u4_tms_5__FF_INPUT) );
  AND2X2 AND2X2_2732 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf2), .B(u0_u4__abc_44844_n246_1), .Y(u0_u4__abc_44844_n247) );
  AND2X2 AND2X2_2733 ( .A(u0_u4__abc_44844_n248_1), .B(u0_u4__abc_44844_n209_1_bF_buf1), .Y(u0_u4__abc_44844_n249_1) );
  AND2X2 AND2X2_2734 ( .A(u0_u4__abc_44844_n249_1), .B(u0_u4__abc_44844_n245_1), .Y(u0_u4_tms_6__FF_INPUT) );
  AND2X2 AND2X2_2735 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf0), .B(u0_u4__abc_44844_n252_1), .Y(u0_u4__abc_44844_n253) );
  AND2X2 AND2X2_2736 ( .A(u0_u4__abc_44844_n254), .B(u0_u4__abc_44844_n209_1_bF_buf0), .Y(u0_u4__abc_44844_n255) );
  AND2X2 AND2X2_2737 ( .A(u0_u4__abc_44844_n255), .B(u0_u4__abc_44844_n251_1), .Y(u0_u4_tms_7__FF_INPUT) );
  AND2X2 AND2X2_2738 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf6), .B(u0_u4__abc_44844_n258_1), .Y(u0_u4__abc_44844_n259_1) );
  AND2X2 AND2X2_2739 ( .A(u0_u4__abc_44844_n260_1), .B(u0_u4__abc_44844_n209_1_bF_buf7), .Y(u0_u4__abc_44844_n261_1) );
  AND2X2 AND2X2_274 ( .A(spec_req_cs_5_bF_buf2), .B(u0_tms5_12_), .Y(u0__abc_49347_n1473) );
  AND2X2 AND2X2_2740 ( .A(u0_u4__abc_44844_n261_1), .B(u0_u4__abc_44844_n257), .Y(u0_u4_tms_8__FF_INPUT) );
  AND2X2 AND2X2_2741 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf4), .B(u0_u4__abc_44844_n264), .Y(u0_u4__abc_44844_n265) );
  AND2X2 AND2X2_2742 ( .A(u0_u4__abc_44844_n266), .B(u0_u4__abc_44844_n209_1_bF_buf6), .Y(u0_u4__abc_44844_n267) );
  AND2X2 AND2X2_2743 ( .A(u0_u4__abc_44844_n267), .B(u0_u4__abc_44844_n263_1), .Y(u0_u4_tms_9__FF_INPUT) );
  AND2X2 AND2X2_2744 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf2), .B(u0_u4__abc_44844_n270_1), .Y(u0_u4__abc_44844_n271) );
  AND2X2 AND2X2_2745 ( .A(u0_u4__abc_44844_n272), .B(u0_u4__abc_44844_n209_1_bF_buf5), .Y(u0_u4__abc_44844_n273) );
  AND2X2 AND2X2_2746 ( .A(u0_u4__abc_44844_n273), .B(u0_u4__abc_44844_n269), .Y(u0_u4_tms_10__FF_INPUT) );
  AND2X2 AND2X2_2747 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf0), .B(u0_u4__abc_44844_n276_1), .Y(u0_u4__abc_44844_n277) );
  AND2X2 AND2X2_2748 ( .A(u0_u4__abc_44844_n278), .B(u0_u4__abc_44844_n209_1_bF_buf4), .Y(u0_u4__abc_44844_n279) );
  AND2X2 AND2X2_2749 ( .A(u0_u4__abc_44844_n279), .B(u0_u4__abc_44844_n275), .Y(u0_u4_tms_11__FF_INPUT) );
  AND2X2 AND2X2_275 ( .A(u0__abc_49347_n1475), .B(u0__abc_49347_n1185_bF_buf5), .Y(u0__abc_49347_n1476) );
  AND2X2 AND2X2_2750 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf6), .B(u0_u4__abc_44844_n282), .Y(u0_u4__abc_44844_n283_1) );
  AND2X2 AND2X2_2751 ( .A(u0_u4__abc_44844_n284), .B(u0_u4__abc_44844_n209_1_bF_buf3), .Y(u0_u4__abc_44844_n285_1) );
  AND2X2 AND2X2_2752 ( .A(u0_u4__abc_44844_n285_1), .B(u0_u4__abc_44844_n281_1), .Y(u0_u4_tms_12__FF_INPUT) );
  AND2X2 AND2X2_2753 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf4), .B(u0_u4__abc_44844_n288), .Y(u0_u4__abc_44844_n289) );
  AND2X2 AND2X2_2754 ( .A(u0_u4__abc_44844_n290), .B(u0_u4__abc_44844_n209_1_bF_buf2), .Y(u0_u4__abc_44844_n291_1) );
  AND2X2 AND2X2_2755 ( .A(u0_u4__abc_44844_n291_1), .B(u0_u4__abc_44844_n287_1), .Y(u0_u4_tms_13__FF_INPUT) );
  AND2X2 AND2X2_2756 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf2), .B(u0_u4__abc_44844_n294), .Y(u0_u4__abc_44844_n295_1) );
  AND2X2 AND2X2_2757 ( .A(u0_u4__abc_44844_n296), .B(u0_u4__abc_44844_n209_1_bF_buf1), .Y(u0_u4__abc_44844_n297_1) );
  AND2X2 AND2X2_2758 ( .A(u0_u4__abc_44844_n297_1), .B(u0_u4__abc_44844_n293_1), .Y(u0_u4_tms_14__FF_INPUT) );
  AND2X2 AND2X2_2759 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf0), .B(u0_u4__abc_44844_n300), .Y(u0_u4__abc_44844_n301) );
  AND2X2 AND2X2_276 ( .A(u0__abc_49347_n1476), .B(u0__abc_49347_n1474), .Y(u0__abc_49347_n1477) );
  AND2X2 AND2X2_2760 ( .A(u0_u4__abc_44844_n302), .B(u0_u4__abc_44844_n209_1_bF_buf0), .Y(u0_u4__abc_44844_n303) );
  AND2X2 AND2X2_2761 ( .A(u0_u4__abc_44844_n303), .B(u0_u4__abc_44844_n299), .Y(u0_u4_tms_15__FF_INPUT) );
  AND2X2 AND2X2_2762 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf6), .B(u0_u4__abc_44844_n306_1), .Y(u0_u4__abc_44844_n307) );
  AND2X2 AND2X2_2763 ( .A(u0_u4__abc_44844_n308), .B(u0_u4__abc_44844_n209_1_bF_buf7), .Y(u0_u4__abc_44844_n309) );
  AND2X2 AND2X2_2764 ( .A(u0_u4__abc_44844_n309), .B(u0_u4__abc_44844_n305), .Y(u0_u4_tms_16__FF_INPUT) );
  AND2X2 AND2X2_2765 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf4), .B(u0_u4__abc_44844_n312), .Y(u0_u4__abc_44844_n313) );
  AND2X2 AND2X2_2766 ( .A(u0_u4__abc_44844_n314), .B(u0_u4__abc_44844_n209_1_bF_buf6), .Y(u0_u4__abc_44844_n315) );
  AND2X2 AND2X2_2767 ( .A(u0_u4__abc_44844_n315), .B(u0_u4__abc_44844_n311), .Y(u0_u4_tms_17__FF_INPUT) );
  AND2X2 AND2X2_2768 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf2), .B(u0_u4__abc_44844_n318_1), .Y(u0_u4__abc_44844_n319) );
  AND2X2 AND2X2_2769 ( .A(u0_u4__abc_44844_n320_1), .B(u0_u4__abc_44844_n209_1_bF_buf5), .Y(u0_u4__abc_44844_n321) );
  AND2X2 AND2X2_277 ( .A(u0__abc_49347_n1478), .B(u0__abc_49347_n1181_bF_buf5), .Y(u0__abc_49347_n1479_1) );
  AND2X2 AND2X2_2770 ( .A(u0_u4__abc_44844_n321), .B(u0_u4__abc_44844_n317), .Y(u0_u4_tms_18__FF_INPUT) );
  AND2X2 AND2X2_2771 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf0), .B(u0_u4__abc_44844_n324_1), .Y(u0_u4__abc_44844_n325) );
  AND2X2 AND2X2_2772 ( .A(u0_u4__abc_44844_n326), .B(u0_u4__abc_44844_n209_1_bF_buf4), .Y(u0_u4__abc_44844_n327) );
  AND2X2 AND2X2_2773 ( .A(u0_u4__abc_44844_n327), .B(u0_u4__abc_44844_n323_1), .Y(u0_u4_tms_19__FF_INPUT) );
  AND2X2 AND2X2_2774 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf6), .B(u0_u4__abc_44844_n330), .Y(u0_u4__abc_44844_n331) );
  AND2X2 AND2X2_2775 ( .A(u0_u4__abc_44844_n332), .B(u0_u4__abc_44844_n209_1_bF_buf3), .Y(u0_u4__abc_44844_n333) );
  AND2X2 AND2X2_2776 ( .A(u0_u4__abc_44844_n333), .B(u0_u4__abc_44844_n329), .Y(u0_u4_tms_20__FF_INPUT) );
  AND2X2 AND2X2_2777 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf4), .B(u0_u4__abc_44844_n336), .Y(u0_u4__abc_44844_n337) );
  AND2X2 AND2X2_2778 ( .A(u0_u4__abc_44844_n338), .B(u0_u4__abc_44844_n209_1_bF_buf2), .Y(u0_u4__abc_44844_n339) );
  AND2X2 AND2X2_2779 ( .A(u0_u4__abc_44844_n339), .B(u0_u4__abc_44844_n335), .Y(u0_u4_tms_21__FF_INPUT) );
  AND2X2 AND2X2_278 ( .A(spec_req_cs_4_bF_buf2), .B(u0_tms4_12_), .Y(u0__abc_49347_n1480_1) );
  AND2X2 AND2X2_2780 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf2), .B(u0_u4__abc_44844_n342), .Y(u0_u4__abc_44844_n343) );
  AND2X2 AND2X2_2781 ( .A(u0_u4__abc_44844_n344), .B(u0_u4__abc_44844_n209_1_bF_buf1), .Y(u0_u4__abc_44844_n345) );
  AND2X2 AND2X2_2782 ( .A(u0_u4__abc_44844_n345), .B(u0_u4__abc_44844_n341), .Y(u0_u4_tms_22__FF_INPUT) );
  AND2X2 AND2X2_2783 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf0), .B(u0_u4__abc_44844_n348), .Y(u0_u4__abc_44844_n349) );
  AND2X2 AND2X2_2784 ( .A(u0_u4__abc_44844_n350), .B(u0_u4__abc_44844_n209_1_bF_buf0), .Y(u0_u4__abc_44844_n351) );
  AND2X2 AND2X2_2785 ( .A(u0_u4__abc_44844_n351), .B(u0_u4__abc_44844_n347), .Y(u0_u4_tms_23__FF_INPUT) );
  AND2X2 AND2X2_2786 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf6), .B(u0_u4__abc_44844_n354), .Y(u0_u4__abc_44844_n355) );
  AND2X2 AND2X2_2787 ( .A(u0_u4__abc_44844_n356), .B(u0_u4__abc_44844_n209_1_bF_buf7), .Y(u0_u4__abc_44844_n357) );
  AND2X2 AND2X2_2788 ( .A(u0_u4__abc_44844_n357), .B(u0_u4__abc_44844_n353), .Y(u0_u4_tms_24__FF_INPUT) );
  AND2X2 AND2X2_2789 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf4), .B(u0_u4__abc_44844_n360), .Y(u0_u4__abc_44844_n361) );
  AND2X2 AND2X2_279 ( .A(u0__abc_49347_n1481), .B(u0__abc_49347_n1180_1_bF_buf5), .Y(u0__abc_49347_n1482) );
  AND2X2 AND2X2_2790 ( .A(u0_u4__abc_44844_n362), .B(u0_u4__abc_44844_n209_1_bF_buf6), .Y(u0_u4__abc_44844_n363) );
  AND2X2 AND2X2_2791 ( .A(u0_u4__abc_44844_n363), .B(u0_u4__abc_44844_n359), .Y(u0_u4_tms_25__FF_INPUT) );
  AND2X2 AND2X2_2792 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf2), .B(u0_u4__abc_44844_n366), .Y(u0_u4__abc_44844_n367) );
  AND2X2 AND2X2_2793 ( .A(u0_u4__abc_44844_n368), .B(u0_u4__abc_44844_n209_1_bF_buf5), .Y(u0_u4__abc_44844_n369) );
  AND2X2 AND2X2_2794 ( .A(u0_u4__abc_44844_n369), .B(u0_u4__abc_44844_n365), .Y(u0_u4_tms_26__FF_INPUT) );
  AND2X2 AND2X2_2795 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf0), .B(u0_u4__abc_44844_n372), .Y(u0_u4__abc_44844_n373) );
  AND2X2 AND2X2_2796 ( .A(u0_u4__abc_44844_n374), .B(u0_u4__abc_44844_n209_1_bF_buf4), .Y(u0_u4__abc_44844_n375) );
  AND2X2 AND2X2_2797 ( .A(u0_u4__abc_44844_n375), .B(u0_u4__abc_44844_n371), .Y(u0_u4_tms_27__FF_INPUT) );
  AND2X2 AND2X2_2798 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf6), .B(u0_u4__abc_44844_n378), .Y(u0_u4__abc_44844_n379) );
  AND2X2 AND2X2_2799 ( .A(u0_u4__abc_44844_n380), .B(u0_u4__abc_44844_n209_1_bF_buf3), .Y(u0_u4__abc_44844_n381) );
  AND2X2 AND2X2_28 ( .A(_abc_55805_n320), .B(_abc_55805_n321), .Y(tms_s_10_) );
  AND2X2 AND2X2_280 ( .A(spec_req_cs_3_bF_buf2), .B(u0_tms3_12_), .Y(u0__abc_49347_n1483) );
  AND2X2 AND2X2_2800 ( .A(u0_u4__abc_44844_n381), .B(u0_u4__abc_44844_n377), .Y(u0_u4_tms_28__FF_INPUT) );
  AND2X2 AND2X2_2801 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf4), .B(u0_u4__abc_44844_n384), .Y(u0_u4__abc_44844_n385) );
  AND2X2 AND2X2_2802 ( .A(u0_u4__abc_44844_n386), .B(u0_u4__abc_44844_n209_1_bF_buf2), .Y(u0_u4__abc_44844_n387) );
  AND2X2 AND2X2_2803 ( .A(u0_u4__abc_44844_n387), .B(u0_u4__abc_44844_n383), .Y(u0_u4_tms_29__FF_INPUT) );
  AND2X2 AND2X2_2804 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf2), .B(u0_u4__abc_44844_n390), .Y(u0_u4__abc_44844_n391) );
  AND2X2 AND2X2_2805 ( .A(u0_u4__abc_44844_n392), .B(u0_u4__abc_44844_n209_1_bF_buf1), .Y(u0_u4__abc_44844_n393) );
  AND2X2 AND2X2_2806 ( .A(u0_u4__abc_44844_n393), .B(u0_u4__abc_44844_n389), .Y(u0_u4_tms_30__FF_INPUT) );
  AND2X2 AND2X2_2807 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf0), .B(u0_u4__abc_44844_n396), .Y(u0_u4__abc_44844_n397) );
  AND2X2 AND2X2_2808 ( .A(u0_u4__abc_44844_n398), .B(u0_u4__abc_44844_n209_1_bF_buf0), .Y(u0_u4__abc_44844_n399) );
  AND2X2 AND2X2_2809 ( .A(u0_u4__abc_44844_n399), .B(u0_u4__abc_44844_n395), .Y(u0_u4_tms_31__FF_INPUT) );
  AND2X2 AND2X2_281 ( .A(u0__abc_49347_n1484), .B(u0__abc_49347_n1179_bF_buf5), .Y(u0__abc_49347_n1485) );
  AND2X2 AND2X2_2810 ( .A(u0_u4__abc_44844_n403), .B(u0_u4_lmr_req_we), .Y(u0_u4__abc_44844_n404) );
  AND2X2 AND2X2_2811 ( .A(u0_u4__abc_44844_n404), .B(u0_u4_inited), .Y(u0_u4__abc_44844_n405) );
  AND2X2 AND2X2_2812 ( .A(u0_u4__abc_44844_n407), .B(u0_lmr_req4), .Y(u0_u4__abc_44844_n408) );
  AND2X2 AND2X2_2813 ( .A(u0_u4__abc_44844_n406), .B(u0_u4__abc_44844_n408), .Y(u0_u4__abc_44844_n409) );
  AND2X2 AND2X2_2814 ( .A(u0_u4__abc_44844_n206_1), .B(u0_u4__abc_44844_n411), .Y(u0_u4_init_req_we_FF_INPUT) );
  AND2X2 AND2X2_2815 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf6), .B(u0_u4__abc_44844_n210_1), .Y(u0_u4__abc_44844_n414) );
  AND2X2 AND2X2_2816 ( .A(u0_u4__abc_44844_n415), .B(u0_u4__abc_44844_n209_1_bF_buf7), .Y(u0_u4__abc_44844_n416) );
  AND2X2 AND2X2_2817 ( .A(u0_u4__abc_44844_n416), .B(u0_u4__abc_44844_n413), .Y(u0_u4_csc_0__FF_INPUT) );
  AND2X2 AND2X2_2818 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf4), .B(u0_u4__abc_44844_n216_1), .Y(u0_u4__abc_44844_n419) );
  AND2X2 AND2X2_2819 ( .A(u0_u4__abc_44844_n420), .B(u0_u4__abc_44844_n209_1_bF_buf6), .Y(u0_u4__abc_44844_n421) );
  AND2X2 AND2X2_282 ( .A(spec_req_cs_2_bF_buf2), .B(u0_tms2_12_), .Y(u0__abc_49347_n1486) );
  AND2X2 AND2X2_2820 ( .A(u0_u4__abc_44844_n421), .B(u0_u4__abc_44844_n418), .Y(u0_u4_csc_1__FF_INPUT) );
  AND2X2 AND2X2_2821 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf2), .B(u0_u4__abc_44844_n222_1), .Y(u0_u4__abc_44844_n424) );
  AND2X2 AND2X2_2822 ( .A(u0_u4__abc_44844_n425), .B(u0_u4__abc_44844_n209_1_bF_buf5), .Y(u0_u4__abc_44844_n426) );
  AND2X2 AND2X2_2823 ( .A(u0_u4__abc_44844_n426), .B(u0_u4__abc_44844_n423), .Y(u0_u4_csc_2__FF_INPUT) );
  AND2X2 AND2X2_2824 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf0), .B(u0_u4__abc_44844_n228_1), .Y(u0_u4__abc_44844_n429) );
  AND2X2 AND2X2_2825 ( .A(u0_u4__abc_44844_n430), .B(u0_u4__abc_44844_n209_1_bF_buf4), .Y(u0_u4__abc_44844_n431) );
  AND2X2 AND2X2_2826 ( .A(u0_u4__abc_44844_n431), .B(u0_u4__abc_44844_n428), .Y(u0_u4_csc_3__FF_INPUT) );
  AND2X2 AND2X2_2827 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf6), .B(u0_u4__abc_44844_n234_1), .Y(u0_u4__abc_44844_n434) );
  AND2X2 AND2X2_2828 ( .A(u0_u4__abc_44844_n435), .B(u0_u4__abc_44844_n209_1_bF_buf3), .Y(u0_u4__abc_44844_n436) );
  AND2X2 AND2X2_2829 ( .A(u0_u4__abc_44844_n436), .B(u0_u4__abc_44844_n433), .Y(u0_u4_csc_4__FF_INPUT) );
  AND2X2 AND2X2_283 ( .A(u0__abc_49347_n1487), .B(u0__abc_49347_n1178_1_bF_buf5), .Y(u0__abc_49347_n1488_1) );
  AND2X2 AND2X2_2830 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf4), .B(u0_u4__abc_44844_n240_1), .Y(u0_u4__abc_44844_n439) );
  AND2X2 AND2X2_2831 ( .A(u0_u4__abc_44844_n440), .B(u0_u4__abc_44844_n209_1_bF_buf2), .Y(u0_u4__abc_44844_n441) );
  AND2X2 AND2X2_2832 ( .A(u0_u4__abc_44844_n441), .B(u0_u4__abc_44844_n438), .Y(u0_u4_csc_5__FF_INPUT) );
  AND2X2 AND2X2_2833 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf2), .B(u0_u4__abc_44844_n246_1), .Y(u0_u4__abc_44844_n444) );
  AND2X2 AND2X2_2834 ( .A(u0_u4__abc_44844_n445), .B(u0_u4__abc_44844_n209_1_bF_buf1), .Y(u0_u4__abc_44844_n446) );
  AND2X2 AND2X2_2835 ( .A(u0_u4__abc_44844_n446), .B(u0_u4__abc_44844_n443), .Y(u0_u4_csc_6__FF_INPUT) );
  AND2X2 AND2X2_2836 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf0), .B(u0_u4__abc_44844_n252_1), .Y(u0_u4__abc_44844_n449) );
  AND2X2 AND2X2_2837 ( .A(u0_u4__abc_44844_n450), .B(u0_u4__abc_44844_n209_1_bF_buf0), .Y(u0_u4__abc_44844_n451) );
  AND2X2 AND2X2_2838 ( .A(u0_u4__abc_44844_n451), .B(u0_u4__abc_44844_n448), .Y(u0_u4_csc_7__FF_INPUT) );
  AND2X2 AND2X2_2839 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf6), .B(u0_u4__abc_44844_n258_1), .Y(u0_u4__abc_44844_n454) );
  AND2X2 AND2X2_284 ( .A(spec_req_cs_1_bF_buf2), .B(u0_tms1_12_), .Y(u0__abc_49347_n1489_1) );
  AND2X2 AND2X2_2840 ( .A(u0_u4__abc_44844_n455), .B(u0_u4__abc_44844_n209_1_bF_buf7), .Y(u0_u4__abc_44844_n456) );
  AND2X2 AND2X2_2841 ( .A(u0_u4__abc_44844_n456), .B(u0_u4__abc_44844_n453), .Y(u0_u4_csc_8__FF_INPUT) );
  AND2X2 AND2X2_2842 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf4), .B(u0_u4__abc_44844_n264), .Y(u0_u4__abc_44844_n459) );
  AND2X2 AND2X2_2843 ( .A(u0_u4__abc_44844_n460), .B(u0_u4__abc_44844_n209_1_bF_buf6), .Y(u0_u4__abc_44844_n461) );
  AND2X2 AND2X2_2844 ( .A(u0_u4__abc_44844_n461), .B(u0_u4__abc_44844_n458), .Y(u0_u4_csc_9__FF_INPUT) );
  AND2X2 AND2X2_2845 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf2), .B(u0_u4__abc_44844_n270_1), .Y(u0_u4__abc_44844_n464) );
  AND2X2 AND2X2_2846 ( .A(u0_u4__abc_44844_n465), .B(u0_u4__abc_44844_n209_1_bF_buf5), .Y(u0_u4__abc_44844_n466) );
  AND2X2 AND2X2_2847 ( .A(u0_u4__abc_44844_n466), .B(u0_u4__abc_44844_n463), .Y(u0_u4_csc_10__FF_INPUT) );
  AND2X2 AND2X2_2848 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf0), .B(u0_u4__abc_44844_n276_1), .Y(u0_u4__abc_44844_n469) );
  AND2X2 AND2X2_2849 ( .A(u0_u4__abc_44844_n470), .B(u0_u4__abc_44844_n209_1_bF_buf4), .Y(u0_u4__abc_44844_n471) );
  AND2X2 AND2X2_285 ( .A(u0__abc_49347_n1175_bF_buf0), .B(u0__abc_49347_n1492), .Y(u0__abc_49347_n1493) );
  AND2X2 AND2X2_2850 ( .A(u0_u4__abc_44844_n471), .B(u0_u4__abc_44844_n468), .Y(u0_u4_csc_11__FF_INPUT) );
  AND2X2 AND2X2_2851 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf6), .B(u0_u4__abc_44844_n282), .Y(u0_u4__abc_44844_n474) );
  AND2X2 AND2X2_2852 ( .A(u0_u4__abc_44844_n475), .B(u0_u4__abc_44844_n209_1_bF_buf3), .Y(u0_u4__abc_44844_n476) );
  AND2X2 AND2X2_2853 ( .A(u0_u4__abc_44844_n476), .B(u0_u4__abc_44844_n473), .Y(u0_u4_csc_12__FF_INPUT) );
  AND2X2 AND2X2_2854 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf4), .B(u0_u4__abc_44844_n288), .Y(u0_u4__abc_44844_n479) );
  AND2X2 AND2X2_2855 ( .A(u0_u4__abc_44844_n480), .B(u0_u4__abc_44844_n209_1_bF_buf2), .Y(u0_u4__abc_44844_n481) );
  AND2X2 AND2X2_2856 ( .A(u0_u4__abc_44844_n481), .B(u0_u4__abc_44844_n478), .Y(u0_u4_csc_13__FF_INPUT) );
  AND2X2 AND2X2_2857 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf2), .B(u0_u4__abc_44844_n294), .Y(u0_u4__abc_44844_n484) );
  AND2X2 AND2X2_2858 ( .A(u0_u4__abc_44844_n485), .B(u0_u4__abc_44844_n209_1_bF_buf1), .Y(u0_u4__abc_44844_n486) );
  AND2X2 AND2X2_2859 ( .A(u0_u4__abc_44844_n486), .B(u0_u4__abc_44844_n483), .Y(u0_u4_csc_14__FF_INPUT) );
  AND2X2 AND2X2_286 ( .A(u0__abc_49347_n1491), .B(u0__abc_49347_n1493), .Y(u0__abc_49347_n1494) );
  AND2X2 AND2X2_2860 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf0), .B(u0_u4__abc_44844_n300), .Y(u0_u4__abc_44844_n489) );
  AND2X2 AND2X2_2861 ( .A(u0_u4__abc_44844_n490), .B(u0_u4__abc_44844_n209_1_bF_buf0), .Y(u0_u4__abc_44844_n491) );
  AND2X2 AND2X2_2862 ( .A(u0_u4__abc_44844_n491), .B(u0_u4__abc_44844_n488), .Y(u0_u4_csc_15__FF_INPUT) );
  AND2X2 AND2X2_2863 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf6), .B(u0_u4__abc_44844_n306_1), .Y(u0_u4__abc_44844_n494) );
  AND2X2 AND2X2_2864 ( .A(u0_u4__abc_44844_n495), .B(u0_u4__abc_44844_n209_1_bF_buf7), .Y(u0_u4__abc_44844_n496) );
  AND2X2 AND2X2_2865 ( .A(u0_u4__abc_44844_n496), .B(u0_u4__abc_44844_n493), .Y(u0_u4_csc_16__FF_INPUT) );
  AND2X2 AND2X2_2866 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf4), .B(u0_u4__abc_44844_n312), .Y(u0_u4__abc_44844_n499) );
  AND2X2 AND2X2_2867 ( .A(u0_u4__abc_44844_n500), .B(u0_u4__abc_44844_n209_1_bF_buf6), .Y(u0_u4__abc_44844_n501) );
  AND2X2 AND2X2_2868 ( .A(u0_u4__abc_44844_n501), .B(u0_u4__abc_44844_n498), .Y(u0_u4_csc_17__FF_INPUT) );
  AND2X2 AND2X2_2869 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf2), .B(u0_u4__abc_44844_n318_1), .Y(u0_u4__abc_44844_n504) );
  AND2X2 AND2X2_287 ( .A(u0__abc_49347_n1176_1_bF_buf0), .B(sp_tms_13_), .Y(u0__abc_49347_n1496) );
  AND2X2 AND2X2_2870 ( .A(u0_u4__abc_44844_n505), .B(u0_u4__abc_44844_n209_1_bF_buf5), .Y(u0_u4__abc_44844_n506) );
  AND2X2 AND2X2_2871 ( .A(u0_u4__abc_44844_n506), .B(u0_u4__abc_44844_n503), .Y(u0_u4_csc_18__FF_INPUT) );
  AND2X2 AND2X2_2872 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf0), .B(u0_u4__abc_44844_n324_1), .Y(u0_u4__abc_44844_n509) );
  AND2X2 AND2X2_2873 ( .A(u0_u4__abc_44844_n510), .B(u0_u4__abc_44844_n209_1_bF_buf4), .Y(u0_u4__abc_44844_n511) );
  AND2X2 AND2X2_2874 ( .A(u0_u4__abc_44844_n511), .B(u0_u4__abc_44844_n508), .Y(u0_u4_csc_19__FF_INPUT) );
  AND2X2 AND2X2_2875 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf6), .B(u0_u4__abc_44844_n330), .Y(u0_u4__abc_44844_n514) );
  AND2X2 AND2X2_2876 ( .A(u0_u4__abc_44844_n515), .B(u0_u4__abc_44844_n209_1_bF_buf3), .Y(u0_u4__abc_44844_n516) );
  AND2X2 AND2X2_2877 ( .A(u0_u4__abc_44844_n516), .B(u0_u4__abc_44844_n513), .Y(u0_u4_csc_20__FF_INPUT) );
  AND2X2 AND2X2_2878 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf4), .B(u0_u4__abc_44844_n336), .Y(u0_u4__abc_44844_n519) );
  AND2X2 AND2X2_2879 ( .A(u0_u4__abc_44844_n520), .B(u0_u4__abc_44844_n209_1_bF_buf2), .Y(u0_u4__abc_44844_n521) );
  AND2X2 AND2X2_288 ( .A(spec_req_cs_5_bF_buf1), .B(u0_tms5_13_), .Y(u0__abc_49347_n1497_1) );
  AND2X2 AND2X2_2880 ( .A(u0_u4__abc_44844_n521), .B(u0_u4__abc_44844_n518), .Y(u0_u4_csc_21__FF_INPUT) );
  AND2X2 AND2X2_2881 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf2), .B(u0_u4__abc_44844_n342), .Y(u0_u4__abc_44844_n524) );
  AND2X2 AND2X2_2882 ( .A(u0_u4__abc_44844_n525), .B(u0_u4__abc_44844_n209_1_bF_buf1), .Y(u0_u4__abc_44844_n526) );
  AND2X2 AND2X2_2883 ( .A(u0_u4__abc_44844_n526), .B(u0_u4__abc_44844_n523), .Y(u0_u4_csc_22__FF_INPUT) );
  AND2X2 AND2X2_2884 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf0), .B(u0_u4__abc_44844_n348), .Y(u0_u4__abc_44844_n529) );
  AND2X2 AND2X2_2885 ( .A(u0_u4__abc_44844_n530), .B(u0_u4__abc_44844_n209_1_bF_buf0), .Y(u0_u4__abc_44844_n531) );
  AND2X2 AND2X2_2886 ( .A(u0_u4__abc_44844_n531), .B(u0_u4__abc_44844_n528), .Y(u0_u4_csc_23__FF_INPUT) );
  AND2X2 AND2X2_2887 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf6), .B(u0_u4__abc_44844_n354), .Y(u0_u4__abc_44844_n534) );
  AND2X2 AND2X2_2888 ( .A(u0_u4__abc_44844_n535), .B(u0_u4__abc_44844_n209_1_bF_buf7), .Y(u0_u4__abc_44844_n536) );
  AND2X2 AND2X2_2889 ( .A(u0_u4__abc_44844_n536), .B(u0_u4__abc_44844_n533), .Y(u0_u4_csc_24__FF_INPUT) );
  AND2X2 AND2X2_289 ( .A(u0__abc_49347_n1499), .B(u0__abc_49347_n1185_bF_buf4), .Y(u0__abc_49347_n1500) );
  AND2X2 AND2X2_2890 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf4), .B(u0_u4__abc_44844_n360), .Y(u0_u4__abc_44844_n539) );
  AND2X2 AND2X2_2891 ( .A(u0_u4__abc_44844_n540), .B(u0_u4__abc_44844_n209_1_bF_buf6), .Y(u0_u4__abc_44844_n541) );
  AND2X2 AND2X2_2892 ( .A(u0_u4__abc_44844_n541), .B(u0_u4__abc_44844_n538), .Y(u0_u4_csc_25__FF_INPUT) );
  AND2X2 AND2X2_2893 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf2), .B(u0_u4__abc_44844_n366), .Y(u0_u4__abc_44844_n544) );
  AND2X2 AND2X2_2894 ( .A(u0_u4__abc_44844_n545), .B(u0_u4__abc_44844_n209_1_bF_buf5), .Y(u0_u4__abc_44844_n546) );
  AND2X2 AND2X2_2895 ( .A(u0_u4__abc_44844_n546), .B(u0_u4__abc_44844_n543), .Y(u0_u4_csc_26__FF_INPUT) );
  AND2X2 AND2X2_2896 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf0), .B(u0_u4__abc_44844_n372), .Y(u0_u4__abc_44844_n549) );
  AND2X2 AND2X2_2897 ( .A(u0_u4__abc_44844_n550), .B(u0_u4__abc_44844_n209_1_bF_buf4), .Y(u0_u4__abc_44844_n551) );
  AND2X2 AND2X2_2898 ( .A(u0_u4__abc_44844_n551), .B(u0_u4__abc_44844_n548), .Y(u0_u4_csc_27__FF_INPUT) );
  AND2X2 AND2X2_2899 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf6), .B(u0_u4__abc_44844_n378), .Y(u0_u4__abc_44844_n554) );
  AND2X2 AND2X2_29 ( .A(_abc_55805_n323), .B(_abc_55805_n324), .Y(tms_s_11_) );
  AND2X2 AND2X2_290 ( .A(u0__abc_49347_n1500), .B(u0__abc_49347_n1498_1), .Y(u0__abc_49347_n1501) );
  AND2X2 AND2X2_2900 ( .A(u0_u4__abc_44844_n555), .B(u0_u4__abc_44844_n209_1_bF_buf3), .Y(u0_u4__abc_44844_n556) );
  AND2X2 AND2X2_2901 ( .A(u0_u4__abc_44844_n556), .B(u0_u4__abc_44844_n553), .Y(u0_u4_csc_28__FF_INPUT) );
  AND2X2 AND2X2_2902 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf4), .B(u0_u4__abc_44844_n384), .Y(u0_u4__abc_44844_n559) );
  AND2X2 AND2X2_2903 ( .A(u0_u4__abc_44844_n560), .B(u0_u4__abc_44844_n209_1_bF_buf2), .Y(u0_u4__abc_44844_n561) );
  AND2X2 AND2X2_2904 ( .A(u0_u4__abc_44844_n561), .B(u0_u4__abc_44844_n558), .Y(u0_u4_csc_29__FF_INPUT) );
  AND2X2 AND2X2_2905 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf2), .B(u0_u4__abc_44844_n390), .Y(u0_u4__abc_44844_n564) );
  AND2X2 AND2X2_2906 ( .A(u0_u4__abc_44844_n565), .B(u0_u4__abc_44844_n209_1_bF_buf1), .Y(u0_u4__abc_44844_n566) );
  AND2X2 AND2X2_2907 ( .A(u0_u4__abc_44844_n566), .B(u0_u4__abc_44844_n563), .Y(u0_u4_csc_30__FF_INPUT) );
  AND2X2 AND2X2_2908 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf0), .B(u0_u4__abc_44844_n396), .Y(u0_u4__abc_44844_n569) );
  AND2X2 AND2X2_2909 ( .A(u0_u4__abc_44844_n570), .B(u0_u4__abc_44844_n209_1_bF_buf0), .Y(u0_u4__abc_44844_n571) );
  AND2X2 AND2X2_291 ( .A(u0__abc_49347_n1502), .B(u0__abc_49347_n1181_bF_buf4), .Y(u0__abc_49347_n1503) );
  AND2X2 AND2X2_2910 ( .A(u0_u4__abc_44844_n571), .B(u0_u4__abc_44844_n568), .Y(u0_u4_csc_31__FF_INPUT) );
  AND2X2 AND2X2_2911 ( .A(u0_u4__abc_44844_n573), .B(u0_init_req4), .Y(u0_u4__abc_44844_n574) );
  AND2X2 AND2X2_2912 ( .A(u0_u4__abc_44844_n575), .B(u0_csc4_0_), .Y(u0_u4__abc_44844_n576) );
  AND2X2 AND2X2_2913 ( .A(u0_u4__abc_44844_n576), .B(u0_u4_init_req_we), .Y(u0_u4__abc_44844_n577) );
  AND2X2 AND2X2_2914 ( .A(u0_u4__abc_44844_n403), .B(u0_u4__abc_44844_n577), .Y(u0_u4__abc_44844_n578) );
  AND2X2 AND2X2_2915 ( .A(u0_csc4_8_), .B(wb_we_i), .Y(u0_u4__abc_44844_n581) );
  AND2X2 AND2X2_2916 ( .A(u0_csc4_20_), .B(u0_csc_mask_4_), .Y(u0_u4__abc_44844_n582) );
  AND2X2 AND2X2_2917 ( .A(u0_csc_mask_4_), .B(wb_addr_i_25_bF_buf3), .Y(u0_u4__abc_44844_n583) );
  AND2X2 AND2X2_2918 ( .A(u0_csc_mask_3_), .B(\wb_addr_i[24] ), .Y(u0_u4__abc_44844_n586) );
  AND2X2 AND2X2_2919 ( .A(u0_csc4_19_), .B(u0_csc_mask_3_), .Y(u0_u4__abc_44844_n587) );
  AND2X2 AND2X2_292 ( .A(spec_req_cs_4_bF_buf1), .B(u0_tms4_13_), .Y(u0__abc_49347_n1504) );
  AND2X2 AND2X2_2920 ( .A(u0_u4__abc_44844_n585), .B(u0_u4__abc_44844_n589), .Y(u0_u4__abc_44844_n590) );
  AND2X2 AND2X2_2921 ( .A(u0_csc4_18_), .B(u0_csc_mask_2_), .Y(u0_u4__abc_44844_n592) );
  AND2X2 AND2X2_2922 ( .A(u0_u4__abc_44844_n592), .B(u0_u4__abc_44844_n591), .Y(u0_u4__abc_44844_n593) );
  AND2X2 AND2X2_2923 ( .A(u0_u4__abc_44844_n596), .B(u0_u4__abc_44844_n594), .Y(u0_u4__abc_44844_n597) );
  AND2X2 AND2X2_2924 ( .A(u0_u4__abc_44844_n590), .B(u0_u4__abc_44844_n597), .Y(u0_u4__abc_44844_n598) );
  AND2X2 AND2X2_2925 ( .A(u0_csc4_22_), .B(u0_csc_mask_6_), .Y(u0_u4__abc_44844_n599) );
  AND2X2 AND2X2_2926 ( .A(u0_csc_mask_6_), .B(\wb_addr_i[27] ), .Y(u0_u4__abc_44844_n600) );
  AND2X2 AND2X2_2927 ( .A(u0_csc_mask_5_), .B(\wb_addr_i[26] ), .Y(u0_u4__abc_44844_n603) );
  AND2X2 AND2X2_2928 ( .A(u0_csc4_21_), .B(u0_csc_mask_5_), .Y(u0_u4__abc_44844_n604) );
  AND2X2 AND2X2_2929 ( .A(u0_u4__abc_44844_n602), .B(u0_u4__abc_44844_n606), .Y(u0_u4__abc_44844_n607) );
  AND2X2 AND2X2_293 ( .A(u0__abc_49347_n1505), .B(u0__abc_49347_n1180_1_bF_buf4), .Y(u0__abc_49347_n1506_1) );
  AND2X2 AND2X2_2930 ( .A(u0_u4__abc_44844_n582), .B(u0_u4__abc_44844_n608), .Y(u0_u4__abc_44844_n609) );
  AND2X2 AND2X2_2931 ( .A(u0_u4__abc_44844_n612), .B(u0_u4__abc_44844_n610), .Y(u0_u4__abc_44844_n613) );
  AND2X2 AND2X2_2932 ( .A(u0_u4__abc_44844_n607), .B(u0_u4__abc_44844_n613), .Y(u0_u4__abc_44844_n614) );
  AND2X2 AND2X2_2933 ( .A(u0_u4__abc_44844_n598), .B(u0_u4__abc_44844_n614), .Y(u0_u4__abc_44844_n615) );
  AND2X2 AND2X2_2934 ( .A(u0_u4__abc_44844_n601), .B(u0_u4__abc_44844_n599), .Y(u0_u4__abc_44844_n616) );
  AND2X2 AND2X2_2935 ( .A(u0_csc_mask_7_), .B(\wb_addr_i[28] ), .Y(u0_u4__abc_44844_n618) );
  AND2X2 AND2X2_2936 ( .A(u0_csc4_23_), .B(u0_csc_mask_7_), .Y(u0_u4__abc_44844_n620) );
  AND2X2 AND2X2_2937 ( .A(u0_u4__abc_44844_n617), .B(u0_u4__abc_44844_n621), .Y(u0_u4__abc_44844_n622) );
  AND2X2 AND2X2_2938 ( .A(u0_u4__abc_44844_n622), .B(u0_u4__abc_44844_n624), .Y(u0_u4__abc_44844_n625) );
  AND2X2 AND2X2_2939 ( .A(u0_u4__abc_44844_n615), .B(u0_u4__abc_44844_n625), .Y(u0_u4__abc_44844_n626) );
  AND2X2 AND2X2_294 ( .A(spec_req_cs_3_bF_buf1), .B(u0_tms3_13_), .Y(u0__abc_49347_n1507_1) );
  AND2X2 AND2X2_2940 ( .A(u0_csc_mask_2_), .B(wb_addr_i_23_bF_buf2), .Y(u0_u4__abc_44844_n627) );
  AND2X2 AND2X2_2941 ( .A(u0_csc_mask_1_), .B(\wb_addr_i[22] ), .Y(u0_u4__abc_44844_n630) );
  AND2X2 AND2X2_2942 ( .A(u0_csc4_17_), .B(u0_csc_mask_1_), .Y(u0_u4__abc_44844_n631) );
  AND2X2 AND2X2_2943 ( .A(u0_u4__abc_44844_n629), .B(u0_u4__abc_44844_n633), .Y(u0_u4__abc_44844_n634) );
  AND2X2 AND2X2_2944 ( .A(u0_csc_mask_0_), .B(\wb_addr_i[21] ), .Y(u0_u4__abc_44844_n635) );
  AND2X2 AND2X2_2945 ( .A(u0_csc4_16_), .B(u0_csc_mask_0_), .Y(u0_u4__abc_44844_n636) );
  AND2X2 AND2X2_2946 ( .A(u0_u4__abc_44844_n638), .B(u0_u4__abc_44844_n640), .Y(u0_u4__abc_44844_n641) );
  AND2X2 AND2X2_2947 ( .A(u0_u4__abc_44844_n634), .B(u0_u4__abc_44844_n641), .Y(u0_u4__abc_44844_n642) );
  AND2X2 AND2X2_2948 ( .A(u0_u4__abc_44844_n644), .B(u0_csc4_0_), .Y(u0_u4__abc_44844_n645) );
  AND2X2 AND2X2_2949 ( .A(u0_u4__abc_44844_n642), .B(u0_u4__abc_44844_n645), .Y(u0_u4__abc_44844_n646) );
  AND2X2 AND2X2_295 ( .A(u0__abc_49347_n1508), .B(u0__abc_49347_n1179_bF_buf4), .Y(u0__abc_49347_n1509) );
  AND2X2 AND2X2_2950 ( .A(u0_u4__abc_44844_n626), .B(u0_u4__abc_44844_n646), .Y(u0_u4__abc_44844_n647) );
  AND2X2 AND2X2_2951 ( .A(u0_u4__abc_44844_n647), .B(u0_u4__abc_44844_n581), .Y(u0_u4_wp_err) );
  AND2X2 AND2X2_2952 ( .A(u0_u4__abc_44844_n647), .B(u0_u4__abc_44844_n649), .Y(u0_cs4) );
  AND2X2 AND2X2_2953 ( .A(u0_u5__abc_45296_n203), .B(u0_u5_lmr_req_we), .Y(u0_u5__abc_45296_n204_1) );
  AND2X2 AND2X2_2954 ( .A(u0_u5__abc_45296_n204_1), .B(u0_u5_inited), .Y(u0_u5__abc_45296_n205_1) );
  AND2X2 AND2X2_2955 ( .A(u0_u5__abc_45296_n207_1), .B(u0_lmr_req5), .Y(u0_u5__abc_45296_n208_1) );
  AND2X2 AND2X2_2956 ( .A(u0_u5__abc_45296_n206), .B(u0_u5__abc_45296_n208_1), .Y(u0_u5__abc_45296_n209) );
  AND2X2 AND2X2_2957 ( .A(u0_u5__abc_45296_n211_1), .B(u0_u5_addr_r_3_), .Y(u0_u5__abc_45296_n212) );
  AND2X2 AND2X2_2958 ( .A(u0_u5_addr_r_5_), .B(u0_u5_addr_r_4_), .Y(u0_u5__abc_45296_n213_1) );
  AND2X2 AND2X2_2959 ( .A(u0_u5__abc_45296_n213_1), .B(u0_rf_we), .Y(u0_u5__abc_45296_n214_1) );
  AND2X2 AND2X2_296 ( .A(spec_req_cs_2_bF_buf1), .B(u0_tms2_13_), .Y(u0__abc_49347_n1510) );
  AND2X2 AND2X2_2960 ( .A(u0_u5__abc_45296_n214_1), .B(u0_u5__abc_45296_n212), .Y(u0_u5__abc_45296_n215) );
  AND2X2 AND2X2_2961 ( .A(u0_u5__abc_45296_n215), .B(u0_u5_addr_r_2_), .Y(u0_u5_lmr_req_we_FF_INPUT) );
  AND2X2 AND2X2_2962 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf6), .B(u0_u5__abc_45296_n219_1), .Y(u0_u5__abc_45296_n220_1) );
  AND2X2 AND2X2_2963 ( .A(u0_u5__abc_45296_n221), .B(u0_u5__abc_45296_n218_bF_buf7), .Y(u0_u5__abc_45296_n222_1) );
  AND2X2 AND2X2_2964 ( .A(u0_u5__abc_45296_n222_1), .B(u0_u5__abc_45296_n217_1), .Y(u0_u5_tms_0__FF_INPUT) );
  AND2X2 AND2X2_2965 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf4), .B(u0_u5__abc_45296_n225_1), .Y(u0_u5__abc_45296_n226_1) );
  AND2X2 AND2X2_2966 ( .A(u0_u5__abc_45296_n227), .B(u0_u5__abc_45296_n218_bF_buf6), .Y(u0_u5__abc_45296_n228_1) );
  AND2X2 AND2X2_2967 ( .A(u0_u5__abc_45296_n228_1), .B(u0_u5__abc_45296_n224), .Y(u0_u5_tms_1__FF_INPUT) );
  AND2X2 AND2X2_2968 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf2), .B(u0_u5__abc_45296_n231_1), .Y(u0_u5__abc_45296_n232_1) );
  AND2X2 AND2X2_2969 ( .A(u0_u5__abc_45296_n233), .B(u0_u5__abc_45296_n218_bF_buf5), .Y(u0_u5__abc_45296_n234_1) );
  AND2X2 AND2X2_297 ( .A(u0__abc_49347_n1511), .B(u0__abc_49347_n1178_1_bF_buf4), .Y(u0__abc_49347_n1512) );
  AND2X2 AND2X2_2970 ( .A(u0_u5__abc_45296_n234_1), .B(u0_u5__abc_45296_n230), .Y(u0_u5_tms_2__FF_INPUT) );
  AND2X2 AND2X2_2971 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf0), .B(u0_u5__abc_45296_n237_1), .Y(u0_u5__abc_45296_n238_1) );
  AND2X2 AND2X2_2972 ( .A(u0_u5__abc_45296_n239), .B(u0_u5__abc_45296_n218_bF_buf4), .Y(u0_u5__abc_45296_n240_1) );
  AND2X2 AND2X2_2973 ( .A(u0_u5__abc_45296_n240_1), .B(u0_u5__abc_45296_n236), .Y(u0_u5_tms_3__FF_INPUT) );
  AND2X2 AND2X2_2974 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf6), .B(u0_u5__abc_45296_n243_1), .Y(u0_u5__abc_45296_n244_1) );
  AND2X2 AND2X2_2975 ( .A(u0_u5__abc_45296_n245), .B(u0_u5__abc_45296_n218_bF_buf3), .Y(u0_u5__abc_45296_n246_1) );
  AND2X2 AND2X2_2976 ( .A(u0_u5__abc_45296_n246_1), .B(u0_u5__abc_45296_n242), .Y(u0_u5_tms_4__FF_INPUT) );
  AND2X2 AND2X2_2977 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf4), .B(u0_u5__abc_45296_n249_1), .Y(u0_u5__abc_45296_n250_1) );
  AND2X2 AND2X2_2978 ( .A(u0_u5__abc_45296_n251), .B(u0_u5__abc_45296_n218_bF_buf2), .Y(u0_u5__abc_45296_n252_1) );
  AND2X2 AND2X2_2979 ( .A(u0_u5__abc_45296_n252_1), .B(u0_u5__abc_45296_n248), .Y(u0_u5_tms_5__FF_INPUT) );
  AND2X2 AND2X2_298 ( .A(spec_req_cs_1_bF_buf1), .B(u0_tms1_13_), .Y(u0__abc_49347_n1513) );
  AND2X2 AND2X2_2980 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf2), .B(u0_u5__abc_45296_n255_1), .Y(u0_u5__abc_45296_n256) );
  AND2X2 AND2X2_2981 ( .A(u0_u5__abc_45296_n257), .B(u0_u5__abc_45296_n218_bF_buf1), .Y(u0_u5__abc_45296_n258) );
  AND2X2 AND2X2_2982 ( .A(u0_u5__abc_45296_n258), .B(u0_u5__abc_45296_n254), .Y(u0_u5_tms_6__FF_INPUT) );
  AND2X2 AND2X2_2983 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf0), .B(u0_u5__abc_45296_n261), .Y(u0_u5__abc_45296_n262_1) );
  AND2X2 AND2X2_2984 ( .A(u0_u5__abc_45296_n263), .B(u0_u5__abc_45296_n218_bF_buf0), .Y(u0_u5__abc_45296_n264) );
  AND2X2 AND2X2_2985 ( .A(u0_u5__abc_45296_n264), .B(u0_u5__abc_45296_n260_1), .Y(u0_u5_tms_7__FF_INPUT) );
  AND2X2 AND2X2_2986 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf6), .B(u0_u5__abc_45296_n267), .Y(u0_u5__abc_45296_n268_1) );
  AND2X2 AND2X2_2987 ( .A(u0_u5__abc_45296_n269), .B(u0_u5__abc_45296_n218_bF_buf7), .Y(u0_u5__abc_45296_n270) );
  AND2X2 AND2X2_2988 ( .A(u0_u5__abc_45296_n270), .B(u0_u5__abc_45296_n266_1), .Y(u0_u5_tms_8__FF_INPUT) );
  AND2X2 AND2X2_2989 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf4), .B(u0_u5__abc_45296_n273_1), .Y(u0_u5__abc_45296_n274) );
  AND2X2 AND2X2_299 ( .A(u0__abc_49347_n1175_bF_buf6), .B(u0__abc_49347_n1516_1), .Y(u0__abc_49347_n1517) );
  AND2X2 AND2X2_2990 ( .A(u0_u5__abc_45296_n275_1), .B(u0_u5__abc_45296_n218_bF_buf6), .Y(u0_u5__abc_45296_n276) );
  AND2X2 AND2X2_2991 ( .A(u0_u5__abc_45296_n276), .B(u0_u5__abc_45296_n272), .Y(u0_u5_tms_9__FF_INPUT) );
  AND2X2 AND2X2_2992 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf2), .B(u0_u5__abc_45296_n279_1), .Y(u0_u5__abc_45296_n280) );
  AND2X2 AND2X2_2993 ( .A(u0_u5__abc_45296_n281), .B(u0_u5__abc_45296_n218_bF_buf5), .Y(u0_u5__abc_45296_n282) );
  AND2X2 AND2X2_2994 ( .A(u0_u5__abc_45296_n282), .B(u0_u5__abc_45296_n278), .Y(u0_u5_tms_10__FF_INPUT) );
  AND2X2 AND2X2_2995 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf0), .B(u0_u5__abc_45296_n285_1), .Y(u0_u5__abc_45296_n286) );
  AND2X2 AND2X2_2996 ( .A(u0_u5__abc_45296_n287_1), .B(u0_u5__abc_45296_n218_bF_buf4), .Y(u0_u5__abc_45296_n288) );
  AND2X2 AND2X2_2997 ( .A(u0_u5__abc_45296_n288), .B(u0_u5__abc_45296_n284), .Y(u0_u5_tms_11__FF_INPUT) );
  AND2X2 AND2X2_2998 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf6), .B(u0_u5__abc_45296_n291), .Y(u0_u5__abc_45296_n292) );
  AND2X2 AND2X2_2999 ( .A(u0_u5__abc_45296_n293), .B(u0_u5__abc_45296_n218_bF_buf3), .Y(u0_u5__abc_45296_n294) );
  AND2X2 AND2X2_3 ( .A(_abc_55805_n244_1), .B(_abc_55805_n246), .Y(obct_cs_0_) );
  AND2X2 AND2X2_30 ( .A(_abc_55805_n326), .B(_abc_55805_n327), .Y(tms_s_12_) );
  AND2X2 AND2X2_300 ( .A(u0__abc_49347_n1515_1), .B(u0__abc_49347_n1517), .Y(u0__abc_49347_n1518) );
  AND2X2 AND2X2_3000 ( .A(u0_u5__abc_45296_n294), .B(u0_u5__abc_45296_n290), .Y(u0_u5_tms_12__FF_INPUT) );
  AND2X2 AND2X2_3001 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf4), .B(u0_u5__abc_45296_n297), .Y(u0_u5__abc_45296_n298_1) );
  AND2X2 AND2X2_3002 ( .A(u0_u5__abc_45296_n299), .B(u0_u5__abc_45296_n218_bF_buf2), .Y(u0_u5__abc_45296_n300) );
  AND2X2 AND2X2_3003 ( .A(u0_u5__abc_45296_n300), .B(u0_u5__abc_45296_n296_1), .Y(u0_u5_tms_13__FF_INPUT) );
  AND2X2 AND2X2_3004 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf2), .B(u0_u5__abc_45296_n303), .Y(u0_u5__abc_45296_n304) );
  AND2X2 AND2X2_3005 ( .A(u0_u5__abc_45296_n305), .B(u0_u5__abc_45296_n218_bF_buf1), .Y(u0_u5__abc_45296_n306) );
  AND2X2 AND2X2_3006 ( .A(u0_u5__abc_45296_n306), .B(u0_u5__abc_45296_n302), .Y(u0_u5_tms_14__FF_INPUT) );
  AND2X2 AND2X2_3007 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf0), .B(u0_u5__abc_45296_n309), .Y(u0_u5__abc_45296_n310_1) );
  AND2X2 AND2X2_3008 ( .A(u0_u5__abc_45296_n311), .B(u0_u5__abc_45296_n218_bF_buf0), .Y(u0_u5__abc_45296_n312_1) );
  AND2X2 AND2X2_3009 ( .A(u0_u5__abc_45296_n312_1), .B(u0_u5__abc_45296_n308), .Y(u0_u5_tms_15__FF_INPUT) );
  AND2X2 AND2X2_301 ( .A(u0__abc_49347_n1176_1_bF_buf6), .B(sp_tms_14_), .Y(u0__abc_49347_n1520) );
  AND2X2 AND2X2_3010 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf6), .B(u0_u5__abc_45296_n315_1), .Y(u0_u5__abc_45296_n316_1) );
  AND2X2 AND2X2_3011 ( .A(u0_u5__abc_45296_n317_1), .B(u0_u5__abc_45296_n218_bF_buf7), .Y(u0_u5__abc_45296_n318) );
  AND2X2 AND2X2_3012 ( .A(u0_u5__abc_45296_n318), .B(u0_u5__abc_45296_n314_1), .Y(u0_u5_tms_16__FF_INPUT) );
  AND2X2 AND2X2_3013 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf4), .B(u0_u5__abc_45296_n321_1), .Y(u0_u5__abc_45296_n322) );
  AND2X2 AND2X2_3014 ( .A(u0_u5__abc_45296_n323_1), .B(u0_u5__abc_45296_n218_bF_buf6), .Y(u0_u5__abc_45296_n324_1) );
  AND2X2 AND2X2_3015 ( .A(u0_u5__abc_45296_n324_1), .B(u0_u5__abc_45296_n320), .Y(u0_u5_tms_17__FF_INPUT) );
  AND2X2 AND2X2_3016 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf2), .B(u0_u5__abc_45296_n327), .Y(u0_u5__abc_45296_n328) );
  AND2X2 AND2X2_3017 ( .A(u0_u5__abc_45296_n329), .B(u0_u5__abc_45296_n218_bF_buf5), .Y(u0_u5__abc_45296_n330) );
  AND2X2 AND2X2_3018 ( .A(u0_u5__abc_45296_n330), .B(u0_u5__abc_45296_n326), .Y(u0_u5_tms_18__FF_INPUT) );
  AND2X2 AND2X2_3019 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf0), .B(u0_u5__abc_45296_n333), .Y(u0_u5__abc_45296_n334) );
  AND2X2 AND2X2_302 ( .A(spec_req_cs_5_bF_buf0), .B(u0_tms5_14_), .Y(u0__abc_49347_n1521) );
  AND2X2 AND2X2_3020 ( .A(u0_u5__abc_45296_n335), .B(u0_u5__abc_45296_n218_bF_buf4), .Y(u0_u5__abc_45296_n336) );
  AND2X2 AND2X2_3021 ( .A(u0_u5__abc_45296_n336), .B(u0_u5__abc_45296_n332), .Y(u0_u5_tms_19__FF_INPUT) );
  AND2X2 AND2X2_3022 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf6), .B(u0_u5__abc_45296_n339), .Y(u0_u5__abc_45296_n340) );
  AND2X2 AND2X2_3023 ( .A(u0_u5__abc_45296_n341), .B(u0_u5__abc_45296_n218_bF_buf3), .Y(u0_u5__abc_45296_n342) );
  AND2X2 AND2X2_3024 ( .A(u0_u5__abc_45296_n342), .B(u0_u5__abc_45296_n338), .Y(u0_u5_tms_20__FF_INPUT) );
  AND2X2 AND2X2_3025 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf4), .B(u0_u5__abc_45296_n345), .Y(u0_u5__abc_45296_n346) );
  AND2X2 AND2X2_3026 ( .A(u0_u5__abc_45296_n347), .B(u0_u5__abc_45296_n218_bF_buf2), .Y(u0_u5__abc_45296_n348) );
  AND2X2 AND2X2_3027 ( .A(u0_u5__abc_45296_n348), .B(u0_u5__abc_45296_n344), .Y(u0_u5_tms_21__FF_INPUT) );
  AND2X2 AND2X2_3028 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf2), .B(u0_u5__abc_45296_n351), .Y(u0_u5__abc_45296_n352) );
  AND2X2 AND2X2_3029 ( .A(u0_u5__abc_45296_n353), .B(u0_u5__abc_45296_n218_bF_buf1), .Y(u0_u5__abc_45296_n354) );
  AND2X2 AND2X2_303 ( .A(u0__abc_49347_n1523), .B(u0__abc_49347_n1185_bF_buf3), .Y(u0__abc_49347_n1524_1) );
  AND2X2 AND2X2_3030 ( .A(u0_u5__abc_45296_n354), .B(u0_u5__abc_45296_n350), .Y(u0_u5_tms_22__FF_INPUT) );
  AND2X2 AND2X2_3031 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf0), .B(u0_u5__abc_45296_n357), .Y(u0_u5__abc_45296_n358) );
  AND2X2 AND2X2_3032 ( .A(u0_u5__abc_45296_n359), .B(u0_u5__abc_45296_n218_bF_buf0), .Y(u0_u5__abc_45296_n360) );
  AND2X2 AND2X2_3033 ( .A(u0_u5__abc_45296_n360), .B(u0_u5__abc_45296_n356), .Y(u0_u5_tms_23__FF_INPUT) );
  AND2X2 AND2X2_3034 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf6), .B(u0_u5__abc_45296_n363), .Y(u0_u5__abc_45296_n364) );
  AND2X2 AND2X2_3035 ( .A(u0_u5__abc_45296_n365), .B(u0_u5__abc_45296_n218_bF_buf7), .Y(u0_u5__abc_45296_n366) );
  AND2X2 AND2X2_3036 ( .A(u0_u5__abc_45296_n366), .B(u0_u5__abc_45296_n362), .Y(u0_u5_tms_24__FF_INPUT) );
  AND2X2 AND2X2_3037 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf4), .B(u0_u5__abc_45296_n369), .Y(u0_u5__abc_45296_n370) );
  AND2X2 AND2X2_3038 ( .A(u0_u5__abc_45296_n371), .B(u0_u5__abc_45296_n218_bF_buf6), .Y(u0_u5__abc_45296_n372) );
  AND2X2 AND2X2_3039 ( .A(u0_u5__abc_45296_n372), .B(u0_u5__abc_45296_n368), .Y(u0_u5_tms_25__FF_INPUT) );
  AND2X2 AND2X2_304 ( .A(u0__abc_49347_n1524_1), .B(u0__abc_49347_n1522), .Y(u0__abc_49347_n1525_1) );
  AND2X2 AND2X2_3040 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf2), .B(u0_u5__abc_45296_n375), .Y(u0_u5__abc_45296_n376) );
  AND2X2 AND2X2_3041 ( .A(u0_u5__abc_45296_n377), .B(u0_u5__abc_45296_n218_bF_buf5), .Y(u0_u5__abc_45296_n378) );
  AND2X2 AND2X2_3042 ( .A(u0_u5__abc_45296_n378), .B(u0_u5__abc_45296_n374), .Y(u0_u5_tms_26__FF_INPUT) );
  AND2X2 AND2X2_3043 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf0), .B(u0_u5__abc_45296_n381), .Y(u0_u5__abc_45296_n382) );
  AND2X2 AND2X2_3044 ( .A(u0_u5__abc_45296_n383), .B(u0_u5__abc_45296_n218_bF_buf4), .Y(u0_u5__abc_45296_n384) );
  AND2X2 AND2X2_3045 ( .A(u0_u5__abc_45296_n384), .B(u0_u5__abc_45296_n380), .Y(u0_u5_tms_27__FF_INPUT) );
  AND2X2 AND2X2_3046 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf6), .B(u0_u5__abc_45296_n387), .Y(u0_u5__abc_45296_n388) );
  AND2X2 AND2X2_3047 ( .A(u0_u5__abc_45296_n389), .B(u0_u5__abc_45296_n218_bF_buf3), .Y(u0_u5__abc_45296_n390) );
  AND2X2 AND2X2_3048 ( .A(u0_u5__abc_45296_n390), .B(u0_u5__abc_45296_n386), .Y(u0_u5_tms_28__FF_INPUT) );
  AND2X2 AND2X2_3049 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf4), .B(u0_u5__abc_45296_n393), .Y(u0_u5__abc_45296_n394) );
  AND2X2 AND2X2_305 ( .A(u0__abc_49347_n1526), .B(u0__abc_49347_n1181_bF_buf3), .Y(u0__abc_49347_n1527) );
  AND2X2 AND2X2_3050 ( .A(u0_u5__abc_45296_n395), .B(u0_u5__abc_45296_n218_bF_buf2), .Y(u0_u5__abc_45296_n396) );
  AND2X2 AND2X2_3051 ( .A(u0_u5__abc_45296_n396), .B(u0_u5__abc_45296_n392), .Y(u0_u5_tms_29__FF_INPUT) );
  AND2X2 AND2X2_3052 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf2), .B(u0_u5__abc_45296_n399), .Y(u0_u5__abc_45296_n400) );
  AND2X2 AND2X2_3053 ( .A(u0_u5__abc_45296_n401), .B(u0_u5__abc_45296_n218_bF_buf1), .Y(u0_u5__abc_45296_n402) );
  AND2X2 AND2X2_3054 ( .A(u0_u5__abc_45296_n402), .B(u0_u5__abc_45296_n398), .Y(u0_u5_tms_30__FF_INPUT) );
  AND2X2 AND2X2_3055 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf0), .B(u0_u5__abc_45296_n405), .Y(u0_u5__abc_45296_n406) );
  AND2X2 AND2X2_3056 ( .A(u0_u5__abc_45296_n407), .B(u0_u5__abc_45296_n218_bF_buf0), .Y(u0_u5__abc_45296_n408) );
  AND2X2 AND2X2_3057 ( .A(u0_u5__abc_45296_n408), .B(u0_u5__abc_45296_n404), .Y(u0_u5_tms_31__FF_INPUT) );
  AND2X2 AND2X2_3058 ( .A(u0_u5__abc_45296_n215), .B(u0_u5__abc_45296_n410), .Y(u0_u5_init_req_we_FF_INPUT) );
  AND2X2 AND2X2_3059 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf6), .B(u0_u5__abc_45296_n219_1), .Y(u0_u5__abc_45296_n413) );
  AND2X2 AND2X2_306 ( .A(spec_req_cs_4_bF_buf0), .B(u0_tms4_14_), .Y(u0__abc_49347_n1528) );
  AND2X2 AND2X2_3060 ( .A(u0_u5__abc_45296_n414), .B(u0_u5__abc_45296_n218_bF_buf7), .Y(u0_u5__abc_45296_n415) );
  AND2X2 AND2X2_3061 ( .A(u0_u5__abc_45296_n415), .B(u0_u5__abc_45296_n412), .Y(u0_u5_csc_0__FF_INPUT) );
  AND2X2 AND2X2_3062 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf4), .B(u0_u5__abc_45296_n225_1), .Y(u0_u5__abc_45296_n418) );
  AND2X2 AND2X2_3063 ( .A(u0_u5__abc_45296_n419), .B(u0_u5__abc_45296_n218_bF_buf6), .Y(u0_u5__abc_45296_n420) );
  AND2X2 AND2X2_3064 ( .A(u0_u5__abc_45296_n420), .B(u0_u5__abc_45296_n417), .Y(u0_u5_csc_1__FF_INPUT) );
  AND2X2 AND2X2_3065 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf2), .B(u0_u5__abc_45296_n231_1), .Y(u0_u5__abc_45296_n423) );
  AND2X2 AND2X2_3066 ( .A(u0_u5__abc_45296_n424), .B(u0_u5__abc_45296_n218_bF_buf5), .Y(u0_u5__abc_45296_n425) );
  AND2X2 AND2X2_3067 ( .A(u0_u5__abc_45296_n425), .B(u0_u5__abc_45296_n422), .Y(u0_u5_csc_2__FF_INPUT) );
  AND2X2 AND2X2_3068 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf0), .B(u0_u5__abc_45296_n237_1), .Y(u0_u5__abc_45296_n428) );
  AND2X2 AND2X2_3069 ( .A(u0_u5__abc_45296_n429), .B(u0_u5__abc_45296_n218_bF_buf4), .Y(u0_u5__abc_45296_n430) );
  AND2X2 AND2X2_307 ( .A(u0__abc_49347_n1529), .B(u0__abc_49347_n1180_1_bF_buf3), .Y(u0__abc_49347_n1530) );
  AND2X2 AND2X2_3070 ( .A(u0_u5__abc_45296_n430), .B(u0_u5__abc_45296_n427), .Y(u0_u5_csc_3__FF_INPUT) );
  AND2X2 AND2X2_3071 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf6), .B(u0_u5__abc_45296_n243_1), .Y(u0_u5__abc_45296_n433) );
  AND2X2 AND2X2_3072 ( .A(u0_u5__abc_45296_n434), .B(u0_u5__abc_45296_n218_bF_buf3), .Y(u0_u5__abc_45296_n435) );
  AND2X2 AND2X2_3073 ( .A(u0_u5__abc_45296_n435), .B(u0_u5__abc_45296_n432), .Y(u0_u5_csc_4__FF_INPUT) );
  AND2X2 AND2X2_3074 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf4), .B(u0_u5__abc_45296_n249_1), .Y(u0_u5__abc_45296_n438) );
  AND2X2 AND2X2_3075 ( .A(u0_u5__abc_45296_n439), .B(u0_u5__abc_45296_n218_bF_buf2), .Y(u0_u5__abc_45296_n440) );
  AND2X2 AND2X2_3076 ( .A(u0_u5__abc_45296_n440), .B(u0_u5__abc_45296_n437), .Y(u0_u5_csc_5__FF_INPUT) );
  AND2X2 AND2X2_3077 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf2), .B(u0_u5__abc_45296_n255_1), .Y(u0_u5__abc_45296_n443) );
  AND2X2 AND2X2_3078 ( .A(u0_u5__abc_45296_n444), .B(u0_u5__abc_45296_n218_bF_buf1), .Y(u0_u5__abc_45296_n445) );
  AND2X2 AND2X2_3079 ( .A(u0_u5__abc_45296_n445), .B(u0_u5__abc_45296_n442), .Y(u0_u5_csc_6__FF_INPUT) );
  AND2X2 AND2X2_308 ( .A(spec_req_cs_3_bF_buf0), .B(u0_tms3_14_), .Y(u0__abc_49347_n1531) );
  AND2X2 AND2X2_3080 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf0), .B(u0_u5__abc_45296_n261), .Y(u0_u5__abc_45296_n448) );
  AND2X2 AND2X2_3081 ( .A(u0_u5__abc_45296_n449), .B(u0_u5__abc_45296_n218_bF_buf0), .Y(u0_u5__abc_45296_n450) );
  AND2X2 AND2X2_3082 ( .A(u0_u5__abc_45296_n450), .B(u0_u5__abc_45296_n447), .Y(u0_u5_csc_7__FF_INPUT) );
  AND2X2 AND2X2_3083 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf6), .B(u0_u5__abc_45296_n267), .Y(u0_u5__abc_45296_n453) );
  AND2X2 AND2X2_3084 ( .A(u0_u5__abc_45296_n454), .B(u0_u5__abc_45296_n218_bF_buf7), .Y(u0_u5__abc_45296_n455) );
  AND2X2 AND2X2_3085 ( .A(u0_u5__abc_45296_n455), .B(u0_u5__abc_45296_n452), .Y(u0_u5_csc_8__FF_INPUT) );
  AND2X2 AND2X2_3086 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf4), .B(u0_u5__abc_45296_n273_1), .Y(u0_u5__abc_45296_n458) );
  AND2X2 AND2X2_3087 ( .A(u0_u5__abc_45296_n459), .B(u0_u5__abc_45296_n218_bF_buf6), .Y(u0_u5__abc_45296_n460) );
  AND2X2 AND2X2_3088 ( .A(u0_u5__abc_45296_n460), .B(u0_u5__abc_45296_n457), .Y(u0_u5_csc_9__FF_INPUT) );
  AND2X2 AND2X2_3089 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf2), .B(u0_u5__abc_45296_n279_1), .Y(u0_u5__abc_45296_n463) );
  AND2X2 AND2X2_309 ( .A(u0__abc_49347_n1532), .B(u0__abc_49347_n1179_bF_buf3), .Y(u0__abc_49347_n1533_1) );
  AND2X2 AND2X2_3090 ( .A(u0_u5__abc_45296_n464), .B(u0_u5__abc_45296_n218_bF_buf5), .Y(u0_u5__abc_45296_n465) );
  AND2X2 AND2X2_3091 ( .A(u0_u5__abc_45296_n465), .B(u0_u5__abc_45296_n462), .Y(u0_u5_csc_10__FF_INPUT) );
  AND2X2 AND2X2_3092 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf0), .B(u0_u5__abc_45296_n285_1), .Y(u0_u5__abc_45296_n468) );
  AND2X2 AND2X2_3093 ( .A(u0_u5__abc_45296_n469), .B(u0_u5__abc_45296_n218_bF_buf4), .Y(u0_u5__abc_45296_n470) );
  AND2X2 AND2X2_3094 ( .A(u0_u5__abc_45296_n470), .B(u0_u5__abc_45296_n467), .Y(u0_u5_csc_11__FF_INPUT) );
  AND2X2 AND2X2_3095 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf6), .B(u0_u5__abc_45296_n291), .Y(u0_u5__abc_45296_n473) );
  AND2X2 AND2X2_3096 ( .A(u0_u5__abc_45296_n474), .B(u0_u5__abc_45296_n218_bF_buf3), .Y(u0_u5__abc_45296_n475) );
  AND2X2 AND2X2_3097 ( .A(u0_u5__abc_45296_n475), .B(u0_u5__abc_45296_n472), .Y(u0_u5_csc_12__FF_INPUT) );
  AND2X2 AND2X2_3098 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf4), .B(u0_u5__abc_45296_n297), .Y(u0_u5__abc_45296_n478) );
  AND2X2 AND2X2_3099 ( .A(u0_u5__abc_45296_n479), .B(u0_u5__abc_45296_n218_bF_buf2), .Y(u0_u5__abc_45296_n480) );
  AND2X2 AND2X2_31 ( .A(_abc_55805_n329), .B(_abc_55805_n330), .Y(tms_s_13_) );
  AND2X2 AND2X2_310 ( .A(spec_req_cs_2_bF_buf0), .B(u0_tms2_14_), .Y(u0__abc_49347_n1534_1) );
  AND2X2 AND2X2_3100 ( .A(u0_u5__abc_45296_n480), .B(u0_u5__abc_45296_n477), .Y(u0_u5_csc_13__FF_INPUT) );
  AND2X2 AND2X2_3101 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf2), .B(u0_u5__abc_45296_n303), .Y(u0_u5__abc_45296_n483) );
  AND2X2 AND2X2_3102 ( .A(u0_u5__abc_45296_n484), .B(u0_u5__abc_45296_n218_bF_buf1), .Y(u0_u5__abc_45296_n485) );
  AND2X2 AND2X2_3103 ( .A(u0_u5__abc_45296_n485), .B(u0_u5__abc_45296_n482), .Y(u0_u5_csc_14__FF_INPUT) );
  AND2X2 AND2X2_3104 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf0), .B(u0_u5__abc_45296_n309), .Y(u0_u5__abc_45296_n488) );
  AND2X2 AND2X2_3105 ( .A(u0_u5__abc_45296_n489), .B(u0_u5__abc_45296_n218_bF_buf0), .Y(u0_u5__abc_45296_n490) );
  AND2X2 AND2X2_3106 ( .A(u0_u5__abc_45296_n490), .B(u0_u5__abc_45296_n487), .Y(u0_u5_csc_15__FF_INPUT) );
  AND2X2 AND2X2_3107 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf6), .B(u0_u5__abc_45296_n315_1), .Y(u0_u5__abc_45296_n493) );
  AND2X2 AND2X2_3108 ( .A(u0_u5__abc_45296_n494), .B(u0_u5__abc_45296_n218_bF_buf7), .Y(u0_u5__abc_45296_n495) );
  AND2X2 AND2X2_3109 ( .A(u0_u5__abc_45296_n495), .B(u0_u5__abc_45296_n492), .Y(u0_u5_csc_16__FF_INPUT) );
  AND2X2 AND2X2_311 ( .A(u0__abc_49347_n1535), .B(u0__abc_49347_n1178_1_bF_buf3), .Y(u0__abc_49347_n1536) );
  AND2X2 AND2X2_3110 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf4), .B(u0_u5__abc_45296_n321_1), .Y(u0_u5__abc_45296_n498) );
  AND2X2 AND2X2_3111 ( .A(u0_u5__abc_45296_n499), .B(u0_u5__abc_45296_n218_bF_buf6), .Y(u0_u5__abc_45296_n500) );
  AND2X2 AND2X2_3112 ( .A(u0_u5__abc_45296_n500), .B(u0_u5__abc_45296_n497), .Y(u0_u5_csc_17__FF_INPUT) );
  AND2X2 AND2X2_3113 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf2), .B(u0_u5__abc_45296_n327), .Y(u0_u5__abc_45296_n503) );
  AND2X2 AND2X2_3114 ( .A(u0_u5__abc_45296_n504), .B(u0_u5__abc_45296_n218_bF_buf5), .Y(u0_u5__abc_45296_n505) );
  AND2X2 AND2X2_3115 ( .A(u0_u5__abc_45296_n505), .B(u0_u5__abc_45296_n502), .Y(u0_u5_csc_18__FF_INPUT) );
  AND2X2 AND2X2_3116 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf0), .B(u0_u5__abc_45296_n333), .Y(u0_u5__abc_45296_n508) );
  AND2X2 AND2X2_3117 ( .A(u0_u5__abc_45296_n509), .B(u0_u5__abc_45296_n218_bF_buf4), .Y(u0_u5__abc_45296_n510) );
  AND2X2 AND2X2_3118 ( .A(u0_u5__abc_45296_n510), .B(u0_u5__abc_45296_n507), .Y(u0_u5_csc_19__FF_INPUT) );
  AND2X2 AND2X2_3119 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf6), .B(u0_u5__abc_45296_n339), .Y(u0_u5__abc_45296_n513) );
  AND2X2 AND2X2_312 ( .A(spec_req_cs_1_bF_buf0), .B(u0_tms1_14_), .Y(u0__abc_49347_n1537) );
  AND2X2 AND2X2_3120 ( .A(u0_u5__abc_45296_n514), .B(u0_u5__abc_45296_n218_bF_buf3), .Y(u0_u5__abc_45296_n515) );
  AND2X2 AND2X2_3121 ( .A(u0_u5__abc_45296_n515), .B(u0_u5__abc_45296_n512), .Y(u0_u5_csc_20__FF_INPUT) );
  AND2X2 AND2X2_3122 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf4), .B(u0_u5__abc_45296_n345), .Y(u0_u5__abc_45296_n518) );
  AND2X2 AND2X2_3123 ( .A(u0_u5__abc_45296_n519), .B(u0_u5__abc_45296_n218_bF_buf2), .Y(u0_u5__abc_45296_n520) );
  AND2X2 AND2X2_3124 ( .A(u0_u5__abc_45296_n520), .B(u0_u5__abc_45296_n517), .Y(u0_u5_csc_21__FF_INPUT) );
  AND2X2 AND2X2_3125 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf2), .B(u0_u5__abc_45296_n351), .Y(u0_u5__abc_45296_n523) );
  AND2X2 AND2X2_3126 ( .A(u0_u5__abc_45296_n524), .B(u0_u5__abc_45296_n218_bF_buf1), .Y(u0_u5__abc_45296_n525) );
  AND2X2 AND2X2_3127 ( .A(u0_u5__abc_45296_n525), .B(u0_u5__abc_45296_n522), .Y(u0_u5_csc_22__FF_INPUT) );
  AND2X2 AND2X2_3128 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf0), .B(u0_u5__abc_45296_n357), .Y(u0_u5__abc_45296_n528) );
  AND2X2 AND2X2_3129 ( .A(u0_u5__abc_45296_n529), .B(u0_u5__abc_45296_n218_bF_buf0), .Y(u0_u5__abc_45296_n530) );
  AND2X2 AND2X2_313 ( .A(u0__abc_49347_n1175_bF_buf5), .B(u0__abc_49347_n1540), .Y(u0__abc_49347_n1541) );
  AND2X2 AND2X2_3130 ( .A(u0_u5__abc_45296_n530), .B(u0_u5__abc_45296_n527), .Y(u0_u5_csc_23__FF_INPUT) );
  AND2X2 AND2X2_3131 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf6), .B(u0_u5__abc_45296_n363), .Y(u0_u5__abc_45296_n533) );
  AND2X2 AND2X2_3132 ( .A(u0_u5__abc_45296_n534), .B(u0_u5__abc_45296_n218_bF_buf7), .Y(u0_u5__abc_45296_n535) );
  AND2X2 AND2X2_3133 ( .A(u0_u5__abc_45296_n535), .B(u0_u5__abc_45296_n532), .Y(u0_u5_csc_24__FF_INPUT) );
  AND2X2 AND2X2_3134 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf4), .B(u0_u5__abc_45296_n369), .Y(u0_u5__abc_45296_n538) );
  AND2X2 AND2X2_3135 ( .A(u0_u5__abc_45296_n539), .B(u0_u5__abc_45296_n218_bF_buf6), .Y(u0_u5__abc_45296_n540) );
  AND2X2 AND2X2_3136 ( .A(u0_u5__abc_45296_n540), .B(u0_u5__abc_45296_n537), .Y(u0_u5_csc_25__FF_INPUT) );
  AND2X2 AND2X2_3137 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf2), .B(u0_u5__abc_45296_n375), .Y(u0_u5__abc_45296_n543) );
  AND2X2 AND2X2_3138 ( .A(u0_u5__abc_45296_n544), .B(u0_u5__abc_45296_n218_bF_buf5), .Y(u0_u5__abc_45296_n545) );
  AND2X2 AND2X2_3139 ( .A(u0_u5__abc_45296_n545), .B(u0_u5__abc_45296_n542), .Y(u0_u5_csc_26__FF_INPUT) );
  AND2X2 AND2X2_314 ( .A(u0__abc_49347_n1539), .B(u0__abc_49347_n1541), .Y(u0__abc_49347_n1542_1) );
  AND2X2 AND2X2_3140 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf0), .B(u0_u5__abc_45296_n381), .Y(u0_u5__abc_45296_n548) );
  AND2X2 AND2X2_3141 ( .A(u0_u5__abc_45296_n549), .B(u0_u5__abc_45296_n218_bF_buf4), .Y(u0_u5__abc_45296_n550) );
  AND2X2 AND2X2_3142 ( .A(u0_u5__abc_45296_n550), .B(u0_u5__abc_45296_n547), .Y(u0_u5_csc_27__FF_INPUT) );
  AND2X2 AND2X2_3143 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf6), .B(u0_u5__abc_45296_n387), .Y(u0_u5__abc_45296_n553) );
  AND2X2 AND2X2_3144 ( .A(u0_u5__abc_45296_n554), .B(u0_u5__abc_45296_n218_bF_buf3), .Y(u0_u5__abc_45296_n555) );
  AND2X2 AND2X2_3145 ( .A(u0_u5__abc_45296_n555), .B(u0_u5__abc_45296_n552), .Y(u0_u5_csc_28__FF_INPUT) );
  AND2X2 AND2X2_3146 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf4), .B(u0_u5__abc_45296_n393), .Y(u0_u5__abc_45296_n558) );
  AND2X2 AND2X2_3147 ( .A(u0_u5__abc_45296_n559), .B(u0_u5__abc_45296_n218_bF_buf2), .Y(u0_u5__abc_45296_n560) );
  AND2X2 AND2X2_3148 ( .A(u0_u5__abc_45296_n560), .B(u0_u5__abc_45296_n557), .Y(u0_u5_csc_29__FF_INPUT) );
  AND2X2 AND2X2_3149 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf2), .B(u0_u5__abc_45296_n399), .Y(u0_u5__abc_45296_n563) );
  AND2X2 AND2X2_315 ( .A(u0__abc_49347_n1176_1_bF_buf5), .B(sp_tms_15_), .Y(u0__abc_49347_n1544) );
  AND2X2 AND2X2_3150 ( .A(u0_u5__abc_45296_n564), .B(u0_u5__abc_45296_n218_bF_buf1), .Y(u0_u5__abc_45296_n565) );
  AND2X2 AND2X2_3151 ( .A(u0_u5__abc_45296_n565), .B(u0_u5__abc_45296_n562), .Y(u0_u5_csc_30__FF_INPUT) );
  AND2X2 AND2X2_3152 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf0), .B(u0_u5__abc_45296_n405), .Y(u0_u5__abc_45296_n568) );
  AND2X2 AND2X2_3153 ( .A(u0_u5__abc_45296_n569), .B(u0_u5__abc_45296_n218_bF_buf0), .Y(u0_u5__abc_45296_n570) );
  AND2X2 AND2X2_3154 ( .A(u0_u5__abc_45296_n570), .B(u0_u5__abc_45296_n567), .Y(u0_u5_csc_31__FF_INPUT) );
  AND2X2 AND2X2_3155 ( .A(u0_csc5_8_), .B(wb_we_i), .Y(u0_u5__abc_45296_n572) );
  AND2X2 AND2X2_3156 ( .A(u0_csc5_20_), .B(u0_csc_mask_4_), .Y(u0_u5__abc_45296_n573) );
  AND2X2 AND2X2_3157 ( .A(u0_csc_mask_4_), .B(wb_addr_i_25_bF_buf1), .Y(u0_u5__abc_45296_n574) );
  AND2X2 AND2X2_3158 ( .A(u0_csc_mask_3_), .B(\wb_addr_i[24] ), .Y(u0_u5__abc_45296_n577) );
  AND2X2 AND2X2_3159 ( .A(u0_csc5_19_), .B(u0_csc_mask_3_), .Y(u0_u5__abc_45296_n578) );
  AND2X2 AND2X2_316 ( .A(spec_req_cs_5_bF_buf5), .B(u0_tms5_15_), .Y(u0__abc_49347_n1545) );
  AND2X2 AND2X2_3160 ( .A(u0_u5__abc_45296_n576), .B(u0_u5__abc_45296_n580), .Y(u0_u5__abc_45296_n581) );
  AND2X2 AND2X2_3161 ( .A(u0_csc5_18_), .B(u0_csc_mask_2_), .Y(u0_u5__abc_45296_n583) );
  AND2X2 AND2X2_3162 ( .A(u0_u5__abc_45296_n583), .B(u0_u5__abc_45296_n582), .Y(u0_u5__abc_45296_n584) );
  AND2X2 AND2X2_3163 ( .A(u0_u5__abc_45296_n587), .B(u0_u5__abc_45296_n585), .Y(u0_u5__abc_45296_n588) );
  AND2X2 AND2X2_3164 ( .A(u0_u5__abc_45296_n581), .B(u0_u5__abc_45296_n588), .Y(u0_u5__abc_45296_n589) );
  AND2X2 AND2X2_3165 ( .A(u0_csc5_22_), .B(u0_csc_mask_6_), .Y(u0_u5__abc_45296_n590) );
  AND2X2 AND2X2_3166 ( .A(u0_csc_mask_6_), .B(\wb_addr_i[27] ), .Y(u0_u5__abc_45296_n591) );
  AND2X2 AND2X2_3167 ( .A(u0_csc_mask_5_), .B(\wb_addr_i[26] ), .Y(u0_u5__abc_45296_n594) );
  AND2X2 AND2X2_3168 ( .A(u0_csc5_21_), .B(u0_csc_mask_5_), .Y(u0_u5__abc_45296_n595) );
  AND2X2 AND2X2_3169 ( .A(u0_u5__abc_45296_n593), .B(u0_u5__abc_45296_n597), .Y(u0_u5__abc_45296_n598) );
  AND2X2 AND2X2_317 ( .A(u0__abc_49347_n1547), .B(u0__abc_49347_n1185_bF_buf2), .Y(u0__abc_49347_n1548) );
  AND2X2 AND2X2_3170 ( .A(u0_u5__abc_45296_n573), .B(u0_u5__abc_45296_n599), .Y(u0_u5__abc_45296_n600) );
  AND2X2 AND2X2_3171 ( .A(u0_u5__abc_45296_n603), .B(u0_u5__abc_45296_n601), .Y(u0_u5__abc_45296_n604) );
  AND2X2 AND2X2_3172 ( .A(u0_u5__abc_45296_n598), .B(u0_u5__abc_45296_n604), .Y(u0_u5__abc_45296_n605) );
  AND2X2 AND2X2_3173 ( .A(u0_u5__abc_45296_n589), .B(u0_u5__abc_45296_n605), .Y(u0_u5__abc_45296_n606) );
  AND2X2 AND2X2_3174 ( .A(u0_u5__abc_45296_n592), .B(u0_u5__abc_45296_n590), .Y(u0_u5__abc_45296_n607) );
  AND2X2 AND2X2_3175 ( .A(u0_csc_mask_7_), .B(\wb_addr_i[28] ), .Y(u0_u5__abc_45296_n609) );
  AND2X2 AND2X2_3176 ( .A(u0_csc5_23_), .B(u0_csc_mask_7_), .Y(u0_u5__abc_45296_n611) );
  AND2X2 AND2X2_3177 ( .A(u0_u5__abc_45296_n608), .B(u0_u5__abc_45296_n612), .Y(u0_u5__abc_45296_n613) );
  AND2X2 AND2X2_3178 ( .A(u0_u5__abc_45296_n613), .B(u0_u5__abc_45296_n615), .Y(u0_u5__abc_45296_n616) );
  AND2X2 AND2X2_3179 ( .A(u0_u5__abc_45296_n606), .B(u0_u5__abc_45296_n616), .Y(u0_u5__abc_45296_n617) );
  AND2X2 AND2X2_318 ( .A(u0__abc_49347_n1548), .B(u0__abc_49347_n1546), .Y(u0__abc_49347_n1549) );
  AND2X2 AND2X2_3180 ( .A(u0_csc_mask_2_), .B(wb_addr_i_23_bF_buf0), .Y(u0_u5__abc_45296_n618) );
  AND2X2 AND2X2_3181 ( .A(u0_csc_mask_1_), .B(\wb_addr_i[22] ), .Y(u0_u5__abc_45296_n621) );
  AND2X2 AND2X2_3182 ( .A(u0_csc5_17_), .B(u0_csc_mask_1_), .Y(u0_u5__abc_45296_n622) );
  AND2X2 AND2X2_3183 ( .A(u0_u5__abc_45296_n620), .B(u0_u5__abc_45296_n624), .Y(u0_u5__abc_45296_n625) );
  AND2X2 AND2X2_3184 ( .A(u0_csc_mask_0_), .B(\wb_addr_i[21] ), .Y(u0_u5__abc_45296_n626) );
  AND2X2 AND2X2_3185 ( .A(u0_csc5_16_), .B(u0_csc_mask_0_), .Y(u0_u5__abc_45296_n627) );
  AND2X2 AND2X2_3186 ( .A(u0_u5__abc_45296_n629), .B(u0_u5__abc_45296_n631), .Y(u0_u5__abc_45296_n632) );
  AND2X2 AND2X2_3187 ( .A(u0_u5__abc_45296_n625), .B(u0_u5__abc_45296_n632), .Y(u0_u5__abc_45296_n633) );
  AND2X2 AND2X2_3188 ( .A(u0_u5__abc_45296_n635), .B(u0_csc5_0_), .Y(u0_u5__abc_45296_n636) );
  AND2X2 AND2X2_3189 ( .A(u0_u5__abc_45296_n633), .B(u0_u5__abc_45296_n636), .Y(u0_u5__abc_45296_n637) );
  AND2X2 AND2X2_319 ( .A(u0__abc_49347_n1550), .B(u0__abc_49347_n1181_bF_buf2), .Y(u0__abc_49347_n1551_1) );
  AND2X2 AND2X2_3190 ( .A(u0_u5__abc_45296_n617), .B(u0_u5__abc_45296_n637), .Y(u0_u5__abc_45296_n638) );
  AND2X2 AND2X2_3191 ( .A(u0_u5__abc_45296_n638), .B(u0_u5__abc_45296_n572), .Y(u0_u5_wp_err) );
  AND2X2 AND2X2_3192 ( .A(u0_u5__abc_45296_n638), .B(u0_u5__abc_45296_n640), .Y(u0_cs5) );
  AND2X2 AND2X2_3193 ( .A(u0_u5__abc_45296_n643), .B(u0_init_req5), .Y(u0_u5__abc_45296_n644) );
  AND2X2 AND2X2_3194 ( .A(u0_u5__abc_45296_n645), .B(u0_csc5_0_), .Y(u0_u5__abc_45296_n646) );
  AND2X2 AND2X2_3195 ( .A(u0_u5__abc_45296_n646), .B(u0_u5_init_req_we), .Y(u0_u5__abc_45296_n647) );
  AND2X2 AND2X2_3196 ( .A(u0_u5__abc_45296_n203), .B(u0_u5__abc_45296_n647), .Y(u0_u5__abc_45296_n648) );
  AND2X2 AND2X2_3197 ( .A(u1__abc_45852_n258_1), .B(csc_s_6_), .Y(u1__abc_45852_n259_1) );
  AND2X2 AND2X2_3198 ( .A(u1__abc_45852_n261_bF_buf4), .B(u1__abc_45852_n259_1), .Y(u1__abc_45852_n262_1) );
  AND2X2 AND2X2_3199 ( .A(u1__abc_45852_n263), .B(csc_s_7_), .Y(u1__abc_45852_n264) );
  AND2X2 AND2X2_32 ( .A(_abc_55805_n332), .B(_abc_55805_n333), .Y(tms_s_14_) );
  AND2X2 AND2X2_320 ( .A(spec_req_cs_4_bF_buf5), .B(u0_tms4_15_), .Y(u0__abc_49347_n1552_1) );
  AND2X2 AND2X2_3200 ( .A(u1__abc_45852_n261_bF_buf3), .B(u1__abc_45852_n264), .Y(u1__abc_45852_n265_1) );
  AND2X2 AND2X2_3201 ( .A(u1__abc_45852_n271_1), .B(u1__abc_45852_n273_1), .Y(u1__abc_45852_n274) );
  AND2X2 AND2X2_3202 ( .A(u1__abc_45852_n275), .B(csc_s_4_), .Y(u1__abc_45852_n276) );
  AND2X2 AND2X2_3203 ( .A(u1__abc_45852_n264), .B(u1__abc_45852_n276_bF_buf4), .Y(u1__abc_45852_n277) );
  AND2X2 AND2X2_3204 ( .A(u1__abc_45852_n274), .B(u1__abc_45852_n278_1), .Y(u1__abc_45852_n279_1) );
  AND2X2 AND2X2_3205 ( .A(u1__abc_45852_n279_1), .B(u1__abc_45852_n267_1), .Y(page_size_8_) );
  AND2X2 AND2X2_3206 ( .A(u1__abc_45852_n281), .B(bank_adr_0_bF_buf3), .Y(u1__abc_45852_n282) );
  AND2X2 AND2X2_3207 ( .A(page_size_8_), .B(\wb_addr_i[10] ), .Y(u1__abc_45852_n283) );
  AND2X2 AND2X2_3208 ( .A(page_size_9_), .B(\wb_addr_i[11] ), .Y(u1__abc_45852_n285_1) );
  AND2X2 AND2X2_3209 ( .A(page_size_10_bF_buf2), .B(\wb_addr_i[12] ), .Y(u1__abc_45852_n286_1) );
  AND2X2 AND2X2_321 ( .A(u0__abc_49347_n1553), .B(u0__abc_49347_n1180_1_bF_buf2), .Y(u0__abc_49347_n1554) );
  AND2X2 AND2X2_3210 ( .A(u1__abc_45852_n269), .B(csc_s_5_bF_buf1), .Y(u1__abc_45852_n292_1) );
  AND2X2 AND2X2_3211 ( .A(u1__abc_45852_n291), .B(u1__abc_45852_n292_1), .Y(u1__abc_45852_n293_1) );
  AND2X2 AND2X2_3212 ( .A(u1__abc_45852_n259_1), .B(u1__abc_45852_n292_1), .Y(u1__abc_45852_n294_1) );
  AND2X2 AND2X2_3213 ( .A(u1__abc_45852_n291), .B(u1__abc_45852_n276_bF_buf3), .Y(u1__abc_45852_n295) );
  AND2X2 AND2X2_3214 ( .A(u1__abc_45852_n267_1), .B(u1__abc_45852_n278_1), .Y(u1__abc_45852_n299_1) );
  AND2X2 AND2X2_3215 ( .A(u1__abc_45852_n298), .B(u1__abc_45852_n299_1), .Y(u1__abc_45852_n300_1) );
  AND2X2 AND2X2_3216 ( .A(u1__abc_45852_n300_1), .B(wb_addr_i_23_bF_buf3), .Y(u1__abc_45852_n301_1) );
  AND2X2 AND2X2_3217 ( .A(u1__abc_45852_n296), .B(\wb_addr_i[22] ), .Y(u1__abc_45852_n302) );
  AND2X2 AND2X2_3218 ( .A(u1__abc_45852_n303), .B(\wb_addr_i[24] ), .Y(u1__abc_45852_n304) );
  AND2X2 AND2X2_3219 ( .A(u1__abc_45852_n265_1), .B(wb_addr_i_25_bF_buf3), .Y(u1__abc_45852_n305) );
  AND2X2 AND2X2_322 ( .A(spec_req_cs_3_bF_buf5), .B(u0_tms3_15_), .Y(u0__abc_49347_n1555) );
  AND2X2 AND2X2_3220 ( .A(u1__abc_45852_n293_1), .B(\wb_addr_i[21] ), .Y(u1__abc_45852_n306_1) );
  AND2X2 AND2X2_3221 ( .A(u1__abc_45852_n311), .B(cs_le_bF_buf3), .Y(u1__abc_45852_n312) );
  AND2X2 AND2X2_3222 ( .A(u1__abc_45852_n312), .B(u1__abc_45852_n289), .Y(u1__abc_45852_n313_1) );
  AND2X2 AND2X2_3223 ( .A(u1__abc_45852_n281), .B(bank_adr_1_bF_buf3), .Y(u1__abc_45852_n315_1) );
  AND2X2 AND2X2_3224 ( .A(page_size_8_), .B(\wb_addr_i[11] ), .Y(u1__abc_45852_n316) );
  AND2X2 AND2X2_3225 ( .A(page_size_9_), .B(\wb_addr_i[12] ), .Y(u1__abc_45852_n317) );
  AND2X2 AND2X2_3226 ( .A(page_size_10_bF_buf1), .B(\wb_addr_i[13] ), .Y(u1__abc_45852_n318) );
  AND2X2 AND2X2_3227 ( .A(u1__abc_45852_n300_1), .B(\wb_addr_i[24] ), .Y(u1__abc_45852_n322_1) );
  AND2X2 AND2X2_3228 ( .A(u1__abc_45852_n303), .B(wb_addr_i_25_bF_buf2), .Y(u1__abc_45852_n323) );
  AND2X2 AND2X2_3229 ( .A(u1__abc_45852_n296), .B(wb_addr_i_23_bF_buf2), .Y(u1__abc_45852_n324) );
  AND2X2 AND2X2_323 ( .A(u0__abc_49347_n1556), .B(u0__abc_49347_n1179_bF_buf2), .Y(u0__abc_49347_n1557) );
  AND2X2 AND2X2_3230 ( .A(u1__abc_45852_n265_1), .B(\wb_addr_i[26] ), .Y(u1__abc_45852_n325) );
  AND2X2 AND2X2_3231 ( .A(u1__abc_45852_n293_1), .B(\wb_addr_i[22] ), .Y(u1__abc_45852_n326) );
  AND2X2 AND2X2_3232 ( .A(u1__abc_45852_n331), .B(cs_le_bF_buf2), .Y(u1__abc_45852_n332) );
  AND2X2 AND2X2_3233 ( .A(u1__abc_45852_n332), .B(u1__abc_45852_n321_1), .Y(u1__abc_45852_n333_1) );
  AND2X2 AND2X2_3234 ( .A(u1__abc_45852_n281), .B(row_adr_0_bF_buf6), .Y(u1__abc_45852_n335_1) );
  AND2X2 AND2X2_3235 ( .A(page_size_8_), .B(\wb_addr_i[12] ), .Y(u1__abc_45852_n336) );
  AND2X2 AND2X2_3236 ( .A(page_size_10_bF_buf0), .B(\wb_addr_i[14] ), .Y(u1__abc_45852_n337) );
  AND2X2 AND2X2_3237 ( .A(page_size_9_), .B(\wb_addr_i[13] ), .Y(u1__abc_45852_n338) );
  AND2X2 AND2X2_3238 ( .A(u1__abc_45852_n342), .B(cs_le_bF_buf1), .Y(u1__abc_45852_n343) );
  AND2X2 AND2X2_3239 ( .A(u1__abc_45852_n343), .B(u1__abc_45852_n341_1), .Y(u1__abc_45852_n344) );
  AND2X2 AND2X2_324 ( .A(spec_req_cs_2_bF_buf5), .B(u0_tms2_15_), .Y(u0__abc_49347_n1558) );
  AND2X2 AND2X2_3240 ( .A(u1__abc_45852_n281), .B(row_adr_1_bF_buf6), .Y(u1__abc_45852_n346_1) );
  AND2X2 AND2X2_3241 ( .A(page_size_8_), .B(\wb_addr_i[13] ), .Y(u1__abc_45852_n347_1) );
  AND2X2 AND2X2_3242 ( .A(page_size_10_bF_buf3), .B(\wb_addr_i[15] ), .Y(u1__abc_45852_n348) );
  AND2X2 AND2X2_3243 ( .A(page_size_9_), .B(\wb_addr_i[14] ), .Y(u1__abc_45852_n349) );
  AND2X2 AND2X2_3244 ( .A(u1__abc_45852_n353_1), .B(cs_le_bF_buf0), .Y(u1__abc_45852_n354) );
  AND2X2 AND2X2_3245 ( .A(u1__abc_45852_n354), .B(u1__abc_45852_n352_1), .Y(u1__abc_45852_n355) );
  AND2X2 AND2X2_3246 ( .A(u1__abc_45852_n281), .B(row_adr_2_bF_buf6), .Y(u1__abc_45852_n357_1) );
  AND2X2 AND2X2_3247 ( .A(page_size_8_), .B(u1__abc_45852_n298), .Y(u1__abc_45852_n358_1) );
  AND2X2 AND2X2_3248 ( .A(u1__abc_45852_n358_1), .B(\wb_addr_i[14] ), .Y(u1__abc_45852_n359_1) );
  AND2X2 AND2X2_3249 ( .A(u1__abc_45852_n296), .B(\wb_addr_i[14] ), .Y(u1__abc_45852_n360) );
  AND2X2 AND2X2_325 ( .A(u0__abc_49347_n1559), .B(u0__abc_49347_n1178_1_bF_buf2), .Y(u0__abc_49347_n1560_1) );
  AND2X2 AND2X2_3250 ( .A(u1__abc_45852_n259_1), .B(u1__abc_45852_n276_bF_buf2), .Y(u1__abc_45852_n361) );
  AND2X2 AND2X2_3251 ( .A(u1__abc_45852_n363_1), .B(\wb_addr_i[15] ), .Y(u1__abc_45852_n364_1) );
  AND2X2 AND2X2_3252 ( .A(page_size_10_bF_buf2), .B(\wb_addr_i[16] ), .Y(u1__abc_45852_n366) );
  AND2X2 AND2X2_3253 ( .A(u1__abc_45852_n293_1), .B(\wb_addr_i[14] ), .Y(u1__abc_45852_n367) );
  AND2X2 AND2X2_3254 ( .A(u1__abc_45852_n277), .B(\wb_addr_i[15] ), .Y(u1__abc_45852_n368) );
  AND2X2 AND2X2_3255 ( .A(u1__abc_45852_n374), .B(cs_le_bF_buf4), .Y(u1__abc_45852_n375_1) );
  AND2X2 AND2X2_3256 ( .A(u1__abc_45852_n375_1), .B(u1__abc_45852_n373), .Y(u1__abc_45852_n376_1) );
  AND2X2 AND2X2_3257 ( .A(u1__abc_45852_n281), .B(row_adr_3_bF_buf6), .Y(u1__abc_45852_n378) );
  AND2X2 AND2X2_3258 ( .A(u1__abc_45852_n358_1), .B(\wb_addr_i[15] ), .Y(u1__abc_45852_n379) );
  AND2X2 AND2X2_3259 ( .A(page_size_9_), .B(\wb_addr_i[16] ), .Y(u1__abc_45852_n380) );
  AND2X2 AND2X2_326 ( .A(spec_req_cs_1_bF_buf5), .B(u0_tms1_15_), .Y(u0__abc_49347_n1561_1) );
  AND2X2 AND2X2_3260 ( .A(page_size_10_bF_buf1), .B(\wb_addr_i[17] ), .Y(u1__abc_45852_n381_1) );
  AND2X2 AND2X2_3261 ( .A(u1__abc_45852_n297), .B(\wb_addr_i[15] ), .Y(u1__abc_45852_n382_1) );
  AND2X2 AND2X2_3262 ( .A(u1__abc_45852_n387_1), .B(cs_le_bF_buf3), .Y(u1__abc_45852_n388_1) );
  AND2X2 AND2X2_3263 ( .A(u1__abc_45852_n388_1), .B(u1__abc_45852_n386), .Y(u1__abc_45852_n389_1) );
  AND2X2 AND2X2_3264 ( .A(u1__abc_45852_n281), .B(row_adr_4_bF_buf6), .Y(u1__abc_45852_n391) );
  AND2X2 AND2X2_3265 ( .A(u1__abc_45852_n358_1), .B(\wb_addr_i[16] ), .Y(u1__abc_45852_n392) );
  AND2X2 AND2X2_3266 ( .A(u1__abc_45852_n296), .B(\wb_addr_i[16] ), .Y(u1__abc_45852_n393_1) );
  AND2X2 AND2X2_3267 ( .A(u1__abc_45852_n363_1), .B(\wb_addr_i[17] ), .Y(u1__abc_45852_n394_1) );
  AND2X2 AND2X2_3268 ( .A(page_size_10_bF_buf0), .B(\wb_addr_i[18] ), .Y(u1__abc_45852_n396) );
  AND2X2 AND2X2_3269 ( .A(u1__abc_45852_n293_1), .B(\wb_addr_i[16] ), .Y(u1__abc_45852_n397) );
  AND2X2 AND2X2_327 ( .A(u0__abc_49347_n1175_bF_buf4), .B(u0__abc_49347_n1564), .Y(u0__abc_49347_n1565) );
  AND2X2 AND2X2_3270 ( .A(u1__abc_45852_n277), .B(\wb_addr_i[17] ), .Y(u1__abc_45852_n398) );
  AND2X2 AND2X2_3271 ( .A(u1__abc_45852_n404), .B(cs_le_bF_buf2), .Y(u1__abc_45852_n405_1) );
  AND2X2 AND2X2_3272 ( .A(u1__abc_45852_n405_1), .B(u1__abc_45852_n403), .Y(u1__abc_45852_n406_1) );
  AND2X2 AND2X2_3273 ( .A(u1__abc_45852_n281), .B(row_adr_5_bF_buf6), .Y(u1__abc_45852_n408) );
  AND2X2 AND2X2_3274 ( .A(u1__abc_45852_n358_1), .B(\wb_addr_i[17] ), .Y(u1__abc_45852_n410) );
  AND2X2 AND2X2_3275 ( .A(u1__abc_45852_n296), .B(\wb_addr_i[17] ), .Y(u1__abc_45852_n411_1) );
  AND2X2 AND2X2_3276 ( .A(u1__abc_45852_n363_1), .B(\wb_addr_i[18] ), .Y(u1__abc_45852_n412_1) );
  AND2X2 AND2X2_3277 ( .A(page_size_10_bF_buf3), .B(\wb_addr_i[19] ), .Y(u1__abc_45852_n414) );
  AND2X2 AND2X2_3278 ( .A(u1__abc_45852_n293_1), .B(\wb_addr_i[17] ), .Y(u1__abc_45852_n415) );
  AND2X2 AND2X2_3279 ( .A(u1__abc_45852_n277), .B(\wb_addr_i[18] ), .Y(u1__abc_45852_n416) );
  AND2X2 AND2X2_328 ( .A(u0__abc_49347_n1563), .B(u0__abc_49347_n1565), .Y(u0__abc_49347_n1566) );
  AND2X2 AND2X2_3280 ( .A(u1__abc_45852_n421_1), .B(cs_le_bF_buf1), .Y(u1__abc_45852_n422_1) );
  AND2X2 AND2X2_3281 ( .A(u1__abc_45852_n422_1), .B(u1__abc_45852_n409), .Y(u1__abc_45852_n423_1) );
  AND2X2 AND2X2_3282 ( .A(u1__abc_45852_n281), .B(row_adr_6_bF_buf6), .Y(u1__abc_45852_n425_1) );
  AND2X2 AND2X2_3283 ( .A(page_size_8_), .B(\wb_addr_i[18] ), .Y(u1__abc_45852_n426_1) );
  AND2X2 AND2X2_3284 ( .A(page_size_10_bF_buf2), .B(\wb_addr_i[20] ), .Y(u1__abc_45852_n427_1) );
  AND2X2 AND2X2_3285 ( .A(page_size_9_), .B(\wb_addr_i[19] ), .Y(u1__abc_45852_n428_1) );
  AND2X2 AND2X2_3286 ( .A(u1__abc_45852_n432_1), .B(cs_le_bF_buf0), .Y(u1__abc_45852_n433_1) );
  AND2X2 AND2X2_3287 ( .A(u1__abc_45852_n433_1), .B(u1__abc_45852_n431_1), .Y(u1__abc_45852_n434_1) );
  AND2X2 AND2X2_3288 ( .A(u1__abc_45852_n281), .B(row_adr_7_bF_buf6), .Y(u1__abc_45852_n436_1) );
  AND2X2 AND2X2_3289 ( .A(page_size_8_), .B(\wb_addr_i[19] ), .Y(u1__abc_45852_n438_1) );
  AND2X2 AND2X2_329 ( .A(u0__abc_49347_n1176_1_bF_buf4), .B(sp_tms_16_), .Y(u0__abc_49347_n1568) );
  AND2X2 AND2X2_3290 ( .A(page_size_10_bF_buf1), .B(\wb_addr_i[21] ), .Y(u1__abc_45852_n439_1) );
  AND2X2 AND2X2_3291 ( .A(page_size_9_), .B(\wb_addr_i[20] ), .Y(u1__abc_45852_n440_1) );
  AND2X2 AND2X2_3292 ( .A(u1__abc_45852_n443_1), .B(cs_le_bF_buf4), .Y(u1__abc_45852_n444_1) );
  AND2X2 AND2X2_3293 ( .A(u1__abc_45852_n444_1), .B(u1__abc_45852_n437_1), .Y(u1__abc_45852_n445_1) );
  AND2X2 AND2X2_3294 ( .A(u1__abc_45852_n281), .B(row_adr_8_bF_buf6), .Y(u1__abc_45852_n447_1) );
  AND2X2 AND2X2_3295 ( .A(u1__abc_45852_n358_1), .B(\wb_addr_i[20] ), .Y(u1__abc_45852_n448_1) );
  AND2X2 AND2X2_3296 ( .A(page_size_9_), .B(\wb_addr_i[21] ), .Y(u1__abc_45852_n449_1) );
  AND2X2 AND2X2_3297 ( .A(page_size_10_bF_buf0), .B(\wb_addr_i[22] ), .Y(u1__abc_45852_n450_1) );
  AND2X2 AND2X2_3298 ( .A(u1__abc_45852_n297), .B(\wb_addr_i[20] ), .Y(u1__abc_45852_n451_1) );
  AND2X2 AND2X2_3299 ( .A(u1__abc_45852_n456_1), .B(cs_le_bF_buf3), .Y(u1__abc_45852_n457_1) );
  AND2X2 AND2X2_33 ( .A(_abc_55805_n335), .B(_abc_55805_n336), .Y(tms_s_15_) );
  AND2X2 AND2X2_330 ( .A(spec_req_cs_5_bF_buf4), .B(u0_tms5_16_), .Y(u0__abc_49347_n1569_1) );
  AND2X2 AND2X2_3300 ( .A(u1__abc_45852_n457_1), .B(u1__abc_45852_n455_1), .Y(u1__abc_45852_n458_1) );
  AND2X2 AND2X2_3301 ( .A(u1__abc_45852_n281), .B(row_adr_9_bF_buf6), .Y(u1__abc_45852_n460_1) );
  AND2X2 AND2X2_3302 ( .A(u1__abc_45852_n358_1), .B(\wb_addr_i[21] ), .Y(u1__abc_45852_n462_1) );
  AND2X2 AND2X2_3303 ( .A(page_size_9_), .B(\wb_addr_i[22] ), .Y(u1__abc_45852_n463_1) );
  AND2X2 AND2X2_3304 ( .A(page_size_10_bF_buf3), .B(wb_addr_i_23_bF_buf1), .Y(u1__abc_45852_n464_1) );
  AND2X2 AND2X2_3305 ( .A(u1__abc_45852_n296), .B(\wb_addr_i[21] ), .Y(u1__abc_45852_n465_1) );
  AND2X2 AND2X2_3306 ( .A(u1__abc_45852_n470_1), .B(cs_le_bF_buf2), .Y(u1__abc_45852_n471) );
  AND2X2 AND2X2_3307 ( .A(u1__abc_45852_n471), .B(u1__abc_45852_n461_1), .Y(u1__abc_45852_n472_1) );
  AND2X2 AND2X2_3308 ( .A(u1__abc_45852_n281), .B(row_adr_10_bF_buf6), .Y(u1__abc_45852_n474_1) );
  AND2X2 AND2X2_3309 ( .A(u1__abc_45852_n358_1), .B(\wb_addr_i[22] ), .Y(u1__abc_45852_n476_1) );
  AND2X2 AND2X2_331 ( .A(u0__abc_49347_n1571), .B(u0__abc_49347_n1185_bF_buf1), .Y(u0__abc_49347_n1572) );
  AND2X2 AND2X2_3310 ( .A(u1__abc_45852_n276_bF_buf1), .B(wb_addr_i_23_bF_buf0), .Y(u1__abc_45852_n477_1) );
  AND2X2 AND2X2_3311 ( .A(u1__abc_45852_n477_1), .B(u1__abc_45852_n264), .Y(u1__abc_45852_n478) );
  AND2X2 AND2X2_3312 ( .A(u1__abc_45852_n363_1), .B(wb_addr_i_23_bF_buf3), .Y(u1__abc_45852_n481) );
  AND2X2 AND2X2_3313 ( .A(page_size_10_bF_buf2), .B(\wb_addr_i[24] ), .Y(u1__abc_45852_n483_1) );
  AND2X2 AND2X2_3314 ( .A(u1__abc_45852_n486), .B(cs_le_bF_buf1), .Y(u1__abc_45852_n487) );
  AND2X2 AND2X2_3315 ( .A(u1__abc_45852_n487), .B(u1__abc_45852_n475), .Y(u1__abc_45852_n488_1) );
  AND2X2 AND2X2_3316 ( .A(u1__abc_45852_n281), .B(row_adr_11_bF_buf6), .Y(u1__abc_45852_n490_1) );
  AND2X2 AND2X2_3317 ( .A(u1__abc_45852_n358_1), .B(wb_addr_i_23_bF_buf2), .Y(u1__abc_45852_n493) );
  AND2X2 AND2X2_3318 ( .A(page_size_9_), .B(\wb_addr_i[24] ), .Y(u1__abc_45852_n494_1) );
  AND2X2 AND2X2_3319 ( .A(page_size_10_bF_buf1), .B(wb_addr_i_25_bF_buf1), .Y(u1__abc_45852_n495) );
  AND2X2 AND2X2_332 ( .A(u0__abc_49347_n1572), .B(u0__abc_49347_n1570_1), .Y(u0__abc_49347_n1573) );
  AND2X2 AND2X2_3320 ( .A(u1__abc_45852_n499), .B(cs_le_bF_buf0), .Y(u1__abc_45852_n500_1) );
  AND2X2 AND2X2_3321 ( .A(u1__abc_45852_n500_1), .B(u1__abc_45852_n492), .Y(u1__abc_45852_n501) );
  AND2X2 AND2X2_3322 ( .A(u1__abc_45852_n281), .B(row_adr_12_bF_buf6), .Y(u1__abc_45852_n503) );
  AND2X2 AND2X2_3323 ( .A(u1__abc_45852_n265_1), .B(\wb_addr_i[24] ), .Y(u1__abc_45852_n504) );
  AND2X2 AND2X2_3324 ( .A(u1__abc_45852_n358_1), .B(\wb_addr_i[24] ), .Y(u1__abc_45852_n508_1) );
  AND2X2 AND2X2_3325 ( .A(u1__abc_45852_n277), .B(wb_addr_i_25_bF_buf0), .Y(u1__abc_45852_n509) );
  AND2X2 AND2X2_3326 ( .A(u1__abc_45852_n512_1), .B(cs_le_bF_buf4), .Y(u1__abc_45852_n513) );
  AND2X2 AND2X2_3327 ( .A(u1__abc_45852_n513), .B(u1__abc_45852_n507), .Y(u1__abc_45852_n514_1) );
  AND2X2 AND2X2_3328 ( .A(u1__abc_45852_n516), .B(wb_stb_i_bF_buf3), .Y(u1__abc_45852_n517) );
  AND2X2 AND2X2_3329 ( .A(mem_ack_r), .B(u1_wr_cycle), .Y(u1__abc_45852_n518_1) );
  AND2X2 AND2X2_333 ( .A(u0__abc_49347_n1574), .B(u0__abc_49347_n1181_bF_buf1), .Y(u0__abc_49347_n1575) );
  AND2X2 AND2X2_3330 ( .A(u1__abc_45852_n521), .B(u1__abc_45852_n522), .Y(u1_col_adr_0__FF_INPUT) );
  AND2X2 AND2X2_3331 ( .A(u1__abc_45852_n524_1), .B(u1__abc_45852_n525), .Y(u1_col_adr_1__FF_INPUT) );
  AND2X2 AND2X2_3332 ( .A(u1__abc_45852_n527), .B(u1__abc_45852_n528), .Y(u1_col_adr_2__FF_INPUT) );
  AND2X2 AND2X2_3333 ( .A(u1__abc_45852_n530_1), .B(u1__abc_45852_n531), .Y(u1_col_adr_3__FF_INPUT) );
  AND2X2 AND2X2_3334 ( .A(u1__abc_45852_n533), .B(u1__abc_45852_n534), .Y(u1_col_adr_4__FF_INPUT) );
  AND2X2 AND2X2_3335 ( .A(u1__abc_45852_n536_1), .B(u1__abc_45852_n537), .Y(u1_col_adr_5__FF_INPUT) );
  AND2X2 AND2X2_3336 ( .A(u1__abc_45852_n539), .B(u1__abc_45852_n540), .Y(u1_col_adr_6__FF_INPUT) );
  AND2X2 AND2X2_3337 ( .A(u1__abc_45852_n542_1), .B(u1__abc_45852_n543), .Y(u1_col_adr_7__FF_INPUT) );
  AND2X2 AND2X2_3338 ( .A(u1__abc_45852_n520_1), .B(u1_col_adr_8_), .Y(u1__abc_45852_n545) );
  AND2X2 AND2X2_3339 ( .A(u1__abc_45852_n519), .B(\wb_addr_i[10] ), .Y(u1__abc_45852_n547) );
  AND2X2 AND2X2_334 ( .A(spec_req_cs_4_bF_buf4), .B(u0_tms4_16_), .Y(u0__abc_49347_n1576) );
  AND2X2 AND2X2_3340 ( .A(u1__abc_45852_n546), .B(u1__abc_45852_n547), .Y(u1__abc_45852_n548_1) );
  AND2X2 AND2X2_3341 ( .A(u1__abc_45852_n520_1), .B(u1_col_adr_9_), .Y(u1__abc_45852_n550_1) );
  AND2X2 AND2X2_3342 ( .A(u1__abc_45852_n519), .B(\wb_addr_i[11] ), .Y(u1__abc_45852_n551) );
  AND2X2 AND2X2_3343 ( .A(page_size_10_bF_buf0), .B(u1__abc_45852_n551), .Y(u1__abc_45852_n552) );
  AND2X2 AND2X2_3344 ( .A(u1__abc_45852_n557_1), .B(u1__abc_45852_n555), .Y(u1__abc_45852_n558) );
  AND2X2 AND2X2_3345 ( .A(u1__abc_45852_n276_bF_buf0), .B(\wb_addr_i[1] ), .Y(u1__abc_45852_n560_1) );
  AND2X2 AND2X2_3346 ( .A(u1__abc_45852_n261_bF_buf2), .B(\wb_addr_i[0] ), .Y(u1__abc_45852_n561) );
  AND2X2 AND2X2_3347 ( .A(csc_s_5_bF_buf0), .B(\wb_addr_i[2] ), .Y(u1__abc_45852_n563) );
  AND2X2 AND2X2_3348 ( .A(u1__abc_45852_n566), .B(u1__abc_45852_n559), .Y(u1_acs_addr_0__FF_INPUT) );
  AND2X2 AND2X2_3349 ( .A(u1__abc_45852_n569), .B(u1__abc_45852_n568), .Y(u1__abc_45852_n570_1) );
  AND2X2 AND2X2_335 ( .A(u0__abc_49347_n1577), .B(u0__abc_49347_n1180_1_bF_buf1), .Y(u0__abc_49347_n1578_1) );
  AND2X2 AND2X2_3350 ( .A(u1__abc_45852_n276_bF_buf4), .B(\wb_addr_i[2] ), .Y(u1__abc_45852_n572) );
  AND2X2 AND2X2_3351 ( .A(u1__abc_45852_n261_bF_buf1), .B(\wb_addr_i[1] ), .Y(u1__abc_45852_n573_1) );
  AND2X2 AND2X2_3352 ( .A(csc_s_5_bF_buf4), .B(\wb_addr_i[3] ), .Y(u1__abc_45852_n574) );
  AND2X2 AND2X2_3353 ( .A(u1__abc_45852_n577), .B(u1__abc_45852_n571), .Y(u1_acs_addr_1__FF_INPUT) );
  AND2X2 AND2X2_3354 ( .A(u1__abc_45852_n580), .B(u1__abc_45852_n579_1), .Y(u1__abc_45852_n581) );
  AND2X2 AND2X2_3355 ( .A(u1__abc_45852_n276_bF_buf3), .B(\wb_addr_i[3] ), .Y(u1__abc_45852_n583) );
  AND2X2 AND2X2_3356 ( .A(u1__abc_45852_n261_bF_buf0), .B(\wb_addr_i[2] ), .Y(u1__abc_45852_n584) );
  AND2X2 AND2X2_3357 ( .A(csc_s_5_bF_buf3), .B(\wb_addr_i[4] ), .Y(u1__abc_45852_n585_1) );
  AND2X2 AND2X2_3358 ( .A(u1__abc_45852_n588_1), .B(u1__abc_45852_n582_1), .Y(u1_acs_addr_2__FF_INPUT) );
  AND2X2 AND2X2_3359 ( .A(u1__abc_45852_n591), .B(u1__abc_45852_n590_1), .Y(u1__abc_45852_n592) );
  AND2X2 AND2X2_336 ( .A(spec_req_cs_3_bF_buf4), .B(u0_tms3_16_), .Y(u0__abc_49347_n1579_1) );
  AND2X2 AND2X2_3360 ( .A(u1__abc_45852_n276_bF_buf2), .B(\wb_addr_i[4] ), .Y(u1__abc_45852_n594) );
  AND2X2 AND2X2_3361 ( .A(u1__abc_45852_n261_bF_buf4), .B(\wb_addr_i[3] ), .Y(u1__abc_45852_n595_1) );
  AND2X2 AND2X2_3362 ( .A(csc_s_5_bF_buf2), .B(\wb_addr_i[5] ), .Y(u1__abc_45852_n596) );
  AND2X2 AND2X2_3363 ( .A(u1__abc_45852_n599_1), .B(u1__abc_45852_n593), .Y(u1_acs_addr_3__FF_INPUT) );
  AND2X2 AND2X2_3364 ( .A(u1__abc_45852_n602), .B(u1__abc_45852_n601_1), .Y(u1__abc_45852_n603) );
  AND2X2 AND2X2_3365 ( .A(u1__abc_45852_n276_bF_buf1), .B(\wb_addr_i[5] ), .Y(u1__abc_45852_n605) );
  AND2X2 AND2X2_3366 ( .A(u1__abc_45852_n261_bF_buf3), .B(\wb_addr_i[4] ), .Y(u1__abc_45852_n606) );
  AND2X2 AND2X2_3367 ( .A(csc_s_5_bF_buf1), .B(\wb_addr_i[6] ), .Y(u1__abc_45852_n607) );
  AND2X2 AND2X2_3368 ( .A(u1__abc_45852_n610), .B(u1__abc_45852_n604), .Y(u1_acs_addr_4__FF_INPUT) );
  AND2X2 AND2X2_3369 ( .A(u1__abc_45852_n613), .B(u1__abc_45852_n612), .Y(u1__abc_45852_n614) );
  AND2X2 AND2X2_337 ( .A(u0__abc_49347_n1580), .B(u0__abc_49347_n1179_bF_buf1), .Y(u0__abc_49347_n1581) );
  AND2X2 AND2X2_3370 ( .A(u1__abc_45852_n276_bF_buf0), .B(\wb_addr_i[6] ), .Y(u1__abc_45852_n616) );
  AND2X2 AND2X2_3371 ( .A(u1__abc_45852_n261_bF_buf2), .B(\wb_addr_i[5] ), .Y(u1__abc_45852_n617) );
  AND2X2 AND2X2_3372 ( .A(csc_s_5_bF_buf0), .B(\wb_addr_i[7] ), .Y(u1__abc_45852_n618) );
  AND2X2 AND2X2_3373 ( .A(u1__abc_45852_n621), .B(u1__abc_45852_n615), .Y(u1_acs_addr_5__FF_INPUT) );
  AND2X2 AND2X2_3374 ( .A(u1__abc_45852_n624), .B(u1__abc_45852_n623), .Y(u1__abc_45852_n625) );
  AND2X2 AND2X2_3375 ( .A(u1__abc_45852_n276_bF_buf4), .B(\wb_addr_i[7] ), .Y(u1__abc_45852_n627) );
  AND2X2 AND2X2_3376 ( .A(u1__abc_45852_n261_bF_buf1), .B(\wb_addr_i[6] ), .Y(u1__abc_45852_n628) );
  AND2X2 AND2X2_3377 ( .A(csc_s_5_bF_buf4), .B(\wb_addr_i[8] ), .Y(u1__abc_45852_n629) );
  AND2X2 AND2X2_3378 ( .A(u1__abc_45852_n632), .B(u1__abc_45852_n626), .Y(u1_acs_addr_6__FF_INPUT) );
  AND2X2 AND2X2_3379 ( .A(u1__abc_45852_n635), .B(u1__abc_45852_n634), .Y(u1__abc_45852_n636) );
  AND2X2 AND2X2_338 ( .A(spec_req_cs_2_bF_buf4), .B(u0_tms2_16_), .Y(u0__abc_49347_n1582) );
  AND2X2 AND2X2_3380 ( .A(u1__abc_45852_n276_bF_buf3), .B(\wb_addr_i[8] ), .Y(u1__abc_45852_n638) );
  AND2X2 AND2X2_3381 ( .A(u1__abc_45852_n261_bF_buf0), .B(\wb_addr_i[7] ), .Y(u1__abc_45852_n639) );
  AND2X2 AND2X2_3382 ( .A(csc_s_5_bF_buf3), .B(\wb_addr_i[9] ), .Y(u1__abc_45852_n640) );
  AND2X2 AND2X2_3383 ( .A(u1__abc_45852_n643), .B(u1__abc_45852_n637), .Y(u1_acs_addr_7__FF_INPUT) );
  AND2X2 AND2X2_3384 ( .A(u1__abc_45852_n646), .B(u1__abc_45852_n645), .Y(u1__abc_45852_n647) );
  AND2X2 AND2X2_3385 ( .A(u1__abc_45852_n276_bF_buf2), .B(\wb_addr_i[9] ), .Y(u1__abc_45852_n649) );
  AND2X2 AND2X2_3386 ( .A(u1__abc_45852_n261_bF_buf4), .B(\wb_addr_i[8] ), .Y(u1__abc_45852_n650) );
  AND2X2 AND2X2_3387 ( .A(csc_s_5_bF_buf2), .B(\wb_addr_i[10] ), .Y(u1__abc_45852_n651) );
  AND2X2 AND2X2_3388 ( .A(u1__abc_45852_n654), .B(u1__abc_45852_n648), .Y(u1_acs_addr_8__FF_INPUT) );
  AND2X2 AND2X2_3389 ( .A(u1__abc_45852_n657), .B(u1__abc_45852_n656), .Y(u1__abc_45852_n658) );
  AND2X2 AND2X2_339 ( .A(u0__abc_49347_n1583), .B(u0__abc_49347_n1178_1_bF_buf1), .Y(u0__abc_49347_n1584) );
  AND2X2 AND2X2_3390 ( .A(u1__abc_45852_n276_bF_buf1), .B(\wb_addr_i[10] ), .Y(u1__abc_45852_n660) );
  AND2X2 AND2X2_3391 ( .A(u1__abc_45852_n261_bF_buf3), .B(\wb_addr_i[9] ), .Y(u1__abc_45852_n661) );
  AND2X2 AND2X2_3392 ( .A(csc_s_5_bF_buf1), .B(\wb_addr_i[11] ), .Y(u1__abc_45852_n662) );
  AND2X2 AND2X2_3393 ( .A(u1__abc_45852_n665), .B(u1__abc_45852_n659), .Y(u1_acs_addr_9__FF_INPUT) );
  AND2X2 AND2X2_3394 ( .A(u1__abc_45852_n668), .B(u1__abc_45852_n667), .Y(u1__abc_45852_n669) );
  AND2X2 AND2X2_3395 ( .A(u1__abc_45852_n276_bF_buf0), .B(\wb_addr_i[11] ), .Y(u1__abc_45852_n671) );
  AND2X2 AND2X2_3396 ( .A(u1__abc_45852_n261_bF_buf2), .B(\wb_addr_i[10] ), .Y(u1__abc_45852_n672) );
  AND2X2 AND2X2_3397 ( .A(csc_s_5_bF_buf0), .B(\wb_addr_i[12] ), .Y(u1__abc_45852_n673) );
  AND2X2 AND2X2_3398 ( .A(u1__abc_45852_n676), .B(u1__abc_45852_n670), .Y(u1_acs_addr_10__FF_INPUT) );
  AND2X2 AND2X2_3399 ( .A(u1__abc_45852_n679), .B(u1__abc_45852_n678), .Y(u1__abc_45852_n680) );
  AND2X2 AND2X2_34 ( .A(_abc_55805_n338), .B(_abc_55805_n339), .Y(tms_s_16_) );
  AND2X2 AND2X2_340 ( .A(spec_req_cs_1_bF_buf4), .B(u0_tms1_16_), .Y(u0__abc_49347_n1585) );
  AND2X2 AND2X2_3400 ( .A(u1__abc_45852_n276_bF_buf4), .B(\wb_addr_i[12] ), .Y(u1__abc_45852_n682) );
  AND2X2 AND2X2_3401 ( .A(u1__abc_45852_n261_bF_buf1), .B(\wb_addr_i[11] ), .Y(u1__abc_45852_n683) );
  AND2X2 AND2X2_3402 ( .A(csc_s_5_bF_buf4), .B(\wb_addr_i[13] ), .Y(u1__abc_45852_n684) );
  AND2X2 AND2X2_3403 ( .A(u1__abc_45852_n687), .B(u1__abc_45852_n681), .Y(u1_acs_addr_11__FF_INPUT) );
  AND2X2 AND2X2_3404 ( .A(u1__abc_45852_n690), .B(u1__abc_45852_n689), .Y(u1__abc_45852_n691) );
  AND2X2 AND2X2_3405 ( .A(u1__abc_45852_n276_bF_buf3), .B(\wb_addr_i[13] ), .Y(u1__abc_45852_n693) );
  AND2X2 AND2X2_3406 ( .A(u1__abc_45852_n261_bF_buf0), .B(\wb_addr_i[12] ), .Y(u1__abc_45852_n694) );
  AND2X2 AND2X2_3407 ( .A(csc_s_5_bF_buf3), .B(\wb_addr_i[14] ), .Y(u1__abc_45852_n695) );
  AND2X2 AND2X2_3408 ( .A(u1__abc_45852_n698), .B(u1__abc_45852_n692), .Y(u1_acs_addr_12__FF_INPUT) );
  AND2X2 AND2X2_3409 ( .A(u1__abc_45852_n701), .B(u1__abc_45852_n700), .Y(u1__abc_45852_n702) );
  AND2X2 AND2X2_341 ( .A(u0__abc_49347_n1175_bF_buf3), .B(u0__abc_49347_n1588_1), .Y(u0__abc_49347_n1589) );
  AND2X2 AND2X2_3410 ( .A(u1__abc_45852_n276_bF_buf2), .B(\wb_addr_i[14] ), .Y(u1__abc_45852_n704) );
  AND2X2 AND2X2_3411 ( .A(u1__abc_45852_n261_bF_buf4), .B(\wb_addr_i[13] ), .Y(u1__abc_45852_n705) );
  AND2X2 AND2X2_3412 ( .A(csc_s_5_bF_buf2), .B(\wb_addr_i[15] ), .Y(u1__abc_45852_n706) );
  AND2X2 AND2X2_3413 ( .A(u1__abc_45852_n709), .B(u1__abc_45852_n703), .Y(u1_acs_addr_13__FF_INPUT) );
  AND2X2 AND2X2_3414 ( .A(u1__abc_45852_n712), .B(u1__abc_45852_n711), .Y(u1__abc_45852_n713) );
  AND2X2 AND2X2_3415 ( .A(u1__abc_45852_n276_bF_buf1), .B(\wb_addr_i[15] ), .Y(u1__abc_45852_n715) );
  AND2X2 AND2X2_3416 ( .A(u1__abc_45852_n261_bF_buf3), .B(\wb_addr_i[14] ), .Y(u1__abc_45852_n716) );
  AND2X2 AND2X2_3417 ( .A(csc_s_5_bF_buf1), .B(\wb_addr_i[16] ), .Y(u1__abc_45852_n717) );
  AND2X2 AND2X2_3418 ( .A(u1__abc_45852_n720), .B(u1__abc_45852_n714), .Y(u1_acs_addr_14__FF_INPUT) );
  AND2X2 AND2X2_3419 ( .A(u1__abc_45852_n723), .B(u1__abc_45852_n722), .Y(u1__abc_45852_n724) );
  AND2X2 AND2X2_342 ( .A(u0__abc_49347_n1587_1), .B(u0__abc_49347_n1589), .Y(u0__abc_49347_n1590) );
  AND2X2 AND2X2_3420 ( .A(u1__abc_45852_n276_bF_buf0), .B(\wb_addr_i[16] ), .Y(u1__abc_45852_n726) );
  AND2X2 AND2X2_3421 ( .A(u1__abc_45852_n261_bF_buf2), .B(\wb_addr_i[15] ), .Y(u1__abc_45852_n727) );
  AND2X2 AND2X2_3422 ( .A(csc_s_5_bF_buf0), .B(\wb_addr_i[17] ), .Y(u1__abc_45852_n728) );
  AND2X2 AND2X2_3423 ( .A(u1__abc_45852_n731), .B(u1__abc_45852_n725), .Y(u1_acs_addr_15__FF_INPUT) );
  AND2X2 AND2X2_3424 ( .A(u1__abc_45852_n734), .B(u1__abc_45852_n733), .Y(u1__abc_45852_n735) );
  AND2X2 AND2X2_3425 ( .A(u1__abc_45852_n276_bF_buf4), .B(\wb_addr_i[17] ), .Y(u1__abc_45852_n737) );
  AND2X2 AND2X2_3426 ( .A(u1__abc_45852_n261_bF_buf1), .B(\wb_addr_i[16] ), .Y(u1__abc_45852_n738) );
  AND2X2 AND2X2_3427 ( .A(csc_s_5_bF_buf4), .B(\wb_addr_i[18] ), .Y(u1__abc_45852_n739) );
  AND2X2 AND2X2_3428 ( .A(u1__abc_45852_n742), .B(u1__abc_45852_n736), .Y(u1_acs_addr_16__FF_INPUT) );
  AND2X2 AND2X2_3429 ( .A(u1__abc_45852_n745), .B(u1__abc_45852_n744), .Y(u1__abc_45852_n746) );
  AND2X2 AND2X2_343 ( .A(u0__abc_49347_n1176_1_bF_buf3), .B(sp_tms_17_), .Y(u0__abc_49347_n1592) );
  AND2X2 AND2X2_3430 ( .A(u1__abc_45852_n276_bF_buf3), .B(\wb_addr_i[18] ), .Y(u1__abc_45852_n748) );
  AND2X2 AND2X2_3431 ( .A(u1__abc_45852_n261_bF_buf0), .B(\wb_addr_i[17] ), .Y(u1__abc_45852_n749) );
  AND2X2 AND2X2_3432 ( .A(csc_s_5_bF_buf3), .B(\wb_addr_i[19] ), .Y(u1__abc_45852_n750) );
  AND2X2 AND2X2_3433 ( .A(u1__abc_45852_n753), .B(u1__abc_45852_n747), .Y(u1_acs_addr_17__FF_INPUT) );
  AND2X2 AND2X2_3434 ( .A(u1__abc_45852_n756), .B(u1__abc_45852_n755), .Y(u1__abc_45852_n757) );
  AND2X2 AND2X2_3435 ( .A(u1__abc_45852_n276_bF_buf2), .B(\wb_addr_i[19] ), .Y(u1__abc_45852_n759) );
  AND2X2 AND2X2_3436 ( .A(u1__abc_45852_n261_bF_buf4), .B(\wb_addr_i[18] ), .Y(u1__abc_45852_n760) );
  AND2X2 AND2X2_3437 ( .A(csc_s_5_bF_buf2), .B(\wb_addr_i[20] ), .Y(u1__abc_45852_n761) );
  AND2X2 AND2X2_3438 ( .A(u1__abc_45852_n764), .B(u1__abc_45852_n758), .Y(u1_acs_addr_18__FF_INPUT) );
  AND2X2 AND2X2_3439 ( .A(u1__abc_45852_n767), .B(u1__abc_45852_n766), .Y(u1__abc_45852_n768) );
  AND2X2 AND2X2_344 ( .A(spec_req_cs_5_bF_buf3), .B(u0_tms5_17_), .Y(u0__abc_49347_n1593) );
  AND2X2 AND2X2_3440 ( .A(u1__abc_45852_n276_bF_buf1), .B(\wb_addr_i[20] ), .Y(u1__abc_45852_n770) );
  AND2X2 AND2X2_3441 ( .A(u1__abc_45852_n261_bF_buf3), .B(\wb_addr_i[19] ), .Y(u1__abc_45852_n771) );
  AND2X2 AND2X2_3442 ( .A(csc_s_5_bF_buf1), .B(\wb_addr_i[21] ), .Y(u1__abc_45852_n772) );
  AND2X2 AND2X2_3443 ( .A(u1__abc_45852_n775), .B(u1__abc_45852_n769), .Y(u1_acs_addr_19__FF_INPUT) );
  AND2X2 AND2X2_3444 ( .A(u1__abc_45852_n778), .B(u1__abc_45852_n777), .Y(u1__abc_45852_n779) );
  AND2X2 AND2X2_3445 ( .A(u1__abc_45852_n276_bF_buf0), .B(\wb_addr_i[21] ), .Y(u1__abc_45852_n781) );
  AND2X2 AND2X2_3446 ( .A(u1__abc_45852_n261_bF_buf2), .B(\wb_addr_i[20] ), .Y(u1__abc_45852_n782) );
  AND2X2 AND2X2_3447 ( .A(csc_s_5_bF_buf0), .B(\wb_addr_i[22] ), .Y(u1__abc_45852_n783) );
  AND2X2 AND2X2_3448 ( .A(u1__abc_45852_n786), .B(u1__abc_45852_n780), .Y(u1_acs_addr_20__FF_INPUT) );
  AND2X2 AND2X2_3449 ( .A(u1__abc_45852_n789), .B(u1__abc_45852_n788), .Y(u1__abc_45852_n790) );
  AND2X2 AND2X2_345 ( .A(u0__abc_49347_n1595), .B(u0__abc_49347_n1185_bF_buf0), .Y(u0__abc_49347_n1596_1) );
  AND2X2 AND2X2_3450 ( .A(u1__abc_45852_n276_bF_buf4), .B(\wb_addr_i[22] ), .Y(u1__abc_45852_n792) );
  AND2X2 AND2X2_3451 ( .A(u1__abc_45852_n261_bF_buf1), .B(\wb_addr_i[21] ), .Y(u1__abc_45852_n793) );
  AND2X2 AND2X2_3452 ( .A(csc_s_5_bF_buf4), .B(wb_addr_i_23_bF_buf1), .Y(u1__abc_45852_n794) );
  AND2X2 AND2X2_3453 ( .A(u1__abc_45852_n797), .B(u1__abc_45852_n791), .Y(u1_acs_addr_21__FF_INPUT) );
  AND2X2 AND2X2_3454 ( .A(u1__abc_45852_n800), .B(u1__abc_45852_n799), .Y(u1__abc_45852_n801) );
  AND2X2 AND2X2_3455 ( .A(u1__abc_45852_n261_bF_buf0), .B(\wb_addr_i[22] ), .Y(u1__abc_45852_n803) );
  AND2X2 AND2X2_3456 ( .A(csc_s_5_bF_buf3), .B(\wb_addr_i[24] ), .Y(u1__abc_45852_n804) );
  AND2X2 AND2X2_3457 ( .A(u1__abc_45852_n807), .B(u1__abc_45852_n802), .Y(u1_acs_addr_22__FF_INPUT) );
  AND2X2 AND2X2_3458 ( .A(u1__abc_45852_n810), .B(u1__abc_45852_n809), .Y(u1__abc_45852_n811) );
  AND2X2 AND2X2_3459 ( .A(u1__abc_45852_n276_bF_buf3), .B(\wb_addr_i[24] ), .Y(u1__abc_45852_n813) );
  AND2X2 AND2X2_346 ( .A(u0__abc_49347_n1596_1), .B(u0__abc_49347_n1594), .Y(u0__abc_49347_n1597_1) );
  AND2X2 AND2X2_3460 ( .A(u1__abc_45852_n261_bF_buf4), .B(wb_addr_i_23_bF_buf0), .Y(u1__abc_45852_n814) );
  AND2X2 AND2X2_3461 ( .A(csc_s_5_bF_buf2), .B(wb_addr_i_25_bF_buf3), .Y(u1__abc_45852_n815) );
  AND2X2 AND2X2_3462 ( .A(u1__abc_45852_n818), .B(u1__abc_45852_n812), .Y(u1_acs_addr_23__FF_INPUT) );
  AND2X2 AND2X2_3463 ( .A(u1__abc_45852_n822), .B(u1__abc_45852_n820), .Y(u1_sram_addr_0__FF_INPUT) );
  AND2X2 AND2X2_3464 ( .A(u1__abc_45852_n825), .B(u1__abc_45852_n824), .Y(u1_sram_addr_1__FF_INPUT) );
  AND2X2 AND2X2_3465 ( .A(u1__abc_45852_n828), .B(u1__abc_45852_n827), .Y(u1_sram_addr_2__FF_INPUT) );
  AND2X2 AND2X2_3466 ( .A(u1__abc_45852_n831), .B(u1__abc_45852_n830), .Y(u1_sram_addr_3__FF_INPUT) );
  AND2X2 AND2X2_3467 ( .A(u1__abc_45852_n834), .B(u1__abc_45852_n833), .Y(u1_sram_addr_4__FF_INPUT) );
  AND2X2 AND2X2_3468 ( .A(u1__abc_45852_n837), .B(u1__abc_45852_n836), .Y(u1_sram_addr_5__FF_INPUT) );
  AND2X2 AND2X2_3469 ( .A(u1__abc_45852_n840), .B(u1__abc_45852_n839), .Y(u1_sram_addr_6__FF_INPUT) );
  AND2X2 AND2X2_347 ( .A(u0__abc_49347_n1598), .B(u0__abc_49347_n1181_bF_buf0), .Y(u0__abc_49347_n1599) );
  AND2X2 AND2X2_3470 ( .A(u1__abc_45852_n843), .B(u1__abc_45852_n842), .Y(u1_sram_addr_7__FF_INPUT) );
  AND2X2 AND2X2_3471 ( .A(u1__abc_45852_n846), .B(u1__abc_45852_n845), .Y(u1_sram_addr_8__FF_INPUT) );
  AND2X2 AND2X2_3472 ( .A(u1__abc_45852_n849), .B(u1__abc_45852_n848), .Y(u1_sram_addr_9__FF_INPUT) );
  AND2X2 AND2X2_3473 ( .A(u1__abc_45852_n852), .B(u1__abc_45852_n851), .Y(u1_sram_addr_10__FF_INPUT) );
  AND2X2 AND2X2_3474 ( .A(u1__abc_45852_n855), .B(u1__abc_45852_n854), .Y(u1_sram_addr_11__FF_INPUT) );
  AND2X2 AND2X2_3475 ( .A(u1__abc_45852_n858), .B(u1__abc_45852_n857), .Y(u1_sram_addr_12__FF_INPUT) );
  AND2X2 AND2X2_3476 ( .A(u1__abc_45852_n861), .B(u1__abc_45852_n860), .Y(u1_sram_addr_13__FF_INPUT) );
  AND2X2 AND2X2_3477 ( .A(u1__abc_45852_n864), .B(u1__abc_45852_n863), .Y(u1_sram_addr_14__FF_INPUT) );
  AND2X2 AND2X2_3478 ( .A(u1__abc_45852_n867), .B(u1__abc_45852_n866), .Y(u1_sram_addr_15__FF_INPUT) );
  AND2X2 AND2X2_3479 ( .A(u1__abc_45852_n870), .B(u1__abc_45852_n869), .Y(u1_sram_addr_16__FF_INPUT) );
  AND2X2 AND2X2_348 ( .A(spec_req_cs_4_bF_buf3), .B(u0_tms4_17_), .Y(u0__abc_49347_n1600) );
  AND2X2 AND2X2_3480 ( .A(u1__abc_45852_n873), .B(u1__abc_45852_n872), .Y(u1_sram_addr_17__FF_INPUT) );
  AND2X2 AND2X2_3481 ( .A(u1__abc_45852_n876), .B(u1__abc_45852_n875), .Y(u1_sram_addr_18__FF_INPUT) );
  AND2X2 AND2X2_3482 ( .A(u1__abc_45852_n879), .B(u1__abc_45852_n878), .Y(u1_sram_addr_19__FF_INPUT) );
  AND2X2 AND2X2_3483 ( .A(u1__abc_45852_n882), .B(u1__abc_45852_n881), .Y(u1_sram_addr_20__FF_INPUT) );
  AND2X2 AND2X2_3484 ( .A(u1__abc_45852_n885), .B(u1__abc_45852_n884), .Y(u1_sram_addr_21__FF_INPUT) );
  AND2X2 AND2X2_3485 ( .A(u1__abc_45852_n888), .B(u1__abc_45852_n887), .Y(u1_sram_addr_22__FF_INPUT) );
  AND2X2 AND2X2_3486 ( .A(u1__abc_45852_n891), .B(u1__abc_45852_n890), .Y(u1_sram_addr_23__FF_INPUT) );
  AND2X2 AND2X2_3487 ( .A(u1_acs_addr_0_), .B(csc_s_2_bF_buf4), .Y(u1__abc_45852_n894) );
  AND2X2 AND2X2_3488 ( .A(u1__abc_45852_n896), .B(csc_s_2_bF_buf3), .Y(u1__abc_45852_n897) );
  AND2X2 AND2X2_3489 ( .A(csc_s_1_), .B(u1_wr_hold), .Y(u1__abc_45852_n900) );
  AND2X2 AND2X2_349 ( .A(u0__abc_49347_n1601), .B(u0__abc_49347_n1180_1_bF_buf0), .Y(u0__abc_49347_n1602) );
  AND2X2 AND2X2_3490 ( .A(u1__abc_45852_n899), .B(u1__abc_45852_n900), .Y(u1__abc_45852_n901) );
  AND2X2 AND2X2_3491 ( .A(u1__abc_45852_n901_bF_buf4), .B(u1_sram_addr_0_), .Y(u1__abc_45852_n902) );
  AND2X2 AND2X2_3492 ( .A(u1__abc_45852_n903_bF_buf3), .B(\wb_addr_i[2] ), .Y(u1__abc_45852_n904) );
  AND2X2 AND2X2_3493 ( .A(u1__abc_45852_n906), .B(u1__abc_45852_n895), .Y(u1__abc_45852_n907) );
  AND2X2 AND2X2_3494 ( .A(u1__abc_45852_n908), .B(lmr_sel_bF_buf3), .Y(u1__abc_45852_n909) );
  AND2X2 AND2X2_3495 ( .A(u1__abc_45852_n911), .B(u1__abc_45852_n912), .Y(u1__abc_45852_n913) );
  AND2X2 AND2X2_3496 ( .A(u1__abc_45852_n896), .B(u1__abc_45852_n915), .Y(u1__abc_45852_n916) );
  AND2X2 AND2X2_3497 ( .A(u1__abc_45852_n918), .B(u1__abc_45852_n916), .Y(u1__abc_45852_n919) );
  AND2X2 AND2X2_3498 ( .A(u1__abc_45852_n919), .B(u1__abc_45852_n914), .Y(u1__abc_45852_n920) );
  AND2X2 AND2X2_3499 ( .A(u1_acs_addr_1_), .B(csc_s_2_bF_buf0), .Y(u1__abc_45852_n922) );
  AND2X2 AND2X2_35 ( .A(_abc_55805_n341), .B(_abc_55805_n342), .Y(tms_s_17_) );
  AND2X2 AND2X2_350 ( .A(spec_req_cs_3_bF_buf3), .B(u0_tms3_17_), .Y(u0__abc_49347_n1603) );
  AND2X2 AND2X2_3500 ( .A(u1__abc_45852_n901_bF_buf2), .B(u1_sram_addr_1_), .Y(u1__abc_45852_n924) );
  AND2X2 AND2X2_3501 ( .A(u1__abc_45852_n903_bF_buf2), .B(\wb_addr_i[3] ), .Y(u1__abc_45852_n925) );
  AND2X2 AND2X2_3502 ( .A(u1__abc_45852_n927), .B(u1__abc_45852_n923), .Y(u1__abc_45852_n928) );
  AND2X2 AND2X2_3503 ( .A(u1__abc_45852_n929), .B(u1__abc_45852_n930), .Y(u1__abc_45852_n931) );
  AND2X2 AND2X2_3504 ( .A(u1__abc_45852_n933), .B(u1__abc_45852_n916), .Y(u1__abc_45852_n934) );
  AND2X2 AND2X2_3505 ( .A(u1__abc_45852_n934), .B(u1__abc_45852_n932), .Y(u1__abc_45852_n935) );
  AND2X2 AND2X2_3506 ( .A(u1_acs_addr_2_), .B(csc_s_2_bF_buf4), .Y(u1__abc_45852_n937) );
  AND2X2 AND2X2_3507 ( .A(u1__abc_45852_n901_bF_buf1), .B(u1_sram_addr_2_), .Y(u1__abc_45852_n939) );
  AND2X2 AND2X2_3508 ( .A(u1__abc_45852_n903_bF_buf1), .B(\wb_addr_i[4] ), .Y(u1__abc_45852_n940) );
  AND2X2 AND2X2_3509 ( .A(u1__abc_45852_n942), .B(u1__abc_45852_n938), .Y(u1__abc_45852_n943) );
  AND2X2 AND2X2_351 ( .A(u0__abc_49347_n1604), .B(u0__abc_49347_n1179_bF_buf0), .Y(u0__abc_49347_n1605_1) );
  AND2X2 AND2X2_3510 ( .A(u1__abc_45852_n944), .B(u1__abc_45852_n945), .Y(u1__abc_45852_n946) );
  AND2X2 AND2X2_3511 ( .A(u1__abc_45852_n948), .B(u1__abc_45852_n916), .Y(u1__abc_45852_n949) );
  AND2X2 AND2X2_3512 ( .A(u1__abc_45852_n949), .B(u1__abc_45852_n947), .Y(u1__abc_45852_n950) );
  AND2X2 AND2X2_3513 ( .A(u1_acs_addr_3_), .B(csc_s_2_bF_buf3), .Y(u1__abc_45852_n952) );
  AND2X2 AND2X2_3514 ( .A(u1__abc_45852_n901_bF_buf0), .B(u1_sram_addr_3_), .Y(u1__abc_45852_n954) );
  AND2X2 AND2X2_3515 ( .A(u1__abc_45852_n903_bF_buf0), .B(\wb_addr_i[5] ), .Y(u1__abc_45852_n955) );
  AND2X2 AND2X2_3516 ( .A(u1__abc_45852_n957), .B(u1__abc_45852_n953), .Y(u1__abc_45852_n958) );
  AND2X2 AND2X2_3517 ( .A(u1__abc_45852_n959), .B(u1__abc_45852_n960), .Y(u1__abc_45852_n961) );
  AND2X2 AND2X2_3518 ( .A(u1__abc_45852_n963), .B(u1__abc_45852_n916), .Y(u1__abc_45852_n964) );
  AND2X2 AND2X2_3519 ( .A(u1__abc_45852_n964), .B(u1__abc_45852_n962), .Y(u1__abc_45852_n965) );
  AND2X2 AND2X2_352 ( .A(spec_req_cs_2_bF_buf3), .B(u0_tms2_17_), .Y(u0__abc_49347_n1606_1) );
  AND2X2 AND2X2_3520 ( .A(u1_acs_addr_4_), .B(csc_s_2_bF_buf2), .Y(u1__abc_45852_n967) );
  AND2X2 AND2X2_3521 ( .A(u1__abc_45852_n901_bF_buf4), .B(u1_sram_addr_4_), .Y(u1__abc_45852_n969) );
  AND2X2 AND2X2_3522 ( .A(u1__abc_45852_n903_bF_buf3), .B(\wb_addr_i[6] ), .Y(u1__abc_45852_n970) );
  AND2X2 AND2X2_3523 ( .A(u1__abc_45852_n972), .B(u1__abc_45852_n968), .Y(u1__abc_45852_n973) );
  AND2X2 AND2X2_3524 ( .A(u1__abc_45852_n974), .B(u1__abc_45852_n975), .Y(u1__abc_45852_n976) );
  AND2X2 AND2X2_3525 ( .A(u1__abc_45852_n978), .B(u1__abc_45852_n916), .Y(u1__abc_45852_n979) );
  AND2X2 AND2X2_3526 ( .A(u1__abc_45852_n979), .B(u1__abc_45852_n977), .Y(u1__abc_45852_n980) );
  AND2X2 AND2X2_3527 ( .A(u1_acs_addr_5_), .B(csc_s_2_bF_buf1), .Y(u1__abc_45852_n982) );
  AND2X2 AND2X2_3528 ( .A(u1__abc_45852_n901_bF_buf3), .B(u1_sram_addr_5_), .Y(u1__abc_45852_n984) );
  AND2X2 AND2X2_3529 ( .A(u1__abc_45852_n903_bF_buf2), .B(\wb_addr_i[7] ), .Y(u1__abc_45852_n985) );
  AND2X2 AND2X2_353 ( .A(u0__abc_49347_n1607), .B(u0__abc_49347_n1178_1_bF_buf0), .Y(u0__abc_49347_n1608) );
  AND2X2 AND2X2_3530 ( .A(u1__abc_45852_n987), .B(u1__abc_45852_n983), .Y(u1__abc_45852_n988) );
  AND2X2 AND2X2_3531 ( .A(u1__abc_45852_n989), .B(u1__abc_45852_n990), .Y(u1__abc_45852_n991) );
  AND2X2 AND2X2_3532 ( .A(u1__abc_45852_n993), .B(u1__abc_45852_n916), .Y(u1__abc_45852_n994) );
  AND2X2 AND2X2_3533 ( .A(u1__abc_45852_n994), .B(u1__abc_45852_n992), .Y(u1__abc_45852_n995) );
  AND2X2 AND2X2_3534 ( .A(u1_acs_addr_6_), .B(csc_s_2_bF_buf0), .Y(u1__abc_45852_n997) );
  AND2X2 AND2X2_3535 ( .A(u1__abc_45852_n901_bF_buf2), .B(u1_sram_addr_6_), .Y(u1__abc_45852_n999) );
  AND2X2 AND2X2_3536 ( .A(u1__abc_45852_n903_bF_buf1), .B(\wb_addr_i[8] ), .Y(u1__abc_45852_n1000) );
  AND2X2 AND2X2_3537 ( .A(u1__abc_45852_n1002), .B(u1__abc_45852_n998), .Y(u1__abc_45852_n1003) );
  AND2X2 AND2X2_3538 ( .A(u1__abc_45852_n1004), .B(u1__abc_45852_n1005), .Y(u1__abc_45852_n1006) );
  AND2X2 AND2X2_3539 ( .A(u1__abc_45852_n1008), .B(u1__abc_45852_n916), .Y(u1__abc_45852_n1009) );
  AND2X2 AND2X2_354 ( .A(spec_req_cs_1_bF_buf3), .B(u0_tms1_17_), .Y(u0__abc_49347_n1609) );
  AND2X2 AND2X2_3540 ( .A(u1__abc_45852_n1009), .B(u1__abc_45852_n1007), .Y(u1__abc_45852_n1010) );
  AND2X2 AND2X2_3541 ( .A(u1_acs_addr_7_), .B(csc_s_2_bF_buf4), .Y(u1__abc_45852_n1012) );
  AND2X2 AND2X2_3542 ( .A(u1__abc_45852_n901_bF_buf1), .B(u1_sram_addr_7_), .Y(u1__abc_45852_n1014) );
  AND2X2 AND2X2_3543 ( .A(u1__abc_45852_n903_bF_buf0), .B(\wb_addr_i[9] ), .Y(u1__abc_45852_n1015) );
  AND2X2 AND2X2_3544 ( .A(u1__abc_45852_n1017), .B(u1__abc_45852_n1013), .Y(u1__abc_45852_n1018) );
  AND2X2 AND2X2_3545 ( .A(u1__abc_45852_n1019), .B(u1__abc_45852_n1020), .Y(u1__abc_45852_n1021) );
  AND2X2 AND2X2_3546 ( .A(u1__abc_45852_n1023), .B(u1__abc_45852_n916), .Y(u1__abc_45852_n1024) );
  AND2X2 AND2X2_3547 ( .A(u1__abc_45852_n1024), .B(u1__abc_45852_n1022), .Y(u1__abc_45852_n1025) );
  AND2X2 AND2X2_3548 ( .A(u1_acs_addr_8_), .B(csc_s_2_bF_buf3), .Y(u1__abc_45852_n1027) );
  AND2X2 AND2X2_3549 ( .A(u1__abc_45852_n901_bF_buf0), .B(u1_sram_addr_8_), .Y(u1__abc_45852_n1029) );
  AND2X2 AND2X2_355 ( .A(u0__abc_49347_n1175_bF_buf2), .B(u0__abc_49347_n1612), .Y(u0__abc_49347_n1613) );
  AND2X2 AND2X2_3550 ( .A(u1__abc_45852_n903_bF_buf3), .B(\wb_addr_i[10] ), .Y(u1__abc_45852_n1030) );
  AND2X2 AND2X2_3551 ( .A(u1__abc_45852_n1032), .B(u1__abc_45852_n1028), .Y(u1__abc_45852_n1033) );
  AND2X2 AND2X2_3552 ( .A(u1__abc_45852_n1034), .B(u1__abc_45852_n1035), .Y(u1__abc_45852_n1036) );
  AND2X2 AND2X2_3553 ( .A(u1__abc_45852_n1038), .B(u1__abc_45852_n916), .Y(u1__abc_45852_n1039) );
  AND2X2 AND2X2_3554 ( .A(u1__abc_45852_n1039), .B(u1__abc_45852_n1037), .Y(u1__abc_45852_n1040) );
  AND2X2 AND2X2_3555 ( .A(u1_acs_addr_9_), .B(csc_s_2_bF_buf2), .Y(u1__abc_45852_n1042) );
  AND2X2 AND2X2_3556 ( .A(u1__abc_45852_n901_bF_buf4), .B(u1_sram_addr_9_), .Y(u1__abc_45852_n1044) );
  AND2X2 AND2X2_3557 ( .A(u1__abc_45852_n903_bF_buf2), .B(\wb_addr_i[11] ), .Y(u1__abc_45852_n1045) );
  AND2X2 AND2X2_3558 ( .A(u1__abc_45852_n1047), .B(u1__abc_45852_n1043), .Y(u1__abc_45852_n1048) );
  AND2X2 AND2X2_3559 ( .A(u1__abc_45852_n1049), .B(u1__abc_45852_n1050), .Y(u1__abc_45852_n1051) );
  AND2X2 AND2X2_356 ( .A(u0__abc_49347_n1611), .B(u0__abc_49347_n1613), .Y(u0__abc_49347_n1614_1) );
  AND2X2 AND2X2_3560 ( .A(u1__abc_45852_n1053), .B(u1__abc_45852_n916), .Y(u1__abc_45852_n1054) );
  AND2X2 AND2X2_3561 ( .A(u1__abc_45852_n1054), .B(u1__abc_45852_n1052), .Y(u1__abc_45852_n1055) );
  AND2X2 AND2X2_3562 ( .A(row_adr_11_bF_buf5), .B(row_sel), .Y(u1__abc_45852_n1058) );
  AND2X2 AND2X2_3563 ( .A(u1__abc_45852_n916), .B(u1__abc_45852_n1059), .Y(u1__abc_45852_n1060) );
  AND2X2 AND2X2_3564 ( .A(u1__abc_45852_n1060), .B(u1__abc_45852_n1057), .Y(u1__abc_45852_n1061) );
  AND2X2 AND2X2_3565 ( .A(u1_acs_addr_11_), .B(csc_s_2_bF_buf1), .Y(u1__abc_45852_n1062) );
  AND2X2 AND2X2_3566 ( .A(u1__abc_45852_n1064), .B(u1__abc_45852_n1065), .Y(u1__abc_45852_n1066) );
  AND2X2 AND2X2_3567 ( .A(u1__abc_45852_n1067), .B(u1__abc_45852_n1063), .Y(u1__abc_45852_n1068) );
  AND2X2 AND2X2_3568 ( .A(row_adr_12_bF_buf5), .B(row_sel), .Y(u1__abc_45852_n1071) );
  AND2X2 AND2X2_3569 ( .A(u1__abc_45852_n916), .B(u1__abc_45852_n1072), .Y(u1__abc_45852_n1073) );
  AND2X2 AND2X2_357 ( .A(u0__abc_49347_n1176_1_bF_buf2), .B(sp_tms_18_), .Y(u0__abc_49347_n1616) );
  AND2X2 AND2X2_3570 ( .A(u1__abc_45852_n1073), .B(u1__abc_45852_n1070), .Y(u1__abc_45852_n1074) );
  AND2X2 AND2X2_3571 ( .A(u1_acs_addr_12_), .B(csc_s_2_bF_buf0), .Y(u1__abc_45852_n1075) );
  AND2X2 AND2X2_3572 ( .A(u1__abc_45852_n1077), .B(u1__abc_45852_n1078), .Y(u1__abc_45852_n1079) );
  AND2X2 AND2X2_3573 ( .A(u1__abc_45852_n1080), .B(u1__abc_45852_n1076), .Y(u1__abc_45852_n1081) );
  AND2X2 AND2X2_3574 ( .A(u1__abc_45852_n916), .B(bank_adr_0_bF_buf2), .Y(u1__abc_45852_n1083) );
  AND2X2 AND2X2_3575 ( .A(u1_acs_addr_13_), .B(csc_s_2_bF_buf4), .Y(u1__abc_45852_n1084) );
  AND2X2 AND2X2_3576 ( .A(u1__abc_45852_n1086), .B(u1__abc_45852_n1087), .Y(u1__abc_45852_n1088) );
  AND2X2 AND2X2_3577 ( .A(u1__abc_45852_n1089), .B(u1__abc_45852_n1085), .Y(u1__abc_45852_n1090) );
  AND2X2 AND2X2_3578 ( .A(u1__abc_45852_n916), .B(bank_adr_1_bF_buf2), .Y(u1__abc_45852_n1092) );
  AND2X2 AND2X2_3579 ( .A(u1_acs_addr_14_), .B(csc_s_2_bF_buf3), .Y(u1__abc_45852_n1093) );
  AND2X2 AND2X2_358 ( .A(spec_req_cs_5_bF_buf2), .B(u0_tms5_18_), .Y(u0__abc_49347_n1617) );
  AND2X2 AND2X2_3580 ( .A(u1__abc_45852_n1095), .B(u1__abc_45852_n1096), .Y(u1__abc_45852_n1097) );
  AND2X2 AND2X2_3581 ( .A(u1__abc_45852_n1098), .B(u1__abc_45852_n1094), .Y(u1__abc_45852_n1099) );
  AND2X2 AND2X2_3582 ( .A(u1_acs_addr_15_), .B(csc_s_2_bF_buf2), .Y(u1__abc_45852_n1101) );
  AND2X2 AND2X2_3583 ( .A(u1__abc_45852_n903_bF_buf1), .B(\wb_addr_i[17] ), .Y(u1__abc_45852_n1103) );
  AND2X2 AND2X2_3584 ( .A(u1__abc_45852_n901_bF_buf4), .B(u1_sram_addr_15_), .Y(u1__abc_45852_n1104) );
  AND2X2 AND2X2_3585 ( .A(u1__abc_45852_n1106), .B(u1__abc_45852_n1102), .Y(mc_addr_d_15_) );
  AND2X2 AND2X2_3586 ( .A(u1_acs_addr_16_), .B(csc_s_2_bF_buf1), .Y(u1__abc_45852_n1108) );
  AND2X2 AND2X2_3587 ( .A(u1__abc_45852_n901_bF_buf3), .B(u1_sram_addr_16_), .Y(u1__abc_45852_n1110) );
  AND2X2 AND2X2_3588 ( .A(u1__abc_45852_n903_bF_buf0), .B(\wb_addr_i[18] ), .Y(u1__abc_45852_n1111) );
  AND2X2 AND2X2_3589 ( .A(u1__abc_45852_n1113), .B(u1__abc_45852_n1109), .Y(mc_addr_d_16_) );
  AND2X2 AND2X2_359 ( .A(u0__abc_49347_n1619), .B(u0__abc_49347_n1185_bF_buf5), .Y(u0__abc_49347_n1620) );
  AND2X2 AND2X2_3590 ( .A(u1_acs_addr_17_), .B(csc_s_2_bF_buf0), .Y(u1__abc_45852_n1115) );
  AND2X2 AND2X2_3591 ( .A(u1__abc_45852_n901_bF_buf2), .B(u1_sram_addr_17_), .Y(u1__abc_45852_n1117) );
  AND2X2 AND2X2_3592 ( .A(u1__abc_45852_n903_bF_buf3), .B(\wb_addr_i[19] ), .Y(u1__abc_45852_n1118) );
  AND2X2 AND2X2_3593 ( .A(u1__abc_45852_n1120), .B(u1__abc_45852_n1116), .Y(mc_addr_d_17_) );
  AND2X2 AND2X2_3594 ( .A(u1_acs_addr_18_), .B(csc_s_2_bF_buf4), .Y(u1__abc_45852_n1122) );
  AND2X2 AND2X2_3595 ( .A(u1__abc_45852_n901_bF_buf1), .B(u1_sram_addr_18_), .Y(u1__abc_45852_n1124) );
  AND2X2 AND2X2_3596 ( .A(u1__abc_45852_n903_bF_buf2), .B(\wb_addr_i[20] ), .Y(u1__abc_45852_n1125) );
  AND2X2 AND2X2_3597 ( .A(u1__abc_45852_n1127), .B(u1__abc_45852_n1123), .Y(mc_addr_d_18_) );
  AND2X2 AND2X2_3598 ( .A(u1_acs_addr_19_), .B(csc_s_2_bF_buf3), .Y(u1__abc_45852_n1129) );
  AND2X2 AND2X2_3599 ( .A(u1__abc_45852_n901_bF_buf0), .B(u1_sram_addr_19_), .Y(u1__abc_45852_n1131) );
  AND2X2 AND2X2_36 ( .A(_abc_55805_n344), .B(_abc_55805_n345), .Y(tms_s_18_) );
  AND2X2 AND2X2_360 ( .A(u0__abc_49347_n1620), .B(u0__abc_49347_n1618), .Y(u0__abc_49347_n1621) );
  AND2X2 AND2X2_3600 ( .A(u1__abc_45852_n903_bF_buf1), .B(\wb_addr_i[21] ), .Y(u1__abc_45852_n1132) );
  AND2X2 AND2X2_3601 ( .A(u1__abc_45852_n1134), .B(u1__abc_45852_n1130), .Y(mc_addr_d_19_) );
  AND2X2 AND2X2_3602 ( .A(u1_acs_addr_20_), .B(csc_s_2_bF_buf2), .Y(u1__abc_45852_n1136) );
  AND2X2 AND2X2_3603 ( .A(u1__abc_45852_n901_bF_buf4), .B(u1_sram_addr_20_), .Y(u1__abc_45852_n1138) );
  AND2X2 AND2X2_3604 ( .A(u1__abc_45852_n903_bF_buf0), .B(\wb_addr_i[22] ), .Y(u1__abc_45852_n1139) );
  AND2X2 AND2X2_3605 ( .A(u1__abc_45852_n1141), .B(u1__abc_45852_n1137), .Y(mc_addr_d_20_) );
  AND2X2 AND2X2_3606 ( .A(u1_acs_addr_21_), .B(csc_s_2_bF_buf1), .Y(u1__abc_45852_n1143) );
  AND2X2 AND2X2_3607 ( .A(u1__abc_45852_n901_bF_buf3), .B(u1_sram_addr_21_), .Y(u1__abc_45852_n1145) );
  AND2X2 AND2X2_3608 ( .A(u1__abc_45852_n903_bF_buf3), .B(wb_addr_i_23_bF_buf2), .Y(u1__abc_45852_n1146) );
  AND2X2 AND2X2_3609 ( .A(u1__abc_45852_n1148), .B(u1__abc_45852_n1144), .Y(mc_addr_d_21_) );
  AND2X2 AND2X2_361 ( .A(u0__abc_49347_n1622), .B(u0__abc_49347_n1181_bF_buf5), .Y(u0__abc_49347_n1623_1) );
  AND2X2 AND2X2_3610 ( .A(u1_acs_addr_22_), .B(csc_s_2_bF_buf0), .Y(u1__abc_45852_n1150) );
  AND2X2 AND2X2_3611 ( .A(u1__abc_45852_n901_bF_buf2), .B(u1_sram_addr_22_), .Y(u1__abc_45852_n1152) );
  AND2X2 AND2X2_3612 ( .A(u1__abc_45852_n903_bF_buf2), .B(\wb_addr_i[24] ), .Y(u1__abc_45852_n1153) );
  AND2X2 AND2X2_3613 ( .A(u1__abc_45852_n1155), .B(u1__abc_45852_n1151), .Y(mc_addr_d_22_) );
  AND2X2 AND2X2_3614 ( .A(u1_acs_addr_23_), .B(csc_s_2_bF_buf4), .Y(u1__abc_45852_n1157) );
  AND2X2 AND2X2_3615 ( .A(u1__abc_45852_n901_bF_buf1), .B(u1_sram_addr_23_), .Y(u1__abc_45852_n1159) );
  AND2X2 AND2X2_3616 ( .A(u1__abc_45852_n903_bF_buf1), .B(wb_addr_i_25_bF_buf1), .Y(u1__abc_45852_n1160) );
  AND2X2 AND2X2_3617 ( .A(u1__abc_45852_n1162), .B(u1__abc_45852_n1158), .Y(mc_addr_d_23_) );
  AND2X2 AND2X2_3618 ( .A(u1__abc_45852_n1165), .B(u1__abc_45852_n1164), .Y(u1__abc_45852_n1166) );
  AND2X2 AND2X2_3619 ( .A(u1_acs_addr_10_), .B(csc_s_2_bF_buf3), .Y(u1__abc_45852_n1168) );
  AND2X2 AND2X2_362 ( .A(spec_req_cs_4_bF_buf2), .B(u0_tms4_18_), .Y(u0__abc_49347_n1624_1) );
  AND2X2 AND2X2_3620 ( .A(u1__abc_45852_n1167), .B(u1__abc_45852_n1169), .Y(u1__abc_45852_n1170) );
  AND2X2 AND2X2_3621 ( .A(u1__abc_45852_n1172), .B(u1__abc_45852_n1171), .Y(u1__abc_45852_n1173) );
  AND2X2 AND2X2_3622 ( .A(u1__abc_45852_n1175), .B(u1__abc_45852_n916), .Y(u1__abc_45852_n1176) );
  AND2X2 AND2X2_3623 ( .A(u1__abc_45852_n1176), .B(u1__abc_45852_n1174), .Y(u1__abc_45852_n1177) );
  AND2X2 AND2X2_3624 ( .A(u1_u0_inc_next), .B(u1_acs_addr_12_), .Y(u1_u0__abc_45749_n51) );
  AND2X2 AND2X2_3625 ( .A(u1_u0__abc_45749_n51), .B(u1_acs_addr_13_), .Y(u1_u0__abc_45749_n52_1) );
  AND2X2 AND2X2_3626 ( .A(u1_u0__abc_45749_n53_1), .B(u1_u0__abc_45749_n54), .Y(u1_acs_addr_pl1_13_) );
  AND2X2 AND2X2_3627 ( .A(u1_u0__abc_45749_n52_1), .B(u1_acs_addr_14_), .Y(u1_u0__abc_45749_n56_1) );
  AND2X2 AND2X2_3628 ( .A(u1_u0__abc_45749_n57), .B(u1_u0__abc_45749_n58), .Y(u1_acs_addr_pl1_14_) );
  AND2X2 AND2X2_3629 ( .A(u1_acs_addr_14_), .B(u1_acs_addr_15_), .Y(u1_u0__abc_45749_n61) );
  AND2X2 AND2X2_363 ( .A(u0__abc_49347_n1625), .B(u0__abc_49347_n1180_1_bF_buf5), .Y(u0__abc_49347_n1626) );
  AND2X2 AND2X2_3630 ( .A(u1_u0__abc_45749_n52_1), .B(u1_u0__abc_45749_n61), .Y(u1_u0__abc_45749_n62_1) );
  AND2X2 AND2X2_3631 ( .A(u1_u0__abc_45749_n60_1), .B(u1_u0__abc_45749_n63_1), .Y(u1_acs_addr_pl1_15_) );
  AND2X2 AND2X2_3632 ( .A(u1_u0__abc_45749_n62_1), .B(u1_acs_addr_16_), .Y(u1_u0__abc_45749_n65) );
  AND2X2 AND2X2_3633 ( .A(u1_u0__abc_45749_n66), .B(u1_u0__abc_45749_n67_1), .Y(u1_acs_addr_pl1_16_) );
  AND2X2 AND2X2_3634 ( .A(u1_acs_addr_16_), .B(u1_acs_addr_17_), .Y(u1_u0__abc_45749_n70_1) );
  AND2X2 AND2X2_3635 ( .A(u1_u0__abc_45749_n62_1), .B(u1_u0__abc_45749_n70_1), .Y(u1_u0__abc_45749_n71_1) );
  AND2X2 AND2X2_3636 ( .A(u1_u0__abc_45749_n69), .B(u1_u0__abc_45749_n72), .Y(u1_acs_addr_pl1_17_) );
  AND2X2 AND2X2_3637 ( .A(u1_u0__abc_45749_n71_1), .B(u1_acs_addr_18_), .Y(u1_u0__abc_45749_n74_1) );
  AND2X2 AND2X2_3638 ( .A(u1_u0__abc_45749_n75_1), .B(u1_u0__abc_45749_n76), .Y(u1_acs_addr_pl1_18_) );
  AND2X2 AND2X2_3639 ( .A(u1_acs_addr_18_), .B(u1_acs_addr_19_), .Y(u1_u0__abc_45749_n79_1) );
  AND2X2 AND2X2_364 ( .A(spec_req_cs_3_bF_buf2), .B(u0_tms3_18_), .Y(u0__abc_49347_n1627) );
  AND2X2 AND2X2_3640 ( .A(u1_u0__abc_45749_n70_1), .B(u1_u0__abc_45749_n79_1), .Y(u1_u0__abc_45749_n80) );
  AND2X2 AND2X2_3641 ( .A(u1_u0__abc_45749_n62_1), .B(u1_u0__abc_45749_n80), .Y(u1_u0__abc_45749_n81) );
  AND2X2 AND2X2_3642 ( .A(u1_u0__abc_45749_n78_1), .B(u1_u0__abc_45749_n82_1), .Y(u1_acs_addr_pl1_19_) );
  AND2X2 AND2X2_3643 ( .A(u1_u0__abc_45749_n81), .B(u1_acs_addr_20_), .Y(u1_u0__abc_45749_n84) );
  AND2X2 AND2X2_3644 ( .A(u1_u0__abc_45749_n85), .B(u1_u0__abc_45749_n86), .Y(u1_acs_addr_pl1_20_) );
  AND2X2 AND2X2_3645 ( .A(u1_acs_addr_20_), .B(u1_acs_addr_21_), .Y(u1_u0__abc_45749_n89) );
  AND2X2 AND2X2_3646 ( .A(u1_u0__abc_45749_n81), .B(u1_u0__abc_45749_n89), .Y(u1_u0__abc_45749_n90) );
  AND2X2 AND2X2_3647 ( .A(u1_u0__abc_45749_n88), .B(u1_u0__abc_45749_n91), .Y(u1_acs_addr_pl1_21_) );
  AND2X2 AND2X2_3648 ( .A(u1_u0__abc_45749_n90), .B(u1_acs_addr_22_), .Y(u1_u0__abc_45749_n93) );
  AND2X2 AND2X2_3649 ( .A(u1_u0__abc_45749_n94), .B(u1_u0__abc_45749_n95), .Y(u1_acs_addr_pl1_22_) );
  AND2X2 AND2X2_365 ( .A(u0__abc_49347_n1628), .B(u0__abc_49347_n1179_bF_buf5), .Y(u0__abc_49347_n1629) );
  AND2X2 AND2X2_3650 ( .A(u1_u0__abc_45749_n93), .B(u1_acs_addr_23_), .Y(u1_u0__abc_45749_n98) );
  AND2X2 AND2X2_3651 ( .A(u1_u0__abc_45749_n99), .B(u1_u0__abc_45749_n97), .Y(u1_acs_addr_pl1_23_) );
  AND2X2 AND2X2_3652 ( .A(u1_u0__abc_45749_n101), .B(u1_u0__abc_45749_n102), .Y(u1_acs_addr_pl1_12_) );
  AND2X2 AND2X2_3653 ( .A(u1_acs_addr_0_), .B(u1_acs_addr_1_), .Y(u1_u0__abc_45749_n104) );
  AND2X2 AND2X2_3654 ( .A(u1_u0__abc_45749_n105), .B(u1_u0__abc_45749_n106), .Y(u1_u0_out_r_1__FF_INPUT) );
  AND2X2 AND2X2_3655 ( .A(u1_u0__abc_45749_n104), .B(u1_acs_addr_2_), .Y(u1_u0__abc_45749_n108) );
  AND2X2 AND2X2_3656 ( .A(u1_u0__abc_45749_n109), .B(u1_u0__abc_45749_n110), .Y(u1_u0_out_r_2__FF_INPUT) );
  AND2X2 AND2X2_3657 ( .A(u1_u0__abc_45749_n108), .B(u1_acs_addr_3_), .Y(u1_u0__abc_45749_n112) );
  AND2X2 AND2X2_3658 ( .A(u1_u0__abc_45749_n113), .B(u1_u0__abc_45749_n114), .Y(u1_u0_out_r_3__FF_INPUT) );
  AND2X2 AND2X2_3659 ( .A(u1_u0__abc_45749_n112), .B(u1_acs_addr_4_), .Y(u1_u0__abc_45749_n116) );
  AND2X2 AND2X2_366 ( .A(spec_req_cs_2_bF_buf2), .B(u0_tms2_18_), .Y(u0__abc_49347_n1630) );
  AND2X2 AND2X2_3660 ( .A(u1_u0__abc_45749_n117), .B(u1_u0__abc_45749_n118), .Y(u1_u0_out_r_4__FF_INPUT) );
  AND2X2 AND2X2_3661 ( .A(u1_acs_addr_4_), .B(u1_acs_addr_5_), .Y(u1_u0__abc_45749_n121) );
  AND2X2 AND2X2_3662 ( .A(u1_u0__abc_45749_n112), .B(u1_u0__abc_45749_n121), .Y(u1_u0__abc_45749_n122) );
  AND2X2 AND2X2_3663 ( .A(u1_u0__abc_45749_n120), .B(u1_u0__abc_45749_n123), .Y(u1_u0_out_r_5__FF_INPUT) );
  AND2X2 AND2X2_3664 ( .A(u1_u0__abc_45749_n122), .B(u1_acs_addr_6_), .Y(u1_u0__abc_45749_n125) );
  AND2X2 AND2X2_3665 ( .A(u1_u0__abc_45749_n126), .B(u1_u0__abc_45749_n127), .Y(u1_u0_out_r_6__FF_INPUT) );
  AND2X2 AND2X2_3666 ( .A(u1_acs_addr_6_), .B(u1_acs_addr_7_), .Y(u1_u0__abc_45749_n130) );
  AND2X2 AND2X2_3667 ( .A(u1_u0__abc_45749_n121), .B(u1_u0__abc_45749_n130), .Y(u1_u0__abc_45749_n131) );
  AND2X2 AND2X2_3668 ( .A(u1_u0__abc_45749_n112), .B(u1_u0__abc_45749_n131), .Y(u1_u0__abc_45749_n132) );
  AND2X2 AND2X2_3669 ( .A(u1_u0__abc_45749_n129), .B(u1_u0__abc_45749_n133), .Y(u1_u0_out_r_7__FF_INPUT) );
  AND2X2 AND2X2_367 ( .A(u0__abc_49347_n1631), .B(u0__abc_49347_n1178_1_bF_buf5), .Y(u0__abc_49347_n1632_1) );
  AND2X2 AND2X2_3670 ( .A(u1_u0__abc_45749_n132), .B(u1_acs_addr_8_), .Y(u1_u0__abc_45749_n135) );
  AND2X2 AND2X2_3671 ( .A(u1_u0__abc_45749_n136), .B(u1_u0__abc_45749_n137), .Y(u1_u0_out_r_8__FF_INPUT) );
  AND2X2 AND2X2_3672 ( .A(u1_acs_addr_8_), .B(u1_acs_addr_9_), .Y(u1_u0__abc_45749_n140) );
  AND2X2 AND2X2_3673 ( .A(u1_u0__abc_45749_n132), .B(u1_u0__abc_45749_n140), .Y(u1_u0__abc_45749_n141) );
  AND2X2 AND2X2_3674 ( .A(u1_u0__abc_45749_n139), .B(u1_u0__abc_45749_n142), .Y(u1_u0_out_r_9__FF_INPUT) );
  AND2X2 AND2X2_3675 ( .A(u1_u0__abc_45749_n141), .B(u1_acs_addr_10_), .Y(u1_u0__abc_45749_n144) );
  AND2X2 AND2X2_3676 ( .A(u1_u0__abc_45749_n145), .B(u1_u0__abc_45749_n146), .Y(u1_u0_out_r_10__FF_INPUT) );
  AND2X2 AND2X2_3677 ( .A(u1_u0__abc_45749_n144), .B(u1_acs_addr_11_), .Y(u1_u0_out_r_12__FF_INPUT) );
  AND2X2 AND2X2_3678 ( .A(u1_u0__abc_45749_n149), .B(u1_u0__abc_45749_n150), .Y(u1_u0_out_r_11__FF_INPUT) );
  AND2X2 AND2X2_3679 ( .A(bank_set), .B(obct_cs_0_), .Y(u2_bank_set_0) );
  AND2X2 AND2X2_368 ( .A(spec_req_cs_1_bF_buf2), .B(u0_tms1_18_), .Y(u0__abc_49347_n1633_1) );
  AND2X2 AND2X2_3680 ( .A(bank_set), .B(obct_cs_1_), .Y(u2_bank_set_1) );
  AND2X2 AND2X2_3681 ( .A(bank_set), .B(obct_cs_2_), .Y(u2_bank_set_2) );
  AND2X2 AND2X2_3682 ( .A(bank_set), .B(obct_cs_3_), .Y(u2_bank_set_3) );
  AND2X2 AND2X2_3683 ( .A(bank_set), .B(obct_cs_4_), .Y(u2_bank_set_4) );
  AND2X2 AND2X2_3684 ( .A(bank_set), .B(obct_cs_5_), .Y(u2_bank_set_5) );
  AND2X2 AND2X2_3685 ( .A(obct_cs_0_), .B(bank_clr), .Y(u2_bank_clr_0) );
  AND2X2 AND2X2_3686 ( .A(obct_cs_1_), .B(bank_clr), .Y(u2_bank_clr_1) );
  AND2X2 AND2X2_3687 ( .A(obct_cs_2_), .B(bank_clr), .Y(u2_bank_clr_2) );
  AND2X2 AND2X2_3688 ( .A(obct_cs_3_), .B(bank_clr), .Y(u2_bank_clr_3) );
  AND2X2 AND2X2_3689 ( .A(obct_cs_4_), .B(bank_clr), .Y(u2_bank_clr_4) );
  AND2X2 AND2X2_369 ( .A(u0__abc_49347_n1175_bF_buf1), .B(u0__abc_49347_n1636), .Y(u0__abc_49347_n1637) );
  AND2X2 AND2X2_3690 ( .A(obct_cs_5_), .B(bank_clr), .Y(u2_bank_clr_5) );
  AND2X2 AND2X2_3691 ( .A(obct_cs_0_), .B(bank_clr_all), .Y(u2__abc_48153_n80) );
  AND2X2 AND2X2_3692 ( .A(obct_cs_1_), .B(bank_clr_all), .Y(u2__abc_48153_n82_1) );
  AND2X2 AND2X2_3693 ( .A(obct_cs_2_), .B(bank_clr_all), .Y(u2__abc_48153_n84_1) );
  AND2X2 AND2X2_3694 ( .A(obct_cs_3_), .B(bank_clr_all), .Y(u2__abc_48153_n86) );
  AND2X2 AND2X2_3695 ( .A(obct_cs_4_), .B(bank_clr_all), .Y(u2__abc_48153_n88_1) );
  AND2X2 AND2X2_3696 ( .A(obct_cs_5_), .B(bank_clr_all), .Y(u2__abc_48153_n90) );
  AND2X2 AND2X2_3697 ( .A(obct_cs_1_), .B(u2_bank_open_1), .Y(u2__abc_48153_n96) );
  AND2X2 AND2X2_3698 ( .A(obct_cs_0_), .B(u2_bank_open_0), .Y(u2__abc_48153_n97) );
  AND2X2 AND2X2_3699 ( .A(obct_cs_5_), .B(u2_bank_open_5), .Y(u2__abc_48153_n99) );
  AND2X2 AND2X2_37 ( .A(_abc_55805_n347), .B(_abc_55805_n348), .Y(tms_s_19_) );
  AND2X2 AND2X2_370 ( .A(u0__abc_49347_n1635), .B(u0__abc_49347_n1637), .Y(u0__abc_49347_n1638) );
  AND2X2 AND2X2_3700 ( .A(obct_cs_4_), .B(u2_bank_open_4), .Y(u2__abc_48153_n100) );
  AND2X2 AND2X2_3701 ( .A(obct_cs_3_), .B(u2_bank_open_3), .Y(u2__abc_48153_n103) );
  AND2X2 AND2X2_3702 ( .A(obct_cs_2_), .B(u2_bank_open_2), .Y(u2__abc_48153_n104) );
  AND2X2 AND2X2_3703 ( .A(obct_cs_7_), .B(1'b0), .Y(u2__abc_48153_n106) );
  AND2X2 AND2X2_3704 ( .A(obct_cs_6_), .B(1'b0), .Y(u2__abc_48153_n107) );
  AND2X2 AND2X2_3705 ( .A(obct_cs_1_), .B(u2_row_same_1), .Y(u2__abc_48153_n111) );
  AND2X2 AND2X2_3706 ( .A(obct_cs_0_), .B(u2_row_same_0), .Y(u2__abc_48153_n112) );
  AND2X2 AND2X2_3707 ( .A(obct_cs_5_), .B(u2_row_same_5), .Y(u2__abc_48153_n114) );
  AND2X2 AND2X2_3708 ( .A(obct_cs_4_), .B(u2_row_same_4), .Y(u2__abc_48153_n115) );
  AND2X2 AND2X2_3709 ( .A(obct_cs_3_), .B(u2_row_same_3), .Y(u2__abc_48153_n118) );
  AND2X2 AND2X2_371 ( .A(u0__abc_49347_n1176_1_bF_buf1), .B(sp_tms_19_), .Y(u0__abc_49347_n1640) );
  AND2X2 AND2X2_3710 ( .A(obct_cs_2_), .B(u2_row_same_2), .Y(u2__abc_48153_n119) );
  AND2X2 AND2X2_3711 ( .A(obct_cs_7_), .B(1'b0), .Y(u2__abc_48153_n121) );
  AND2X2 AND2X2_3712 ( .A(obct_cs_6_), .B(1'b0), .Y(u2__abc_48153_n122) );
  AND2X2 AND2X2_3713 ( .A(bank_adr_0_bF_buf1), .B(bank_adr_1_bF_buf1), .Y(u2_u0__abc_47660_n136) );
  AND2X2 AND2X2_3714 ( .A(u2_u0__abc_47660_n136), .B(u2_bank_set_0), .Y(u2_u0__abc_47660_n137) );
  AND2X2 AND2X2_3715 ( .A(u2_u0__abc_47660_n137_bF_buf3), .B(u2_u0__abc_47660_n139), .Y(u2_u0__abc_47660_n140) );
  AND2X2 AND2X2_3716 ( .A(u2_u0__abc_47660_n141), .B(u2_u0__abc_47660_n138), .Y(u2_u0_b3_last_row_0__FF_INPUT) );
  AND2X2 AND2X2_3717 ( .A(u2_u0__abc_47660_n137_bF_buf1), .B(u2_u0__abc_47660_n144), .Y(u2_u0__abc_47660_n145) );
  AND2X2 AND2X2_3718 ( .A(u2_u0__abc_47660_n146), .B(u2_u0__abc_47660_n143), .Y(u2_u0_b3_last_row_1__FF_INPUT) );
  AND2X2 AND2X2_3719 ( .A(u2_u0__abc_47660_n137_bF_buf4), .B(u2_u0__abc_47660_n149), .Y(u2_u0__abc_47660_n150) );
  AND2X2 AND2X2_372 ( .A(spec_req_cs_5_bF_buf1), .B(u0_tms5_19_), .Y(u0__abc_49347_n1641_1) );
  AND2X2 AND2X2_3720 ( .A(u2_u0__abc_47660_n151), .B(u2_u0__abc_47660_n148), .Y(u2_u0_b3_last_row_2__FF_INPUT) );
  AND2X2 AND2X2_3721 ( .A(u2_u0__abc_47660_n137_bF_buf2), .B(u2_u0__abc_47660_n154), .Y(u2_u0__abc_47660_n155) );
  AND2X2 AND2X2_3722 ( .A(u2_u0__abc_47660_n156), .B(u2_u0__abc_47660_n153), .Y(u2_u0_b3_last_row_3__FF_INPUT) );
  AND2X2 AND2X2_3723 ( .A(u2_u0__abc_47660_n137_bF_buf0), .B(u2_u0__abc_47660_n159), .Y(u2_u0__abc_47660_n160) );
  AND2X2 AND2X2_3724 ( .A(u2_u0__abc_47660_n161), .B(u2_u0__abc_47660_n158), .Y(u2_u0_b3_last_row_4__FF_INPUT) );
  AND2X2 AND2X2_3725 ( .A(u2_u0__abc_47660_n137_bF_buf3), .B(u2_u0__abc_47660_n164), .Y(u2_u0__abc_47660_n165) );
  AND2X2 AND2X2_3726 ( .A(u2_u0__abc_47660_n166), .B(u2_u0__abc_47660_n163), .Y(u2_u0_b3_last_row_5__FF_INPUT) );
  AND2X2 AND2X2_3727 ( .A(u2_u0__abc_47660_n137_bF_buf1), .B(u2_u0__abc_47660_n169), .Y(u2_u0__abc_47660_n170) );
  AND2X2 AND2X2_3728 ( .A(u2_u0__abc_47660_n171), .B(u2_u0__abc_47660_n168), .Y(u2_u0_b3_last_row_6__FF_INPUT) );
  AND2X2 AND2X2_3729 ( .A(u2_u0__abc_47660_n137_bF_buf4), .B(u2_u0__abc_47660_n174), .Y(u2_u0__abc_47660_n175) );
  AND2X2 AND2X2_373 ( .A(u0__abc_49347_n1643), .B(u0__abc_49347_n1185_bF_buf4), .Y(u0__abc_49347_n1644) );
  AND2X2 AND2X2_3730 ( .A(u2_u0__abc_47660_n176), .B(u2_u0__abc_47660_n173), .Y(u2_u0_b3_last_row_7__FF_INPUT) );
  AND2X2 AND2X2_3731 ( .A(u2_u0__abc_47660_n137_bF_buf2), .B(u2_u0__abc_47660_n179), .Y(u2_u0__abc_47660_n180) );
  AND2X2 AND2X2_3732 ( .A(u2_u0__abc_47660_n181), .B(u2_u0__abc_47660_n178), .Y(u2_u0_b3_last_row_8__FF_INPUT) );
  AND2X2 AND2X2_3733 ( .A(u2_u0__abc_47660_n137_bF_buf0), .B(u2_u0__abc_47660_n184), .Y(u2_u0__abc_47660_n185) );
  AND2X2 AND2X2_3734 ( .A(u2_u0__abc_47660_n186), .B(u2_u0__abc_47660_n183), .Y(u2_u0_b3_last_row_9__FF_INPUT) );
  AND2X2 AND2X2_3735 ( .A(u2_u0__abc_47660_n137_bF_buf3), .B(u2_u0__abc_47660_n189), .Y(u2_u0__abc_47660_n190) );
  AND2X2 AND2X2_3736 ( .A(u2_u0__abc_47660_n191), .B(u2_u0__abc_47660_n188), .Y(u2_u0_b3_last_row_10__FF_INPUT) );
  AND2X2 AND2X2_3737 ( .A(u2_u0__abc_47660_n137_bF_buf1), .B(u2_u0__abc_47660_n194), .Y(u2_u0__abc_47660_n195) );
  AND2X2 AND2X2_3738 ( .A(u2_u0__abc_47660_n196), .B(u2_u0__abc_47660_n193), .Y(u2_u0_b3_last_row_11__FF_INPUT) );
  AND2X2 AND2X2_3739 ( .A(u2_u0__abc_47660_n137_bF_buf4), .B(u2_u0__abc_47660_n199), .Y(u2_u0__abc_47660_n200) );
  AND2X2 AND2X2_374 ( .A(u0__abc_49347_n1644), .B(u0__abc_49347_n1642_1), .Y(u0__abc_49347_n1645) );
  AND2X2 AND2X2_3740 ( .A(u2_u0__abc_47660_n201), .B(u2_u0__abc_47660_n198), .Y(u2_u0_b3_last_row_12__FF_INPUT) );
  AND2X2 AND2X2_3741 ( .A(u2_u0__abc_47660_n203), .B(bank_adr_1_bF_buf0), .Y(u2_u0__abc_47660_n204) );
  AND2X2 AND2X2_3742 ( .A(u2_u0__abc_47660_n204), .B(u2_bank_set_0), .Y(u2_u0__abc_47660_n205) );
  AND2X2 AND2X2_3743 ( .A(u2_u0__abc_47660_n208), .B(u2_u0__abc_47660_n206), .Y(u2_u0_b2_last_row_0__FF_INPUT) );
  AND2X2 AND2X2_3744 ( .A(u2_u0__abc_47660_n211), .B(u2_u0__abc_47660_n210), .Y(u2_u0_b2_last_row_1__FF_INPUT) );
  AND2X2 AND2X2_3745 ( .A(u2_u0__abc_47660_n214), .B(u2_u0__abc_47660_n213), .Y(u2_u0_b2_last_row_2__FF_INPUT) );
  AND2X2 AND2X2_3746 ( .A(u2_u0__abc_47660_n217), .B(u2_u0__abc_47660_n216), .Y(u2_u0_b2_last_row_3__FF_INPUT) );
  AND2X2 AND2X2_3747 ( .A(u2_u0__abc_47660_n220), .B(u2_u0__abc_47660_n219), .Y(u2_u0_b2_last_row_4__FF_INPUT) );
  AND2X2 AND2X2_3748 ( .A(u2_u0__abc_47660_n223), .B(u2_u0__abc_47660_n222), .Y(u2_u0_b2_last_row_5__FF_INPUT) );
  AND2X2 AND2X2_3749 ( .A(u2_u0__abc_47660_n226), .B(u2_u0__abc_47660_n225), .Y(u2_u0_b2_last_row_6__FF_INPUT) );
  AND2X2 AND2X2_375 ( .A(u0__abc_49347_n1646), .B(u0__abc_49347_n1181_bF_buf4), .Y(u0__abc_49347_n1647) );
  AND2X2 AND2X2_3750 ( .A(u2_u0__abc_47660_n229), .B(u2_u0__abc_47660_n228), .Y(u2_u0_b2_last_row_7__FF_INPUT) );
  AND2X2 AND2X2_3751 ( .A(u2_u0__abc_47660_n232), .B(u2_u0__abc_47660_n231), .Y(u2_u0_b2_last_row_8__FF_INPUT) );
  AND2X2 AND2X2_3752 ( .A(u2_u0__abc_47660_n235), .B(u2_u0__abc_47660_n234), .Y(u2_u0_b2_last_row_9__FF_INPUT) );
  AND2X2 AND2X2_3753 ( .A(u2_u0__abc_47660_n238), .B(u2_u0__abc_47660_n237), .Y(u2_u0_b2_last_row_10__FF_INPUT) );
  AND2X2 AND2X2_3754 ( .A(u2_u0__abc_47660_n241), .B(u2_u0__abc_47660_n240), .Y(u2_u0_b2_last_row_11__FF_INPUT) );
  AND2X2 AND2X2_3755 ( .A(u2_u0__abc_47660_n244), .B(u2_u0__abc_47660_n243), .Y(u2_u0_b2_last_row_12__FF_INPUT) );
  AND2X2 AND2X2_3756 ( .A(u2_u0__abc_47660_n246), .B(bank_adr_0_bF_buf3), .Y(u2_u0__abc_47660_n247) );
  AND2X2 AND2X2_3757 ( .A(u2_u0__abc_47660_n247), .B(u2_bank_set_0), .Y(u2_u0__abc_47660_n248) );
  AND2X2 AND2X2_3758 ( .A(u2_u0__abc_47660_n251), .B(u2_u0__abc_47660_n249), .Y(u2_u0_b1_last_row_0__FF_INPUT) );
  AND2X2 AND2X2_3759 ( .A(u2_u0__abc_47660_n254), .B(u2_u0__abc_47660_n253), .Y(u2_u0_b1_last_row_1__FF_INPUT) );
  AND2X2 AND2X2_376 ( .A(spec_req_cs_4_bF_buf1), .B(u0_tms4_19_), .Y(u0__abc_49347_n1648) );
  AND2X2 AND2X2_3760 ( .A(u2_u0__abc_47660_n257), .B(u2_u0__abc_47660_n256), .Y(u2_u0_b1_last_row_2__FF_INPUT) );
  AND2X2 AND2X2_3761 ( .A(u2_u0__abc_47660_n260), .B(u2_u0__abc_47660_n259), .Y(u2_u0_b1_last_row_3__FF_INPUT) );
  AND2X2 AND2X2_3762 ( .A(u2_u0__abc_47660_n263), .B(u2_u0__abc_47660_n262), .Y(u2_u0_b1_last_row_4__FF_INPUT) );
  AND2X2 AND2X2_3763 ( .A(u2_u0__abc_47660_n266), .B(u2_u0__abc_47660_n265), .Y(u2_u0_b1_last_row_5__FF_INPUT) );
  AND2X2 AND2X2_3764 ( .A(u2_u0__abc_47660_n269), .B(u2_u0__abc_47660_n268), .Y(u2_u0_b1_last_row_6__FF_INPUT) );
  AND2X2 AND2X2_3765 ( .A(u2_u0__abc_47660_n272), .B(u2_u0__abc_47660_n271), .Y(u2_u0_b1_last_row_7__FF_INPUT) );
  AND2X2 AND2X2_3766 ( .A(u2_u0__abc_47660_n275_1), .B(u2_u0__abc_47660_n274), .Y(u2_u0_b1_last_row_8__FF_INPUT) );
  AND2X2 AND2X2_3767 ( .A(u2_u0__abc_47660_n278_1), .B(u2_u0__abc_47660_n277), .Y(u2_u0_b1_last_row_9__FF_INPUT) );
  AND2X2 AND2X2_3768 ( .A(u2_u0__abc_47660_n281), .B(u2_u0__abc_47660_n280), .Y(u2_u0_b1_last_row_10__FF_INPUT) );
  AND2X2 AND2X2_3769 ( .A(u2_u0__abc_47660_n284), .B(u2_u0__abc_47660_n283_1), .Y(u2_u0_b1_last_row_11__FF_INPUT) );
  AND2X2 AND2X2_377 ( .A(u0__abc_49347_n1649), .B(u0__abc_49347_n1180_1_bF_buf4), .Y(u0__abc_49347_n1650_1) );
  AND2X2 AND2X2_3770 ( .A(u2_u0__abc_47660_n287_1), .B(u2_u0__abc_47660_n286_1), .Y(u2_u0_b1_last_row_12__FF_INPUT) );
  AND2X2 AND2X2_3771 ( .A(u2_u0__abc_47660_n203), .B(u2_u0__abc_47660_n246), .Y(u2_u0__abc_47660_n289) );
  AND2X2 AND2X2_3772 ( .A(u2_u0__abc_47660_n289), .B(u2_bank_set_0), .Y(u2_u0__abc_47660_n290_1) );
  AND2X2 AND2X2_3773 ( .A(u2_u0__abc_47660_n293), .B(u2_u0__abc_47660_n291), .Y(u2_u0_b0_last_row_0__FF_INPUT) );
  AND2X2 AND2X2_3774 ( .A(u2_u0__abc_47660_n296_1), .B(u2_u0__abc_47660_n295), .Y(u2_u0_b0_last_row_1__FF_INPUT) );
  AND2X2 AND2X2_3775 ( .A(u2_u0__abc_47660_n299), .B(u2_u0__abc_47660_n298), .Y(u2_u0_b0_last_row_2__FF_INPUT) );
  AND2X2 AND2X2_3776 ( .A(u2_u0__abc_47660_n302), .B(u2_u0__abc_47660_n301), .Y(u2_u0_b0_last_row_3__FF_INPUT) );
  AND2X2 AND2X2_3777 ( .A(u2_u0__abc_47660_n305_1), .B(u2_u0__abc_47660_n304_1), .Y(u2_u0_b0_last_row_4__FF_INPUT) );
  AND2X2 AND2X2_3778 ( .A(u2_u0__abc_47660_n308), .B(u2_u0__abc_47660_n307), .Y(u2_u0_b0_last_row_5__FF_INPUT) );
  AND2X2 AND2X2_3779 ( .A(u2_u0__abc_47660_n311), .B(u2_u0__abc_47660_n310), .Y(u2_u0_b0_last_row_6__FF_INPUT) );
  AND2X2 AND2X2_378 ( .A(spec_req_cs_3_bF_buf1), .B(u0_tms3_19_), .Y(u0__abc_49347_n1651_1) );
  AND2X2 AND2X2_3780 ( .A(u2_u0__abc_47660_n314), .B(u2_u0__abc_47660_n313), .Y(u2_u0_b0_last_row_7__FF_INPUT) );
  AND2X2 AND2X2_3781 ( .A(u2_u0__abc_47660_n317), .B(u2_u0__abc_47660_n316), .Y(u2_u0_b0_last_row_8__FF_INPUT) );
  AND2X2 AND2X2_3782 ( .A(u2_u0__abc_47660_n320), .B(u2_u0__abc_47660_n319), .Y(u2_u0_b0_last_row_9__FF_INPUT) );
  AND2X2 AND2X2_3783 ( .A(u2_u0__abc_47660_n323), .B(u2_u0__abc_47660_n322), .Y(u2_u0_b0_last_row_10__FF_INPUT) );
  AND2X2 AND2X2_3784 ( .A(u2_u0__abc_47660_n326), .B(u2_u0__abc_47660_n325), .Y(u2_u0_b0_last_row_11__FF_INPUT) );
  AND2X2 AND2X2_3785 ( .A(u2_u0__abc_47660_n329), .B(u2_u0__abc_47660_n328), .Y(u2_u0_b0_last_row_12__FF_INPUT) );
  AND2X2 AND2X2_3786 ( .A(u2_u0__abc_47660_n334), .B(u2_u0__abc_47660_n335), .Y(u2_u0__abc_47660_n336) );
  AND2X2 AND2X2_3787 ( .A(u2_u0__abc_47660_n336), .B(u2_u0__abc_47660_n332), .Y(u2_u0__abc_47660_n337) );
  AND2X2 AND2X2_3788 ( .A(u2_u0__abc_47660_n338), .B(u2_u0__abc_47660_n340), .Y(u2_u0__abc_47660_n341) );
  AND2X2 AND2X2_3789 ( .A(u2_u0__abc_47660_n342), .B(u2_u0__abc_47660_n344), .Y(u2_u0__abc_47660_n345) );
  AND2X2 AND2X2_379 ( .A(u0__abc_49347_n1652), .B(u0__abc_49347_n1179_bF_buf4), .Y(u0__abc_49347_n1653) );
  AND2X2 AND2X2_3790 ( .A(u2_u0__abc_47660_n341), .B(u2_u0__abc_47660_n345), .Y(u2_u0__abc_47660_n346) );
  AND2X2 AND2X2_3791 ( .A(u2_u0__abc_47660_n346), .B(u2_u0__abc_47660_n337), .Y(u2_u0__abc_47660_n347) );
  AND2X2 AND2X2_3792 ( .A(u2_u0__abc_47660_n348), .B(u2_u0__abc_47660_n289), .Y(u2_u0__abc_47660_n349) );
  AND2X2 AND2X2_3793 ( .A(u2_u0__abc_47660_n350), .B(u2_u0__abc_47660_n352), .Y(u2_u0__abc_47660_n353) );
  AND2X2 AND2X2_3794 ( .A(u2_u0__abc_47660_n353), .B(u2_u0__abc_47660_n349), .Y(u2_u0__abc_47660_n354) );
  AND2X2 AND2X2_3795 ( .A(u2_u0__abc_47660_n356), .B(u2_u0__abc_47660_n357), .Y(u2_u0__abc_47660_n358) );
  AND2X2 AND2X2_3796 ( .A(u2_u0__abc_47660_n359), .B(u2_u0__abc_47660_n361), .Y(u2_u0__abc_47660_n362) );
  AND2X2 AND2X2_3797 ( .A(u2_u0__abc_47660_n358), .B(u2_u0__abc_47660_n362), .Y(u2_u0__abc_47660_n363) );
  AND2X2 AND2X2_3798 ( .A(u2_u0__abc_47660_n363), .B(u2_u0__abc_47660_n354), .Y(u2_u0__abc_47660_n364) );
  AND2X2 AND2X2_3799 ( .A(u2_u0__abc_47660_n347), .B(u2_u0__abc_47660_n364), .Y(u2_u0__abc_47660_n365) );
  AND2X2 AND2X2_38 ( .A(_abc_55805_n350), .B(_abc_55805_n351), .Y(tms_s_20_) );
  AND2X2 AND2X2_380 ( .A(spec_req_cs_2_bF_buf1), .B(u0_tms2_19_), .Y(u0__abc_49347_n1654) );
  AND2X2 AND2X2_3800 ( .A(u2_u0__abc_47660_n367), .B(u2_u0__abc_47660_n368), .Y(u2_u0__abc_47660_n369) );
  AND2X2 AND2X2_3801 ( .A(row_adr_8_bF_buf0), .B(u2_u0_b0_last_row_8_), .Y(u2_u0__abc_47660_n370) );
  AND2X2 AND2X2_3802 ( .A(u2_u0__abc_47660_n179), .B(u2_u0__abc_47660_n371), .Y(u2_u0__abc_47660_n372) );
  AND2X2 AND2X2_3803 ( .A(u2_u0__abc_47660_n369), .B(u2_u0__abc_47660_n373), .Y(u2_u0__abc_47660_n374) );
  AND2X2 AND2X2_3804 ( .A(u2_u0__abc_47660_n375), .B(u2_u0__abc_47660_n377), .Y(u2_u0__abc_47660_n378) );
  AND2X2 AND2X2_3805 ( .A(u2_u0__abc_47660_n380), .B(u2_u0__abc_47660_n381), .Y(u2_u0__abc_47660_n382) );
  AND2X2 AND2X2_3806 ( .A(u2_u0__abc_47660_n378), .B(u2_u0__abc_47660_n382), .Y(u2_u0__abc_47660_n383) );
  AND2X2 AND2X2_3807 ( .A(u2_u0__abc_47660_n385), .B(u2_u0__abc_47660_n386), .Y(u2_u0__abc_47660_n387) );
  AND2X2 AND2X2_3808 ( .A(row_adr_6_bF_buf0), .B(u2_u0_b0_last_row_6_), .Y(u2_u0__abc_47660_n388) );
  AND2X2 AND2X2_3809 ( .A(u2_u0__abc_47660_n169), .B(u2_u0__abc_47660_n389), .Y(u2_u0__abc_47660_n390) );
  AND2X2 AND2X2_381 ( .A(u0__abc_49347_n1655), .B(u0__abc_49347_n1178_1_bF_buf4), .Y(u0__abc_49347_n1656) );
  AND2X2 AND2X2_3810 ( .A(u2_u0__abc_47660_n387), .B(u2_u0__abc_47660_n391), .Y(u2_u0__abc_47660_n392) );
  AND2X2 AND2X2_3811 ( .A(u2_u0__abc_47660_n383), .B(u2_u0__abc_47660_n392), .Y(u2_u0__abc_47660_n393) );
  AND2X2 AND2X2_3812 ( .A(u2_u0__abc_47660_n393), .B(u2_u0__abc_47660_n374), .Y(u2_u0__abc_47660_n394) );
  AND2X2 AND2X2_3813 ( .A(u2_u0__abc_47660_n365), .B(u2_u0__abc_47660_n394), .Y(u2_u0__abc_47660_n395) );
  AND2X2 AND2X2_3814 ( .A(u2_u0__abc_47660_n399), .B(u2_u0__abc_47660_n400), .Y(u2_u0__abc_47660_n401) );
  AND2X2 AND2X2_3815 ( .A(u2_u0__abc_47660_n401), .B(u2_u0__abc_47660_n397), .Y(u2_u0__abc_47660_n402) );
  AND2X2 AND2X2_3816 ( .A(u2_u0__abc_47660_n403), .B(u2_u0__abc_47660_n405), .Y(u2_u0__abc_47660_n406) );
  AND2X2 AND2X2_3817 ( .A(u2_u0__abc_47660_n407), .B(u2_u0__abc_47660_n409), .Y(u2_u0__abc_47660_n410) );
  AND2X2 AND2X2_3818 ( .A(u2_u0__abc_47660_n406), .B(u2_u0__abc_47660_n410), .Y(u2_u0__abc_47660_n411) );
  AND2X2 AND2X2_3819 ( .A(u2_u0__abc_47660_n411), .B(u2_u0__abc_47660_n402), .Y(u2_u0__abc_47660_n412) );
  AND2X2 AND2X2_382 ( .A(spec_req_cs_1_bF_buf1), .B(u0_tms1_19_), .Y(u0__abc_49347_n1657) );
  AND2X2 AND2X2_3820 ( .A(u2_u0__abc_47660_n413), .B(u2_u0__abc_47660_n204), .Y(u2_u0__abc_47660_n414) );
  AND2X2 AND2X2_3821 ( .A(u2_u0__abc_47660_n415), .B(u2_u0__abc_47660_n417), .Y(u2_u0__abc_47660_n418) );
  AND2X2 AND2X2_3822 ( .A(u2_u0__abc_47660_n418), .B(u2_u0__abc_47660_n414), .Y(u2_u0__abc_47660_n419) );
  AND2X2 AND2X2_3823 ( .A(u2_u0__abc_47660_n421), .B(u2_u0__abc_47660_n422), .Y(u2_u0__abc_47660_n423) );
  AND2X2 AND2X2_3824 ( .A(u2_u0__abc_47660_n424), .B(u2_u0__abc_47660_n426), .Y(u2_u0__abc_47660_n427) );
  AND2X2 AND2X2_3825 ( .A(u2_u0__abc_47660_n423), .B(u2_u0__abc_47660_n427), .Y(u2_u0__abc_47660_n428) );
  AND2X2 AND2X2_3826 ( .A(u2_u0__abc_47660_n428), .B(u2_u0__abc_47660_n419), .Y(u2_u0__abc_47660_n429) );
  AND2X2 AND2X2_3827 ( .A(u2_u0__abc_47660_n412), .B(u2_u0__abc_47660_n429), .Y(u2_u0__abc_47660_n430) );
  AND2X2 AND2X2_3828 ( .A(u2_u0__abc_47660_n432), .B(u2_u0__abc_47660_n433), .Y(u2_u0__abc_47660_n434) );
  AND2X2 AND2X2_3829 ( .A(row_adr_8_bF_buf6), .B(u2_u0_b2_last_row_8_), .Y(u2_u0__abc_47660_n435) );
  AND2X2 AND2X2_383 ( .A(u0__abc_49347_n1175_bF_buf0), .B(u0__abc_49347_n1660_1), .Y(u0__abc_49347_n1661) );
  AND2X2 AND2X2_3830 ( .A(u2_u0__abc_47660_n179), .B(u2_u0__abc_47660_n436), .Y(u2_u0__abc_47660_n437) );
  AND2X2 AND2X2_3831 ( .A(u2_u0__abc_47660_n434), .B(u2_u0__abc_47660_n438), .Y(u2_u0__abc_47660_n439) );
  AND2X2 AND2X2_3832 ( .A(u2_u0__abc_47660_n440), .B(u2_u0__abc_47660_n442), .Y(u2_u0__abc_47660_n443) );
  AND2X2 AND2X2_3833 ( .A(u2_u0__abc_47660_n445), .B(u2_u0__abc_47660_n446), .Y(u2_u0__abc_47660_n447) );
  AND2X2 AND2X2_3834 ( .A(u2_u0__abc_47660_n443), .B(u2_u0__abc_47660_n447), .Y(u2_u0__abc_47660_n448) );
  AND2X2 AND2X2_3835 ( .A(u2_u0__abc_47660_n450), .B(u2_u0__abc_47660_n451), .Y(u2_u0__abc_47660_n452) );
  AND2X2 AND2X2_3836 ( .A(row_adr_6_bF_buf6), .B(u2_u0_b2_last_row_6_), .Y(u2_u0__abc_47660_n453) );
  AND2X2 AND2X2_3837 ( .A(u2_u0__abc_47660_n169), .B(u2_u0__abc_47660_n454), .Y(u2_u0__abc_47660_n455) );
  AND2X2 AND2X2_3838 ( .A(u2_u0__abc_47660_n452), .B(u2_u0__abc_47660_n456), .Y(u2_u0__abc_47660_n457) );
  AND2X2 AND2X2_3839 ( .A(u2_u0__abc_47660_n448), .B(u2_u0__abc_47660_n457), .Y(u2_u0__abc_47660_n458) );
  AND2X2 AND2X2_384 ( .A(u0__abc_49347_n1659_1), .B(u0__abc_49347_n1661), .Y(u0__abc_49347_n1662) );
  AND2X2 AND2X2_3840 ( .A(u2_u0__abc_47660_n458), .B(u2_u0__abc_47660_n439), .Y(u2_u0__abc_47660_n459) );
  AND2X2 AND2X2_3841 ( .A(u2_u0__abc_47660_n430), .B(u2_u0__abc_47660_n459), .Y(u2_u0__abc_47660_n460) );
  AND2X2 AND2X2_3842 ( .A(u2_u0__abc_47660_n465), .B(u2_u0__abc_47660_n466), .Y(u2_u0__abc_47660_n467) );
  AND2X2 AND2X2_3843 ( .A(u2_u0__abc_47660_n467), .B(u2_u0__abc_47660_n463), .Y(u2_u0__abc_47660_n468) );
  AND2X2 AND2X2_3844 ( .A(u2_u0__abc_47660_n469), .B(u2_u0__abc_47660_n471), .Y(u2_u0__abc_47660_n472) );
  AND2X2 AND2X2_3845 ( .A(u2_u0__abc_47660_n473), .B(u2_u0__abc_47660_n475), .Y(u2_u0__abc_47660_n476) );
  AND2X2 AND2X2_3846 ( .A(u2_u0__abc_47660_n472), .B(u2_u0__abc_47660_n476), .Y(u2_u0__abc_47660_n477) );
  AND2X2 AND2X2_3847 ( .A(u2_u0__abc_47660_n477), .B(u2_u0__abc_47660_n468), .Y(u2_u0__abc_47660_n478) );
  AND2X2 AND2X2_3848 ( .A(u2_u0__abc_47660_n479), .B(u2_u0__abc_47660_n247), .Y(u2_u0__abc_47660_n480) );
  AND2X2 AND2X2_3849 ( .A(u2_u0__abc_47660_n481), .B(u2_u0__abc_47660_n483), .Y(u2_u0__abc_47660_n484) );
  AND2X2 AND2X2_385 ( .A(u0__abc_49347_n1176_1_bF_buf0), .B(sp_tms_20_), .Y(u0__abc_49347_n1664) );
  AND2X2 AND2X2_3850 ( .A(u2_u0__abc_47660_n484), .B(u2_u0__abc_47660_n480), .Y(u2_u0__abc_47660_n485) );
  AND2X2 AND2X2_3851 ( .A(u2_u0__abc_47660_n487), .B(u2_u0__abc_47660_n488), .Y(u2_u0__abc_47660_n489) );
  AND2X2 AND2X2_3852 ( .A(u2_u0__abc_47660_n490), .B(u2_u0__abc_47660_n492), .Y(u2_u0__abc_47660_n493) );
  AND2X2 AND2X2_3853 ( .A(u2_u0__abc_47660_n489), .B(u2_u0__abc_47660_n493), .Y(u2_u0__abc_47660_n494) );
  AND2X2 AND2X2_3854 ( .A(u2_u0__abc_47660_n494), .B(u2_u0__abc_47660_n485), .Y(u2_u0__abc_47660_n495) );
  AND2X2 AND2X2_3855 ( .A(u2_u0__abc_47660_n478), .B(u2_u0__abc_47660_n495), .Y(u2_u0__abc_47660_n496) );
  AND2X2 AND2X2_3856 ( .A(u2_u0__abc_47660_n498), .B(u2_u0__abc_47660_n499), .Y(u2_u0__abc_47660_n500) );
  AND2X2 AND2X2_3857 ( .A(row_adr_8_bF_buf5), .B(u2_u0_b1_last_row_8_), .Y(u2_u0__abc_47660_n501) );
  AND2X2 AND2X2_3858 ( .A(u2_u0__abc_47660_n179), .B(u2_u0__abc_47660_n502), .Y(u2_u0__abc_47660_n503) );
  AND2X2 AND2X2_3859 ( .A(u2_u0__abc_47660_n500), .B(u2_u0__abc_47660_n504), .Y(u2_u0__abc_47660_n505) );
  AND2X2 AND2X2_386 ( .A(spec_req_cs_5_bF_buf0), .B(u0_tms5_20_), .Y(u0__abc_49347_n1665) );
  AND2X2 AND2X2_3860 ( .A(u2_u0__abc_47660_n506), .B(u2_u0__abc_47660_n508), .Y(u2_u0__abc_47660_n509) );
  AND2X2 AND2X2_3861 ( .A(u2_u0__abc_47660_n511), .B(u2_u0__abc_47660_n512), .Y(u2_u0__abc_47660_n513) );
  AND2X2 AND2X2_3862 ( .A(u2_u0__abc_47660_n509), .B(u2_u0__abc_47660_n513), .Y(u2_u0__abc_47660_n514) );
  AND2X2 AND2X2_3863 ( .A(u2_u0__abc_47660_n516), .B(u2_u0__abc_47660_n517), .Y(u2_u0__abc_47660_n518) );
  AND2X2 AND2X2_3864 ( .A(row_adr_6_bF_buf5), .B(u2_u0_b1_last_row_6_), .Y(u2_u0__abc_47660_n519) );
  AND2X2 AND2X2_3865 ( .A(u2_u0__abc_47660_n169), .B(u2_u0__abc_47660_n520), .Y(u2_u0__abc_47660_n521) );
  AND2X2 AND2X2_3866 ( .A(u2_u0__abc_47660_n518), .B(u2_u0__abc_47660_n522), .Y(u2_u0__abc_47660_n523) );
  AND2X2 AND2X2_3867 ( .A(u2_u0__abc_47660_n514), .B(u2_u0__abc_47660_n523), .Y(u2_u0__abc_47660_n524) );
  AND2X2 AND2X2_3868 ( .A(u2_u0__abc_47660_n524), .B(u2_u0__abc_47660_n505), .Y(u2_u0__abc_47660_n525) );
  AND2X2 AND2X2_3869 ( .A(u2_u0__abc_47660_n496), .B(u2_u0__abc_47660_n525), .Y(u2_u0__abc_47660_n526) );
  AND2X2 AND2X2_387 ( .A(u0__abc_49347_n1667), .B(u0__abc_49347_n1185_bF_buf3), .Y(u0__abc_49347_n1668_1) );
  AND2X2 AND2X2_3870 ( .A(u2_u0__abc_47660_n529), .B(u2_u0__abc_47660_n530), .Y(u2_u0__abc_47660_n531) );
  AND2X2 AND2X2_3871 ( .A(u2_u0__abc_47660_n531), .B(u2_u0__abc_47660_n528), .Y(u2_u0__abc_47660_n532) );
  AND2X2 AND2X2_3872 ( .A(u2_u0__abc_47660_n533), .B(u2_u0__abc_47660_n535), .Y(u2_u0__abc_47660_n536) );
  AND2X2 AND2X2_3873 ( .A(u2_u0__abc_47660_n537), .B(u2_u0__abc_47660_n539), .Y(u2_u0__abc_47660_n540) );
  AND2X2 AND2X2_3874 ( .A(u2_u0__abc_47660_n536), .B(u2_u0__abc_47660_n540), .Y(u2_u0__abc_47660_n541) );
  AND2X2 AND2X2_3875 ( .A(u2_u0__abc_47660_n541), .B(u2_u0__abc_47660_n532), .Y(u2_u0__abc_47660_n542) );
  AND2X2 AND2X2_3876 ( .A(u2_u0__abc_47660_n543), .B(u2_u0__abc_47660_n545), .Y(u2_u0__abc_47660_n546) );
  AND2X2 AND2X2_3877 ( .A(u2_u0__abc_47660_n548), .B(u2_u0__abc_47660_n136), .Y(u2_u0__abc_47660_n549) );
  AND2X2 AND2X2_3878 ( .A(u2_u0__abc_47660_n546), .B(u2_u0__abc_47660_n549), .Y(u2_u0__abc_47660_n550) );
  AND2X2 AND2X2_3879 ( .A(u2_u0__abc_47660_n552), .B(u2_u0__abc_47660_n553), .Y(u2_u0__abc_47660_n554) );
  AND2X2 AND2X2_388 ( .A(u0__abc_49347_n1668_1), .B(u0__abc_49347_n1666), .Y(u0__abc_49347_n1669_1) );
  AND2X2 AND2X2_3880 ( .A(u2_u0__abc_47660_n556), .B(u2_u0__abc_47660_n557), .Y(u2_u0__abc_47660_n558) );
  AND2X2 AND2X2_3881 ( .A(u2_u0__abc_47660_n554), .B(u2_u0__abc_47660_n558), .Y(u2_u0__abc_47660_n559) );
  AND2X2 AND2X2_3882 ( .A(u2_u0__abc_47660_n559), .B(u2_u0__abc_47660_n550), .Y(u2_u0__abc_47660_n560) );
  AND2X2 AND2X2_3883 ( .A(u2_u0__abc_47660_n542), .B(u2_u0__abc_47660_n560), .Y(u2_u0__abc_47660_n561) );
  AND2X2 AND2X2_3884 ( .A(u2_u0__abc_47660_n562), .B(u2_u0__abc_47660_n564), .Y(u2_u0__abc_47660_n565) );
  AND2X2 AND2X2_3885 ( .A(u2_u0__abc_47660_n567), .B(u2_u0__abc_47660_n568), .Y(u2_u0__abc_47660_n569) );
  AND2X2 AND2X2_3886 ( .A(u2_u0__abc_47660_n565), .B(u2_u0__abc_47660_n569), .Y(u2_u0__abc_47660_n570) );
  AND2X2 AND2X2_3887 ( .A(u2_u0__abc_47660_n571), .B(u2_u0__abc_47660_n573), .Y(u2_u0__abc_47660_n574) );
  AND2X2 AND2X2_3888 ( .A(u2_u0__abc_47660_n576), .B(u2_u0__abc_47660_n577), .Y(u2_u0__abc_47660_n578) );
  AND2X2 AND2X2_3889 ( .A(u2_u0__abc_47660_n574), .B(u2_u0__abc_47660_n578), .Y(u2_u0__abc_47660_n579) );
  AND2X2 AND2X2_389 ( .A(u0__abc_49347_n1670), .B(u0__abc_49347_n1181_bF_buf3), .Y(u0__abc_49347_n1671) );
  AND2X2 AND2X2_3890 ( .A(u2_u0__abc_47660_n580), .B(u2_u0__abc_47660_n582), .Y(u2_u0__abc_47660_n583) );
  AND2X2 AND2X2_3891 ( .A(u2_u0__abc_47660_n584), .B(u2_u0__abc_47660_n586), .Y(u2_u0__abc_47660_n587) );
  AND2X2 AND2X2_3892 ( .A(u2_u0__abc_47660_n583), .B(u2_u0__abc_47660_n587), .Y(u2_u0__abc_47660_n588) );
  AND2X2 AND2X2_3893 ( .A(u2_u0__abc_47660_n579), .B(u2_u0__abc_47660_n588), .Y(u2_u0__abc_47660_n589) );
  AND2X2 AND2X2_3894 ( .A(u2_u0__abc_47660_n589), .B(u2_u0__abc_47660_n570), .Y(u2_u0__abc_47660_n590) );
  AND2X2 AND2X2_3895 ( .A(u2_u0__abc_47660_n561), .B(u2_u0__abc_47660_n590), .Y(u2_u0__abc_47660_n591) );
  AND2X2 AND2X2_3896 ( .A(u2_u0__abc_47660_n289), .B(u2_u0_bank0_open), .Y(u2_u0__abc_47660_n594) );
  AND2X2 AND2X2_3897 ( .A(u2_u0__abc_47660_n204), .B(u2_u0_bank2_open), .Y(u2_u0__abc_47660_n595) );
  AND2X2 AND2X2_3898 ( .A(u2_u0__abc_47660_n136), .B(u2_u0_bank3_open), .Y(u2_u0__abc_47660_n597) );
  AND2X2 AND2X2_3899 ( .A(u2_u0__abc_47660_n247), .B(u2_u0_bank1_open), .Y(u2_u0__abc_47660_n598) );
  AND2X2 AND2X2_39 ( .A(_abc_55805_n353), .B(_abc_55805_n354), .Y(tms_s_21_) );
  AND2X2 AND2X2_390 ( .A(spec_req_cs_4_bF_buf0), .B(u0_tms4_20_), .Y(u0__abc_49347_n1672) );
  AND2X2 AND2X2_3900 ( .A(u2_u0__abc_47660_n136), .B(u2_bank_clr_0), .Y(u2_u0__abc_47660_n604) );
  AND2X2 AND2X2_3901 ( .A(u2_u0__abc_47660_n606), .B(u2_u0_bank3_open), .Y(u2_u0__abc_47660_n607) );
  AND2X2 AND2X2_3902 ( .A(u2_u0__abc_47660_n605), .B(u2_u0__abc_47660_n607), .Y(u2_u0__abc_47660_n608) );
  AND2X2 AND2X2_3903 ( .A(u2_u0__abc_47660_n606), .B(u2_u0_bank2_open), .Y(u2_u0__abc_47660_n613) );
  AND2X2 AND2X2_3904 ( .A(u2_u0__abc_47660_n612), .B(u2_u0__abc_47660_n613), .Y(u2_u0__abc_47660_n614) );
  AND2X2 AND2X2_3905 ( .A(u2_u0__abc_47660_n606), .B(u2_u0_bank1_open), .Y(u2_u0__abc_47660_n618) );
  AND2X2 AND2X2_3906 ( .A(u2_u0__abc_47660_n617), .B(u2_u0__abc_47660_n618), .Y(u2_u0__abc_47660_n619) );
  AND2X2 AND2X2_3907 ( .A(u2_u0__abc_47660_n606), .B(u2_u0_bank0_open), .Y(u2_u0__abc_47660_n623) );
  AND2X2 AND2X2_3908 ( .A(u2_u0__abc_47660_n622), .B(u2_u0__abc_47660_n623), .Y(u2_u0__abc_47660_n624) );
  AND2X2 AND2X2_3909 ( .A(bank_adr_0_bF_buf2), .B(bank_adr_1_bF_buf2), .Y(u2_u1__abc_47660_n136) );
  AND2X2 AND2X2_391 ( .A(u0__abc_49347_n1673), .B(u0__abc_49347_n1180_1_bF_buf3), .Y(u0__abc_49347_n1674) );
  AND2X2 AND2X2_3910 ( .A(u2_u1__abc_47660_n136), .B(u2_bank_set_1), .Y(u2_u1__abc_47660_n137) );
  AND2X2 AND2X2_3911 ( .A(u2_u1__abc_47660_n137_bF_buf3), .B(u2_u1__abc_47660_n139), .Y(u2_u1__abc_47660_n140) );
  AND2X2 AND2X2_3912 ( .A(u2_u1__abc_47660_n141), .B(u2_u1__abc_47660_n138), .Y(u2_u1_b3_last_row_0__FF_INPUT) );
  AND2X2 AND2X2_3913 ( .A(u2_u1__abc_47660_n137_bF_buf1), .B(u2_u1__abc_47660_n144), .Y(u2_u1__abc_47660_n145) );
  AND2X2 AND2X2_3914 ( .A(u2_u1__abc_47660_n146), .B(u2_u1__abc_47660_n143), .Y(u2_u1_b3_last_row_1__FF_INPUT) );
  AND2X2 AND2X2_3915 ( .A(u2_u1__abc_47660_n137_bF_buf4), .B(u2_u1__abc_47660_n149), .Y(u2_u1__abc_47660_n150) );
  AND2X2 AND2X2_3916 ( .A(u2_u1__abc_47660_n151), .B(u2_u1__abc_47660_n148), .Y(u2_u1_b3_last_row_2__FF_INPUT) );
  AND2X2 AND2X2_3917 ( .A(u2_u1__abc_47660_n137_bF_buf2), .B(u2_u1__abc_47660_n154), .Y(u2_u1__abc_47660_n155) );
  AND2X2 AND2X2_3918 ( .A(u2_u1__abc_47660_n156), .B(u2_u1__abc_47660_n153), .Y(u2_u1_b3_last_row_3__FF_INPUT) );
  AND2X2 AND2X2_3919 ( .A(u2_u1__abc_47660_n137_bF_buf0), .B(u2_u1__abc_47660_n159), .Y(u2_u1__abc_47660_n160) );
  AND2X2 AND2X2_392 ( .A(spec_req_cs_3_bF_buf0), .B(u0_tms3_20_), .Y(u0__abc_49347_n1675) );
  AND2X2 AND2X2_3920 ( .A(u2_u1__abc_47660_n161), .B(u2_u1__abc_47660_n158), .Y(u2_u1_b3_last_row_4__FF_INPUT) );
  AND2X2 AND2X2_3921 ( .A(u2_u1__abc_47660_n137_bF_buf3), .B(u2_u1__abc_47660_n164), .Y(u2_u1__abc_47660_n165) );
  AND2X2 AND2X2_3922 ( .A(u2_u1__abc_47660_n166), .B(u2_u1__abc_47660_n163), .Y(u2_u1_b3_last_row_5__FF_INPUT) );
  AND2X2 AND2X2_3923 ( .A(u2_u1__abc_47660_n137_bF_buf1), .B(u2_u1__abc_47660_n169), .Y(u2_u1__abc_47660_n170) );
  AND2X2 AND2X2_3924 ( .A(u2_u1__abc_47660_n171), .B(u2_u1__abc_47660_n168), .Y(u2_u1_b3_last_row_6__FF_INPUT) );
  AND2X2 AND2X2_3925 ( .A(u2_u1__abc_47660_n137_bF_buf4), .B(u2_u1__abc_47660_n174), .Y(u2_u1__abc_47660_n175) );
  AND2X2 AND2X2_3926 ( .A(u2_u1__abc_47660_n176), .B(u2_u1__abc_47660_n173), .Y(u2_u1_b3_last_row_7__FF_INPUT) );
  AND2X2 AND2X2_3927 ( .A(u2_u1__abc_47660_n137_bF_buf2), .B(u2_u1__abc_47660_n179), .Y(u2_u1__abc_47660_n180) );
  AND2X2 AND2X2_3928 ( .A(u2_u1__abc_47660_n181), .B(u2_u1__abc_47660_n178), .Y(u2_u1_b3_last_row_8__FF_INPUT) );
  AND2X2 AND2X2_3929 ( .A(u2_u1__abc_47660_n137_bF_buf0), .B(u2_u1__abc_47660_n184), .Y(u2_u1__abc_47660_n185) );
  AND2X2 AND2X2_393 ( .A(u0__abc_49347_n1676), .B(u0__abc_49347_n1179_bF_buf3), .Y(u0__abc_49347_n1677_1) );
  AND2X2 AND2X2_3930 ( .A(u2_u1__abc_47660_n186), .B(u2_u1__abc_47660_n183), .Y(u2_u1_b3_last_row_9__FF_INPUT) );
  AND2X2 AND2X2_3931 ( .A(u2_u1__abc_47660_n137_bF_buf3), .B(u2_u1__abc_47660_n189), .Y(u2_u1__abc_47660_n190) );
  AND2X2 AND2X2_3932 ( .A(u2_u1__abc_47660_n191), .B(u2_u1__abc_47660_n188), .Y(u2_u1_b3_last_row_10__FF_INPUT) );
  AND2X2 AND2X2_3933 ( .A(u2_u1__abc_47660_n137_bF_buf1), .B(u2_u1__abc_47660_n194), .Y(u2_u1__abc_47660_n195) );
  AND2X2 AND2X2_3934 ( .A(u2_u1__abc_47660_n196), .B(u2_u1__abc_47660_n193), .Y(u2_u1_b3_last_row_11__FF_INPUT) );
  AND2X2 AND2X2_3935 ( .A(u2_u1__abc_47660_n137_bF_buf4), .B(u2_u1__abc_47660_n199), .Y(u2_u1__abc_47660_n200) );
  AND2X2 AND2X2_3936 ( .A(u2_u1__abc_47660_n201), .B(u2_u1__abc_47660_n198), .Y(u2_u1_b3_last_row_12__FF_INPUT) );
  AND2X2 AND2X2_3937 ( .A(u2_u1__abc_47660_n203), .B(bank_adr_1_bF_buf1), .Y(u2_u1__abc_47660_n204) );
  AND2X2 AND2X2_3938 ( .A(u2_u1__abc_47660_n204), .B(u2_bank_set_1), .Y(u2_u1__abc_47660_n205) );
  AND2X2 AND2X2_3939 ( .A(u2_u1__abc_47660_n208), .B(u2_u1__abc_47660_n206), .Y(u2_u1_b2_last_row_0__FF_INPUT) );
  AND2X2 AND2X2_394 ( .A(spec_req_cs_2_bF_buf0), .B(u0_tms2_20_), .Y(u0__abc_49347_n1678_1) );
  AND2X2 AND2X2_3940 ( .A(u2_u1__abc_47660_n211), .B(u2_u1__abc_47660_n210), .Y(u2_u1_b2_last_row_1__FF_INPUT) );
  AND2X2 AND2X2_3941 ( .A(u2_u1__abc_47660_n214), .B(u2_u1__abc_47660_n213), .Y(u2_u1_b2_last_row_2__FF_INPUT) );
  AND2X2 AND2X2_3942 ( .A(u2_u1__abc_47660_n217), .B(u2_u1__abc_47660_n216), .Y(u2_u1_b2_last_row_3__FF_INPUT) );
  AND2X2 AND2X2_3943 ( .A(u2_u1__abc_47660_n220), .B(u2_u1__abc_47660_n219), .Y(u2_u1_b2_last_row_4__FF_INPUT) );
  AND2X2 AND2X2_3944 ( .A(u2_u1__abc_47660_n223), .B(u2_u1__abc_47660_n222), .Y(u2_u1_b2_last_row_5__FF_INPUT) );
  AND2X2 AND2X2_3945 ( .A(u2_u1__abc_47660_n226), .B(u2_u1__abc_47660_n225), .Y(u2_u1_b2_last_row_6__FF_INPUT) );
  AND2X2 AND2X2_3946 ( .A(u2_u1__abc_47660_n229), .B(u2_u1__abc_47660_n228), .Y(u2_u1_b2_last_row_7__FF_INPUT) );
  AND2X2 AND2X2_3947 ( .A(u2_u1__abc_47660_n232), .B(u2_u1__abc_47660_n231), .Y(u2_u1_b2_last_row_8__FF_INPUT) );
  AND2X2 AND2X2_3948 ( .A(u2_u1__abc_47660_n235), .B(u2_u1__abc_47660_n234), .Y(u2_u1_b2_last_row_9__FF_INPUT) );
  AND2X2 AND2X2_3949 ( .A(u2_u1__abc_47660_n238), .B(u2_u1__abc_47660_n237), .Y(u2_u1_b2_last_row_10__FF_INPUT) );
  AND2X2 AND2X2_395 ( .A(u0__abc_49347_n1679), .B(u0__abc_49347_n1178_1_bF_buf3), .Y(u0__abc_49347_n1680) );
  AND2X2 AND2X2_3950 ( .A(u2_u1__abc_47660_n241), .B(u2_u1__abc_47660_n240), .Y(u2_u1_b2_last_row_11__FF_INPUT) );
  AND2X2 AND2X2_3951 ( .A(u2_u1__abc_47660_n244), .B(u2_u1__abc_47660_n243), .Y(u2_u1_b2_last_row_12__FF_INPUT) );
  AND2X2 AND2X2_3952 ( .A(u2_u1__abc_47660_n246), .B(bank_adr_0_bF_buf0), .Y(u2_u1__abc_47660_n247) );
  AND2X2 AND2X2_3953 ( .A(u2_u1__abc_47660_n247), .B(u2_bank_set_1), .Y(u2_u1__abc_47660_n248) );
  AND2X2 AND2X2_3954 ( .A(u2_u1__abc_47660_n251), .B(u2_u1__abc_47660_n249), .Y(u2_u1_b1_last_row_0__FF_INPUT) );
  AND2X2 AND2X2_3955 ( .A(u2_u1__abc_47660_n254), .B(u2_u1__abc_47660_n253), .Y(u2_u1_b1_last_row_1__FF_INPUT) );
  AND2X2 AND2X2_3956 ( .A(u2_u1__abc_47660_n257), .B(u2_u1__abc_47660_n256), .Y(u2_u1_b1_last_row_2__FF_INPUT) );
  AND2X2 AND2X2_3957 ( .A(u2_u1__abc_47660_n260), .B(u2_u1__abc_47660_n259), .Y(u2_u1_b1_last_row_3__FF_INPUT) );
  AND2X2 AND2X2_3958 ( .A(u2_u1__abc_47660_n263), .B(u2_u1__abc_47660_n262), .Y(u2_u1_b1_last_row_4__FF_INPUT) );
  AND2X2 AND2X2_3959 ( .A(u2_u1__abc_47660_n266), .B(u2_u1__abc_47660_n265), .Y(u2_u1_b1_last_row_5__FF_INPUT) );
  AND2X2 AND2X2_396 ( .A(spec_req_cs_1_bF_buf0), .B(u0_tms1_20_), .Y(u0__abc_49347_n1681) );
  AND2X2 AND2X2_3960 ( .A(u2_u1__abc_47660_n269), .B(u2_u1__abc_47660_n268), .Y(u2_u1_b1_last_row_6__FF_INPUT) );
  AND2X2 AND2X2_3961 ( .A(u2_u1__abc_47660_n272), .B(u2_u1__abc_47660_n271), .Y(u2_u1_b1_last_row_7__FF_INPUT) );
  AND2X2 AND2X2_3962 ( .A(u2_u1__abc_47660_n275_1), .B(u2_u1__abc_47660_n274), .Y(u2_u1_b1_last_row_8__FF_INPUT) );
  AND2X2 AND2X2_3963 ( .A(u2_u1__abc_47660_n278_1), .B(u2_u1__abc_47660_n277), .Y(u2_u1_b1_last_row_9__FF_INPUT) );
  AND2X2 AND2X2_3964 ( .A(u2_u1__abc_47660_n281), .B(u2_u1__abc_47660_n280), .Y(u2_u1_b1_last_row_10__FF_INPUT) );
  AND2X2 AND2X2_3965 ( .A(u2_u1__abc_47660_n284), .B(u2_u1__abc_47660_n283_1), .Y(u2_u1_b1_last_row_11__FF_INPUT) );
  AND2X2 AND2X2_3966 ( .A(u2_u1__abc_47660_n287_1), .B(u2_u1__abc_47660_n286_1), .Y(u2_u1_b1_last_row_12__FF_INPUT) );
  AND2X2 AND2X2_3967 ( .A(u2_u1__abc_47660_n203), .B(u2_u1__abc_47660_n246), .Y(u2_u1__abc_47660_n289) );
  AND2X2 AND2X2_3968 ( .A(u2_u1__abc_47660_n289), .B(u2_bank_set_1), .Y(u2_u1__abc_47660_n290_1) );
  AND2X2 AND2X2_3969 ( .A(u2_u1__abc_47660_n293), .B(u2_u1__abc_47660_n291), .Y(u2_u1_b0_last_row_0__FF_INPUT) );
  AND2X2 AND2X2_397 ( .A(u0__abc_49347_n1175_bF_buf6), .B(u0__abc_49347_n1684), .Y(u0__abc_49347_n1685) );
  AND2X2 AND2X2_3970 ( .A(u2_u1__abc_47660_n296_1), .B(u2_u1__abc_47660_n295), .Y(u2_u1_b0_last_row_1__FF_INPUT) );
  AND2X2 AND2X2_3971 ( .A(u2_u1__abc_47660_n299), .B(u2_u1__abc_47660_n298), .Y(u2_u1_b0_last_row_2__FF_INPUT) );
  AND2X2 AND2X2_3972 ( .A(u2_u1__abc_47660_n302), .B(u2_u1__abc_47660_n301), .Y(u2_u1_b0_last_row_3__FF_INPUT) );
  AND2X2 AND2X2_3973 ( .A(u2_u1__abc_47660_n305_1), .B(u2_u1__abc_47660_n304_1), .Y(u2_u1_b0_last_row_4__FF_INPUT) );
  AND2X2 AND2X2_3974 ( .A(u2_u1__abc_47660_n308), .B(u2_u1__abc_47660_n307), .Y(u2_u1_b0_last_row_5__FF_INPUT) );
  AND2X2 AND2X2_3975 ( .A(u2_u1__abc_47660_n311), .B(u2_u1__abc_47660_n310), .Y(u2_u1_b0_last_row_6__FF_INPUT) );
  AND2X2 AND2X2_3976 ( .A(u2_u1__abc_47660_n314), .B(u2_u1__abc_47660_n313), .Y(u2_u1_b0_last_row_7__FF_INPUT) );
  AND2X2 AND2X2_3977 ( .A(u2_u1__abc_47660_n317), .B(u2_u1__abc_47660_n316), .Y(u2_u1_b0_last_row_8__FF_INPUT) );
  AND2X2 AND2X2_3978 ( .A(u2_u1__abc_47660_n320), .B(u2_u1__abc_47660_n319), .Y(u2_u1_b0_last_row_9__FF_INPUT) );
  AND2X2 AND2X2_3979 ( .A(u2_u1__abc_47660_n323), .B(u2_u1__abc_47660_n322), .Y(u2_u1_b0_last_row_10__FF_INPUT) );
  AND2X2 AND2X2_398 ( .A(u0__abc_49347_n1683), .B(u0__abc_49347_n1685), .Y(u0__abc_49347_n1686_1) );
  AND2X2 AND2X2_3980 ( .A(u2_u1__abc_47660_n326), .B(u2_u1__abc_47660_n325), .Y(u2_u1_b0_last_row_11__FF_INPUT) );
  AND2X2 AND2X2_3981 ( .A(u2_u1__abc_47660_n329), .B(u2_u1__abc_47660_n328), .Y(u2_u1_b0_last_row_12__FF_INPUT) );
  AND2X2 AND2X2_3982 ( .A(u2_u1__abc_47660_n334), .B(u2_u1__abc_47660_n335), .Y(u2_u1__abc_47660_n336) );
  AND2X2 AND2X2_3983 ( .A(u2_u1__abc_47660_n336), .B(u2_u1__abc_47660_n332), .Y(u2_u1__abc_47660_n337) );
  AND2X2 AND2X2_3984 ( .A(u2_u1__abc_47660_n338), .B(u2_u1__abc_47660_n340), .Y(u2_u1__abc_47660_n341) );
  AND2X2 AND2X2_3985 ( .A(u2_u1__abc_47660_n342), .B(u2_u1__abc_47660_n344), .Y(u2_u1__abc_47660_n345) );
  AND2X2 AND2X2_3986 ( .A(u2_u1__abc_47660_n341), .B(u2_u1__abc_47660_n345), .Y(u2_u1__abc_47660_n346) );
  AND2X2 AND2X2_3987 ( .A(u2_u1__abc_47660_n346), .B(u2_u1__abc_47660_n337), .Y(u2_u1__abc_47660_n347) );
  AND2X2 AND2X2_3988 ( .A(u2_u1__abc_47660_n348), .B(u2_u1__abc_47660_n289), .Y(u2_u1__abc_47660_n349) );
  AND2X2 AND2X2_3989 ( .A(u2_u1__abc_47660_n350), .B(u2_u1__abc_47660_n352), .Y(u2_u1__abc_47660_n353) );
  AND2X2 AND2X2_399 ( .A(u0__abc_49347_n1176_1_bF_buf6), .B(sp_tms_21_), .Y(u0__abc_49347_n1688) );
  AND2X2 AND2X2_3990 ( .A(u2_u1__abc_47660_n353), .B(u2_u1__abc_47660_n349), .Y(u2_u1__abc_47660_n354) );
  AND2X2 AND2X2_3991 ( .A(u2_u1__abc_47660_n356), .B(u2_u1__abc_47660_n357), .Y(u2_u1__abc_47660_n358) );
  AND2X2 AND2X2_3992 ( .A(u2_u1__abc_47660_n359), .B(u2_u1__abc_47660_n361), .Y(u2_u1__abc_47660_n362) );
  AND2X2 AND2X2_3993 ( .A(u2_u1__abc_47660_n358), .B(u2_u1__abc_47660_n362), .Y(u2_u1__abc_47660_n363) );
  AND2X2 AND2X2_3994 ( .A(u2_u1__abc_47660_n363), .B(u2_u1__abc_47660_n354), .Y(u2_u1__abc_47660_n364) );
  AND2X2 AND2X2_3995 ( .A(u2_u1__abc_47660_n347), .B(u2_u1__abc_47660_n364), .Y(u2_u1__abc_47660_n365) );
  AND2X2 AND2X2_3996 ( .A(u2_u1__abc_47660_n367), .B(u2_u1__abc_47660_n368), .Y(u2_u1__abc_47660_n369) );
  AND2X2 AND2X2_3997 ( .A(row_adr_8_bF_buf6), .B(u2_u1_b0_last_row_8_), .Y(u2_u1__abc_47660_n370) );
  AND2X2 AND2X2_3998 ( .A(u2_u1__abc_47660_n179), .B(u2_u1__abc_47660_n371), .Y(u2_u1__abc_47660_n372) );
  AND2X2 AND2X2_3999 ( .A(u2_u1__abc_47660_n369), .B(u2_u1__abc_47660_n373), .Y(u2_u1__abc_47660_n374) );
  AND2X2 AND2X2_4 ( .A(_abc_55805_n248), .B(_abc_55805_n249), .Y(_abc_55805_n250) );
  AND2X2 AND2X2_40 ( .A(_abc_55805_n356), .B(_abc_55805_n357), .Y(tms_s_22_) );
  AND2X2 AND2X2_400 ( .A(spec_req_cs_5_bF_buf5), .B(u0_tms5_21_), .Y(u0__abc_49347_n1689) );
  AND2X2 AND2X2_4000 ( .A(u2_u1__abc_47660_n375), .B(u2_u1__abc_47660_n377), .Y(u2_u1__abc_47660_n378) );
  AND2X2 AND2X2_4001 ( .A(u2_u1__abc_47660_n380), .B(u2_u1__abc_47660_n381), .Y(u2_u1__abc_47660_n382) );
  AND2X2 AND2X2_4002 ( .A(u2_u1__abc_47660_n378), .B(u2_u1__abc_47660_n382), .Y(u2_u1__abc_47660_n383) );
  AND2X2 AND2X2_4003 ( .A(u2_u1__abc_47660_n385), .B(u2_u1__abc_47660_n386), .Y(u2_u1__abc_47660_n387) );
  AND2X2 AND2X2_4004 ( .A(row_adr_6_bF_buf6), .B(u2_u1_b0_last_row_6_), .Y(u2_u1__abc_47660_n388) );
  AND2X2 AND2X2_4005 ( .A(u2_u1__abc_47660_n169), .B(u2_u1__abc_47660_n389), .Y(u2_u1__abc_47660_n390) );
  AND2X2 AND2X2_4006 ( .A(u2_u1__abc_47660_n387), .B(u2_u1__abc_47660_n391), .Y(u2_u1__abc_47660_n392) );
  AND2X2 AND2X2_4007 ( .A(u2_u1__abc_47660_n383), .B(u2_u1__abc_47660_n392), .Y(u2_u1__abc_47660_n393) );
  AND2X2 AND2X2_4008 ( .A(u2_u1__abc_47660_n393), .B(u2_u1__abc_47660_n374), .Y(u2_u1__abc_47660_n394) );
  AND2X2 AND2X2_4009 ( .A(u2_u1__abc_47660_n365), .B(u2_u1__abc_47660_n394), .Y(u2_u1__abc_47660_n395) );
  AND2X2 AND2X2_401 ( .A(u0__abc_49347_n1691), .B(u0__abc_49347_n1185_bF_buf2), .Y(u0__abc_49347_n1692) );
  AND2X2 AND2X2_4010 ( .A(u2_u1__abc_47660_n399), .B(u2_u1__abc_47660_n400), .Y(u2_u1__abc_47660_n401) );
  AND2X2 AND2X2_4011 ( .A(u2_u1__abc_47660_n401), .B(u2_u1__abc_47660_n397), .Y(u2_u1__abc_47660_n402) );
  AND2X2 AND2X2_4012 ( .A(u2_u1__abc_47660_n403), .B(u2_u1__abc_47660_n405), .Y(u2_u1__abc_47660_n406) );
  AND2X2 AND2X2_4013 ( .A(u2_u1__abc_47660_n407), .B(u2_u1__abc_47660_n409), .Y(u2_u1__abc_47660_n410) );
  AND2X2 AND2X2_4014 ( .A(u2_u1__abc_47660_n406), .B(u2_u1__abc_47660_n410), .Y(u2_u1__abc_47660_n411) );
  AND2X2 AND2X2_4015 ( .A(u2_u1__abc_47660_n411), .B(u2_u1__abc_47660_n402), .Y(u2_u1__abc_47660_n412) );
  AND2X2 AND2X2_4016 ( .A(u2_u1__abc_47660_n413), .B(u2_u1__abc_47660_n204), .Y(u2_u1__abc_47660_n414) );
  AND2X2 AND2X2_4017 ( .A(u2_u1__abc_47660_n415), .B(u2_u1__abc_47660_n417), .Y(u2_u1__abc_47660_n418) );
  AND2X2 AND2X2_4018 ( .A(u2_u1__abc_47660_n418), .B(u2_u1__abc_47660_n414), .Y(u2_u1__abc_47660_n419) );
  AND2X2 AND2X2_4019 ( .A(u2_u1__abc_47660_n421), .B(u2_u1__abc_47660_n422), .Y(u2_u1__abc_47660_n423) );
  AND2X2 AND2X2_402 ( .A(u0__abc_49347_n1692), .B(u0__abc_49347_n1690), .Y(u0__abc_49347_n1693) );
  AND2X2 AND2X2_4020 ( .A(u2_u1__abc_47660_n424), .B(u2_u1__abc_47660_n426), .Y(u2_u1__abc_47660_n427) );
  AND2X2 AND2X2_4021 ( .A(u2_u1__abc_47660_n423), .B(u2_u1__abc_47660_n427), .Y(u2_u1__abc_47660_n428) );
  AND2X2 AND2X2_4022 ( .A(u2_u1__abc_47660_n428), .B(u2_u1__abc_47660_n419), .Y(u2_u1__abc_47660_n429) );
  AND2X2 AND2X2_4023 ( .A(u2_u1__abc_47660_n412), .B(u2_u1__abc_47660_n429), .Y(u2_u1__abc_47660_n430) );
  AND2X2 AND2X2_4024 ( .A(u2_u1__abc_47660_n432), .B(u2_u1__abc_47660_n433), .Y(u2_u1__abc_47660_n434) );
  AND2X2 AND2X2_4025 ( .A(row_adr_8_bF_buf5), .B(u2_u1_b2_last_row_8_), .Y(u2_u1__abc_47660_n435) );
  AND2X2 AND2X2_4026 ( .A(u2_u1__abc_47660_n179), .B(u2_u1__abc_47660_n436), .Y(u2_u1__abc_47660_n437) );
  AND2X2 AND2X2_4027 ( .A(u2_u1__abc_47660_n434), .B(u2_u1__abc_47660_n438), .Y(u2_u1__abc_47660_n439) );
  AND2X2 AND2X2_4028 ( .A(u2_u1__abc_47660_n440), .B(u2_u1__abc_47660_n442), .Y(u2_u1__abc_47660_n443) );
  AND2X2 AND2X2_4029 ( .A(u2_u1__abc_47660_n445), .B(u2_u1__abc_47660_n446), .Y(u2_u1__abc_47660_n447) );
  AND2X2 AND2X2_403 ( .A(u0__abc_49347_n1694), .B(u0__abc_49347_n1181_bF_buf2), .Y(u0__abc_49347_n1695_1) );
  AND2X2 AND2X2_4030 ( .A(u2_u1__abc_47660_n443), .B(u2_u1__abc_47660_n447), .Y(u2_u1__abc_47660_n448) );
  AND2X2 AND2X2_4031 ( .A(u2_u1__abc_47660_n450), .B(u2_u1__abc_47660_n451), .Y(u2_u1__abc_47660_n452) );
  AND2X2 AND2X2_4032 ( .A(row_adr_6_bF_buf5), .B(u2_u1_b2_last_row_6_), .Y(u2_u1__abc_47660_n453) );
  AND2X2 AND2X2_4033 ( .A(u2_u1__abc_47660_n169), .B(u2_u1__abc_47660_n454), .Y(u2_u1__abc_47660_n455) );
  AND2X2 AND2X2_4034 ( .A(u2_u1__abc_47660_n452), .B(u2_u1__abc_47660_n456), .Y(u2_u1__abc_47660_n457) );
  AND2X2 AND2X2_4035 ( .A(u2_u1__abc_47660_n448), .B(u2_u1__abc_47660_n457), .Y(u2_u1__abc_47660_n458) );
  AND2X2 AND2X2_4036 ( .A(u2_u1__abc_47660_n458), .B(u2_u1__abc_47660_n439), .Y(u2_u1__abc_47660_n459) );
  AND2X2 AND2X2_4037 ( .A(u2_u1__abc_47660_n430), .B(u2_u1__abc_47660_n459), .Y(u2_u1__abc_47660_n460) );
  AND2X2 AND2X2_4038 ( .A(u2_u1__abc_47660_n465), .B(u2_u1__abc_47660_n466), .Y(u2_u1__abc_47660_n467) );
  AND2X2 AND2X2_4039 ( .A(u2_u1__abc_47660_n467), .B(u2_u1__abc_47660_n463), .Y(u2_u1__abc_47660_n468) );
  AND2X2 AND2X2_404 ( .A(spec_req_cs_4_bF_buf5), .B(u0_tms4_21_), .Y(u0__abc_49347_n1696_1) );
  AND2X2 AND2X2_4040 ( .A(u2_u1__abc_47660_n469), .B(u2_u1__abc_47660_n471), .Y(u2_u1__abc_47660_n472) );
  AND2X2 AND2X2_4041 ( .A(u2_u1__abc_47660_n473), .B(u2_u1__abc_47660_n475), .Y(u2_u1__abc_47660_n476) );
  AND2X2 AND2X2_4042 ( .A(u2_u1__abc_47660_n472), .B(u2_u1__abc_47660_n476), .Y(u2_u1__abc_47660_n477) );
  AND2X2 AND2X2_4043 ( .A(u2_u1__abc_47660_n477), .B(u2_u1__abc_47660_n468), .Y(u2_u1__abc_47660_n478) );
  AND2X2 AND2X2_4044 ( .A(u2_u1__abc_47660_n479), .B(u2_u1__abc_47660_n247), .Y(u2_u1__abc_47660_n480) );
  AND2X2 AND2X2_4045 ( .A(u2_u1__abc_47660_n481), .B(u2_u1__abc_47660_n483), .Y(u2_u1__abc_47660_n484) );
  AND2X2 AND2X2_4046 ( .A(u2_u1__abc_47660_n484), .B(u2_u1__abc_47660_n480), .Y(u2_u1__abc_47660_n485) );
  AND2X2 AND2X2_4047 ( .A(u2_u1__abc_47660_n487), .B(u2_u1__abc_47660_n488), .Y(u2_u1__abc_47660_n489) );
  AND2X2 AND2X2_4048 ( .A(u2_u1__abc_47660_n490), .B(u2_u1__abc_47660_n492), .Y(u2_u1__abc_47660_n493) );
  AND2X2 AND2X2_4049 ( .A(u2_u1__abc_47660_n489), .B(u2_u1__abc_47660_n493), .Y(u2_u1__abc_47660_n494) );
  AND2X2 AND2X2_405 ( .A(u0__abc_49347_n1697), .B(u0__abc_49347_n1180_1_bF_buf2), .Y(u0__abc_49347_n1698) );
  AND2X2 AND2X2_4050 ( .A(u2_u1__abc_47660_n494), .B(u2_u1__abc_47660_n485), .Y(u2_u1__abc_47660_n495) );
  AND2X2 AND2X2_4051 ( .A(u2_u1__abc_47660_n478), .B(u2_u1__abc_47660_n495), .Y(u2_u1__abc_47660_n496) );
  AND2X2 AND2X2_4052 ( .A(u2_u1__abc_47660_n498), .B(u2_u1__abc_47660_n499), .Y(u2_u1__abc_47660_n500) );
  AND2X2 AND2X2_4053 ( .A(row_adr_8_bF_buf4), .B(u2_u1_b1_last_row_8_), .Y(u2_u1__abc_47660_n501) );
  AND2X2 AND2X2_4054 ( .A(u2_u1__abc_47660_n179), .B(u2_u1__abc_47660_n502), .Y(u2_u1__abc_47660_n503) );
  AND2X2 AND2X2_4055 ( .A(u2_u1__abc_47660_n500), .B(u2_u1__abc_47660_n504), .Y(u2_u1__abc_47660_n505) );
  AND2X2 AND2X2_4056 ( .A(u2_u1__abc_47660_n506), .B(u2_u1__abc_47660_n508), .Y(u2_u1__abc_47660_n509) );
  AND2X2 AND2X2_4057 ( .A(u2_u1__abc_47660_n511), .B(u2_u1__abc_47660_n512), .Y(u2_u1__abc_47660_n513) );
  AND2X2 AND2X2_4058 ( .A(u2_u1__abc_47660_n509), .B(u2_u1__abc_47660_n513), .Y(u2_u1__abc_47660_n514) );
  AND2X2 AND2X2_4059 ( .A(u2_u1__abc_47660_n516), .B(u2_u1__abc_47660_n517), .Y(u2_u1__abc_47660_n518) );
  AND2X2 AND2X2_406 ( .A(spec_req_cs_3_bF_buf5), .B(u0_tms3_21_), .Y(u0__abc_49347_n1699) );
  AND2X2 AND2X2_4060 ( .A(row_adr_6_bF_buf4), .B(u2_u1_b1_last_row_6_), .Y(u2_u1__abc_47660_n519) );
  AND2X2 AND2X2_4061 ( .A(u2_u1__abc_47660_n169), .B(u2_u1__abc_47660_n520), .Y(u2_u1__abc_47660_n521) );
  AND2X2 AND2X2_4062 ( .A(u2_u1__abc_47660_n518), .B(u2_u1__abc_47660_n522), .Y(u2_u1__abc_47660_n523) );
  AND2X2 AND2X2_4063 ( .A(u2_u1__abc_47660_n514), .B(u2_u1__abc_47660_n523), .Y(u2_u1__abc_47660_n524) );
  AND2X2 AND2X2_4064 ( .A(u2_u1__abc_47660_n524), .B(u2_u1__abc_47660_n505), .Y(u2_u1__abc_47660_n525) );
  AND2X2 AND2X2_4065 ( .A(u2_u1__abc_47660_n496), .B(u2_u1__abc_47660_n525), .Y(u2_u1__abc_47660_n526) );
  AND2X2 AND2X2_4066 ( .A(u2_u1__abc_47660_n529), .B(u2_u1__abc_47660_n530), .Y(u2_u1__abc_47660_n531) );
  AND2X2 AND2X2_4067 ( .A(u2_u1__abc_47660_n531), .B(u2_u1__abc_47660_n528), .Y(u2_u1__abc_47660_n532) );
  AND2X2 AND2X2_4068 ( .A(u2_u1__abc_47660_n533), .B(u2_u1__abc_47660_n535), .Y(u2_u1__abc_47660_n536) );
  AND2X2 AND2X2_4069 ( .A(u2_u1__abc_47660_n537), .B(u2_u1__abc_47660_n539), .Y(u2_u1__abc_47660_n540) );
  AND2X2 AND2X2_407 ( .A(u0__abc_49347_n1700), .B(u0__abc_49347_n1179_bF_buf2), .Y(u0__abc_49347_n1701) );
  AND2X2 AND2X2_4070 ( .A(u2_u1__abc_47660_n536), .B(u2_u1__abc_47660_n540), .Y(u2_u1__abc_47660_n541) );
  AND2X2 AND2X2_4071 ( .A(u2_u1__abc_47660_n541), .B(u2_u1__abc_47660_n532), .Y(u2_u1__abc_47660_n542) );
  AND2X2 AND2X2_4072 ( .A(u2_u1__abc_47660_n543), .B(u2_u1__abc_47660_n545), .Y(u2_u1__abc_47660_n546) );
  AND2X2 AND2X2_4073 ( .A(u2_u1__abc_47660_n548), .B(u2_u1__abc_47660_n136), .Y(u2_u1__abc_47660_n549) );
  AND2X2 AND2X2_4074 ( .A(u2_u1__abc_47660_n546), .B(u2_u1__abc_47660_n549), .Y(u2_u1__abc_47660_n550) );
  AND2X2 AND2X2_4075 ( .A(u2_u1__abc_47660_n552), .B(u2_u1__abc_47660_n553), .Y(u2_u1__abc_47660_n554) );
  AND2X2 AND2X2_4076 ( .A(u2_u1__abc_47660_n556), .B(u2_u1__abc_47660_n557), .Y(u2_u1__abc_47660_n558) );
  AND2X2 AND2X2_4077 ( .A(u2_u1__abc_47660_n554), .B(u2_u1__abc_47660_n558), .Y(u2_u1__abc_47660_n559) );
  AND2X2 AND2X2_4078 ( .A(u2_u1__abc_47660_n559), .B(u2_u1__abc_47660_n550), .Y(u2_u1__abc_47660_n560) );
  AND2X2 AND2X2_4079 ( .A(u2_u1__abc_47660_n542), .B(u2_u1__abc_47660_n560), .Y(u2_u1__abc_47660_n561) );
  AND2X2 AND2X2_408 ( .A(spec_req_cs_2_bF_buf5), .B(u0_tms2_21_), .Y(u0__abc_49347_n1702) );
  AND2X2 AND2X2_4080 ( .A(u2_u1__abc_47660_n562), .B(u2_u1__abc_47660_n564), .Y(u2_u1__abc_47660_n565) );
  AND2X2 AND2X2_4081 ( .A(u2_u1__abc_47660_n567), .B(u2_u1__abc_47660_n568), .Y(u2_u1__abc_47660_n569) );
  AND2X2 AND2X2_4082 ( .A(u2_u1__abc_47660_n565), .B(u2_u1__abc_47660_n569), .Y(u2_u1__abc_47660_n570) );
  AND2X2 AND2X2_4083 ( .A(u2_u1__abc_47660_n571), .B(u2_u1__abc_47660_n573), .Y(u2_u1__abc_47660_n574) );
  AND2X2 AND2X2_4084 ( .A(u2_u1__abc_47660_n576), .B(u2_u1__abc_47660_n577), .Y(u2_u1__abc_47660_n578) );
  AND2X2 AND2X2_4085 ( .A(u2_u1__abc_47660_n574), .B(u2_u1__abc_47660_n578), .Y(u2_u1__abc_47660_n579) );
  AND2X2 AND2X2_4086 ( .A(u2_u1__abc_47660_n580), .B(u2_u1__abc_47660_n582), .Y(u2_u1__abc_47660_n583) );
  AND2X2 AND2X2_4087 ( .A(u2_u1__abc_47660_n584), .B(u2_u1__abc_47660_n586), .Y(u2_u1__abc_47660_n587) );
  AND2X2 AND2X2_4088 ( .A(u2_u1__abc_47660_n583), .B(u2_u1__abc_47660_n587), .Y(u2_u1__abc_47660_n588) );
  AND2X2 AND2X2_4089 ( .A(u2_u1__abc_47660_n579), .B(u2_u1__abc_47660_n588), .Y(u2_u1__abc_47660_n589) );
  AND2X2 AND2X2_409 ( .A(u0__abc_49347_n1703), .B(u0__abc_49347_n1178_1_bF_buf2), .Y(u0__abc_49347_n1704_1) );
  AND2X2 AND2X2_4090 ( .A(u2_u1__abc_47660_n589), .B(u2_u1__abc_47660_n570), .Y(u2_u1__abc_47660_n590) );
  AND2X2 AND2X2_4091 ( .A(u2_u1__abc_47660_n561), .B(u2_u1__abc_47660_n590), .Y(u2_u1__abc_47660_n591) );
  AND2X2 AND2X2_4092 ( .A(u2_u1__abc_47660_n289), .B(u2_u1_bank0_open), .Y(u2_u1__abc_47660_n594) );
  AND2X2 AND2X2_4093 ( .A(u2_u1__abc_47660_n204), .B(u2_u1_bank2_open), .Y(u2_u1__abc_47660_n595) );
  AND2X2 AND2X2_4094 ( .A(u2_u1__abc_47660_n136), .B(u2_u1_bank3_open), .Y(u2_u1__abc_47660_n597) );
  AND2X2 AND2X2_4095 ( .A(u2_u1__abc_47660_n247), .B(u2_u1_bank1_open), .Y(u2_u1__abc_47660_n598) );
  AND2X2 AND2X2_4096 ( .A(u2_u1__abc_47660_n136), .B(u2_bank_clr_1), .Y(u2_u1__abc_47660_n604) );
  AND2X2 AND2X2_4097 ( .A(u2_u1__abc_47660_n606), .B(u2_u1_bank3_open), .Y(u2_u1__abc_47660_n607) );
  AND2X2 AND2X2_4098 ( .A(u2_u1__abc_47660_n605), .B(u2_u1__abc_47660_n607), .Y(u2_u1__abc_47660_n608) );
  AND2X2 AND2X2_4099 ( .A(u2_u1__abc_47660_n606), .B(u2_u1_bank2_open), .Y(u2_u1__abc_47660_n613) );
  AND2X2 AND2X2_41 ( .A(_abc_55805_n359), .B(_abc_55805_n360), .Y(tms_s_23_) );
  AND2X2 AND2X2_410 ( .A(spec_req_cs_1_bF_buf5), .B(u0_tms1_21_), .Y(u0__abc_49347_n1705_1) );
  AND2X2 AND2X2_4100 ( .A(u2_u1__abc_47660_n612), .B(u2_u1__abc_47660_n613), .Y(u2_u1__abc_47660_n614) );
  AND2X2 AND2X2_4101 ( .A(u2_u1__abc_47660_n606), .B(u2_u1_bank1_open), .Y(u2_u1__abc_47660_n618) );
  AND2X2 AND2X2_4102 ( .A(u2_u1__abc_47660_n617), .B(u2_u1__abc_47660_n618), .Y(u2_u1__abc_47660_n619) );
  AND2X2 AND2X2_4103 ( .A(u2_u1__abc_47660_n606), .B(u2_u1_bank0_open), .Y(u2_u1__abc_47660_n623) );
  AND2X2 AND2X2_4104 ( .A(u2_u1__abc_47660_n622), .B(u2_u1__abc_47660_n623), .Y(u2_u1__abc_47660_n624) );
  AND2X2 AND2X2_4105 ( .A(bank_adr_0_bF_buf3), .B(bank_adr_1_bF_buf3), .Y(u2_u2__abc_47660_n136) );
  AND2X2 AND2X2_4106 ( .A(u2_u2__abc_47660_n136), .B(u2_bank_set_2), .Y(u2_u2__abc_47660_n137) );
  AND2X2 AND2X2_4107 ( .A(u2_u2__abc_47660_n137_bF_buf3), .B(u2_u2__abc_47660_n139), .Y(u2_u2__abc_47660_n140) );
  AND2X2 AND2X2_4108 ( .A(u2_u2__abc_47660_n141), .B(u2_u2__abc_47660_n138), .Y(u2_u2_b3_last_row_0__FF_INPUT) );
  AND2X2 AND2X2_4109 ( .A(u2_u2__abc_47660_n137_bF_buf1), .B(u2_u2__abc_47660_n144), .Y(u2_u2__abc_47660_n145) );
  AND2X2 AND2X2_411 ( .A(u0__abc_49347_n1175_bF_buf5), .B(u0__abc_49347_n1708), .Y(u0__abc_49347_n1709) );
  AND2X2 AND2X2_4110 ( .A(u2_u2__abc_47660_n146), .B(u2_u2__abc_47660_n143), .Y(u2_u2_b3_last_row_1__FF_INPUT) );
  AND2X2 AND2X2_4111 ( .A(u2_u2__abc_47660_n137_bF_buf4), .B(u2_u2__abc_47660_n149), .Y(u2_u2__abc_47660_n150) );
  AND2X2 AND2X2_4112 ( .A(u2_u2__abc_47660_n151), .B(u2_u2__abc_47660_n148), .Y(u2_u2_b3_last_row_2__FF_INPUT) );
  AND2X2 AND2X2_4113 ( .A(u2_u2__abc_47660_n137_bF_buf2), .B(u2_u2__abc_47660_n154), .Y(u2_u2__abc_47660_n155) );
  AND2X2 AND2X2_4114 ( .A(u2_u2__abc_47660_n156), .B(u2_u2__abc_47660_n153), .Y(u2_u2_b3_last_row_3__FF_INPUT) );
  AND2X2 AND2X2_4115 ( .A(u2_u2__abc_47660_n137_bF_buf0), .B(u2_u2__abc_47660_n159), .Y(u2_u2__abc_47660_n160) );
  AND2X2 AND2X2_4116 ( .A(u2_u2__abc_47660_n161), .B(u2_u2__abc_47660_n158), .Y(u2_u2_b3_last_row_4__FF_INPUT) );
  AND2X2 AND2X2_4117 ( .A(u2_u2__abc_47660_n137_bF_buf3), .B(u2_u2__abc_47660_n164), .Y(u2_u2__abc_47660_n165) );
  AND2X2 AND2X2_4118 ( .A(u2_u2__abc_47660_n166), .B(u2_u2__abc_47660_n163), .Y(u2_u2_b3_last_row_5__FF_INPUT) );
  AND2X2 AND2X2_4119 ( .A(u2_u2__abc_47660_n137_bF_buf1), .B(u2_u2__abc_47660_n169), .Y(u2_u2__abc_47660_n170) );
  AND2X2 AND2X2_412 ( .A(u0__abc_49347_n1707), .B(u0__abc_49347_n1709), .Y(u0__abc_49347_n1710) );
  AND2X2 AND2X2_4120 ( .A(u2_u2__abc_47660_n171), .B(u2_u2__abc_47660_n168), .Y(u2_u2_b3_last_row_6__FF_INPUT) );
  AND2X2 AND2X2_4121 ( .A(u2_u2__abc_47660_n137_bF_buf4), .B(u2_u2__abc_47660_n174), .Y(u2_u2__abc_47660_n175) );
  AND2X2 AND2X2_4122 ( .A(u2_u2__abc_47660_n176), .B(u2_u2__abc_47660_n173), .Y(u2_u2_b3_last_row_7__FF_INPUT) );
  AND2X2 AND2X2_4123 ( .A(u2_u2__abc_47660_n137_bF_buf2), .B(u2_u2__abc_47660_n179), .Y(u2_u2__abc_47660_n180) );
  AND2X2 AND2X2_4124 ( .A(u2_u2__abc_47660_n181), .B(u2_u2__abc_47660_n178), .Y(u2_u2_b3_last_row_8__FF_INPUT) );
  AND2X2 AND2X2_4125 ( .A(u2_u2__abc_47660_n137_bF_buf0), .B(u2_u2__abc_47660_n184), .Y(u2_u2__abc_47660_n185) );
  AND2X2 AND2X2_4126 ( .A(u2_u2__abc_47660_n186), .B(u2_u2__abc_47660_n183), .Y(u2_u2_b3_last_row_9__FF_INPUT) );
  AND2X2 AND2X2_4127 ( .A(u2_u2__abc_47660_n137_bF_buf3), .B(u2_u2__abc_47660_n189), .Y(u2_u2__abc_47660_n190) );
  AND2X2 AND2X2_4128 ( .A(u2_u2__abc_47660_n191), .B(u2_u2__abc_47660_n188), .Y(u2_u2_b3_last_row_10__FF_INPUT) );
  AND2X2 AND2X2_4129 ( .A(u2_u2__abc_47660_n137_bF_buf1), .B(u2_u2__abc_47660_n194), .Y(u2_u2__abc_47660_n195) );
  AND2X2 AND2X2_413 ( .A(u0__abc_49347_n1176_1_bF_buf5), .B(sp_tms_22_), .Y(u0__abc_49347_n1712) );
  AND2X2 AND2X2_4130 ( .A(u2_u2__abc_47660_n196), .B(u2_u2__abc_47660_n193), .Y(u2_u2_b3_last_row_11__FF_INPUT) );
  AND2X2 AND2X2_4131 ( .A(u2_u2__abc_47660_n137_bF_buf4), .B(u2_u2__abc_47660_n199), .Y(u2_u2__abc_47660_n200) );
  AND2X2 AND2X2_4132 ( .A(u2_u2__abc_47660_n201), .B(u2_u2__abc_47660_n198), .Y(u2_u2_b3_last_row_12__FF_INPUT) );
  AND2X2 AND2X2_4133 ( .A(u2_u2__abc_47660_n203), .B(bank_adr_1_bF_buf2), .Y(u2_u2__abc_47660_n204) );
  AND2X2 AND2X2_4134 ( .A(u2_u2__abc_47660_n204), .B(u2_bank_set_2), .Y(u2_u2__abc_47660_n205) );
  AND2X2 AND2X2_4135 ( .A(u2_u2__abc_47660_n208), .B(u2_u2__abc_47660_n206), .Y(u2_u2_b2_last_row_0__FF_INPUT) );
  AND2X2 AND2X2_4136 ( .A(u2_u2__abc_47660_n211), .B(u2_u2__abc_47660_n210), .Y(u2_u2_b2_last_row_1__FF_INPUT) );
  AND2X2 AND2X2_4137 ( .A(u2_u2__abc_47660_n214), .B(u2_u2__abc_47660_n213), .Y(u2_u2_b2_last_row_2__FF_INPUT) );
  AND2X2 AND2X2_4138 ( .A(u2_u2__abc_47660_n217), .B(u2_u2__abc_47660_n216), .Y(u2_u2_b2_last_row_3__FF_INPUT) );
  AND2X2 AND2X2_4139 ( .A(u2_u2__abc_47660_n220), .B(u2_u2__abc_47660_n219), .Y(u2_u2_b2_last_row_4__FF_INPUT) );
  AND2X2 AND2X2_414 ( .A(spec_req_cs_5_bF_buf4), .B(u0_tms5_22_), .Y(u0__abc_49347_n1713_1) );
  AND2X2 AND2X2_4140 ( .A(u2_u2__abc_47660_n223), .B(u2_u2__abc_47660_n222), .Y(u2_u2_b2_last_row_5__FF_INPUT) );
  AND2X2 AND2X2_4141 ( .A(u2_u2__abc_47660_n226), .B(u2_u2__abc_47660_n225), .Y(u2_u2_b2_last_row_6__FF_INPUT) );
  AND2X2 AND2X2_4142 ( .A(u2_u2__abc_47660_n229), .B(u2_u2__abc_47660_n228), .Y(u2_u2_b2_last_row_7__FF_INPUT) );
  AND2X2 AND2X2_4143 ( .A(u2_u2__abc_47660_n232), .B(u2_u2__abc_47660_n231), .Y(u2_u2_b2_last_row_8__FF_INPUT) );
  AND2X2 AND2X2_4144 ( .A(u2_u2__abc_47660_n235), .B(u2_u2__abc_47660_n234), .Y(u2_u2_b2_last_row_9__FF_INPUT) );
  AND2X2 AND2X2_4145 ( .A(u2_u2__abc_47660_n238), .B(u2_u2__abc_47660_n237), .Y(u2_u2_b2_last_row_10__FF_INPUT) );
  AND2X2 AND2X2_4146 ( .A(u2_u2__abc_47660_n241), .B(u2_u2__abc_47660_n240), .Y(u2_u2_b2_last_row_11__FF_INPUT) );
  AND2X2 AND2X2_4147 ( .A(u2_u2__abc_47660_n244), .B(u2_u2__abc_47660_n243), .Y(u2_u2_b2_last_row_12__FF_INPUT) );
  AND2X2 AND2X2_4148 ( .A(u2_u2__abc_47660_n246), .B(bank_adr_0_bF_buf1), .Y(u2_u2__abc_47660_n247) );
  AND2X2 AND2X2_4149 ( .A(u2_u2__abc_47660_n247), .B(u2_bank_set_2), .Y(u2_u2__abc_47660_n248) );
  AND2X2 AND2X2_415 ( .A(u0__abc_49347_n1715), .B(u0__abc_49347_n1185_bF_buf1), .Y(u0__abc_49347_n1716) );
  AND2X2 AND2X2_4150 ( .A(u2_u2__abc_47660_n251), .B(u2_u2__abc_47660_n249), .Y(u2_u2_b1_last_row_0__FF_INPUT) );
  AND2X2 AND2X2_4151 ( .A(u2_u2__abc_47660_n254), .B(u2_u2__abc_47660_n253), .Y(u2_u2_b1_last_row_1__FF_INPUT) );
  AND2X2 AND2X2_4152 ( .A(u2_u2__abc_47660_n257), .B(u2_u2__abc_47660_n256), .Y(u2_u2_b1_last_row_2__FF_INPUT) );
  AND2X2 AND2X2_4153 ( .A(u2_u2__abc_47660_n260), .B(u2_u2__abc_47660_n259), .Y(u2_u2_b1_last_row_3__FF_INPUT) );
  AND2X2 AND2X2_4154 ( .A(u2_u2__abc_47660_n263), .B(u2_u2__abc_47660_n262), .Y(u2_u2_b1_last_row_4__FF_INPUT) );
  AND2X2 AND2X2_4155 ( .A(u2_u2__abc_47660_n266), .B(u2_u2__abc_47660_n265), .Y(u2_u2_b1_last_row_5__FF_INPUT) );
  AND2X2 AND2X2_4156 ( .A(u2_u2__abc_47660_n269), .B(u2_u2__abc_47660_n268), .Y(u2_u2_b1_last_row_6__FF_INPUT) );
  AND2X2 AND2X2_4157 ( .A(u2_u2__abc_47660_n272), .B(u2_u2__abc_47660_n271), .Y(u2_u2_b1_last_row_7__FF_INPUT) );
  AND2X2 AND2X2_4158 ( .A(u2_u2__abc_47660_n275_1), .B(u2_u2__abc_47660_n274), .Y(u2_u2_b1_last_row_8__FF_INPUT) );
  AND2X2 AND2X2_4159 ( .A(u2_u2__abc_47660_n278_1), .B(u2_u2__abc_47660_n277), .Y(u2_u2_b1_last_row_9__FF_INPUT) );
  AND2X2 AND2X2_416 ( .A(u0__abc_49347_n1716), .B(u0__abc_49347_n1714_1), .Y(u0__abc_49347_n1717) );
  AND2X2 AND2X2_4160 ( .A(u2_u2__abc_47660_n281), .B(u2_u2__abc_47660_n280), .Y(u2_u2_b1_last_row_10__FF_INPUT) );
  AND2X2 AND2X2_4161 ( .A(u2_u2__abc_47660_n284), .B(u2_u2__abc_47660_n283_1), .Y(u2_u2_b1_last_row_11__FF_INPUT) );
  AND2X2 AND2X2_4162 ( .A(u2_u2__abc_47660_n287_1), .B(u2_u2__abc_47660_n286_1), .Y(u2_u2_b1_last_row_12__FF_INPUT) );
  AND2X2 AND2X2_4163 ( .A(u2_u2__abc_47660_n203), .B(u2_u2__abc_47660_n246), .Y(u2_u2__abc_47660_n289) );
  AND2X2 AND2X2_4164 ( .A(u2_u2__abc_47660_n289), .B(u2_bank_set_2), .Y(u2_u2__abc_47660_n290_1) );
  AND2X2 AND2X2_4165 ( .A(u2_u2__abc_47660_n293), .B(u2_u2__abc_47660_n291), .Y(u2_u2_b0_last_row_0__FF_INPUT) );
  AND2X2 AND2X2_4166 ( .A(u2_u2__abc_47660_n296_1), .B(u2_u2__abc_47660_n295), .Y(u2_u2_b0_last_row_1__FF_INPUT) );
  AND2X2 AND2X2_4167 ( .A(u2_u2__abc_47660_n299), .B(u2_u2__abc_47660_n298), .Y(u2_u2_b0_last_row_2__FF_INPUT) );
  AND2X2 AND2X2_4168 ( .A(u2_u2__abc_47660_n302), .B(u2_u2__abc_47660_n301), .Y(u2_u2_b0_last_row_3__FF_INPUT) );
  AND2X2 AND2X2_4169 ( .A(u2_u2__abc_47660_n305_1), .B(u2_u2__abc_47660_n304_1), .Y(u2_u2_b0_last_row_4__FF_INPUT) );
  AND2X2 AND2X2_417 ( .A(u0__abc_49347_n1718), .B(u0__abc_49347_n1181_bF_buf1), .Y(u0__abc_49347_n1719) );
  AND2X2 AND2X2_4170 ( .A(u2_u2__abc_47660_n308), .B(u2_u2__abc_47660_n307), .Y(u2_u2_b0_last_row_5__FF_INPUT) );
  AND2X2 AND2X2_4171 ( .A(u2_u2__abc_47660_n311), .B(u2_u2__abc_47660_n310), .Y(u2_u2_b0_last_row_6__FF_INPUT) );
  AND2X2 AND2X2_4172 ( .A(u2_u2__abc_47660_n314), .B(u2_u2__abc_47660_n313), .Y(u2_u2_b0_last_row_7__FF_INPUT) );
  AND2X2 AND2X2_4173 ( .A(u2_u2__abc_47660_n317), .B(u2_u2__abc_47660_n316), .Y(u2_u2_b0_last_row_8__FF_INPUT) );
  AND2X2 AND2X2_4174 ( .A(u2_u2__abc_47660_n320), .B(u2_u2__abc_47660_n319), .Y(u2_u2_b0_last_row_9__FF_INPUT) );
  AND2X2 AND2X2_4175 ( .A(u2_u2__abc_47660_n323), .B(u2_u2__abc_47660_n322), .Y(u2_u2_b0_last_row_10__FF_INPUT) );
  AND2X2 AND2X2_4176 ( .A(u2_u2__abc_47660_n326), .B(u2_u2__abc_47660_n325), .Y(u2_u2_b0_last_row_11__FF_INPUT) );
  AND2X2 AND2X2_4177 ( .A(u2_u2__abc_47660_n329), .B(u2_u2__abc_47660_n328), .Y(u2_u2_b0_last_row_12__FF_INPUT) );
  AND2X2 AND2X2_4178 ( .A(u2_u2__abc_47660_n334), .B(u2_u2__abc_47660_n335), .Y(u2_u2__abc_47660_n336) );
  AND2X2 AND2X2_4179 ( .A(u2_u2__abc_47660_n336), .B(u2_u2__abc_47660_n332), .Y(u2_u2__abc_47660_n337) );
  AND2X2 AND2X2_418 ( .A(spec_req_cs_4_bF_buf4), .B(u0_tms4_22_), .Y(u0__abc_49347_n1720) );
  AND2X2 AND2X2_4180 ( .A(u2_u2__abc_47660_n338), .B(u2_u2__abc_47660_n340), .Y(u2_u2__abc_47660_n341) );
  AND2X2 AND2X2_4181 ( .A(u2_u2__abc_47660_n342), .B(u2_u2__abc_47660_n344), .Y(u2_u2__abc_47660_n345) );
  AND2X2 AND2X2_4182 ( .A(u2_u2__abc_47660_n341), .B(u2_u2__abc_47660_n345), .Y(u2_u2__abc_47660_n346) );
  AND2X2 AND2X2_4183 ( .A(u2_u2__abc_47660_n346), .B(u2_u2__abc_47660_n337), .Y(u2_u2__abc_47660_n347) );
  AND2X2 AND2X2_4184 ( .A(u2_u2__abc_47660_n348), .B(u2_u2__abc_47660_n289), .Y(u2_u2__abc_47660_n349) );
  AND2X2 AND2X2_4185 ( .A(u2_u2__abc_47660_n350), .B(u2_u2__abc_47660_n352), .Y(u2_u2__abc_47660_n353) );
  AND2X2 AND2X2_4186 ( .A(u2_u2__abc_47660_n353), .B(u2_u2__abc_47660_n349), .Y(u2_u2__abc_47660_n354) );
  AND2X2 AND2X2_4187 ( .A(u2_u2__abc_47660_n356), .B(u2_u2__abc_47660_n357), .Y(u2_u2__abc_47660_n358) );
  AND2X2 AND2X2_4188 ( .A(u2_u2__abc_47660_n359), .B(u2_u2__abc_47660_n361), .Y(u2_u2__abc_47660_n362) );
  AND2X2 AND2X2_4189 ( .A(u2_u2__abc_47660_n358), .B(u2_u2__abc_47660_n362), .Y(u2_u2__abc_47660_n363) );
  AND2X2 AND2X2_419 ( .A(u0__abc_49347_n1721), .B(u0__abc_49347_n1180_1_bF_buf1), .Y(u0__abc_49347_n1722_1) );
  AND2X2 AND2X2_4190 ( .A(u2_u2__abc_47660_n363), .B(u2_u2__abc_47660_n354), .Y(u2_u2__abc_47660_n364) );
  AND2X2 AND2X2_4191 ( .A(u2_u2__abc_47660_n347), .B(u2_u2__abc_47660_n364), .Y(u2_u2__abc_47660_n365) );
  AND2X2 AND2X2_4192 ( .A(u2_u2__abc_47660_n367), .B(u2_u2__abc_47660_n368), .Y(u2_u2__abc_47660_n369) );
  AND2X2 AND2X2_4193 ( .A(row_adr_8_bF_buf5), .B(u2_u2_b0_last_row_8_), .Y(u2_u2__abc_47660_n370) );
  AND2X2 AND2X2_4194 ( .A(u2_u2__abc_47660_n179), .B(u2_u2__abc_47660_n371), .Y(u2_u2__abc_47660_n372) );
  AND2X2 AND2X2_4195 ( .A(u2_u2__abc_47660_n369), .B(u2_u2__abc_47660_n373), .Y(u2_u2__abc_47660_n374) );
  AND2X2 AND2X2_4196 ( .A(u2_u2__abc_47660_n375), .B(u2_u2__abc_47660_n377), .Y(u2_u2__abc_47660_n378) );
  AND2X2 AND2X2_4197 ( .A(u2_u2__abc_47660_n380), .B(u2_u2__abc_47660_n381), .Y(u2_u2__abc_47660_n382) );
  AND2X2 AND2X2_4198 ( .A(u2_u2__abc_47660_n378), .B(u2_u2__abc_47660_n382), .Y(u2_u2__abc_47660_n383) );
  AND2X2 AND2X2_4199 ( .A(u2_u2__abc_47660_n385), .B(u2_u2__abc_47660_n386), .Y(u2_u2__abc_47660_n387) );
  AND2X2 AND2X2_42 ( .A(_abc_55805_n362), .B(_abc_55805_n363), .Y(tms_s_24_) );
  AND2X2 AND2X2_420 ( .A(spec_req_cs_3_bF_buf4), .B(u0_tms3_22_), .Y(u0__abc_49347_n1723_1) );
  AND2X2 AND2X2_4200 ( .A(row_adr_6_bF_buf5), .B(u2_u2_b0_last_row_6_), .Y(u2_u2__abc_47660_n388) );
  AND2X2 AND2X2_4201 ( .A(u2_u2__abc_47660_n169), .B(u2_u2__abc_47660_n389), .Y(u2_u2__abc_47660_n390) );
  AND2X2 AND2X2_4202 ( .A(u2_u2__abc_47660_n387), .B(u2_u2__abc_47660_n391), .Y(u2_u2__abc_47660_n392) );
  AND2X2 AND2X2_4203 ( .A(u2_u2__abc_47660_n383), .B(u2_u2__abc_47660_n392), .Y(u2_u2__abc_47660_n393) );
  AND2X2 AND2X2_4204 ( .A(u2_u2__abc_47660_n393), .B(u2_u2__abc_47660_n374), .Y(u2_u2__abc_47660_n394) );
  AND2X2 AND2X2_4205 ( .A(u2_u2__abc_47660_n365), .B(u2_u2__abc_47660_n394), .Y(u2_u2__abc_47660_n395) );
  AND2X2 AND2X2_4206 ( .A(u2_u2__abc_47660_n399), .B(u2_u2__abc_47660_n400), .Y(u2_u2__abc_47660_n401) );
  AND2X2 AND2X2_4207 ( .A(u2_u2__abc_47660_n401), .B(u2_u2__abc_47660_n397), .Y(u2_u2__abc_47660_n402) );
  AND2X2 AND2X2_4208 ( .A(u2_u2__abc_47660_n403), .B(u2_u2__abc_47660_n405), .Y(u2_u2__abc_47660_n406) );
  AND2X2 AND2X2_4209 ( .A(u2_u2__abc_47660_n407), .B(u2_u2__abc_47660_n409), .Y(u2_u2__abc_47660_n410) );
  AND2X2 AND2X2_421 ( .A(u0__abc_49347_n1724), .B(u0__abc_49347_n1179_bF_buf1), .Y(u0__abc_49347_n1725) );
  AND2X2 AND2X2_4210 ( .A(u2_u2__abc_47660_n406), .B(u2_u2__abc_47660_n410), .Y(u2_u2__abc_47660_n411) );
  AND2X2 AND2X2_4211 ( .A(u2_u2__abc_47660_n411), .B(u2_u2__abc_47660_n402), .Y(u2_u2__abc_47660_n412) );
  AND2X2 AND2X2_4212 ( .A(u2_u2__abc_47660_n413), .B(u2_u2__abc_47660_n204), .Y(u2_u2__abc_47660_n414) );
  AND2X2 AND2X2_4213 ( .A(u2_u2__abc_47660_n415), .B(u2_u2__abc_47660_n417), .Y(u2_u2__abc_47660_n418) );
  AND2X2 AND2X2_4214 ( .A(u2_u2__abc_47660_n418), .B(u2_u2__abc_47660_n414), .Y(u2_u2__abc_47660_n419) );
  AND2X2 AND2X2_4215 ( .A(u2_u2__abc_47660_n421), .B(u2_u2__abc_47660_n422), .Y(u2_u2__abc_47660_n423) );
  AND2X2 AND2X2_4216 ( .A(u2_u2__abc_47660_n424), .B(u2_u2__abc_47660_n426), .Y(u2_u2__abc_47660_n427) );
  AND2X2 AND2X2_4217 ( .A(u2_u2__abc_47660_n423), .B(u2_u2__abc_47660_n427), .Y(u2_u2__abc_47660_n428) );
  AND2X2 AND2X2_4218 ( .A(u2_u2__abc_47660_n428), .B(u2_u2__abc_47660_n419), .Y(u2_u2__abc_47660_n429) );
  AND2X2 AND2X2_4219 ( .A(u2_u2__abc_47660_n412), .B(u2_u2__abc_47660_n429), .Y(u2_u2__abc_47660_n430) );
  AND2X2 AND2X2_422 ( .A(spec_req_cs_2_bF_buf4), .B(u0_tms2_22_), .Y(u0__abc_49347_n1726) );
  AND2X2 AND2X2_4220 ( .A(u2_u2__abc_47660_n432), .B(u2_u2__abc_47660_n433), .Y(u2_u2__abc_47660_n434) );
  AND2X2 AND2X2_4221 ( .A(row_adr_8_bF_buf4), .B(u2_u2_b2_last_row_8_), .Y(u2_u2__abc_47660_n435) );
  AND2X2 AND2X2_4222 ( .A(u2_u2__abc_47660_n179), .B(u2_u2__abc_47660_n436), .Y(u2_u2__abc_47660_n437) );
  AND2X2 AND2X2_4223 ( .A(u2_u2__abc_47660_n434), .B(u2_u2__abc_47660_n438), .Y(u2_u2__abc_47660_n439) );
  AND2X2 AND2X2_4224 ( .A(u2_u2__abc_47660_n440), .B(u2_u2__abc_47660_n442), .Y(u2_u2__abc_47660_n443) );
  AND2X2 AND2X2_4225 ( .A(u2_u2__abc_47660_n445), .B(u2_u2__abc_47660_n446), .Y(u2_u2__abc_47660_n447) );
  AND2X2 AND2X2_4226 ( .A(u2_u2__abc_47660_n443), .B(u2_u2__abc_47660_n447), .Y(u2_u2__abc_47660_n448) );
  AND2X2 AND2X2_4227 ( .A(u2_u2__abc_47660_n450), .B(u2_u2__abc_47660_n451), .Y(u2_u2__abc_47660_n452) );
  AND2X2 AND2X2_4228 ( .A(row_adr_6_bF_buf4), .B(u2_u2_b2_last_row_6_), .Y(u2_u2__abc_47660_n453) );
  AND2X2 AND2X2_4229 ( .A(u2_u2__abc_47660_n169), .B(u2_u2__abc_47660_n454), .Y(u2_u2__abc_47660_n455) );
  AND2X2 AND2X2_423 ( .A(u0__abc_49347_n1727), .B(u0__abc_49347_n1178_1_bF_buf1), .Y(u0__abc_49347_n1728) );
  AND2X2 AND2X2_4230 ( .A(u2_u2__abc_47660_n452), .B(u2_u2__abc_47660_n456), .Y(u2_u2__abc_47660_n457) );
  AND2X2 AND2X2_4231 ( .A(u2_u2__abc_47660_n448), .B(u2_u2__abc_47660_n457), .Y(u2_u2__abc_47660_n458) );
  AND2X2 AND2X2_4232 ( .A(u2_u2__abc_47660_n458), .B(u2_u2__abc_47660_n439), .Y(u2_u2__abc_47660_n459) );
  AND2X2 AND2X2_4233 ( .A(u2_u2__abc_47660_n430), .B(u2_u2__abc_47660_n459), .Y(u2_u2__abc_47660_n460) );
  AND2X2 AND2X2_4234 ( .A(u2_u2__abc_47660_n465), .B(u2_u2__abc_47660_n466), .Y(u2_u2__abc_47660_n467) );
  AND2X2 AND2X2_4235 ( .A(u2_u2__abc_47660_n467), .B(u2_u2__abc_47660_n463), .Y(u2_u2__abc_47660_n468) );
  AND2X2 AND2X2_4236 ( .A(u2_u2__abc_47660_n469), .B(u2_u2__abc_47660_n471), .Y(u2_u2__abc_47660_n472) );
  AND2X2 AND2X2_4237 ( .A(u2_u2__abc_47660_n473), .B(u2_u2__abc_47660_n475), .Y(u2_u2__abc_47660_n476) );
  AND2X2 AND2X2_4238 ( .A(u2_u2__abc_47660_n472), .B(u2_u2__abc_47660_n476), .Y(u2_u2__abc_47660_n477) );
  AND2X2 AND2X2_4239 ( .A(u2_u2__abc_47660_n477), .B(u2_u2__abc_47660_n468), .Y(u2_u2__abc_47660_n478) );
  AND2X2 AND2X2_424 ( .A(spec_req_cs_1_bF_buf4), .B(u0_tms1_22_), .Y(u0__abc_49347_n1729) );
  AND2X2 AND2X2_4240 ( .A(u2_u2__abc_47660_n479), .B(u2_u2__abc_47660_n247), .Y(u2_u2__abc_47660_n480) );
  AND2X2 AND2X2_4241 ( .A(u2_u2__abc_47660_n481), .B(u2_u2__abc_47660_n483), .Y(u2_u2__abc_47660_n484) );
  AND2X2 AND2X2_4242 ( .A(u2_u2__abc_47660_n484), .B(u2_u2__abc_47660_n480), .Y(u2_u2__abc_47660_n485) );
  AND2X2 AND2X2_4243 ( .A(u2_u2__abc_47660_n487), .B(u2_u2__abc_47660_n488), .Y(u2_u2__abc_47660_n489) );
  AND2X2 AND2X2_4244 ( .A(u2_u2__abc_47660_n490), .B(u2_u2__abc_47660_n492), .Y(u2_u2__abc_47660_n493) );
  AND2X2 AND2X2_4245 ( .A(u2_u2__abc_47660_n489), .B(u2_u2__abc_47660_n493), .Y(u2_u2__abc_47660_n494) );
  AND2X2 AND2X2_4246 ( .A(u2_u2__abc_47660_n494), .B(u2_u2__abc_47660_n485), .Y(u2_u2__abc_47660_n495) );
  AND2X2 AND2X2_4247 ( .A(u2_u2__abc_47660_n478), .B(u2_u2__abc_47660_n495), .Y(u2_u2__abc_47660_n496) );
  AND2X2 AND2X2_4248 ( .A(u2_u2__abc_47660_n498), .B(u2_u2__abc_47660_n499), .Y(u2_u2__abc_47660_n500) );
  AND2X2 AND2X2_4249 ( .A(row_adr_8_bF_buf3), .B(u2_u2_b1_last_row_8_), .Y(u2_u2__abc_47660_n501) );
  AND2X2 AND2X2_425 ( .A(u0__abc_49347_n1175_bF_buf4), .B(u0__abc_49347_n1732_1), .Y(u0__abc_49347_n1733) );
  AND2X2 AND2X2_4250 ( .A(u2_u2__abc_47660_n179), .B(u2_u2__abc_47660_n502), .Y(u2_u2__abc_47660_n503) );
  AND2X2 AND2X2_4251 ( .A(u2_u2__abc_47660_n500), .B(u2_u2__abc_47660_n504), .Y(u2_u2__abc_47660_n505) );
  AND2X2 AND2X2_4252 ( .A(u2_u2__abc_47660_n506), .B(u2_u2__abc_47660_n508), .Y(u2_u2__abc_47660_n509) );
  AND2X2 AND2X2_4253 ( .A(u2_u2__abc_47660_n511), .B(u2_u2__abc_47660_n512), .Y(u2_u2__abc_47660_n513) );
  AND2X2 AND2X2_4254 ( .A(u2_u2__abc_47660_n509), .B(u2_u2__abc_47660_n513), .Y(u2_u2__abc_47660_n514) );
  AND2X2 AND2X2_4255 ( .A(u2_u2__abc_47660_n516), .B(u2_u2__abc_47660_n517), .Y(u2_u2__abc_47660_n518) );
  AND2X2 AND2X2_4256 ( .A(row_adr_6_bF_buf3), .B(u2_u2_b1_last_row_6_), .Y(u2_u2__abc_47660_n519) );
  AND2X2 AND2X2_4257 ( .A(u2_u2__abc_47660_n169), .B(u2_u2__abc_47660_n520), .Y(u2_u2__abc_47660_n521) );
  AND2X2 AND2X2_4258 ( .A(u2_u2__abc_47660_n518), .B(u2_u2__abc_47660_n522), .Y(u2_u2__abc_47660_n523) );
  AND2X2 AND2X2_4259 ( .A(u2_u2__abc_47660_n514), .B(u2_u2__abc_47660_n523), .Y(u2_u2__abc_47660_n524) );
  AND2X2 AND2X2_426 ( .A(u0__abc_49347_n1731_1), .B(u0__abc_49347_n1733), .Y(u0__abc_49347_n1734) );
  AND2X2 AND2X2_4260 ( .A(u2_u2__abc_47660_n524), .B(u2_u2__abc_47660_n505), .Y(u2_u2__abc_47660_n525) );
  AND2X2 AND2X2_4261 ( .A(u2_u2__abc_47660_n496), .B(u2_u2__abc_47660_n525), .Y(u2_u2__abc_47660_n526) );
  AND2X2 AND2X2_4262 ( .A(u2_u2__abc_47660_n529), .B(u2_u2__abc_47660_n530), .Y(u2_u2__abc_47660_n531) );
  AND2X2 AND2X2_4263 ( .A(u2_u2__abc_47660_n531), .B(u2_u2__abc_47660_n528), .Y(u2_u2__abc_47660_n532) );
  AND2X2 AND2X2_4264 ( .A(u2_u2__abc_47660_n533), .B(u2_u2__abc_47660_n535), .Y(u2_u2__abc_47660_n536) );
  AND2X2 AND2X2_4265 ( .A(u2_u2__abc_47660_n537), .B(u2_u2__abc_47660_n539), .Y(u2_u2__abc_47660_n540) );
  AND2X2 AND2X2_4266 ( .A(u2_u2__abc_47660_n536), .B(u2_u2__abc_47660_n540), .Y(u2_u2__abc_47660_n541) );
  AND2X2 AND2X2_4267 ( .A(u2_u2__abc_47660_n541), .B(u2_u2__abc_47660_n532), .Y(u2_u2__abc_47660_n542) );
  AND2X2 AND2X2_4268 ( .A(u2_u2__abc_47660_n543), .B(u2_u2__abc_47660_n545), .Y(u2_u2__abc_47660_n546) );
  AND2X2 AND2X2_4269 ( .A(u2_u2__abc_47660_n548), .B(u2_u2__abc_47660_n136), .Y(u2_u2__abc_47660_n549) );
  AND2X2 AND2X2_427 ( .A(u0__abc_49347_n1176_1_bF_buf4), .B(sp_tms_23_), .Y(u0__abc_49347_n1736) );
  AND2X2 AND2X2_4270 ( .A(u2_u2__abc_47660_n546), .B(u2_u2__abc_47660_n549), .Y(u2_u2__abc_47660_n550) );
  AND2X2 AND2X2_4271 ( .A(u2_u2__abc_47660_n552), .B(u2_u2__abc_47660_n553), .Y(u2_u2__abc_47660_n554) );
  AND2X2 AND2X2_4272 ( .A(u2_u2__abc_47660_n556), .B(u2_u2__abc_47660_n557), .Y(u2_u2__abc_47660_n558) );
  AND2X2 AND2X2_4273 ( .A(u2_u2__abc_47660_n554), .B(u2_u2__abc_47660_n558), .Y(u2_u2__abc_47660_n559) );
  AND2X2 AND2X2_4274 ( .A(u2_u2__abc_47660_n559), .B(u2_u2__abc_47660_n550), .Y(u2_u2__abc_47660_n560) );
  AND2X2 AND2X2_4275 ( .A(u2_u2__abc_47660_n542), .B(u2_u2__abc_47660_n560), .Y(u2_u2__abc_47660_n561) );
  AND2X2 AND2X2_4276 ( .A(u2_u2__abc_47660_n562), .B(u2_u2__abc_47660_n564), .Y(u2_u2__abc_47660_n565) );
  AND2X2 AND2X2_4277 ( .A(u2_u2__abc_47660_n567), .B(u2_u2__abc_47660_n568), .Y(u2_u2__abc_47660_n569) );
  AND2X2 AND2X2_4278 ( .A(u2_u2__abc_47660_n565), .B(u2_u2__abc_47660_n569), .Y(u2_u2__abc_47660_n570) );
  AND2X2 AND2X2_4279 ( .A(u2_u2__abc_47660_n571), .B(u2_u2__abc_47660_n573), .Y(u2_u2__abc_47660_n574) );
  AND2X2 AND2X2_428 ( .A(spec_req_cs_5_bF_buf3), .B(u0_tms5_23_), .Y(u0__abc_49347_n1737) );
  AND2X2 AND2X2_4280 ( .A(u2_u2__abc_47660_n576), .B(u2_u2__abc_47660_n577), .Y(u2_u2__abc_47660_n578) );
  AND2X2 AND2X2_4281 ( .A(u2_u2__abc_47660_n574), .B(u2_u2__abc_47660_n578), .Y(u2_u2__abc_47660_n579) );
  AND2X2 AND2X2_4282 ( .A(u2_u2__abc_47660_n580), .B(u2_u2__abc_47660_n582), .Y(u2_u2__abc_47660_n583) );
  AND2X2 AND2X2_4283 ( .A(u2_u2__abc_47660_n584), .B(u2_u2__abc_47660_n586), .Y(u2_u2__abc_47660_n587) );
  AND2X2 AND2X2_4284 ( .A(u2_u2__abc_47660_n583), .B(u2_u2__abc_47660_n587), .Y(u2_u2__abc_47660_n588) );
  AND2X2 AND2X2_4285 ( .A(u2_u2__abc_47660_n579), .B(u2_u2__abc_47660_n588), .Y(u2_u2__abc_47660_n589) );
  AND2X2 AND2X2_4286 ( .A(u2_u2__abc_47660_n589), .B(u2_u2__abc_47660_n570), .Y(u2_u2__abc_47660_n590) );
  AND2X2 AND2X2_4287 ( .A(u2_u2__abc_47660_n561), .B(u2_u2__abc_47660_n590), .Y(u2_u2__abc_47660_n591) );
  AND2X2 AND2X2_4288 ( .A(u2_u2__abc_47660_n289), .B(u2_u2_bank0_open), .Y(u2_u2__abc_47660_n594) );
  AND2X2 AND2X2_4289 ( .A(u2_u2__abc_47660_n204), .B(u2_u2_bank2_open), .Y(u2_u2__abc_47660_n595) );
  AND2X2 AND2X2_429 ( .A(u0__abc_49347_n1739), .B(u0__abc_49347_n1185_bF_buf0), .Y(u0__abc_49347_n1740_1) );
  AND2X2 AND2X2_4290 ( .A(u2_u2__abc_47660_n136), .B(u2_u2_bank3_open), .Y(u2_u2__abc_47660_n597) );
  AND2X2 AND2X2_4291 ( .A(u2_u2__abc_47660_n247), .B(u2_u2_bank1_open), .Y(u2_u2__abc_47660_n598) );
  AND2X2 AND2X2_4292 ( .A(u2_u2__abc_47660_n136), .B(u2_bank_clr_2), .Y(u2_u2__abc_47660_n604) );
  AND2X2 AND2X2_4293 ( .A(u2_u2__abc_47660_n606), .B(u2_u2_bank3_open), .Y(u2_u2__abc_47660_n607) );
  AND2X2 AND2X2_4294 ( .A(u2_u2__abc_47660_n605), .B(u2_u2__abc_47660_n607), .Y(u2_u2__abc_47660_n608) );
  AND2X2 AND2X2_4295 ( .A(u2_u2__abc_47660_n606), .B(u2_u2_bank2_open), .Y(u2_u2__abc_47660_n613) );
  AND2X2 AND2X2_4296 ( .A(u2_u2__abc_47660_n612), .B(u2_u2__abc_47660_n613), .Y(u2_u2__abc_47660_n614) );
  AND2X2 AND2X2_4297 ( .A(u2_u2__abc_47660_n606), .B(u2_u2_bank1_open), .Y(u2_u2__abc_47660_n618) );
  AND2X2 AND2X2_4298 ( .A(u2_u2__abc_47660_n617), .B(u2_u2__abc_47660_n618), .Y(u2_u2__abc_47660_n619) );
  AND2X2 AND2X2_4299 ( .A(u2_u2__abc_47660_n606), .B(u2_u2_bank0_open), .Y(u2_u2__abc_47660_n623) );
  AND2X2 AND2X2_43 ( .A(_abc_55805_n365), .B(_abc_55805_n366), .Y(tms_s_25_) );
  AND2X2 AND2X2_430 ( .A(u0__abc_49347_n1740_1), .B(u0__abc_49347_n1738), .Y(u0__abc_49347_n1741_1) );
  AND2X2 AND2X2_4300 ( .A(u2_u2__abc_47660_n622), .B(u2_u2__abc_47660_n623), .Y(u2_u2__abc_47660_n624) );
  AND2X2 AND2X2_4301 ( .A(bank_adr_0_bF_buf0), .B(bank_adr_1_bF_buf0), .Y(u2_u3__abc_47660_n136) );
  AND2X2 AND2X2_4302 ( .A(u2_u3__abc_47660_n136), .B(u2_bank_set_3), .Y(u2_u3__abc_47660_n137) );
  AND2X2 AND2X2_4303 ( .A(u2_u3__abc_47660_n137_bF_buf3), .B(u2_u3__abc_47660_n139), .Y(u2_u3__abc_47660_n140) );
  AND2X2 AND2X2_4304 ( .A(u2_u3__abc_47660_n141), .B(u2_u3__abc_47660_n138), .Y(u2_u3_b3_last_row_0__FF_INPUT) );
  AND2X2 AND2X2_4305 ( .A(u2_u3__abc_47660_n137_bF_buf1), .B(u2_u3__abc_47660_n144), .Y(u2_u3__abc_47660_n145) );
  AND2X2 AND2X2_4306 ( .A(u2_u3__abc_47660_n146), .B(u2_u3__abc_47660_n143), .Y(u2_u3_b3_last_row_1__FF_INPUT) );
  AND2X2 AND2X2_4307 ( .A(u2_u3__abc_47660_n137_bF_buf4), .B(u2_u3__abc_47660_n149), .Y(u2_u3__abc_47660_n150) );
  AND2X2 AND2X2_4308 ( .A(u2_u3__abc_47660_n151), .B(u2_u3__abc_47660_n148), .Y(u2_u3_b3_last_row_2__FF_INPUT) );
  AND2X2 AND2X2_4309 ( .A(u2_u3__abc_47660_n137_bF_buf2), .B(u2_u3__abc_47660_n154), .Y(u2_u3__abc_47660_n155) );
  AND2X2 AND2X2_431 ( .A(u0__abc_49347_n1742), .B(u0__abc_49347_n1181_bF_buf0), .Y(u0__abc_49347_n1743) );
  AND2X2 AND2X2_4310 ( .A(u2_u3__abc_47660_n156), .B(u2_u3__abc_47660_n153), .Y(u2_u3_b3_last_row_3__FF_INPUT) );
  AND2X2 AND2X2_4311 ( .A(u2_u3__abc_47660_n137_bF_buf0), .B(u2_u3__abc_47660_n159), .Y(u2_u3__abc_47660_n160) );
  AND2X2 AND2X2_4312 ( .A(u2_u3__abc_47660_n161), .B(u2_u3__abc_47660_n158), .Y(u2_u3_b3_last_row_4__FF_INPUT) );
  AND2X2 AND2X2_4313 ( .A(u2_u3__abc_47660_n137_bF_buf3), .B(u2_u3__abc_47660_n164), .Y(u2_u3__abc_47660_n165) );
  AND2X2 AND2X2_4314 ( .A(u2_u3__abc_47660_n166), .B(u2_u3__abc_47660_n163), .Y(u2_u3_b3_last_row_5__FF_INPUT) );
  AND2X2 AND2X2_4315 ( .A(u2_u3__abc_47660_n137_bF_buf1), .B(u2_u3__abc_47660_n169), .Y(u2_u3__abc_47660_n170) );
  AND2X2 AND2X2_4316 ( .A(u2_u3__abc_47660_n171), .B(u2_u3__abc_47660_n168), .Y(u2_u3_b3_last_row_6__FF_INPUT) );
  AND2X2 AND2X2_4317 ( .A(u2_u3__abc_47660_n137_bF_buf4), .B(u2_u3__abc_47660_n174), .Y(u2_u3__abc_47660_n175) );
  AND2X2 AND2X2_4318 ( .A(u2_u3__abc_47660_n176), .B(u2_u3__abc_47660_n173), .Y(u2_u3_b3_last_row_7__FF_INPUT) );
  AND2X2 AND2X2_4319 ( .A(u2_u3__abc_47660_n137_bF_buf2), .B(u2_u3__abc_47660_n179), .Y(u2_u3__abc_47660_n180) );
  AND2X2 AND2X2_432 ( .A(spec_req_cs_4_bF_buf3), .B(u0_tms4_23_), .Y(u0__abc_49347_n1744) );
  AND2X2 AND2X2_4320 ( .A(u2_u3__abc_47660_n181), .B(u2_u3__abc_47660_n178), .Y(u2_u3_b3_last_row_8__FF_INPUT) );
  AND2X2 AND2X2_4321 ( .A(u2_u3__abc_47660_n137_bF_buf0), .B(u2_u3__abc_47660_n184), .Y(u2_u3__abc_47660_n185) );
  AND2X2 AND2X2_4322 ( .A(u2_u3__abc_47660_n186), .B(u2_u3__abc_47660_n183), .Y(u2_u3_b3_last_row_9__FF_INPUT) );
  AND2X2 AND2X2_4323 ( .A(u2_u3__abc_47660_n137_bF_buf3), .B(u2_u3__abc_47660_n189), .Y(u2_u3__abc_47660_n190) );
  AND2X2 AND2X2_4324 ( .A(u2_u3__abc_47660_n191), .B(u2_u3__abc_47660_n188), .Y(u2_u3_b3_last_row_10__FF_INPUT) );
  AND2X2 AND2X2_4325 ( .A(u2_u3__abc_47660_n137_bF_buf1), .B(u2_u3__abc_47660_n194), .Y(u2_u3__abc_47660_n195) );
  AND2X2 AND2X2_4326 ( .A(u2_u3__abc_47660_n196), .B(u2_u3__abc_47660_n193), .Y(u2_u3_b3_last_row_11__FF_INPUT) );
  AND2X2 AND2X2_4327 ( .A(u2_u3__abc_47660_n137_bF_buf4), .B(u2_u3__abc_47660_n199), .Y(u2_u3__abc_47660_n200) );
  AND2X2 AND2X2_4328 ( .A(u2_u3__abc_47660_n201), .B(u2_u3__abc_47660_n198), .Y(u2_u3_b3_last_row_12__FF_INPUT) );
  AND2X2 AND2X2_4329 ( .A(u2_u3__abc_47660_n203), .B(bank_adr_1_bF_buf3), .Y(u2_u3__abc_47660_n204) );
  AND2X2 AND2X2_433 ( .A(u0__abc_49347_n1745), .B(u0__abc_49347_n1180_1_bF_buf0), .Y(u0__abc_49347_n1746) );
  AND2X2 AND2X2_4330 ( .A(u2_u3__abc_47660_n204), .B(u2_bank_set_3), .Y(u2_u3__abc_47660_n205) );
  AND2X2 AND2X2_4331 ( .A(u2_u3__abc_47660_n208), .B(u2_u3__abc_47660_n206), .Y(u2_u3_b2_last_row_0__FF_INPUT) );
  AND2X2 AND2X2_4332 ( .A(u2_u3__abc_47660_n211), .B(u2_u3__abc_47660_n210), .Y(u2_u3_b2_last_row_1__FF_INPUT) );
  AND2X2 AND2X2_4333 ( .A(u2_u3__abc_47660_n214), .B(u2_u3__abc_47660_n213), .Y(u2_u3_b2_last_row_2__FF_INPUT) );
  AND2X2 AND2X2_4334 ( .A(u2_u3__abc_47660_n217), .B(u2_u3__abc_47660_n216), .Y(u2_u3_b2_last_row_3__FF_INPUT) );
  AND2X2 AND2X2_4335 ( .A(u2_u3__abc_47660_n220), .B(u2_u3__abc_47660_n219), .Y(u2_u3_b2_last_row_4__FF_INPUT) );
  AND2X2 AND2X2_4336 ( .A(u2_u3__abc_47660_n223), .B(u2_u3__abc_47660_n222), .Y(u2_u3_b2_last_row_5__FF_INPUT) );
  AND2X2 AND2X2_4337 ( .A(u2_u3__abc_47660_n226), .B(u2_u3__abc_47660_n225), .Y(u2_u3_b2_last_row_6__FF_INPUT) );
  AND2X2 AND2X2_4338 ( .A(u2_u3__abc_47660_n229), .B(u2_u3__abc_47660_n228), .Y(u2_u3_b2_last_row_7__FF_INPUT) );
  AND2X2 AND2X2_4339 ( .A(u2_u3__abc_47660_n232), .B(u2_u3__abc_47660_n231), .Y(u2_u3_b2_last_row_8__FF_INPUT) );
  AND2X2 AND2X2_434 ( .A(spec_req_cs_3_bF_buf3), .B(u0_tms3_23_), .Y(u0__abc_49347_n1747) );
  AND2X2 AND2X2_4340 ( .A(u2_u3__abc_47660_n235), .B(u2_u3__abc_47660_n234), .Y(u2_u3_b2_last_row_9__FF_INPUT) );
  AND2X2 AND2X2_4341 ( .A(u2_u3__abc_47660_n238), .B(u2_u3__abc_47660_n237), .Y(u2_u3_b2_last_row_10__FF_INPUT) );
  AND2X2 AND2X2_4342 ( .A(u2_u3__abc_47660_n241), .B(u2_u3__abc_47660_n240), .Y(u2_u3_b2_last_row_11__FF_INPUT) );
  AND2X2 AND2X2_4343 ( .A(u2_u3__abc_47660_n244), .B(u2_u3__abc_47660_n243), .Y(u2_u3_b2_last_row_12__FF_INPUT) );
  AND2X2 AND2X2_4344 ( .A(u2_u3__abc_47660_n246), .B(bank_adr_0_bF_buf2), .Y(u2_u3__abc_47660_n247) );
  AND2X2 AND2X2_4345 ( .A(u2_u3__abc_47660_n247), .B(u2_bank_set_3), .Y(u2_u3__abc_47660_n248) );
  AND2X2 AND2X2_4346 ( .A(u2_u3__abc_47660_n251), .B(u2_u3__abc_47660_n249), .Y(u2_u3_b1_last_row_0__FF_INPUT) );
  AND2X2 AND2X2_4347 ( .A(u2_u3__abc_47660_n254), .B(u2_u3__abc_47660_n253), .Y(u2_u3_b1_last_row_1__FF_INPUT) );
  AND2X2 AND2X2_4348 ( .A(u2_u3__abc_47660_n257), .B(u2_u3__abc_47660_n256), .Y(u2_u3_b1_last_row_2__FF_INPUT) );
  AND2X2 AND2X2_4349 ( .A(u2_u3__abc_47660_n260), .B(u2_u3__abc_47660_n259), .Y(u2_u3_b1_last_row_3__FF_INPUT) );
  AND2X2 AND2X2_435 ( .A(u0__abc_49347_n1748), .B(u0__abc_49347_n1179_bF_buf0), .Y(u0__abc_49347_n1749_1) );
  AND2X2 AND2X2_4350 ( .A(u2_u3__abc_47660_n263), .B(u2_u3__abc_47660_n262), .Y(u2_u3_b1_last_row_4__FF_INPUT) );
  AND2X2 AND2X2_4351 ( .A(u2_u3__abc_47660_n266), .B(u2_u3__abc_47660_n265), .Y(u2_u3_b1_last_row_5__FF_INPUT) );
  AND2X2 AND2X2_4352 ( .A(u2_u3__abc_47660_n269), .B(u2_u3__abc_47660_n268), .Y(u2_u3_b1_last_row_6__FF_INPUT) );
  AND2X2 AND2X2_4353 ( .A(u2_u3__abc_47660_n272), .B(u2_u3__abc_47660_n271), .Y(u2_u3_b1_last_row_7__FF_INPUT) );
  AND2X2 AND2X2_4354 ( .A(u2_u3__abc_47660_n275_1), .B(u2_u3__abc_47660_n274), .Y(u2_u3_b1_last_row_8__FF_INPUT) );
  AND2X2 AND2X2_4355 ( .A(u2_u3__abc_47660_n278_1), .B(u2_u3__abc_47660_n277), .Y(u2_u3_b1_last_row_9__FF_INPUT) );
  AND2X2 AND2X2_4356 ( .A(u2_u3__abc_47660_n281), .B(u2_u3__abc_47660_n280), .Y(u2_u3_b1_last_row_10__FF_INPUT) );
  AND2X2 AND2X2_4357 ( .A(u2_u3__abc_47660_n284), .B(u2_u3__abc_47660_n283_1), .Y(u2_u3_b1_last_row_11__FF_INPUT) );
  AND2X2 AND2X2_4358 ( .A(u2_u3__abc_47660_n287_1), .B(u2_u3__abc_47660_n286_1), .Y(u2_u3_b1_last_row_12__FF_INPUT) );
  AND2X2 AND2X2_4359 ( .A(u2_u3__abc_47660_n203), .B(u2_u3__abc_47660_n246), .Y(u2_u3__abc_47660_n289) );
  AND2X2 AND2X2_436 ( .A(spec_req_cs_2_bF_buf3), .B(u0_tms2_23_), .Y(u0__abc_49347_n1750_1) );
  AND2X2 AND2X2_4360 ( .A(u2_u3__abc_47660_n289), .B(u2_bank_set_3), .Y(u2_u3__abc_47660_n290_1) );
  AND2X2 AND2X2_4361 ( .A(u2_u3__abc_47660_n293), .B(u2_u3__abc_47660_n291), .Y(u2_u3_b0_last_row_0__FF_INPUT) );
  AND2X2 AND2X2_4362 ( .A(u2_u3__abc_47660_n296_1), .B(u2_u3__abc_47660_n295), .Y(u2_u3_b0_last_row_1__FF_INPUT) );
  AND2X2 AND2X2_4363 ( .A(u2_u3__abc_47660_n299), .B(u2_u3__abc_47660_n298), .Y(u2_u3_b0_last_row_2__FF_INPUT) );
  AND2X2 AND2X2_4364 ( .A(u2_u3__abc_47660_n302), .B(u2_u3__abc_47660_n301), .Y(u2_u3_b0_last_row_3__FF_INPUT) );
  AND2X2 AND2X2_4365 ( .A(u2_u3__abc_47660_n305_1), .B(u2_u3__abc_47660_n304_1), .Y(u2_u3_b0_last_row_4__FF_INPUT) );
  AND2X2 AND2X2_4366 ( .A(u2_u3__abc_47660_n308), .B(u2_u3__abc_47660_n307), .Y(u2_u3_b0_last_row_5__FF_INPUT) );
  AND2X2 AND2X2_4367 ( .A(u2_u3__abc_47660_n311), .B(u2_u3__abc_47660_n310), .Y(u2_u3_b0_last_row_6__FF_INPUT) );
  AND2X2 AND2X2_4368 ( .A(u2_u3__abc_47660_n314), .B(u2_u3__abc_47660_n313), .Y(u2_u3_b0_last_row_7__FF_INPUT) );
  AND2X2 AND2X2_4369 ( .A(u2_u3__abc_47660_n317), .B(u2_u3__abc_47660_n316), .Y(u2_u3_b0_last_row_8__FF_INPUT) );
  AND2X2 AND2X2_437 ( .A(u0__abc_49347_n1751_1), .B(u0__abc_49347_n1178_1_bF_buf0), .Y(u0__abc_49347_n1752) );
  AND2X2 AND2X2_4370 ( .A(u2_u3__abc_47660_n320), .B(u2_u3__abc_47660_n319), .Y(u2_u3_b0_last_row_9__FF_INPUT) );
  AND2X2 AND2X2_4371 ( .A(u2_u3__abc_47660_n323), .B(u2_u3__abc_47660_n322), .Y(u2_u3_b0_last_row_10__FF_INPUT) );
  AND2X2 AND2X2_4372 ( .A(u2_u3__abc_47660_n326), .B(u2_u3__abc_47660_n325), .Y(u2_u3_b0_last_row_11__FF_INPUT) );
  AND2X2 AND2X2_4373 ( .A(u2_u3__abc_47660_n329), .B(u2_u3__abc_47660_n328), .Y(u2_u3_b0_last_row_12__FF_INPUT) );
  AND2X2 AND2X2_4374 ( .A(u2_u3__abc_47660_n334), .B(u2_u3__abc_47660_n335), .Y(u2_u3__abc_47660_n336) );
  AND2X2 AND2X2_4375 ( .A(u2_u3__abc_47660_n336), .B(u2_u3__abc_47660_n332), .Y(u2_u3__abc_47660_n337) );
  AND2X2 AND2X2_4376 ( .A(u2_u3__abc_47660_n338), .B(u2_u3__abc_47660_n340), .Y(u2_u3__abc_47660_n341) );
  AND2X2 AND2X2_4377 ( .A(u2_u3__abc_47660_n342), .B(u2_u3__abc_47660_n344), .Y(u2_u3__abc_47660_n345) );
  AND2X2 AND2X2_4378 ( .A(u2_u3__abc_47660_n341), .B(u2_u3__abc_47660_n345), .Y(u2_u3__abc_47660_n346) );
  AND2X2 AND2X2_4379 ( .A(u2_u3__abc_47660_n346), .B(u2_u3__abc_47660_n337), .Y(u2_u3__abc_47660_n347) );
  AND2X2 AND2X2_438 ( .A(spec_req_cs_1_bF_buf3), .B(u0_tms1_23_), .Y(u0__abc_49347_n1753) );
  AND2X2 AND2X2_4380 ( .A(u2_u3__abc_47660_n348), .B(u2_u3__abc_47660_n289), .Y(u2_u3__abc_47660_n349) );
  AND2X2 AND2X2_4381 ( .A(u2_u3__abc_47660_n350), .B(u2_u3__abc_47660_n352), .Y(u2_u3__abc_47660_n353) );
  AND2X2 AND2X2_4382 ( .A(u2_u3__abc_47660_n353), .B(u2_u3__abc_47660_n349), .Y(u2_u3__abc_47660_n354) );
  AND2X2 AND2X2_4383 ( .A(u2_u3__abc_47660_n356), .B(u2_u3__abc_47660_n357), .Y(u2_u3__abc_47660_n358) );
  AND2X2 AND2X2_4384 ( .A(u2_u3__abc_47660_n359), .B(u2_u3__abc_47660_n361), .Y(u2_u3__abc_47660_n362) );
  AND2X2 AND2X2_4385 ( .A(u2_u3__abc_47660_n358), .B(u2_u3__abc_47660_n362), .Y(u2_u3__abc_47660_n363) );
  AND2X2 AND2X2_4386 ( .A(u2_u3__abc_47660_n363), .B(u2_u3__abc_47660_n354), .Y(u2_u3__abc_47660_n364) );
  AND2X2 AND2X2_4387 ( .A(u2_u3__abc_47660_n347), .B(u2_u3__abc_47660_n364), .Y(u2_u3__abc_47660_n365) );
  AND2X2 AND2X2_4388 ( .A(u2_u3__abc_47660_n367), .B(u2_u3__abc_47660_n368), .Y(u2_u3__abc_47660_n369) );
  AND2X2 AND2X2_4389 ( .A(row_adr_8_bF_buf4), .B(u2_u3_b0_last_row_8_), .Y(u2_u3__abc_47660_n370) );
  AND2X2 AND2X2_439 ( .A(u0__abc_49347_n1175_bF_buf3), .B(u0__abc_49347_n1756_1), .Y(u0__abc_49347_n1757_1) );
  AND2X2 AND2X2_4390 ( .A(u2_u3__abc_47660_n179), .B(u2_u3__abc_47660_n371), .Y(u2_u3__abc_47660_n372) );
  AND2X2 AND2X2_4391 ( .A(u2_u3__abc_47660_n369), .B(u2_u3__abc_47660_n373), .Y(u2_u3__abc_47660_n374) );
  AND2X2 AND2X2_4392 ( .A(u2_u3__abc_47660_n375), .B(u2_u3__abc_47660_n377), .Y(u2_u3__abc_47660_n378) );
  AND2X2 AND2X2_4393 ( .A(u2_u3__abc_47660_n380), .B(u2_u3__abc_47660_n381), .Y(u2_u3__abc_47660_n382) );
  AND2X2 AND2X2_4394 ( .A(u2_u3__abc_47660_n378), .B(u2_u3__abc_47660_n382), .Y(u2_u3__abc_47660_n383) );
  AND2X2 AND2X2_4395 ( .A(u2_u3__abc_47660_n385), .B(u2_u3__abc_47660_n386), .Y(u2_u3__abc_47660_n387) );
  AND2X2 AND2X2_4396 ( .A(row_adr_6_bF_buf4), .B(u2_u3_b0_last_row_6_), .Y(u2_u3__abc_47660_n388) );
  AND2X2 AND2X2_4397 ( .A(u2_u3__abc_47660_n169), .B(u2_u3__abc_47660_n389), .Y(u2_u3__abc_47660_n390) );
  AND2X2 AND2X2_4398 ( .A(u2_u3__abc_47660_n387), .B(u2_u3__abc_47660_n391), .Y(u2_u3__abc_47660_n392) );
  AND2X2 AND2X2_4399 ( .A(u2_u3__abc_47660_n383), .B(u2_u3__abc_47660_n392), .Y(u2_u3__abc_47660_n393) );
  AND2X2 AND2X2_44 ( .A(_abc_55805_n368), .B(_abc_55805_n369), .Y(tms_s_26_) );
  AND2X2 AND2X2_440 ( .A(u0__abc_49347_n1755), .B(u0__abc_49347_n1757_1), .Y(u0__abc_49347_n1758) );
  AND2X2 AND2X2_4400 ( .A(u2_u3__abc_47660_n393), .B(u2_u3__abc_47660_n374), .Y(u2_u3__abc_47660_n394) );
  AND2X2 AND2X2_4401 ( .A(u2_u3__abc_47660_n365), .B(u2_u3__abc_47660_n394), .Y(u2_u3__abc_47660_n395) );
  AND2X2 AND2X2_4402 ( .A(u2_u3__abc_47660_n399), .B(u2_u3__abc_47660_n400), .Y(u2_u3__abc_47660_n401) );
  AND2X2 AND2X2_4403 ( .A(u2_u3__abc_47660_n401), .B(u2_u3__abc_47660_n397), .Y(u2_u3__abc_47660_n402) );
  AND2X2 AND2X2_4404 ( .A(u2_u3__abc_47660_n403), .B(u2_u3__abc_47660_n405), .Y(u2_u3__abc_47660_n406) );
  AND2X2 AND2X2_4405 ( .A(u2_u3__abc_47660_n407), .B(u2_u3__abc_47660_n409), .Y(u2_u3__abc_47660_n410) );
  AND2X2 AND2X2_4406 ( .A(u2_u3__abc_47660_n406), .B(u2_u3__abc_47660_n410), .Y(u2_u3__abc_47660_n411) );
  AND2X2 AND2X2_4407 ( .A(u2_u3__abc_47660_n411), .B(u2_u3__abc_47660_n402), .Y(u2_u3__abc_47660_n412) );
  AND2X2 AND2X2_4408 ( .A(u2_u3__abc_47660_n413), .B(u2_u3__abc_47660_n204), .Y(u2_u3__abc_47660_n414) );
  AND2X2 AND2X2_4409 ( .A(u2_u3__abc_47660_n415), .B(u2_u3__abc_47660_n417), .Y(u2_u3__abc_47660_n418) );
  AND2X2 AND2X2_441 ( .A(u0__abc_49347_n1176_1_bF_buf3), .B(sp_tms_24_), .Y(u0__abc_49347_n1760_1) );
  AND2X2 AND2X2_4410 ( .A(u2_u3__abc_47660_n418), .B(u2_u3__abc_47660_n414), .Y(u2_u3__abc_47660_n419) );
  AND2X2 AND2X2_4411 ( .A(u2_u3__abc_47660_n421), .B(u2_u3__abc_47660_n422), .Y(u2_u3__abc_47660_n423) );
  AND2X2 AND2X2_4412 ( .A(u2_u3__abc_47660_n424), .B(u2_u3__abc_47660_n426), .Y(u2_u3__abc_47660_n427) );
  AND2X2 AND2X2_4413 ( .A(u2_u3__abc_47660_n423), .B(u2_u3__abc_47660_n427), .Y(u2_u3__abc_47660_n428) );
  AND2X2 AND2X2_4414 ( .A(u2_u3__abc_47660_n428), .B(u2_u3__abc_47660_n419), .Y(u2_u3__abc_47660_n429) );
  AND2X2 AND2X2_4415 ( .A(u2_u3__abc_47660_n412), .B(u2_u3__abc_47660_n429), .Y(u2_u3__abc_47660_n430) );
  AND2X2 AND2X2_4416 ( .A(u2_u3__abc_47660_n432), .B(u2_u3__abc_47660_n433), .Y(u2_u3__abc_47660_n434) );
  AND2X2 AND2X2_4417 ( .A(row_adr_8_bF_buf3), .B(u2_u3_b2_last_row_8_), .Y(u2_u3__abc_47660_n435) );
  AND2X2 AND2X2_4418 ( .A(u2_u3__abc_47660_n179), .B(u2_u3__abc_47660_n436), .Y(u2_u3__abc_47660_n437) );
  AND2X2 AND2X2_4419 ( .A(u2_u3__abc_47660_n434), .B(u2_u3__abc_47660_n438), .Y(u2_u3__abc_47660_n439) );
  AND2X2 AND2X2_442 ( .A(spec_req_cs_5_bF_buf2), .B(u0_tms5_24_), .Y(u0__abc_49347_n1761) );
  AND2X2 AND2X2_4420 ( .A(u2_u3__abc_47660_n440), .B(u2_u3__abc_47660_n442), .Y(u2_u3__abc_47660_n443) );
  AND2X2 AND2X2_4421 ( .A(u2_u3__abc_47660_n445), .B(u2_u3__abc_47660_n446), .Y(u2_u3__abc_47660_n447) );
  AND2X2 AND2X2_4422 ( .A(u2_u3__abc_47660_n443), .B(u2_u3__abc_47660_n447), .Y(u2_u3__abc_47660_n448) );
  AND2X2 AND2X2_4423 ( .A(u2_u3__abc_47660_n450), .B(u2_u3__abc_47660_n451), .Y(u2_u3__abc_47660_n452) );
  AND2X2 AND2X2_4424 ( .A(row_adr_6_bF_buf3), .B(u2_u3_b2_last_row_6_), .Y(u2_u3__abc_47660_n453) );
  AND2X2 AND2X2_4425 ( .A(u2_u3__abc_47660_n169), .B(u2_u3__abc_47660_n454), .Y(u2_u3__abc_47660_n455) );
  AND2X2 AND2X2_4426 ( .A(u2_u3__abc_47660_n452), .B(u2_u3__abc_47660_n456), .Y(u2_u3__abc_47660_n457) );
  AND2X2 AND2X2_4427 ( .A(u2_u3__abc_47660_n448), .B(u2_u3__abc_47660_n457), .Y(u2_u3__abc_47660_n458) );
  AND2X2 AND2X2_4428 ( .A(u2_u3__abc_47660_n458), .B(u2_u3__abc_47660_n439), .Y(u2_u3__abc_47660_n459) );
  AND2X2 AND2X2_4429 ( .A(u2_u3__abc_47660_n430), .B(u2_u3__abc_47660_n459), .Y(u2_u3__abc_47660_n460) );
  AND2X2 AND2X2_443 ( .A(u0__abc_49347_n1763_1), .B(u0__abc_49347_n1185_bF_buf5), .Y(u0__abc_49347_n1764_1) );
  AND2X2 AND2X2_4430 ( .A(u2_u3__abc_47660_n465), .B(u2_u3__abc_47660_n466), .Y(u2_u3__abc_47660_n467) );
  AND2X2 AND2X2_4431 ( .A(u2_u3__abc_47660_n467), .B(u2_u3__abc_47660_n463), .Y(u2_u3__abc_47660_n468) );
  AND2X2 AND2X2_4432 ( .A(u2_u3__abc_47660_n469), .B(u2_u3__abc_47660_n471), .Y(u2_u3__abc_47660_n472) );
  AND2X2 AND2X2_4433 ( .A(u2_u3__abc_47660_n473), .B(u2_u3__abc_47660_n475), .Y(u2_u3__abc_47660_n476) );
  AND2X2 AND2X2_4434 ( .A(u2_u3__abc_47660_n472), .B(u2_u3__abc_47660_n476), .Y(u2_u3__abc_47660_n477) );
  AND2X2 AND2X2_4435 ( .A(u2_u3__abc_47660_n477), .B(u2_u3__abc_47660_n468), .Y(u2_u3__abc_47660_n478) );
  AND2X2 AND2X2_4436 ( .A(u2_u3__abc_47660_n479), .B(u2_u3__abc_47660_n247), .Y(u2_u3__abc_47660_n480) );
  AND2X2 AND2X2_4437 ( .A(u2_u3__abc_47660_n481), .B(u2_u3__abc_47660_n483), .Y(u2_u3__abc_47660_n484) );
  AND2X2 AND2X2_4438 ( .A(u2_u3__abc_47660_n484), .B(u2_u3__abc_47660_n480), .Y(u2_u3__abc_47660_n485) );
  AND2X2 AND2X2_4439 ( .A(u2_u3__abc_47660_n487), .B(u2_u3__abc_47660_n488), .Y(u2_u3__abc_47660_n489) );
  AND2X2 AND2X2_444 ( .A(u0__abc_49347_n1764_1), .B(u0__abc_49347_n1762), .Y(u0__abc_49347_n1765) );
  AND2X2 AND2X2_4440 ( .A(u2_u3__abc_47660_n490), .B(u2_u3__abc_47660_n492), .Y(u2_u3__abc_47660_n493) );
  AND2X2 AND2X2_4441 ( .A(u2_u3__abc_47660_n489), .B(u2_u3__abc_47660_n493), .Y(u2_u3__abc_47660_n494) );
  AND2X2 AND2X2_4442 ( .A(u2_u3__abc_47660_n494), .B(u2_u3__abc_47660_n485), .Y(u2_u3__abc_47660_n495) );
  AND2X2 AND2X2_4443 ( .A(u2_u3__abc_47660_n478), .B(u2_u3__abc_47660_n495), .Y(u2_u3__abc_47660_n496) );
  AND2X2 AND2X2_4444 ( .A(u2_u3__abc_47660_n498), .B(u2_u3__abc_47660_n499), .Y(u2_u3__abc_47660_n500) );
  AND2X2 AND2X2_4445 ( .A(row_adr_8_bF_buf2), .B(u2_u3_b1_last_row_8_), .Y(u2_u3__abc_47660_n501) );
  AND2X2 AND2X2_4446 ( .A(u2_u3__abc_47660_n179), .B(u2_u3__abc_47660_n502), .Y(u2_u3__abc_47660_n503) );
  AND2X2 AND2X2_4447 ( .A(u2_u3__abc_47660_n500), .B(u2_u3__abc_47660_n504), .Y(u2_u3__abc_47660_n505) );
  AND2X2 AND2X2_4448 ( .A(u2_u3__abc_47660_n506), .B(u2_u3__abc_47660_n508), .Y(u2_u3__abc_47660_n509) );
  AND2X2 AND2X2_4449 ( .A(u2_u3__abc_47660_n511), .B(u2_u3__abc_47660_n512), .Y(u2_u3__abc_47660_n513) );
  AND2X2 AND2X2_445 ( .A(u0__abc_49347_n1766_1), .B(u0__abc_49347_n1181_bF_buf5), .Y(u0__abc_49347_n1767_1) );
  AND2X2 AND2X2_4450 ( .A(u2_u3__abc_47660_n509), .B(u2_u3__abc_47660_n513), .Y(u2_u3__abc_47660_n514) );
  AND2X2 AND2X2_4451 ( .A(u2_u3__abc_47660_n516), .B(u2_u3__abc_47660_n517), .Y(u2_u3__abc_47660_n518) );
  AND2X2 AND2X2_4452 ( .A(row_adr_6_bF_buf2), .B(u2_u3_b1_last_row_6_), .Y(u2_u3__abc_47660_n519) );
  AND2X2 AND2X2_4453 ( .A(u2_u3__abc_47660_n169), .B(u2_u3__abc_47660_n520), .Y(u2_u3__abc_47660_n521) );
  AND2X2 AND2X2_4454 ( .A(u2_u3__abc_47660_n518), .B(u2_u3__abc_47660_n522), .Y(u2_u3__abc_47660_n523) );
  AND2X2 AND2X2_4455 ( .A(u2_u3__abc_47660_n514), .B(u2_u3__abc_47660_n523), .Y(u2_u3__abc_47660_n524) );
  AND2X2 AND2X2_4456 ( .A(u2_u3__abc_47660_n524), .B(u2_u3__abc_47660_n505), .Y(u2_u3__abc_47660_n525) );
  AND2X2 AND2X2_4457 ( .A(u2_u3__abc_47660_n496), .B(u2_u3__abc_47660_n525), .Y(u2_u3__abc_47660_n526) );
  AND2X2 AND2X2_4458 ( .A(u2_u3__abc_47660_n529), .B(u2_u3__abc_47660_n530), .Y(u2_u3__abc_47660_n531) );
  AND2X2 AND2X2_4459 ( .A(u2_u3__abc_47660_n531), .B(u2_u3__abc_47660_n528), .Y(u2_u3__abc_47660_n532) );
  AND2X2 AND2X2_446 ( .A(spec_req_cs_4_bF_buf2), .B(u0_tms4_24_), .Y(u0__abc_49347_n1768) );
  AND2X2 AND2X2_4460 ( .A(u2_u3__abc_47660_n533), .B(u2_u3__abc_47660_n535), .Y(u2_u3__abc_47660_n536) );
  AND2X2 AND2X2_4461 ( .A(u2_u3__abc_47660_n537), .B(u2_u3__abc_47660_n539), .Y(u2_u3__abc_47660_n540) );
  AND2X2 AND2X2_4462 ( .A(u2_u3__abc_47660_n536), .B(u2_u3__abc_47660_n540), .Y(u2_u3__abc_47660_n541) );
  AND2X2 AND2X2_4463 ( .A(u2_u3__abc_47660_n541), .B(u2_u3__abc_47660_n532), .Y(u2_u3__abc_47660_n542) );
  AND2X2 AND2X2_4464 ( .A(u2_u3__abc_47660_n543), .B(u2_u3__abc_47660_n545), .Y(u2_u3__abc_47660_n546) );
  AND2X2 AND2X2_4465 ( .A(u2_u3__abc_47660_n548), .B(u2_u3__abc_47660_n136), .Y(u2_u3__abc_47660_n549) );
  AND2X2 AND2X2_4466 ( .A(u2_u3__abc_47660_n546), .B(u2_u3__abc_47660_n549), .Y(u2_u3__abc_47660_n550) );
  AND2X2 AND2X2_4467 ( .A(u2_u3__abc_47660_n552), .B(u2_u3__abc_47660_n553), .Y(u2_u3__abc_47660_n554) );
  AND2X2 AND2X2_4468 ( .A(u2_u3__abc_47660_n556), .B(u2_u3__abc_47660_n557), .Y(u2_u3__abc_47660_n558) );
  AND2X2 AND2X2_4469 ( .A(u2_u3__abc_47660_n554), .B(u2_u3__abc_47660_n558), .Y(u2_u3__abc_47660_n559) );
  AND2X2 AND2X2_447 ( .A(u0__abc_49347_n1769), .B(u0__abc_49347_n1180_1_bF_buf5), .Y(u0__abc_49347_n1770) );
  AND2X2 AND2X2_4470 ( .A(u2_u3__abc_47660_n559), .B(u2_u3__abc_47660_n550), .Y(u2_u3__abc_47660_n560) );
  AND2X2 AND2X2_4471 ( .A(u2_u3__abc_47660_n542), .B(u2_u3__abc_47660_n560), .Y(u2_u3__abc_47660_n561) );
  AND2X2 AND2X2_4472 ( .A(u2_u3__abc_47660_n562), .B(u2_u3__abc_47660_n564), .Y(u2_u3__abc_47660_n565) );
  AND2X2 AND2X2_4473 ( .A(u2_u3__abc_47660_n567), .B(u2_u3__abc_47660_n568), .Y(u2_u3__abc_47660_n569) );
  AND2X2 AND2X2_4474 ( .A(u2_u3__abc_47660_n565), .B(u2_u3__abc_47660_n569), .Y(u2_u3__abc_47660_n570) );
  AND2X2 AND2X2_4475 ( .A(u2_u3__abc_47660_n571), .B(u2_u3__abc_47660_n573), .Y(u2_u3__abc_47660_n574) );
  AND2X2 AND2X2_4476 ( .A(u2_u3__abc_47660_n576), .B(u2_u3__abc_47660_n577), .Y(u2_u3__abc_47660_n578) );
  AND2X2 AND2X2_4477 ( .A(u2_u3__abc_47660_n574), .B(u2_u3__abc_47660_n578), .Y(u2_u3__abc_47660_n579) );
  AND2X2 AND2X2_4478 ( .A(u2_u3__abc_47660_n580), .B(u2_u3__abc_47660_n582), .Y(u2_u3__abc_47660_n583) );
  AND2X2 AND2X2_4479 ( .A(u2_u3__abc_47660_n584), .B(u2_u3__abc_47660_n586), .Y(u2_u3__abc_47660_n587) );
  AND2X2 AND2X2_448 ( .A(spec_req_cs_3_bF_buf2), .B(u0_tms3_24_), .Y(u0__abc_49347_n1771_1) );
  AND2X2 AND2X2_4480 ( .A(u2_u3__abc_47660_n583), .B(u2_u3__abc_47660_n587), .Y(u2_u3__abc_47660_n588) );
  AND2X2 AND2X2_4481 ( .A(u2_u3__abc_47660_n579), .B(u2_u3__abc_47660_n588), .Y(u2_u3__abc_47660_n589) );
  AND2X2 AND2X2_4482 ( .A(u2_u3__abc_47660_n589), .B(u2_u3__abc_47660_n570), .Y(u2_u3__abc_47660_n590) );
  AND2X2 AND2X2_4483 ( .A(u2_u3__abc_47660_n561), .B(u2_u3__abc_47660_n590), .Y(u2_u3__abc_47660_n591) );
  AND2X2 AND2X2_4484 ( .A(u2_u3__abc_47660_n289), .B(u2_u3_bank0_open), .Y(u2_u3__abc_47660_n594) );
  AND2X2 AND2X2_4485 ( .A(u2_u3__abc_47660_n204), .B(u2_u3_bank2_open), .Y(u2_u3__abc_47660_n595) );
  AND2X2 AND2X2_4486 ( .A(u2_u3__abc_47660_n136), .B(u2_u3_bank3_open), .Y(u2_u3__abc_47660_n597) );
  AND2X2 AND2X2_4487 ( .A(u2_u3__abc_47660_n247), .B(u2_u3_bank1_open), .Y(u2_u3__abc_47660_n598) );
  AND2X2 AND2X2_4488 ( .A(u2_u3__abc_47660_n136), .B(u2_bank_clr_3), .Y(u2_u3__abc_47660_n604) );
  AND2X2 AND2X2_4489 ( .A(u2_u3__abc_47660_n606), .B(u2_u3_bank3_open), .Y(u2_u3__abc_47660_n607) );
  AND2X2 AND2X2_449 ( .A(u0__abc_49347_n1772_1), .B(u0__abc_49347_n1179_bF_buf5), .Y(u0__abc_49347_n1773_1) );
  AND2X2 AND2X2_4490 ( .A(u2_u3__abc_47660_n605), .B(u2_u3__abc_47660_n607), .Y(u2_u3__abc_47660_n608) );
  AND2X2 AND2X2_4491 ( .A(u2_u3__abc_47660_n606), .B(u2_u3_bank2_open), .Y(u2_u3__abc_47660_n613) );
  AND2X2 AND2X2_4492 ( .A(u2_u3__abc_47660_n612), .B(u2_u3__abc_47660_n613), .Y(u2_u3__abc_47660_n614) );
  AND2X2 AND2X2_4493 ( .A(u2_u3__abc_47660_n606), .B(u2_u3_bank1_open), .Y(u2_u3__abc_47660_n618) );
  AND2X2 AND2X2_4494 ( .A(u2_u3__abc_47660_n617), .B(u2_u3__abc_47660_n618), .Y(u2_u3__abc_47660_n619) );
  AND2X2 AND2X2_4495 ( .A(u2_u3__abc_47660_n606), .B(u2_u3_bank0_open), .Y(u2_u3__abc_47660_n623) );
  AND2X2 AND2X2_4496 ( .A(u2_u3__abc_47660_n622), .B(u2_u3__abc_47660_n623), .Y(u2_u3__abc_47660_n624) );
  AND2X2 AND2X2_4497 ( .A(bank_adr_0_bF_buf1), .B(bank_adr_1_bF_buf1), .Y(u2_u4__abc_47660_n136) );
  AND2X2 AND2X2_4498 ( .A(u2_u4__abc_47660_n136), .B(u2_bank_set_4), .Y(u2_u4__abc_47660_n137) );
  AND2X2 AND2X2_4499 ( .A(u2_u4__abc_47660_n137_bF_buf3), .B(u2_u4__abc_47660_n139), .Y(u2_u4__abc_47660_n140) );
  AND2X2 AND2X2_45 ( .A(_abc_55805_n371), .B(_abc_55805_n372), .Y(tms_s_27_) );
  AND2X2 AND2X2_450 ( .A(spec_req_cs_2_bF_buf2), .B(u0_tms2_24_), .Y(u0__abc_49347_n1774_1) );
  AND2X2 AND2X2_4500 ( .A(u2_u4__abc_47660_n141), .B(u2_u4__abc_47660_n138), .Y(u2_u4_b3_last_row_0__FF_INPUT) );
  AND2X2 AND2X2_4501 ( .A(u2_u4__abc_47660_n137_bF_buf1), .B(u2_u4__abc_47660_n144), .Y(u2_u4__abc_47660_n145) );
  AND2X2 AND2X2_4502 ( .A(u2_u4__abc_47660_n146), .B(u2_u4__abc_47660_n143), .Y(u2_u4_b3_last_row_1__FF_INPUT) );
  AND2X2 AND2X2_4503 ( .A(u2_u4__abc_47660_n137_bF_buf4), .B(u2_u4__abc_47660_n149), .Y(u2_u4__abc_47660_n150) );
  AND2X2 AND2X2_4504 ( .A(u2_u4__abc_47660_n151), .B(u2_u4__abc_47660_n148), .Y(u2_u4_b3_last_row_2__FF_INPUT) );
  AND2X2 AND2X2_4505 ( .A(u2_u4__abc_47660_n137_bF_buf2), .B(u2_u4__abc_47660_n154), .Y(u2_u4__abc_47660_n155) );
  AND2X2 AND2X2_4506 ( .A(u2_u4__abc_47660_n156), .B(u2_u4__abc_47660_n153), .Y(u2_u4_b3_last_row_3__FF_INPUT) );
  AND2X2 AND2X2_4507 ( .A(u2_u4__abc_47660_n137_bF_buf0), .B(u2_u4__abc_47660_n159), .Y(u2_u4__abc_47660_n160) );
  AND2X2 AND2X2_4508 ( .A(u2_u4__abc_47660_n161), .B(u2_u4__abc_47660_n158), .Y(u2_u4_b3_last_row_4__FF_INPUT) );
  AND2X2 AND2X2_4509 ( .A(u2_u4__abc_47660_n137_bF_buf3), .B(u2_u4__abc_47660_n164), .Y(u2_u4__abc_47660_n165) );
  AND2X2 AND2X2_451 ( .A(u0__abc_49347_n1775_1), .B(u0__abc_49347_n1178_1_bF_buf5), .Y(u0__abc_49347_n1776_1) );
  AND2X2 AND2X2_4510 ( .A(u2_u4__abc_47660_n166), .B(u2_u4__abc_47660_n163), .Y(u2_u4_b3_last_row_5__FF_INPUT) );
  AND2X2 AND2X2_4511 ( .A(u2_u4__abc_47660_n137_bF_buf1), .B(u2_u4__abc_47660_n169), .Y(u2_u4__abc_47660_n170) );
  AND2X2 AND2X2_4512 ( .A(u2_u4__abc_47660_n171), .B(u2_u4__abc_47660_n168), .Y(u2_u4_b3_last_row_6__FF_INPUT) );
  AND2X2 AND2X2_4513 ( .A(u2_u4__abc_47660_n137_bF_buf4), .B(u2_u4__abc_47660_n174), .Y(u2_u4__abc_47660_n175) );
  AND2X2 AND2X2_4514 ( .A(u2_u4__abc_47660_n176), .B(u2_u4__abc_47660_n173), .Y(u2_u4_b3_last_row_7__FF_INPUT) );
  AND2X2 AND2X2_4515 ( .A(u2_u4__abc_47660_n137_bF_buf2), .B(u2_u4__abc_47660_n179), .Y(u2_u4__abc_47660_n180) );
  AND2X2 AND2X2_4516 ( .A(u2_u4__abc_47660_n181), .B(u2_u4__abc_47660_n178), .Y(u2_u4_b3_last_row_8__FF_INPUT) );
  AND2X2 AND2X2_4517 ( .A(u2_u4__abc_47660_n137_bF_buf0), .B(u2_u4__abc_47660_n184), .Y(u2_u4__abc_47660_n185) );
  AND2X2 AND2X2_4518 ( .A(u2_u4__abc_47660_n186), .B(u2_u4__abc_47660_n183), .Y(u2_u4_b3_last_row_9__FF_INPUT) );
  AND2X2 AND2X2_4519 ( .A(u2_u4__abc_47660_n137_bF_buf3), .B(u2_u4__abc_47660_n189), .Y(u2_u4__abc_47660_n190) );
  AND2X2 AND2X2_452 ( .A(spec_req_cs_1_bF_buf2), .B(u0_tms1_24_), .Y(u0__abc_49347_n1777_1) );
  AND2X2 AND2X2_4520 ( .A(u2_u4__abc_47660_n191), .B(u2_u4__abc_47660_n188), .Y(u2_u4_b3_last_row_10__FF_INPUT) );
  AND2X2 AND2X2_4521 ( .A(u2_u4__abc_47660_n137_bF_buf1), .B(u2_u4__abc_47660_n194), .Y(u2_u4__abc_47660_n195) );
  AND2X2 AND2X2_4522 ( .A(u2_u4__abc_47660_n196), .B(u2_u4__abc_47660_n193), .Y(u2_u4_b3_last_row_11__FF_INPUT) );
  AND2X2 AND2X2_4523 ( .A(u2_u4__abc_47660_n137_bF_buf4), .B(u2_u4__abc_47660_n199), .Y(u2_u4__abc_47660_n200) );
  AND2X2 AND2X2_4524 ( .A(u2_u4__abc_47660_n201), .B(u2_u4__abc_47660_n198), .Y(u2_u4_b3_last_row_12__FF_INPUT) );
  AND2X2 AND2X2_4525 ( .A(u2_u4__abc_47660_n203), .B(bank_adr_1_bF_buf0), .Y(u2_u4__abc_47660_n204) );
  AND2X2 AND2X2_4526 ( .A(u2_u4__abc_47660_n204), .B(u2_bank_set_4), .Y(u2_u4__abc_47660_n205) );
  AND2X2 AND2X2_4527 ( .A(u2_u4__abc_47660_n208), .B(u2_u4__abc_47660_n206), .Y(u2_u4_b2_last_row_0__FF_INPUT) );
  AND2X2 AND2X2_4528 ( .A(u2_u4__abc_47660_n211), .B(u2_u4__abc_47660_n210), .Y(u2_u4_b2_last_row_1__FF_INPUT) );
  AND2X2 AND2X2_4529 ( .A(u2_u4__abc_47660_n214), .B(u2_u4__abc_47660_n213), .Y(u2_u4_b2_last_row_2__FF_INPUT) );
  AND2X2 AND2X2_453 ( .A(u0__abc_49347_n1175_bF_buf2), .B(u0__abc_49347_n1780_1), .Y(u0__abc_49347_n1781_1) );
  AND2X2 AND2X2_4530 ( .A(u2_u4__abc_47660_n217), .B(u2_u4__abc_47660_n216), .Y(u2_u4_b2_last_row_3__FF_INPUT) );
  AND2X2 AND2X2_4531 ( .A(u2_u4__abc_47660_n220), .B(u2_u4__abc_47660_n219), .Y(u2_u4_b2_last_row_4__FF_INPUT) );
  AND2X2 AND2X2_4532 ( .A(u2_u4__abc_47660_n223), .B(u2_u4__abc_47660_n222), .Y(u2_u4_b2_last_row_5__FF_INPUT) );
  AND2X2 AND2X2_4533 ( .A(u2_u4__abc_47660_n226), .B(u2_u4__abc_47660_n225), .Y(u2_u4_b2_last_row_6__FF_INPUT) );
  AND2X2 AND2X2_4534 ( .A(u2_u4__abc_47660_n229), .B(u2_u4__abc_47660_n228), .Y(u2_u4_b2_last_row_7__FF_INPUT) );
  AND2X2 AND2X2_4535 ( .A(u2_u4__abc_47660_n232), .B(u2_u4__abc_47660_n231), .Y(u2_u4_b2_last_row_8__FF_INPUT) );
  AND2X2 AND2X2_4536 ( .A(u2_u4__abc_47660_n235), .B(u2_u4__abc_47660_n234), .Y(u2_u4_b2_last_row_9__FF_INPUT) );
  AND2X2 AND2X2_4537 ( .A(u2_u4__abc_47660_n238), .B(u2_u4__abc_47660_n237), .Y(u2_u4_b2_last_row_10__FF_INPUT) );
  AND2X2 AND2X2_4538 ( .A(u2_u4__abc_47660_n241), .B(u2_u4__abc_47660_n240), .Y(u2_u4_b2_last_row_11__FF_INPUT) );
  AND2X2 AND2X2_4539 ( .A(u2_u4__abc_47660_n244), .B(u2_u4__abc_47660_n243), .Y(u2_u4_b2_last_row_12__FF_INPUT) );
  AND2X2 AND2X2_454 ( .A(u0__abc_49347_n1779_1), .B(u0__abc_49347_n1781_1), .Y(u0__abc_49347_n1782_1) );
  AND2X2 AND2X2_4540 ( .A(u2_u4__abc_47660_n246), .B(bank_adr_0_bF_buf3), .Y(u2_u4__abc_47660_n247) );
  AND2X2 AND2X2_4541 ( .A(u2_u4__abc_47660_n247), .B(u2_bank_set_4), .Y(u2_u4__abc_47660_n248) );
  AND2X2 AND2X2_4542 ( .A(u2_u4__abc_47660_n251), .B(u2_u4__abc_47660_n249), .Y(u2_u4_b1_last_row_0__FF_INPUT) );
  AND2X2 AND2X2_4543 ( .A(u2_u4__abc_47660_n254), .B(u2_u4__abc_47660_n253), .Y(u2_u4_b1_last_row_1__FF_INPUT) );
  AND2X2 AND2X2_4544 ( .A(u2_u4__abc_47660_n257), .B(u2_u4__abc_47660_n256), .Y(u2_u4_b1_last_row_2__FF_INPUT) );
  AND2X2 AND2X2_4545 ( .A(u2_u4__abc_47660_n260), .B(u2_u4__abc_47660_n259), .Y(u2_u4_b1_last_row_3__FF_INPUT) );
  AND2X2 AND2X2_4546 ( .A(u2_u4__abc_47660_n263), .B(u2_u4__abc_47660_n262), .Y(u2_u4_b1_last_row_4__FF_INPUT) );
  AND2X2 AND2X2_4547 ( .A(u2_u4__abc_47660_n266), .B(u2_u4__abc_47660_n265), .Y(u2_u4_b1_last_row_5__FF_INPUT) );
  AND2X2 AND2X2_4548 ( .A(u2_u4__abc_47660_n269), .B(u2_u4__abc_47660_n268), .Y(u2_u4_b1_last_row_6__FF_INPUT) );
  AND2X2 AND2X2_4549 ( .A(u2_u4__abc_47660_n272), .B(u2_u4__abc_47660_n271), .Y(u2_u4_b1_last_row_7__FF_INPUT) );
  AND2X2 AND2X2_455 ( .A(u0__abc_49347_n1176_1_bF_buf2), .B(sp_tms_25_), .Y(u0__abc_49347_n1784_1) );
  AND2X2 AND2X2_4550 ( .A(u2_u4__abc_47660_n275_1), .B(u2_u4__abc_47660_n274), .Y(u2_u4_b1_last_row_8__FF_INPUT) );
  AND2X2 AND2X2_4551 ( .A(u2_u4__abc_47660_n278_1), .B(u2_u4__abc_47660_n277), .Y(u2_u4_b1_last_row_9__FF_INPUT) );
  AND2X2 AND2X2_4552 ( .A(u2_u4__abc_47660_n281), .B(u2_u4__abc_47660_n280), .Y(u2_u4_b1_last_row_10__FF_INPUT) );
  AND2X2 AND2X2_4553 ( .A(u2_u4__abc_47660_n284), .B(u2_u4__abc_47660_n283_1), .Y(u2_u4_b1_last_row_11__FF_INPUT) );
  AND2X2 AND2X2_4554 ( .A(u2_u4__abc_47660_n287_1), .B(u2_u4__abc_47660_n286_1), .Y(u2_u4_b1_last_row_12__FF_INPUT) );
  AND2X2 AND2X2_4555 ( .A(u2_u4__abc_47660_n203), .B(u2_u4__abc_47660_n246), .Y(u2_u4__abc_47660_n289) );
  AND2X2 AND2X2_4556 ( .A(u2_u4__abc_47660_n289), .B(u2_bank_set_4), .Y(u2_u4__abc_47660_n290_1) );
  AND2X2 AND2X2_4557 ( .A(u2_u4__abc_47660_n293), .B(u2_u4__abc_47660_n291), .Y(u2_u4_b0_last_row_0__FF_INPUT) );
  AND2X2 AND2X2_4558 ( .A(u2_u4__abc_47660_n296_1), .B(u2_u4__abc_47660_n295), .Y(u2_u4_b0_last_row_1__FF_INPUT) );
  AND2X2 AND2X2_4559 ( .A(u2_u4__abc_47660_n299), .B(u2_u4__abc_47660_n298), .Y(u2_u4_b0_last_row_2__FF_INPUT) );
  AND2X2 AND2X2_456 ( .A(spec_req_cs_5_bF_buf1), .B(u0_tms5_25_), .Y(u0__abc_49347_n1785_1) );
  AND2X2 AND2X2_4560 ( .A(u2_u4__abc_47660_n302), .B(u2_u4__abc_47660_n301), .Y(u2_u4_b0_last_row_3__FF_INPUT) );
  AND2X2 AND2X2_4561 ( .A(u2_u4__abc_47660_n305_1), .B(u2_u4__abc_47660_n304_1), .Y(u2_u4_b0_last_row_4__FF_INPUT) );
  AND2X2 AND2X2_4562 ( .A(u2_u4__abc_47660_n308), .B(u2_u4__abc_47660_n307), .Y(u2_u4_b0_last_row_5__FF_INPUT) );
  AND2X2 AND2X2_4563 ( .A(u2_u4__abc_47660_n311), .B(u2_u4__abc_47660_n310), .Y(u2_u4_b0_last_row_6__FF_INPUT) );
  AND2X2 AND2X2_4564 ( .A(u2_u4__abc_47660_n314), .B(u2_u4__abc_47660_n313), .Y(u2_u4_b0_last_row_7__FF_INPUT) );
  AND2X2 AND2X2_4565 ( .A(u2_u4__abc_47660_n317), .B(u2_u4__abc_47660_n316), .Y(u2_u4_b0_last_row_8__FF_INPUT) );
  AND2X2 AND2X2_4566 ( .A(u2_u4__abc_47660_n320), .B(u2_u4__abc_47660_n319), .Y(u2_u4_b0_last_row_9__FF_INPUT) );
  AND2X2 AND2X2_4567 ( .A(u2_u4__abc_47660_n323), .B(u2_u4__abc_47660_n322), .Y(u2_u4_b0_last_row_10__FF_INPUT) );
  AND2X2 AND2X2_4568 ( .A(u2_u4__abc_47660_n326), .B(u2_u4__abc_47660_n325), .Y(u2_u4_b0_last_row_11__FF_INPUT) );
  AND2X2 AND2X2_4569 ( .A(u2_u4__abc_47660_n329), .B(u2_u4__abc_47660_n328), .Y(u2_u4_b0_last_row_12__FF_INPUT) );
  AND2X2 AND2X2_457 ( .A(u0__abc_49347_n1787_1), .B(u0__abc_49347_n1185_bF_buf4), .Y(u0__abc_49347_n1788_1) );
  AND2X2 AND2X2_4570 ( .A(u2_u4__abc_47660_n334), .B(u2_u4__abc_47660_n335), .Y(u2_u4__abc_47660_n336) );
  AND2X2 AND2X2_4571 ( .A(u2_u4__abc_47660_n336), .B(u2_u4__abc_47660_n332), .Y(u2_u4__abc_47660_n337) );
  AND2X2 AND2X2_4572 ( .A(u2_u4__abc_47660_n338), .B(u2_u4__abc_47660_n340), .Y(u2_u4__abc_47660_n341) );
  AND2X2 AND2X2_4573 ( .A(u2_u4__abc_47660_n342), .B(u2_u4__abc_47660_n344), .Y(u2_u4__abc_47660_n345) );
  AND2X2 AND2X2_4574 ( .A(u2_u4__abc_47660_n341), .B(u2_u4__abc_47660_n345), .Y(u2_u4__abc_47660_n346) );
  AND2X2 AND2X2_4575 ( .A(u2_u4__abc_47660_n346), .B(u2_u4__abc_47660_n337), .Y(u2_u4__abc_47660_n347) );
  AND2X2 AND2X2_4576 ( .A(u2_u4__abc_47660_n348), .B(u2_u4__abc_47660_n289), .Y(u2_u4__abc_47660_n349) );
  AND2X2 AND2X2_4577 ( .A(u2_u4__abc_47660_n350), .B(u2_u4__abc_47660_n352), .Y(u2_u4__abc_47660_n353) );
  AND2X2 AND2X2_4578 ( .A(u2_u4__abc_47660_n353), .B(u2_u4__abc_47660_n349), .Y(u2_u4__abc_47660_n354) );
  AND2X2 AND2X2_4579 ( .A(u2_u4__abc_47660_n356), .B(u2_u4__abc_47660_n357), .Y(u2_u4__abc_47660_n358) );
  AND2X2 AND2X2_458 ( .A(u0__abc_49347_n1788_1), .B(u0__abc_49347_n1786_1), .Y(u0__abc_49347_n1789_1) );
  AND2X2 AND2X2_4580 ( .A(u2_u4__abc_47660_n359), .B(u2_u4__abc_47660_n361), .Y(u2_u4__abc_47660_n362) );
  AND2X2 AND2X2_4581 ( .A(u2_u4__abc_47660_n358), .B(u2_u4__abc_47660_n362), .Y(u2_u4__abc_47660_n363) );
  AND2X2 AND2X2_4582 ( .A(u2_u4__abc_47660_n363), .B(u2_u4__abc_47660_n354), .Y(u2_u4__abc_47660_n364) );
  AND2X2 AND2X2_4583 ( .A(u2_u4__abc_47660_n347), .B(u2_u4__abc_47660_n364), .Y(u2_u4__abc_47660_n365) );
  AND2X2 AND2X2_4584 ( .A(u2_u4__abc_47660_n367), .B(u2_u4__abc_47660_n368), .Y(u2_u4__abc_47660_n369) );
  AND2X2 AND2X2_4585 ( .A(row_adr_8_bF_buf3), .B(u2_u4_b0_last_row_8_), .Y(u2_u4__abc_47660_n370) );
  AND2X2 AND2X2_4586 ( .A(u2_u4__abc_47660_n179), .B(u2_u4__abc_47660_n371), .Y(u2_u4__abc_47660_n372) );
  AND2X2 AND2X2_4587 ( .A(u2_u4__abc_47660_n369), .B(u2_u4__abc_47660_n373), .Y(u2_u4__abc_47660_n374) );
  AND2X2 AND2X2_4588 ( .A(u2_u4__abc_47660_n375), .B(u2_u4__abc_47660_n377), .Y(u2_u4__abc_47660_n378) );
  AND2X2 AND2X2_4589 ( .A(u2_u4__abc_47660_n380), .B(u2_u4__abc_47660_n381), .Y(u2_u4__abc_47660_n382) );
  AND2X2 AND2X2_459 ( .A(u0__abc_49347_n1790_1), .B(u0__abc_49347_n1181_bF_buf4), .Y(u0__abc_49347_n1791_1) );
  AND2X2 AND2X2_4590 ( .A(u2_u4__abc_47660_n378), .B(u2_u4__abc_47660_n382), .Y(u2_u4__abc_47660_n383) );
  AND2X2 AND2X2_4591 ( .A(u2_u4__abc_47660_n385), .B(u2_u4__abc_47660_n386), .Y(u2_u4__abc_47660_n387) );
  AND2X2 AND2X2_4592 ( .A(row_adr_6_bF_buf3), .B(u2_u4_b0_last_row_6_), .Y(u2_u4__abc_47660_n388) );
  AND2X2 AND2X2_4593 ( .A(u2_u4__abc_47660_n169), .B(u2_u4__abc_47660_n389), .Y(u2_u4__abc_47660_n390) );
  AND2X2 AND2X2_4594 ( .A(u2_u4__abc_47660_n387), .B(u2_u4__abc_47660_n391), .Y(u2_u4__abc_47660_n392) );
  AND2X2 AND2X2_4595 ( .A(u2_u4__abc_47660_n383), .B(u2_u4__abc_47660_n392), .Y(u2_u4__abc_47660_n393) );
  AND2X2 AND2X2_4596 ( .A(u2_u4__abc_47660_n393), .B(u2_u4__abc_47660_n374), .Y(u2_u4__abc_47660_n394) );
  AND2X2 AND2X2_4597 ( .A(u2_u4__abc_47660_n365), .B(u2_u4__abc_47660_n394), .Y(u2_u4__abc_47660_n395) );
  AND2X2 AND2X2_4598 ( .A(u2_u4__abc_47660_n399), .B(u2_u4__abc_47660_n400), .Y(u2_u4__abc_47660_n401) );
  AND2X2 AND2X2_4599 ( .A(u2_u4__abc_47660_n401), .B(u2_u4__abc_47660_n397), .Y(u2_u4__abc_47660_n402) );
  AND2X2 AND2X2_46 ( .A(_abc_55805_n389), .B(_abc_55805_n390), .Y(csc_s_1_) );
  AND2X2 AND2X2_460 ( .A(spec_req_cs_4_bF_buf1), .B(u0_tms4_25_), .Y(u0__abc_49347_n1792_1) );
  AND2X2 AND2X2_4600 ( .A(u2_u4__abc_47660_n403), .B(u2_u4__abc_47660_n405), .Y(u2_u4__abc_47660_n406) );
  AND2X2 AND2X2_4601 ( .A(u2_u4__abc_47660_n407), .B(u2_u4__abc_47660_n409), .Y(u2_u4__abc_47660_n410) );
  AND2X2 AND2X2_4602 ( .A(u2_u4__abc_47660_n406), .B(u2_u4__abc_47660_n410), .Y(u2_u4__abc_47660_n411) );
  AND2X2 AND2X2_4603 ( .A(u2_u4__abc_47660_n411), .B(u2_u4__abc_47660_n402), .Y(u2_u4__abc_47660_n412) );
  AND2X2 AND2X2_4604 ( .A(u2_u4__abc_47660_n413), .B(u2_u4__abc_47660_n204), .Y(u2_u4__abc_47660_n414) );
  AND2X2 AND2X2_4605 ( .A(u2_u4__abc_47660_n415), .B(u2_u4__abc_47660_n417), .Y(u2_u4__abc_47660_n418) );
  AND2X2 AND2X2_4606 ( .A(u2_u4__abc_47660_n418), .B(u2_u4__abc_47660_n414), .Y(u2_u4__abc_47660_n419) );
  AND2X2 AND2X2_4607 ( .A(u2_u4__abc_47660_n421), .B(u2_u4__abc_47660_n422), .Y(u2_u4__abc_47660_n423) );
  AND2X2 AND2X2_4608 ( .A(u2_u4__abc_47660_n424), .B(u2_u4__abc_47660_n426), .Y(u2_u4__abc_47660_n427) );
  AND2X2 AND2X2_4609 ( .A(u2_u4__abc_47660_n423), .B(u2_u4__abc_47660_n427), .Y(u2_u4__abc_47660_n428) );
  AND2X2 AND2X2_461 ( .A(u0__abc_49347_n1793_1), .B(u0__abc_49347_n1180_1_bF_buf4), .Y(u0__abc_49347_n1794_1) );
  AND2X2 AND2X2_4610 ( .A(u2_u4__abc_47660_n428), .B(u2_u4__abc_47660_n419), .Y(u2_u4__abc_47660_n429) );
  AND2X2 AND2X2_4611 ( .A(u2_u4__abc_47660_n412), .B(u2_u4__abc_47660_n429), .Y(u2_u4__abc_47660_n430) );
  AND2X2 AND2X2_4612 ( .A(u2_u4__abc_47660_n432), .B(u2_u4__abc_47660_n433), .Y(u2_u4__abc_47660_n434) );
  AND2X2 AND2X2_4613 ( .A(row_adr_8_bF_buf2), .B(u2_u4_b2_last_row_8_), .Y(u2_u4__abc_47660_n435) );
  AND2X2 AND2X2_4614 ( .A(u2_u4__abc_47660_n179), .B(u2_u4__abc_47660_n436), .Y(u2_u4__abc_47660_n437) );
  AND2X2 AND2X2_4615 ( .A(u2_u4__abc_47660_n434), .B(u2_u4__abc_47660_n438), .Y(u2_u4__abc_47660_n439) );
  AND2X2 AND2X2_4616 ( .A(u2_u4__abc_47660_n440), .B(u2_u4__abc_47660_n442), .Y(u2_u4__abc_47660_n443) );
  AND2X2 AND2X2_4617 ( .A(u2_u4__abc_47660_n445), .B(u2_u4__abc_47660_n446), .Y(u2_u4__abc_47660_n447) );
  AND2X2 AND2X2_4618 ( .A(u2_u4__abc_47660_n443), .B(u2_u4__abc_47660_n447), .Y(u2_u4__abc_47660_n448) );
  AND2X2 AND2X2_4619 ( .A(u2_u4__abc_47660_n450), .B(u2_u4__abc_47660_n451), .Y(u2_u4__abc_47660_n452) );
  AND2X2 AND2X2_462 ( .A(spec_req_cs_3_bF_buf1), .B(u0_tms3_25_), .Y(u0__abc_49347_n1795_1) );
  AND2X2 AND2X2_4620 ( .A(row_adr_6_bF_buf2), .B(u2_u4_b2_last_row_6_), .Y(u2_u4__abc_47660_n453) );
  AND2X2 AND2X2_4621 ( .A(u2_u4__abc_47660_n169), .B(u2_u4__abc_47660_n454), .Y(u2_u4__abc_47660_n455) );
  AND2X2 AND2X2_4622 ( .A(u2_u4__abc_47660_n452), .B(u2_u4__abc_47660_n456), .Y(u2_u4__abc_47660_n457) );
  AND2X2 AND2X2_4623 ( .A(u2_u4__abc_47660_n448), .B(u2_u4__abc_47660_n457), .Y(u2_u4__abc_47660_n458) );
  AND2X2 AND2X2_4624 ( .A(u2_u4__abc_47660_n458), .B(u2_u4__abc_47660_n439), .Y(u2_u4__abc_47660_n459) );
  AND2X2 AND2X2_4625 ( .A(u2_u4__abc_47660_n430), .B(u2_u4__abc_47660_n459), .Y(u2_u4__abc_47660_n460) );
  AND2X2 AND2X2_4626 ( .A(u2_u4__abc_47660_n465), .B(u2_u4__abc_47660_n466), .Y(u2_u4__abc_47660_n467) );
  AND2X2 AND2X2_4627 ( .A(u2_u4__abc_47660_n467), .B(u2_u4__abc_47660_n463), .Y(u2_u4__abc_47660_n468) );
  AND2X2 AND2X2_4628 ( .A(u2_u4__abc_47660_n469), .B(u2_u4__abc_47660_n471), .Y(u2_u4__abc_47660_n472) );
  AND2X2 AND2X2_4629 ( .A(u2_u4__abc_47660_n473), .B(u2_u4__abc_47660_n475), .Y(u2_u4__abc_47660_n476) );
  AND2X2 AND2X2_463 ( .A(u0__abc_49347_n1796_1), .B(u0__abc_49347_n1179_bF_buf4), .Y(u0__abc_49347_n1797_1) );
  AND2X2 AND2X2_4630 ( .A(u2_u4__abc_47660_n472), .B(u2_u4__abc_47660_n476), .Y(u2_u4__abc_47660_n477) );
  AND2X2 AND2X2_4631 ( .A(u2_u4__abc_47660_n477), .B(u2_u4__abc_47660_n468), .Y(u2_u4__abc_47660_n478) );
  AND2X2 AND2X2_4632 ( .A(u2_u4__abc_47660_n479), .B(u2_u4__abc_47660_n247), .Y(u2_u4__abc_47660_n480) );
  AND2X2 AND2X2_4633 ( .A(u2_u4__abc_47660_n481), .B(u2_u4__abc_47660_n483), .Y(u2_u4__abc_47660_n484) );
  AND2X2 AND2X2_4634 ( .A(u2_u4__abc_47660_n484), .B(u2_u4__abc_47660_n480), .Y(u2_u4__abc_47660_n485) );
  AND2X2 AND2X2_4635 ( .A(u2_u4__abc_47660_n487), .B(u2_u4__abc_47660_n488), .Y(u2_u4__abc_47660_n489) );
  AND2X2 AND2X2_4636 ( .A(u2_u4__abc_47660_n490), .B(u2_u4__abc_47660_n492), .Y(u2_u4__abc_47660_n493) );
  AND2X2 AND2X2_4637 ( .A(u2_u4__abc_47660_n489), .B(u2_u4__abc_47660_n493), .Y(u2_u4__abc_47660_n494) );
  AND2X2 AND2X2_4638 ( .A(u2_u4__abc_47660_n494), .B(u2_u4__abc_47660_n485), .Y(u2_u4__abc_47660_n495) );
  AND2X2 AND2X2_4639 ( .A(u2_u4__abc_47660_n478), .B(u2_u4__abc_47660_n495), .Y(u2_u4__abc_47660_n496) );
  AND2X2 AND2X2_464 ( .A(spec_req_cs_2_bF_buf1), .B(u0_tms2_25_), .Y(u0__abc_49347_n1798_1) );
  AND2X2 AND2X2_4640 ( .A(u2_u4__abc_47660_n498), .B(u2_u4__abc_47660_n499), .Y(u2_u4__abc_47660_n500) );
  AND2X2 AND2X2_4641 ( .A(row_adr_8_bF_buf1), .B(u2_u4_b1_last_row_8_), .Y(u2_u4__abc_47660_n501) );
  AND2X2 AND2X2_4642 ( .A(u2_u4__abc_47660_n179), .B(u2_u4__abc_47660_n502), .Y(u2_u4__abc_47660_n503) );
  AND2X2 AND2X2_4643 ( .A(u2_u4__abc_47660_n500), .B(u2_u4__abc_47660_n504), .Y(u2_u4__abc_47660_n505) );
  AND2X2 AND2X2_4644 ( .A(u2_u4__abc_47660_n506), .B(u2_u4__abc_47660_n508), .Y(u2_u4__abc_47660_n509) );
  AND2X2 AND2X2_4645 ( .A(u2_u4__abc_47660_n511), .B(u2_u4__abc_47660_n512), .Y(u2_u4__abc_47660_n513) );
  AND2X2 AND2X2_4646 ( .A(u2_u4__abc_47660_n509), .B(u2_u4__abc_47660_n513), .Y(u2_u4__abc_47660_n514) );
  AND2X2 AND2X2_4647 ( .A(u2_u4__abc_47660_n516), .B(u2_u4__abc_47660_n517), .Y(u2_u4__abc_47660_n518) );
  AND2X2 AND2X2_4648 ( .A(row_adr_6_bF_buf1), .B(u2_u4_b1_last_row_6_), .Y(u2_u4__abc_47660_n519) );
  AND2X2 AND2X2_4649 ( .A(u2_u4__abc_47660_n169), .B(u2_u4__abc_47660_n520), .Y(u2_u4__abc_47660_n521) );
  AND2X2 AND2X2_465 ( .A(u0__abc_49347_n1799_1), .B(u0__abc_49347_n1178_1_bF_buf4), .Y(u0__abc_49347_n1800_1) );
  AND2X2 AND2X2_4650 ( .A(u2_u4__abc_47660_n518), .B(u2_u4__abc_47660_n522), .Y(u2_u4__abc_47660_n523) );
  AND2X2 AND2X2_4651 ( .A(u2_u4__abc_47660_n514), .B(u2_u4__abc_47660_n523), .Y(u2_u4__abc_47660_n524) );
  AND2X2 AND2X2_4652 ( .A(u2_u4__abc_47660_n524), .B(u2_u4__abc_47660_n505), .Y(u2_u4__abc_47660_n525) );
  AND2X2 AND2X2_4653 ( .A(u2_u4__abc_47660_n496), .B(u2_u4__abc_47660_n525), .Y(u2_u4__abc_47660_n526) );
  AND2X2 AND2X2_4654 ( .A(u2_u4__abc_47660_n529), .B(u2_u4__abc_47660_n530), .Y(u2_u4__abc_47660_n531) );
  AND2X2 AND2X2_4655 ( .A(u2_u4__abc_47660_n531), .B(u2_u4__abc_47660_n528), .Y(u2_u4__abc_47660_n532) );
  AND2X2 AND2X2_4656 ( .A(u2_u4__abc_47660_n533), .B(u2_u4__abc_47660_n535), .Y(u2_u4__abc_47660_n536) );
  AND2X2 AND2X2_4657 ( .A(u2_u4__abc_47660_n537), .B(u2_u4__abc_47660_n539), .Y(u2_u4__abc_47660_n540) );
  AND2X2 AND2X2_4658 ( .A(u2_u4__abc_47660_n536), .B(u2_u4__abc_47660_n540), .Y(u2_u4__abc_47660_n541) );
  AND2X2 AND2X2_4659 ( .A(u2_u4__abc_47660_n541), .B(u2_u4__abc_47660_n532), .Y(u2_u4__abc_47660_n542) );
  AND2X2 AND2X2_466 ( .A(spec_req_cs_1_bF_buf1), .B(u0_tms1_25_), .Y(u0__abc_49347_n1801_1) );
  AND2X2 AND2X2_4660 ( .A(u2_u4__abc_47660_n543), .B(u2_u4__abc_47660_n545), .Y(u2_u4__abc_47660_n546) );
  AND2X2 AND2X2_4661 ( .A(u2_u4__abc_47660_n548), .B(u2_u4__abc_47660_n136), .Y(u2_u4__abc_47660_n549) );
  AND2X2 AND2X2_4662 ( .A(u2_u4__abc_47660_n546), .B(u2_u4__abc_47660_n549), .Y(u2_u4__abc_47660_n550) );
  AND2X2 AND2X2_4663 ( .A(u2_u4__abc_47660_n552), .B(u2_u4__abc_47660_n553), .Y(u2_u4__abc_47660_n554) );
  AND2X2 AND2X2_4664 ( .A(u2_u4__abc_47660_n556), .B(u2_u4__abc_47660_n557), .Y(u2_u4__abc_47660_n558) );
  AND2X2 AND2X2_4665 ( .A(u2_u4__abc_47660_n554), .B(u2_u4__abc_47660_n558), .Y(u2_u4__abc_47660_n559) );
  AND2X2 AND2X2_4666 ( .A(u2_u4__abc_47660_n559), .B(u2_u4__abc_47660_n550), .Y(u2_u4__abc_47660_n560) );
  AND2X2 AND2X2_4667 ( .A(u2_u4__abc_47660_n542), .B(u2_u4__abc_47660_n560), .Y(u2_u4__abc_47660_n561) );
  AND2X2 AND2X2_4668 ( .A(u2_u4__abc_47660_n562), .B(u2_u4__abc_47660_n564), .Y(u2_u4__abc_47660_n565) );
  AND2X2 AND2X2_4669 ( .A(u2_u4__abc_47660_n567), .B(u2_u4__abc_47660_n568), .Y(u2_u4__abc_47660_n569) );
  AND2X2 AND2X2_467 ( .A(u0__abc_49347_n1175_bF_buf1), .B(u0__abc_49347_n1804_1), .Y(u0__abc_49347_n1805_1) );
  AND2X2 AND2X2_4670 ( .A(u2_u4__abc_47660_n565), .B(u2_u4__abc_47660_n569), .Y(u2_u4__abc_47660_n570) );
  AND2X2 AND2X2_4671 ( .A(u2_u4__abc_47660_n571), .B(u2_u4__abc_47660_n573), .Y(u2_u4__abc_47660_n574) );
  AND2X2 AND2X2_4672 ( .A(u2_u4__abc_47660_n576), .B(u2_u4__abc_47660_n577), .Y(u2_u4__abc_47660_n578) );
  AND2X2 AND2X2_4673 ( .A(u2_u4__abc_47660_n574), .B(u2_u4__abc_47660_n578), .Y(u2_u4__abc_47660_n579) );
  AND2X2 AND2X2_4674 ( .A(u2_u4__abc_47660_n580), .B(u2_u4__abc_47660_n582), .Y(u2_u4__abc_47660_n583) );
  AND2X2 AND2X2_4675 ( .A(u2_u4__abc_47660_n584), .B(u2_u4__abc_47660_n586), .Y(u2_u4__abc_47660_n587) );
  AND2X2 AND2X2_4676 ( .A(u2_u4__abc_47660_n583), .B(u2_u4__abc_47660_n587), .Y(u2_u4__abc_47660_n588) );
  AND2X2 AND2X2_4677 ( .A(u2_u4__abc_47660_n579), .B(u2_u4__abc_47660_n588), .Y(u2_u4__abc_47660_n589) );
  AND2X2 AND2X2_4678 ( .A(u2_u4__abc_47660_n589), .B(u2_u4__abc_47660_n570), .Y(u2_u4__abc_47660_n590) );
  AND2X2 AND2X2_4679 ( .A(u2_u4__abc_47660_n561), .B(u2_u4__abc_47660_n590), .Y(u2_u4__abc_47660_n591) );
  AND2X2 AND2X2_468 ( .A(u0__abc_49347_n1803_1), .B(u0__abc_49347_n1805_1), .Y(u0__abc_49347_n1806_1) );
  AND2X2 AND2X2_4680 ( .A(u2_u4__abc_47660_n289), .B(u2_u4_bank0_open), .Y(u2_u4__abc_47660_n594) );
  AND2X2 AND2X2_4681 ( .A(u2_u4__abc_47660_n204), .B(u2_u4_bank2_open), .Y(u2_u4__abc_47660_n595) );
  AND2X2 AND2X2_4682 ( .A(u2_u4__abc_47660_n136), .B(u2_u4_bank3_open), .Y(u2_u4__abc_47660_n597) );
  AND2X2 AND2X2_4683 ( .A(u2_u4__abc_47660_n247), .B(u2_u4_bank1_open), .Y(u2_u4__abc_47660_n598) );
  AND2X2 AND2X2_4684 ( .A(u2_u4__abc_47660_n136), .B(u2_bank_clr_4), .Y(u2_u4__abc_47660_n604) );
  AND2X2 AND2X2_4685 ( .A(u2_u4__abc_47660_n606), .B(u2_u4_bank3_open), .Y(u2_u4__abc_47660_n607) );
  AND2X2 AND2X2_4686 ( .A(u2_u4__abc_47660_n605), .B(u2_u4__abc_47660_n607), .Y(u2_u4__abc_47660_n608) );
  AND2X2 AND2X2_4687 ( .A(u2_u4__abc_47660_n606), .B(u2_u4_bank2_open), .Y(u2_u4__abc_47660_n613) );
  AND2X2 AND2X2_4688 ( .A(u2_u4__abc_47660_n612), .B(u2_u4__abc_47660_n613), .Y(u2_u4__abc_47660_n614) );
  AND2X2 AND2X2_4689 ( .A(u2_u4__abc_47660_n606), .B(u2_u4_bank1_open), .Y(u2_u4__abc_47660_n618) );
  AND2X2 AND2X2_469 ( .A(u0__abc_49347_n1176_1_bF_buf1), .B(sp_tms_26_), .Y(u0__abc_49347_n1808_1) );
  AND2X2 AND2X2_4690 ( .A(u2_u4__abc_47660_n617), .B(u2_u4__abc_47660_n618), .Y(u2_u4__abc_47660_n619) );
  AND2X2 AND2X2_4691 ( .A(u2_u4__abc_47660_n606), .B(u2_u4_bank0_open), .Y(u2_u4__abc_47660_n623) );
  AND2X2 AND2X2_4692 ( .A(u2_u4__abc_47660_n622), .B(u2_u4__abc_47660_n623), .Y(u2_u4__abc_47660_n624) );
  AND2X2 AND2X2_4693 ( .A(bank_adr_0_bF_buf2), .B(bank_adr_1_bF_buf2), .Y(u2_u5__abc_47660_n136) );
  AND2X2 AND2X2_4694 ( .A(u2_u5__abc_47660_n136), .B(u2_bank_set_5), .Y(u2_u5__abc_47660_n137) );
  AND2X2 AND2X2_4695 ( .A(u2_u5__abc_47660_n137_bF_buf3), .B(u2_u5__abc_47660_n139), .Y(u2_u5__abc_47660_n140) );
  AND2X2 AND2X2_4696 ( .A(u2_u5__abc_47660_n141), .B(u2_u5__abc_47660_n138), .Y(u2_u5_b3_last_row_0__FF_INPUT) );
  AND2X2 AND2X2_4697 ( .A(u2_u5__abc_47660_n137_bF_buf1), .B(u2_u5__abc_47660_n144), .Y(u2_u5__abc_47660_n145) );
  AND2X2 AND2X2_4698 ( .A(u2_u5__abc_47660_n146), .B(u2_u5__abc_47660_n143), .Y(u2_u5_b3_last_row_1__FF_INPUT) );
  AND2X2 AND2X2_4699 ( .A(u2_u5__abc_47660_n137_bF_buf4), .B(u2_u5__abc_47660_n149), .Y(u2_u5__abc_47660_n150) );
  AND2X2 AND2X2_47 ( .A(_abc_55805_n392), .B(_abc_55805_n393), .Y(csc_s_2_) );
  AND2X2 AND2X2_470 ( .A(spec_req_cs_5_bF_buf0), .B(u0_tms5_26_), .Y(u0__abc_49347_n1809_1) );
  AND2X2 AND2X2_4700 ( .A(u2_u5__abc_47660_n151), .B(u2_u5__abc_47660_n148), .Y(u2_u5_b3_last_row_2__FF_INPUT) );
  AND2X2 AND2X2_4701 ( .A(u2_u5__abc_47660_n137_bF_buf2), .B(u2_u5__abc_47660_n154), .Y(u2_u5__abc_47660_n155) );
  AND2X2 AND2X2_4702 ( .A(u2_u5__abc_47660_n156), .B(u2_u5__abc_47660_n153), .Y(u2_u5_b3_last_row_3__FF_INPUT) );
  AND2X2 AND2X2_4703 ( .A(u2_u5__abc_47660_n137_bF_buf0), .B(u2_u5__abc_47660_n159), .Y(u2_u5__abc_47660_n160) );
  AND2X2 AND2X2_4704 ( .A(u2_u5__abc_47660_n161), .B(u2_u5__abc_47660_n158), .Y(u2_u5_b3_last_row_4__FF_INPUT) );
  AND2X2 AND2X2_4705 ( .A(u2_u5__abc_47660_n137_bF_buf3), .B(u2_u5__abc_47660_n164), .Y(u2_u5__abc_47660_n165) );
  AND2X2 AND2X2_4706 ( .A(u2_u5__abc_47660_n166), .B(u2_u5__abc_47660_n163), .Y(u2_u5_b3_last_row_5__FF_INPUT) );
  AND2X2 AND2X2_4707 ( .A(u2_u5__abc_47660_n137_bF_buf1), .B(u2_u5__abc_47660_n169), .Y(u2_u5__abc_47660_n170) );
  AND2X2 AND2X2_4708 ( .A(u2_u5__abc_47660_n171), .B(u2_u5__abc_47660_n168), .Y(u2_u5_b3_last_row_6__FF_INPUT) );
  AND2X2 AND2X2_4709 ( .A(u2_u5__abc_47660_n137_bF_buf4), .B(u2_u5__abc_47660_n174), .Y(u2_u5__abc_47660_n175) );
  AND2X2 AND2X2_471 ( .A(u0__abc_49347_n1811_1), .B(u0__abc_49347_n1185_bF_buf3), .Y(u0__abc_49347_n1812_1) );
  AND2X2 AND2X2_4710 ( .A(u2_u5__abc_47660_n176), .B(u2_u5__abc_47660_n173), .Y(u2_u5_b3_last_row_7__FF_INPUT) );
  AND2X2 AND2X2_4711 ( .A(u2_u5__abc_47660_n137_bF_buf2), .B(u2_u5__abc_47660_n179), .Y(u2_u5__abc_47660_n180) );
  AND2X2 AND2X2_4712 ( .A(u2_u5__abc_47660_n181), .B(u2_u5__abc_47660_n178), .Y(u2_u5_b3_last_row_8__FF_INPUT) );
  AND2X2 AND2X2_4713 ( .A(u2_u5__abc_47660_n137_bF_buf0), .B(u2_u5__abc_47660_n184), .Y(u2_u5__abc_47660_n185) );
  AND2X2 AND2X2_4714 ( .A(u2_u5__abc_47660_n186), .B(u2_u5__abc_47660_n183), .Y(u2_u5_b3_last_row_9__FF_INPUT) );
  AND2X2 AND2X2_4715 ( .A(u2_u5__abc_47660_n137_bF_buf3), .B(u2_u5__abc_47660_n189), .Y(u2_u5__abc_47660_n190) );
  AND2X2 AND2X2_4716 ( .A(u2_u5__abc_47660_n191), .B(u2_u5__abc_47660_n188), .Y(u2_u5_b3_last_row_10__FF_INPUT) );
  AND2X2 AND2X2_4717 ( .A(u2_u5__abc_47660_n137_bF_buf1), .B(u2_u5__abc_47660_n194), .Y(u2_u5__abc_47660_n195) );
  AND2X2 AND2X2_4718 ( .A(u2_u5__abc_47660_n196), .B(u2_u5__abc_47660_n193), .Y(u2_u5_b3_last_row_11__FF_INPUT) );
  AND2X2 AND2X2_4719 ( .A(u2_u5__abc_47660_n137_bF_buf4), .B(u2_u5__abc_47660_n199), .Y(u2_u5__abc_47660_n200) );
  AND2X2 AND2X2_472 ( .A(u0__abc_49347_n1812_1), .B(u0__abc_49347_n1810_1), .Y(u0__abc_49347_n1813_1) );
  AND2X2 AND2X2_4720 ( .A(u2_u5__abc_47660_n201), .B(u2_u5__abc_47660_n198), .Y(u2_u5_b3_last_row_12__FF_INPUT) );
  AND2X2 AND2X2_4721 ( .A(u2_u5__abc_47660_n203), .B(bank_adr_1_bF_buf1), .Y(u2_u5__abc_47660_n204) );
  AND2X2 AND2X2_4722 ( .A(u2_u5__abc_47660_n204), .B(u2_bank_set_5), .Y(u2_u5__abc_47660_n205) );
  AND2X2 AND2X2_4723 ( .A(u2_u5__abc_47660_n208), .B(u2_u5__abc_47660_n206), .Y(u2_u5_b2_last_row_0__FF_INPUT) );
  AND2X2 AND2X2_4724 ( .A(u2_u5__abc_47660_n211), .B(u2_u5__abc_47660_n210), .Y(u2_u5_b2_last_row_1__FF_INPUT) );
  AND2X2 AND2X2_4725 ( .A(u2_u5__abc_47660_n214), .B(u2_u5__abc_47660_n213), .Y(u2_u5_b2_last_row_2__FF_INPUT) );
  AND2X2 AND2X2_4726 ( .A(u2_u5__abc_47660_n217), .B(u2_u5__abc_47660_n216), .Y(u2_u5_b2_last_row_3__FF_INPUT) );
  AND2X2 AND2X2_4727 ( .A(u2_u5__abc_47660_n220), .B(u2_u5__abc_47660_n219), .Y(u2_u5_b2_last_row_4__FF_INPUT) );
  AND2X2 AND2X2_4728 ( .A(u2_u5__abc_47660_n223), .B(u2_u5__abc_47660_n222), .Y(u2_u5_b2_last_row_5__FF_INPUT) );
  AND2X2 AND2X2_4729 ( .A(u2_u5__abc_47660_n226), .B(u2_u5__abc_47660_n225), .Y(u2_u5_b2_last_row_6__FF_INPUT) );
  AND2X2 AND2X2_473 ( .A(u0__abc_49347_n1814_1), .B(u0__abc_49347_n1181_bF_buf3), .Y(u0__abc_49347_n1815_1) );
  AND2X2 AND2X2_4730 ( .A(u2_u5__abc_47660_n229), .B(u2_u5__abc_47660_n228), .Y(u2_u5_b2_last_row_7__FF_INPUT) );
  AND2X2 AND2X2_4731 ( .A(u2_u5__abc_47660_n232), .B(u2_u5__abc_47660_n231), .Y(u2_u5_b2_last_row_8__FF_INPUT) );
  AND2X2 AND2X2_4732 ( .A(u2_u5__abc_47660_n235), .B(u2_u5__abc_47660_n234), .Y(u2_u5_b2_last_row_9__FF_INPUT) );
  AND2X2 AND2X2_4733 ( .A(u2_u5__abc_47660_n238), .B(u2_u5__abc_47660_n237), .Y(u2_u5_b2_last_row_10__FF_INPUT) );
  AND2X2 AND2X2_4734 ( .A(u2_u5__abc_47660_n241), .B(u2_u5__abc_47660_n240), .Y(u2_u5_b2_last_row_11__FF_INPUT) );
  AND2X2 AND2X2_4735 ( .A(u2_u5__abc_47660_n244), .B(u2_u5__abc_47660_n243), .Y(u2_u5_b2_last_row_12__FF_INPUT) );
  AND2X2 AND2X2_4736 ( .A(u2_u5__abc_47660_n246), .B(bank_adr_0_bF_buf0), .Y(u2_u5__abc_47660_n247) );
  AND2X2 AND2X2_4737 ( .A(u2_u5__abc_47660_n247), .B(u2_bank_set_5), .Y(u2_u5__abc_47660_n248) );
  AND2X2 AND2X2_4738 ( .A(u2_u5__abc_47660_n251), .B(u2_u5__abc_47660_n249), .Y(u2_u5_b1_last_row_0__FF_INPUT) );
  AND2X2 AND2X2_4739 ( .A(u2_u5__abc_47660_n254), .B(u2_u5__abc_47660_n253), .Y(u2_u5_b1_last_row_1__FF_INPUT) );
  AND2X2 AND2X2_474 ( .A(spec_req_cs_4_bF_buf0), .B(u0_tms4_26_), .Y(u0__abc_49347_n1816_1) );
  AND2X2 AND2X2_4740 ( .A(u2_u5__abc_47660_n257), .B(u2_u5__abc_47660_n256), .Y(u2_u5_b1_last_row_2__FF_INPUT) );
  AND2X2 AND2X2_4741 ( .A(u2_u5__abc_47660_n260), .B(u2_u5__abc_47660_n259), .Y(u2_u5_b1_last_row_3__FF_INPUT) );
  AND2X2 AND2X2_4742 ( .A(u2_u5__abc_47660_n263), .B(u2_u5__abc_47660_n262), .Y(u2_u5_b1_last_row_4__FF_INPUT) );
  AND2X2 AND2X2_4743 ( .A(u2_u5__abc_47660_n266), .B(u2_u5__abc_47660_n265), .Y(u2_u5_b1_last_row_5__FF_INPUT) );
  AND2X2 AND2X2_4744 ( .A(u2_u5__abc_47660_n269), .B(u2_u5__abc_47660_n268), .Y(u2_u5_b1_last_row_6__FF_INPUT) );
  AND2X2 AND2X2_4745 ( .A(u2_u5__abc_47660_n272), .B(u2_u5__abc_47660_n271), .Y(u2_u5_b1_last_row_7__FF_INPUT) );
  AND2X2 AND2X2_4746 ( .A(u2_u5__abc_47660_n275_1), .B(u2_u5__abc_47660_n274), .Y(u2_u5_b1_last_row_8__FF_INPUT) );
  AND2X2 AND2X2_4747 ( .A(u2_u5__abc_47660_n278_1), .B(u2_u5__abc_47660_n277), .Y(u2_u5_b1_last_row_9__FF_INPUT) );
  AND2X2 AND2X2_4748 ( .A(u2_u5__abc_47660_n281), .B(u2_u5__abc_47660_n280), .Y(u2_u5_b1_last_row_10__FF_INPUT) );
  AND2X2 AND2X2_4749 ( .A(u2_u5__abc_47660_n284), .B(u2_u5__abc_47660_n283_1), .Y(u2_u5_b1_last_row_11__FF_INPUT) );
  AND2X2 AND2X2_475 ( .A(u0__abc_49347_n1817_1), .B(u0__abc_49347_n1180_1_bF_buf3), .Y(u0__abc_49347_n1818_1) );
  AND2X2 AND2X2_4750 ( .A(u2_u5__abc_47660_n287_1), .B(u2_u5__abc_47660_n286_1), .Y(u2_u5_b1_last_row_12__FF_INPUT) );
  AND2X2 AND2X2_4751 ( .A(u2_u5__abc_47660_n203), .B(u2_u5__abc_47660_n246), .Y(u2_u5__abc_47660_n289) );
  AND2X2 AND2X2_4752 ( .A(u2_u5__abc_47660_n289), .B(u2_bank_set_5), .Y(u2_u5__abc_47660_n290_1) );
  AND2X2 AND2X2_4753 ( .A(u2_u5__abc_47660_n293), .B(u2_u5__abc_47660_n291), .Y(u2_u5_b0_last_row_0__FF_INPUT) );
  AND2X2 AND2X2_4754 ( .A(u2_u5__abc_47660_n296_1), .B(u2_u5__abc_47660_n295), .Y(u2_u5_b0_last_row_1__FF_INPUT) );
  AND2X2 AND2X2_4755 ( .A(u2_u5__abc_47660_n299), .B(u2_u5__abc_47660_n298), .Y(u2_u5_b0_last_row_2__FF_INPUT) );
  AND2X2 AND2X2_4756 ( .A(u2_u5__abc_47660_n302), .B(u2_u5__abc_47660_n301), .Y(u2_u5_b0_last_row_3__FF_INPUT) );
  AND2X2 AND2X2_4757 ( .A(u2_u5__abc_47660_n305_1), .B(u2_u5__abc_47660_n304_1), .Y(u2_u5_b0_last_row_4__FF_INPUT) );
  AND2X2 AND2X2_4758 ( .A(u2_u5__abc_47660_n308), .B(u2_u5__abc_47660_n307), .Y(u2_u5_b0_last_row_5__FF_INPUT) );
  AND2X2 AND2X2_4759 ( .A(u2_u5__abc_47660_n311), .B(u2_u5__abc_47660_n310), .Y(u2_u5_b0_last_row_6__FF_INPUT) );
  AND2X2 AND2X2_476 ( .A(spec_req_cs_3_bF_buf0), .B(u0_tms3_26_), .Y(u0__abc_49347_n1819_1) );
  AND2X2 AND2X2_4760 ( .A(u2_u5__abc_47660_n314), .B(u2_u5__abc_47660_n313), .Y(u2_u5_b0_last_row_7__FF_INPUT) );
  AND2X2 AND2X2_4761 ( .A(u2_u5__abc_47660_n317), .B(u2_u5__abc_47660_n316), .Y(u2_u5_b0_last_row_8__FF_INPUT) );
  AND2X2 AND2X2_4762 ( .A(u2_u5__abc_47660_n320), .B(u2_u5__abc_47660_n319), .Y(u2_u5_b0_last_row_9__FF_INPUT) );
  AND2X2 AND2X2_4763 ( .A(u2_u5__abc_47660_n323), .B(u2_u5__abc_47660_n322), .Y(u2_u5_b0_last_row_10__FF_INPUT) );
  AND2X2 AND2X2_4764 ( .A(u2_u5__abc_47660_n326), .B(u2_u5__abc_47660_n325), .Y(u2_u5_b0_last_row_11__FF_INPUT) );
  AND2X2 AND2X2_4765 ( .A(u2_u5__abc_47660_n329), .B(u2_u5__abc_47660_n328), .Y(u2_u5_b0_last_row_12__FF_INPUT) );
  AND2X2 AND2X2_4766 ( .A(u2_u5__abc_47660_n334), .B(u2_u5__abc_47660_n335), .Y(u2_u5__abc_47660_n336) );
  AND2X2 AND2X2_4767 ( .A(u2_u5__abc_47660_n336), .B(u2_u5__abc_47660_n332), .Y(u2_u5__abc_47660_n337) );
  AND2X2 AND2X2_4768 ( .A(u2_u5__abc_47660_n338), .B(u2_u5__abc_47660_n340), .Y(u2_u5__abc_47660_n341) );
  AND2X2 AND2X2_4769 ( .A(u2_u5__abc_47660_n342), .B(u2_u5__abc_47660_n344), .Y(u2_u5__abc_47660_n345) );
  AND2X2 AND2X2_477 ( .A(u0__abc_49347_n1820_1), .B(u0__abc_49347_n1179_bF_buf3), .Y(u0__abc_49347_n1821_1) );
  AND2X2 AND2X2_4770 ( .A(u2_u5__abc_47660_n341), .B(u2_u5__abc_47660_n345), .Y(u2_u5__abc_47660_n346) );
  AND2X2 AND2X2_4771 ( .A(u2_u5__abc_47660_n346), .B(u2_u5__abc_47660_n337), .Y(u2_u5__abc_47660_n347) );
  AND2X2 AND2X2_4772 ( .A(u2_u5__abc_47660_n348), .B(u2_u5__abc_47660_n289), .Y(u2_u5__abc_47660_n349) );
  AND2X2 AND2X2_4773 ( .A(u2_u5__abc_47660_n350), .B(u2_u5__abc_47660_n352), .Y(u2_u5__abc_47660_n353) );
  AND2X2 AND2X2_4774 ( .A(u2_u5__abc_47660_n353), .B(u2_u5__abc_47660_n349), .Y(u2_u5__abc_47660_n354) );
  AND2X2 AND2X2_4775 ( .A(u2_u5__abc_47660_n356), .B(u2_u5__abc_47660_n357), .Y(u2_u5__abc_47660_n358) );
  AND2X2 AND2X2_4776 ( .A(u2_u5__abc_47660_n359), .B(u2_u5__abc_47660_n361), .Y(u2_u5__abc_47660_n362) );
  AND2X2 AND2X2_4777 ( .A(u2_u5__abc_47660_n358), .B(u2_u5__abc_47660_n362), .Y(u2_u5__abc_47660_n363) );
  AND2X2 AND2X2_4778 ( .A(u2_u5__abc_47660_n363), .B(u2_u5__abc_47660_n354), .Y(u2_u5__abc_47660_n364) );
  AND2X2 AND2X2_4779 ( .A(u2_u5__abc_47660_n347), .B(u2_u5__abc_47660_n364), .Y(u2_u5__abc_47660_n365) );
  AND2X2 AND2X2_478 ( .A(spec_req_cs_2_bF_buf0), .B(u0_tms2_26_), .Y(u0__abc_49347_n1822_1) );
  AND2X2 AND2X2_4780 ( .A(u2_u5__abc_47660_n367), .B(u2_u5__abc_47660_n368), .Y(u2_u5__abc_47660_n369) );
  AND2X2 AND2X2_4781 ( .A(row_adr_8_bF_buf2), .B(u2_u5_b0_last_row_8_), .Y(u2_u5__abc_47660_n370) );
  AND2X2 AND2X2_4782 ( .A(u2_u5__abc_47660_n179), .B(u2_u5__abc_47660_n371), .Y(u2_u5__abc_47660_n372) );
  AND2X2 AND2X2_4783 ( .A(u2_u5__abc_47660_n369), .B(u2_u5__abc_47660_n373), .Y(u2_u5__abc_47660_n374) );
  AND2X2 AND2X2_4784 ( .A(u2_u5__abc_47660_n375), .B(u2_u5__abc_47660_n377), .Y(u2_u5__abc_47660_n378) );
  AND2X2 AND2X2_4785 ( .A(u2_u5__abc_47660_n380), .B(u2_u5__abc_47660_n381), .Y(u2_u5__abc_47660_n382) );
  AND2X2 AND2X2_4786 ( .A(u2_u5__abc_47660_n378), .B(u2_u5__abc_47660_n382), .Y(u2_u5__abc_47660_n383) );
  AND2X2 AND2X2_4787 ( .A(u2_u5__abc_47660_n385), .B(u2_u5__abc_47660_n386), .Y(u2_u5__abc_47660_n387) );
  AND2X2 AND2X2_4788 ( .A(row_adr_6_bF_buf2), .B(u2_u5_b0_last_row_6_), .Y(u2_u5__abc_47660_n388) );
  AND2X2 AND2X2_4789 ( .A(u2_u5__abc_47660_n169), .B(u2_u5__abc_47660_n389), .Y(u2_u5__abc_47660_n390) );
  AND2X2 AND2X2_479 ( .A(u0__abc_49347_n1823_1), .B(u0__abc_49347_n1178_1_bF_buf3), .Y(u0__abc_49347_n1824_1) );
  AND2X2 AND2X2_4790 ( .A(u2_u5__abc_47660_n387), .B(u2_u5__abc_47660_n391), .Y(u2_u5__abc_47660_n392) );
  AND2X2 AND2X2_4791 ( .A(u2_u5__abc_47660_n383), .B(u2_u5__abc_47660_n392), .Y(u2_u5__abc_47660_n393) );
  AND2X2 AND2X2_4792 ( .A(u2_u5__abc_47660_n393), .B(u2_u5__abc_47660_n374), .Y(u2_u5__abc_47660_n394) );
  AND2X2 AND2X2_4793 ( .A(u2_u5__abc_47660_n365), .B(u2_u5__abc_47660_n394), .Y(u2_u5__abc_47660_n395) );
  AND2X2 AND2X2_4794 ( .A(u2_u5__abc_47660_n399), .B(u2_u5__abc_47660_n400), .Y(u2_u5__abc_47660_n401) );
  AND2X2 AND2X2_4795 ( .A(u2_u5__abc_47660_n401), .B(u2_u5__abc_47660_n397), .Y(u2_u5__abc_47660_n402) );
  AND2X2 AND2X2_4796 ( .A(u2_u5__abc_47660_n403), .B(u2_u5__abc_47660_n405), .Y(u2_u5__abc_47660_n406) );
  AND2X2 AND2X2_4797 ( .A(u2_u5__abc_47660_n407), .B(u2_u5__abc_47660_n409), .Y(u2_u5__abc_47660_n410) );
  AND2X2 AND2X2_4798 ( .A(u2_u5__abc_47660_n406), .B(u2_u5__abc_47660_n410), .Y(u2_u5__abc_47660_n411) );
  AND2X2 AND2X2_4799 ( .A(u2_u5__abc_47660_n411), .B(u2_u5__abc_47660_n402), .Y(u2_u5__abc_47660_n412) );
  AND2X2 AND2X2_48 ( .A(_abc_55805_n395), .B(_abc_55805_n396), .Y(csc_s_3_) );
  AND2X2 AND2X2_480 ( .A(spec_req_cs_1_bF_buf0), .B(u0_tms1_26_), .Y(u0__abc_49347_n1825_1) );
  AND2X2 AND2X2_4800 ( .A(u2_u5__abc_47660_n413), .B(u2_u5__abc_47660_n204), .Y(u2_u5__abc_47660_n414) );
  AND2X2 AND2X2_4801 ( .A(u2_u5__abc_47660_n415), .B(u2_u5__abc_47660_n417), .Y(u2_u5__abc_47660_n418) );
  AND2X2 AND2X2_4802 ( .A(u2_u5__abc_47660_n418), .B(u2_u5__abc_47660_n414), .Y(u2_u5__abc_47660_n419) );
  AND2X2 AND2X2_4803 ( .A(u2_u5__abc_47660_n421), .B(u2_u5__abc_47660_n422), .Y(u2_u5__abc_47660_n423) );
  AND2X2 AND2X2_4804 ( .A(u2_u5__abc_47660_n424), .B(u2_u5__abc_47660_n426), .Y(u2_u5__abc_47660_n427) );
  AND2X2 AND2X2_4805 ( .A(u2_u5__abc_47660_n423), .B(u2_u5__abc_47660_n427), .Y(u2_u5__abc_47660_n428) );
  AND2X2 AND2X2_4806 ( .A(u2_u5__abc_47660_n428), .B(u2_u5__abc_47660_n419), .Y(u2_u5__abc_47660_n429) );
  AND2X2 AND2X2_4807 ( .A(u2_u5__abc_47660_n412), .B(u2_u5__abc_47660_n429), .Y(u2_u5__abc_47660_n430) );
  AND2X2 AND2X2_4808 ( .A(u2_u5__abc_47660_n432), .B(u2_u5__abc_47660_n433), .Y(u2_u5__abc_47660_n434) );
  AND2X2 AND2X2_4809 ( .A(row_adr_8_bF_buf1), .B(u2_u5_b2_last_row_8_), .Y(u2_u5__abc_47660_n435) );
  AND2X2 AND2X2_481 ( .A(u0__abc_49347_n1175_bF_buf0), .B(u0__abc_49347_n1828_1), .Y(u0__abc_49347_n1829_1) );
  AND2X2 AND2X2_4810 ( .A(u2_u5__abc_47660_n179), .B(u2_u5__abc_47660_n436), .Y(u2_u5__abc_47660_n437) );
  AND2X2 AND2X2_4811 ( .A(u2_u5__abc_47660_n434), .B(u2_u5__abc_47660_n438), .Y(u2_u5__abc_47660_n439) );
  AND2X2 AND2X2_4812 ( .A(u2_u5__abc_47660_n440), .B(u2_u5__abc_47660_n442), .Y(u2_u5__abc_47660_n443) );
  AND2X2 AND2X2_4813 ( .A(u2_u5__abc_47660_n445), .B(u2_u5__abc_47660_n446), .Y(u2_u5__abc_47660_n447) );
  AND2X2 AND2X2_4814 ( .A(u2_u5__abc_47660_n443), .B(u2_u5__abc_47660_n447), .Y(u2_u5__abc_47660_n448) );
  AND2X2 AND2X2_4815 ( .A(u2_u5__abc_47660_n450), .B(u2_u5__abc_47660_n451), .Y(u2_u5__abc_47660_n452) );
  AND2X2 AND2X2_4816 ( .A(row_adr_6_bF_buf1), .B(u2_u5_b2_last_row_6_), .Y(u2_u5__abc_47660_n453) );
  AND2X2 AND2X2_4817 ( .A(u2_u5__abc_47660_n169), .B(u2_u5__abc_47660_n454), .Y(u2_u5__abc_47660_n455) );
  AND2X2 AND2X2_4818 ( .A(u2_u5__abc_47660_n452), .B(u2_u5__abc_47660_n456), .Y(u2_u5__abc_47660_n457) );
  AND2X2 AND2X2_4819 ( .A(u2_u5__abc_47660_n448), .B(u2_u5__abc_47660_n457), .Y(u2_u5__abc_47660_n458) );
  AND2X2 AND2X2_482 ( .A(u0__abc_49347_n1827_1), .B(u0__abc_49347_n1829_1), .Y(u0__abc_49347_n1830_1) );
  AND2X2 AND2X2_4820 ( .A(u2_u5__abc_47660_n458), .B(u2_u5__abc_47660_n439), .Y(u2_u5__abc_47660_n459) );
  AND2X2 AND2X2_4821 ( .A(u2_u5__abc_47660_n430), .B(u2_u5__abc_47660_n459), .Y(u2_u5__abc_47660_n460) );
  AND2X2 AND2X2_4822 ( .A(u2_u5__abc_47660_n465), .B(u2_u5__abc_47660_n466), .Y(u2_u5__abc_47660_n467) );
  AND2X2 AND2X2_4823 ( .A(u2_u5__abc_47660_n467), .B(u2_u5__abc_47660_n463), .Y(u2_u5__abc_47660_n468) );
  AND2X2 AND2X2_4824 ( .A(u2_u5__abc_47660_n469), .B(u2_u5__abc_47660_n471), .Y(u2_u5__abc_47660_n472) );
  AND2X2 AND2X2_4825 ( .A(u2_u5__abc_47660_n473), .B(u2_u5__abc_47660_n475), .Y(u2_u5__abc_47660_n476) );
  AND2X2 AND2X2_4826 ( .A(u2_u5__abc_47660_n472), .B(u2_u5__abc_47660_n476), .Y(u2_u5__abc_47660_n477) );
  AND2X2 AND2X2_4827 ( .A(u2_u5__abc_47660_n477), .B(u2_u5__abc_47660_n468), .Y(u2_u5__abc_47660_n478) );
  AND2X2 AND2X2_4828 ( .A(u2_u5__abc_47660_n479), .B(u2_u5__abc_47660_n247), .Y(u2_u5__abc_47660_n480) );
  AND2X2 AND2X2_4829 ( .A(u2_u5__abc_47660_n481), .B(u2_u5__abc_47660_n483), .Y(u2_u5__abc_47660_n484) );
  AND2X2 AND2X2_483 ( .A(u0__abc_49347_n1176_1_bF_buf0), .B(sp_tms_27_), .Y(u0__abc_49347_n1832_1) );
  AND2X2 AND2X2_4830 ( .A(u2_u5__abc_47660_n484), .B(u2_u5__abc_47660_n480), .Y(u2_u5__abc_47660_n485) );
  AND2X2 AND2X2_4831 ( .A(u2_u5__abc_47660_n487), .B(u2_u5__abc_47660_n488), .Y(u2_u5__abc_47660_n489) );
  AND2X2 AND2X2_4832 ( .A(u2_u5__abc_47660_n490), .B(u2_u5__abc_47660_n492), .Y(u2_u5__abc_47660_n493) );
  AND2X2 AND2X2_4833 ( .A(u2_u5__abc_47660_n489), .B(u2_u5__abc_47660_n493), .Y(u2_u5__abc_47660_n494) );
  AND2X2 AND2X2_4834 ( .A(u2_u5__abc_47660_n494), .B(u2_u5__abc_47660_n485), .Y(u2_u5__abc_47660_n495) );
  AND2X2 AND2X2_4835 ( .A(u2_u5__abc_47660_n478), .B(u2_u5__abc_47660_n495), .Y(u2_u5__abc_47660_n496) );
  AND2X2 AND2X2_4836 ( .A(u2_u5__abc_47660_n498), .B(u2_u5__abc_47660_n499), .Y(u2_u5__abc_47660_n500) );
  AND2X2 AND2X2_4837 ( .A(row_adr_8_bF_buf0), .B(u2_u5_b1_last_row_8_), .Y(u2_u5__abc_47660_n501) );
  AND2X2 AND2X2_4838 ( .A(u2_u5__abc_47660_n179), .B(u2_u5__abc_47660_n502), .Y(u2_u5__abc_47660_n503) );
  AND2X2 AND2X2_4839 ( .A(u2_u5__abc_47660_n500), .B(u2_u5__abc_47660_n504), .Y(u2_u5__abc_47660_n505) );
  AND2X2 AND2X2_484 ( .A(spec_req_cs_5_bF_buf5), .B(u0_tms5_27_), .Y(u0__abc_49347_n1833_1) );
  AND2X2 AND2X2_4840 ( .A(u2_u5__abc_47660_n506), .B(u2_u5__abc_47660_n508), .Y(u2_u5__abc_47660_n509) );
  AND2X2 AND2X2_4841 ( .A(u2_u5__abc_47660_n511), .B(u2_u5__abc_47660_n512), .Y(u2_u5__abc_47660_n513) );
  AND2X2 AND2X2_4842 ( .A(u2_u5__abc_47660_n509), .B(u2_u5__abc_47660_n513), .Y(u2_u5__abc_47660_n514) );
  AND2X2 AND2X2_4843 ( .A(u2_u5__abc_47660_n516), .B(u2_u5__abc_47660_n517), .Y(u2_u5__abc_47660_n518) );
  AND2X2 AND2X2_4844 ( .A(row_adr_6_bF_buf0), .B(u2_u5_b1_last_row_6_), .Y(u2_u5__abc_47660_n519) );
  AND2X2 AND2X2_4845 ( .A(u2_u5__abc_47660_n169), .B(u2_u5__abc_47660_n520), .Y(u2_u5__abc_47660_n521) );
  AND2X2 AND2X2_4846 ( .A(u2_u5__abc_47660_n518), .B(u2_u5__abc_47660_n522), .Y(u2_u5__abc_47660_n523) );
  AND2X2 AND2X2_4847 ( .A(u2_u5__abc_47660_n514), .B(u2_u5__abc_47660_n523), .Y(u2_u5__abc_47660_n524) );
  AND2X2 AND2X2_4848 ( .A(u2_u5__abc_47660_n524), .B(u2_u5__abc_47660_n505), .Y(u2_u5__abc_47660_n525) );
  AND2X2 AND2X2_4849 ( .A(u2_u5__abc_47660_n496), .B(u2_u5__abc_47660_n525), .Y(u2_u5__abc_47660_n526) );
  AND2X2 AND2X2_485 ( .A(u0__abc_49347_n1835_1), .B(u0__abc_49347_n1185_bF_buf2), .Y(u0__abc_49347_n1836_1) );
  AND2X2 AND2X2_4850 ( .A(u2_u5__abc_47660_n529), .B(u2_u5__abc_47660_n530), .Y(u2_u5__abc_47660_n531) );
  AND2X2 AND2X2_4851 ( .A(u2_u5__abc_47660_n531), .B(u2_u5__abc_47660_n528), .Y(u2_u5__abc_47660_n532) );
  AND2X2 AND2X2_4852 ( .A(u2_u5__abc_47660_n533), .B(u2_u5__abc_47660_n535), .Y(u2_u5__abc_47660_n536) );
  AND2X2 AND2X2_4853 ( .A(u2_u5__abc_47660_n537), .B(u2_u5__abc_47660_n539), .Y(u2_u5__abc_47660_n540) );
  AND2X2 AND2X2_4854 ( .A(u2_u5__abc_47660_n536), .B(u2_u5__abc_47660_n540), .Y(u2_u5__abc_47660_n541) );
  AND2X2 AND2X2_4855 ( .A(u2_u5__abc_47660_n541), .B(u2_u5__abc_47660_n532), .Y(u2_u5__abc_47660_n542) );
  AND2X2 AND2X2_4856 ( .A(u2_u5__abc_47660_n543), .B(u2_u5__abc_47660_n545), .Y(u2_u5__abc_47660_n546) );
  AND2X2 AND2X2_4857 ( .A(u2_u5__abc_47660_n548), .B(u2_u5__abc_47660_n136), .Y(u2_u5__abc_47660_n549) );
  AND2X2 AND2X2_4858 ( .A(u2_u5__abc_47660_n546), .B(u2_u5__abc_47660_n549), .Y(u2_u5__abc_47660_n550) );
  AND2X2 AND2X2_4859 ( .A(u2_u5__abc_47660_n552), .B(u2_u5__abc_47660_n553), .Y(u2_u5__abc_47660_n554) );
  AND2X2 AND2X2_486 ( .A(u0__abc_49347_n1836_1), .B(u0__abc_49347_n1834_1), .Y(u0__abc_49347_n1837_1) );
  AND2X2 AND2X2_4860 ( .A(u2_u5__abc_47660_n556), .B(u2_u5__abc_47660_n557), .Y(u2_u5__abc_47660_n558) );
  AND2X2 AND2X2_4861 ( .A(u2_u5__abc_47660_n554), .B(u2_u5__abc_47660_n558), .Y(u2_u5__abc_47660_n559) );
  AND2X2 AND2X2_4862 ( .A(u2_u5__abc_47660_n559), .B(u2_u5__abc_47660_n550), .Y(u2_u5__abc_47660_n560) );
  AND2X2 AND2X2_4863 ( .A(u2_u5__abc_47660_n542), .B(u2_u5__abc_47660_n560), .Y(u2_u5__abc_47660_n561) );
  AND2X2 AND2X2_4864 ( .A(u2_u5__abc_47660_n562), .B(u2_u5__abc_47660_n564), .Y(u2_u5__abc_47660_n565) );
  AND2X2 AND2X2_4865 ( .A(u2_u5__abc_47660_n567), .B(u2_u5__abc_47660_n568), .Y(u2_u5__abc_47660_n569) );
  AND2X2 AND2X2_4866 ( .A(u2_u5__abc_47660_n565), .B(u2_u5__abc_47660_n569), .Y(u2_u5__abc_47660_n570) );
  AND2X2 AND2X2_4867 ( .A(u2_u5__abc_47660_n571), .B(u2_u5__abc_47660_n573), .Y(u2_u5__abc_47660_n574) );
  AND2X2 AND2X2_4868 ( .A(u2_u5__abc_47660_n576), .B(u2_u5__abc_47660_n577), .Y(u2_u5__abc_47660_n578) );
  AND2X2 AND2X2_4869 ( .A(u2_u5__abc_47660_n574), .B(u2_u5__abc_47660_n578), .Y(u2_u5__abc_47660_n579) );
  AND2X2 AND2X2_487 ( .A(u0__abc_49347_n1838_1), .B(u0__abc_49347_n1181_bF_buf2), .Y(u0__abc_49347_n1839_1) );
  AND2X2 AND2X2_4870 ( .A(u2_u5__abc_47660_n580), .B(u2_u5__abc_47660_n582), .Y(u2_u5__abc_47660_n583) );
  AND2X2 AND2X2_4871 ( .A(u2_u5__abc_47660_n584), .B(u2_u5__abc_47660_n586), .Y(u2_u5__abc_47660_n587) );
  AND2X2 AND2X2_4872 ( .A(u2_u5__abc_47660_n583), .B(u2_u5__abc_47660_n587), .Y(u2_u5__abc_47660_n588) );
  AND2X2 AND2X2_4873 ( .A(u2_u5__abc_47660_n579), .B(u2_u5__abc_47660_n588), .Y(u2_u5__abc_47660_n589) );
  AND2X2 AND2X2_4874 ( .A(u2_u5__abc_47660_n589), .B(u2_u5__abc_47660_n570), .Y(u2_u5__abc_47660_n590) );
  AND2X2 AND2X2_4875 ( .A(u2_u5__abc_47660_n561), .B(u2_u5__abc_47660_n590), .Y(u2_u5__abc_47660_n591) );
  AND2X2 AND2X2_4876 ( .A(u2_u5__abc_47660_n289), .B(u2_u5_bank0_open), .Y(u2_u5__abc_47660_n594) );
  AND2X2 AND2X2_4877 ( .A(u2_u5__abc_47660_n204), .B(u2_u5_bank2_open), .Y(u2_u5__abc_47660_n595) );
  AND2X2 AND2X2_4878 ( .A(u2_u5__abc_47660_n136), .B(u2_u5_bank3_open), .Y(u2_u5__abc_47660_n597) );
  AND2X2 AND2X2_4879 ( .A(u2_u5__abc_47660_n247), .B(u2_u5_bank1_open), .Y(u2_u5__abc_47660_n598) );
  AND2X2 AND2X2_488 ( .A(spec_req_cs_4_bF_buf5), .B(u0_tms4_27_), .Y(u0__abc_49347_n1840_1) );
  AND2X2 AND2X2_4880 ( .A(u2_u5__abc_47660_n136), .B(u2_bank_clr_5), .Y(u2_u5__abc_47660_n604) );
  AND2X2 AND2X2_4881 ( .A(u2_u5__abc_47660_n606), .B(u2_u5_bank3_open), .Y(u2_u5__abc_47660_n607) );
  AND2X2 AND2X2_4882 ( .A(u2_u5__abc_47660_n605), .B(u2_u5__abc_47660_n607), .Y(u2_u5__abc_47660_n608) );
  AND2X2 AND2X2_4883 ( .A(u2_u5__abc_47660_n606), .B(u2_u5_bank2_open), .Y(u2_u5__abc_47660_n613) );
  AND2X2 AND2X2_4884 ( .A(u2_u5__abc_47660_n612), .B(u2_u5__abc_47660_n613), .Y(u2_u5__abc_47660_n614) );
  AND2X2 AND2X2_4885 ( .A(u2_u5__abc_47660_n606), .B(u2_u5_bank1_open), .Y(u2_u5__abc_47660_n618) );
  AND2X2 AND2X2_4886 ( .A(u2_u5__abc_47660_n617), .B(u2_u5__abc_47660_n618), .Y(u2_u5__abc_47660_n619) );
  AND2X2 AND2X2_4887 ( .A(u2_u5__abc_47660_n606), .B(u2_u5_bank0_open), .Y(u2_u5__abc_47660_n623) );
  AND2X2 AND2X2_4888 ( .A(u2_u5__abc_47660_n622), .B(u2_u5__abc_47660_n623), .Y(u2_u5__abc_47660_n624) );
  AND2X2 AND2X2_4889 ( .A(\wb_data_i[3] ), .B(\wb_data_i[2] ), .Y(u3__abc_46775_n281_1) );
  AND2X2 AND2X2_489 ( .A(u0__abc_49347_n1841_1), .B(u0__abc_49347_n1180_1_bF_buf2), .Y(u0__abc_49347_n1842_1) );
  AND2X2 AND2X2_4890 ( .A(u3__abc_46775_n282_1), .B(u3__abc_46775_n280), .Y(u3__abc_46775_n283) );
  AND2X2 AND2X2_4891 ( .A(u3__abc_46775_n286_1), .B(u3__abc_46775_n288), .Y(u3__abc_46775_n289) );
  AND2X2 AND2X2_4892 ( .A(u3__abc_46775_n284), .B(u3__abc_46775_n289), .Y(u3__abc_46775_n290_1) );
  AND2X2 AND2X2_4893 ( .A(u3__abc_46775_n291_1), .B(u3__abc_46775_n292_1), .Y(u3__abc_46775_n293) );
  AND2X2 AND2X2_4894 ( .A(\wb_data_i[7] ), .B(\wb_data_i[6] ), .Y(u3__abc_46775_n296_1) );
  AND2X2 AND2X2_4895 ( .A(u3__abc_46775_n297_1), .B(u3__abc_46775_n295_1), .Y(u3__abc_46775_n298) );
  AND2X2 AND2X2_4896 ( .A(u3__abc_46775_n301_1), .B(u3__abc_46775_n303), .Y(u3__abc_46775_n304) );
  AND2X2 AND2X2_4897 ( .A(u3__abc_46775_n305_1), .B(u3__abc_46775_n299), .Y(u3__abc_46775_n306_1) );
  AND2X2 AND2X2_4898 ( .A(u3__abc_46775_n304), .B(u3__abc_46775_n298), .Y(u3__abc_46775_n307_1) );
  AND2X2 AND2X2_4899 ( .A(u3__abc_46775_n310_1), .B(u3__abc_46775_n311_1), .Y(u3__abc_46775_n312_1) );
  AND2X2 AND2X2_49 ( .A(_abc_55805_n398), .B(_abc_55805_n399), .Y(csc_s_4_) );
  AND2X2 AND2X2_490 ( .A(spec_req_cs_3_bF_buf5), .B(u0_tms3_27_), .Y(u0__abc_49347_n1843_1) );
  AND2X2 AND2X2_4900 ( .A(u3__abc_46775_n313), .B(u3__abc_46775_n278_1), .Y(u3_mc_dp_o_0__FF_INPUT) );
  AND2X2 AND2X2_4901 ( .A(\wb_data_i[11] ), .B(\wb_data_i[10] ), .Y(u3__abc_46775_n317_1) );
  AND2X2 AND2X2_4902 ( .A(u3__abc_46775_n318), .B(u3__abc_46775_n316_1), .Y(u3__abc_46775_n319) );
  AND2X2 AND2X2_4903 ( .A(u3__abc_46775_n321_1), .B(u3__abc_46775_n323), .Y(u3__abc_46775_n324) );
  AND2X2 AND2X2_4904 ( .A(u3__abc_46775_n325_1), .B(u3__abc_46775_n319), .Y(u3__abc_46775_n326_1) );
  AND2X2 AND2X2_4905 ( .A(u3__abc_46775_n327_1), .B(u3__abc_46775_n328), .Y(u3__abc_46775_n329) );
  AND2X2 AND2X2_4906 ( .A(\wb_data_i[15] ), .B(\wb_data_i[14] ), .Y(u3__abc_46775_n332_1) );
  AND2X2 AND2X2_4907 ( .A(u3__abc_46775_n333), .B(u3__abc_46775_n331_1), .Y(u3__abc_46775_n334) );
  AND2X2 AND2X2_4908 ( .A(u3__abc_46775_n337_1), .B(u3__abc_46775_n339), .Y(u3__abc_46775_n340_1) );
  AND2X2 AND2X2_4909 ( .A(u3__abc_46775_n341_1), .B(u3__abc_46775_n335_1), .Y(u3__abc_46775_n342_1) );
  AND2X2 AND2X2_491 ( .A(u0__abc_49347_n1844_1), .B(u0__abc_49347_n1179_bF_buf2), .Y(u0__abc_49347_n1845_1) );
  AND2X2 AND2X2_4910 ( .A(u3__abc_46775_n340_1), .B(u3__abc_46775_n334), .Y(u3__abc_46775_n343) );
  AND2X2 AND2X2_4911 ( .A(u3__abc_46775_n346_1), .B(u3__abc_46775_n347_1), .Y(u3__abc_46775_n348) );
  AND2X2 AND2X2_4912 ( .A(u3__abc_46775_n349), .B(u3__abc_46775_n315_1), .Y(u3_mc_dp_o_1__FF_INPUT) );
  AND2X2 AND2X2_4913 ( .A(\wb_data_i[19] ), .B(\wb_data_i[18] ), .Y(u3__abc_46775_n352_1) );
  AND2X2 AND2X2_4914 ( .A(u3__abc_46775_n353), .B(u3__abc_46775_n351_1), .Y(u3__abc_46775_n354) );
  AND2X2 AND2X2_4915 ( .A(u3__abc_46775_n356_1), .B(u3__abc_46775_n358), .Y(u3__abc_46775_n359) );
  AND2X2 AND2X2_4916 ( .A(u3__abc_46775_n360_1), .B(u3__abc_46775_n354), .Y(u3__abc_46775_n361_1) );
  AND2X2 AND2X2_4917 ( .A(u3__abc_46775_n362_1), .B(u3__abc_46775_n363), .Y(u3__abc_46775_n364) );
  AND2X2 AND2X2_4918 ( .A(\wb_data_i[23] ), .B(\wb_data_i[22] ), .Y(u3__abc_46775_n366_1) );
  AND2X2 AND2X2_4919 ( .A(u3__abc_46775_n367_1), .B(u3__abc_46775_n365_1), .Y(u3__abc_46775_n368_1) );
  AND2X2 AND2X2_492 ( .A(spec_req_cs_2_bF_buf5), .B(u0_tms2_27_), .Y(u0__abc_49347_n1846_1) );
  AND2X2 AND2X2_4920 ( .A(u3__abc_46775_n371_1), .B(u3__abc_46775_n373_1), .Y(u3__abc_46775_n374) );
  AND2X2 AND2X2_4921 ( .A(u3__abc_46775_n375), .B(u3__abc_46775_n369), .Y(u3__abc_46775_n376) );
  AND2X2 AND2X2_4922 ( .A(u3__abc_46775_n374), .B(u3__abc_46775_n368_1), .Y(u3__abc_46775_n377) );
  AND2X2 AND2X2_4923 ( .A(u3__abc_46775_n379), .B(u3__abc_46775_n364), .Y(u3__abc_46775_n380) );
  AND2X2 AND2X2_4924 ( .A(u3__abc_46775_n381_1), .B(u3__abc_46775_n378), .Y(u3__abc_46775_n382) );
  AND2X2 AND2X2_4925 ( .A(u3__abc_46775_n383), .B(u3__abc_46775_n277_1_bF_buf2), .Y(u3__abc_46775_n384) );
  AND2X2 AND2X2_4926 ( .A(u3__abc_46775_n279_bF_buf3), .B(mc_dp_od_2_), .Y(u3__abc_46775_n385) );
  AND2X2 AND2X2_4927 ( .A(\wb_data_i[27] ), .B(\wb_data_i[26] ), .Y(u3__abc_46775_n388) );
  AND2X2 AND2X2_4928 ( .A(u3__abc_46775_n389), .B(u3__abc_46775_n387), .Y(u3__abc_46775_n390_1) );
  AND2X2 AND2X2_4929 ( .A(u3__abc_46775_n392_1), .B(u3__abc_46775_n394), .Y(u3__abc_46775_n395) );
  AND2X2 AND2X2_493 ( .A(u0__abc_49347_n1847_1), .B(u0__abc_49347_n1178_1_bF_buf2), .Y(u0__abc_49347_n1848_1) );
  AND2X2 AND2X2_4930 ( .A(u3__abc_46775_n396), .B(u3__abc_46775_n390_1), .Y(u3__abc_46775_n397) );
  AND2X2 AND2X2_4931 ( .A(u3__abc_46775_n398), .B(u3__abc_46775_n399), .Y(u3__abc_46775_n400) );
  AND2X2 AND2X2_4932 ( .A(\wb_data_i[31] ), .B(\wb_data_i[30] ), .Y(u3__abc_46775_n402_1) );
  AND2X2 AND2X2_4933 ( .A(u3__abc_46775_n403), .B(u3__abc_46775_n401), .Y(u3__abc_46775_n404) );
  AND2X2 AND2X2_4934 ( .A(u3__abc_46775_n407), .B(u3__abc_46775_n409), .Y(u3__abc_46775_n410) );
  AND2X2 AND2X2_4935 ( .A(u3__abc_46775_n411_1), .B(u3__abc_46775_n405), .Y(u3__abc_46775_n412) );
  AND2X2 AND2X2_4936 ( .A(u3__abc_46775_n410), .B(u3__abc_46775_n404), .Y(u3__abc_46775_n413_1) );
  AND2X2 AND2X2_4937 ( .A(u3__abc_46775_n415), .B(u3__abc_46775_n400), .Y(u3__abc_46775_n416_1) );
  AND2X2 AND2X2_4938 ( .A(u3__abc_46775_n417), .B(u3__abc_46775_n414_1), .Y(u3__abc_46775_n418) );
  AND2X2 AND2X2_4939 ( .A(u3__abc_46775_n419_1), .B(u3__abc_46775_n277_1_bF_buf1), .Y(u3__abc_46775_n420) );
  AND2X2 AND2X2_494 ( .A(spec_req_cs_1_bF_buf5), .B(u0_tms1_27_), .Y(u0__abc_49347_n1849_1) );
  AND2X2 AND2X2_4940 ( .A(u3__abc_46775_n279_bF_buf2), .B(mc_dp_od_3_), .Y(u3__abc_46775_n421_1) );
  AND2X2 AND2X2_4941 ( .A(u3__abc_46775_n425), .B(u3__abc_46775_n423), .Y(u3_byte2_0__FF_INPUT) );
  AND2X2 AND2X2_4942 ( .A(u3__abc_46775_n428), .B(u3__abc_46775_n427), .Y(u3_byte2_1__FF_INPUT) );
  AND2X2 AND2X2_4943 ( .A(u3__abc_46775_n431), .B(u3__abc_46775_n430), .Y(u3_byte2_2__FF_INPUT) );
  AND2X2 AND2X2_4944 ( .A(u3__abc_46775_n434), .B(u3__abc_46775_n433), .Y(u3_byte2_3__FF_INPUT) );
  AND2X2 AND2X2_4945 ( .A(u3__abc_46775_n437), .B(u3__abc_46775_n436), .Y(u3_byte2_4__FF_INPUT) );
  AND2X2 AND2X2_4946 ( .A(u3__abc_46775_n440), .B(u3__abc_46775_n439), .Y(u3_byte2_5__FF_INPUT) );
  AND2X2 AND2X2_4947 ( .A(u3__abc_46775_n443), .B(u3__abc_46775_n442), .Y(u3_byte2_6__FF_INPUT) );
  AND2X2 AND2X2_4948 ( .A(u3__abc_46775_n446), .B(u3__abc_46775_n445), .Y(u3_byte2_7__FF_INPUT) );
  AND2X2 AND2X2_4949 ( .A(u3__abc_46775_n448_bF_buf3), .B(u3__abc_46775_n449), .Y(u3__abc_46775_n450) );
  AND2X2 AND2X2_495 ( .A(u0__abc_49347_n1175_bF_buf6), .B(u0__abc_49347_n1852_1), .Y(u0__abc_49347_n1853_1) );
  AND2X2 AND2X2_4950 ( .A(u3__abc_46775_n450_bF_buf3), .B(pack_le1), .Y(u3__abc_46775_n451) );
  AND2X2 AND2X2_4951 ( .A(u3__abc_46775_n448_bF_buf2), .B(csc_4_), .Y(u3__abc_46775_n452) );
  AND2X2 AND2X2_4952 ( .A(u3__abc_46775_n452_bF_buf3), .B(pack_le0), .Y(u3__abc_46775_n453) );
  AND2X2 AND2X2_4953 ( .A(u3__abc_46775_n455), .B(u3__abc_46775_n456), .Y(u3__abc_46775_n457) );
  AND2X2 AND2X2_4954 ( .A(u3__abc_46775_n458), .B(u3__abc_46775_n460), .Y(u3_byte1_0__FF_INPUT) );
  AND2X2 AND2X2_4955 ( .A(u3__abc_46775_n462), .B(u3__abc_46775_n463), .Y(u3__abc_46775_n464) );
  AND2X2 AND2X2_4956 ( .A(u3__abc_46775_n465), .B(u3__abc_46775_n466), .Y(u3_byte1_1__FF_INPUT) );
  AND2X2 AND2X2_4957 ( .A(u3__abc_46775_n468), .B(u3__abc_46775_n469), .Y(u3__abc_46775_n470) );
  AND2X2 AND2X2_4958 ( .A(u3__abc_46775_n471), .B(u3__abc_46775_n472), .Y(u3_byte1_2__FF_INPUT) );
  AND2X2 AND2X2_4959 ( .A(u3__abc_46775_n474), .B(u3__abc_46775_n475), .Y(u3__abc_46775_n476) );
  AND2X2 AND2X2_496 ( .A(u0__abc_49347_n1851_1), .B(u0__abc_49347_n1853_1), .Y(u0__abc_49347_n1854_1) );
  AND2X2 AND2X2_4960 ( .A(u3__abc_46775_n477), .B(u3__abc_46775_n478), .Y(u3_byte1_3__FF_INPUT) );
  AND2X2 AND2X2_4961 ( .A(u3__abc_46775_n480), .B(u3__abc_46775_n481), .Y(u3__abc_46775_n482) );
  AND2X2 AND2X2_4962 ( .A(u3__abc_46775_n483), .B(u3__abc_46775_n484), .Y(u3_byte1_4__FF_INPUT) );
  AND2X2 AND2X2_4963 ( .A(u3__abc_46775_n486), .B(u3__abc_46775_n487), .Y(u3__abc_46775_n488) );
  AND2X2 AND2X2_4964 ( .A(u3__abc_46775_n489), .B(u3__abc_46775_n490), .Y(u3_byte1_5__FF_INPUT) );
  AND2X2 AND2X2_4965 ( .A(u3__abc_46775_n492), .B(u3__abc_46775_n493), .Y(u3__abc_46775_n494) );
  AND2X2 AND2X2_4966 ( .A(u3__abc_46775_n495), .B(u3__abc_46775_n496), .Y(u3_byte1_6__FF_INPUT) );
  AND2X2 AND2X2_4967 ( .A(u3__abc_46775_n498), .B(u3__abc_46775_n499), .Y(u3__abc_46775_n500) );
  AND2X2 AND2X2_4968 ( .A(u3__abc_46775_n501), .B(u3__abc_46775_n502), .Y(u3_byte1_7__FF_INPUT) );
  AND2X2 AND2X2_4969 ( .A(u3__abc_46775_n506), .B(u3__abc_46775_n504), .Y(u3_byte0_0__FF_INPUT) );
  AND2X2 AND2X2_497 ( .A(u0__abc_49347_n1173), .B(cs_le_d), .Y(u0__abc_49347_n1952_1) );
  AND2X2 AND2X2_4970 ( .A(u3__abc_46775_n509), .B(u3__abc_46775_n508), .Y(u3_byte0_1__FF_INPUT) );
  AND2X2 AND2X2_4971 ( .A(u3__abc_46775_n512), .B(u3__abc_46775_n511), .Y(u3_byte0_2__FF_INPUT) );
  AND2X2 AND2X2_4972 ( .A(u3__abc_46775_n515), .B(u3__abc_46775_n514), .Y(u3_byte0_3__FF_INPUT) );
  AND2X2 AND2X2_4973 ( .A(u3__abc_46775_n518), .B(u3__abc_46775_n517), .Y(u3_byte0_4__FF_INPUT) );
  AND2X2 AND2X2_4974 ( .A(u3__abc_46775_n521), .B(u3__abc_46775_n520), .Y(u3_byte0_5__FF_INPUT) );
  AND2X2 AND2X2_4975 ( .A(u3__abc_46775_n524), .B(u3__abc_46775_n523), .Y(u3_byte0_6__FF_INPUT) );
  AND2X2 AND2X2_4976 ( .A(u3__abc_46775_n527), .B(u3__abc_46775_n526), .Y(u3_byte0_7__FF_INPUT) );
  AND2X2 AND2X2_4977 ( .A(u3__abc_46775_n529), .B(u3__abc_46775_n530), .Y(u3_mc_data_o_0__FF_INPUT) );
  AND2X2 AND2X2_4978 ( .A(u3__abc_46775_n532), .B(u3__abc_46775_n533), .Y(u3_mc_data_o_1__FF_INPUT) );
  AND2X2 AND2X2_4979 ( .A(u3__abc_46775_n535), .B(u3__abc_46775_n536), .Y(u3_mc_data_o_2__FF_INPUT) );
  AND2X2 AND2X2_498 ( .A(u0__abc_49347_n1953_1_bF_buf3), .B(sp_csc_1_), .Y(u0__abc_49347_n1978) );
  AND2X2 AND2X2_4980 ( .A(u3__abc_46775_n538), .B(u3__abc_46775_n539), .Y(u3_mc_data_o_3__FF_INPUT) );
  AND2X2 AND2X2_4981 ( .A(u3__abc_46775_n541), .B(u3__abc_46775_n542), .Y(u3_mc_data_o_4__FF_INPUT) );
  AND2X2 AND2X2_4982 ( .A(u3__abc_46775_n544), .B(u3__abc_46775_n545), .Y(u3_mc_data_o_5__FF_INPUT) );
  AND2X2 AND2X2_4983 ( .A(u3__abc_46775_n547), .B(u3__abc_46775_n548), .Y(u3_mc_data_o_6__FF_INPUT) );
  AND2X2 AND2X2_4984 ( .A(u3__abc_46775_n550), .B(u3__abc_46775_n551), .Y(u3_mc_data_o_7__FF_INPUT) );
  AND2X2 AND2X2_4985 ( .A(u3__abc_46775_n553), .B(u3__abc_46775_n554), .Y(u3_mc_data_o_8__FF_INPUT) );
  AND2X2 AND2X2_4986 ( .A(u3__abc_46775_n556), .B(u3__abc_46775_n557), .Y(u3_mc_data_o_9__FF_INPUT) );
  AND2X2 AND2X2_4987 ( .A(u3__abc_46775_n559), .B(u3__abc_46775_n560), .Y(u3_mc_data_o_10__FF_INPUT) );
  AND2X2 AND2X2_4988 ( .A(u3__abc_46775_n562), .B(u3__abc_46775_n563), .Y(u3_mc_data_o_11__FF_INPUT) );
  AND2X2 AND2X2_4989 ( .A(u3__abc_46775_n565), .B(u3__abc_46775_n566), .Y(u3_mc_data_o_12__FF_INPUT) );
  AND2X2 AND2X2_499 ( .A(spec_req_cs_5_bF_buf4), .B(u0_csc5_1_), .Y(u0__abc_49347_n1979_1) );
  AND2X2 AND2X2_4990 ( .A(u3__abc_46775_n568), .B(u3__abc_46775_n569), .Y(u3_mc_data_o_13__FF_INPUT) );
  AND2X2 AND2X2_4991 ( .A(u3__abc_46775_n571), .B(u3__abc_46775_n572), .Y(u3_mc_data_o_14__FF_INPUT) );
  AND2X2 AND2X2_4992 ( .A(u3__abc_46775_n574), .B(u3__abc_46775_n575), .Y(u3_mc_data_o_15__FF_INPUT) );
  AND2X2 AND2X2_4993 ( .A(u3__abc_46775_n577), .B(u3__abc_46775_n578), .Y(u3_mc_data_o_16__FF_INPUT) );
  AND2X2 AND2X2_4994 ( .A(u3__abc_46775_n580), .B(u3__abc_46775_n581), .Y(u3_mc_data_o_17__FF_INPUT) );
  AND2X2 AND2X2_4995 ( .A(u3__abc_46775_n583), .B(u3__abc_46775_n584), .Y(u3_mc_data_o_18__FF_INPUT) );
  AND2X2 AND2X2_4996 ( .A(u3__abc_46775_n586), .B(u3__abc_46775_n587), .Y(u3_mc_data_o_19__FF_INPUT) );
  AND2X2 AND2X2_4997 ( .A(u3__abc_46775_n589), .B(u3__abc_46775_n590), .Y(u3_mc_data_o_20__FF_INPUT) );
  AND2X2 AND2X2_4998 ( .A(u3__abc_46775_n592), .B(u3__abc_46775_n593), .Y(u3_mc_data_o_21__FF_INPUT) );
  AND2X2 AND2X2_4999 ( .A(u3__abc_46775_n595), .B(u3__abc_46775_n596), .Y(u3_mc_data_o_22__FF_INPUT) );
  AND2X2 AND2X2_5 ( .A(_abc_55805_n251), .B(_abc_55805_n252), .Y(obct_cs_1_) );
  AND2X2 AND2X2_50 ( .A(_abc_55805_n401), .B(_abc_55805_n402), .Y(csc_s_5_) );
  AND2X2 AND2X2_500 ( .A(u0__abc_49347_n1981_1), .B(u0__abc_49347_n1185_bF_buf1), .Y(u0__abc_49347_n1982) );
  AND2X2 AND2X2_5000 ( .A(u3__abc_46775_n598), .B(u3__abc_46775_n599), .Y(u3_mc_data_o_23__FF_INPUT) );
  AND2X2 AND2X2_5001 ( .A(u3__abc_46775_n601), .B(u3__abc_46775_n602), .Y(u3_mc_data_o_24__FF_INPUT) );
  AND2X2 AND2X2_5002 ( .A(u3__abc_46775_n604), .B(u3__abc_46775_n605), .Y(u3_mc_data_o_25__FF_INPUT) );
  AND2X2 AND2X2_5003 ( .A(u3__abc_46775_n607), .B(u3__abc_46775_n608), .Y(u3_mc_data_o_26__FF_INPUT) );
  AND2X2 AND2X2_5004 ( .A(u3__abc_46775_n610), .B(u3__abc_46775_n611), .Y(u3_mc_data_o_27__FF_INPUT) );
  AND2X2 AND2X2_5005 ( .A(u3__abc_46775_n613), .B(u3__abc_46775_n614), .Y(u3_mc_data_o_28__FF_INPUT) );
  AND2X2 AND2X2_5006 ( .A(u3__abc_46775_n616), .B(u3__abc_46775_n617), .Y(u3_mc_data_o_29__FF_INPUT) );
  AND2X2 AND2X2_5007 ( .A(u3__abc_46775_n619), .B(u3__abc_46775_n620), .Y(u3_mc_data_o_30__FF_INPUT) );
  AND2X2 AND2X2_5008 ( .A(u3__abc_46775_n622), .B(u3__abc_46775_n623), .Y(u3_mc_data_o_31__FF_INPUT) );
  AND2X2 AND2X2_5009 ( .A(u3__abc_46775_n627), .B(u3__abc_46775_n626), .Y(u3__abc_46775_n628) );
  AND2X2 AND2X2_501 ( .A(u0__abc_49347_n1982), .B(u0__abc_49347_n1980), .Y(u0__abc_49347_n1983_1) );
  AND2X2 AND2X2_5010 ( .A(u3__abc_46775_n629), .B(u3__abc_46775_n630), .Y(mem_dout_0_) );
  AND2X2 AND2X2_5011 ( .A(u3__abc_46775_n633), .B(u3__abc_46775_n632), .Y(u3__abc_46775_n634) );
  AND2X2 AND2X2_5012 ( .A(u3__abc_46775_n635), .B(u3__abc_46775_n636), .Y(mem_dout_1_) );
  AND2X2 AND2X2_5013 ( .A(u3__abc_46775_n639), .B(u3__abc_46775_n638), .Y(u3__abc_46775_n640) );
  AND2X2 AND2X2_5014 ( .A(u3__abc_46775_n641), .B(u3__abc_46775_n642), .Y(mem_dout_2_) );
  AND2X2 AND2X2_5015 ( .A(u3__abc_46775_n645), .B(u3__abc_46775_n644), .Y(u3__abc_46775_n646) );
  AND2X2 AND2X2_5016 ( .A(u3__abc_46775_n647), .B(u3__abc_46775_n648), .Y(mem_dout_3_) );
  AND2X2 AND2X2_5017 ( .A(u3__abc_46775_n651), .B(u3__abc_46775_n650), .Y(u3__abc_46775_n652) );
  AND2X2 AND2X2_5018 ( .A(u3__abc_46775_n653), .B(u3__abc_46775_n654), .Y(mem_dout_4_) );
  AND2X2 AND2X2_5019 ( .A(u3__abc_46775_n657), .B(u3__abc_46775_n656), .Y(u3__abc_46775_n658) );
  AND2X2 AND2X2_502 ( .A(u0__abc_49347_n1984_1), .B(u0__abc_49347_n1181_bF_buf1), .Y(u0__abc_49347_n1985) );
  AND2X2 AND2X2_5020 ( .A(u3__abc_46775_n659), .B(u3__abc_46775_n660), .Y(mem_dout_5_) );
  AND2X2 AND2X2_5021 ( .A(u3__abc_46775_n663), .B(u3__abc_46775_n662), .Y(u3__abc_46775_n664) );
  AND2X2 AND2X2_5022 ( .A(u3__abc_46775_n665), .B(u3__abc_46775_n666), .Y(mem_dout_6_) );
  AND2X2 AND2X2_5023 ( .A(u3__abc_46775_n669), .B(u3__abc_46775_n668), .Y(u3__abc_46775_n670) );
  AND2X2 AND2X2_5024 ( .A(u3__abc_46775_n671), .B(u3__abc_46775_n672), .Y(mem_dout_7_) );
  AND2X2 AND2X2_5025 ( .A(u3__abc_46775_n675), .B(u3__abc_46775_n674), .Y(u3__abc_46775_n676) );
  AND2X2 AND2X2_5026 ( .A(u3__abc_46775_n677), .B(u3__abc_46775_n678), .Y(mem_dout_8_) );
  AND2X2 AND2X2_5027 ( .A(u3__abc_46775_n681), .B(u3__abc_46775_n680), .Y(u3__abc_46775_n682) );
  AND2X2 AND2X2_5028 ( .A(u3__abc_46775_n683), .B(u3__abc_46775_n684), .Y(mem_dout_9_) );
  AND2X2 AND2X2_5029 ( .A(u3__abc_46775_n687), .B(u3__abc_46775_n686), .Y(u3__abc_46775_n688) );
  AND2X2 AND2X2_503 ( .A(spec_req_cs_4_bF_buf4), .B(u0_csc4_1_), .Y(u0__abc_49347_n1986) );
  AND2X2 AND2X2_5030 ( .A(u3__abc_46775_n689), .B(u3__abc_46775_n690), .Y(mem_dout_10_) );
  AND2X2 AND2X2_5031 ( .A(u3__abc_46775_n693), .B(u3__abc_46775_n692), .Y(u3__abc_46775_n694) );
  AND2X2 AND2X2_5032 ( .A(u3__abc_46775_n695), .B(u3__abc_46775_n696), .Y(mem_dout_11_) );
  AND2X2 AND2X2_5033 ( .A(u3__abc_46775_n699), .B(u3__abc_46775_n698), .Y(u3__abc_46775_n700) );
  AND2X2 AND2X2_5034 ( .A(u3__abc_46775_n701), .B(u3__abc_46775_n702), .Y(mem_dout_12_) );
  AND2X2 AND2X2_5035 ( .A(u3__abc_46775_n705), .B(u3__abc_46775_n704), .Y(u3__abc_46775_n706) );
  AND2X2 AND2X2_5036 ( .A(u3__abc_46775_n707), .B(u3__abc_46775_n708), .Y(mem_dout_13_) );
  AND2X2 AND2X2_5037 ( .A(u3__abc_46775_n711), .B(u3__abc_46775_n710), .Y(u3__abc_46775_n712) );
  AND2X2 AND2X2_5038 ( .A(u3__abc_46775_n713), .B(u3__abc_46775_n714), .Y(mem_dout_14_) );
  AND2X2 AND2X2_5039 ( .A(u3__abc_46775_n717), .B(u3__abc_46775_n716), .Y(u3__abc_46775_n718) );
  AND2X2 AND2X2_504 ( .A(u0__abc_49347_n1987), .B(u0__abc_49347_n1180_1_bF_buf1), .Y(u0__abc_49347_n1988) );
  AND2X2 AND2X2_5040 ( .A(u3__abc_46775_n719), .B(u3__abc_46775_n720), .Y(mem_dout_15_) );
  AND2X2 AND2X2_5041 ( .A(u3__abc_46775_n452_bF_buf2), .B(mc_data_ir_0_), .Y(u3__abc_46775_n722) );
  AND2X2 AND2X2_5042 ( .A(csc_5_bF_buf0), .B(mc_data_ir_16_), .Y(u3__abc_46775_n723) );
  AND2X2 AND2X2_5043 ( .A(u3__abc_46775_n450_bF_buf2), .B(u3_byte2_0_), .Y(u3__abc_46775_n725) );
  AND2X2 AND2X2_5044 ( .A(u3__abc_46775_n727), .B(u3__abc_46775_n728), .Y(mem_dout_16_) );
  AND2X2 AND2X2_5045 ( .A(u3__abc_46775_n452_bF_buf1), .B(mc_data_ir_1_), .Y(u3__abc_46775_n730) );
  AND2X2 AND2X2_5046 ( .A(csc_5_bF_buf4), .B(mc_data_ir_17_), .Y(u3__abc_46775_n731) );
  AND2X2 AND2X2_5047 ( .A(u3__abc_46775_n450_bF_buf1), .B(u3_byte2_1_), .Y(u3__abc_46775_n733) );
  AND2X2 AND2X2_5048 ( .A(u3__abc_46775_n735), .B(u3__abc_46775_n736), .Y(mem_dout_17_) );
  AND2X2 AND2X2_5049 ( .A(u3__abc_46775_n452_bF_buf0), .B(mc_data_ir_2_), .Y(u3__abc_46775_n738) );
  AND2X2 AND2X2_505 ( .A(spec_req_cs_3_bF_buf4), .B(u0_csc3_1_), .Y(u0__abc_49347_n1989) );
  AND2X2 AND2X2_5050 ( .A(csc_5_bF_buf3), .B(mc_data_ir_18_), .Y(u3__abc_46775_n739) );
  AND2X2 AND2X2_5051 ( .A(u3__abc_46775_n450_bF_buf0), .B(u3_byte2_2_), .Y(u3__abc_46775_n741) );
  AND2X2 AND2X2_5052 ( .A(u3__abc_46775_n743), .B(u3__abc_46775_n744), .Y(mem_dout_18_) );
  AND2X2 AND2X2_5053 ( .A(u3__abc_46775_n452_bF_buf3), .B(mc_data_ir_3_), .Y(u3__abc_46775_n746) );
  AND2X2 AND2X2_5054 ( .A(csc_5_bF_buf2), .B(mc_data_ir_19_), .Y(u3__abc_46775_n747) );
  AND2X2 AND2X2_5055 ( .A(u3__abc_46775_n450_bF_buf3), .B(u3_byte2_3_), .Y(u3__abc_46775_n749) );
  AND2X2 AND2X2_5056 ( .A(u3__abc_46775_n751), .B(u3__abc_46775_n752), .Y(mem_dout_19_) );
  AND2X2 AND2X2_5057 ( .A(u3__abc_46775_n452_bF_buf2), .B(mc_data_ir_4_), .Y(u3__abc_46775_n754) );
  AND2X2 AND2X2_5058 ( .A(csc_5_bF_buf1), .B(mc_data_ir_20_), .Y(u3__abc_46775_n755) );
  AND2X2 AND2X2_5059 ( .A(u3__abc_46775_n450_bF_buf2), .B(u3_byte2_4_), .Y(u3__abc_46775_n757) );
  AND2X2 AND2X2_506 ( .A(u0__abc_49347_n1990), .B(u0__abc_49347_n1179_bF_buf1), .Y(u0__abc_49347_n1991) );
  AND2X2 AND2X2_5060 ( .A(u3__abc_46775_n759), .B(u3__abc_46775_n760), .Y(mem_dout_20_) );
  AND2X2 AND2X2_5061 ( .A(u3__abc_46775_n452_bF_buf1), .B(mc_data_ir_5_), .Y(u3__abc_46775_n762) );
  AND2X2 AND2X2_5062 ( .A(csc_5_bF_buf0), .B(mc_data_ir_21_), .Y(u3__abc_46775_n763) );
  AND2X2 AND2X2_5063 ( .A(u3__abc_46775_n450_bF_buf1), .B(u3_byte2_5_), .Y(u3__abc_46775_n765) );
  AND2X2 AND2X2_5064 ( .A(u3__abc_46775_n767), .B(u3__abc_46775_n768), .Y(mem_dout_21_) );
  AND2X2 AND2X2_5065 ( .A(u3__abc_46775_n452_bF_buf0), .B(mc_data_ir_6_), .Y(u3__abc_46775_n770) );
  AND2X2 AND2X2_5066 ( .A(csc_5_bF_buf4), .B(mc_data_ir_22_), .Y(u3__abc_46775_n771) );
  AND2X2 AND2X2_5067 ( .A(u3__abc_46775_n450_bF_buf0), .B(u3_byte2_6_), .Y(u3__abc_46775_n773) );
  AND2X2 AND2X2_5068 ( .A(u3__abc_46775_n775), .B(u3__abc_46775_n776), .Y(mem_dout_22_) );
  AND2X2 AND2X2_5069 ( .A(u3__abc_46775_n452_bF_buf3), .B(mc_data_ir_7_), .Y(u3__abc_46775_n778) );
  AND2X2 AND2X2_507 ( .A(spec_req_cs_2_bF_buf4), .B(u0_csc2_1_), .Y(u0__abc_49347_n1992) );
  AND2X2 AND2X2_5070 ( .A(csc_5_bF_buf3), .B(mc_data_ir_23_), .Y(u3__abc_46775_n779) );
  AND2X2 AND2X2_5071 ( .A(u3__abc_46775_n450_bF_buf3), .B(u3_byte2_7_), .Y(u3__abc_46775_n781) );
  AND2X2 AND2X2_5072 ( .A(u3__abc_46775_n783), .B(u3__abc_46775_n784), .Y(mem_dout_23_) );
  AND2X2 AND2X2_5073 ( .A(u3__abc_46775_n452_bF_buf2), .B(mc_data_ir_8_), .Y(u3__abc_46775_n786) );
  AND2X2 AND2X2_5074 ( .A(csc_5_bF_buf2), .B(mc_data_ir_24_), .Y(u3__abc_46775_n787) );
  AND2X2 AND2X2_5075 ( .A(u3__abc_46775_n450_bF_buf2), .B(mc_data_ir_0_), .Y(u3__abc_46775_n789) );
  AND2X2 AND2X2_5076 ( .A(u3__abc_46775_n791), .B(u3__abc_46775_n792), .Y(mem_dout_24_) );
  AND2X2 AND2X2_5077 ( .A(u3__abc_46775_n452_bF_buf1), .B(mc_data_ir_9_), .Y(u3__abc_46775_n794) );
  AND2X2 AND2X2_5078 ( .A(csc_5_bF_buf1), .B(mc_data_ir_25_), .Y(u3__abc_46775_n795) );
  AND2X2 AND2X2_5079 ( .A(u3__abc_46775_n450_bF_buf1), .B(mc_data_ir_1_), .Y(u3__abc_46775_n797) );
  AND2X2 AND2X2_508 ( .A(u0__abc_49347_n1993), .B(u0__abc_49347_n1178_1_bF_buf1), .Y(u0__abc_49347_n1994) );
  AND2X2 AND2X2_5080 ( .A(u3__abc_46775_n799), .B(u3__abc_46775_n800), .Y(mem_dout_25_) );
  AND2X2 AND2X2_5081 ( .A(u3__abc_46775_n452_bF_buf0), .B(mc_data_ir_10_), .Y(u3__abc_46775_n802) );
  AND2X2 AND2X2_5082 ( .A(csc_5_bF_buf0), .B(mc_data_ir_26_), .Y(u3__abc_46775_n803) );
  AND2X2 AND2X2_5083 ( .A(u3__abc_46775_n450_bF_buf0), .B(mc_data_ir_2_), .Y(u3__abc_46775_n805) );
  AND2X2 AND2X2_5084 ( .A(u3__abc_46775_n807), .B(u3__abc_46775_n808), .Y(mem_dout_26_) );
  AND2X2 AND2X2_5085 ( .A(u3__abc_46775_n452_bF_buf3), .B(mc_data_ir_11_), .Y(u3__abc_46775_n810) );
  AND2X2 AND2X2_5086 ( .A(csc_5_bF_buf4), .B(mc_data_ir_27_), .Y(u3__abc_46775_n811) );
  AND2X2 AND2X2_5087 ( .A(u3__abc_46775_n450_bF_buf3), .B(mc_data_ir_3_), .Y(u3__abc_46775_n813) );
  AND2X2 AND2X2_5088 ( .A(u3__abc_46775_n815), .B(u3__abc_46775_n816), .Y(mem_dout_27_) );
  AND2X2 AND2X2_5089 ( .A(u3__abc_46775_n452_bF_buf2), .B(mc_data_ir_12_), .Y(u3__abc_46775_n818) );
  AND2X2 AND2X2_509 ( .A(spec_req_cs_1_bF_buf4), .B(u0_csc1_1_), .Y(u0__abc_49347_n1995) );
  AND2X2 AND2X2_5090 ( .A(csc_5_bF_buf3), .B(mc_data_ir_28_), .Y(u3__abc_46775_n819) );
  AND2X2 AND2X2_5091 ( .A(u3__abc_46775_n450_bF_buf2), .B(mc_data_ir_4_), .Y(u3__abc_46775_n821) );
  AND2X2 AND2X2_5092 ( .A(u3__abc_46775_n823), .B(u3__abc_46775_n824), .Y(mem_dout_28_) );
  AND2X2 AND2X2_5093 ( .A(u3__abc_46775_n452_bF_buf1), .B(mc_data_ir_13_), .Y(u3__abc_46775_n826) );
  AND2X2 AND2X2_5094 ( .A(csc_5_bF_buf2), .B(mc_data_ir_29_), .Y(u3__abc_46775_n827) );
  AND2X2 AND2X2_5095 ( .A(u3__abc_46775_n450_bF_buf1), .B(mc_data_ir_5_), .Y(u3__abc_46775_n829) );
  AND2X2 AND2X2_5096 ( .A(u3__abc_46775_n831), .B(u3__abc_46775_n832), .Y(mem_dout_29_) );
  AND2X2 AND2X2_5097 ( .A(u3__abc_46775_n452_bF_buf0), .B(mc_data_ir_14_), .Y(u3__abc_46775_n834) );
  AND2X2 AND2X2_5098 ( .A(csc_5_bF_buf1), .B(mc_data_ir_30_), .Y(u3__abc_46775_n835) );
  AND2X2 AND2X2_5099 ( .A(u3__abc_46775_n450_bF_buf0), .B(mc_data_ir_6_), .Y(u3__abc_46775_n837) );
  AND2X2 AND2X2_51 ( .A(_abc_55805_n404), .B(_abc_55805_n405), .Y(csc_s_6_) );
  AND2X2 AND2X2_510 ( .A(u0__abc_49347_n1952_1_bF_buf2), .B(u0__abc_49347_n1998), .Y(u0__abc_49347_n1999) );
  AND2X2 AND2X2_5100 ( .A(u3__abc_46775_n839), .B(u3__abc_46775_n840), .Y(mem_dout_30_) );
  AND2X2 AND2X2_5101 ( .A(u3__abc_46775_n452_bF_buf3), .B(mc_data_ir_15_), .Y(u3__abc_46775_n842) );
  AND2X2 AND2X2_5102 ( .A(csc_5_bF_buf0), .B(mc_data_ir_31_), .Y(u3__abc_46775_n843) );
  AND2X2 AND2X2_5103 ( .A(u3__abc_46775_n450_bF_buf3), .B(mc_data_ir_7_), .Y(u3__abc_46775_n845) );
  AND2X2 AND2X2_5104 ( .A(u3__abc_46775_n847), .B(u3__abc_46775_n848), .Y(mem_dout_31_) );
  AND2X2 AND2X2_5105 ( .A(wb_stb_i_bF_buf1), .B(wb_we_i), .Y(u3__abc_46775_n851) );
  AND2X2 AND2X2_5106 ( .A(mem_ack_r), .B(u3_wb_read_go), .Y(u3_re) );
  AND2X2 AND2X2_5107 ( .A(u3_rd_fifo_out_14_), .B(u3_rd_fifo_out_15_), .Y(u3__abc_46775_n855) );
  AND2X2 AND2X2_5108 ( .A(u3__abc_46775_n856), .B(u3__abc_46775_n854), .Y(u3__abc_46775_n857) );
  AND2X2 AND2X2_5109 ( .A(u3__abc_46775_n860), .B(u3_rd_fifo_out_8_), .Y(u3__abc_46775_n861) );
  AND2X2 AND2X2_511 ( .A(u0__abc_49347_n1997), .B(u0__abc_49347_n1999), .Y(u0__abc_49347_n2000) );
  AND2X2 AND2X2_5110 ( .A(u3__abc_46775_n862), .B(u3_rd_fifo_out_9_), .Y(u3__abc_46775_n863) );
  AND2X2 AND2X2_5111 ( .A(u3__abc_46775_n866), .B(u3__abc_46775_n867), .Y(u3__abc_46775_n868) );
  AND2X2 AND2X2_5112 ( .A(u3__abc_46775_n865), .B(u3__abc_46775_n869), .Y(u3__abc_46775_n870) );
  AND2X2 AND2X2_5113 ( .A(u3__abc_46775_n873), .B(u3__abc_46775_n872), .Y(u3__abc_46775_n874) );
  AND2X2 AND2X2_5114 ( .A(u3__abc_46775_n871), .B(u3__abc_46775_n875), .Y(u3__abc_46775_n876) );
  AND2X2 AND2X2_5115 ( .A(u3_rd_fifo_out_12_), .B(u3_rd_fifo_out_13_), .Y(u3__abc_46775_n879) );
  AND2X2 AND2X2_5116 ( .A(u3__abc_46775_n880), .B(u3__abc_46775_n878), .Y(u3__abc_46775_n881) );
  AND2X2 AND2X2_5117 ( .A(u3__abc_46775_n883), .B(u3_rd_fifo_out_10_), .Y(u3__abc_46775_n884) );
  AND2X2 AND2X2_5118 ( .A(u3__abc_46775_n885), .B(u3__abc_46775_n886), .Y(u3__abc_46775_n887) );
  AND2X2 AND2X2_5119 ( .A(u3__abc_46775_n888), .B(u3__abc_46775_n882), .Y(u3__abc_46775_n889) );
  AND2X2 AND2X2_512 ( .A(u0__abc_49347_n1953_1_bF_buf2), .B(sp_csc_2_), .Y(u0__abc_49347_n2002) );
  AND2X2 AND2X2_5120 ( .A(u3__abc_46775_n887), .B(u3__abc_46775_n881), .Y(u3__abc_46775_n890) );
  AND2X2 AND2X2_5121 ( .A(u3__abc_46775_n894), .B(\wb_sel_i[1] ), .Y(u3__abc_46775_n895) );
  AND2X2 AND2X2_5122 ( .A(u3__abc_46775_n895), .B(u3__abc_46775_n893), .Y(u3__abc_46775_n896) );
  AND2X2 AND2X2_5123 ( .A(u3_rd_fifo_out_22_), .B(u3_rd_fifo_out_23_), .Y(u3__abc_46775_n898) );
  AND2X2 AND2X2_5124 ( .A(u3__abc_46775_n899), .B(u3__abc_46775_n897), .Y(u3__abc_46775_n900) );
  AND2X2 AND2X2_5125 ( .A(u3_rd_fifo_out_16_), .B(u3_rd_fifo_out_17_), .Y(u3__abc_46775_n904) );
  AND2X2 AND2X2_5126 ( .A(u3__abc_46775_n905), .B(u3__abc_46775_n903), .Y(u3__abc_46775_n906) );
  AND2X2 AND2X2_5127 ( .A(u3__abc_46775_n908), .B(u3__abc_46775_n909), .Y(u3__abc_46775_n910) );
  AND2X2 AND2X2_5128 ( .A(u3__abc_46775_n912), .B(u3__abc_46775_n907), .Y(u3__abc_46775_n913) );
  AND2X2 AND2X2_5129 ( .A(u3__abc_46775_n911), .B(u3_rd_fifo_out_34_), .Y(u3__abc_46775_n915) );
  AND2X2 AND2X2_513 ( .A(spec_req_cs_5_bF_buf3), .B(u0_csc5_2_), .Y(u0__abc_49347_n2003) );
  AND2X2 AND2X2_5130 ( .A(u3__abc_46775_n906), .B(u3__abc_46775_n902), .Y(u3__abc_46775_n916) );
  AND2X2 AND2X2_5131 ( .A(u3__abc_46775_n914), .B(u3__abc_46775_n918), .Y(u3__abc_46775_n919) );
  AND2X2 AND2X2_5132 ( .A(u3_rd_fifo_out_20_), .B(u3_rd_fifo_out_21_), .Y(u3__abc_46775_n922) );
  AND2X2 AND2X2_5133 ( .A(u3__abc_46775_n923), .B(u3__abc_46775_n921), .Y(u3__abc_46775_n924) );
  AND2X2 AND2X2_5134 ( .A(u3__abc_46775_n926), .B(u3_rd_fifo_out_18_), .Y(u3__abc_46775_n927) );
  AND2X2 AND2X2_5135 ( .A(u3__abc_46775_n928), .B(u3__abc_46775_n929), .Y(u3__abc_46775_n930) );
  AND2X2 AND2X2_5136 ( .A(u3__abc_46775_n931), .B(u3__abc_46775_n925), .Y(u3__abc_46775_n932) );
  AND2X2 AND2X2_5137 ( .A(u3__abc_46775_n930), .B(u3__abc_46775_n924), .Y(u3__abc_46775_n933) );
  AND2X2 AND2X2_5138 ( .A(u3__abc_46775_n937), .B(\wb_sel_i[2] ), .Y(u3__abc_46775_n938) );
  AND2X2 AND2X2_5139 ( .A(u3__abc_46775_n938), .B(u3__abc_46775_n936), .Y(u3__abc_46775_n939) );
  AND2X2 AND2X2_514 ( .A(u0__abc_49347_n2005), .B(u0__abc_49347_n1185_bF_buf0), .Y(u0__abc_49347_n2006) );
  AND2X2 AND2X2_5140 ( .A(u3_rd_fifo_out_6_), .B(u3_rd_fifo_out_7_), .Y(u3__abc_46775_n942) );
  AND2X2 AND2X2_5141 ( .A(u3__abc_46775_n943), .B(u3__abc_46775_n941), .Y(u3__abc_46775_n944) );
  AND2X2 AND2X2_5142 ( .A(u3_rd_fifo_out_0_), .B(u3_rd_fifo_out_1_), .Y(u3__abc_46775_n948) );
  AND2X2 AND2X2_5143 ( .A(u3__abc_46775_n949), .B(u3__abc_46775_n947), .Y(u3__abc_46775_n950) );
  AND2X2 AND2X2_5144 ( .A(u3__abc_46775_n952), .B(u3__abc_46775_n953), .Y(u3__abc_46775_n954) );
  AND2X2 AND2X2_5145 ( .A(u3__abc_46775_n956), .B(u3__abc_46775_n951), .Y(u3__abc_46775_n957) );
  AND2X2 AND2X2_5146 ( .A(u3__abc_46775_n955), .B(u3_rd_fifo_out_32_), .Y(u3__abc_46775_n959) );
  AND2X2 AND2X2_5147 ( .A(u3__abc_46775_n950), .B(u3__abc_46775_n946), .Y(u3__abc_46775_n960) );
  AND2X2 AND2X2_5148 ( .A(u3__abc_46775_n958), .B(u3__abc_46775_n962), .Y(u3__abc_46775_n963) );
  AND2X2 AND2X2_5149 ( .A(u3_rd_fifo_out_4_), .B(u3_rd_fifo_out_5_), .Y(u3__abc_46775_n966) );
  AND2X2 AND2X2_515 ( .A(u0__abc_49347_n2006), .B(u0__abc_49347_n2004), .Y(u0__abc_49347_n2007) );
  AND2X2 AND2X2_5150 ( .A(u3__abc_46775_n967), .B(u3__abc_46775_n965), .Y(u3__abc_46775_n968) );
  AND2X2 AND2X2_5151 ( .A(u3__abc_46775_n970), .B(u3_rd_fifo_out_2_), .Y(u3__abc_46775_n971) );
  AND2X2 AND2X2_5152 ( .A(u3__abc_46775_n972), .B(u3__abc_46775_n973), .Y(u3__abc_46775_n974) );
  AND2X2 AND2X2_5153 ( .A(u3__abc_46775_n975), .B(u3__abc_46775_n969), .Y(u3__abc_46775_n976) );
  AND2X2 AND2X2_5154 ( .A(u3__abc_46775_n974), .B(u3__abc_46775_n968), .Y(u3__abc_46775_n977) );
  AND2X2 AND2X2_5155 ( .A(u3__abc_46775_n981), .B(\wb_sel_i[0] ), .Y(u3__abc_46775_n982) );
  AND2X2 AND2X2_5156 ( .A(u3__abc_46775_n982), .B(u3__abc_46775_n980), .Y(u3__abc_46775_n983) );
  AND2X2 AND2X2_5157 ( .A(u3_rd_fifo_out_30_), .B(u3_rd_fifo_out_31_), .Y(u3__abc_46775_n985) );
  AND2X2 AND2X2_5158 ( .A(u3__abc_46775_n986), .B(u3__abc_46775_n984), .Y(u3__abc_46775_n987) );
  AND2X2 AND2X2_5159 ( .A(u3_rd_fifo_out_24_), .B(u3_rd_fifo_out_25_), .Y(u3__abc_46775_n991) );
  AND2X2 AND2X2_516 ( .A(u0__abc_49347_n2008), .B(u0__abc_49347_n1181_bF_buf0), .Y(u0__abc_49347_n2009) );
  AND2X2 AND2X2_5160 ( .A(u3__abc_46775_n992), .B(u3__abc_46775_n990), .Y(u3__abc_46775_n993) );
  AND2X2 AND2X2_5161 ( .A(u3__abc_46775_n996), .B(u3__abc_46775_n998), .Y(u3__abc_46775_n999) );
  AND2X2 AND2X2_5162 ( .A(u3__abc_46775_n1000), .B(u3__abc_46775_n994), .Y(u3__abc_46775_n1001) );
  AND2X2 AND2X2_5163 ( .A(u3__abc_46775_n999), .B(u3_rd_fifo_out_35_), .Y(u3__abc_46775_n1003) );
  AND2X2 AND2X2_5164 ( .A(u3__abc_46775_n993), .B(u3__abc_46775_n989), .Y(u3__abc_46775_n1004) );
  AND2X2 AND2X2_5165 ( .A(u3__abc_46775_n1002), .B(u3__abc_46775_n1006), .Y(u3__abc_46775_n1007) );
  AND2X2 AND2X2_5166 ( .A(u3_rd_fifo_out_28_), .B(u3_rd_fifo_out_29_), .Y(u3__abc_46775_n1010) );
  AND2X2 AND2X2_5167 ( .A(u3__abc_46775_n1011), .B(u3__abc_46775_n1009), .Y(u3__abc_46775_n1012) );
  AND2X2 AND2X2_5168 ( .A(u3__abc_46775_n1014), .B(u3_rd_fifo_out_26_), .Y(u3__abc_46775_n1015) );
  AND2X2 AND2X2_5169 ( .A(u3__abc_46775_n1016), .B(u3__abc_46775_n1017), .Y(u3__abc_46775_n1018) );
  AND2X2 AND2X2_517 ( .A(spec_req_cs_4_bF_buf3), .B(u0_csc4_2_), .Y(u0__abc_49347_n2010) );
  AND2X2 AND2X2_5170 ( .A(u3__abc_46775_n1019), .B(u3__abc_46775_n1013), .Y(u3__abc_46775_n1020) );
  AND2X2 AND2X2_5171 ( .A(u3__abc_46775_n1018), .B(u3__abc_46775_n1012), .Y(u3__abc_46775_n1021) );
  AND2X2 AND2X2_5172 ( .A(u3__abc_46775_n1025), .B(\wb_sel_i[3] ), .Y(u3__abc_46775_n1026) );
  AND2X2 AND2X2_5173 ( .A(u3__abc_46775_n1026), .B(u3__abc_46775_n1024), .Y(u3__abc_46775_n1027) );
  AND2X2 AND2X2_5174 ( .A(u3__abc_46775_n1030), .B(mem_ack), .Y(u3__abc_46775_n1031) );
  AND2X2 AND2X2_5175 ( .A(u3__abc_46775_n1031), .B(u3_pen), .Y(u3__abc_46775_n1032) );
  AND2X2 AND2X2_5176 ( .A(u3__abc_46775_n1029), .B(u3__abc_46775_n1032), .Y(par_err) );
  AND2X2 AND2X2_5177 ( .A(dv), .B(u3_u0_wr_adr_3_), .Y(u3_u0__abc_48231_n382) );
  AND2X2 AND2X2_5178 ( .A(u3_u0__abc_48231_n382_bF_buf6), .B(u3_u0__abc_48231_n384_1), .Y(u3_u0__abc_48231_n385) );
  AND2X2 AND2X2_5179 ( .A(u3_u0__abc_48231_n386), .B(u3_u0__abc_48231_n383), .Y(u3_u0_r3_0__FF_INPUT) );
  AND2X2 AND2X2_518 ( .A(u0__abc_49347_n2011), .B(u0__abc_49347_n1180_1_bF_buf0), .Y(u0__abc_49347_n2012) );
  AND2X2 AND2X2_5180 ( .A(u3_u0__abc_48231_n382_bF_buf4), .B(u3_u0__abc_48231_n389), .Y(u3_u0__abc_48231_n390) );
  AND2X2 AND2X2_5181 ( .A(u3_u0__abc_48231_n391), .B(u3_u0__abc_48231_n388_1), .Y(u3_u0_r3_1__FF_INPUT) );
  AND2X2 AND2X2_5182 ( .A(u3_u0__abc_48231_n382_bF_buf2), .B(u3_u0__abc_48231_n394), .Y(u3_u0__abc_48231_n395) );
  AND2X2 AND2X2_5183 ( .A(u3_u0__abc_48231_n396_1), .B(u3_u0__abc_48231_n393), .Y(u3_u0_r3_2__FF_INPUT) );
  AND2X2 AND2X2_5184 ( .A(u3_u0__abc_48231_n382_bF_buf0), .B(u3_u0__abc_48231_n399), .Y(u3_u0__abc_48231_n400_1) );
  AND2X2 AND2X2_5185 ( .A(u3_u0__abc_48231_n401), .B(u3_u0__abc_48231_n398), .Y(u3_u0_r3_3__FF_INPUT) );
  AND2X2 AND2X2_5186 ( .A(u3_u0__abc_48231_n382_bF_buf6), .B(u3_u0__abc_48231_n404_1), .Y(u3_u0__abc_48231_n405) );
  AND2X2 AND2X2_5187 ( .A(u3_u0__abc_48231_n406), .B(u3_u0__abc_48231_n403), .Y(u3_u0_r3_4__FF_INPUT) );
  AND2X2 AND2X2_5188 ( .A(u3_u0__abc_48231_n382_bF_buf4), .B(u3_u0__abc_48231_n409), .Y(u3_u0__abc_48231_n410) );
  AND2X2 AND2X2_5189 ( .A(u3_u0__abc_48231_n411), .B(u3_u0__abc_48231_n408_1), .Y(u3_u0_r3_5__FF_INPUT) );
  AND2X2 AND2X2_519 ( .A(spec_req_cs_3_bF_buf3), .B(u0_csc3_2_), .Y(u0__abc_49347_n2013) );
  AND2X2 AND2X2_5190 ( .A(u3_u0__abc_48231_n382_bF_buf2), .B(u3_u0__abc_48231_n414), .Y(u3_u0__abc_48231_n415) );
  AND2X2 AND2X2_5191 ( .A(u3_u0__abc_48231_n416_1), .B(u3_u0__abc_48231_n413), .Y(u3_u0_r3_6__FF_INPUT) );
  AND2X2 AND2X2_5192 ( .A(u3_u0__abc_48231_n382_bF_buf0), .B(u3_u0__abc_48231_n419), .Y(u3_u0__abc_48231_n420_1) );
  AND2X2 AND2X2_5193 ( .A(u3_u0__abc_48231_n421), .B(u3_u0__abc_48231_n418), .Y(u3_u0_r3_7__FF_INPUT) );
  AND2X2 AND2X2_5194 ( .A(u3_u0__abc_48231_n382_bF_buf6), .B(u3_u0__abc_48231_n424_1), .Y(u3_u0__abc_48231_n425) );
  AND2X2 AND2X2_5195 ( .A(u3_u0__abc_48231_n426), .B(u3_u0__abc_48231_n423), .Y(u3_u0_r3_8__FF_INPUT) );
  AND2X2 AND2X2_5196 ( .A(u3_u0__abc_48231_n382_bF_buf4), .B(u3_u0__abc_48231_n429), .Y(u3_u0__abc_48231_n430) );
  AND2X2 AND2X2_5197 ( .A(u3_u0__abc_48231_n431), .B(u3_u0__abc_48231_n428_1), .Y(u3_u0_r3_9__FF_INPUT) );
  AND2X2 AND2X2_5198 ( .A(u3_u0__abc_48231_n382_bF_buf2), .B(u3_u0__abc_48231_n434), .Y(u3_u0__abc_48231_n435) );
  AND2X2 AND2X2_5199 ( .A(u3_u0__abc_48231_n436_1), .B(u3_u0__abc_48231_n433), .Y(u3_u0_r3_10__FF_INPUT) );
  AND2X2 AND2X2_52 ( .A(_abc_55805_n407), .B(_abc_55805_n408), .Y(csc_s_7_) );
  AND2X2 AND2X2_520 ( .A(u0__abc_49347_n2014), .B(u0__abc_49347_n1179_bF_buf0), .Y(u0__abc_49347_n2015) );
  AND2X2 AND2X2_5200 ( .A(u3_u0__abc_48231_n382_bF_buf0), .B(u3_u0__abc_48231_n439), .Y(u3_u0__abc_48231_n440_1) );
  AND2X2 AND2X2_5201 ( .A(u3_u0__abc_48231_n441), .B(u3_u0__abc_48231_n438), .Y(u3_u0_r3_11__FF_INPUT) );
  AND2X2 AND2X2_5202 ( .A(u3_u0__abc_48231_n382_bF_buf6), .B(u3_u0__abc_48231_n444_1), .Y(u3_u0__abc_48231_n445) );
  AND2X2 AND2X2_5203 ( .A(u3_u0__abc_48231_n446), .B(u3_u0__abc_48231_n443), .Y(u3_u0_r3_12__FF_INPUT) );
  AND2X2 AND2X2_5204 ( .A(u3_u0__abc_48231_n382_bF_buf4), .B(u3_u0__abc_48231_n449), .Y(u3_u0__abc_48231_n450) );
  AND2X2 AND2X2_5205 ( .A(u3_u0__abc_48231_n451), .B(u3_u0__abc_48231_n448_1), .Y(u3_u0_r3_13__FF_INPUT) );
  AND2X2 AND2X2_5206 ( .A(u3_u0__abc_48231_n382_bF_buf2), .B(u3_u0__abc_48231_n454), .Y(u3_u0__abc_48231_n455) );
  AND2X2 AND2X2_5207 ( .A(u3_u0__abc_48231_n456_1), .B(u3_u0__abc_48231_n453), .Y(u3_u0_r3_14__FF_INPUT) );
  AND2X2 AND2X2_5208 ( .A(u3_u0__abc_48231_n382_bF_buf0), .B(u3_u0__abc_48231_n459), .Y(u3_u0__abc_48231_n460_1) );
  AND2X2 AND2X2_5209 ( .A(u3_u0__abc_48231_n461), .B(u3_u0__abc_48231_n458), .Y(u3_u0_r3_15__FF_INPUT) );
  AND2X2 AND2X2_521 ( .A(spec_req_cs_2_bF_buf3), .B(u0_csc2_2_), .Y(u0__abc_49347_n2016) );
  AND2X2 AND2X2_5210 ( .A(u3_u0__abc_48231_n382_bF_buf6), .B(u3_u0__abc_48231_n464_1), .Y(u3_u0__abc_48231_n465) );
  AND2X2 AND2X2_5211 ( .A(u3_u0__abc_48231_n466), .B(u3_u0__abc_48231_n463), .Y(u3_u0_r3_16__FF_INPUT) );
  AND2X2 AND2X2_5212 ( .A(u3_u0__abc_48231_n382_bF_buf4), .B(u3_u0__abc_48231_n469), .Y(u3_u0__abc_48231_n470) );
  AND2X2 AND2X2_5213 ( .A(u3_u0__abc_48231_n471), .B(u3_u0__abc_48231_n468_1), .Y(u3_u0_r3_17__FF_INPUT) );
  AND2X2 AND2X2_5214 ( .A(u3_u0__abc_48231_n382_bF_buf2), .B(u3_u0__abc_48231_n474), .Y(u3_u0__abc_48231_n475) );
  AND2X2 AND2X2_5215 ( .A(u3_u0__abc_48231_n476_1), .B(u3_u0__abc_48231_n473), .Y(u3_u0_r3_18__FF_INPUT) );
  AND2X2 AND2X2_5216 ( .A(u3_u0__abc_48231_n382_bF_buf0), .B(u3_u0__abc_48231_n479), .Y(u3_u0__abc_48231_n480_1) );
  AND2X2 AND2X2_5217 ( .A(u3_u0__abc_48231_n481), .B(u3_u0__abc_48231_n478), .Y(u3_u0_r3_19__FF_INPUT) );
  AND2X2 AND2X2_5218 ( .A(u3_u0__abc_48231_n382_bF_buf6), .B(u3_u0__abc_48231_n484_1), .Y(u3_u0__abc_48231_n485) );
  AND2X2 AND2X2_5219 ( .A(u3_u0__abc_48231_n486), .B(u3_u0__abc_48231_n483), .Y(u3_u0_r3_20__FF_INPUT) );
  AND2X2 AND2X2_522 ( .A(u0__abc_49347_n2017), .B(u0__abc_49347_n1178_1_bF_buf0), .Y(u0__abc_49347_n2018) );
  AND2X2 AND2X2_5220 ( .A(u3_u0__abc_48231_n382_bF_buf4), .B(u3_u0__abc_48231_n489), .Y(u3_u0__abc_48231_n490) );
  AND2X2 AND2X2_5221 ( .A(u3_u0__abc_48231_n491), .B(u3_u0__abc_48231_n488_1), .Y(u3_u0_r3_21__FF_INPUT) );
  AND2X2 AND2X2_5222 ( .A(u3_u0__abc_48231_n382_bF_buf2), .B(u3_u0__abc_48231_n494), .Y(u3_u0__abc_48231_n495) );
  AND2X2 AND2X2_5223 ( .A(u3_u0__abc_48231_n496_1), .B(u3_u0__abc_48231_n493), .Y(u3_u0_r3_22__FF_INPUT) );
  AND2X2 AND2X2_5224 ( .A(u3_u0__abc_48231_n382_bF_buf0), .B(u3_u0__abc_48231_n499), .Y(u3_u0__abc_48231_n500_1) );
  AND2X2 AND2X2_5225 ( .A(u3_u0__abc_48231_n501), .B(u3_u0__abc_48231_n498), .Y(u3_u0_r3_23__FF_INPUT) );
  AND2X2 AND2X2_5226 ( .A(u3_u0__abc_48231_n382_bF_buf6), .B(u3_u0__abc_48231_n504_1), .Y(u3_u0__abc_48231_n505) );
  AND2X2 AND2X2_5227 ( .A(u3_u0__abc_48231_n506), .B(u3_u0__abc_48231_n503), .Y(u3_u0_r3_24__FF_INPUT) );
  AND2X2 AND2X2_5228 ( .A(u3_u0__abc_48231_n382_bF_buf4), .B(u3_u0__abc_48231_n509), .Y(u3_u0__abc_48231_n510) );
  AND2X2 AND2X2_5229 ( .A(u3_u0__abc_48231_n511), .B(u3_u0__abc_48231_n508_1), .Y(u3_u0_r3_25__FF_INPUT) );
  AND2X2 AND2X2_523 ( .A(spec_req_cs_1_bF_buf3), .B(u0_csc1_2_), .Y(u0__abc_49347_n2019) );
  AND2X2 AND2X2_5230 ( .A(u3_u0__abc_48231_n382_bF_buf2), .B(u3_u0__abc_48231_n514_1), .Y(u3_u0__abc_48231_n515) );
  AND2X2 AND2X2_5231 ( .A(u3_u0__abc_48231_n516), .B(u3_u0__abc_48231_n513_1), .Y(u3_u0_r3_26__FF_INPUT) );
  AND2X2 AND2X2_5232 ( .A(u3_u0__abc_48231_n382_bF_buf0), .B(u3_u0__abc_48231_n519), .Y(u3_u0__abc_48231_n520) );
  AND2X2 AND2X2_5233 ( .A(u3_u0__abc_48231_n521), .B(u3_u0__abc_48231_n518), .Y(u3_u0_r3_27__FF_INPUT) );
  AND2X2 AND2X2_5234 ( .A(u3_u0__abc_48231_n382_bF_buf6), .B(u3_u0__abc_48231_n524), .Y(u3_u0__abc_48231_n525) );
  AND2X2 AND2X2_5235 ( .A(u3_u0__abc_48231_n526), .B(u3_u0__abc_48231_n523), .Y(u3_u0_r3_28__FF_INPUT) );
  AND2X2 AND2X2_5236 ( .A(u3_u0__abc_48231_n382_bF_buf4), .B(u3_u0__abc_48231_n529), .Y(u3_u0__abc_48231_n530) );
  AND2X2 AND2X2_5237 ( .A(u3_u0__abc_48231_n531), .B(u3_u0__abc_48231_n528), .Y(u3_u0_r3_29__FF_INPUT) );
  AND2X2 AND2X2_5238 ( .A(u3_u0__abc_48231_n382_bF_buf2), .B(u3_u0__abc_48231_n534), .Y(u3_u0__abc_48231_n535) );
  AND2X2 AND2X2_5239 ( .A(u3_u0__abc_48231_n536), .B(u3_u0__abc_48231_n533), .Y(u3_u0_r3_30__FF_INPUT) );
  AND2X2 AND2X2_524 ( .A(u0__abc_49347_n1952_1_bF_buf1), .B(u0__abc_49347_n2022), .Y(u0__abc_49347_n2023) );
  AND2X2 AND2X2_5240 ( .A(u3_u0__abc_48231_n382_bF_buf0), .B(u3_u0__abc_48231_n539), .Y(u3_u0__abc_48231_n540) );
  AND2X2 AND2X2_5241 ( .A(u3_u0__abc_48231_n541), .B(u3_u0__abc_48231_n538), .Y(u3_u0_r3_31__FF_INPUT) );
  AND2X2 AND2X2_5242 ( .A(u3_u0__abc_48231_n382_bF_buf6), .B(u3_u0__abc_48231_n544), .Y(u3_u0__abc_48231_n545) );
  AND2X2 AND2X2_5243 ( .A(u3_u0__abc_48231_n546), .B(u3_u0__abc_48231_n543), .Y(u3_u0_r3_32__FF_INPUT) );
  AND2X2 AND2X2_5244 ( .A(u3_u0__abc_48231_n382_bF_buf4), .B(u3_u0__abc_48231_n549), .Y(u3_u0__abc_48231_n550) );
  AND2X2 AND2X2_5245 ( .A(u3_u0__abc_48231_n551), .B(u3_u0__abc_48231_n548), .Y(u3_u0_r3_33__FF_INPUT) );
  AND2X2 AND2X2_5246 ( .A(u3_u0__abc_48231_n382_bF_buf2), .B(u3_u0__abc_48231_n554), .Y(u3_u0__abc_48231_n555) );
  AND2X2 AND2X2_5247 ( .A(u3_u0__abc_48231_n556), .B(u3_u0__abc_48231_n553), .Y(u3_u0_r3_34__FF_INPUT) );
  AND2X2 AND2X2_5248 ( .A(u3_u0__abc_48231_n382_bF_buf0), .B(u3_u0__abc_48231_n559), .Y(u3_u0__abc_48231_n560) );
  AND2X2 AND2X2_5249 ( .A(u3_u0__abc_48231_n561), .B(u3_u0__abc_48231_n558), .Y(u3_u0_r3_35__FF_INPUT) );
  AND2X2 AND2X2_525 ( .A(u0__abc_49347_n2021), .B(u0__abc_49347_n2023), .Y(u0__abc_49347_n2024) );
  AND2X2 AND2X2_5250 ( .A(dv), .B(u3_u0_wr_adr_2_), .Y(u3_u0__abc_48231_n563) );
  AND2X2 AND2X2_5251 ( .A(u3_u0__abc_48231_n563_bF_buf6), .B(u3_u0__abc_48231_n384_1), .Y(u3_u0__abc_48231_n565) );
  AND2X2 AND2X2_5252 ( .A(u3_u0__abc_48231_n566), .B(u3_u0__abc_48231_n564), .Y(u3_u0_r2_0__FF_INPUT) );
  AND2X2 AND2X2_5253 ( .A(u3_u0__abc_48231_n563_bF_buf4), .B(u3_u0__abc_48231_n389), .Y(u3_u0__abc_48231_n569) );
  AND2X2 AND2X2_5254 ( .A(u3_u0__abc_48231_n570), .B(u3_u0__abc_48231_n568), .Y(u3_u0_r2_1__FF_INPUT) );
  AND2X2 AND2X2_5255 ( .A(u3_u0__abc_48231_n563_bF_buf2), .B(u3_u0__abc_48231_n394), .Y(u3_u0__abc_48231_n573) );
  AND2X2 AND2X2_5256 ( .A(u3_u0__abc_48231_n574), .B(u3_u0__abc_48231_n572), .Y(u3_u0_r2_2__FF_INPUT) );
  AND2X2 AND2X2_5257 ( .A(u3_u0__abc_48231_n563_bF_buf0), .B(u3_u0__abc_48231_n399), .Y(u3_u0__abc_48231_n577) );
  AND2X2 AND2X2_5258 ( .A(u3_u0__abc_48231_n578), .B(u3_u0__abc_48231_n576), .Y(u3_u0_r2_3__FF_INPUT) );
  AND2X2 AND2X2_5259 ( .A(u3_u0__abc_48231_n563_bF_buf6), .B(u3_u0__abc_48231_n404_1), .Y(u3_u0__abc_48231_n581) );
  AND2X2 AND2X2_526 ( .A(u0__abc_49347_n1953_1_bF_buf1), .B(sp_csc_3_), .Y(u0__abc_49347_n2026) );
  AND2X2 AND2X2_5260 ( .A(u3_u0__abc_48231_n582), .B(u3_u0__abc_48231_n580), .Y(u3_u0_r2_4__FF_INPUT) );
  AND2X2 AND2X2_5261 ( .A(u3_u0__abc_48231_n563_bF_buf4), .B(u3_u0__abc_48231_n409), .Y(u3_u0__abc_48231_n585) );
  AND2X2 AND2X2_5262 ( .A(u3_u0__abc_48231_n586), .B(u3_u0__abc_48231_n584), .Y(u3_u0_r2_5__FF_INPUT) );
  AND2X2 AND2X2_5263 ( .A(u3_u0__abc_48231_n563_bF_buf2), .B(u3_u0__abc_48231_n414), .Y(u3_u0__abc_48231_n589) );
  AND2X2 AND2X2_5264 ( .A(u3_u0__abc_48231_n590), .B(u3_u0__abc_48231_n588), .Y(u3_u0_r2_6__FF_INPUT) );
  AND2X2 AND2X2_5265 ( .A(u3_u0__abc_48231_n563_bF_buf0), .B(u3_u0__abc_48231_n419), .Y(u3_u0__abc_48231_n593) );
  AND2X2 AND2X2_5266 ( .A(u3_u0__abc_48231_n594), .B(u3_u0__abc_48231_n592), .Y(u3_u0_r2_7__FF_INPUT) );
  AND2X2 AND2X2_5267 ( .A(u3_u0__abc_48231_n563_bF_buf6), .B(u3_u0__abc_48231_n424_1), .Y(u3_u0__abc_48231_n597) );
  AND2X2 AND2X2_5268 ( .A(u3_u0__abc_48231_n598), .B(u3_u0__abc_48231_n596), .Y(u3_u0_r2_8__FF_INPUT) );
  AND2X2 AND2X2_5269 ( .A(u3_u0__abc_48231_n563_bF_buf4), .B(u3_u0__abc_48231_n429), .Y(u3_u0__abc_48231_n601) );
  AND2X2 AND2X2_527 ( .A(spec_req_cs_5_bF_buf2), .B(u0_csc5_3_), .Y(u0__abc_49347_n2027) );
  AND2X2 AND2X2_5270 ( .A(u3_u0__abc_48231_n602), .B(u3_u0__abc_48231_n600), .Y(u3_u0_r2_9__FF_INPUT) );
  AND2X2 AND2X2_5271 ( .A(u3_u0__abc_48231_n563_bF_buf2), .B(u3_u0__abc_48231_n434), .Y(u3_u0__abc_48231_n605) );
  AND2X2 AND2X2_5272 ( .A(u3_u0__abc_48231_n606), .B(u3_u0__abc_48231_n604), .Y(u3_u0_r2_10__FF_INPUT) );
  AND2X2 AND2X2_5273 ( .A(u3_u0__abc_48231_n563_bF_buf0), .B(u3_u0__abc_48231_n439), .Y(u3_u0__abc_48231_n609) );
  AND2X2 AND2X2_5274 ( .A(u3_u0__abc_48231_n610), .B(u3_u0__abc_48231_n608), .Y(u3_u0_r2_11__FF_INPUT) );
  AND2X2 AND2X2_5275 ( .A(u3_u0__abc_48231_n563_bF_buf6), .B(u3_u0__abc_48231_n444_1), .Y(u3_u0__abc_48231_n613) );
  AND2X2 AND2X2_5276 ( .A(u3_u0__abc_48231_n614), .B(u3_u0__abc_48231_n612), .Y(u3_u0_r2_12__FF_INPUT) );
  AND2X2 AND2X2_5277 ( .A(u3_u0__abc_48231_n563_bF_buf4), .B(u3_u0__abc_48231_n449), .Y(u3_u0__abc_48231_n617) );
  AND2X2 AND2X2_5278 ( .A(u3_u0__abc_48231_n618), .B(u3_u0__abc_48231_n616), .Y(u3_u0_r2_13__FF_INPUT) );
  AND2X2 AND2X2_5279 ( .A(u3_u0__abc_48231_n563_bF_buf2), .B(u3_u0__abc_48231_n454), .Y(u3_u0__abc_48231_n621) );
  AND2X2 AND2X2_528 ( .A(u0__abc_49347_n2029), .B(u0__abc_49347_n1185_bF_buf5), .Y(u0__abc_49347_n2030) );
  AND2X2 AND2X2_5280 ( .A(u3_u0__abc_48231_n622), .B(u3_u0__abc_48231_n620), .Y(u3_u0_r2_14__FF_INPUT) );
  AND2X2 AND2X2_5281 ( .A(u3_u0__abc_48231_n563_bF_buf0), .B(u3_u0__abc_48231_n459), .Y(u3_u0__abc_48231_n625) );
  AND2X2 AND2X2_5282 ( .A(u3_u0__abc_48231_n626), .B(u3_u0__abc_48231_n624), .Y(u3_u0_r2_15__FF_INPUT) );
  AND2X2 AND2X2_5283 ( .A(u3_u0__abc_48231_n563_bF_buf6), .B(u3_u0__abc_48231_n464_1), .Y(u3_u0__abc_48231_n629) );
  AND2X2 AND2X2_5284 ( .A(u3_u0__abc_48231_n630), .B(u3_u0__abc_48231_n628), .Y(u3_u0_r2_16__FF_INPUT) );
  AND2X2 AND2X2_5285 ( .A(u3_u0__abc_48231_n563_bF_buf4), .B(u3_u0__abc_48231_n469), .Y(u3_u0__abc_48231_n633) );
  AND2X2 AND2X2_5286 ( .A(u3_u0__abc_48231_n634), .B(u3_u0__abc_48231_n632), .Y(u3_u0_r2_17__FF_INPUT) );
  AND2X2 AND2X2_5287 ( .A(u3_u0__abc_48231_n563_bF_buf2), .B(u3_u0__abc_48231_n474), .Y(u3_u0__abc_48231_n637) );
  AND2X2 AND2X2_5288 ( .A(u3_u0__abc_48231_n638), .B(u3_u0__abc_48231_n636), .Y(u3_u0_r2_18__FF_INPUT) );
  AND2X2 AND2X2_5289 ( .A(u3_u0__abc_48231_n563_bF_buf0), .B(u3_u0__abc_48231_n479), .Y(u3_u0__abc_48231_n641) );
  AND2X2 AND2X2_529 ( .A(u0__abc_49347_n2030), .B(u0__abc_49347_n2028), .Y(u0__abc_49347_n2031) );
  AND2X2 AND2X2_5290 ( .A(u3_u0__abc_48231_n642), .B(u3_u0__abc_48231_n640), .Y(u3_u0_r2_19__FF_INPUT) );
  AND2X2 AND2X2_5291 ( .A(u3_u0__abc_48231_n563_bF_buf6), .B(u3_u0__abc_48231_n484_1), .Y(u3_u0__abc_48231_n645) );
  AND2X2 AND2X2_5292 ( .A(u3_u0__abc_48231_n646), .B(u3_u0__abc_48231_n644), .Y(u3_u0_r2_20__FF_INPUT) );
  AND2X2 AND2X2_5293 ( .A(u3_u0__abc_48231_n563_bF_buf4), .B(u3_u0__abc_48231_n489), .Y(u3_u0__abc_48231_n649) );
  AND2X2 AND2X2_5294 ( .A(u3_u0__abc_48231_n650), .B(u3_u0__abc_48231_n648), .Y(u3_u0_r2_21__FF_INPUT) );
  AND2X2 AND2X2_5295 ( .A(u3_u0__abc_48231_n563_bF_buf2), .B(u3_u0__abc_48231_n494), .Y(u3_u0__abc_48231_n653) );
  AND2X2 AND2X2_5296 ( .A(u3_u0__abc_48231_n654), .B(u3_u0__abc_48231_n652), .Y(u3_u0_r2_22__FF_INPUT) );
  AND2X2 AND2X2_5297 ( .A(u3_u0__abc_48231_n563_bF_buf0), .B(u3_u0__abc_48231_n499), .Y(u3_u0__abc_48231_n657) );
  AND2X2 AND2X2_5298 ( .A(u3_u0__abc_48231_n658), .B(u3_u0__abc_48231_n656), .Y(u3_u0_r2_23__FF_INPUT) );
  AND2X2 AND2X2_5299 ( .A(u3_u0__abc_48231_n563_bF_buf6), .B(u3_u0__abc_48231_n504_1), .Y(u3_u0__abc_48231_n661) );
  AND2X2 AND2X2_53 ( .A(_abc_55805_n413), .B(_abc_55805_n414), .Y(u1_bas) );
  AND2X2 AND2X2_530 ( .A(u0__abc_49347_n2032), .B(u0__abc_49347_n1181_bF_buf5), .Y(u0__abc_49347_n2033) );
  AND2X2 AND2X2_5300 ( .A(u3_u0__abc_48231_n662), .B(u3_u0__abc_48231_n660), .Y(u3_u0_r2_24__FF_INPUT) );
  AND2X2 AND2X2_5301 ( .A(u3_u0__abc_48231_n563_bF_buf4), .B(u3_u0__abc_48231_n509), .Y(u3_u0__abc_48231_n665) );
  AND2X2 AND2X2_5302 ( .A(u3_u0__abc_48231_n666), .B(u3_u0__abc_48231_n664), .Y(u3_u0_r2_25__FF_INPUT) );
  AND2X2 AND2X2_5303 ( .A(u3_u0__abc_48231_n563_bF_buf2), .B(u3_u0__abc_48231_n514_1), .Y(u3_u0__abc_48231_n669) );
  AND2X2 AND2X2_5304 ( .A(u3_u0__abc_48231_n670), .B(u3_u0__abc_48231_n668), .Y(u3_u0_r2_26__FF_INPUT) );
  AND2X2 AND2X2_5305 ( .A(u3_u0__abc_48231_n563_bF_buf0), .B(u3_u0__abc_48231_n519), .Y(u3_u0__abc_48231_n673) );
  AND2X2 AND2X2_5306 ( .A(u3_u0__abc_48231_n674), .B(u3_u0__abc_48231_n672), .Y(u3_u0_r2_27__FF_INPUT) );
  AND2X2 AND2X2_5307 ( .A(u3_u0__abc_48231_n563_bF_buf6), .B(u3_u0__abc_48231_n524), .Y(u3_u0__abc_48231_n677) );
  AND2X2 AND2X2_5308 ( .A(u3_u0__abc_48231_n678), .B(u3_u0__abc_48231_n676), .Y(u3_u0_r2_28__FF_INPUT) );
  AND2X2 AND2X2_5309 ( .A(u3_u0__abc_48231_n563_bF_buf4), .B(u3_u0__abc_48231_n529), .Y(u3_u0__abc_48231_n681) );
  AND2X2 AND2X2_531 ( .A(spec_req_cs_4_bF_buf2), .B(u0_csc4_3_), .Y(u0__abc_49347_n2034) );
  AND2X2 AND2X2_5310 ( .A(u3_u0__abc_48231_n682), .B(u3_u0__abc_48231_n680), .Y(u3_u0_r2_29__FF_INPUT) );
  AND2X2 AND2X2_5311 ( .A(u3_u0__abc_48231_n563_bF_buf2), .B(u3_u0__abc_48231_n534), .Y(u3_u0__abc_48231_n685) );
  AND2X2 AND2X2_5312 ( .A(u3_u0__abc_48231_n686), .B(u3_u0__abc_48231_n684), .Y(u3_u0_r2_30__FF_INPUT) );
  AND2X2 AND2X2_5313 ( .A(u3_u0__abc_48231_n563_bF_buf0), .B(u3_u0__abc_48231_n539), .Y(u3_u0__abc_48231_n689) );
  AND2X2 AND2X2_5314 ( .A(u3_u0__abc_48231_n690), .B(u3_u0__abc_48231_n688), .Y(u3_u0_r2_31__FF_INPUT) );
  AND2X2 AND2X2_5315 ( .A(u3_u0__abc_48231_n563_bF_buf6), .B(u3_u0__abc_48231_n544), .Y(u3_u0__abc_48231_n693) );
  AND2X2 AND2X2_5316 ( .A(u3_u0__abc_48231_n694), .B(u3_u0__abc_48231_n692), .Y(u3_u0_r2_32__FF_INPUT) );
  AND2X2 AND2X2_5317 ( .A(u3_u0__abc_48231_n563_bF_buf4), .B(u3_u0__abc_48231_n549), .Y(u3_u0__abc_48231_n697) );
  AND2X2 AND2X2_5318 ( .A(u3_u0__abc_48231_n698), .B(u3_u0__abc_48231_n696), .Y(u3_u0_r2_33__FF_INPUT) );
  AND2X2 AND2X2_5319 ( .A(u3_u0__abc_48231_n563_bF_buf2), .B(u3_u0__abc_48231_n554), .Y(u3_u0__abc_48231_n701) );
  AND2X2 AND2X2_532 ( .A(u0__abc_49347_n2035), .B(u0__abc_49347_n1180_1_bF_buf5), .Y(u0__abc_49347_n2036) );
  AND2X2 AND2X2_5320 ( .A(u3_u0__abc_48231_n702), .B(u3_u0__abc_48231_n700), .Y(u3_u0_r2_34__FF_INPUT) );
  AND2X2 AND2X2_5321 ( .A(u3_u0__abc_48231_n563_bF_buf0), .B(u3_u0__abc_48231_n559), .Y(u3_u0__abc_48231_n705) );
  AND2X2 AND2X2_5322 ( .A(u3_u0__abc_48231_n706), .B(u3_u0__abc_48231_n704), .Y(u3_u0_r2_35__FF_INPUT) );
  AND2X2 AND2X2_5323 ( .A(dv), .B(u3_u0_wr_adr_1_), .Y(u3_u0__abc_48231_n708) );
  AND2X2 AND2X2_5324 ( .A(u3_u0__abc_48231_n708_bF_buf6), .B(u3_u0__abc_48231_n384_1), .Y(u3_u0__abc_48231_n710) );
  AND2X2 AND2X2_5325 ( .A(u3_u0__abc_48231_n711), .B(u3_u0__abc_48231_n709), .Y(u3_u0_r1_0__FF_INPUT) );
  AND2X2 AND2X2_5326 ( .A(u3_u0__abc_48231_n708_bF_buf4), .B(u3_u0__abc_48231_n389), .Y(u3_u0__abc_48231_n714) );
  AND2X2 AND2X2_5327 ( .A(u3_u0__abc_48231_n715), .B(u3_u0__abc_48231_n713), .Y(u3_u0_r1_1__FF_INPUT) );
  AND2X2 AND2X2_5328 ( .A(u3_u0__abc_48231_n708_bF_buf2), .B(u3_u0__abc_48231_n394), .Y(u3_u0__abc_48231_n718) );
  AND2X2 AND2X2_5329 ( .A(u3_u0__abc_48231_n719), .B(u3_u0__abc_48231_n717), .Y(u3_u0_r1_2__FF_INPUT) );
  AND2X2 AND2X2_533 ( .A(spec_req_cs_3_bF_buf2), .B(u0_csc3_3_), .Y(u0__abc_49347_n2037) );
  AND2X2 AND2X2_5330 ( .A(u3_u0__abc_48231_n708_bF_buf0), .B(u3_u0__abc_48231_n399), .Y(u3_u0__abc_48231_n722) );
  AND2X2 AND2X2_5331 ( .A(u3_u0__abc_48231_n723), .B(u3_u0__abc_48231_n721), .Y(u3_u0_r1_3__FF_INPUT) );
  AND2X2 AND2X2_5332 ( .A(u3_u0__abc_48231_n708_bF_buf6), .B(u3_u0__abc_48231_n404_1), .Y(u3_u0__abc_48231_n726) );
  AND2X2 AND2X2_5333 ( .A(u3_u0__abc_48231_n727), .B(u3_u0__abc_48231_n725), .Y(u3_u0_r1_4__FF_INPUT) );
  AND2X2 AND2X2_5334 ( .A(u3_u0__abc_48231_n708_bF_buf4), .B(u3_u0__abc_48231_n409), .Y(u3_u0__abc_48231_n730) );
  AND2X2 AND2X2_5335 ( .A(u3_u0__abc_48231_n731), .B(u3_u0__abc_48231_n729), .Y(u3_u0_r1_5__FF_INPUT) );
  AND2X2 AND2X2_5336 ( .A(u3_u0__abc_48231_n708_bF_buf2), .B(u3_u0__abc_48231_n414), .Y(u3_u0__abc_48231_n734) );
  AND2X2 AND2X2_5337 ( .A(u3_u0__abc_48231_n735), .B(u3_u0__abc_48231_n733), .Y(u3_u0_r1_6__FF_INPUT) );
  AND2X2 AND2X2_5338 ( .A(u3_u0__abc_48231_n708_bF_buf0), .B(u3_u0__abc_48231_n419), .Y(u3_u0__abc_48231_n738) );
  AND2X2 AND2X2_5339 ( .A(u3_u0__abc_48231_n739), .B(u3_u0__abc_48231_n737), .Y(u3_u0_r1_7__FF_INPUT) );
  AND2X2 AND2X2_534 ( .A(u0__abc_49347_n2038), .B(u0__abc_49347_n1179_bF_buf5), .Y(u0__abc_49347_n2039) );
  AND2X2 AND2X2_5340 ( .A(u3_u0__abc_48231_n708_bF_buf6), .B(u3_u0__abc_48231_n424_1), .Y(u3_u0__abc_48231_n742) );
  AND2X2 AND2X2_5341 ( .A(u3_u0__abc_48231_n743), .B(u3_u0__abc_48231_n741), .Y(u3_u0_r1_8__FF_INPUT) );
  AND2X2 AND2X2_5342 ( .A(u3_u0__abc_48231_n708_bF_buf4), .B(u3_u0__abc_48231_n429), .Y(u3_u0__abc_48231_n746) );
  AND2X2 AND2X2_5343 ( .A(u3_u0__abc_48231_n747), .B(u3_u0__abc_48231_n745), .Y(u3_u0_r1_9__FF_INPUT) );
  AND2X2 AND2X2_5344 ( .A(u3_u0__abc_48231_n708_bF_buf2), .B(u3_u0__abc_48231_n434), .Y(u3_u0__abc_48231_n750) );
  AND2X2 AND2X2_5345 ( .A(u3_u0__abc_48231_n751), .B(u3_u0__abc_48231_n749), .Y(u3_u0_r1_10__FF_INPUT) );
  AND2X2 AND2X2_5346 ( .A(u3_u0__abc_48231_n708_bF_buf0), .B(u3_u0__abc_48231_n439), .Y(u3_u0__abc_48231_n754) );
  AND2X2 AND2X2_5347 ( .A(u3_u0__abc_48231_n755), .B(u3_u0__abc_48231_n753), .Y(u3_u0_r1_11__FF_INPUT) );
  AND2X2 AND2X2_5348 ( .A(u3_u0__abc_48231_n708_bF_buf6), .B(u3_u0__abc_48231_n444_1), .Y(u3_u0__abc_48231_n758) );
  AND2X2 AND2X2_5349 ( .A(u3_u0__abc_48231_n759), .B(u3_u0__abc_48231_n757), .Y(u3_u0_r1_12__FF_INPUT) );
  AND2X2 AND2X2_535 ( .A(spec_req_cs_2_bF_buf2), .B(u0_csc2_3_), .Y(u0__abc_49347_n2040) );
  AND2X2 AND2X2_5350 ( .A(u3_u0__abc_48231_n708_bF_buf4), .B(u3_u0__abc_48231_n449), .Y(u3_u0__abc_48231_n762) );
  AND2X2 AND2X2_5351 ( .A(u3_u0__abc_48231_n763), .B(u3_u0__abc_48231_n761), .Y(u3_u0_r1_13__FF_INPUT) );
  AND2X2 AND2X2_5352 ( .A(u3_u0__abc_48231_n708_bF_buf2), .B(u3_u0__abc_48231_n454), .Y(u3_u0__abc_48231_n766) );
  AND2X2 AND2X2_5353 ( .A(u3_u0__abc_48231_n767), .B(u3_u0__abc_48231_n765), .Y(u3_u0_r1_14__FF_INPUT) );
  AND2X2 AND2X2_5354 ( .A(u3_u0__abc_48231_n708_bF_buf0), .B(u3_u0__abc_48231_n459), .Y(u3_u0__abc_48231_n770) );
  AND2X2 AND2X2_5355 ( .A(u3_u0__abc_48231_n771), .B(u3_u0__abc_48231_n769), .Y(u3_u0_r1_15__FF_INPUT) );
  AND2X2 AND2X2_5356 ( .A(u3_u0__abc_48231_n708_bF_buf6), .B(u3_u0__abc_48231_n464_1), .Y(u3_u0__abc_48231_n774) );
  AND2X2 AND2X2_5357 ( .A(u3_u0__abc_48231_n775), .B(u3_u0__abc_48231_n773), .Y(u3_u0_r1_16__FF_INPUT) );
  AND2X2 AND2X2_5358 ( .A(u3_u0__abc_48231_n708_bF_buf4), .B(u3_u0__abc_48231_n469), .Y(u3_u0__abc_48231_n778) );
  AND2X2 AND2X2_5359 ( .A(u3_u0__abc_48231_n779), .B(u3_u0__abc_48231_n777), .Y(u3_u0_r1_17__FF_INPUT) );
  AND2X2 AND2X2_536 ( .A(u0__abc_49347_n2041), .B(u0__abc_49347_n1178_1_bF_buf5), .Y(u0__abc_49347_n2042) );
  AND2X2 AND2X2_5360 ( .A(u3_u0__abc_48231_n708_bF_buf2), .B(u3_u0__abc_48231_n474), .Y(u3_u0__abc_48231_n782) );
  AND2X2 AND2X2_5361 ( .A(u3_u0__abc_48231_n783), .B(u3_u0__abc_48231_n781), .Y(u3_u0_r1_18__FF_INPUT) );
  AND2X2 AND2X2_5362 ( .A(u3_u0__abc_48231_n708_bF_buf0), .B(u3_u0__abc_48231_n479), .Y(u3_u0__abc_48231_n786) );
  AND2X2 AND2X2_5363 ( .A(u3_u0__abc_48231_n787), .B(u3_u0__abc_48231_n785), .Y(u3_u0_r1_19__FF_INPUT) );
  AND2X2 AND2X2_5364 ( .A(u3_u0__abc_48231_n708_bF_buf6), .B(u3_u0__abc_48231_n484_1), .Y(u3_u0__abc_48231_n790) );
  AND2X2 AND2X2_5365 ( .A(u3_u0__abc_48231_n791), .B(u3_u0__abc_48231_n789), .Y(u3_u0_r1_20__FF_INPUT) );
  AND2X2 AND2X2_5366 ( .A(u3_u0__abc_48231_n708_bF_buf4), .B(u3_u0__abc_48231_n489), .Y(u3_u0__abc_48231_n794) );
  AND2X2 AND2X2_5367 ( .A(u3_u0__abc_48231_n795), .B(u3_u0__abc_48231_n793), .Y(u3_u0_r1_21__FF_INPUT) );
  AND2X2 AND2X2_5368 ( .A(u3_u0__abc_48231_n708_bF_buf2), .B(u3_u0__abc_48231_n494), .Y(u3_u0__abc_48231_n798) );
  AND2X2 AND2X2_5369 ( .A(u3_u0__abc_48231_n799), .B(u3_u0__abc_48231_n797), .Y(u3_u0_r1_22__FF_INPUT) );
  AND2X2 AND2X2_537 ( .A(spec_req_cs_1_bF_buf2), .B(u0_csc1_3_), .Y(u0__abc_49347_n2043) );
  AND2X2 AND2X2_5370 ( .A(u3_u0__abc_48231_n708_bF_buf0), .B(u3_u0__abc_48231_n499), .Y(u3_u0__abc_48231_n802) );
  AND2X2 AND2X2_5371 ( .A(u3_u0__abc_48231_n803), .B(u3_u0__abc_48231_n801), .Y(u3_u0_r1_23__FF_INPUT) );
  AND2X2 AND2X2_5372 ( .A(u3_u0__abc_48231_n708_bF_buf6), .B(u3_u0__abc_48231_n504_1), .Y(u3_u0__abc_48231_n806) );
  AND2X2 AND2X2_5373 ( .A(u3_u0__abc_48231_n807), .B(u3_u0__abc_48231_n805), .Y(u3_u0_r1_24__FF_INPUT) );
  AND2X2 AND2X2_5374 ( .A(u3_u0__abc_48231_n708_bF_buf4), .B(u3_u0__abc_48231_n509), .Y(u3_u0__abc_48231_n810) );
  AND2X2 AND2X2_5375 ( .A(u3_u0__abc_48231_n811), .B(u3_u0__abc_48231_n809), .Y(u3_u0_r1_25__FF_INPUT) );
  AND2X2 AND2X2_5376 ( .A(u3_u0__abc_48231_n708_bF_buf2), .B(u3_u0__abc_48231_n514_1), .Y(u3_u0__abc_48231_n814) );
  AND2X2 AND2X2_5377 ( .A(u3_u0__abc_48231_n815), .B(u3_u0__abc_48231_n813), .Y(u3_u0_r1_26__FF_INPUT) );
  AND2X2 AND2X2_5378 ( .A(u3_u0__abc_48231_n708_bF_buf0), .B(u3_u0__abc_48231_n519), .Y(u3_u0__abc_48231_n818) );
  AND2X2 AND2X2_5379 ( .A(u3_u0__abc_48231_n819), .B(u3_u0__abc_48231_n817), .Y(u3_u0_r1_27__FF_INPUT) );
  AND2X2 AND2X2_538 ( .A(u0__abc_49347_n1952_1_bF_buf0), .B(u0__abc_49347_n2046), .Y(u0__abc_49347_n2047) );
  AND2X2 AND2X2_5380 ( .A(u3_u0__abc_48231_n708_bF_buf6), .B(u3_u0__abc_48231_n524), .Y(u3_u0__abc_48231_n822) );
  AND2X2 AND2X2_5381 ( .A(u3_u0__abc_48231_n823), .B(u3_u0__abc_48231_n821), .Y(u3_u0_r1_28__FF_INPUT) );
  AND2X2 AND2X2_5382 ( .A(u3_u0__abc_48231_n708_bF_buf4), .B(u3_u0__abc_48231_n529), .Y(u3_u0__abc_48231_n826) );
  AND2X2 AND2X2_5383 ( .A(u3_u0__abc_48231_n827), .B(u3_u0__abc_48231_n825), .Y(u3_u0_r1_29__FF_INPUT) );
  AND2X2 AND2X2_5384 ( .A(u3_u0__abc_48231_n708_bF_buf2), .B(u3_u0__abc_48231_n534), .Y(u3_u0__abc_48231_n830) );
  AND2X2 AND2X2_5385 ( .A(u3_u0__abc_48231_n831), .B(u3_u0__abc_48231_n829), .Y(u3_u0_r1_30__FF_INPUT) );
  AND2X2 AND2X2_5386 ( .A(u3_u0__abc_48231_n708_bF_buf0), .B(u3_u0__abc_48231_n539), .Y(u3_u0__abc_48231_n834) );
  AND2X2 AND2X2_5387 ( .A(u3_u0__abc_48231_n835), .B(u3_u0__abc_48231_n833), .Y(u3_u0_r1_31__FF_INPUT) );
  AND2X2 AND2X2_5388 ( .A(u3_u0__abc_48231_n708_bF_buf6), .B(u3_u0__abc_48231_n544), .Y(u3_u0__abc_48231_n838) );
  AND2X2 AND2X2_5389 ( .A(u3_u0__abc_48231_n839), .B(u3_u0__abc_48231_n837), .Y(u3_u0_r1_32__FF_INPUT) );
  AND2X2 AND2X2_539 ( .A(u0__abc_49347_n2045), .B(u0__abc_49347_n2047), .Y(u0__abc_49347_n2048) );
  AND2X2 AND2X2_5390 ( .A(u3_u0__abc_48231_n708_bF_buf4), .B(u3_u0__abc_48231_n549), .Y(u3_u0__abc_48231_n842) );
  AND2X2 AND2X2_5391 ( .A(u3_u0__abc_48231_n843), .B(u3_u0__abc_48231_n841), .Y(u3_u0_r1_33__FF_INPUT) );
  AND2X2 AND2X2_5392 ( .A(u3_u0__abc_48231_n708_bF_buf2), .B(u3_u0__abc_48231_n554), .Y(u3_u0__abc_48231_n846) );
  AND2X2 AND2X2_5393 ( .A(u3_u0__abc_48231_n847), .B(u3_u0__abc_48231_n845), .Y(u3_u0_r1_34__FF_INPUT) );
  AND2X2 AND2X2_5394 ( .A(u3_u0__abc_48231_n708_bF_buf0), .B(u3_u0__abc_48231_n559), .Y(u3_u0__abc_48231_n850) );
  AND2X2 AND2X2_5395 ( .A(u3_u0__abc_48231_n851), .B(u3_u0__abc_48231_n849), .Y(u3_u0_r1_35__FF_INPUT) );
  AND2X2 AND2X2_5396 ( .A(dv), .B(u3_u0_wr_adr_0_), .Y(u3_u0__abc_48231_n853) );
  AND2X2 AND2X2_5397 ( .A(u3_u0__abc_48231_n853_bF_buf6), .B(u3_u0__abc_48231_n384_1), .Y(u3_u0__abc_48231_n855) );
  AND2X2 AND2X2_5398 ( .A(u3_u0__abc_48231_n856), .B(u3_u0__abc_48231_n854), .Y(u3_u0_r0_0__FF_INPUT) );
  AND2X2 AND2X2_5399 ( .A(u3_u0__abc_48231_n853_bF_buf4), .B(u3_u0__abc_48231_n389), .Y(u3_u0__abc_48231_n859) );
  AND2X2 AND2X2_54 ( .A(_abc_55805_n416), .B(_abc_55805_n417), .Y(u5_kro) );
  AND2X2 AND2X2_540 ( .A(u0__abc_49347_n1953_1_bF_buf0), .B(sp_csc_4_), .Y(u0__abc_49347_n2050) );
  AND2X2 AND2X2_5400 ( .A(u3_u0__abc_48231_n860), .B(u3_u0__abc_48231_n858), .Y(u3_u0_r0_1__FF_INPUT) );
  AND2X2 AND2X2_5401 ( .A(u3_u0__abc_48231_n853_bF_buf2), .B(u3_u0__abc_48231_n394), .Y(u3_u0__abc_48231_n863) );
  AND2X2 AND2X2_5402 ( .A(u3_u0__abc_48231_n864), .B(u3_u0__abc_48231_n862), .Y(u3_u0_r0_2__FF_INPUT) );
  AND2X2 AND2X2_5403 ( .A(u3_u0__abc_48231_n853_bF_buf0), .B(u3_u0__abc_48231_n399), .Y(u3_u0__abc_48231_n867) );
  AND2X2 AND2X2_5404 ( .A(u3_u0__abc_48231_n868), .B(u3_u0__abc_48231_n866), .Y(u3_u0_r0_3__FF_INPUT) );
  AND2X2 AND2X2_5405 ( .A(u3_u0__abc_48231_n853_bF_buf6), .B(u3_u0__abc_48231_n404_1), .Y(u3_u0__abc_48231_n871) );
  AND2X2 AND2X2_5406 ( .A(u3_u0__abc_48231_n872), .B(u3_u0__abc_48231_n870), .Y(u3_u0_r0_4__FF_INPUT) );
  AND2X2 AND2X2_5407 ( .A(u3_u0__abc_48231_n853_bF_buf4), .B(u3_u0__abc_48231_n409), .Y(u3_u0__abc_48231_n875) );
  AND2X2 AND2X2_5408 ( .A(u3_u0__abc_48231_n876), .B(u3_u0__abc_48231_n874), .Y(u3_u0_r0_5__FF_INPUT) );
  AND2X2 AND2X2_5409 ( .A(u3_u0__abc_48231_n853_bF_buf2), .B(u3_u0__abc_48231_n414), .Y(u3_u0__abc_48231_n879) );
  AND2X2 AND2X2_541 ( .A(spec_req_cs_5_bF_buf1), .B(u0_csc5_4_), .Y(u0__abc_49347_n2051_1) );
  AND2X2 AND2X2_5410 ( .A(u3_u0__abc_48231_n880), .B(u3_u0__abc_48231_n878), .Y(u3_u0_r0_6__FF_INPUT) );
  AND2X2 AND2X2_5411 ( .A(u3_u0__abc_48231_n853_bF_buf0), .B(u3_u0__abc_48231_n419), .Y(u3_u0__abc_48231_n883) );
  AND2X2 AND2X2_5412 ( .A(u3_u0__abc_48231_n884), .B(u3_u0__abc_48231_n882), .Y(u3_u0_r0_7__FF_INPUT) );
  AND2X2 AND2X2_5413 ( .A(u3_u0__abc_48231_n853_bF_buf6), .B(u3_u0__abc_48231_n424_1), .Y(u3_u0__abc_48231_n887) );
  AND2X2 AND2X2_5414 ( .A(u3_u0__abc_48231_n888), .B(u3_u0__abc_48231_n886), .Y(u3_u0_r0_8__FF_INPUT) );
  AND2X2 AND2X2_5415 ( .A(u3_u0__abc_48231_n853_bF_buf4), .B(u3_u0__abc_48231_n429), .Y(u3_u0__abc_48231_n891) );
  AND2X2 AND2X2_5416 ( .A(u3_u0__abc_48231_n892), .B(u3_u0__abc_48231_n890), .Y(u3_u0_r0_9__FF_INPUT) );
  AND2X2 AND2X2_5417 ( .A(u3_u0__abc_48231_n853_bF_buf2), .B(u3_u0__abc_48231_n434), .Y(u3_u0__abc_48231_n895) );
  AND2X2 AND2X2_5418 ( .A(u3_u0__abc_48231_n896), .B(u3_u0__abc_48231_n894), .Y(u3_u0_r0_10__FF_INPUT) );
  AND2X2 AND2X2_5419 ( .A(u3_u0__abc_48231_n853_bF_buf0), .B(u3_u0__abc_48231_n439), .Y(u3_u0__abc_48231_n899) );
  AND2X2 AND2X2_542 ( .A(u0__abc_49347_n2053), .B(u0__abc_49347_n1185_bF_buf4), .Y(u0__abc_49347_n2054) );
  AND2X2 AND2X2_5420 ( .A(u3_u0__abc_48231_n900), .B(u3_u0__abc_48231_n898), .Y(u3_u0_r0_11__FF_INPUT) );
  AND2X2 AND2X2_5421 ( .A(u3_u0__abc_48231_n853_bF_buf6), .B(u3_u0__abc_48231_n444_1), .Y(u3_u0__abc_48231_n903) );
  AND2X2 AND2X2_5422 ( .A(u3_u0__abc_48231_n904), .B(u3_u0__abc_48231_n902), .Y(u3_u0_r0_12__FF_INPUT) );
  AND2X2 AND2X2_5423 ( .A(u3_u0__abc_48231_n853_bF_buf4), .B(u3_u0__abc_48231_n449), .Y(u3_u0__abc_48231_n907) );
  AND2X2 AND2X2_5424 ( .A(u3_u0__abc_48231_n908), .B(u3_u0__abc_48231_n906), .Y(u3_u0_r0_13__FF_INPUT) );
  AND2X2 AND2X2_5425 ( .A(u3_u0__abc_48231_n853_bF_buf2), .B(u3_u0__abc_48231_n454), .Y(u3_u0__abc_48231_n911) );
  AND2X2 AND2X2_5426 ( .A(u3_u0__abc_48231_n912), .B(u3_u0__abc_48231_n910), .Y(u3_u0_r0_14__FF_INPUT) );
  AND2X2 AND2X2_5427 ( .A(u3_u0__abc_48231_n853_bF_buf0), .B(u3_u0__abc_48231_n459), .Y(u3_u0__abc_48231_n915) );
  AND2X2 AND2X2_5428 ( .A(u3_u0__abc_48231_n916), .B(u3_u0__abc_48231_n914), .Y(u3_u0_r0_15__FF_INPUT) );
  AND2X2 AND2X2_5429 ( .A(u3_u0__abc_48231_n853_bF_buf6), .B(u3_u0__abc_48231_n464_1), .Y(u3_u0__abc_48231_n919) );
  AND2X2 AND2X2_543 ( .A(u0__abc_49347_n2054), .B(u0__abc_49347_n2052), .Y(u0__abc_49347_n2055) );
  AND2X2 AND2X2_5430 ( .A(u3_u0__abc_48231_n920), .B(u3_u0__abc_48231_n918), .Y(u3_u0_r0_16__FF_INPUT) );
  AND2X2 AND2X2_5431 ( .A(u3_u0__abc_48231_n853_bF_buf4), .B(u3_u0__abc_48231_n469), .Y(u3_u0__abc_48231_n923) );
  AND2X2 AND2X2_5432 ( .A(u3_u0__abc_48231_n924), .B(u3_u0__abc_48231_n922), .Y(u3_u0_r0_17__FF_INPUT) );
  AND2X2 AND2X2_5433 ( .A(u3_u0__abc_48231_n853_bF_buf2), .B(u3_u0__abc_48231_n474), .Y(u3_u0__abc_48231_n927) );
  AND2X2 AND2X2_5434 ( .A(u3_u0__abc_48231_n928), .B(u3_u0__abc_48231_n926), .Y(u3_u0_r0_18__FF_INPUT) );
  AND2X2 AND2X2_5435 ( .A(u3_u0__abc_48231_n853_bF_buf0), .B(u3_u0__abc_48231_n479), .Y(u3_u0__abc_48231_n931) );
  AND2X2 AND2X2_5436 ( .A(u3_u0__abc_48231_n932), .B(u3_u0__abc_48231_n930), .Y(u3_u0_r0_19__FF_INPUT) );
  AND2X2 AND2X2_5437 ( .A(u3_u0__abc_48231_n853_bF_buf6), .B(u3_u0__abc_48231_n484_1), .Y(u3_u0__abc_48231_n935) );
  AND2X2 AND2X2_5438 ( .A(u3_u0__abc_48231_n936), .B(u3_u0__abc_48231_n934), .Y(u3_u0_r0_20__FF_INPUT) );
  AND2X2 AND2X2_5439 ( .A(u3_u0__abc_48231_n853_bF_buf4), .B(u3_u0__abc_48231_n489), .Y(u3_u0__abc_48231_n939) );
  AND2X2 AND2X2_544 ( .A(u0__abc_49347_n2056), .B(u0__abc_49347_n1181_bF_buf4), .Y(u0__abc_49347_n2057) );
  AND2X2 AND2X2_5440 ( .A(u3_u0__abc_48231_n940), .B(u3_u0__abc_48231_n938), .Y(u3_u0_r0_21__FF_INPUT) );
  AND2X2 AND2X2_5441 ( .A(u3_u0__abc_48231_n853_bF_buf2), .B(u3_u0__abc_48231_n494), .Y(u3_u0__abc_48231_n943) );
  AND2X2 AND2X2_5442 ( .A(u3_u0__abc_48231_n944), .B(u3_u0__abc_48231_n942), .Y(u3_u0_r0_22__FF_INPUT) );
  AND2X2 AND2X2_5443 ( .A(u3_u0__abc_48231_n853_bF_buf0), .B(u3_u0__abc_48231_n499), .Y(u3_u0__abc_48231_n947) );
  AND2X2 AND2X2_5444 ( .A(u3_u0__abc_48231_n948), .B(u3_u0__abc_48231_n946), .Y(u3_u0_r0_23__FF_INPUT) );
  AND2X2 AND2X2_5445 ( .A(u3_u0__abc_48231_n853_bF_buf6), .B(u3_u0__abc_48231_n504_1), .Y(u3_u0__abc_48231_n951) );
  AND2X2 AND2X2_5446 ( .A(u3_u0__abc_48231_n952), .B(u3_u0__abc_48231_n950), .Y(u3_u0_r0_24__FF_INPUT) );
  AND2X2 AND2X2_5447 ( .A(u3_u0__abc_48231_n853_bF_buf4), .B(u3_u0__abc_48231_n509), .Y(u3_u0__abc_48231_n955) );
  AND2X2 AND2X2_5448 ( .A(u3_u0__abc_48231_n956), .B(u3_u0__abc_48231_n954), .Y(u3_u0_r0_25__FF_INPUT) );
  AND2X2 AND2X2_5449 ( .A(u3_u0__abc_48231_n853_bF_buf2), .B(u3_u0__abc_48231_n514_1), .Y(u3_u0__abc_48231_n959) );
  AND2X2 AND2X2_545 ( .A(spec_req_cs_4_bF_buf1), .B(u0_csc4_4_), .Y(u0__abc_49347_n2058) );
  AND2X2 AND2X2_5450 ( .A(u3_u0__abc_48231_n960), .B(u3_u0__abc_48231_n958), .Y(u3_u0_r0_26__FF_INPUT) );
  AND2X2 AND2X2_5451 ( .A(u3_u0__abc_48231_n853_bF_buf0), .B(u3_u0__abc_48231_n519), .Y(u3_u0__abc_48231_n963) );
  AND2X2 AND2X2_5452 ( .A(u3_u0__abc_48231_n964), .B(u3_u0__abc_48231_n962), .Y(u3_u0_r0_27__FF_INPUT) );
  AND2X2 AND2X2_5453 ( .A(u3_u0__abc_48231_n853_bF_buf6), .B(u3_u0__abc_48231_n524), .Y(u3_u0__abc_48231_n967) );
  AND2X2 AND2X2_5454 ( .A(u3_u0__abc_48231_n968), .B(u3_u0__abc_48231_n966), .Y(u3_u0_r0_28__FF_INPUT) );
  AND2X2 AND2X2_5455 ( .A(u3_u0__abc_48231_n853_bF_buf4), .B(u3_u0__abc_48231_n529), .Y(u3_u0__abc_48231_n971) );
  AND2X2 AND2X2_5456 ( .A(u3_u0__abc_48231_n972), .B(u3_u0__abc_48231_n970), .Y(u3_u0_r0_29__FF_INPUT) );
  AND2X2 AND2X2_5457 ( .A(u3_u0__abc_48231_n853_bF_buf2), .B(u3_u0__abc_48231_n534), .Y(u3_u0__abc_48231_n975) );
  AND2X2 AND2X2_5458 ( .A(u3_u0__abc_48231_n976), .B(u3_u0__abc_48231_n974), .Y(u3_u0_r0_30__FF_INPUT) );
  AND2X2 AND2X2_5459 ( .A(u3_u0__abc_48231_n853_bF_buf0), .B(u3_u0__abc_48231_n539), .Y(u3_u0__abc_48231_n979) );
  AND2X2 AND2X2_546 ( .A(u0__abc_49347_n2059), .B(u0__abc_49347_n1180_1_bF_buf4), .Y(u0__abc_49347_n2060) );
  AND2X2 AND2X2_5460 ( .A(u3_u0__abc_48231_n980), .B(u3_u0__abc_48231_n978), .Y(u3_u0_r0_31__FF_INPUT) );
  AND2X2 AND2X2_5461 ( .A(u3_u0__abc_48231_n853_bF_buf6), .B(u3_u0__abc_48231_n544), .Y(u3_u0__abc_48231_n983) );
  AND2X2 AND2X2_5462 ( .A(u3_u0__abc_48231_n984), .B(u3_u0__abc_48231_n982), .Y(u3_u0_r0_32__FF_INPUT) );
  AND2X2 AND2X2_5463 ( .A(u3_u0__abc_48231_n853_bF_buf4), .B(u3_u0__abc_48231_n549), .Y(u3_u0__abc_48231_n987) );
  AND2X2 AND2X2_5464 ( .A(u3_u0__abc_48231_n988), .B(u3_u0__abc_48231_n986), .Y(u3_u0_r0_33__FF_INPUT) );
  AND2X2 AND2X2_5465 ( .A(u3_u0__abc_48231_n853_bF_buf2), .B(u3_u0__abc_48231_n554), .Y(u3_u0__abc_48231_n991) );
  AND2X2 AND2X2_5466 ( .A(u3_u0__abc_48231_n992), .B(u3_u0__abc_48231_n990), .Y(u3_u0_r0_34__FF_INPUT) );
  AND2X2 AND2X2_5467 ( .A(u3_u0__abc_48231_n853_bF_buf0), .B(u3_u0__abc_48231_n559), .Y(u3_u0__abc_48231_n995) );
  AND2X2 AND2X2_5468 ( .A(u3_u0__abc_48231_n996), .B(u3_u0__abc_48231_n994), .Y(u3_u0_r0_35__FF_INPUT) );
  AND2X2 AND2X2_5469 ( .A(u3_u0__abc_48231_n998), .B(u3_u0_wr_adr_0_), .Y(u3_u0__abc_48231_n999) );
  AND2X2 AND2X2_547 ( .A(spec_req_cs_3_bF_buf1), .B(u0_csc3_4_), .Y(u0__abc_49347_n2061) );
  AND2X2 AND2X2_5470 ( .A(u3_u0__abc_48231_n998), .B(u3_u0_wr_adr_1_), .Y(u3_u0__abc_48231_n1003) );
  AND2X2 AND2X2_5471 ( .A(u3_u0__abc_48231_n1004), .B(u3_u0__abc_48231_n1002), .Y(u3_u0_wr_adr_1__FF_INPUT) );
  AND2X2 AND2X2_5472 ( .A(u3_u0__abc_48231_n998), .B(u3_u0_wr_adr_2_), .Y(u3_u0__abc_48231_n1006) );
  AND2X2 AND2X2_5473 ( .A(u3_u0__abc_48231_n1007), .B(u3_u0__abc_48231_n1002), .Y(u3_u0_wr_adr_2__FF_INPUT) );
  AND2X2 AND2X2_5474 ( .A(u3_u0__abc_48231_n998), .B(u3_u0_wr_adr_3_), .Y(u3_u0__abc_48231_n1009) );
  AND2X2 AND2X2_5475 ( .A(u3_u0__abc_48231_n1010), .B(u3_u0__abc_48231_n1002), .Y(u3_u0_wr_adr_3__FF_INPUT) );
  AND2X2 AND2X2_5476 ( .A(u3_u0__abc_48231_n1012), .B(u3_u0_rd_adr_0_), .Y(u3_u0__abc_48231_n1013) );
  AND2X2 AND2X2_5477 ( .A(u3_u0_rd_adr_3_), .B(u3_re), .Y(u3_u0__abc_48231_n1014) );
  AND2X2 AND2X2_5478 ( .A(u3_u0_rd_adr_0_), .B(u3_re), .Y(u3_u0__abc_48231_n1017) );
  AND2X2 AND2X2_5479 ( .A(u3_u0__abc_48231_n1012), .B(u3_u0_rd_adr_1_), .Y(u3_u0__abc_48231_n1018) );
  AND2X2 AND2X2_548 ( .A(u0__abc_49347_n2062), .B(u0__abc_49347_n1179_bF_buf4), .Y(u0__abc_49347_n2063) );
  AND2X2 AND2X2_5480 ( .A(u3_u0__abc_48231_n1019), .B(u3_u0__abc_48231_n1002), .Y(u3_u0_rd_adr_1__FF_INPUT) );
  AND2X2 AND2X2_5481 ( .A(u3_re), .B(u3_u0_rd_adr_1_), .Y(u3_u0__abc_48231_n1021) );
  AND2X2 AND2X2_5482 ( .A(u3_u0__abc_48231_n1012), .B(u3_u0_rd_adr_2_), .Y(u3_u0__abc_48231_n1022) );
  AND2X2 AND2X2_5483 ( .A(u3_u0__abc_48231_n1023), .B(u3_u0__abc_48231_n1002), .Y(u3_u0_rd_adr_2__FF_INPUT) );
  AND2X2 AND2X2_5484 ( .A(u3_re), .B(u3_u0_rd_adr_2_), .Y(u3_u0__abc_48231_n1025) );
  AND2X2 AND2X2_5485 ( .A(u3_u0__abc_48231_n1012), .B(u3_u0_rd_adr_3_), .Y(u3_u0__abc_48231_n1026) );
  AND2X2 AND2X2_5486 ( .A(u3_u0__abc_48231_n1027), .B(u3_u0__abc_48231_n1002), .Y(u3_u0_rd_adr_3__FF_INPUT) );
  AND2X2 AND2X2_5487 ( .A(u3_u0__abc_48231_n1029), .B(u3_u0__abc_48231_n1030), .Y(u3_u0__abc_48231_n1031) );
  AND2X2 AND2X2_5488 ( .A(u3_u0__abc_48231_n1032), .B(u3_u0_rd_adr_1_), .Y(u3_u0__abc_48231_n1033) );
  AND2X2 AND2X2_5489 ( .A(u3_u0__abc_48231_n1031), .B(u3_u0__abc_48231_n1033), .Y(u3_u0__abc_48231_n1034) );
  AND2X2 AND2X2_549 ( .A(spec_req_cs_2_bF_buf1), .B(u0_csc2_4_), .Y(u0__abc_49347_n2064) );
  AND2X2 AND2X2_5490 ( .A(u3_u0__abc_48231_n1038), .B(u3_u0__abc_48231_n1040), .Y(u3_u0__abc_48231_n1041) );
  AND2X2 AND2X2_5491 ( .A(u3_u0__abc_48231_n1041), .B(u3_u0__abc_48231_n1035), .Y(u3_u0__abc_48231_n1042) );
  AND2X2 AND2X2_5492 ( .A(u3_u0__abc_48231_n1042_bF_buf5), .B(u3_u0_r3_0_), .Y(u3_u0__abc_48231_n1043) );
  AND2X2 AND2X2_5493 ( .A(u3_u0__abc_48231_n1029), .B(u3_u0__abc_48231_n1044), .Y(u3_u0__abc_48231_n1045) );
  AND2X2 AND2X2_5494 ( .A(u3_u0__abc_48231_n1032), .B(u3_u0_rd_adr_2_), .Y(u3_u0__abc_48231_n1046) );
  AND2X2 AND2X2_5495 ( .A(u3_u0__abc_48231_n1045), .B(u3_u0__abc_48231_n1046), .Y(u3_u0__abc_48231_n1047) );
  AND2X2 AND2X2_5496 ( .A(u3_u0__abc_48231_n1047_bF_buf5), .B(u3_u0_r2_0_), .Y(u3_u0__abc_48231_n1048) );
  AND2X2 AND2X2_5497 ( .A(u3_u0__abc_48231_n1044), .B(u3_u0_rd_adr_0_), .Y(u3_u0__abc_48231_n1049) );
  AND2X2 AND2X2_5498 ( .A(u3_u0__abc_48231_n1031), .B(u3_u0__abc_48231_n1049), .Y(u3_u0__abc_48231_n1050) );
  AND2X2 AND2X2_5499 ( .A(u3_u0__abc_48231_n1050_bF_buf5), .B(u3_u0_r0_0_), .Y(u3_u0__abc_48231_n1051) );
  AND2X2 AND2X2_55 ( .A(wb_stb_i_bF_buf5), .B(wb_cyc_i), .Y(_abc_55805_n484) );
  AND2X2 AND2X2_550 ( .A(u0__abc_49347_n2065), .B(u0__abc_49347_n1178_1_bF_buf4), .Y(u0__abc_49347_n2066) );
  AND2X2 AND2X2_5500 ( .A(u3_u0__abc_48231_n1034_bF_buf4), .B(u3_u0_r1_0_), .Y(u3_u0__abc_48231_n1052) );
  AND2X2 AND2X2_5501 ( .A(u3_u0__abc_48231_n1042_bF_buf4), .B(u3_u0_r3_1_), .Y(u3_u0__abc_48231_n1056) );
  AND2X2 AND2X2_5502 ( .A(u3_u0__abc_48231_n1034_bF_buf3), .B(u3_u0_r1_1_), .Y(u3_u0__abc_48231_n1057) );
  AND2X2 AND2X2_5503 ( .A(u3_u0__abc_48231_n1050_bF_buf4), .B(u3_u0_r0_1_), .Y(u3_u0__abc_48231_n1058) );
  AND2X2 AND2X2_5504 ( .A(u3_u0__abc_48231_n1047_bF_buf4), .B(u3_u0_r2_1_), .Y(u3_u0__abc_48231_n1059) );
  AND2X2 AND2X2_5505 ( .A(u3_u0__abc_48231_n1042_bF_buf3), .B(u3_u0_r3_2_), .Y(u3_u0__abc_48231_n1063) );
  AND2X2 AND2X2_5506 ( .A(u3_u0__abc_48231_n1034_bF_buf2), .B(u3_u0_r1_2_), .Y(u3_u0__abc_48231_n1064) );
  AND2X2 AND2X2_5507 ( .A(u3_u0__abc_48231_n1050_bF_buf3), .B(u3_u0_r0_2_), .Y(u3_u0__abc_48231_n1065) );
  AND2X2 AND2X2_5508 ( .A(u3_u0__abc_48231_n1047_bF_buf3), .B(u3_u0_r2_2_), .Y(u3_u0__abc_48231_n1066) );
  AND2X2 AND2X2_5509 ( .A(u3_u0__abc_48231_n1042_bF_buf2), .B(u3_u0_r3_3_), .Y(u3_u0__abc_48231_n1070) );
  AND2X2 AND2X2_551 ( .A(spec_req_cs_1_bF_buf1), .B(u0_csc1_4_), .Y(u0__abc_49347_n2067) );
  AND2X2 AND2X2_5510 ( .A(u3_u0__abc_48231_n1034_bF_buf1), .B(u3_u0_r1_3_), .Y(u3_u0__abc_48231_n1071) );
  AND2X2 AND2X2_5511 ( .A(u3_u0__abc_48231_n1050_bF_buf2), .B(u3_u0_r0_3_), .Y(u3_u0__abc_48231_n1072) );
  AND2X2 AND2X2_5512 ( .A(u3_u0__abc_48231_n1047_bF_buf2), .B(u3_u0_r2_3_), .Y(u3_u0__abc_48231_n1073) );
  AND2X2 AND2X2_5513 ( .A(u3_u0__abc_48231_n1042_bF_buf1), .B(u3_u0_r3_4_), .Y(u3_u0__abc_48231_n1077) );
  AND2X2 AND2X2_5514 ( .A(u3_u0__abc_48231_n1047_bF_buf1), .B(u3_u0_r2_4_), .Y(u3_u0__abc_48231_n1078) );
  AND2X2 AND2X2_5515 ( .A(u3_u0__abc_48231_n1050_bF_buf1), .B(u3_u0_r0_4_), .Y(u3_u0__abc_48231_n1079) );
  AND2X2 AND2X2_5516 ( .A(u3_u0__abc_48231_n1034_bF_buf0), .B(u3_u0_r1_4_), .Y(u3_u0__abc_48231_n1080) );
  AND2X2 AND2X2_5517 ( .A(u3_u0__abc_48231_n1042_bF_buf0), .B(u3_u0_r3_5_), .Y(u3_u0__abc_48231_n1084) );
  AND2X2 AND2X2_5518 ( .A(u3_u0__abc_48231_n1034_bF_buf5), .B(u3_u0_r1_5_), .Y(u3_u0__abc_48231_n1085) );
  AND2X2 AND2X2_5519 ( .A(u3_u0__abc_48231_n1050_bF_buf0), .B(u3_u0_r0_5_), .Y(u3_u0__abc_48231_n1086) );
  AND2X2 AND2X2_552 ( .A(u0__abc_49347_n1952_1_bF_buf3), .B(u0__abc_49347_n2070), .Y(u0__abc_49347_n2071) );
  AND2X2 AND2X2_5520 ( .A(u3_u0__abc_48231_n1047_bF_buf0), .B(u3_u0_r2_5_), .Y(u3_u0__abc_48231_n1087) );
  AND2X2 AND2X2_5521 ( .A(u3_u0__abc_48231_n1042_bF_buf5), .B(u3_u0_r3_6_), .Y(u3_u0__abc_48231_n1091) );
  AND2X2 AND2X2_5522 ( .A(u3_u0__abc_48231_n1034_bF_buf4), .B(u3_u0_r1_6_), .Y(u3_u0__abc_48231_n1092) );
  AND2X2 AND2X2_5523 ( .A(u3_u0__abc_48231_n1050_bF_buf5), .B(u3_u0_r0_6_), .Y(u3_u0__abc_48231_n1093) );
  AND2X2 AND2X2_5524 ( .A(u3_u0__abc_48231_n1047_bF_buf5), .B(u3_u0_r2_6_), .Y(u3_u0__abc_48231_n1094) );
  AND2X2 AND2X2_5525 ( .A(u3_u0__abc_48231_n1042_bF_buf4), .B(u3_u0_r3_7_), .Y(u3_u0__abc_48231_n1098) );
  AND2X2 AND2X2_5526 ( .A(u3_u0__abc_48231_n1034_bF_buf3), .B(u3_u0_r1_7_), .Y(u3_u0__abc_48231_n1099) );
  AND2X2 AND2X2_5527 ( .A(u3_u0__abc_48231_n1050_bF_buf4), .B(u3_u0_r0_7_), .Y(u3_u0__abc_48231_n1100) );
  AND2X2 AND2X2_5528 ( .A(u3_u0__abc_48231_n1047_bF_buf4), .B(u3_u0_r2_7_), .Y(u3_u0__abc_48231_n1101) );
  AND2X2 AND2X2_5529 ( .A(u3_u0__abc_48231_n1042_bF_buf3), .B(u3_u0_r3_8_), .Y(u3_u0__abc_48231_n1105) );
  AND2X2 AND2X2_553 ( .A(u0__abc_49347_n2069), .B(u0__abc_49347_n2071), .Y(u0__abc_49347_n2072_1) );
  AND2X2 AND2X2_5530 ( .A(u3_u0__abc_48231_n1034_bF_buf2), .B(u3_u0_r1_8_), .Y(u3_u0__abc_48231_n1106) );
  AND2X2 AND2X2_5531 ( .A(u3_u0__abc_48231_n1050_bF_buf3), .B(u3_u0_r0_8_), .Y(u3_u0__abc_48231_n1107) );
  AND2X2 AND2X2_5532 ( .A(u3_u0__abc_48231_n1047_bF_buf3), .B(u3_u0_r2_8_), .Y(u3_u0__abc_48231_n1108) );
  AND2X2 AND2X2_5533 ( .A(u3_u0__abc_48231_n1042_bF_buf2), .B(u3_u0_r3_9_), .Y(u3_u0__abc_48231_n1112) );
  AND2X2 AND2X2_5534 ( .A(u3_u0__abc_48231_n1034_bF_buf1), .B(u3_u0_r1_9_), .Y(u3_u0__abc_48231_n1113) );
  AND2X2 AND2X2_5535 ( .A(u3_u0__abc_48231_n1050_bF_buf2), .B(u3_u0_r0_9_), .Y(u3_u0__abc_48231_n1114) );
  AND2X2 AND2X2_5536 ( .A(u3_u0__abc_48231_n1047_bF_buf2), .B(u3_u0_r2_9_), .Y(u3_u0__abc_48231_n1115) );
  AND2X2 AND2X2_5537 ( .A(u3_u0__abc_48231_n1042_bF_buf1), .B(u3_u0_r3_10_), .Y(u3_u0__abc_48231_n1119) );
  AND2X2 AND2X2_5538 ( .A(u3_u0__abc_48231_n1034_bF_buf0), .B(u3_u0_r1_10_), .Y(u3_u0__abc_48231_n1120) );
  AND2X2 AND2X2_5539 ( .A(u3_u0__abc_48231_n1050_bF_buf1), .B(u3_u0_r0_10_), .Y(u3_u0__abc_48231_n1121) );
  AND2X2 AND2X2_554 ( .A(u0__abc_49347_n1953_1_bF_buf3), .B(sp_csc_5_), .Y(u0__abc_49347_n2074) );
  AND2X2 AND2X2_5540 ( .A(u3_u0__abc_48231_n1047_bF_buf1), .B(u3_u0_r2_10_), .Y(u3_u0__abc_48231_n1122) );
  AND2X2 AND2X2_5541 ( .A(u3_u0__abc_48231_n1042_bF_buf0), .B(u3_u0_r3_11_), .Y(u3_u0__abc_48231_n1126) );
  AND2X2 AND2X2_5542 ( .A(u3_u0__abc_48231_n1034_bF_buf5), .B(u3_u0_r1_11_), .Y(u3_u0__abc_48231_n1127) );
  AND2X2 AND2X2_5543 ( .A(u3_u0__abc_48231_n1050_bF_buf0), .B(u3_u0_r0_11_), .Y(u3_u0__abc_48231_n1128) );
  AND2X2 AND2X2_5544 ( .A(u3_u0__abc_48231_n1047_bF_buf0), .B(u3_u0_r2_11_), .Y(u3_u0__abc_48231_n1129) );
  AND2X2 AND2X2_5545 ( .A(u3_u0__abc_48231_n1042_bF_buf5), .B(u3_u0_r3_12_), .Y(u3_u0__abc_48231_n1133) );
  AND2X2 AND2X2_5546 ( .A(u3_u0__abc_48231_n1047_bF_buf5), .B(u3_u0_r2_12_), .Y(u3_u0__abc_48231_n1134) );
  AND2X2 AND2X2_5547 ( .A(u3_u0__abc_48231_n1050_bF_buf5), .B(u3_u0_r0_12_), .Y(u3_u0__abc_48231_n1135) );
  AND2X2 AND2X2_5548 ( .A(u3_u0__abc_48231_n1034_bF_buf4), .B(u3_u0_r1_12_), .Y(u3_u0__abc_48231_n1136) );
  AND2X2 AND2X2_5549 ( .A(u3_u0__abc_48231_n1042_bF_buf4), .B(u3_u0_r3_13_), .Y(u3_u0__abc_48231_n1140) );
  AND2X2 AND2X2_555 ( .A(spec_req_cs_5_bF_buf0), .B(u0_csc5_5_), .Y(u0__abc_49347_n2075) );
  AND2X2 AND2X2_5550 ( .A(u3_u0__abc_48231_n1034_bF_buf3), .B(u3_u0_r1_13_), .Y(u3_u0__abc_48231_n1141) );
  AND2X2 AND2X2_5551 ( .A(u3_u0__abc_48231_n1050_bF_buf4), .B(u3_u0_r0_13_), .Y(u3_u0__abc_48231_n1142) );
  AND2X2 AND2X2_5552 ( .A(u3_u0__abc_48231_n1047_bF_buf4), .B(u3_u0_r2_13_), .Y(u3_u0__abc_48231_n1143) );
  AND2X2 AND2X2_5553 ( .A(u3_u0__abc_48231_n1042_bF_buf3), .B(u3_u0_r3_14_), .Y(u3_u0__abc_48231_n1147) );
  AND2X2 AND2X2_5554 ( .A(u3_u0__abc_48231_n1047_bF_buf3), .B(u3_u0_r2_14_), .Y(u3_u0__abc_48231_n1148) );
  AND2X2 AND2X2_5555 ( .A(u3_u0__abc_48231_n1050_bF_buf3), .B(u3_u0_r0_14_), .Y(u3_u0__abc_48231_n1149) );
  AND2X2 AND2X2_5556 ( .A(u3_u0__abc_48231_n1034_bF_buf2), .B(u3_u0_r1_14_), .Y(u3_u0__abc_48231_n1150) );
  AND2X2 AND2X2_5557 ( .A(u3_u0__abc_48231_n1042_bF_buf2), .B(u3_u0_r3_15_), .Y(u3_u0__abc_48231_n1154) );
  AND2X2 AND2X2_5558 ( .A(u3_u0__abc_48231_n1034_bF_buf1), .B(u3_u0_r1_15_), .Y(u3_u0__abc_48231_n1155) );
  AND2X2 AND2X2_5559 ( .A(u3_u0__abc_48231_n1050_bF_buf2), .B(u3_u0_r0_15_), .Y(u3_u0__abc_48231_n1156) );
  AND2X2 AND2X2_556 ( .A(u0__abc_49347_n2077), .B(u0__abc_49347_n1185_bF_buf3), .Y(u0__abc_49347_n2078) );
  AND2X2 AND2X2_5560 ( .A(u3_u0__abc_48231_n1047_bF_buf2), .B(u3_u0_r2_15_), .Y(u3_u0__abc_48231_n1157) );
  AND2X2 AND2X2_5561 ( .A(u3_u0__abc_48231_n1042_bF_buf1), .B(u3_u0_r3_16_), .Y(u3_u0__abc_48231_n1161) );
  AND2X2 AND2X2_5562 ( .A(u3_u0__abc_48231_n1034_bF_buf0), .B(u3_u0_r1_16_), .Y(u3_u0__abc_48231_n1162) );
  AND2X2 AND2X2_5563 ( .A(u3_u0__abc_48231_n1050_bF_buf1), .B(u3_u0_r0_16_), .Y(u3_u0__abc_48231_n1163) );
  AND2X2 AND2X2_5564 ( .A(u3_u0__abc_48231_n1047_bF_buf1), .B(u3_u0_r2_16_), .Y(u3_u0__abc_48231_n1164) );
  AND2X2 AND2X2_5565 ( .A(u3_u0__abc_48231_n1042_bF_buf0), .B(u3_u0_r3_17_), .Y(u3_u0__abc_48231_n1168) );
  AND2X2 AND2X2_5566 ( .A(u3_u0__abc_48231_n1034_bF_buf5), .B(u3_u0_r1_17_), .Y(u3_u0__abc_48231_n1169) );
  AND2X2 AND2X2_5567 ( .A(u3_u0__abc_48231_n1050_bF_buf0), .B(u3_u0_r0_17_), .Y(u3_u0__abc_48231_n1170) );
  AND2X2 AND2X2_5568 ( .A(u3_u0__abc_48231_n1047_bF_buf0), .B(u3_u0_r2_17_), .Y(u3_u0__abc_48231_n1171) );
  AND2X2 AND2X2_5569 ( .A(u3_u0__abc_48231_n1042_bF_buf5), .B(u3_u0_r3_18_), .Y(u3_u0__abc_48231_n1175) );
  AND2X2 AND2X2_557 ( .A(u0__abc_49347_n2078), .B(u0__abc_49347_n2076), .Y(u0__abc_49347_n2079) );
  AND2X2 AND2X2_5570 ( .A(u3_u0__abc_48231_n1034_bF_buf4), .B(u3_u0_r1_18_), .Y(u3_u0__abc_48231_n1176) );
  AND2X2 AND2X2_5571 ( .A(u3_u0__abc_48231_n1050_bF_buf5), .B(u3_u0_r0_18_), .Y(u3_u0__abc_48231_n1177) );
  AND2X2 AND2X2_5572 ( .A(u3_u0__abc_48231_n1047_bF_buf5), .B(u3_u0_r2_18_), .Y(u3_u0__abc_48231_n1178) );
  AND2X2 AND2X2_5573 ( .A(u3_u0__abc_48231_n1042_bF_buf4), .B(u3_u0_r3_19_), .Y(u3_u0__abc_48231_n1182) );
  AND2X2 AND2X2_5574 ( .A(u3_u0__abc_48231_n1034_bF_buf3), .B(u3_u0_r1_19_), .Y(u3_u0__abc_48231_n1183) );
  AND2X2 AND2X2_5575 ( .A(u3_u0__abc_48231_n1050_bF_buf4), .B(u3_u0_r0_19_), .Y(u3_u0__abc_48231_n1184) );
  AND2X2 AND2X2_5576 ( .A(u3_u0__abc_48231_n1047_bF_buf4), .B(u3_u0_r2_19_), .Y(u3_u0__abc_48231_n1185) );
  AND2X2 AND2X2_5577 ( .A(u3_u0__abc_48231_n1042_bF_buf3), .B(u3_u0_r3_20_), .Y(u3_u0__abc_48231_n1189) );
  AND2X2 AND2X2_5578 ( .A(u3_u0__abc_48231_n1047_bF_buf3), .B(u3_u0_r2_20_), .Y(u3_u0__abc_48231_n1190) );
  AND2X2 AND2X2_5579 ( .A(u3_u0__abc_48231_n1050_bF_buf3), .B(u3_u0_r0_20_), .Y(u3_u0__abc_48231_n1191) );
  AND2X2 AND2X2_558 ( .A(u0__abc_49347_n2080), .B(u0__abc_49347_n1181_bF_buf3), .Y(u0__abc_49347_n2081) );
  AND2X2 AND2X2_5580 ( .A(u3_u0__abc_48231_n1034_bF_buf2), .B(u3_u0_r1_20_), .Y(u3_u0__abc_48231_n1192) );
  AND2X2 AND2X2_5581 ( .A(u3_u0__abc_48231_n1042_bF_buf2), .B(u3_u0_r3_21_), .Y(u3_u0__abc_48231_n1196) );
  AND2X2 AND2X2_5582 ( .A(u3_u0__abc_48231_n1034_bF_buf1), .B(u3_u0_r1_21_), .Y(u3_u0__abc_48231_n1197) );
  AND2X2 AND2X2_5583 ( .A(u3_u0__abc_48231_n1050_bF_buf2), .B(u3_u0_r0_21_), .Y(u3_u0__abc_48231_n1198) );
  AND2X2 AND2X2_5584 ( .A(u3_u0__abc_48231_n1047_bF_buf2), .B(u3_u0_r2_21_), .Y(u3_u0__abc_48231_n1199) );
  AND2X2 AND2X2_5585 ( .A(u3_u0__abc_48231_n1042_bF_buf1), .B(u3_u0_r3_22_), .Y(u3_u0__abc_48231_n1203) );
  AND2X2 AND2X2_5586 ( .A(u3_u0__abc_48231_n1034_bF_buf0), .B(u3_u0_r1_22_), .Y(u3_u0__abc_48231_n1204) );
  AND2X2 AND2X2_5587 ( .A(u3_u0__abc_48231_n1050_bF_buf1), .B(u3_u0_r0_22_), .Y(u3_u0__abc_48231_n1205) );
  AND2X2 AND2X2_5588 ( .A(u3_u0__abc_48231_n1047_bF_buf1), .B(u3_u0_r2_22_), .Y(u3_u0__abc_48231_n1206) );
  AND2X2 AND2X2_5589 ( .A(u3_u0__abc_48231_n1042_bF_buf0), .B(u3_u0_r3_23_), .Y(u3_u0__abc_48231_n1210) );
  AND2X2 AND2X2_559 ( .A(spec_req_cs_4_bF_buf0), .B(u0_csc4_5_), .Y(u0__abc_49347_n2082) );
  AND2X2 AND2X2_5590 ( .A(u3_u0__abc_48231_n1034_bF_buf5), .B(u3_u0_r1_23_), .Y(u3_u0__abc_48231_n1211) );
  AND2X2 AND2X2_5591 ( .A(u3_u0__abc_48231_n1050_bF_buf0), .B(u3_u0_r0_23_), .Y(u3_u0__abc_48231_n1212) );
  AND2X2 AND2X2_5592 ( .A(u3_u0__abc_48231_n1047_bF_buf0), .B(u3_u0_r2_23_), .Y(u3_u0__abc_48231_n1213) );
  AND2X2 AND2X2_5593 ( .A(u3_u0__abc_48231_n1042_bF_buf5), .B(u3_u0_r3_24_), .Y(u3_u0__abc_48231_n1217) );
  AND2X2 AND2X2_5594 ( .A(u3_u0__abc_48231_n1047_bF_buf5), .B(u3_u0_r2_24_), .Y(u3_u0__abc_48231_n1218) );
  AND2X2 AND2X2_5595 ( .A(u3_u0__abc_48231_n1050_bF_buf5), .B(u3_u0_r0_24_), .Y(u3_u0__abc_48231_n1219) );
  AND2X2 AND2X2_5596 ( .A(u3_u0__abc_48231_n1034_bF_buf4), .B(u3_u0_r1_24_), .Y(u3_u0__abc_48231_n1220) );
  AND2X2 AND2X2_5597 ( .A(u3_u0__abc_48231_n1042_bF_buf4), .B(u3_u0_r3_25_), .Y(u3_u0__abc_48231_n1224) );
  AND2X2 AND2X2_5598 ( .A(u3_u0__abc_48231_n1034_bF_buf3), .B(u3_u0_r1_25_), .Y(u3_u0__abc_48231_n1225) );
  AND2X2 AND2X2_5599 ( .A(u3_u0__abc_48231_n1050_bF_buf4), .B(u3_u0_r0_25_), .Y(u3_u0__abc_48231_n1226) );
  AND2X2 AND2X2_56 ( .A(_abc_55805_n483), .B(_abc_55805_n484), .Y(not_mem_cyc) );
  AND2X2 AND2X2_560 ( .A(u0__abc_49347_n2083), .B(u0__abc_49347_n1180_1_bF_buf3), .Y(u0__abc_49347_n2084) );
  AND2X2 AND2X2_5600 ( .A(u3_u0__abc_48231_n1047_bF_buf4), .B(u3_u0_r2_25_), .Y(u3_u0__abc_48231_n1227) );
  AND2X2 AND2X2_5601 ( .A(u3_u0__abc_48231_n1042_bF_buf3), .B(u3_u0_r3_26_), .Y(u3_u0__abc_48231_n1231) );
  AND2X2 AND2X2_5602 ( .A(u3_u0__abc_48231_n1034_bF_buf2), .B(u3_u0_r1_26_), .Y(u3_u0__abc_48231_n1232) );
  AND2X2 AND2X2_5603 ( .A(u3_u0__abc_48231_n1050_bF_buf3), .B(u3_u0_r0_26_), .Y(u3_u0__abc_48231_n1233) );
  AND2X2 AND2X2_5604 ( .A(u3_u0__abc_48231_n1047_bF_buf3), .B(u3_u0_r2_26_), .Y(u3_u0__abc_48231_n1234) );
  AND2X2 AND2X2_5605 ( .A(u3_u0__abc_48231_n1042_bF_buf2), .B(u3_u0_r3_27_), .Y(u3_u0__abc_48231_n1238) );
  AND2X2 AND2X2_5606 ( .A(u3_u0__abc_48231_n1034_bF_buf1), .B(u3_u0_r1_27_), .Y(u3_u0__abc_48231_n1239) );
  AND2X2 AND2X2_5607 ( .A(u3_u0__abc_48231_n1050_bF_buf2), .B(u3_u0_r0_27_), .Y(u3_u0__abc_48231_n1240) );
  AND2X2 AND2X2_5608 ( .A(u3_u0__abc_48231_n1047_bF_buf2), .B(u3_u0_r2_27_), .Y(u3_u0__abc_48231_n1241) );
  AND2X2 AND2X2_5609 ( .A(u3_u0__abc_48231_n1042_bF_buf1), .B(u3_u0_r3_28_), .Y(u3_u0__abc_48231_n1245) );
  AND2X2 AND2X2_561 ( .A(spec_req_cs_3_bF_buf0), .B(u0_csc3_5_), .Y(u0__abc_49347_n2085) );
  AND2X2 AND2X2_5610 ( .A(u3_u0__abc_48231_n1034_bF_buf0), .B(u3_u0_r1_28_), .Y(u3_u0__abc_48231_n1246) );
  AND2X2 AND2X2_5611 ( .A(u3_u0__abc_48231_n1050_bF_buf1), .B(u3_u0_r0_28_), .Y(u3_u0__abc_48231_n1247) );
  AND2X2 AND2X2_5612 ( .A(u3_u0__abc_48231_n1047_bF_buf1), .B(u3_u0_r2_28_), .Y(u3_u0__abc_48231_n1248) );
  AND2X2 AND2X2_5613 ( .A(u3_u0__abc_48231_n1042_bF_buf0), .B(u3_u0_r3_29_), .Y(u3_u0__abc_48231_n1252) );
  AND2X2 AND2X2_5614 ( .A(u3_u0__abc_48231_n1034_bF_buf5), .B(u3_u0_r1_29_), .Y(u3_u0__abc_48231_n1253) );
  AND2X2 AND2X2_5615 ( .A(u3_u0__abc_48231_n1050_bF_buf0), .B(u3_u0_r0_29_), .Y(u3_u0__abc_48231_n1254) );
  AND2X2 AND2X2_5616 ( .A(u3_u0__abc_48231_n1047_bF_buf0), .B(u3_u0_r2_29_), .Y(u3_u0__abc_48231_n1255) );
  AND2X2 AND2X2_5617 ( .A(u3_u0__abc_48231_n1042_bF_buf5), .B(u3_u0_r3_30_), .Y(u3_u0__abc_48231_n1259) );
  AND2X2 AND2X2_5618 ( .A(u3_u0__abc_48231_n1034_bF_buf4), .B(u3_u0_r1_30_), .Y(u3_u0__abc_48231_n1260) );
  AND2X2 AND2X2_5619 ( .A(u3_u0__abc_48231_n1050_bF_buf5), .B(u3_u0_r0_30_), .Y(u3_u0__abc_48231_n1261) );
  AND2X2 AND2X2_562 ( .A(u0__abc_49347_n2086), .B(u0__abc_49347_n1179_bF_buf3), .Y(u0__abc_49347_n2087) );
  AND2X2 AND2X2_5620 ( .A(u3_u0__abc_48231_n1047_bF_buf5), .B(u3_u0_r2_30_), .Y(u3_u0__abc_48231_n1262) );
  AND2X2 AND2X2_5621 ( .A(u3_u0__abc_48231_n1042_bF_buf4), .B(u3_u0_r3_31_), .Y(u3_u0__abc_48231_n1266) );
  AND2X2 AND2X2_5622 ( .A(u3_u0__abc_48231_n1034_bF_buf3), .B(u3_u0_r1_31_), .Y(u3_u0__abc_48231_n1267) );
  AND2X2 AND2X2_5623 ( .A(u3_u0__abc_48231_n1050_bF_buf4), .B(u3_u0_r0_31_), .Y(u3_u0__abc_48231_n1268) );
  AND2X2 AND2X2_5624 ( .A(u3_u0__abc_48231_n1047_bF_buf4), .B(u3_u0_r2_31_), .Y(u3_u0__abc_48231_n1269) );
  AND2X2 AND2X2_5625 ( .A(u3_u0__abc_48231_n1042_bF_buf3), .B(u3_u0_r3_32_), .Y(u3_u0__abc_48231_n1273) );
  AND2X2 AND2X2_5626 ( .A(u3_u0__abc_48231_n1034_bF_buf2), .B(u3_u0_r1_32_), .Y(u3_u0__abc_48231_n1274) );
  AND2X2 AND2X2_5627 ( .A(u3_u0__abc_48231_n1050_bF_buf3), .B(u3_u0_r0_32_), .Y(u3_u0__abc_48231_n1275) );
  AND2X2 AND2X2_5628 ( .A(u3_u0__abc_48231_n1047_bF_buf3), .B(u3_u0_r2_32_), .Y(u3_u0__abc_48231_n1276) );
  AND2X2 AND2X2_5629 ( .A(u3_u0__abc_48231_n1042_bF_buf2), .B(u3_u0_r3_33_), .Y(u3_u0__abc_48231_n1280) );
  AND2X2 AND2X2_563 ( .A(spec_req_cs_2_bF_buf0), .B(u0_csc2_5_), .Y(u0__abc_49347_n2088) );
  AND2X2 AND2X2_5630 ( .A(u3_u0__abc_48231_n1034_bF_buf1), .B(u3_u0_r1_33_), .Y(u3_u0__abc_48231_n1281) );
  AND2X2 AND2X2_5631 ( .A(u3_u0__abc_48231_n1050_bF_buf2), .B(u3_u0_r0_33_), .Y(u3_u0__abc_48231_n1282) );
  AND2X2 AND2X2_5632 ( .A(u3_u0__abc_48231_n1047_bF_buf2), .B(u3_u0_r2_33_), .Y(u3_u0__abc_48231_n1283) );
  AND2X2 AND2X2_5633 ( .A(u3_u0__abc_48231_n1042_bF_buf1), .B(u3_u0_r3_34_), .Y(u3_u0__abc_48231_n1287) );
  AND2X2 AND2X2_5634 ( .A(u3_u0__abc_48231_n1034_bF_buf0), .B(u3_u0_r1_34_), .Y(u3_u0__abc_48231_n1288) );
  AND2X2 AND2X2_5635 ( .A(u3_u0__abc_48231_n1050_bF_buf1), .B(u3_u0_r0_34_), .Y(u3_u0__abc_48231_n1289) );
  AND2X2 AND2X2_5636 ( .A(u3_u0__abc_48231_n1047_bF_buf1), .B(u3_u0_r2_34_), .Y(u3_u0__abc_48231_n1290) );
  AND2X2 AND2X2_5637 ( .A(u3_u0__abc_48231_n1042_bF_buf0), .B(u3_u0_r3_35_), .Y(u3_u0__abc_48231_n1294) );
  AND2X2 AND2X2_5638 ( .A(u3_u0__abc_48231_n1034_bF_buf5), .B(u3_u0_r1_35_), .Y(u3_u0__abc_48231_n1295) );
  AND2X2 AND2X2_5639 ( .A(u3_u0__abc_48231_n1050_bF_buf0), .B(u3_u0_r0_35_), .Y(u3_u0__abc_48231_n1296) );
  AND2X2 AND2X2_564 ( .A(u0__abc_49347_n2089), .B(u0__abc_49347_n1178_1_bF_buf3), .Y(u0__abc_49347_n2090) );
  AND2X2 AND2X2_5640 ( .A(u3_u0__abc_48231_n1047_bF_buf0), .B(u3_u0_r2_35_), .Y(u3_u0__abc_48231_n1297) );
  AND2X2 AND2X2_5641 ( .A(u4__abc_49152_n72), .B(u4_ps_cnt_5_), .Y(u4__abc_49152_n73_1) );
  AND2X2 AND2X2_5642 ( .A(u4__abc_49152_n74), .B(rfr_ps_val_5_), .Y(u4__abc_49152_n75) );
  AND2X2 AND2X2_5643 ( .A(u4__abc_49152_n77), .B(u4_ps_cnt_4_), .Y(u4__abc_49152_n78) );
  AND2X2 AND2X2_5644 ( .A(u4__abc_49152_n79_1), .B(rfr_ps_val_4_), .Y(u4__abc_49152_n80) );
  AND2X2 AND2X2_5645 ( .A(u4__abc_49152_n83), .B(u4_ps_cnt_6_), .Y(u4__abc_49152_n84) );
  AND2X2 AND2X2_5646 ( .A(u4__abc_49152_n85_1), .B(rfr_ps_val_6_), .Y(u4__abc_49152_n86) );
  AND2X2 AND2X2_5647 ( .A(u4__abc_49152_n88_1), .B(u4_ps_cnt_7_), .Y(u4__abc_49152_n89) );
  AND2X2 AND2X2_5648 ( .A(u4__abc_49152_n90_1), .B(rfr_ps_val_7_), .Y(u4__abc_49152_n91) );
  AND2X2 AND2X2_5649 ( .A(u4__abc_49152_n95), .B(u4_ps_cnt_0_), .Y(u4__abc_49152_n96) );
  AND2X2 AND2X2_565 ( .A(spec_req_cs_1_bF_buf0), .B(u0_csc1_5_), .Y(u0__abc_49347_n2091) );
  AND2X2 AND2X2_5650 ( .A(u4__abc_49152_n97), .B(rfr_ps_val_0_), .Y(u4__abc_49152_n98) );
  AND2X2 AND2X2_5651 ( .A(u4__abc_49152_n100), .B(u4_ps_cnt_1_), .Y(u4__abc_49152_n101_1) );
  AND2X2 AND2X2_5652 ( .A(u4__abc_49152_n102_1), .B(rfr_ps_val_1_), .Y(u4__abc_49152_n103) );
  AND2X2 AND2X2_5653 ( .A(u4__abc_49152_n106), .B(u4_ps_cnt_2_), .Y(u4__abc_49152_n107) );
  AND2X2 AND2X2_5654 ( .A(u4__abc_49152_n108_1), .B(rfr_ps_val_2_), .Y(u4__abc_49152_n109) );
  AND2X2 AND2X2_5655 ( .A(u4_ps_cnt_3_), .B(rfr_ps_val_3_), .Y(u4__abc_49152_n112) );
  AND2X2 AND2X2_5656 ( .A(u4__abc_49152_n113_1), .B(u4__abc_49152_n111), .Y(u4__abc_49152_n114) );
  AND2X2 AND2X2_5657 ( .A(u4__abc_49152_n120), .B(u4__abc_49152_n119), .Y(u4_rfr_req_FF_INPUT) );
  AND2X2 AND2X2_5658 ( .A(u4_rfr_ce), .B(u4_rfr_cnt_0_), .Y(u4__abc_49152_n122) );
  AND2X2 AND2X2_5659 ( .A(u4__abc_49152_n124_1), .B(u4__abc_49152_n119), .Y(u4__abc_49152_n125) );
  AND2X2 AND2X2_566 ( .A(u0__abc_49347_n1952_1_bF_buf2), .B(u0__abc_49347_n2094), .Y(u0__abc_49347_n2095) );
  AND2X2 AND2X2_5660 ( .A(u4__abc_49152_n125), .B(u4__abc_49152_n123), .Y(u4_rfr_cnt_0__FF_INPUT) );
  AND2X2 AND2X2_5661 ( .A(u4_rfr_cnt_0_), .B(u4_rfr_cnt_1_), .Y(u4__abc_49152_n127) );
  AND2X2 AND2X2_5662 ( .A(u4__abc_49152_n127), .B(u4_rfr_ce), .Y(u4__abc_49152_n128) );
  AND2X2 AND2X2_5663 ( .A(u4__abc_49152_n130), .B(u4__abc_49152_n119), .Y(u4__abc_49152_n131) );
  AND2X2 AND2X2_5664 ( .A(u4__abc_49152_n131), .B(u4__abc_49152_n129_1), .Y(u4_rfr_cnt_1__FF_INPUT) );
  AND2X2 AND2X2_5665 ( .A(u4_rfr_cnt_1_), .B(u4_rfr_cnt_2_), .Y(u4__abc_49152_n134_1) );
  AND2X2 AND2X2_5666 ( .A(u4__abc_49152_n122), .B(u4__abc_49152_n134_1), .Y(u4__abc_49152_n135) );
  AND2X2 AND2X2_5667 ( .A(u4__abc_49152_n136), .B(u4__abc_49152_n119), .Y(u4__abc_49152_n137) );
  AND2X2 AND2X2_5668 ( .A(u4__abc_49152_n137), .B(u4__abc_49152_n133), .Y(u4_rfr_cnt_2__FF_INPUT) );
  AND2X2 AND2X2_5669 ( .A(u4_rfr_cnt_2_), .B(u4_rfr_cnt_3_), .Y(u4__abc_49152_n139_1) );
  AND2X2 AND2X2_567 ( .A(u0__abc_49347_n2093), .B(u0__abc_49347_n2095), .Y(u0__abc_49347_n2096) );
  AND2X2 AND2X2_5670 ( .A(u4__abc_49152_n128), .B(u4__abc_49152_n139_1), .Y(u4__abc_49152_n140) );
  AND2X2 AND2X2_5671 ( .A(u4__abc_49152_n142), .B(u4__abc_49152_n119), .Y(u4__abc_49152_n143_1) );
  AND2X2 AND2X2_5672 ( .A(u4__abc_49152_n143_1), .B(u4__abc_49152_n141_1), .Y(u4_rfr_cnt_3__FF_INPUT) );
  AND2X2 AND2X2_5673 ( .A(u4__abc_49152_n140), .B(u4_rfr_cnt_4_), .Y(u4__abc_49152_n145) );
  AND2X2 AND2X2_5674 ( .A(u4__abc_49152_n147), .B(u4__abc_49152_n119), .Y(u4__abc_49152_n148) );
  AND2X2 AND2X2_5675 ( .A(u4__abc_49152_n148), .B(u4__abc_49152_n146), .Y(u4_rfr_cnt_4__FF_INPUT) );
  AND2X2 AND2X2_5676 ( .A(u4_rfr_cnt_4_), .B(u4_rfr_cnt_5_), .Y(u4__abc_49152_n151) );
  AND2X2 AND2X2_5677 ( .A(u4__abc_49152_n140), .B(u4__abc_49152_n151), .Y(u4__abc_49152_n152) );
  AND2X2 AND2X2_5678 ( .A(u4__abc_49152_n153), .B(u4__abc_49152_n119), .Y(u4__abc_49152_n154) );
  AND2X2 AND2X2_5679 ( .A(u4__abc_49152_n154), .B(u4__abc_49152_n150), .Y(u4_rfr_cnt_5__FF_INPUT) );
  AND2X2 AND2X2_568 ( .A(u0__abc_49347_n1953_1_bF_buf2), .B(sp_csc_6_), .Y(u0__abc_49347_n2098) );
  AND2X2 AND2X2_5680 ( .A(u4__abc_49152_n152), .B(u4_rfr_cnt_6_), .Y(u4__abc_49152_n156) );
  AND2X2 AND2X2_5681 ( .A(u4__abc_49152_n158), .B(u4__abc_49152_n119), .Y(u4__abc_49152_n159_1) );
  AND2X2 AND2X2_5682 ( .A(u4__abc_49152_n159_1), .B(u4__abc_49152_n157), .Y(u4_rfr_cnt_6__FF_INPUT) );
  AND2X2 AND2X2_5683 ( .A(u4_rfr_cnt_6_), .B(u4_rfr_cnt_7_), .Y(u4__abc_49152_n162) );
  AND2X2 AND2X2_5684 ( .A(u4__abc_49152_n152), .B(u4__abc_49152_n162), .Y(u4__abc_49152_n163) );
  AND2X2 AND2X2_5685 ( .A(u4__abc_49152_n164), .B(u4__abc_49152_n119), .Y(u4__abc_49152_n165) );
  AND2X2 AND2X2_5686 ( .A(u4__abc_49152_n165), .B(u4__abc_49152_n161), .Y(u4_rfr_cnt_7__FF_INPUT) );
  AND2X2 AND2X2_5687 ( .A(u4__abc_49152_n83), .B(u4__abc_49152_n88_1), .Y(u4__abc_49152_n167) );
  AND2X2 AND2X2_5688 ( .A(u4__abc_49152_n77), .B(u4__abc_49152_n72), .Y(u4__abc_49152_n168) );
  AND2X2 AND2X2_5689 ( .A(u4__abc_49152_n167), .B(u4__abc_49152_n168), .Y(u4__abc_49152_n169) );
  AND2X2 AND2X2_569 ( .A(spec_req_cs_5_bF_buf5), .B(u0_csc5_6_), .Y(u0__abc_49347_n2099) );
  AND2X2 AND2X2_5690 ( .A(u4__abc_49152_n106), .B(u4__abc_49152_n170), .Y(u4__abc_49152_n171) );
  AND2X2 AND2X2_5691 ( .A(u4__abc_49152_n95), .B(u4__abc_49152_n100), .Y(u4__abc_49152_n172) );
  AND2X2 AND2X2_5692 ( .A(u4__abc_49152_n171), .B(u4__abc_49152_n172), .Y(u4__abc_49152_n173) );
  AND2X2 AND2X2_5693 ( .A(u4__abc_49152_n169), .B(u4__abc_49152_n173), .Y(u4__abc_49152_n174) );
  AND2X2 AND2X2_5694 ( .A(u4_ps_cnt_0_), .B(u4_rfr_en), .Y(u4__abc_49152_n178) );
  AND2X2 AND2X2_5695 ( .A(u4__abc_49152_n179), .B(u4__abc_49152_n177), .Y(u4__abc_49152_n180) );
  AND2X2 AND2X2_5696 ( .A(u4__abc_49152_n175), .B(u4__abc_49152_n180), .Y(u4_ps_cnt_0__FF_INPUT) );
  AND2X2 AND2X2_5697 ( .A(u4__abc_49152_n178), .B(u4_ps_cnt_1_), .Y(u4__abc_49152_n183) );
  AND2X2 AND2X2_5698 ( .A(u4__abc_49152_n184), .B(u4__abc_49152_n182), .Y(u4__abc_49152_n185) );
  AND2X2 AND2X2_5699 ( .A(u4__abc_49152_n175), .B(u4__abc_49152_n185), .Y(u4_ps_cnt_1__FF_INPUT) );
  AND2X2 AND2X2_57 ( .A(u0__abc_49347_n1100_1), .B(u0_lmr_req0), .Y(u0__abc_49347_n1101_1) );
  AND2X2 AND2X2_570 ( .A(u0__abc_49347_n2101), .B(u0__abc_49347_n1185_bF_buf2), .Y(u0__abc_49347_n2102) );
  AND2X2 AND2X2_5700 ( .A(u4__abc_49152_n184), .B(u4_ps_cnt_2_), .Y(u4__abc_49152_n187) );
  AND2X2 AND2X2_5701 ( .A(u4__abc_49152_n183), .B(u4__abc_49152_n108_1), .Y(u4__abc_49152_n188) );
  AND2X2 AND2X2_5702 ( .A(u4__abc_49152_n175), .B(u4__abc_49152_n189_1), .Y(u4_ps_cnt_2__FF_INPUT) );
  AND2X2 AND2X2_5703 ( .A(u4_ps_cnt_2_), .B(u4_ps_cnt_1_), .Y(u4__abc_49152_n191_1) );
  AND2X2 AND2X2_5704 ( .A(u4__abc_49152_n178), .B(u4__abc_49152_n191_1), .Y(u4__abc_49152_n192) );
  AND2X2 AND2X2_5705 ( .A(u4__abc_49152_n192), .B(u4_ps_cnt_3_), .Y(u4__abc_49152_n194) );
  AND2X2 AND2X2_5706 ( .A(u4__abc_49152_n195), .B(u4__abc_49152_n193), .Y(u4__abc_49152_n196) );
  AND2X2 AND2X2_5707 ( .A(u4__abc_49152_n175), .B(u4__abc_49152_n196), .Y(u4_ps_cnt_3__FF_INPUT) );
  AND2X2 AND2X2_5708 ( .A(u4_ps_cnt_3_), .B(u4_ps_cnt_4_), .Y(u4__abc_49152_n199) );
  AND2X2 AND2X2_5709 ( .A(u4__abc_49152_n192), .B(u4__abc_49152_n199), .Y(u4__abc_49152_n200) );
  AND2X2 AND2X2_571 ( .A(u0__abc_49347_n2102), .B(u0__abc_49347_n2100), .Y(u0__abc_49347_n2103) );
  AND2X2 AND2X2_5710 ( .A(u4__abc_49152_n198), .B(u4__abc_49152_n201), .Y(u4__abc_49152_n202) );
  AND2X2 AND2X2_5711 ( .A(u4__abc_49152_n175), .B(u4__abc_49152_n202), .Y(u4_ps_cnt_4__FF_INPUT) );
  AND2X2 AND2X2_5712 ( .A(u4__abc_49152_n200), .B(u4_ps_cnt_5_), .Y(u4__abc_49152_n205) );
  AND2X2 AND2X2_5713 ( .A(u4__abc_49152_n206), .B(u4__abc_49152_n204), .Y(u4__abc_49152_n207) );
  AND2X2 AND2X2_5714 ( .A(u4__abc_49152_n175), .B(u4__abc_49152_n207), .Y(u4_ps_cnt_5__FF_INPUT) );
  AND2X2 AND2X2_5715 ( .A(u4__abc_49152_n191_1), .B(u4_ps_cnt_0_), .Y(u4__abc_49152_n210) );
  AND2X2 AND2X2_5716 ( .A(u4_ps_cnt_4_), .B(u4_ps_cnt_5_), .Y(u4__abc_49152_n211) );
  AND2X2 AND2X2_5717 ( .A(u4__abc_49152_n211), .B(u4_ps_cnt_3_), .Y(u4__abc_49152_n212) );
  AND2X2 AND2X2_5718 ( .A(u4__abc_49152_n210), .B(u4__abc_49152_n212), .Y(u4__abc_49152_n213) );
  AND2X2 AND2X2_5719 ( .A(u4__abc_49152_n213), .B(u4_rfr_en), .Y(u4__abc_49152_n214) );
  AND2X2 AND2X2_572 ( .A(u0__abc_49347_n2104), .B(u0__abc_49347_n1181_bF_buf2), .Y(u0__abc_49347_n2105) );
  AND2X2 AND2X2_5720 ( .A(u4__abc_49152_n214), .B(u4_ps_cnt_6_), .Y(u4__abc_49152_n215) );
  AND2X2 AND2X2_5721 ( .A(u4__abc_49152_n216), .B(u4__abc_49152_n209), .Y(u4__abc_49152_n217) );
  AND2X2 AND2X2_5722 ( .A(u4__abc_49152_n175), .B(u4__abc_49152_n217), .Y(u4_ps_cnt_6__FF_INPUT) );
  AND2X2 AND2X2_5723 ( .A(u4__abc_49152_n215), .B(u4_ps_cnt_7_), .Y(u4__abc_49152_n219) );
  AND2X2 AND2X2_5724 ( .A(u4__abc_49152_n220), .B(u4__abc_49152_n221), .Y(u4__abc_49152_n222) );
  AND2X2 AND2X2_5725 ( .A(u4__abc_49152_n222), .B(u4__abc_49152_n175), .Y(u4_ps_cnt_7__FF_INPUT) );
  AND2X2 AND2X2_5726 ( .A(u4__abc_49152_n127), .B(u4_rfr_early), .Y(u4__abc_49152_n224) );
  AND2X2 AND2X2_5727 ( .A(u4__abc_49152_n224), .B(u4__abc_49152_n139_1), .Y(u4__abc_49152_n225) );
  AND2X2 AND2X2_5728 ( .A(ref_int_0_), .B(ref_int_1_), .Y(u4__abc_49152_n226) );
  AND2X2 AND2X2_5729 ( .A(u4__abc_49152_n225), .B(u4__abc_49152_n226), .Y(u4__abc_49152_n227) );
  AND2X2 AND2X2_573 ( .A(spec_req_cs_4_bF_buf5), .B(u0_csc4_6_), .Y(u0__abc_49347_n2106) );
  AND2X2 AND2X2_5730 ( .A(u4__abc_49152_n228), .B(u4_rfr_early), .Y(u4__abc_49152_n229) );
  AND2X2 AND2X2_5731 ( .A(u4_rfr_cnt_2_), .B(ref_int_1_), .Y(u4__abc_49152_n230) );
  AND2X2 AND2X2_5732 ( .A(u4__abc_49152_n127), .B(u4__abc_49152_n230), .Y(u4__abc_49152_n231) );
  AND2X2 AND2X2_5733 ( .A(u4__abc_49152_n231), .B(u4__abc_49152_n229), .Y(u4__abc_49152_n232) );
  AND2X2 AND2X2_5734 ( .A(u4__abc_49152_n234), .B(ref_int_0_), .Y(u4__abc_49152_n235) );
  AND2X2 AND2X2_5735 ( .A(u4__abc_49152_n224), .B(u4__abc_49152_n235), .Y(u4__abc_49152_n236) );
  AND2X2 AND2X2_5736 ( .A(u4__abc_49152_n234), .B(u4_rfr_cnt_0_), .Y(u4__abc_49152_n237) );
  AND2X2 AND2X2_5737 ( .A(u4__abc_49152_n229), .B(u4__abc_49152_n237), .Y(u4__abc_49152_n238) );
  AND2X2 AND2X2_5738 ( .A(u4__abc_49152_n151), .B(ref_int_0_), .Y(u4__abc_49152_n243) );
  AND2X2 AND2X2_5739 ( .A(u4__abc_49152_n242), .B(u4__abc_49152_n243), .Y(u4__abc_49152_n244) );
  AND2X2 AND2X2_574 ( .A(u0__abc_49347_n2107), .B(u0__abc_49347_n1180_1_bF_buf2), .Y(u0__abc_49347_n2108_1) );
  AND2X2 AND2X2_5740 ( .A(u4__abc_49152_n244), .B(u4__abc_49152_n225), .Y(u4__abc_49152_n245) );
  AND2X2 AND2X2_5741 ( .A(u4_rfr_cnt_3_), .B(u4_rfr_cnt_4_), .Y(u4__abc_49152_n247) );
  AND2X2 AND2X2_5742 ( .A(u4__abc_49152_n134_1), .B(u4__abc_49152_n247), .Y(u4__abc_49152_n248) );
  AND2X2 AND2X2_5743 ( .A(u4__abc_49152_n238), .B(u4__abc_49152_n248), .Y(u4__abc_49152_n249) );
  AND2X2 AND2X2_5744 ( .A(u4__abc_49152_n241), .B(u4__abc_49152_n251), .Y(u4__abc_49152_n252) );
  AND2X2 AND2X2_5745 ( .A(u4_rfr_cnt_5_), .B(u4_rfr_cnt_6_), .Y(u4__abc_49152_n253) );
  AND2X2 AND2X2_5746 ( .A(u4__abc_49152_n253), .B(ref_int_2_), .Y(u4__abc_49152_n254) );
  AND2X2 AND2X2_5747 ( .A(u4__abc_49152_n254), .B(u4__abc_49152_n247), .Y(u4__abc_49152_n255) );
  AND2X2 AND2X2_5748 ( .A(u4__abc_49152_n232), .B(u4__abc_49152_n255), .Y(u4__abc_49152_n256) );
  AND2X2 AND2X2_5749 ( .A(u5__abc_54027_n253_1), .B(u5__abc_54027_n249_1), .Y(u5__abc_54027_n254) );
  AND2X2 AND2X2_575 ( .A(spec_req_cs_3_bF_buf5), .B(u0_csc3_6_), .Y(u0__abc_49347_n2109) );
  AND2X2 AND2X2_5750 ( .A(u5__abc_54027_n254), .B(u5__abc_54027_n248_1), .Y(u5__abc_54027_n255_1) );
  AND2X2 AND2X2_5751 ( .A(u5__abc_54027_n257), .B(u5__abc_54027_n258), .Y(u5__abc_54027_n259_1) );
  AND2X2 AND2X2_5752 ( .A(u5__abc_54027_n260_1), .B(u5__abc_54027_n261), .Y(u5__abc_54027_n262) );
  AND2X2 AND2X2_5753 ( .A(u5__abc_54027_n259_1), .B(u5__abc_54027_n262), .Y(u5__abc_54027_n263) );
  AND2X2 AND2X2_5754 ( .A(u5__abc_54027_n263), .B(u5__abc_54027_n256_1), .Y(u5__abc_54027_n264_1) );
  AND2X2 AND2X2_5755 ( .A(u5__abc_54027_n255_1), .B(u5__abc_54027_n264_1), .Y(u5__abc_54027_n265) );
  AND2X2 AND2X2_5756 ( .A(u5__abc_54027_n268_1), .B(u5_state_4_), .Y(u5__abc_54027_n269) );
  AND2X2 AND2X2_5757 ( .A(u5__abc_54027_n269), .B(u5__abc_54027_n267), .Y(u5__abc_54027_n270) );
  AND2X2 AND2X2_5758 ( .A(u5__abc_54027_n271), .B(u5_state_2_), .Y(u5__abc_54027_n272) );
  AND2X2 AND2X2_5759 ( .A(u5_state_0_), .B(u5_state_1_), .Y(u5__abc_54027_n273) );
  AND2X2 AND2X2_576 ( .A(u0__abc_49347_n2110), .B(u0__abc_49347_n1179_bF_buf2), .Y(u0__abc_49347_n2111) );
  AND2X2 AND2X2_5760 ( .A(u5__abc_54027_n272), .B(u5__abc_54027_n273), .Y(u5__abc_54027_n274) );
  AND2X2 AND2X2_5761 ( .A(u5__abc_54027_n270), .B(u5__abc_54027_n274), .Y(u5_pack_le1_d) );
  AND2X2 AND2X2_5762 ( .A(u5__abc_54027_n268_1), .B(u5__abc_54027_n276), .Y(u5__abc_54027_n277) );
  AND2X2 AND2X2_5763 ( .A(u5__abc_54027_n277), .B(u5__abc_54027_n267), .Y(u5__abc_54027_n278) );
  AND2X2 AND2X2_5764 ( .A(u5__abc_54027_n279), .B(u5__abc_54027_n271), .Y(u5__abc_54027_n280) );
  AND2X2 AND2X2_5765 ( .A(u5__abc_54027_n281), .B(u5_state_0_), .Y(u5__abc_54027_n282) );
  AND2X2 AND2X2_5766 ( .A(u5__abc_54027_n280), .B(u5__abc_54027_n282), .Y(u5__abc_54027_n283) );
  AND2X2 AND2X2_5767 ( .A(u5__abc_54027_n278), .B(u5__abc_54027_n283), .Y(err) );
  AND2X2 AND2X2_5768 ( .A(u5_state_2_), .B(u5_state_3_), .Y(u5__abc_54027_n285_1) );
  AND2X2 AND2X2_5769 ( .A(u5__abc_54027_n286), .B(u5__abc_54027_n281), .Y(u5__abc_54027_n287) );
  AND2X2 AND2X2_577 ( .A(spec_req_cs_2_bF_buf5), .B(u0_csc2_6_), .Y(u0__abc_49347_n2112) );
  AND2X2 AND2X2_5770 ( .A(u5__abc_54027_n287), .B(u5__abc_54027_n285_1), .Y(u5__abc_54027_n288_1) );
  AND2X2 AND2X2_5771 ( .A(u5__abc_54027_n267), .B(u5_state_5_), .Y(u5__abc_54027_n289) );
  AND2X2 AND2X2_5772 ( .A(u5__abc_54027_n289), .B(u5__abc_54027_n276), .Y(u5__abc_54027_n290_1) );
  AND2X2 AND2X2_5773 ( .A(u5__abc_54027_n288_1), .B(u5__abc_54027_n290_1), .Y(u5__abc_54027_n291) );
  AND2X2 AND2X2_5774 ( .A(u5__abc_54027_n279), .B(u5_state_3_), .Y(u5__abc_54027_n292) );
  AND2X2 AND2X2_5775 ( .A(u5__abc_54027_n282), .B(u5__abc_54027_n292), .Y(u5__abc_54027_n293) );
  AND2X2 AND2X2_5776 ( .A(u5__abc_54027_n293), .B(u5__abc_54027_n290_1), .Y(u5__abc_54027_n294) );
  AND2X2 AND2X2_5777 ( .A(u5__abc_54027_n292), .B(u5__abc_54027_n273), .Y(u5__abc_54027_n296) );
  AND2X2 AND2X2_5778 ( .A(u5__abc_54027_n290_1), .B(u5__abc_54027_n296), .Y(u5__abc_54027_n297) );
  AND2X2 AND2X2_5779 ( .A(u5__abc_54027_n286), .B(u5_state_1_), .Y(u5__abc_54027_n299_1) );
  AND2X2 AND2X2_578 ( .A(u0__abc_49347_n2113), .B(u0__abc_49347_n1178_1_bF_buf2), .Y(u0__abc_49347_n2114) );
  AND2X2 AND2X2_5780 ( .A(u5__abc_54027_n292), .B(u5__abc_54027_n299_1), .Y(u5__abc_54027_n300_1) );
  AND2X2 AND2X2_5781 ( .A(u5__abc_54027_n300_1), .B(u5__abc_54027_n290_1), .Y(u5__abc_54027_n301_1) );
  AND2X2 AND2X2_5782 ( .A(u5__abc_54027_n287), .B(u5__abc_54027_n292), .Y(u5__abc_54027_n303) );
  AND2X2 AND2X2_5783 ( .A(u5__abc_54027_n303), .B(u5__abc_54027_n290_1), .Y(u5__abc_54027_n304) );
  AND2X2 AND2X2_5784 ( .A(u5__abc_54027_n302), .B(u5__abc_54027_n305), .Y(u5__abc_54027_n306) );
  AND2X2 AND2X2_5785 ( .A(u5__abc_54027_n306), .B(u5__abc_54027_n298_1), .Y(u5__abc_54027_n307) );
  AND2X2 AND2X2_5786 ( .A(u5__abc_54027_n307), .B(u5__abc_54027_n295), .Y(u5__abc_54027_n308) );
  AND2X2 AND2X2_5787 ( .A(u5_state_5_), .B(u5_state_4_), .Y(u5__abc_54027_n311_1) );
  AND2X2 AND2X2_5788 ( .A(u5__abc_54027_n311_1), .B(u5__abc_54027_n267), .Y(u5__abc_54027_n312_1) );
  AND2X2 AND2X2_5789 ( .A(u5__abc_54027_n274), .B(u5__abc_54027_n312_1), .Y(u5__abc_54027_n313_1) );
  AND2X2 AND2X2_579 ( .A(spec_req_cs_1_bF_buf5), .B(u0_csc1_6_), .Y(u0__abc_49347_n2115) );
  AND2X2 AND2X2_5790 ( .A(u5__abc_54027_n314), .B(u5_wb_cycle), .Y(u5__abc_54027_n315) );
  AND2X2 AND2X2_5791 ( .A(u5_cke_o_del), .B(u5_burst_act_rd), .Y(u5__abc_54027_n316_1) );
  AND2X2 AND2X2_5792 ( .A(u5__abc_54027_n315), .B(u5__abc_54027_n316_1), .Y(u5__abc_54027_n317) );
  AND2X2 AND2X2_5793 ( .A(u5__abc_54027_n313_1), .B(u5__abc_54027_n317), .Y(u5__abc_54027_n318) );
  AND2X2 AND2X2_5794 ( .A(u5__abc_54027_n278), .B(u5__abc_54027_n288_1), .Y(u5__abc_54027_n319) );
  AND2X2 AND2X2_5795 ( .A(u5__abc_54027_n320), .B(u5_mc_adv_r), .Y(u5__abc_54027_n321_1) );
  AND2X2 AND2X2_5796 ( .A(u5__abc_54027_n319), .B(u5__abc_54027_n321_1), .Y(u5__abc_54027_n322_1) );
  AND2X2 AND2X2_5797 ( .A(u5__abc_54027_n327), .B(u5__abc_54027_n328_1), .Y(u5__abc_54027_n329) );
  AND2X2 AND2X2_5798 ( .A(u5__abc_54027_n326), .B(u5__abc_54027_n329), .Y(u5__abc_54027_n330_1) );
  AND2X2 AND2X2_5799 ( .A(u5__abc_54027_n334), .B(u5__abc_54027_n330_1), .Y(u5_timer_is_zero) );
  AND2X2 AND2X2_58 ( .A(u0_init_req0), .B(init_req), .Y(u0__abc_49347_n1102) );
  AND2X2 AND2X2_580 ( .A(u0__abc_49347_n1952_1_bF_buf1), .B(u0__abc_49347_n2118), .Y(u0__abc_49347_n2119) );
  AND2X2 AND2X2_5800 ( .A(u5__abc_54027_n336), .B(u5__abc_54027_n337), .Y(u5__abc_54027_n338) );
  AND2X2 AND2X2_5801 ( .A(u5__abc_54027_n339), .B(u5__abc_54027_n340), .Y(u5__abc_54027_n341) );
  AND2X2 AND2X2_5802 ( .A(u5__abc_54027_n338), .B(u5__abc_54027_n341), .Y(u5_ir_cnt_done_FF_INPUT) );
  AND2X2 AND2X2_5803 ( .A(u5__abc_54027_n282), .B(u5__abc_54027_n285_1), .Y(u5__abc_54027_n343) );
  AND2X2 AND2X2_5804 ( .A(u5__abc_54027_n343), .B(u5__abc_54027_n312_1), .Y(u5__abc_54027_n344_1) );
  AND2X2 AND2X2_5805 ( .A(u5__abc_54027_n344_1), .B(rfr_ack), .Y(u5__abc_54027_n345) );
  AND2X2 AND2X2_5806 ( .A(u5__abc_54027_n299_1), .B(u5__abc_54027_n285_1), .Y(u5__abc_54027_n346) );
  AND2X2 AND2X2_5807 ( .A(u5__abc_54027_n346), .B(u5__abc_54027_n312_1), .Y(u5__abc_54027_n347) );
  AND2X2 AND2X2_5808 ( .A(u5__abc_54027_n347), .B(rfr_ack), .Y(u5__abc_54027_n348) );
  AND2X2 AND2X2_5809 ( .A(u5__abc_54027_n277), .B(u5_state_6_), .Y(u5__abc_54027_n350) );
  AND2X2 AND2X2_581 ( .A(u0__abc_49347_n2117), .B(u0__abc_49347_n2119), .Y(u0__abc_49347_n2120) );
  AND2X2 AND2X2_5810 ( .A(u5__abc_54027_n283), .B(u5__abc_54027_n350), .Y(u5__abc_54027_n351) );
  AND2X2 AND2X2_5811 ( .A(u5__abc_54027_n351_bF_buf3), .B(rfr_req), .Y(u5__abc_54027_n352) );
  AND2X2 AND2X2_5812 ( .A(u5__abc_54027_n272), .B(u5__abc_54027_n282), .Y(u5__abc_54027_n353) );
  AND2X2 AND2X2_5813 ( .A(u5__abc_54027_n353), .B(u5__abc_54027_n290_1), .Y(u5__abc_54027_n354) );
  AND2X2 AND2X2_5814 ( .A(u5__abc_54027_n283), .B(u5__abc_54027_n312_1), .Y(u5__abc_54027_n355) );
  AND2X2 AND2X2_5815 ( .A(u5__abc_54027_n280), .B(u5__abc_54027_n287), .Y(u5__abc_54027_n359) );
  AND2X2 AND2X2_5816 ( .A(u5__abc_54027_n359), .B(u5__abc_54027_n270), .Y(u5__abc_54027_n360) );
  AND2X2 AND2X2_5817 ( .A(u5__abc_54027_n288_1), .B(u5__abc_54027_n312_1), .Y(u5__abc_54027_n362) );
  AND2X2 AND2X2_5818 ( .A(u5__abc_54027_n361), .B(u5__abc_54027_n363), .Y(u5__abc_54027_n364) );
  AND2X2 AND2X2_5819 ( .A(u5__abc_54027_n270), .B(u5__abc_54027_n346), .Y(u5__abc_54027_n366_1) );
  AND2X2 AND2X2_582 ( .A(u0__abc_49347_n1953_1_bF_buf1), .B(sp_csc_7_), .Y(u0__abc_49347_n2122) );
  AND2X2 AND2X2_5820 ( .A(u5__abc_54027_n365_1), .B(u5__abc_54027_n367_1), .Y(u5__abc_54027_n368) );
  AND2X2 AND2X2_5821 ( .A(u5__abc_54027_n278), .B(u5__abc_54027_n346), .Y(u5__abc_54027_n369) );
  AND2X2 AND2X2_5822 ( .A(u5__abc_54027_n278), .B(u5__abc_54027_n353), .Y(u5__abc_54027_n371) );
  AND2X2 AND2X2_5823 ( .A(u5__abc_54027_n372), .B(u5__abc_54027_n370), .Y(u5__abc_54027_n373) );
  AND2X2 AND2X2_5824 ( .A(u5__abc_54027_n272), .B(u5__abc_54027_n299_1), .Y(u5__abc_54027_n374) );
  AND2X2 AND2X2_5825 ( .A(u5__abc_54027_n278), .B(u5__abc_54027_n374), .Y(u5__abc_54027_n375) );
  AND2X2 AND2X2_5826 ( .A(u5__abc_54027_n270), .B(u5__abc_54027_n343), .Y(u5__abc_54027_n377) );
  AND2X2 AND2X2_5827 ( .A(u5__abc_54027_n376), .B(u5__abc_54027_n378), .Y(u5__abc_54027_n379) );
  AND2X2 AND2X2_5828 ( .A(u5__abc_54027_n373), .B(u5__abc_54027_n379), .Y(u5__abc_54027_n380) );
  AND2X2 AND2X2_5829 ( .A(u5__abc_54027_n380), .B(u5__abc_54027_n368), .Y(u5__abc_54027_n381) );
  AND2X2 AND2X2_583 ( .A(spec_req_cs_5_bF_buf4), .B(u0_csc5_7_), .Y(u0__abc_49347_n2123) );
  AND2X2 AND2X2_5830 ( .A(u5__abc_54027_n374), .B(u5__abc_54027_n270), .Y(u5__abc_54027_n382) );
  AND2X2 AND2X2_5831 ( .A(u5__abc_54027_n303), .B(u5__abc_54027_n270), .Y(u5__abc_54027_n384) );
  AND2X2 AND2X2_5832 ( .A(u5__abc_54027_n383), .B(u5__abc_54027_n385), .Y(u5__abc_54027_n386_1) );
  AND2X2 AND2X2_5833 ( .A(u5__abc_54027_n353), .B(u5__abc_54027_n270), .Y(u5__abc_54027_n387_1) );
  AND2X2 AND2X2_5834 ( .A(u5__abc_54027_n287), .B(u5__abc_54027_n272), .Y(u5__abc_54027_n389_1) );
  AND2X2 AND2X2_5835 ( .A(u5__abc_54027_n389_1), .B(u5__abc_54027_n270), .Y(u5__abc_54027_n390_1) );
  AND2X2 AND2X2_5836 ( .A(u5__abc_54027_n388_1), .B(u5__abc_54027_n391), .Y(u5__abc_54027_n392) );
  AND2X2 AND2X2_5837 ( .A(u5__abc_54027_n386_1), .B(u5__abc_54027_n392), .Y(u5__abc_54027_n393) );
  AND2X2 AND2X2_5838 ( .A(u5__abc_54027_n293), .B(u5__abc_54027_n270), .Y(u5__abc_54027_n397) );
  AND2X2 AND2X2_5839 ( .A(u5__abc_54027_n400), .B(u5__abc_54027_n398), .Y(u5__abc_54027_n401) );
  AND2X2 AND2X2_584 ( .A(u0__abc_49347_n2125), .B(u0__abc_49347_n1185_bF_buf1), .Y(u0__abc_49347_n2126) );
  AND2X2 AND2X2_5840 ( .A(u5__abc_54027_n401), .B(u5__abc_54027_n396), .Y(u5__abc_54027_n402) );
  AND2X2 AND2X2_5841 ( .A(u5__abc_54027_n402), .B(u5__abc_54027_n393), .Y(u5__abc_54027_n403) );
  AND2X2 AND2X2_5842 ( .A(u5__abc_54027_n403), .B(u5__abc_54027_n381), .Y(u5__abc_54027_n404) );
  AND2X2 AND2X2_5843 ( .A(u5__abc_54027_n283), .B(u5__abc_54027_n270), .Y(u5__abc_54027_n405) );
  AND2X2 AND2X2_5844 ( .A(u5__abc_54027_n404), .B(u5__abc_54027_n406), .Y(u5__abc_54027_n407) );
  AND2X2 AND2X2_5845 ( .A(u5__abc_54027_n407), .B(u5__abc_54027_n364), .Y(u5__abc_54027_n408) );
  AND2X2 AND2X2_5846 ( .A(u5__abc_54027_n280), .B(u5__abc_54027_n299_1), .Y(u5__abc_54027_n415) );
  AND2X2 AND2X2_5847 ( .A(u5__abc_54027_n278), .B(u5__abc_54027_n415), .Y(u5__abc_54027_n416) );
  AND2X2 AND2X2_5848 ( .A(u5__abc_54027_n417), .B(u5__abc_54027_n414), .Y(u5__abc_54027_n418) );
  AND2X2 AND2X2_5849 ( .A(u5__abc_54027_n408), .B(u5__abc_54027_n418), .Y(u5__abc_54027_n419) );
  AND2X2 AND2X2_585 ( .A(u0__abc_49347_n2126), .B(u0__abc_49347_n2124), .Y(u0__abc_49347_n2127) );
  AND2X2 AND2X2_5850 ( .A(u5__abc_54027_n389_1), .B(u5__abc_54027_n312_1), .Y(u5__abc_54027_n420) );
  AND2X2 AND2X2_5851 ( .A(u5__abc_54027_n353), .B(u5__abc_54027_n312_1), .Y(u5__abc_54027_n422) );
  AND2X2 AND2X2_5852 ( .A(u5__abc_54027_n423), .B(u5__abc_54027_n421), .Y(u5__abc_54027_n424) );
  AND2X2 AND2X2_5853 ( .A(u5__abc_54027_n293), .B(u5__abc_54027_n312_1), .Y(u5__abc_54027_n425) );
  AND2X2 AND2X2_5854 ( .A(u5__abc_54027_n280), .B(u5__abc_54027_n273), .Y(u5__abc_54027_n427) );
  AND2X2 AND2X2_5855 ( .A(u5__abc_54027_n427), .B(u5__abc_54027_n312_1), .Y(u5__abc_54027_n428) );
  AND2X2 AND2X2_5856 ( .A(u5__abc_54027_n415), .B(u5__abc_54027_n270), .Y(u5__abc_54027_n430_1) );
  AND2X2 AND2X2_5857 ( .A(u5__abc_54027_n427), .B(u5__abc_54027_n270), .Y(u5__abc_54027_n432_1) );
  AND2X2 AND2X2_5858 ( .A(u5__abc_54027_n431), .B(u5__abc_54027_n433_1), .Y(u5__abc_54027_n434) );
  AND2X2 AND2X2_5859 ( .A(u5__abc_54027_n278), .B(u5__abc_54027_n427), .Y(u5__abc_54027_n435) );
  AND2X2 AND2X2_586 ( .A(u0__abc_49347_n2128), .B(u0__abc_49347_n1181_bF_buf1), .Y(u0__abc_49347_n2129) );
  AND2X2 AND2X2_5860 ( .A(u5__abc_54027_n278), .B(u5__abc_54027_n303), .Y(u5__abc_54027_n437_1) );
  AND2X2 AND2X2_5861 ( .A(u5__abc_54027_n438_1), .B(u5__abc_54027_n436), .Y(u5__abc_54027_n439) );
  AND2X2 AND2X2_5862 ( .A(u5__abc_54027_n439), .B(u5__abc_54027_n434), .Y(u5__abc_54027_n440) );
  AND2X2 AND2X2_5863 ( .A(u5__abc_54027_n440), .B(u5__abc_54027_n429_1), .Y(u5__abc_54027_n441) );
  AND2X2 AND2X2_5864 ( .A(u5__abc_54027_n441), .B(u5__abc_54027_n426), .Y(u5__abc_54027_n442) );
  AND2X2 AND2X2_5865 ( .A(u5__abc_54027_n442), .B(u5__abc_54027_n424), .Y(u5__abc_54027_n443) );
  AND2X2 AND2X2_5866 ( .A(u5__abc_54027_n359), .B(u5__abc_54027_n312_1), .Y(u5__abc_54027_n445) );
  AND2X2 AND2X2_5867 ( .A(u5__abc_54027_n274), .B(u5__abc_54027_n290_1), .Y(u5__abc_54027_n447_1) );
  AND2X2 AND2X2_5868 ( .A(u5__abc_54027_n446_1), .B(u5__abc_54027_n448), .Y(u5__abc_54027_n449_1) );
  AND2X2 AND2X2_5869 ( .A(u5__abc_54027_n449_1), .B(u5__abc_54027_n444), .Y(u5__abc_54027_n450) );
  AND2X2 AND2X2_587 ( .A(spec_req_cs_4_bF_buf4), .B(u0_csc4_7_), .Y(u0__abc_49347_n2130) );
  AND2X2 AND2X2_5870 ( .A(u5__abc_54027_n415), .B(u5__abc_54027_n312_1), .Y(u5__abc_54027_n452_1) );
  AND2X2 AND2X2_5871 ( .A(u5__abc_54027_n453), .B(u5__abc_54027_n451_1), .Y(u5__abc_54027_n454) );
  AND2X2 AND2X2_5872 ( .A(u5__abc_54027_n450), .B(u5__abc_54027_n454), .Y(u5__abc_54027_n455) );
  AND2X2 AND2X2_5873 ( .A(u5__abc_54027_n456), .B(u5__abc_54027_n457), .Y(u5__abc_54027_n458) );
  AND2X2 AND2X2_5874 ( .A(u5__abc_54027_n458), .B(u5__abc_54027_n302), .Y(u5__abc_54027_n459) );
  AND2X2 AND2X2_5875 ( .A(u5__abc_54027_n290_1), .B(u5__abc_54027_n346), .Y(u5__abc_54027_n460) );
  AND2X2 AND2X2_5876 ( .A(u5__abc_54027_n459), .B(u5__abc_54027_n462), .Y(u5__abc_54027_n463_1) );
  AND2X2 AND2X2_5877 ( .A(u5__abc_54027_n455), .B(u5__abc_54027_n463_1), .Y(u5__abc_54027_n464) );
  AND2X2 AND2X2_5878 ( .A(u5__abc_54027_n443), .B(u5__abc_54027_n464), .Y(u5__abc_54027_n465) );
  AND2X2 AND2X2_5879 ( .A(u5__abc_54027_n419), .B(u5__abc_54027_n465), .Y(u5__abc_54027_n466) );
  AND2X2 AND2X2_588 ( .A(u0__abc_49347_n2131), .B(u0__abc_49347_n1180_1_bF_buf1), .Y(u0__abc_49347_n2132) );
  AND2X2 AND2X2_5880 ( .A(u5__abc_54027_n469), .B(u5__abc_54027_n470_1), .Y(u5__abc_54027_n471) );
  AND2X2 AND2X2_5881 ( .A(u5__abc_54027_n471), .B(u5__abc_54027_n468_1), .Y(u5__abc_54027_n472) );
  AND2X2 AND2X2_5882 ( .A(u5_burst_act_rd_FF_INPUT), .B(u5__abc_54027_n474), .Y(u5__abc_54027_n475_1) );
  AND2X2 AND2X2_5883 ( .A(u5__abc_54027_n475_1), .B(u5__abc_54027_n467), .Y(u5__abc_54027_n476) );
  AND2X2 AND2X2_5884 ( .A(u5__abc_54027_n314), .B(u5__abc_54027_n477), .Y(u5__abc_54027_n478_1) );
  AND2X2 AND2X2_5885 ( .A(u5_cnt), .B(u5_cke_r), .Y(u5__abc_54027_n479) );
  AND2X2 AND2X2_5886 ( .A(u5__abc_54027_n482), .B(u5__abc_54027_n481), .Y(u5__abc_54027_n483) );
  AND2X2 AND2X2_5887 ( .A(u5__abc_54027_n476), .B(u5__abc_54027_n483), .Y(u5__abc_54027_n484_1) );
  AND2X2 AND2X2_5888 ( .A(u5__abc_54027_n473), .B(u5_wb_cycle), .Y(u5__abc_54027_n485) );
  AND2X2 AND2X2_5889 ( .A(u5__abc_54027_n488), .B(csc_s_2_bF_buf2), .Y(u5__abc_54027_n489) );
  AND2X2 AND2X2_589 ( .A(spec_req_cs_3_bF_buf4), .B(u0_csc3_7_), .Y(u0__abc_49347_n2133) );
  AND2X2 AND2X2_5890 ( .A(u5__abc_54027_n489), .B(csc_s_1_), .Y(u5__abc_54027_n490) );
  AND2X2 AND2X2_5891 ( .A(u5__abc_54027_n477), .B(u1_wb_write_go), .Y(u5__abc_54027_n491) );
  AND2X2 AND2X2_5892 ( .A(u5__abc_54027_n490), .B(u5__abc_54027_n491), .Y(u5__abc_54027_n492) );
  AND2X2 AND2X2_5893 ( .A(u5__abc_54027_n500), .B(u5__abc_54027_n501), .Y(u5_no_wb_cycle_FF_INPUT) );
  AND2X2 AND2X2_5894 ( .A(u5__abc_54027_n503), .B(u5_lookup_ready2), .Y(u5__abc_54027_n504_1) );
  AND2X2 AND2X2_5895 ( .A(u5__abc_54027_n499), .B(u5__abc_54027_n504_1), .Y(u5__abc_54027_n505_1) );
  AND2X2 AND2X2_5896 ( .A(u5__abc_54027_n506), .B(u5_susp_req_r), .Y(u5__abc_54027_n507) );
  AND2X2 AND2X2_5897 ( .A(u5_lookup_ready2), .B(lmr_req), .Y(u5__abc_54027_n509) );
  AND2X2 AND2X2_5898 ( .A(u5__abc_54027_n511), .B(u5__abc_54027_n512_1), .Y(u5__abc_54027_n513_1) );
  AND2X2 AND2X2_5899 ( .A(u5__abc_54027_n510), .B(u5__abc_54027_n513_1), .Y(u5__abc_54027_n514) );
  AND2X2 AND2X2_59 ( .A(u0__abc_49347_n1104), .B(u0_sreq_cs_le), .Y(u0__abc_49347_n1105_1) );
  AND2X2 AND2X2_590 ( .A(u0__abc_49347_n2134), .B(u0__abc_49347_n1179_bF_buf1), .Y(u0__abc_49347_n2135) );
  AND2X2 AND2X2_5900 ( .A(u5__abc_54027_n514), .B(u5__abc_54027_n508), .Y(u5__abc_54027_n515) );
  AND2X2 AND2X2_5901 ( .A(u5__abc_54027_n505_1), .B(u5__abc_54027_n515), .Y(u5__abc_54027_n516) );
  AND2X2 AND2X2_5902 ( .A(u5__abc_54027_n516), .B(u5__abc_54027_n492), .Y(u5__abc_54027_n517) );
  AND2X2 AND2X2_5903 ( .A(u5__abc_54027_n519), .B(u5_tmr_done), .Y(u5__abc_54027_n520) );
  AND2X2 AND2X2_5904 ( .A(u5__abc_54027_n416), .B(u5_tmr_done), .Y(u5__abc_54027_n522) );
  AND2X2 AND2X2_5905 ( .A(u5__abc_54027_n523_1), .B(u5__abc_54027_n426), .Y(u5__abc_54027_n524_1) );
  AND2X2 AND2X2_5906 ( .A(u5__abc_54027_n524_1), .B(u5__abc_54027_n521), .Y(u5__abc_54027_n525) );
  AND2X2 AND2X2_5907 ( .A(u5__abc_54027_n525), .B(u5__abc_54027_n459), .Y(u5__abc_54027_n526) );
  AND2X2 AND2X2_5908 ( .A(u5__abc_54027_n526), .B(u5__abc_54027_n518), .Y(u5__abc_54027_n527) );
  AND2X2 AND2X2_5909 ( .A(u5__abc_54027_n408), .B(u5__abc_54027_n527), .Y(u5__abc_54027_n528) );
  AND2X2 AND2X2_591 ( .A(spec_req_cs_2_bF_buf4), .B(u0_csc2_7_), .Y(u0__abc_49347_n2136) );
  AND2X2 AND2X2_5910 ( .A(u5__abc_54027_n487), .B(u5__abc_54027_n528), .Y(u5__abc_54027_n529) );
  AND2X2 AND2X2_5911 ( .A(u5_cmd_del_0_), .B(u1_wr_cycle), .Y(u5__abc_54027_n532_1) );
  AND2X2 AND2X2_5912 ( .A(u5_cmd_0_), .B(u5__abc_54027_n533), .Y(u5__abc_54027_n534) );
  AND2X2 AND2X2_5913 ( .A(u5__abc_54027_n441), .B(u5__abc_54027_n486_1), .Y(u5__abc_54027_n536) );
  AND2X2 AND2X2_5914 ( .A(u5__abc_54027_n536), .B(u5__abc_54027_n455), .Y(u5__abc_54027_n537) );
  AND2X2 AND2X2_5915 ( .A(u5__abc_54027_n419), .B(u5__abc_54027_n537), .Y(u5__abc_54027_n538) );
  AND2X2 AND2X2_5916 ( .A(u1_wr_cycle), .B(u5_cmd_del_1_), .Y(u5__abc_54027_n541) );
  AND2X2 AND2X2_5917 ( .A(u5_cmd_1_), .B(u5__abc_54027_n533), .Y(u5__abc_54027_n542) );
  AND2X2 AND2X2_5918 ( .A(u5__abc_54027_n418), .B(u5__abc_54027_n361), .Y(u5__abc_54027_n544_1) );
  AND2X2 AND2X2_5919 ( .A(u5__abc_54027_n521), .B(u5__abc_54027_n546), .Y(u5__abc_54027_n547) );
  AND2X2 AND2X2_592 ( .A(u0__abc_49347_n2137), .B(u0__abc_49347_n1178_1_bF_buf1), .Y(u0__abc_49347_n2138) );
  AND2X2 AND2X2_5920 ( .A(u5__abc_54027_n547), .B(u5__abc_54027_n544_1), .Y(u5__abc_54027_n548) );
  AND2X2 AND2X2_5921 ( .A(u5__abc_54027_n443), .B(u5__abc_54027_n548), .Y(u5__abc_54027_n549) );
  AND2X2 AND2X2_5922 ( .A(u5__abc_54027_n549), .B(u5__abc_54027_n407), .Y(u5__abc_54027_n550) );
  AND2X2 AND2X2_5923 ( .A(u1_wr_cycle), .B(u5_cmd_del_2_), .Y(u5__abc_54027_n553_1) );
  AND2X2 AND2X2_5924 ( .A(u5_cmd_2_), .B(u5__abc_54027_n533), .Y(u5__abc_54027_n554) );
  AND2X2 AND2X2_5925 ( .A(u5__abc_54027_n556), .B(u5__abc_54027_n557), .Y(u5__abc_54027_n558) );
  AND2X2 AND2X2_5926 ( .A(u5__abc_54027_n561), .B(mc_c_oe_d), .Y(u5__abc_54027_n562) );
  AND2X2 AND2X2_5927 ( .A(u5__abc_54027_n562), .B(u5__abc_54027_n560), .Y(u5__abc_54027_n563_1) );
  AND2X2 AND2X2_5928 ( .A(u5__abc_54027_n569_1), .B(u5__abc_54027_n405), .Y(u5__abc_54027_n570) );
  AND2X2 AND2X2_5929 ( .A(u5__abc_54027_n452_1), .B(u5_tmr_done), .Y(u5__abc_54027_n572_1) );
  AND2X2 AND2X2_593 ( .A(spec_req_cs_1_bF_buf4), .B(u0_csc1_7_), .Y(u0__abc_49347_n2139) );
  AND2X2 AND2X2_5930 ( .A(u5__abc_54027_n572_1), .B(u5__abc_54027_n519), .Y(u5__abc_54027_n573) );
  AND2X2 AND2X2_5931 ( .A(u5__abc_54027_n462), .B(u5__abc_54027_n423), .Y(u5__abc_54027_n575) );
  AND2X2 AND2X2_5932 ( .A(u5__abc_54027_n575), .B(u5__abc_54027_n459), .Y(u5__abc_54027_n576) );
  AND2X2 AND2X2_5933 ( .A(u5__abc_54027_n576), .B(u5__abc_54027_n574), .Y(u5__abc_54027_n577_1) );
  AND2X2 AND2X2_5934 ( .A(u5__abc_54027_n450), .B(u5__abc_54027_n451_1), .Y(u5__abc_54027_n578) );
  AND2X2 AND2X2_5935 ( .A(u5__abc_54027_n579_1), .B(u5__abc_54027_n580), .Y(u5__abc_54027_n581) );
  AND2X2 AND2X2_5936 ( .A(u5__abc_54027_n362), .B(u5__abc_54027_n545_1), .Y(u5__abc_54027_n582) );
  AND2X2 AND2X2_5937 ( .A(u5__abc_54027_n581), .B(u5__abc_54027_n583), .Y(u5__abc_54027_n584) );
  AND2X2 AND2X2_5938 ( .A(u5__abc_54027_n584), .B(u5__abc_54027_n578), .Y(u5__abc_54027_n585) );
  AND2X2 AND2X2_5939 ( .A(u5__abc_54027_n577_1), .B(u5__abc_54027_n585), .Y(u5__abc_54027_n586) );
  AND2X2 AND2X2_594 ( .A(u0__abc_49347_n1952_1_bF_buf0), .B(u0__abc_49347_n2142), .Y(u0__abc_49347_n2143) );
  AND2X2 AND2X2_5940 ( .A(u5__abc_54027_n351_bF_buf2), .B(u5__abc_54027_n515), .Y(u5__abc_54027_n587) );
  AND2X2 AND2X2_5941 ( .A(u5__abc_54027_n587), .B(u5__abc_54027_n505_1), .Y(u5__abc_54027_n588) );
  AND2X2 AND2X2_5942 ( .A(u5__abc_54027_n490), .B(u5__abc_54027_n477), .Y(u5__abc_54027_n589) );
  AND2X2 AND2X2_5943 ( .A(u5__abc_54027_n489), .B(u5__abc_54027_n590), .Y(u5__abc_54027_n591) );
  AND2X2 AND2X2_5944 ( .A(u5__abc_54027_n594), .B(u5__abc_54027_n590), .Y(u5__abc_54027_n595) );
  AND2X2 AND2X2_5945 ( .A(u5__abc_54027_n596), .B(u5__abc_54027_n592_1), .Y(u5__abc_54027_n597) );
  AND2X2 AND2X2_5946 ( .A(u5__abc_54027_n477), .B(u5__abc_54027_n501), .Y(u5__abc_54027_n598) );
  AND2X2 AND2X2_5947 ( .A(u5__abc_54027_n597), .B(u5__abc_54027_n598), .Y(u5__abc_54027_n599) );
  AND2X2 AND2X2_5948 ( .A(u5__abc_54027_n600), .B(u5__abc_54027_n588), .Y(u5__abc_54027_n601_1) );
  AND2X2 AND2X2_5949 ( .A(u5__abc_54027_n404), .B(u5__abc_54027_n442), .Y(u5__abc_54027_n603) );
  AND2X2 AND2X2_595 ( .A(u0__abc_49347_n2141), .B(u0__abc_49347_n2143), .Y(u0__abc_49347_n2144_1) );
  AND2X2 AND2X2_5950 ( .A(u5__abc_54027_n603), .B(u5__abc_54027_n602), .Y(u5__abc_54027_n604) );
  AND2X2 AND2X2_5951 ( .A(u5__abc_54027_n604), .B(u5__abc_54027_n586), .Y(u5__abc_54027_n605_1) );
  AND2X2 AND2X2_5952 ( .A(u5__abc_54027_n571), .B(u5__abc_54027_n605_1), .Y(u5__abc_54027_n606) );
  AND2X2 AND2X2_5953 ( .A(u5__abc_54027_n559), .B(u5__abc_54027_n606), .Y(u5__abc_54027_n607) );
  AND2X2 AND2X2_5954 ( .A(u1_wr_cycle), .B(u5_cmd_del_3_), .Y(u5__abc_54027_n609) );
  AND2X2 AND2X2_5955 ( .A(u5_cmd_3_), .B(u5__abc_54027_n533), .Y(u5__abc_54027_n610) );
  AND2X2 AND2X2_5956 ( .A(u5__abc_54027_n588), .B(u5__abc_54027_n491), .Y(u5__abc_54027_n612) );
  AND2X2 AND2X2_5957 ( .A(u5__abc_54027_n612), .B(u5__abc_54027_n596), .Y(u5__abc_54027_n613) );
  AND2X2 AND2X2_5958 ( .A(u5__abc_54027_n300_1), .B(u5__abc_54027_n312_1), .Y(u5__abc_54027_n615) );
  AND2X2 AND2X2_5959 ( .A(u5__abc_54027_n615), .B(u5__abc_54027_n491), .Y(u5__abc_54027_n616) );
  AND2X2 AND2X2_596 ( .A(u0__abc_49347_n1953_1_bF_buf0), .B(sp_csc_9_), .Y(u0__abc_49347_n2170) );
  AND2X2 AND2X2_5960 ( .A(u5__abc_54027_n278), .B(u5__abc_54027_n274), .Y(u5__abc_54027_n619) );
  AND2X2 AND2X2_5961 ( .A(u5__abc_54027_n619), .B(u5__abc_54027_n491), .Y(u5__abc_54027_n620_1) );
  AND2X2 AND2X2_5962 ( .A(u1_wr_cycle), .B(u5_data_oe_r2), .Y(u5__abc_54027_n626) );
  AND2X2 AND2X2_5963 ( .A(u5_data_oe_d), .B(u5__abc_54027_n533), .Y(u5__abc_54027_n627) );
  AND2X2 AND2X2_5964 ( .A(u5__abc_54027_n477), .B(u5__abc_54027_n629), .Y(u5__abc_54027_n630_1) );
  AND2X2 AND2X2_5965 ( .A(wb_we_i), .B(wb_stb_i_bF_buf0), .Y(u5__abc_54027_n632_1) );
  AND2X2 AND2X2_5966 ( .A(u5__abc_54027_n636), .B(u5__abc_54027_n637), .Y(u5__abc_54027_n638_1) );
  AND2X2 AND2X2_5967 ( .A(u5__abc_54027_n638_1), .B(u5__abc_54027_n635), .Y(u5__abc_54027_n639) );
  AND2X2 AND2X2_5968 ( .A(u5__abc_54027_n437_1), .B(u5_cmd_asserted_bF_buf3), .Y(u5__abc_54027_n644) );
  AND2X2 AND2X2_5969 ( .A(u5__abc_54027_n644), .B(u5__abc_54027_n491), .Y(u5__abc_54027_n645) );
  AND2X2 AND2X2_597 ( .A(spec_req_cs_5_bF_buf3), .B(u0_csc5_9_), .Y(u0__abc_49347_n2171) );
  AND2X2 AND2X2_5970 ( .A(u5__abc_54027_n296), .B(u5__abc_54027_n312_1), .Y(u5__abc_54027_n646) );
  AND2X2 AND2X2_5971 ( .A(u1_wb_write_go), .B(u5_tmr_done), .Y(u5__abc_54027_n647) );
  AND2X2 AND2X2_5972 ( .A(u5__abc_54027_n646), .B(u5__abc_54027_n647), .Y(u5__abc_54027_n648) );
  AND2X2 AND2X2_5973 ( .A(u5__abc_54027_n650), .B(u5__abc_54027_n629), .Y(u5__abc_54027_n651) );
  AND2X2 AND2X2_5974 ( .A(u5__abc_54027_n300_1), .B(u5__abc_54027_n270), .Y(u5__abc_54027_n654_1) );
  AND2X2 AND2X2_5975 ( .A(u5__abc_54027_n273), .B(u5__abc_54027_n285_1), .Y(u5__abc_54027_n656) );
  AND2X2 AND2X2_5976 ( .A(u5__abc_54027_n278), .B(u5__abc_54027_n656), .Y(u5__abc_54027_n657_1) );
  AND2X2 AND2X2_5977 ( .A(u5__abc_54027_n655), .B(u5__abc_54027_n658), .Y(u5__abc_54027_n659) );
  AND2X2 AND2X2_5978 ( .A(u5__abc_54027_n659), .B(u5__abc_54027_n653), .Y(u5__abc_54027_n660) );
  AND2X2 AND2X2_5979 ( .A(u5__abc_54027_n371), .B(u5_tmr_done), .Y(u5__abc_54027_n661) );
  AND2X2 AND2X2_598 ( .A(u0__abc_49347_n2173), .B(u0__abc_49347_n1185_bF_buf0), .Y(u0__abc_49347_n2174) );
  AND2X2 AND2X2_5980 ( .A(u5__abc_54027_n662), .B(u5__abc_54027_n523_1), .Y(u5__abc_54027_n663) );
  AND2X2 AND2X2_5981 ( .A(u5__abc_54027_n663), .B(u5__abc_54027_n660), .Y(u5__abc_54027_n664) );
  AND2X2 AND2X2_5982 ( .A(u5__abc_54027_n652), .B(u5__abc_54027_n664), .Y(u5__abc_54027_n665) );
  AND2X2 AND2X2_5983 ( .A(u5__abc_54027_n613), .B(u5__abc_54027_n666_1), .Y(u5__abc_54027_n667) );
  AND2X2 AND2X2_5984 ( .A(u5__abc_54027_n665), .B(u5__abc_54027_n668), .Y(u5__abc_54027_n669) );
  AND2X2 AND2X2_5985 ( .A(u5__abc_54027_n670), .B(u5__abc_54027_n671), .Y(u5__abc_54027_n672_1) );
  AND2X2 AND2X2_5986 ( .A(u5__abc_54027_n673), .B(u5__abc_54027_n458), .Y(u5__abc_54027_n674) );
  AND2X2 AND2X2_5987 ( .A(u5__abc_54027_n674), .B(u5__abc_54027_n672_1), .Y(u5__abc_54027_n675) );
  AND2X2 AND2X2_5988 ( .A(u5__abc_54027_n675), .B(u5__abc_54027_n563_1), .Y(u5__abc_54027_n676) );
  AND2X2 AND2X2_5989 ( .A(u5__abc_54027_n676), .B(u5__abc_54027_n472), .Y(u5__abc_54027_n677) );
  AND2X2 AND2X2_599 ( .A(u0__abc_49347_n2174), .B(u0__abc_49347_n2172), .Y(u0__abc_49347_n2175) );
  AND2X2 AND2X2_5990 ( .A(u5__abc_54027_n491), .B(u5__abc_54027_n629), .Y(u5__abc_54027_n679) );
  AND2X2 AND2X2_5991 ( .A(u5__abc_54027_n422), .B(u5_cmd_asserted_bF_buf2), .Y(u5__abc_54027_n680) );
  AND2X2 AND2X2_5992 ( .A(u5__abc_54027_n680), .B(u5_wb_cycle), .Y(u5__abc_54027_n681_1) );
  AND2X2 AND2X2_5993 ( .A(u5__abc_54027_n420), .B(u1_wr_cycle), .Y(u5__abc_54027_n682) );
  AND2X2 AND2X2_5994 ( .A(u5__abc_54027_n683), .B(u5__abc_54027_n679), .Y(u5__abc_54027_n684) );
  AND2X2 AND2X2_5995 ( .A(u5__abc_54027_n686), .B(u5__abc_54027_n669), .Y(u5__abc_54027_n687_1) );
  AND2X2 AND2X2_5996 ( .A(u5__abc_54027_n687_1), .B(u5__abc_54027_n643_1), .Y(u5__abc_54027_n688) );
  AND2X2 AND2X2_5997 ( .A(wb_stb_i_bF_buf5), .B(u5_wb_first), .Y(u5__abc_54027_n691) );
  AND2X2 AND2X2_5998 ( .A(u5__abc_54027_n689), .B(u5__abc_54027_n692), .Y(u5_wb_stb_first_FF_INPUT) );
  AND2X2 AND2X2_5999 ( .A(u5__abc_54027_n414), .B(u5_ap_en), .Y(u5__abc_54027_n694_1) );
  AND2X2 AND2X2_6 ( .A(_abc_55805_n254), .B(_abc_55805_n255), .Y(_abc_55805_n256) );
  AND2X2 AND2X2_60 ( .A(u0__abc_49347_n1106), .B(u0__abc_49347_n1107_1), .Y(u0_spec_req_cs_0__FF_INPUT) );
  AND2X2 AND2X2_600 ( .A(u0__abc_49347_n2176), .B(u0__abc_49347_n1181_bF_buf0), .Y(u0__abc_49347_n2177) );
  AND2X2 AND2X2_6000 ( .A(u5__abc_54027_n351_bF_buf1), .B(u5__abc_54027_n519), .Y(u5__abc_54027_n695) );
  AND2X2 AND2X2_6001 ( .A(u5__abc_54027_n677), .B(u5__abc_54027_n695), .Y(u5__abc_54027_n696) );
  AND2X2 AND2X2_6002 ( .A(dv), .B(u5__abc_54027_n533), .Y(u5__abc_54027_n700) );
  AND2X2 AND2X2_6003 ( .A(u5__abc_54027_n699_1), .B(u5__abc_54027_n701), .Y(u5__abc_54027_n702) );
  AND2X2 AND2X2_6004 ( .A(u5__abc_54027_n703), .B(u5__abc_54027_n698), .Y(u5__abc_54027_n704) );
  AND2X2 AND2X2_6005 ( .A(u5__abc_54027_n702), .B(u5_burst_cnt_0_), .Y(u5__abc_54027_n705_1) );
  AND2X2 AND2X2_6006 ( .A(u5__abc_54027_n676), .B(u5__abc_54027_n469), .Y(u5__abc_54027_n708) );
  AND2X2 AND2X2_6007 ( .A(u5__abc_54027_n709_1), .B(1'b0), .Y(u5__abc_54027_n710) );
  AND2X2 AND2X2_6008 ( .A(u5__abc_54027_n712), .B(u5__abc_54027_n370), .Y(u5__abc_54027_n713_1) );
  AND2X2 AND2X2_6009 ( .A(u5__abc_54027_n707), .B(u5__abc_54027_n713_1), .Y(u5_burst_cnt_0__FF_INPUT) );
  AND2X2 AND2X2_601 ( .A(spec_req_cs_4_bF_buf3), .B(u0_csc4_9_), .Y(u0__abc_49347_n2178) );
  AND2X2 AND2X2_6010 ( .A(u5__abc_54027_n715), .B(u5_burst_cnt_1_), .Y(u5__abc_54027_n716) );
  AND2X2 AND2X2_6011 ( .A(u5__abc_54027_n704), .B(u5__abc_54027_n717), .Y(u5__abc_54027_n718) );
  AND2X2 AND2X2_6012 ( .A(u5__abc_54027_n709_1), .B(1'b0), .Y(u5__abc_54027_n721) );
  AND2X2 AND2X2_6013 ( .A(u5__abc_54027_n470_1), .B(tms_s_0_), .Y(u5__abc_54027_n722) );
  AND2X2 AND2X2_6014 ( .A(u5__abc_54027_n708), .B(u5__abc_54027_n722), .Y(u5__abc_54027_n723) );
  AND2X2 AND2X2_6015 ( .A(u5__abc_54027_n725), .B(u5__abc_54027_n370), .Y(u5__abc_54027_n726) );
  AND2X2 AND2X2_6016 ( .A(u5__abc_54027_n720), .B(u5__abc_54027_n726), .Y(u5_burst_cnt_1__FF_INPUT) );
  AND2X2 AND2X2_6017 ( .A(u5__abc_54027_n718), .B(u5__abc_54027_n728), .Y(u5__abc_54027_n729_1) );
  AND2X2 AND2X2_6018 ( .A(u5__abc_54027_n730), .B(u5_burst_cnt_2_), .Y(u5__abc_54027_n731) );
  AND2X2 AND2X2_6019 ( .A(u5__abc_54027_n732), .B(u5__abc_54027_n414), .Y(u5__abc_54027_n733) );
  AND2X2 AND2X2_602 ( .A(u0__abc_49347_n2179), .B(u0__abc_49347_n1180_1_bF_buf0), .Y(u0__abc_49347_n2180_1) );
  AND2X2 AND2X2_6020 ( .A(u5__abc_54027_n708), .B(tms_s_1_), .Y(u5__abc_54027_n734) );
  AND2X2 AND2X2_6021 ( .A(u5__abc_54027_n734), .B(u5__abc_54027_n468_1), .Y(u5__abc_54027_n735) );
  AND2X2 AND2X2_6022 ( .A(u5__abc_54027_n709_1), .B(1'b0), .Y(u5__abc_54027_n736) );
  AND2X2 AND2X2_6023 ( .A(u5__abc_54027_n737_1), .B(u5__abc_54027_n351_bF_buf2), .Y(u5__abc_54027_n738) );
  AND2X2 AND2X2_6024 ( .A(u5__abc_54027_n741), .B(u5_burst_cnt_3_), .Y(u5__abc_54027_n742) );
  AND2X2 AND2X2_6025 ( .A(u5__abc_54027_n703), .B(u5__abc_54027_n253_1), .Y(u5__abc_54027_n743) );
  AND2X2 AND2X2_6026 ( .A(u5__abc_54027_n734), .B(tms_s_0_), .Y(u5__abc_54027_n746) );
  AND2X2 AND2X2_6027 ( .A(u5__abc_54027_n709_1), .B(1'b0), .Y(u5__abc_54027_n747_1) );
  AND2X2 AND2X2_6028 ( .A(u5__abc_54027_n749), .B(u5__abc_54027_n370), .Y(u5__abc_54027_n750) );
  AND2X2 AND2X2_6029 ( .A(u5__abc_54027_n745), .B(u5__abc_54027_n750), .Y(u5_burst_cnt_3__FF_INPUT) );
  AND2X2 AND2X2_603 ( .A(spec_req_cs_3_bF_buf3), .B(u0_csc3_9_), .Y(u0__abc_49347_n2181) );
  AND2X2 AND2X2_6030 ( .A(u5__abc_54027_n752_1), .B(u5_burst_cnt_4_), .Y(u5__abc_54027_n753) );
  AND2X2 AND2X2_6031 ( .A(u5__abc_54027_n703), .B(u5__abc_54027_n254), .Y(u5__abc_54027_n754) );
  AND2X2 AND2X2_6032 ( .A(u5__abc_54027_n755_1), .B(u5__abc_54027_n414), .Y(u5__abc_54027_n756) );
  AND2X2 AND2X2_6033 ( .A(u5__abc_54027_n351_bF_buf0), .B(1'b0), .Y(u5__abc_54027_n757) );
  AND2X2 AND2X2_6034 ( .A(u5__abc_54027_n709_1), .B(u5__abc_54027_n757), .Y(u5__abc_54027_n758) );
  AND2X2 AND2X2_6035 ( .A(u5__abc_54027_n759_1), .B(u5__abc_54027_n370), .Y(u5_burst_cnt_4__FF_INPUT) );
  AND2X2 AND2X2_6036 ( .A(u5__abc_54027_n761), .B(u5_burst_cnt_5_), .Y(u5__abc_54027_n762_1) );
  AND2X2 AND2X2_6037 ( .A(u5__abc_54027_n703), .B(u5__abc_54027_n255_1), .Y(u5__abc_54027_n763_1) );
  AND2X2 AND2X2_6038 ( .A(u5__abc_54027_n709_1), .B(1'b0), .Y(u5__abc_54027_n766_1) );
  AND2X2 AND2X2_6039 ( .A(u5__abc_54027_n767_1), .B(u5__abc_54027_n370), .Y(u5__abc_54027_n768) );
  AND2X2 AND2X2_604 ( .A(u0__abc_49347_n2182), .B(u0__abc_49347_n1179_bF_buf0), .Y(u0__abc_49347_n2183) );
  AND2X2 AND2X2_6040 ( .A(u5__abc_54027_n765), .B(u5__abc_54027_n768), .Y(u5_burst_cnt_5__FF_INPUT) );
  AND2X2 AND2X2_6041 ( .A(u5__abc_54027_n770), .B(u5_burst_cnt_6_), .Y(u5__abc_54027_n771_1) );
  AND2X2 AND2X2_6042 ( .A(u5__abc_54027_n763_1), .B(u5__abc_54027_n260_1), .Y(u5__abc_54027_n772_1) );
  AND2X2 AND2X2_6043 ( .A(u5__abc_54027_n773), .B(u5__abc_54027_n414), .Y(u5__abc_54027_n774) );
  AND2X2 AND2X2_6044 ( .A(u5__abc_54027_n351_bF_buf2), .B(1'b0), .Y(u5__abc_54027_n775) );
  AND2X2 AND2X2_6045 ( .A(u5__abc_54027_n709_1), .B(u5__abc_54027_n775), .Y(u5__abc_54027_n776) );
  AND2X2 AND2X2_6046 ( .A(u5__abc_54027_n777), .B(u5__abc_54027_n370), .Y(u5_burst_cnt_6__FF_INPUT) );
  AND2X2 AND2X2_6047 ( .A(u5__abc_54027_n779), .B(u5_burst_cnt_7_), .Y(u5__abc_54027_n780) );
  AND2X2 AND2X2_6048 ( .A(u5__abc_54027_n772_1), .B(u5__abc_54027_n261), .Y(u5__abc_54027_n781) );
  AND2X2 AND2X2_6049 ( .A(u5__abc_54027_n709_1), .B(1'b0), .Y(u5__abc_54027_n784) );
  AND2X2 AND2X2_605 ( .A(spec_req_cs_2_bF_buf3), .B(u0_csc2_9_), .Y(u0__abc_49347_n2184) );
  AND2X2 AND2X2_6050 ( .A(u5__abc_54027_n785), .B(u5__abc_54027_n370), .Y(u5__abc_54027_n786) );
  AND2X2 AND2X2_6051 ( .A(u5__abc_54027_n783), .B(u5__abc_54027_n786), .Y(u5_burst_cnt_7__FF_INPUT) );
  AND2X2 AND2X2_6052 ( .A(u5__abc_54027_n781), .B(u5__abc_54027_n258), .Y(u5__abc_54027_n788) );
  AND2X2 AND2X2_6053 ( .A(u5__abc_54027_n255_1), .B(u5__abc_54027_n262), .Y(u5__abc_54027_n789) );
  AND2X2 AND2X2_6054 ( .A(u5__abc_54027_n791_1), .B(u5_burst_cnt_8_), .Y(u5__abc_54027_n792) );
  AND2X2 AND2X2_6055 ( .A(u5__abc_54027_n709_1), .B(page_size_8_), .Y(u5__abc_54027_n795) );
  AND2X2 AND2X2_6056 ( .A(u5__abc_54027_n796), .B(u5__abc_54027_n370), .Y(u5__abc_54027_n797) );
  AND2X2 AND2X2_6057 ( .A(u5__abc_54027_n794), .B(u5__abc_54027_n797), .Y(u5_burst_cnt_8__FF_INPUT) );
  AND2X2 AND2X2_6058 ( .A(u5__abc_54027_n789), .B(u5__abc_54027_n258), .Y(u5__abc_54027_n799) );
  AND2X2 AND2X2_6059 ( .A(u5__abc_54027_n802), .B(u5__abc_54027_n800), .Y(u5__abc_54027_n803) );
  AND2X2 AND2X2_606 ( .A(u0__abc_49347_n2185), .B(u0__abc_49347_n1178_1_bF_buf0), .Y(u0__abc_49347_n2186) );
  AND2X2 AND2X2_6060 ( .A(u5__abc_54027_n805), .B(u5__abc_54027_n804), .Y(u5__abc_54027_n806) );
  AND2X2 AND2X2_6061 ( .A(u5__abc_54027_n806), .B(u5__abc_54027_n414), .Y(u5__abc_54027_n807) );
  AND2X2 AND2X2_6062 ( .A(u5__abc_54027_n351_bF_buf3), .B(page_size_9_), .Y(u5__abc_54027_n808) );
  AND2X2 AND2X2_6063 ( .A(u5__abc_54027_n709_1), .B(u5__abc_54027_n808), .Y(u5__abc_54027_n809) );
  AND2X2 AND2X2_6064 ( .A(u5__abc_54027_n810_1), .B(u5__abc_54027_n370), .Y(u5_burst_cnt_9__FF_INPUT) );
  AND2X2 AND2X2_6065 ( .A(u5__abc_54027_n789), .B(u5__abc_54027_n259_1), .Y(u5__abc_54027_n812) );
  AND2X2 AND2X2_6066 ( .A(u5__abc_54027_n815), .B(u5__abc_54027_n813), .Y(u5__abc_54027_n816) );
  AND2X2 AND2X2_6067 ( .A(u5__abc_54027_n818), .B(u5__abc_54027_n817), .Y(u5__abc_54027_n819) );
  AND2X2 AND2X2_6068 ( .A(u5__abc_54027_n819), .B(u5__abc_54027_n414), .Y(u5__abc_54027_n820) );
  AND2X2 AND2X2_6069 ( .A(u5__abc_54027_n351_bF_buf2), .B(page_size_10_bF_buf3), .Y(u5__abc_54027_n821_1) );
  AND2X2 AND2X2_607 ( .A(spec_req_cs_1_bF_buf3), .B(u0_csc1_9_), .Y(u0__abc_49347_n2187) );
  AND2X2 AND2X2_6070 ( .A(u5__abc_54027_n709_1), .B(u5__abc_54027_n821_1), .Y(u5__abc_54027_n822) );
  AND2X2 AND2X2_6071 ( .A(u5__abc_54027_n823), .B(u5__abc_54027_n370), .Y(u5_burst_cnt_10__FF_INPUT) );
  AND2X2 AND2X2_6072 ( .A(u5__abc_54027_n301_1), .B(u5_cmd_asserted_bF_buf1), .Y(u5__abc_54027_n825) );
  AND2X2 AND2X2_6073 ( .A(u5__abc_54027_n826), .B(u5_ir_cnt_0_), .Y(u5__abc_54027_n827) );
  AND2X2 AND2X2_6074 ( .A(u5__abc_54027_n825), .B(u5__abc_54027_n337), .Y(u5__abc_54027_n828) );
  AND2X2 AND2X2_6075 ( .A(u5__abc_54027_n829), .B(u5__abc_54027_n444), .Y(u5_ir_cnt_0__FF_INPUT) );
  AND2X2 AND2X2_6076 ( .A(u5__abc_54027_n831), .B(u5_ir_cnt_1_), .Y(u5__abc_54027_n832) );
  AND2X2 AND2X2_6077 ( .A(u5__abc_54027_n828), .B(u5__abc_54027_n336), .Y(u5__abc_54027_n833_1) );
  AND2X2 AND2X2_6078 ( .A(u5__abc_54027_n836), .B(u5_ir_cnt_2_), .Y(u5__abc_54027_n837) );
  AND2X2 AND2X2_6079 ( .A(u5__abc_54027_n833_1), .B(u5__abc_54027_n340), .Y(u5__abc_54027_n838) );
  AND2X2 AND2X2_608 ( .A(u0__abc_49347_n1952_1_bF_buf3), .B(u0__abc_49347_n2190), .Y(u0__abc_49347_n2191) );
  AND2X2 AND2X2_6080 ( .A(u5__abc_54027_n839), .B(u5__abc_54027_n444), .Y(u5_ir_cnt_2__FF_INPUT) );
  AND2X2 AND2X2_6081 ( .A(u5__abc_54027_n841), .B(u5_ir_cnt_3_), .Y(u5__abc_54027_n842) );
  AND2X2 AND2X2_6082 ( .A(u5__abc_54027_n838), .B(u5__abc_54027_n339), .Y(u5__abc_54027_n843_1) );
  AND2X2 AND2X2_6083 ( .A(u5__abc_54027_n844), .B(u5__abc_54027_n444), .Y(u5_ir_cnt_3__FF_INPUT) );
  AND2X2 AND2X2_6084 ( .A(u5__abc_54027_n490), .B(u5__abc_54027_n598), .Y(u5__abc_54027_n847) );
  AND2X2 AND2X2_6085 ( .A(u5__abc_54027_n588), .B(u5__abc_54027_n847), .Y(u5__abc_54027_n848) );
  AND2X2 AND2X2_6086 ( .A(u5__abc_54027_n849), .B(u5__abc_54027_n376), .Y(u5__abc_54027_n850) );
  AND2X2 AND2X2_6087 ( .A(u5__abc_54027_n278), .B(u5__abc_54027_n389_1), .Y(u5__abc_54027_n852) );
  AND2X2 AND2X2_6088 ( .A(u5__abc_54027_n662), .B(u5__abc_54027_n853), .Y(u5__abc_54027_n854) );
  AND2X2 AND2X2_6089 ( .A(u5__abc_54027_n855_1), .B(u5__abc_54027_n425), .Y(u5__abc_54027_n856) );
  AND2X2 AND2X2_609 ( .A(u0__abc_49347_n2189), .B(u0__abc_49347_n2191), .Y(u0__abc_49347_n2192) );
  AND2X2 AND2X2_6090 ( .A(u5__abc_54027_n862), .B(u5_timer_0_), .Y(u5__abc_54027_n865) );
  AND2X2 AND2X2_6091 ( .A(u5__abc_54027_n427), .B(u5__abc_54027_n290_1), .Y(u5__abc_54027_n867) );
  AND2X2 AND2X2_6092 ( .A(u5__abc_54027_n389_1), .B(u5__abc_54027_n290_1), .Y(u5__abc_54027_n869_1) );
  AND2X2 AND2X2_6093 ( .A(u5__abc_54027_n870), .B(u5__abc_54027_n868_1), .Y(u5__abc_54027_n871) );
  AND2X2 AND2X2_6094 ( .A(u5__abc_54027_n270), .B(u5__abc_54027_n656), .Y(u5__abc_54027_n873) );
  AND2X2 AND2X2_6095 ( .A(u5__abc_54027_n876_1), .B(u5__abc_54027_n426), .Y(u5__abc_54027_n877) );
  AND2X2 AND2X2_6096 ( .A(u5__abc_54027_n861_1), .B(u5__abc_54027_n877), .Y(u5__abc_54027_n878) );
  AND2X2 AND2X2_6097 ( .A(u5__abc_54027_n879), .B(u5__abc_54027_n583), .Y(u5__abc_54027_n880) );
  AND2X2 AND2X2_6098 ( .A(u5__abc_54027_n574), .B(u5__abc_54027_n429_1), .Y(u5__abc_54027_n881) );
  AND2X2 AND2X2_6099 ( .A(u5__abc_54027_n578), .B(u5__abc_54027_n881), .Y(u5__abc_54027_n882_1) );
  AND2X2 AND2X2_61 ( .A(u0__abc_49347_n1100_1), .B(u0_lmr_req1), .Y(u0__abc_49347_n1109_1) );
  AND2X2 AND2X2_610 ( .A(u0__abc_49347_n1953_1_bF_buf3), .B(sp_csc_10_), .Y(u0__abc_49347_n2194) );
  AND2X2 AND2X2_6100 ( .A(u5__abc_54027_n884), .B(u5__abc_54027_n582), .Y(u5__abc_54027_n885) );
  AND2X2 AND2X2_6101 ( .A(u5__abc_54027_n889), .B(u5__abc_54027_n424), .Y(u5__abc_54027_n890) );
  AND2X2 AND2X2_6102 ( .A(u5__abc_54027_n887_1), .B(u5__abc_54027_n890), .Y(u5__abc_54027_n891) );
  AND2X2 AND2X2_6103 ( .A(u5__abc_54027_n888), .B(u5__abc_54027_n893), .Y(u5__abc_54027_n894) );
  AND2X2 AND2X2_6104 ( .A(u5__abc_54027_n896_1), .B(u5__abc_54027_n614), .Y(u5__abc_54027_n897_1) );
  AND2X2 AND2X2_6105 ( .A(u5__abc_54027_n897_1), .B(u5__abc_54027_n895_1), .Y(u5__abc_54027_n898_1) );
  AND2X2 AND2X2_6106 ( .A(u5__abc_54027_n900_1), .B(u5__abc_54027_n854), .Y(u5__abc_54027_n901) );
  AND2X2 AND2X2_6107 ( .A(u5__abc_54027_n901), .B(u5__abc_54027_n851), .Y(u5__abc_54027_n902) );
  AND2X2 AND2X2_6108 ( .A(u5__abc_54027_n588), .B(u5__abc_54027_n492), .Y(u5__abc_54027_n903) );
  AND2X2 AND2X2_6109 ( .A(u5__abc_54027_n904), .B(u5__abc_54027_n436), .Y(u5__abc_54027_n905_1) );
  AND2X2 AND2X2_611 ( .A(spec_req_cs_5_bF_buf2), .B(u0_csc5_10_), .Y(u0__abc_49347_n2195) );
  AND2X2 AND2X2_6110 ( .A(u5__abc_54027_n908), .B(u5__abc_54027_n907), .Y(u5__abc_54027_n909) );
  AND2X2 AND2X2_6111 ( .A(u5__abc_54027_n911), .B(u5__abc_54027_n913), .Y(u5_timer_0__FF_INPUT) );
  AND2X2 AND2X2_6112 ( .A(u5__abc_54027_n915), .B(u5__abc_54027_n906_1), .Y(u5__abc_54027_n916) );
  AND2X2 AND2X2_6113 ( .A(u5__abc_54027_n922), .B(u5__abc_54027_n921), .Y(u5__abc_54027_n923) );
  AND2X2 AND2X2_6114 ( .A(u5__abc_54027_n863), .B(u5_timer_1_), .Y(u5__abc_54027_n924) );
  AND2X2 AND2X2_6115 ( .A(u5__abc_54027_n926), .B(u5__abc_54027_n426), .Y(u5__abc_54027_n927) );
  AND2X2 AND2X2_6116 ( .A(u5__abc_54027_n927), .B(u5__abc_54027_n920), .Y(u5__abc_54027_n928) );
  AND2X2 AND2X2_6117 ( .A(u5__abc_54027_n929), .B(u5__abc_54027_n425), .Y(u5__abc_54027_n930) );
  AND2X2 AND2X2_6118 ( .A(u5__abc_54027_n932), .B(u5__abc_54027_n882_1), .Y(u5__abc_54027_n933) );
  AND2X2 AND2X2_6119 ( .A(u5__abc_54027_n933), .B(u5__abc_54027_n918), .Y(u5__abc_54027_n934) );
  AND2X2 AND2X2_612 ( .A(u0__abc_49347_n2197), .B(u0__abc_49347_n1185_bF_buf5), .Y(u0__abc_49347_n2198) );
  AND2X2 AND2X2_6120 ( .A(u5__abc_54027_n935), .B(u5__abc_54027_n883), .Y(u5__abc_54027_n936) );
  AND2X2 AND2X2_6121 ( .A(u5__abc_54027_n939), .B(u5__abc_54027_n935), .Y(u5__abc_54027_n940) );
  AND2X2 AND2X2_6122 ( .A(u5__abc_54027_n676), .B(u5__abc_54027_n942_1), .Y(u5__abc_54027_n943) );
  AND2X2 AND2X2_6123 ( .A(u5__abc_54027_n943), .B(u5__abc_54027_n941), .Y(u5__abc_54027_n944) );
  AND2X2 AND2X2_6124 ( .A(u5__abc_54027_n676), .B(u5__abc_54027_n941), .Y(u5__abc_54027_n947) );
  AND2X2 AND2X2_6125 ( .A(u5__abc_54027_n949), .B(u5__abc_54027_n948), .Y(u5__abc_54027_n950) );
  AND2X2 AND2X2_6126 ( .A(u5__abc_54027_n946), .B(u5__abc_54027_n951), .Y(u5__abc_54027_n952) );
  AND2X2 AND2X2_6127 ( .A(u5__abc_54027_n953_1), .B(u5__abc_54027_n850), .Y(u5__abc_54027_n954) );
  AND2X2 AND2X2_6128 ( .A(u5__abc_54027_n938), .B(u5__abc_54027_n954), .Y(u5__abc_54027_n955) );
  AND2X2 AND2X2_6129 ( .A(u5__abc_54027_n956), .B(u5__abc_54027_n892), .Y(u5__abc_54027_n957) );
  AND2X2 AND2X2_613 ( .A(u0__abc_49347_n2198), .B(u0__abc_49347_n2196), .Y(u0__abc_49347_n2199) );
  AND2X2 AND2X2_6130 ( .A(u5__abc_54027_n905_1), .B(u5__abc_54027_n854), .Y(u5__abc_54027_n960) );
  AND2X2 AND2X2_6131 ( .A(u5__abc_54027_n961), .B(u5__abc_54027_n905_1), .Y(u5__abc_54027_n962) );
  AND2X2 AND2X2_6132 ( .A(u5__abc_54027_n959), .B(u5__abc_54027_n963), .Y(u5__abc_54027_n964) );
  AND2X2 AND2X2_6133 ( .A(u5__abc_54027_n583), .B(u5__abc_54027_n426), .Y(u5__abc_54027_n968) );
  AND2X2 AND2X2_6134 ( .A(u5__abc_54027_n969), .B(u5__abc_54027_n858), .Y(u5__abc_54027_n970) );
  AND2X2 AND2X2_6135 ( .A(u5__abc_54027_n859), .B(u5__abc_54027_n971), .Y(u5__abc_54027_n972) );
  AND2X2 AND2X2_6136 ( .A(u5__abc_54027_n973), .B(u5_timer_2_), .Y(u5__abc_54027_n974) );
  AND2X2 AND2X2_6137 ( .A(u5__abc_54027_n923), .B(u5__abc_54027_n975), .Y(u5__abc_54027_n976) );
  AND2X2 AND2X2_6138 ( .A(u5__abc_54027_n978), .B(u5__abc_54027_n972), .Y(u5__abc_54027_n979) );
  AND2X2 AND2X2_6139 ( .A(u5__abc_54027_n980), .B(u5__abc_54027_n968), .Y(u5__abc_54027_n981) );
  AND2X2 AND2X2_614 ( .A(u0__abc_49347_n2200), .B(u0__abc_49347_n1181_bF_buf5), .Y(u0__abc_49347_n2201) );
  AND2X2 AND2X2_6140 ( .A(u5__abc_54027_n566_1), .B(u5__abc_54027_n582), .Y(u5__abc_54027_n982) );
  AND2X2 AND2X2_6141 ( .A(u5__abc_54027_n984), .B(u5__abc_54027_n967), .Y(u5__abc_54027_n985) );
  AND2X2 AND2X2_6142 ( .A(u5__abc_54027_n985), .B(u5__abc_54027_n424), .Y(u5__abc_54027_n986) );
  AND2X2 AND2X2_6143 ( .A(u5__abc_54027_n946), .B(u5__abc_54027_n948), .Y(u5__abc_54027_n988) );
  AND2X2 AND2X2_6144 ( .A(u5__abc_54027_n950), .B(u5__abc_54027_n894), .Y(u5__abc_54027_n990) );
  AND2X2 AND2X2_6145 ( .A(u5__abc_54027_n992), .B(u5__abc_54027_n614), .Y(u5__abc_54027_n993) );
  AND2X2 AND2X2_6146 ( .A(u5__abc_54027_n993), .B(u5__abc_54027_n989), .Y(u5__abc_54027_n994) );
  AND2X2 AND2X2_6147 ( .A(u5__abc_54027_n997), .B(u5__abc_54027_n854), .Y(u5__abc_54027_n998) );
  AND2X2 AND2X2_6148 ( .A(u5__abc_54027_n996), .B(u5__abc_54027_n998), .Y(u5__abc_54027_n999) );
  AND2X2 AND2X2_6149 ( .A(u5__abc_54027_n1000_1), .B(u5__abc_54027_n907), .Y(u5__abc_54027_n1001) );
  AND2X2 AND2X2_615 ( .A(spec_req_cs_4_bF_buf2), .B(u0_csc4_10_), .Y(u0__abc_49347_n2202) );
  AND2X2 AND2X2_6150 ( .A(u5__abc_54027_n1003), .B(u5__abc_54027_n1005), .Y(u5_timer_2__FF_INPUT) );
  AND2X2 AND2X2_6151 ( .A(u5__abc_54027_n893), .B(u5__abc_54027_n906_1), .Y(u5__abc_54027_n1007) );
  AND2X2 AND2X2_6152 ( .A(u5__abc_54027_n991), .B(u5__abc_54027_n966), .Y(u5__abc_54027_n1008) );
  AND2X2 AND2X2_6153 ( .A(u5__abc_54027_n1008), .B(u5__abc_54027_n1010), .Y(u5__abc_54027_n1011) );
  AND2X2 AND2X2_6154 ( .A(u5__abc_54027_n989), .B(u5__abc_54027_n1009), .Y(u5__abc_54027_n1012) );
  AND2X2 AND2X2_6155 ( .A(u5__abc_54027_n1015), .B(u5__abc_54027_n858), .Y(u5__abc_54027_n1016) );
  AND2X2 AND2X2_6156 ( .A(u5__abc_54027_n923), .B(u5__abc_54027_n326), .Y(u5__abc_54027_n1018) );
  AND2X2 AND2X2_6157 ( .A(u5__abc_54027_n1019), .B(u5_timer_3_), .Y(u5__abc_54027_n1020) );
  AND2X2 AND2X2_6158 ( .A(u5__abc_54027_n1021), .B(u5__abc_54027_n1017), .Y(u5__abc_54027_n1022) );
  AND2X2 AND2X2_6159 ( .A(u5__abc_54027_n882_1), .B(u5__abc_54027_n968), .Y(u5__abc_54027_n1024) );
  AND2X2 AND2X2_616 ( .A(u0__abc_49347_n2203), .B(u0__abc_49347_n1180_1_bF_buf5), .Y(u0__abc_49347_n2204) );
  AND2X2 AND2X2_6160 ( .A(u5__abc_54027_n1023), .B(u5__abc_54027_n1024), .Y(u5__abc_54027_n1025) );
  AND2X2 AND2X2_6161 ( .A(u5__abc_54027_n1009), .B(u5__abc_54027_n883), .Y(u5__abc_54027_n1026) );
  AND2X2 AND2X2_6162 ( .A(u5__abc_54027_n1028), .B(u5__abc_54027_n850), .Y(u5__abc_54027_n1029) );
  AND2X2 AND2X2_6163 ( .A(u5__abc_54027_n1014), .B(u5__abc_54027_n1029), .Y(u5__abc_54027_n1030) );
  AND2X2 AND2X2_6164 ( .A(u5__abc_54027_n1031), .B(u5__abc_54027_n892), .Y(u5__abc_54027_n1032) );
  AND2X2 AND2X2_6165 ( .A(u5__abc_54027_n1035), .B(u5__abc_54027_n905_1), .Y(u5__abc_54027_n1036) );
  AND2X2 AND2X2_6166 ( .A(u5__abc_54027_n1034), .B(u5__abc_54027_n1037), .Y(u5__abc_54027_n1038) );
  AND2X2 AND2X2_6167 ( .A(u5__abc_54027_n326), .B(u5__abc_54027_n921), .Y(u5__abc_54027_n1040) );
  AND2X2 AND2X2_6168 ( .A(u5__abc_54027_n1040), .B(u5__abc_54027_n328_1), .Y(u5__abc_54027_n1041) );
  AND2X2 AND2X2_6169 ( .A(u5__abc_54027_n922), .B(u5__abc_54027_n1041), .Y(u5__abc_54027_n1042) );
  AND2X2 AND2X2_617 ( .A(spec_req_cs_3_bF_buf2), .B(u0_csc3_10_), .Y(u0__abc_49347_n2205) );
  AND2X2 AND2X2_6170 ( .A(u5__abc_54027_n1043), .B(u5_timer_4_), .Y(u5__abc_54027_n1044) );
  AND2X2 AND2X2_6171 ( .A(u5__abc_54027_n426), .B(u5__abc_54027_n971), .Y(u5__abc_54027_n1046) );
  AND2X2 AND2X2_6172 ( .A(u5__abc_54027_n424), .B(u5__abc_54027_n1046), .Y(u5__abc_54027_n1047) );
  AND2X2 AND2X2_6173 ( .A(u5__abc_54027_n871), .B(u5__abc_54027_n583), .Y(u5__abc_54027_n1048) );
  AND2X2 AND2X2_6174 ( .A(u5__abc_54027_n1047), .B(u5__abc_54027_n1048), .Y(u5__abc_54027_n1049) );
  AND2X2 AND2X2_6175 ( .A(u5__abc_54027_n859), .B(u5__abc_54027_n1049), .Y(u5__abc_54027_n1050) );
  AND2X2 AND2X2_6176 ( .A(u5__abc_54027_n1050), .B(u5__abc_54027_n882_1), .Y(u5__abc_54027_n1051) );
  AND2X2 AND2X2_6177 ( .A(u5__abc_54027_n1051), .B(u5__abc_54027_n850), .Y(u5__abc_54027_n1052_1) );
  AND2X2 AND2X2_6178 ( .A(u5__abc_54027_n1052_1), .B(u5__abc_54027_n1045), .Y(u5__abc_54027_n1053_1) );
  AND2X2 AND2X2_6179 ( .A(u5__abc_54027_n855_1), .B(u5__abc_54027_n892), .Y(u5__abc_54027_n1054) );
  AND2X2 AND2X2_618 ( .A(u0__abc_49347_n2206), .B(u0__abc_49347_n1179_bF_buf5), .Y(u0__abc_49347_n2207) );
  AND2X2 AND2X2_6180 ( .A(u5__abc_54027_n1055), .B(u5__abc_54027_n960), .Y(u5_timer_4__FF_INPUT) );
  AND2X2 AND2X2_6181 ( .A(u5__abc_54027_n1042), .B(u5__abc_54027_n327), .Y(u5__abc_54027_n1057) );
  AND2X2 AND2X2_6182 ( .A(u5__abc_54027_n1058_1), .B(u5_timer_5_), .Y(u5__abc_54027_n1059) );
  AND2X2 AND2X2_6183 ( .A(u5__abc_54027_n1052_1), .B(u5__abc_54027_n1060), .Y(u5__abc_54027_n1061) );
  AND2X2 AND2X2_6184 ( .A(u5__abc_54027_n929), .B(u5__abc_54027_n892), .Y(u5__abc_54027_n1062) );
  AND2X2 AND2X2_6185 ( .A(u5__abc_54027_n1063), .B(u5__abc_54027_n960), .Y(u5_timer_5__FF_INPUT) );
  AND2X2 AND2X2_6186 ( .A(u5__abc_54027_n1065), .B(u5__abc_54027_n892), .Y(u5__abc_54027_n1066) );
  AND2X2 AND2X2_6187 ( .A(u5__abc_54027_n1067), .B(u5_timer_6_), .Y(u5__abc_54027_n1068) );
  AND2X2 AND2X2_6188 ( .A(u5__abc_54027_n330_1), .B(u5__abc_54027_n921), .Y(u5__abc_54027_n1070) );
  AND2X2 AND2X2_6189 ( .A(u5__abc_54027_n1070), .B(u5__abc_54027_n1069), .Y(u5__abc_54027_n1071) );
  AND2X2 AND2X2_619 ( .A(spec_req_cs_2_bF_buf2), .B(u0_csc2_10_), .Y(u0__abc_49347_n2208) );
  AND2X2 AND2X2_6190 ( .A(u5__abc_54027_n922), .B(u5__abc_54027_n1071), .Y(u5__abc_54027_n1072) );
  AND2X2 AND2X2_6191 ( .A(u5__abc_54027_n1052_1), .B(u5__abc_54027_n1073), .Y(u5__abc_54027_n1074) );
  AND2X2 AND2X2_6192 ( .A(u5__abc_54027_n1075), .B(u5__abc_54027_n960), .Y(u5_timer_6__FF_INPUT) );
  AND2X2 AND2X2_6193 ( .A(u5__abc_54027_n1077), .B(u5__abc_54027_n892), .Y(u5__abc_54027_n1078) );
  AND2X2 AND2X2_6194 ( .A(u5__abc_54027_n1079), .B(u5_timer_7_), .Y(u5__abc_54027_n1080) );
  AND2X2 AND2X2_6195 ( .A(u5__abc_54027_n1052_1), .B(u5__abc_54027_n1080), .Y(u5__abc_54027_n1081) );
  AND2X2 AND2X2_6196 ( .A(u5__abc_54027_n1082), .B(u5__abc_54027_n960), .Y(u5_timer_7__FF_INPUT) );
  AND2X2 AND2X2_6197 ( .A(u5__abc_54027_n351_bF_buf1), .B(u5__abc_54027_n490), .Y(u5__abc_54027_n1084) );
  AND2X2 AND2X2_6198 ( .A(u5__abc_54027_n939), .B(u5__abc_54027_n1084), .Y(u5__abc_54027_n1085) );
  AND2X2 AND2X2_6199 ( .A(u5__abc_54027_n594), .B(csc_s_1_), .Y(u5__abc_54027_n1086) );
  AND2X2 AND2X2_62 ( .A(init_req), .B(u0_init_req1), .Y(u0__abc_49347_n1110) );
  AND2X2 AND2X2_620 ( .A(u0__abc_49347_n2209), .B(u0__abc_49347_n1178_1_bF_buf5), .Y(u0__abc_49347_n2210) );
  AND2X2 AND2X2_6200 ( .A(u5__abc_54027_n351_bF_buf0), .B(u5__abc_54027_n1086), .Y(u5__abc_54027_n1087) );
  AND2X2 AND2X2_6201 ( .A(u5__abc_54027_n1091), .B(u5__abc_54027_n433_1), .Y(u5__abc_54027_n1092) );
  AND2X2 AND2X2_6202 ( .A(u5__abc_54027_n912), .B(u5__abc_54027_n1093), .Y(u5__abc_54027_n1094) );
  AND2X2 AND2X2_6203 ( .A(u5__abc_54027_n1103), .B(u5__abc_54027_n1095), .Y(u5__abc_54027_n1104) );
  AND2X2 AND2X2_6204 ( .A(u5__abc_54027_n388_1), .B(u5__abc_54027_n398), .Y(u5__abc_54027_n1105) );
  AND2X2 AND2X2_6205 ( .A(u5__abc_54027_n1105), .B(u5__abc_54027_n368), .Y(u5__abc_54027_n1106) );
  AND2X2 AND2X2_6206 ( .A(u5__abc_54027_n1106), .B(u5__abc_54027_n659), .Y(u5__abc_54027_n1107) );
  AND2X2 AND2X2_6207 ( .A(u5__abc_54027_n430_1), .B(u5_tmr2_done), .Y(u5__abc_54027_n1110) );
  AND2X2 AND2X2_6208 ( .A(u5__abc_54027_n1092), .B(u5__abc_54027_n1111), .Y(u5__abc_54027_n1112) );
  AND2X2 AND2X2_6209 ( .A(u5__abc_54027_n1113), .B(u5__abc_54027_n1112), .Y(u5__abc_54027_n1114) );
  AND2X2 AND2X2_621 ( .A(spec_req_cs_1_bF_buf2), .B(u0_csc1_10_), .Y(u0__abc_49347_n2211) );
  AND2X2 AND2X2_6210 ( .A(u5__abc_54027_n1114), .B(u5__abc_54027_n1109), .Y(u5__abc_54027_n1115) );
  AND2X2 AND2X2_6211 ( .A(u5__abc_54027_n1116), .B(u5__abc_54027_n1090), .Y(u5__abc_54027_n1117) );
  AND2X2 AND2X2_6212 ( .A(u5_timer2_1_), .B(u5_timer2_0_), .Y(u5__abc_54027_n1120) );
  AND2X2 AND2X2_6213 ( .A(u5__abc_54027_n1106), .B(u5__abc_54027_n1121), .Y(u5__abc_54027_n1122) );
  AND2X2 AND2X2_6214 ( .A(u5__abc_54027_n1103), .B(u5__abc_54027_n1122), .Y(u5__abc_54027_n1123) );
  AND2X2 AND2X2_6215 ( .A(u5__abc_54027_n846), .B(u5__abc_54027_n1124), .Y(u5__abc_54027_n1125) );
  AND2X2 AND2X2_6216 ( .A(u5__abc_54027_n1127), .B(u5__abc_54027_n1128), .Y(u5__abc_54027_n1129) );
  AND2X2 AND2X2_6217 ( .A(u5__abc_54027_n1130), .B(u5__abc_54027_n1131), .Y(u5__abc_54027_n1132) );
  AND2X2 AND2X2_6218 ( .A(u5__abc_54027_n1133), .B(u5__abc_54027_n1134), .Y(u5__abc_54027_n1135) );
  AND2X2 AND2X2_6219 ( .A(u5__abc_54027_n1137), .B(u5__abc_54027_n1090), .Y(u5__abc_54027_n1138) );
  AND2X2 AND2X2_622 ( .A(u0__abc_49347_n1952_1_bF_buf2), .B(u0__abc_49347_n2214), .Y(u0__abc_49347_n2215) );
  AND2X2 AND2X2_6220 ( .A(u5__abc_54027_n1136), .B(u5__abc_54027_n1138), .Y(u5__abc_54027_n1139) );
  AND2X2 AND2X2_6221 ( .A(u5__abc_54027_n884), .B(u5__abc_54027_n1084), .Y(u5__abc_54027_n1140) );
  AND2X2 AND2X2_6222 ( .A(u5__abc_54027_n956), .B(u5__abc_54027_n1124), .Y(u5__abc_54027_n1144) );
  AND2X2 AND2X2_6223 ( .A(u5__abc_54027_n1096), .B(u5_timer2_2_), .Y(u5__abc_54027_n1146) );
  AND2X2 AND2X2_6224 ( .A(u5__abc_54027_n1106), .B(u5__abc_54027_n1147), .Y(u5__abc_54027_n1148) );
  AND2X2 AND2X2_6225 ( .A(u5__abc_54027_n1103), .B(u5__abc_54027_n1148), .Y(u5__abc_54027_n1149) );
  AND2X2 AND2X2_6226 ( .A(u5__abc_54027_n1150), .B(u5__abc_54027_n655), .Y(u5__abc_54027_n1151) );
  AND2X2 AND2X2_6227 ( .A(u5__abc_54027_n961), .B(u5__abc_54027_n654_1), .Y(u5__abc_54027_n1152) );
  AND2X2 AND2X2_6228 ( .A(u5__abc_54027_n1155), .B(u5__abc_54027_n1111), .Y(u5__abc_54027_n1156) );
  AND2X2 AND2X2_6229 ( .A(u5__abc_54027_n1154), .B(u5__abc_54027_n1156), .Y(u5__abc_54027_n1157) );
  AND2X2 AND2X2_623 ( .A(u0__abc_49347_n2213), .B(u0__abc_49347_n2215), .Y(u0__abc_49347_n2216_1) );
  AND2X2 AND2X2_6230 ( .A(u5__abc_54027_n884), .B(u5__abc_54027_n1110), .Y(u5__abc_54027_n1158) );
  AND2X2 AND2X2_6231 ( .A(u5__abc_54027_n1159), .B(u5__abc_54027_n1092), .Y(u5__abc_54027_n1160) );
  AND2X2 AND2X2_6232 ( .A(u5__abc_54027_n1004), .B(u5__abc_54027_n1093), .Y(u5__abc_54027_n1161) );
  AND2X2 AND2X2_6233 ( .A(u5__abc_54027_n1163), .B(u5__abc_54027_n1143), .Y(u5_timer2_2__FF_INPUT) );
  AND2X2 AND2X2_6234 ( .A(u5__abc_54027_n1097), .B(u5_timer2_3_), .Y(u5__abc_54027_n1166) );
  AND2X2 AND2X2_6235 ( .A(u5__abc_54027_n1106), .B(u5__abc_54027_n1167), .Y(u5__abc_54027_n1168) );
  AND2X2 AND2X2_6236 ( .A(u5__abc_54027_n1103), .B(u5__abc_54027_n1168), .Y(u5__abc_54027_n1169) );
  AND2X2 AND2X2_6237 ( .A(u5__abc_54027_n709_1), .B(u5__abc_54027_n1124), .Y(u5__abc_54027_n1170) );
  AND2X2 AND2X2_6238 ( .A(u5__abc_54027_n1172), .B(u5__abc_54027_n1173), .Y(u5__abc_54027_n1174) );
  AND2X2 AND2X2_6239 ( .A(u5__abc_54027_n1175), .B(u5__abc_54027_n1176), .Y(u5__abc_54027_n1177) );
  AND2X2 AND2X2_624 ( .A(u0__abc_49347_n1176_1_bF_buf6), .B(tms_0_), .Y(u0__abc_49347_n2722) );
  AND2X2 AND2X2_6240 ( .A(u5__abc_54027_n1177), .B(u5__abc_54027_n1111), .Y(u5__abc_54027_n1178) );
  AND2X2 AND2X2_6241 ( .A(u5__abc_54027_n917), .B(u5__abc_54027_n1110), .Y(u5__abc_54027_n1179) );
  AND2X2 AND2X2_6242 ( .A(u5__abc_54027_n1182), .B(u5__abc_54027_n1090), .Y(u5__abc_54027_n1183) );
  AND2X2 AND2X2_6243 ( .A(u5__abc_54027_n1181), .B(u5__abc_54027_n1183), .Y(u5__abc_54027_n1184) );
  AND2X2 AND2X2_6244 ( .A(u5__abc_54027_n566_1), .B(u5__abc_54027_n1084), .Y(u5__abc_54027_n1185) );
  AND2X2 AND2X2_6245 ( .A(u5__abc_54027_n888), .B(u5__abc_54027_n1084), .Y(u5__abc_54027_n1187) );
  AND2X2 AND2X2_6246 ( .A(u5__abc_54027_n1090), .B(u5__abc_54027_n1092), .Y(u5__abc_54027_n1188) );
  AND2X2 AND2X2_6247 ( .A(u5__abc_54027_n1031), .B(u5__abc_54027_n1124), .Y(u5__abc_54027_n1190) );
  AND2X2 AND2X2_6248 ( .A(u5__abc_54027_n1098), .B(u5_timer2_4_), .Y(u5__abc_54027_n1192) );
  AND2X2 AND2X2_6249 ( .A(u5__abc_54027_n1193), .B(u5__abc_54027_n1106), .Y(u5__abc_54027_n1194) );
  AND2X2 AND2X2_625 ( .A(u0_tms5_0_), .B(u0_cs5_bF_buf5), .Y(u0__abc_49347_n2727) );
  AND2X2 AND2X2_6250 ( .A(u5__abc_54027_n1103), .B(u5__abc_54027_n1194), .Y(u5__abc_54027_n1195) );
  AND2X2 AND2X2_6251 ( .A(u5__abc_54027_n1196), .B(u5__abc_54027_n655), .Y(u5__abc_54027_n1197) );
  AND2X2 AND2X2_6252 ( .A(u5__abc_54027_n1035), .B(u5__abc_54027_n654_1), .Y(u5__abc_54027_n1198) );
  AND2X2 AND2X2_6253 ( .A(u5__abc_54027_n1199), .B(u5__abc_54027_n658), .Y(u5__abc_54027_n1200) );
  AND2X2 AND2X2_6254 ( .A(u5__abc_54027_n860), .B(u5__abc_54027_n657_1), .Y(u5__abc_54027_n1201) );
  AND2X2 AND2X2_6255 ( .A(u5__abc_54027_n1203), .B(u5__abc_54027_n1189), .Y(u5__abc_54027_n1204) );
  AND2X2 AND2X2_6256 ( .A(u5__abc_54027_n1204), .B(u5__abc_54027_n1188), .Y(u5__abc_54027_n1205_1) );
  AND2X2 AND2X2_6257 ( .A(u5__abc_54027_n935), .B(u5__abc_54027_n1084), .Y(u5__abc_54027_n1207) );
  AND2X2 AND2X2_6258 ( .A(u5__abc_54027_n919), .B(u5__abc_54027_n657_1), .Y(u5__abc_54027_n1208) );
  AND2X2 AND2X2_6259 ( .A(u5__abc_54027_n1099), .B(u5_timer2_5_), .Y(u5__abc_54027_n1210) );
  AND2X2 AND2X2_626 ( .A(u0__abc_49347_n2731), .B(u0__abc_49347_n2730_bF_buf5), .Y(u0__abc_49347_n2732) );
  AND2X2 AND2X2_6260 ( .A(u5__abc_54027_n1211), .B(u5__abc_54027_n1106), .Y(u5__abc_54027_n1212) );
  AND2X2 AND2X2_6261 ( .A(u5__abc_54027_n1103), .B(u5__abc_54027_n1212), .Y(u5__abc_54027_n1213) );
  AND2X2 AND2X2_6262 ( .A(u5__abc_54027_n855_1), .B(u5__abc_54027_n1124), .Y(u5__abc_54027_n1214) );
  AND2X2 AND2X2_6263 ( .A(u5__abc_54027_n1215), .B(u5__abc_54027_n659), .Y(u5__abc_54027_n1216) );
  AND2X2 AND2X2_6264 ( .A(u5__abc_54027_n1090), .B(u5__abc_54027_n1112), .Y(u5__abc_54027_n1218) );
  AND2X2 AND2X2_6265 ( .A(u5__abc_54027_n1217), .B(u5__abc_54027_n1218), .Y(u5__abc_54027_n1219) );
  AND2X2 AND2X2_6266 ( .A(u5__abc_54027_n966), .B(u5__abc_54027_n1084), .Y(u5__abc_54027_n1221) );
  AND2X2 AND2X2_6267 ( .A(u5__abc_54027_n1100), .B(u5_timer2_6_), .Y(u5__abc_54027_n1223) );
  AND2X2 AND2X2_6268 ( .A(u5__abc_54027_n1103), .B(u5__abc_54027_n1224), .Y(u5__abc_54027_n1225) );
  AND2X2 AND2X2_6269 ( .A(u5__abc_54027_n1218), .B(u5__abc_54027_n659), .Y(u5__abc_54027_n1227) );
  AND2X2 AND2X2_627 ( .A(u0__abc_49347_n2732), .B(u0__abc_49347_n2729), .Y(u0__abc_49347_n2733) );
  AND2X2 AND2X2_6270 ( .A(u5__abc_54027_n1228), .B(u5__abc_54027_n1227), .Y(u5__abc_54027_n1229) );
  AND2X2 AND2X2_6271 ( .A(u5__abc_54027_n1229), .B(u5__abc_54027_n1226), .Y(u5__abc_54027_n1230) );
  AND2X2 AND2X2_6272 ( .A(u5__abc_54027_n1009), .B(u5__abc_54027_n1084), .Y(u5__abc_54027_n1232) );
  AND2X2 AND2X2_6273 ( .A(u5__abc_54027_n1234), .B(u5_timer2_8_), .Y(u5__abc_54027_n1235_1) );
  AND2X2 AND2X2_6274 ( .A(u5__abc_54027_n1101), .B(u5_timer2_7_), .Y(u5__abc_54027_n1236) );
  AND2X2 AND2X2_6275 ( .A(u5__abc_54027_n1238), .B(u5__abc_54027_n1233_1), .Y(u5__abc_54027_n1239) );
  AND2X2 AND2X2_6276 ( .A(u5__abc_54027_n1239), .B(u5__abc_54027_n1227), .Y(u5__abc_54027_n1240) );
  AND2X2 AND2X2_6277 ( .A(u5__abc_54027_n860), .B(u5__abc_54027_n1084), .Y(u5__abc_54027_n1242) );
  AND2X2 AND2X2_6278 ( .A(u5__abc_54027_n1102), .B(u5_timer2_8_), .Y(u5__abc_54027_n1244) );
  AND2X2 AND2X2_6279 ( .A(u5__abc_54027_n1245), .B(u5__abc_54027_n1227), .Y(u5__abc_54027_n1246) );
  AND2X2 AND2X2_628 ( .A(u0__abc_49347_n2734), .B(u0__abc_49347_n2726_bF_buf5), .Y(u0__abc_49347_n2735) );
  AND2X2 AND2X2_6280 ( .A(u5__abc_54027_n1246), .B(u5__abc_54027_n1243), .Y(u5__abc_54027_n1247) );
  AND2X2 AND2X2_6281 ( .A(u5__abc_54027_n643_1), .B(dv), .Y(u5__abc_54027_n1249) );
  AND2X2 AND2X2_6282 ( .A(u5__abc_54027_n1256), .B(u5__abc_54027_n1255), .Y(u5__abc_54027_n1257) );
  AND2X2 AND2X2_6283 ( .A(u5__abc_54027_n1257), .B(u5__abc_54027_n1254), .Y(u5_ack_cnt_0__FF_INPUT) );
  AND2X2 AND2X2_6284 ( .A(u5__abc_54027_n1251), .B(u5__abc_54027_n637), .Y(u5__abc_54027_n1259) );
  AND2X2 AND2X2_6285 ( .A(u5__abc_54027_n1249), .B(u5_ack_cnt_0_), .Y(u5__abc_54027_n1260) );
  AND2X2 AND2X2_6286 ( .A(u5__abc_54027_n1264), .B(u5__abc_54027_n1255), .Y(u5__abc_54027_n1265) );
  AND2X2 AND2X2_6287 ( .A(u5__abc_54027_n1265), .B(u5__abc_54027_n1263), .Y(u5_ack_cnt_1__FF_INPUT) );
  AND2X2 AND2X2_6288 ( .A(u5__abc_54027_n1251), .B(u5__abc_54027_n638_1), .Y(u5__abc_54027_n1267) );
  AND2X2 AND2X2_6289 ( .A(u5_ack_cnt_1_), .B(u5_ack_cnt_0_), .Y(u5__abc_54027_n1268) );
  AND2X2 AND2X2_629 ( .A(u0_tms4_0_), .B(u0_cs4_bF_buf4), .Y(u0__abc_49347_n2736) );
  AND2X2 AND2X2_6290 ( .A(u5__abc_54027_n1249), .B(u5__abc_54027_n1268), .Y(u5__abc_54027_n1269) );
  AND2X2 AND2X2_6291 ( .A(u5__abc_54027_n1273), .B(u5__abc_54027_n1255), .Y(u5__abc_54027_n1274) );
  AND2X2 AND2X2_6292 ( .A(u5__abc_54027_n1274), .B(u5__abc_54027_n1272), .Y(u5_ack_cnt_2__FF_INPUT) );
  AND2X2 AND2X2_6293 ( .A(u5__abc_54027_n1277), .B(u5_ack_cnt_3_), .Y(u5__abc_54027_n1278) );
  AND2X2 AND2X2_6294 ( .A(u5__abc_54027_n1269), .B(u5_ack_cnt_2_), .Y(u5__abc_54027_n1279) );
  AND2X2 AND2X2_6295 ( .A(u5__abc_54027_n1279), .B(u5_ack_cnt_3_), .Y(u5__abc_54027_n1281) );
  AND2X2 AND2X2_6296 ( .A(u5__abc_54027_n1282), .B(u5__abc_54027_n1255), .Y(u5__abc_54027_n1283) );
  AND2X2 AND2X2_6297 ( .A(u5__abc_54027_n1283), .B(u5__abc_54027_n1280), .Y(u5_ack_cnt_3__FF_INPUT) );
  AND2X2 AND2X2_6298 ( .A(u5__abc_54027_n1286), .B(u5__abc_54027_n1285), .Y(u5_cmd_asserted2_FF_INPUT) );
  AND2X2 AND2X2_6299 ( .A(u5_mc_le), .B(u5_cmd_asserted_bF_buf2), .Y(u5__abc_54027_n1288) );
  AND2X2 AND2X2_63 ( .A(u0__abc_49347_n1105_1), .B(u0__abc_49347_n1111_1), .Y(u0__abc_49347_n1112) );
  AND2X2 AND2X2_630 ( .A(u0__abc_49347_n2737), .B(u0__abc_49347_n2725_bF_buf5), .Y(u0__abc_49347_n2738) );
  AND2X2 AND2X2_6300 ( .A(u5_cmd_3_), .B(u5_mc_le_FF_INPUT), .Y(u5__abc_54027_n1289) );
  AND2X2 AND2X2_6301 ( .A(u5__abc_54027_n1292), .B(u5__abc_54027_n1291), .Y(u5_mc_adv_r_FF_INPUT) );
  AND2X2 AND2X2_6302 ( .A(u5__abc_54027_n278), .B(u5__abc_54027_n343), .Y(u5__abc_54027_n1295) );
  AND2X2 AND2X2_6303 ( .A(u5__abc_54027_n1294), .B(u5__abc_54027_n1296), .Y(u5__abc_54027_n1297) );
  AND2X2 AND2X2_6304 ( .A(u5__abc_54027_n1295), .B(u5__abc_54027_n1299), .Y(u5__abc_54027_n1300) );
  AND2X2 AND2X2_6305 ( .A(u5__abc_54027_n1298), .B(u5__abc_54027_n1301), .Y(mc_adv_d) );
  AND2X2 AND2X2_6306 ( .A(u5__abc_54027_n1303), .B(u5__abc_54027_n1304), .Y(u5_mc_adv_r1_FF_INPUT) );
  AND2X2 AND2X2_6307 ( .A(u5_wb_cycle), .B(u1_wb_write_go), .Y(u5__abc_54027_n1308) );
  AND2X2 AND2X2_6308 ( .A(u5__abc_54027_n1307), .B(u5__abc_54027_n1309), .Y(u5__abc_54027_n1310) );
  AND2X2 AND2X2_6309 ( .A(u5__abc_54027_n428), .B(u5__abc_54027_n1312_1), .Y(u5__abc_54027_n1313) );
  AND2X2 AND2X2_631 ( .A(u0_tms3_0_), .B(u0_cs3_bF_buf4), .Y(u0__abc_49347_n2739) );
  AND2X2 AND2X2_6310 ( .A(u5__abc_54027_n1311), .B(u5__abc_54027_n1314), .Y(u5__abc_54027_n1315) );
  AND2X2 AND2X2_6311 ( .A(u5__abc_54027_n473), .B(u5__abc_54027_n506), .Y(u5__abc_54027_n1316) );
  AND2X2 AND2X2_6312 ( .A(u5__abc_54027_n483), .B(u5__abc_54027_n420), .Y(u5__abc_54027_n1318) );
  AND2X2 AND2X2_6313 ( .A(u5__abc_54027_n1318), .B(u5__abc_54027_n1317), .Y(u5__abc_54027_n1319) );
  AND2X2 AND2X2_6314 ( .A(u5__abc_54027_n476), .B(u5__abc_54027_n1319), .Y(u5__abc_54027_n1320) );
  AND2X2 AND2X2_6315 ( .A(u5__abc_54027_n680), .B(u5__abc_54027_n501), .Y(u5__abc_54027_n1321) );
  AND2X2 AND2X2_6316 ( .A(u5__abc_54027_n475_1), .B(u5__abc_54027_n1321), .Y(u5__abc_54027_n1322) );
  AND2X2 AND2X2_6317 ( .A(u5__abc_54027_n1315), .B(u5__abc_54027_n1324), .Y(u5__abc_54027_n1325) );
  AND2X2 AND2X2_6318 ( .A(u5__abc_54027_n1326), .B(u3_wb_read_go), .Y(u5__abc_54027_n1327) );
  AND2X2 AND2X2_6319 ( .A(u5__abc_54027_n1328), .B(u5__abc_54027_n319), .Y(u5__abc_54027_n1329) );
  AND2X2 AND2X2_632 ( .A(u0__abc_49347_n2740), .B(u0__abc_49347_n2724_bF_buf5), .Y(u0__abc_49347_n2741) );
  AND2X2 AND2X2_6320 ( .A(u5__abc_54027_n278), .B(u5__abc_54027_n296), .Y(u5__abc_54027_n1330) );
  AND2X2 AND2X2_6321 ( .A(u5__abc_54027_n641), .B(u3_wb_read_go), .Y(u5__abc_54027_n1331) );
  AND2X2 AND2X2_6322 ( .A(u5__abc_54027_n1331), .B(u5__abc_54027_n1330), .Y(u5__abc_54027_n1332) );
  AND2X2 AND2X2_6323 ( .A(u5__abc_54027_n303), .B(u5__abc_54027_n312_1), .Y(u5__abc_54027_n1335) );
  AND2X2 AND2X2_6324 ( .A(u5__abc_54027_n1335), .B(u5_tmr_done), .Y(u5__abc_54027_n1336) );
  AND2X2 AND2X2_6325 ( .A(u5__abc_54027_n313_1), .B(u5__abc_54027_n1309), .Y(u5__abc_54027_n1338) );
  AND2X2 AND2X2_6326 ( .A(u5__abc_54027_n1338), .B(u5_wb_cycle), .Y(u5__abc_54027_n1339) );
  AND2X2 AND2X2_6327 ( .A(u5__abc_54027_n1341_1), .B(u5__abc_54027_n1337), .Y(u5__abc_54027_n1342) );
  AND2X2 AND2X2_6328 ( .A(u5__abc_54027_n422), .B(u5__abc_54027_n1312_1), .Y(u5__abc_54027_n1343) );
  AND2X2 AND2X2_6329 ( .A(u5__abc_54027_n1346), .B(csc_s_4_), .Y(u5__abc_54027_n1347) );
  AND2X2 AND2X2_633 ( .A(u0_tms2_0_), .B(u0_cs2_bF_buf4), .Y(u0__abc_49347_n2742) );
  AND2X2 AND2X2_6330 ( .A(u5__abc_54027_n377), .B(u5__abc_54027_n1347), .Y(u5__abc_54027_n1348) );
  AND2X2 AND2X2_6331 ( .A(u5__abc_54027_n1349), .B(u5_tmr2_done), .Y(u5__abc_54027_n1350) );
  AND2X2 AND2X2_6332 ( .A(u5__abc_54027_n508), .B(u5__abc_54027_n510), .Y(u5__abc_54027_n1353) );
  AND2X2 AND2X2_6333 ( .A(u5__abc_54027_n1352), .B(u5__abc_54027_n1353), .Y(u5__abc_54027_n1354) );
  AND2X2 AND2X2_6334 ( .A(u5__abc_54027_n351_bF_buf3), .B(u5__abc_54027_n513_1), .Y(u5__abc_54027_n1356) );
  AND2X2 AND2X2_6335 ( .A(u5__abc_54027_n1361), .B(u5__abc_54027_n1351), .Y(u5__abc_54027_n1362) );
  AND2X2 AND2X2_6336 ( .A(u5__abc_54027_n1362), .B(u5__abc_54027_n1345), .Y(u5__abc_54027_n1363) );
  AND2X2 AND2X2_6337 ( .A(u5__abc_54027_n869_1), .B(u5_resume_req_r), .Y(u5__abc_54027_n1364_1) );
  AND2X2 AND2X2_6338 ( .A(u5__abc_54027_n384), .B(u5_tmr2_done), .Y(u5__abc_54027_n1366) );
  AND2X2 AND2X2_6339 ( .A(u5__abc_54027_n1365), .B(u5__abc_54027_n1367), .Y(u5__abc_54027_n1368) );
  AND2X2 AND2X2_634 ( .A(u0__abc_49347_n2743), .B(u0__abc_49347_n2723_bF_buf5), .Y(u0__abc_49347_n2744) );
  AND2X2 AND2X2_6340 ( .A(u5__abc_54027_n377), .B(u5_tmr2_done), .Y(u5__abc_54027_n1370) );
  AND2X2 AND2X2_6341 ( .A(u5__abc_54027_n1372), .B(u5__abc_54027_n1368), .Y(u5__abc_54027_n1373_1) );
  AND2X2 AND2X2_6342 ( .A(u5__abc_54027_n1374), .B(u5__abc_54027_n400), .Y(u5__abc_54027_n1375) );
  AND2X2 AND2X2_6343 ( .A(u5__abc_54027_n369), .B(u5_cmd_asserted_bF_buf0), .Y(u5__abc_54027_n1376) );
  AND2X2 AND2X2_6344 ( .A(u5__abc_54027_n1378_1), .B(u5__abc_54027_n1375), .Y(u5__abc_54027_n1379) );
  AND2X2 AND2X2_6345 ( .A(u5__abc_54027_n1379), .B(u5__abc_54027_n1373_1), .Y(u5__abc_54027_n1380_1) );
  AND2X2 AND2X2_6346 ( .A(u5__abc_54027_n360), .B(u5_tmr2_done), .Y(u5__abc_54027_n1381_1) );
  AND2X2 AND2X2_6347 ( .A(u5__abc_54027_n294), .B(u5__abc_54027_n1383_1), .Y(u5__abc_54027_n1384) );
  AND2X2 AND2X2_6348 ( .A(u5__abc_54027_n511), .B(init_req), .Y(u5__abc_54027_n1386) );
  AND2X2 AND2X2_6349 ( .A(u5__abc_54027_n351_bF_buf2), .B(u5__abc_54027_n1386), .Y(u5__abc_54027_n1387) );
  AND2X2 AND2X2_635 ( .A(u0_tms1_0_), .B(u0_cs1_bF_buf4), .Y(u0__abc_49347_n2745) );
  AND2X2 AND2X2_6350 ( .A(u5__abc_54027_n1388), .B(u5__abc_54027_n1385), .Y(u5__abc_54027_n1389) );
  AND2X2 AND2X2_6351 ( .A(u5__abc_54027_n1389), .B(u5__abc_54027_n1382), .Y(u5__abc_54027_n1390) );
  AND2X2 AND2X2_6352 ( .A(u5__abc_54027_n375), .B(mc_ack_r), .Y(u5__abc_54027_n1391_1) );
  AND2X2 AND2X2_6353 ( .A(u5__abc_54027_n371), .B(u5__abc_54027_n1383_1), .Y(u5__abc_54027_n1392) );
  AND2X2 AND2X2_6354 ( .A(u5__abc_54027_n826), .B(u5__abc_54027_n1111), .Y(u5__abc_54027_n1395) );
  AND2X2 AND2X2_6355 ( .A(u5__abc_54027_n1394), .B(u5__abc_54027_n1395), .Y(u5__abc_54027_n1396_1) );
  AND2X2 AND2X2_6356 ( .A(u5__abc_54027_n1396_1), .B(u5__abc_54027_n1390), .Y(u5__abc_54027_n1397) );
  AND2X2 AND2X2_6357 ( .A(u5__abc_54027_n1397), .B(u5__abc_54027_n1380_1), .Y(u5__abc_54027_n1398) );
  AND2X2 AND2X2_6358 ( .A(u5__abc_54027_n1363), .B(u5__abc_54027_n1398), .Y(u5__abc_54027_n1399) );
  AND2X2 AND2X2_6359 ( .A(u5__abc_54027_n1402), .B(u5_tmr_done), .Y(u5__abc_54027_n1403) );
  AND2X2 AND2X2_636 ( .A(u0__abc_49347_n1175_bF_buf5), .B(u0__abc_49347_n2749), .Y(u0__abc_49347_n2750) );
  AND2X2 AND2X2_6360 ( .A(u5__abc_54027_n1400), .B(u5__abc_54027_n1404), .Y(u5__abc_54027_n1405) );
  AND2X2 AND2X2_6361 ( .A(u5__abc_54027_n598), .B(u5__abc_54027_n519), .Y(u5__abc_54027_n1406) );
  AND2X2 AND2X2_6362 ( .A(u5__abc_54027_n615), .B(u5__abc_54027_n1406), .Y(u5__abc_54027_n1407_1) );
  AND2X2 AND2X2_6363 ( .A(u5__abc_54027_n425), .B(u5__abc_54027_n1312_1), .Y(u5__abc_54027_n1409) );
  AND2X2 AND2X2_6364 ( .A(u5__abc_54027_n1408), .B(u5__abc_54027_n1410), .Y(u5__abc_54027_n1411) );
  AND2X2 AND2X2_6365 ( .A(u5__abc_54027_n1405), .B(u5__abc_54027_n1411), .Y(u5__abc_54027_n1412_1) );
  AND2X2 AND2X2_6366 ( .A(u5__abc_54027_n598), .B(u5_kro), .Y(u5__abc_54027_n1415) );
  AND2X2 AND2X2_6367 ( .A(u5__abc_54027_n615), .B(u5__abc_54027_n1415), .Y(u5__abc_54027_n1416) );
  AND2X2 AND2X2_6368 ( .A(u5__abc_54027_n1414), .B(u5__abc_54027_n1417), .Y(u5__abc_54027_n1418) );
  AND2X2 AND2X2_6369 ( .A(u5__abc_54027_n1419), .B(u5__abc_54027_n1412_1), .Y(u5__abc_54027_n1420) );
  AND2X2 AND2X2_637 ( .A(u0__abc_49347_n2747), .B(u0__abc_49347_n2750), .Y(u0__abc_49347_n2751) );
  AND2X2 AND2X2_6370 ( .A(u5__abc_54027_n1421), .B(u5_wb_wait), .Y(u5__abc_54027_n1422) );
  AND2X2 AND2X2_6371 ( .A(u5__abc_54027_n505_1), .B(u5__abc_54027_n591), .Y(u5__abc_54027_n1427) );
  AND2X2 AND2X2_6372 ( .A(u5__abc_54027_n1429), .B(u5__abc_54027_n1423), .Y(u5__abc_54027_n1430) );
  AND2X2 AND2X2_6373 ( .A(u5__abc_54027_n1430), .B(u5__abc_54027_n1420), .Y(u5__abc_54027_n1431) );
  AND2X2 AND2X2_6374 ( .A(u5__abc_54027_n1399), .B(u5__abc_54027_n1431), .Y(u5__abc_54027_n1432) );
  AND2X2 AND2X2_6375 ( .A(u5__abc_54027_n1299), .B(u5__abc_54027_n1433), .Y(u5__abc_54027_n1434) );
  AND2X2 AND2X2_6376 ( .A(u5__abc_54027_n904), .B(u5__abc_54027_n1436), .Y(u5__abc_54027_n1437) );
  AND2X2 AND2X2_6377 ( .A(u5__abc_54027_n447_1), .B(u5__abc_54027_n1312_1), .Y(u5__abc_54027_n1438_1) );
  AND2X2 AND2X2_6378 ( .A(u5__abc_54027_n510), .B(u5__abc_54027_n507), .Y(u5__abc_54027_n1439) );
  AND2X2 AND2X2_6379 ( .A(u5__abc_54027_n1356), .B(u5__abc_54027_n1439), .Y(u5__abc_54027_n1440) );
  AND2X2 AND2X2_638 ( .A(u0__abc_49347_n1176_1_bF_buf5), .B(tms_1_), .Y(u0__abc_49347_n2753) );
  AND2X2 AND2X2_6380 ( .A(u5__abc_54027_n873), .B(mc_br_r), .Y(u5__abc_54027_n1443) );
  AND2X2 AND2X2_6381 ( .A(u5__abc_54027_n359), .B(u5__abc_54027_n290_1), .Y(u5__abc_54027_n1444) );
  AND2X2 AND2X2_6382 ( .A(u5__abc_54027_n1442), .B(u5__abc_54027_n1446), .Y(u5__abc_54027_n1447) );
  AND2X2 AND2X2_6383 ( .A(u5__abc_54027_n344_1), .B(u5__abc_54027_n1383_1), .Y(u5__abc_54027_n1448_1) );
  AND2X2 AND2X2_6384 ( .A(u5__abc_54027_n347), .B(u5_cmd_asserted_bF_buf3), .Y(u5__abc_54027_n1449) );
  AND2X2 AND2X2_6385 ( .A(u5__abc_54027_n377), .B(u5__abc_54027_n1299), .Y(u5__abc_54027_n1452) );
  AND2X2 AND2X2_6386 ( .A(u5__abc_54027_n1451), .B(u5__abc_54027_n1454_1), .Y(u5__abc_54027_n1455_1) );
  AND2X2 AND2X2_6387 ( .A(u5__abc_54027_n374), .B(u5__abc_54027_n290_1), .Y(u5__abc_54027_n1456) );
  AND2X2 AND2X2_6388 ( .A(u5__abc_54027_n1456), .B(u5_tmr_done), .Y(u5__abc_54027_n1457) );
  AND2X2 AND2X2_6389 ( .A(u5__abc_54027_n354), .B(u5__abc_54027_n1312_1), .Y(u5__abc_54027_n1458) );
  AND2X2 AND2X2_639 ( .A(u0_tms5_1_), .B(u0_cs5_bF_buf3), .Y(u0__abc_49347_n2754) );
  AND2X2 AND2X2_6390 ( .A(u5__abc_54027_n376), .B(u5__abc_54027_n436), .Y(u5__abc_54027_n1461) );
  AND2X2 AND2X2_6391 ( .A(u5__abc_54027_n1460), .B(u5__abc_54027_n1463), .Y(u5__abc_54027_n1464) );
  AND2X2 AND2X2_6392 ( .A(u5__abc_54027_n1464), .B(u5__abc_54027_n1455_1), .Y(u5__abc_54027_n1465) );
  AND2X2 AND2X2_6393 ( .A(u5__abc_54027_n1465), .B(u5__abc_54027_n1447), .Y(u5__abc_54027_n1466) );
  AND2X2 AND2X2_6394 ( .A(u5_wb_cycle), .B(u5_wb_wait), .Y(u5__abc_54027_n1469) );
  AND2X2 AND2X2_6395 ( .A(u5__abc_54027_n1471), .B(u5__abc_54027_n1468), .Y(u5__abc_54027_n1472) );
  AND2X2 AND2X2_6396 ( .A(u5__abc_54027_n656), .B(u5__abc_54027_n312_1), .Y(u5__abc_54027_n1474) );
  AND2X2 AND2X2_6397 ( .A(u5__abc_54027_n1473), .B(u5__abc_54027_n1474), .Y(u5__abc_54027_n1475) );
  AND2X2 AND2X2_6398 ( .A(u5__abc_54027_n290_1), .B(u5__abc_54027_n656), .Y(u5__abc_54027_n1478) );
  AND2X2 AND2X2_6399 ( .A(u5__abc_54027_n1478), .B(u5__abc_54027_n1383_1), .Y(u5__abc_54027_n1479) );
  AND2X2 AND2X2_64 ( .A(u0__abc_49347_n1113_1), .B(spec_req_cs_1_bF_buf4), .Y(u0__abc_49347_n1114) );
  AND2X2 AND2X2_640 ( .A(u0__abc_49347_n2756), .B(u0__abc_49347_n2730_bF_buf4), .Y(u0__abc_49347_n2757) );
  AND2X2 AND2X2_6400 ( .A(u5__abc_54027_n445), .B(u5_cmd_asserted_bF_buf2), .Y(u5__abc_54027_n1480) );
  AND2X2 AND2X2_6401 ( .A(u5__abc_54027_n297), .B(u5__abc_54027_n1383_1), .Y(u5__abc_54027_n1484) );
  AND2X2 AND2X2_6402 ( .A(u5__abc_54027_n1483), .B(u5__abc_54027_n1485), .Y(u5__abc_54027_n1486) );
  AND2X2 AND2X2_6403 ( .A(u5__abc_54027_n1482), .B(u5__abc_54027_n1486), .Y(u5__abc_54027_n1487) );
  AND2X2 AND2X2_6404 ( .A(u5__abc_54027_n1477), .B(u5__abc_54027_n1487), .Y(u5__abc_54027_n1488) );
  AND2X2 AND2X2_6405 ( .A(u5__abc_54027_n278), .B(u5__abc_54027_n300_1), .Y(u5__abc_54027_n1490) );
  AND2X2 AND2X2_6406 ( .A(u5__abc_54027_n1491_1), .B(u5__abc_54027_n1489), .Y(u5__abc_54027_n1492) );
  AND2X2 AND2X2_6407 ( .A(u5__abc_54027_n1496), .B(u5__abc_54027_n1493), .Y(u5__abc_54027_n1497) );
  AND2X2 AND2X2_6408 ( .A(u5__abc_54027_n1488), .B(u5__abc_54027_n1497), .Y(u5__abc_54027_n1498) );
  AND2X2 AND2X2_6409 ( .A(u5__abc_54027_n1498), .B(u5__abc_54027_n1466), .Y(u5__abc_54027_n1499) );
  AND2X2 AND2X2_641 ( .A(u0__abc_49347_n2757), .B(u0__abc_49347_n2755), .Y(u0__abc_49347_n2758) );
  AND2X2 AND2X2_6410 ( .A(u5__abc_54027_n1499), .B(u5__abc_54027_n1437), .Y(u5__abc_54027_n1500) );
  AND2X2 AND2X2_6411 ( .A(u5__abc_54027_n511), .B(u5_wb_wait), .Y(u5__abc_54027_n1501) );
  AND2X2 AND2X2_6412 ( .A(u5__abc_54027_n351_bF_buf1), .B(u5__abc_54027_n1501), .Y(u5__abc_54027_n1502) );
  AND2X2 AND2X2_6413 ( .A(u5__abc_54027_n1353), .B(u5__abc_54027_n512_1), .Y(u5__abc_54027_n1503) );
  AND2X2 AND2X2_6414 ( .A(u5__abc_54027_n1503), .B(u5__abc_54027_n596), .Y(u5__abc_54027_n1504) );
  AND2X2 AND2X2_6415 ( .A(u5__abc_54027_n1504), .B(u5__abc_54027_n1502), .Y(u5__abc_54027_n1505) );
  AND2X2 AND2X2_6416 ( .A(u5__abc_54027_n1505), .B(u5__abc_54027_n505_1), .Y(u5__abc_54027_n1506) );
  AND2X2 AND2X2_6417 ( .A(u5_cmd_asserted2), .B(mc_br_r), .Y(u5__abc_54027_n1507) );
  AND2X2 AND2X2_6418 ( .A(u5__abc_54027_n1356), .B(u5__abc_54027_n1507), .Y(u5__abc_54027_n1508) );
  AND2X2 AND2X2_6419 ( .A(u5__abc_54027_n1354), .B(u5__abc_54027_n1508), .Y(u5__abc_54027_n1509) );
  AND2X2 AND2X2_642 ( .A(u0__abc_49347_n2759), .B(u0__abc_49347_n2726_bF_buf4), .Y(u0__abc_49347_n2760) );
  AND2X2 AND2X2_6420 ( .A(u5__abc_54027_n587), .B(u5__abc_54027_n1358), .Y(u5__abc_54027_n1510) );
  AND2X2 AND2X2_6421 ( .A(u5__abc_54027_n1510), .B(u5__abc_54027_n1352), .Y(u5__abc_54027_n1511) );
  AND2X2 AND2X2_6422 ( .A(u5__abc_54027_n595), .B(u5__abc_54027_n1515), .Y(u5__abc_54027_n1516) );
  AND2X2 AND2X2_6423 ( .A(u5__abc_54027_n588), .B(u5__abc_54027_n1516), .Y(u5__abc_54027_n1517) );
  AND2X2 AND2X2_6424 ( .A(u5__abc_54027_n359), .B(u5__abc_54027_n277), .Y(u5__abc_54027_n1518) );
  AND2X2 AND2X2_6425 ( .A(u5__abc_54027_n1518), .B(u5_tmr_done), .Y(u5__abc_54027_n1519) );
  AND2X2 AND2X2_6426 ( .A(u5__abc_54027_n278), .B(u5__abc_54027_n293), .Y(u5__abc_54027_n1520) );
  AND2X2 AND2X2_6427 ( .A(u5__abc_54027_n1472), .B(u5__abc_54027_n1474), .Y(u5__abc_54027_n1522) );
  AND2X2 AND2X2_6428 ( .A(u5__abc_54027_n452_1), .B(u5_kro), .Y(u5__abc_54027_n1523) );
  AND2X2 AND2X2_6429 ( .A(u5__abc_54027_n1523), .B(u5_tmr_done), .Y(u5__abc_54027_n1524) );
  AND2X2 AND2X2_643 ( .A(u0_tms4_1_), .B(u0_cs4_bF_buf3), .Y(u0__abc_49347_n2761) );
  AND2X2 AND2X2_6430 ( .A(u5__abc_54027_n1530), .B(u5__abc_54027_n1312_1), .Y(u5__abc_54027_n1531) );
  AND2X2 AND2X2_6431 ( .A(u5__abc_54027_n660), .B(u5__abc_54027_n1531), .Y(u5__abc_54027_n1532) );
  AND2X2 AND2X2_6432 ( .A(u5__abc_54027_n415), .B(u5__abc_54027_n290_1), .Y(u5__abc_54027_n1535) );
  AND2X2 AND2X2_6433 ( .A(u5__abc_54027_n670), .B(u5__abc_54027_n1536), .Y(u5__abc_54027_n1537_1) );
  AND2X2 AND2X2_6434 ( .A(u5__abc_54027_n1534), .B(u5__abc_54027_n1538), .Y(u5__abc_54027_n1539) );
  AND2X2 AND2X2_6435 ( .A(u5__abc_54027_n1529), .B(u5__abc_54027_n1539), .Y(u5__abc_54027_n1540_1) );
  AND2X2 AND2X2_6436 ( .A(u5__abc_54027_n1500), .B(u5__abc_54027_n1540_1), .Y(u5__abc_54027_n1541_1) );
  AND2X2 AND2X2_6437 ( .A(u5__abc_54027_n1541_1), .B(u5__abc_54027_n1432), .Y(u5__abc_54027_n1542_1) );
  AND2X2 AND2X2_6438 ( .A(u5__abc_54027_n1542_1), .B(u5__abc_54027_n1342), .Y(u5__abc_54027_n1543) );
  AND2X2 AND2X2_6439 ( .A(u5__abc_54027_n1543), .B(u5__abc_54027_n1334), .Y(u5__abc_54027_n1544_1) );
  AND2X2 AND2X2_644 ( .A(u0__abc_49347_n2762), .B(u0__abc_49347_n2725_bF_buf4), .Y(u0__abc_49347_n2763) );
  AND2X2 AND2X2_6440 ( .A(u5__abc_54027_n1544_1), .B(u5__abc_54027_n1325), .Y(u5__abc_54027_n1545) );
  AND2X2 AND2X2_6441 ( .A(u5__abc_54027_n678), .B(u5__abc_54027_n1338), .Y(u5__abc_54027_n1548) );
  AND2X2 AND2X2_6442 ( .A(u5__abc_54027_n374), .B(u5__abc_54027_n312_1), .Y(u5__abc_54027_n1549) );
  AND2X2 AND2X2_6443 ( .A(u5__abc_54027_n641), .B(u5__abc_54027_n501), .Y(u5__abc_54027_n1550) );
  AND2X2 AND2X2_6444 ( .A(u5__abc_54027_n519), .B(u5__abc_54027_n1551_1), .Y(u5__abc_54027_n1552_1) );
  AND2X2 AND2X2_6445 ( .A(u5__abc_54027_n631), .B(u5__abc_54027_n1553), .Y(u5__abc_54027_n1554_1) );
  AND2X2 AND2X2_6446 ( .A(u5__abc_54027_n1555_1), .B(u5__abc_54027_n1549), .Y(u5__abc_54027_n1556) );
  AND2X2 AND2X2_6447 ( .A(u5__abc_54027_n1560), .B(u5__abc_54027_n477), .Y(u5__abc_54027_n1561_1) );
  AND2X2 AND2X2_6448 ( .A(u5__abc_54027_n505_1), .B(u5__abc_54027_n477), .Y(u5__abc_54027_n1563) );
  AND2X2 AND2X2_6449 ( .A(u5_kro), .B(bank_open), .Y(u5__abc_54027_n1564) );
  AND2X2 AND2X2_645 ( .A(u0_tms3_1_), .B(u0_cs3_bF_buf3), .Y(u0__abc_49347_n2764) );
  AND2X2 AND2X2_6450 ( .A(u5__abc_54027_n595), .B(u5__abc_54027_n1564), .Y(u5__abc_54027_n1565) );
  AND2X2 AND2X2_6451 ( .A(u5__abc_54027_n587), .B(u5__abc_54027_n1565), .Y(u5__abc_54027_n1566) );
  AND2X2 AND2X2_6452 ( .A(u5__abc_54027_n1566), .B(row_same), .Y(u5__abc_54027_n1567) );
  AND2X2 AND2X2_6453 ( .A(u5__abc_54027_n1567), .B(u5__abc_54027_n1563), .Y(u5__abc_54027_n1568) );
  AND2X2 AND2X2_6454 ( .A(u5__abc_54027_n1569), .B(u5__abc_54027_n1562_1), .Y(u5__abc_54027_n1570) );
  AND2X2 AND2X2_6455 ( .A(u5__abc_54027_n1570), .B(u5__abc_54027_n1437), .Y(u5__abc_54027_n1571_1) );
  AND2X2 AND2X2_6456 ( .A(u5__abc_54027_n347), .B(u5__abc_54027_n1312_1), .Y(u5__abc_54027_n1572_1) );
  AND2X2 AND2X2_6457 ( .A(u5__abc_54027_n1566), .B(u5__abc_54027_n1573_1), .Y(u5__abc_54027_n1574_1) );
  AND2X2 AND2X2_6458 ( .A(u5__abc_54027_n1574_1), .B(u5__abc_54027_n1563), .Y(u5__abc_54027_n1575_1) );
  AND2X2 AND2X2_6459 ( .A(u5__abc_54027_n1478), .B(u5_tmr_done), .Y(u5__abc_54027_n1579) );
  AND2X2 AND2X2_646 ( .A(u0__abc_49347_n2765), .B(u0__abc_49347_n2724_bF_buf4), .Y(u0__abc_49347_n2766) );
  AND2X2 AND2X2_6460 ( .A(u5__abc_54027_n1532), .B(u5__abc_54027_n460), .Y(u5__abc_54027_n1580) );
  AND2X2 AND2X2_6461 ( .A(u5__abc_54027_n1578), .B(u5__abc_54027_n1582), .Y(u5__abc_54027_n1583) );
  AND2X2 AND2X2_6462 ( .A(u5__abc_54027_n1583), .B(u5__abc_54027_n1571_1), .Y(u5__abc_54027_n1584) );
  AND2X2 AND2X2_6463 ( .A(u5__abc_54027_n375), .B(u5__abc_54027_n1434), .Y(u5__abc_54027_n1585) );
  AND2X2 AND2X2_6464 ( .A(u5__abc_54027_n849), .B(u5__abc_54027_n1586), .Y(u5__abc_54027_n1587) );
  AND2X2 AND2X2_6465 ( .A(u5__abc_54027_n477), .B(u3_wb_read_go), .Y(u5__abc_54027_n1588) );
  AND2X2 AND2X2_6466 ( .A(u5__abc_54027_n1490), .B(u5__abc_54027_n1588), .Y(u5__abc_54027_n1589) );
  AND2X2 AND2X2_6467 ( .A(u5__abc_54027_n369), .B(u5__abc_54027_n1312_1), .Y(u5__abc_54027_n1590) );
  AND2X2 AND2X2_6468 ( .A(u5__abc_54027_n587), .B(u5__abc_54027_n598), .Y(u5__abc_54027_n1592) );
  AND2X2 AND2X2_6469 ( .A(u5__abc_54027_n596), .B(u5__abc_54027_n666_1), .Y(u5__abc_54027_n1593) );
  AND2X2 AND2X2_647 ( .A(u0_tms2_1_), .B(u0_cs2_bF_buf3), .Y(u0__abc_49347_n2767) );
  AND2X2 AND2X2_6470 ( .A(u5__abc_54027_n505_1), .B(u5__abc_54027_n1593), .Y(u5__abc_54027_n1594) );
  AND2X2 AND2X2_6471 ( .A(u5__abc_54027_n1592), .B(u5__abc_54027_n1594), .Y(u5__abc_54027_n1595) );
  AND2X2 AND2X2_6472 ( .A(u5__abc_54027_n1430), .B(u5__abc_54027_n1597), .Y(u5__abc_54027_n1598) );
  AND2X2 AND2X2_6473 ( .A(u5__abc_54027_n1598), .B(u5__abc_54027_n1587), .Y(u5__abc_54027_n1599) );
  AND2X2 AND2X2_6474 ( .A(u5__abc_54027_n1592), .B(u5__abc_54027_n1427), .Y(u5__abc_54027_n1600) );
  AND2X2 AND2X2_6475 ( .A(u5__abc_54027_n301_1), .B(u5__abc_54027_n1312_1), .Y(u5__abc_54027_n1602) );
  AND2X2 AND2X2_6476 ( .A(u5__abc_54027_n294), .B(u5__abc_54027_n1604), .Y(u5__abc_54027_n1605) );
  AND2X2 AND2X2_6477 ( .A(u5__abc_54027_n1606), .B(u5__abc_54027_n298_1), .Y(u5__abc_54027_n1607) );
  AND2X2 AND2X2_6478 ( .A(u5__abc_54027_n1608), .B(u5__abc_54027_n1603), .Y(u5__abc_54027_n1609) );
  AND2X2 AND2X2_6479 ( .A(u5__abc_54027_n1488), .B(u5__abc_54027_n1609), .Y(u5__abc_54027_n1610) );
  AND2X2 AND2X2_648 ( .A(u0__abc_49347_n2768), .B(u0__abc_49347_n2723_bF_buf4), .Y(u0__abc_49347_n2769) );
  AND2X2 AND2X2_6480 ( .A(u5__abc_54027_n1610), .B(u5__abc_54027_n1601), .Y(u5__abc_54027_n1611) );
  AND2X2 AND2X2_6481 ( .A(u5__abc_54027_n1375), .B(u5__abc_54027_n1368), .Y(u5__abc_54027_n1612) );
  AND2X2 AND2X2_6482 ( .A(u5__abc_54027_n1456), .B(u5__abc_54027_n1383_1), .Y(u5__abc_54027_n1613) );
  AND2X2 AND2X2_6483 ( .A(u5__abc_54027_n447_1), .B(u5_cmd_asserted_bF_buf1), .Y(u5__abc_54027_n1614) );
  AND2X2 AND2X2_6484 ( .A(u5__abc_54027_n1616), .B(u5__abc_54027_n1405), .Y(u5__abc_54027_n1617) );
  AND2X2 AND2X2_6485 ( .A(u5__abc_54027_n1617), .B(u5__abc_54027_n1612), .Y(u5__abc_54027_n1618) );
  AND2X2 AND2X2_6486 ( .A(u5__abc_54027_n1619), .B(u5__abc_54027_n1620), .Y(u5__abc_54027_n1621) );
  AND2X2 AND2X2_6487 ( .A(u5__abc_54027_n579_1), .B(u5__abc_54027_n396), .Y(u5__abc_54027_n1623) );
  AND2X2 AND2X2_6488 ( .A(u5__abc_54027_n1624), .B(u5__abc_54027_n1382), .Y(u5__abc_54027_n1625) );
  AND2X2 AND2X2_6489 ( .A(u5__abc_54027_n1623), .B(u5__abc_54027_n1625), .Y(u5__abc_54027_n1626) );
  AND2X2 AND2X2_649 ( .A(u0_tms1_1_), .B(u0_cs1_bF_buf3), .Y(u0__abc_49347_n2770) );
  AND2X2 AND2X2_6490 ( .A(u5__abc_54027_n1622), .B(u5__abc_54027_n1626), .Y(u5__abc_54027_n1627) );
  AND2X2 AND2X2_6491 ( .A(u5__abc_54027_n1627), .B(u5__abc_54027_n1618), .Y(u5__abc_54027_n1628) );
  AND2X2 AND2X2_6492 ( .A(u5__abc_54027_n382), .B(u5__abc_54027_n1299), .Y(u5__abc_54027_n1629) );
  AND2X2 AND2X2_6493 ( .A(u5__abc_54027_n1632), .B(u5__abc_54027_n433_1), .Y(u5__abc_54027_n1633) );
  AND2X2 AND2X2_6494 ( .A(u5__abc_54027_n1535), .B(u5__abc_54027_n1383_1), .Y(u5__abc_54027_n1634) );
  AND2X2 AND2X2_6495 ( .A(u5__abc_54027_n1635), .B(u5__abc_54027_n868_1), .Y(u5__abc_54027_n1636) );
  AND2X2 AND2X2_6496 ( .A(u5__abc_54027_n1633), .B(u5__abc_54027_n1636), .Y(u5__abc_54027_n1637) );
  AND2X2 AND2X2_6497 ( .A(u5__abc_54027_n1637), .B(u5__abc_54027_n1631), .Y(u5__abc_54027_n1638) );
  AND2X2 AND2X2_6498 ( .A(u5__abc_54027_n1447), .B(u5__abc_54027_n1638), .Y(u5__abc_54027_n1639) );
  AND2X2 AND2X2_6499 ( .A(u5__abc_54027_n1628), .B(u5__abc_54027_n1639), .Y(u5__abc_54027_n1640) );
  AND2X2 AND2X2_65 ( .A(u0__abc_49347_n1113_1), .B(spec_req_cs_2_bF_buf4), .Y(u0__abc_49347_n1116_1) );
  AND2X2 AND2X2_650 ( .A(u0__abc_49347_n1175_bF_buf4), .B(u0__abc_49347_n2773), .Y(u0__abc_49347_n2774) );
  AND2X2 AND2X2_6500 ( .A(u5__abc_54027_n1611), .B(u5__abc_54027_n1640), .Y(u5__abc_54027_n1641) );
  AND2X2 AND2X2_6501 ( .A(u5__abc_54027_n1641), .B(u5__abc_54027_n1599), .Y(u5__abc_54027_n1642) );
  AND2X2 AND2X2_6502 ( .A(u5__abc_54027_n1642), .B(u5__abc_54027_n1584), .Y(u5__abc_54027_n1643) );
  AND2X2 AND2X2_6503 ( .A(u5__abc_54027_n678), .B(u5_wb_cycle), .Y(u5__abc_54027_n1647) );
  AND2X2 AND2X2_6504 ( .A(u5__abc_54027_n1321), .B(u5__abc_54027_n1551_1), .Y(u5__abc_54027_n1650) );
  AND2X2 AND2X2_6505 ( .A(u5__abc_54027_n1649), .B(u5__abc_54027_n1650), .Y(u5__abc_54027_n1651) );
  AND2X2 AND2X2_6506 ( .A(u5__abc_54027_n1648), .B(u5__abc_54027_n1651), .Y(u5__abc_54027_n1652) );
  AND2X2 AND2X2_6507 ( .A(u5__abc_54027_n678), .B(u5__abc_54027_n1551_1), .Y(u5__abc_54027_n1653) );
  AND2X2 AND2X2_6508 ( .A(u5__abc_54027_n1653), .B(u5__abc_54027_n1319), .Y(u5__abc_54027_n1654) );
  AND2X2 AND2X2_6509 ( .A(u5__abc_54027_n429_1), .B(u5_cmd_asserted_bF_buf0), .Y(u5__abc_54027_n1655) );
  AND2X2 AND2X2_651 ( .A(u0__abc_49347_n2772), .B(u0__abc_49347_n2774), .Y(u0__abc_49347_n2775) );
  AND2X2 AND2X2_6510 ( .A(u5__abc_54027_n574), .B(u5__abc_54027_n1312_1), .Y(u5__abc_54027_n1656) );
  AND2X2 AND2X2_6511 ( .A(u5__abc_54027_n452_1), .B(u5__abc_54027_n1383_1), .Y(u5__abc_54027_n1658) );
  AND2X2 AND2X2_6512 ( .A(u5__abc_54027_n1659), .B(u5__abc_54027_n1549), .Y(u5__abc_54027_n1660) );
  AND2X2 AND2X2_6513 ( .A(u5__abc_54027_n1660), .B(u5__abc_54027_n1552_1), .Y(u5__abc_54027_n1661) );
  AND2X2 AND2X2_6514 ( .A(u5__abc_54027_n1663), .B(u5__abc_54027_n1657), .Y(u5__abc_54027_n1664) );
  AND2X2 AND2X2_6515 ( .A(u5__abc_54027_n1325), .B(u5__abc_54027_n1668), .Y(u5__abc_54027_n1669) );
  AND2X2 AND2X2_6516 ( .A(u5__abc_54027_n483), .B(u5__abc_54027_n1317), .Y(u5__abc_54027_n1673) );
  AND2X2 AND2X2_6517 ( .A(u5__abc_54027_n1672), .B(u5__abc_54027_n1673), .Y(u5__abc_54027_n1674) );
  AND2X2 AND2X2_6518 ( .A(u5__abc_54027_n1674), .B(u5__abc_54027_n1326), .Y(u5__abc_54027_n1675) );
  AND2X2 AND2X2_6519 ( .A(u5__abc_54027_n467), .B(u3_wb_read_go), .Y(u5__abc_54027_n1676) );
  AND2X2 AND2X2_652 ( .A(u0__abc_49347_n1176_1_bF_buf4), .B(tms_2_), .Y(u0__abc_49347_n2777) );
  AND2X2 AND2X2_6520 ( .A(u5__abc_54027_n1679), .B(u5__abc_54027_n1675), .Y(u5__abc_54027_n1680) );
  AND2X2 AND2X2_6521 ( .A(u5__abc_54027_n680), .B(u1_wb_write_go), .Y(u5__abc_54027_n1682) );
  AND2X2 AND2X2_6522 ( .A(u5__abc_54027_n1648), .B(u5__abc_54027_n1682), .Y(u5__abc_54027_n1683) );
  AND2X2 AND2X2_6523 ( .A(u5__abc_54027_n1684), .B(u5__abc_54027_n1685), .Y(u5__abc_54027_n1686) );
  AND2X2 AND2X2_6524 ( .A(u5__abc_54027_n1681), .B(u5__abc_54027_n1686), .Y(u5__abc_54027_n1687) );
  AND2X2 AND2X2_6525 ( .A(u5__abc_54027_n1327), .B(u5__abc_54027_n319), .Y(u5__abc_54027_n1690) );
  AND2X2 AND2X2_6526 ( .A(u5__abc_54027_n1295), .B(u5_tmr2_done), .Y(u5__abc_54027_n1691) );
  AND2X2 AND2X2_6527 ( .A(u5__abc_54027_n1477), .B(u5__abc_54027_n1451), .Y(u5__abc_54027_n1694) );
  AND2X2 AND2X2_6528 ( .A(u5__abc_54027_n1578), .B(u5__abc_54027_n1694), .Y(u5__abc_54027_n1695) );
  AND2X2 AND2X2_6529 ( .A(u5__abc_54027_n662), .B(u5__abc_54027_n1367), .Y(u5__abc_54027_n1696) );
  AND2X2 AND2X2_653 ( .A(u0_tms5_2_), .B(u0_cs5_bF_buf2), .Y(u0__abc_49347_n2778) );
  AND2X2 AND2X2_6530 ( .A(u5__abc_54027_n1394), .B(u5__abc_54027_n1696), .Y(u5__abc_54027_n1697) );
  AND2X2 AND2X2_6531 ( .A(u5__abc_54027_n1697), .B(u5__abc_54027_n1423), .Y(u5__abc_54027_n1698) );
  AND2X2 AND2X2_6532 ( .A(u5__abc_54027_n1460), .B(u5__abc_54027_n1616), .Y(u5__abc_54027_n1699) );
  AND2X2 AND2X2_6533 ( .A(u5__abc_54027_n1699), .B(u5__abc_54027_n1442), .Y(u5__abc_54027_n1700) );
  AND2X2 AND2X2_6534 ( .A(u5__abc_54027_n1700), .B(u5__abc_54027_n1698), .Y(u5__abc_54027_n1701) );
  AND2X2 AND2X2_6535 ( .A(u5__abc_54027_n1351), .B(u5__abc_54027_n1631), .Y(u5__abc_54027_n1702) );
  AND2X2 AND2X2_6536 ( .A(u5__abc_54027_n390_1), .B(u5__abc_54027_n1299), .Y(u5__abc_54027_n1703) );
  AND2X2 AND2X2_6537 ( .A(u5__abc_54027_n1706), .B(u5__abc_54027_n1705), .Y(u5__abc_54027_n1707) );
  AND2X2 AND2X2_6538 ( .A(u5__abc_54027_n290_1), .B(u5__abc_54027_n343), .Y(u5__abc_54027_n1708) );
  AND2X2 AND2X2_6539 ( .A(u5__abc_54027_n291), .B(u5__abc_54027_n1312_1), .Y(u5__abc_54027_n1709) );
  AND2X2 AND2X2_654 ( .A(u0__abc_49347_n2780), .B(u0__abc_49347_n2730_bF_buf3), .Y(u0__abc_49347_n2781) );
  AND2X2 AND2X2_6540 ( .A(u5__abc_54027_n869_1), .B(u5__abc_54027_n1712), .Y(u5__abc_54027_n1713) );
  AND2X2 AND2X2_6541 ( .A(u5__abc_54027_n354), .B(u5_cmd_asserted_bF_buf3), .Y(u5__abc_54027_n1714) );
  AND2X2 AND2X2_6542 ( .A(u5__abc_54027_n1716), .B(u5__abc_54027_n1711), .Y(u5__abc_54027_n1717) );
  AND2X2 AND2X2_6543 ( .A(u5__abc_54027_n1717), .B(u5__abc_54027_n1707), .Y(u5__abc_54027_n1718) );
  AND2X2 AND2X2_6544 ( .A(u5__abc_54027_n1718), .B(u5__abc_54027_n1702), .Y(u5__abc_54027_n1719) );
  AND2X2 AND2X2_6545 ( .A(u5__abc_54027_n1701), .B(u5__abc_54027_n1719), .Y(u5__abc_54027_n1720) );
  AND2X2 AND2X2_6546 ( .A(u5__abc_54027_n561), .B(u5_tmr_done), .Y(u5__abc_54027_n1721) );
  AND2X2 AND2X2_6547 ( .A(u5__abc_54027_n344_1), .B(u5__abc_54027_n1721), .Y(u5__abc_54027_n1722) );
  AND2X2 AND2X2_6548 ( .A(u5__abc_54027_n362), .B(u5__abc_54027_n1312_1), .Y(u5__abc_54027_n1723) );
  AND2X2 AND2X2_6549 ( .A(u5__abc_54027_n587), .B(u5__abc_54027_n595), .Y(u5__abc_54027_n1725) );
  AND2X2 AND2X2_655 ( .A(u0__abc_49347_n2781), .B(u0__abc_49347_n2779), .Y(u0__abc_49347_n2782) );
  AND2X2 AND2X2_6550 ( .A(u5__abc_54027_n1563), .B(u5__abc_54027_n1726), .Y(u5__abc_54027_n1727) );
  AND2X2 AND2X2_6551 ( .A(u5__abc_54027_n1727), .B(u5__abc_54027_n1725), .Y(u5__abc_54027_n1728) );
  AND2X2 AND2X2_6552 ( .A(u5__abc_54027_n1454_1), .B(u5__abc_54027_n1446), .Y(u5__abc_54027_n1731) );
  AND2X2 AND2X2_6553 ( .A(u5__abc_54027_n1731), .B(u5__abc_54027_n1601), .Y(u5__abc_54027_n1732) );
  AND2X2 AND2X2_6554 ( .A(u5__abc_54027_n1732), .B(u5__abc_54027_n1587), .Y(u5__abc_54027_n1733) );
  AND2X2 AND2X2_6555 ( .A(u5__abc_54027_n1730), .B(u5__abc_54027_n1733), .Y(u5__abc_54027_n1734) );
  AND2X2 AND2X2_6556 ( .A(u5__abc_54027_n1720), .B(u5__abc_54027_n1734), .Y(u5__abc_54027_n1735) );
  AND2X2 AND2X2_6557 ( .A(u5__abc_54027_n1695), .B(u5__abc_54027_n1735), .Y(u5__abc_54027_n1736) );
  AND2X2 AND2X2_6558 ( .A(u5__abc_54027_n1582), .B(u5__abc_54027_n1388), .Y(u5__abc_54027_n1737) );
  AND2X2 AND2X2_6559 ( .A(u5__abc_54027_n1378_1), .B(u5__abc_54027_n1382), .Y(u5__abc_54027_n1738) );
  AND2X2 AND2X2_656 ( .A(u0__abc_49347_n2783), .B(u0__abc_49347_n2726_bF_buf3), .Y(u0__abc_49347_n2784_1) );
  AND2X2 AND2X2_6560 ( .A(u5__abc_54027_n1738), .B(u5__abc_54027_n1482), .Y(u5__abc_54027_n1739) );
  AND2X2 AND2X2_6561 ( .A(u5__abc_54027_n1597), .B(u5__abc_54027_n1739), .Y(u5__abc_54027_n1740) );
  AND2X2 AND2X2_6562 ( .A(u5__abc_54027_n1737), .B(u5__abc_54027_n1740), .Y(u5__abc_54027_n1741) );
  AND2X2 AND2X2_6563 ( .A(u5__abc_54027_n1736), .B(u5__abc_54027_n1741), .Y(u5__abc_54027_n1742) );
  AND2X2 AND2X2_6564 ( .A(u5__abc_54027_n1570), .B(u5__abc_54027_n1420), .Y(u5__abc_54027_n1747) );
  AND2X2 AND2X2_6565 ( .A(u5__abc_54027_n1747), .B(u5__abc_54027_n1730), .Y(u5__abc_54027_n1748) );
  AND2X2 AND2X2_6566 ( .A(u5__abc_54027_n1695), .B(u5__abc_54027_n1748), .Y(u5__abc_54027_n1749) );
  AND2X2 AND2X2_6567 ( .A(u5__abc_54027_n425), .B(u5_cmd_asserted_bF_buf2), .Y(u5__abc_54027_n1752) );
  AND2X2 AND2X2_6568 ( .A(u5__abc_54027_n1751), .B(u5__abc_54027_n1753), .Y(u5__abc_54027_n1754) );
  AND2X2 AND2X2_6569 ( .A(u5__abc_54027_n1424), .B(u5_cmd_asserted_bF_buf1), .Y(u5__abc_54027_n1756) );
  AND2X2 AND2X2_657 ( .A(u0_tms4_2_), .B(u0_cs4_bF_buf2), .Y(u0__abc_49347_n2785) );
  AND2X2 AND2X2_6570 ( .A(u5__abc_54027_n1757), .B(u5__abc_54027_n1755), .Y(u5__abc_54027_n1758) );
  AND2X2 AND2X2_6571 ( .A(u5__abc_54027_n1759), .B(u5__abc_54027_n398), .Y(u5__abc_54027_n1760) );
  AND2X2 AND2X2_6572 ( .A(u5__abc_54027_n1758), .B(u5__abc_54027_n1760), .Y(u5__abc_54027_n1761) );
  AND2X2 AND2X2_6573 ( .A(u5__abc_54027_n1761), .B(u5__abc_54027_n1754), .Y(u5__abc_54027_n1762) );
  AND2X2 AND2X2_6574 ( .A(u5__abc_54027_n1762), .B(u5__abc_54027_n1622), .Y(u5__abc_54027_n1763) );
  AND2X2 AND2X2_6575 ( .A(u5__abc_54027_n1763), .B(u5__abc_54027_n1497), .Y(u5__abc_54027_n1764) );
  AND2X2 AND2X2_6576 ( .A(u5__abc_54027_n1764), .B(u5__abc_54027_n668), .Y(u5__abc_54027_n1765) );
  AND2X2 AND2X2_6577 ( .A(u5__abc_54027_n1372), .B(u5__abc_54027_n396), .Y(u5__abc_54027_n1766) );
  AND2X2 AND2X2_6578 ( .A(u5__abc_54027_n1766), .B(u5__abc_54027_n1706), .Y(u5__abc_54027_n1767) );
  AND2X2 AND2X2_6579 ( .A(u5__abc_54027_n1767), .B(u5__abc_54027_n1375), .Y(u5__abc_54027_n1768) );
  AND2X2 AND2X2_658 ( .A(u0__abc_49347_n2786), .B(u0__abc_49347_n2725_bF_buf3), .Y(u0__abc_49347_n2787) );
  AND2X2 AND2X2_6580 ( .A(u5__abc_54027_n1768), .B(u5__abc_54027_n1732), .Y(u5__abc_54027_n1769) );
  AND2X2 AND2X2_6581 ( .A(u5__abc_54027_n294), .B(u5__abc_54027_n1771), .Y(u5__abc_54027_n1772) );
  AND2X2 AND2X2_6582 ( .A(u5__abc_54027_n826), .B(u5__abc_54027_n1773), .Y(u5__abc_54027_n1774) );
  AND2X2 AND2X2_6583 ( .A(u5__abc_54027_n1486), .B(u5__abc_54027_n1774), .Y(u5__abc_54027_n1775) );
  AND2X2 AND2X2_6584 ( .A(u5__abc_54027_n1775), .B(u5__abc_54027_n1711), .Y(u5__abc_54027_n1776) );
  AND2X2 AND2X2_6585 ( .A(u5__abc_54027_n1776), .B(u5__abc_54027_n1609), .Y(u5__abc_54027_n1777) );
  AND2X2 AND2X2_6586 ( .A(u5__abc_54027_n1777), .B(u5__abc_54027_n1770), .Y(u5__abc_54027_n1778) );
  AND2X2 AND2X2_6587 ( .A(u5__abc_54027_n1778), .B(u5__abc_54027_n1769), .Y(u5__abc_54027_n1779) );
  AND2X2 AND2X2_6588 ( .A(u5__abc_54027_n1779), .B(u5__abc_54027_n1765), .Y(u5__abc_54027_n1780) );
  AND2X2 AND2X2_6589 ( .A(u5__abc_54027_n1780), .B(u5__abc_54027_n1741), .Y(u5__abc_54027_n1781) );
  AND2X2 AND2X2_659 ( .A(u0_tms3_2_), .B(u0_cs3_bF_buf2), .Y(u0__abc_49347_n2788) );
  AND2X2 AND2X2_6590 ( .A(u5__abc_54027_n1781), .B(u5__abc_54027_n1749), .Y(u5__abc_54027_n1782) );
  AND2X2 AND2X2_6591 ( .A(u5__abc_54027_n1539), .B(u5__abc_54027_n1754), .Y(u5__abc_54027_n1787) );
  AND2X2 AND2X2_6592 ( .A(u5__abc_54027_n1342), .B(u5__abc_54027_n1787), .Y(u5__abc_54027_n1788) );
  AND2X2 AND2X2_6593 ( .A(u5__abc_54027_n1788), .B(u5__abc_54027_n1749), .Y(u5__abc_54027_n1789) );
  AND2X2 AND2X2_6594 ( .A(u5__abc_54027_n1789), .B(u5__abc_54027_n1786), .Y(u5__abc_54027_n1790) );
  AND2X2 AND2X2_6595 ( .A(u5__abc_54027_n1669), .B(u5__abc_54027_n1790), .Y(u5__abc_54027_n1791) );
  AND2X2 AND2X2_6596 ( .A(u5__abc_54027_n1791), .B(u5__abc_54027_n1687), .Y(u5__abc_54027_n1792) );
  AND2X2 AND2X2_6597 ( .A(u5__abc_54027_n1633), .B(u5__abc_54027_n1705), .Y(u5__abc_54027_n1793) );
  AND2X2 AND2X2_6598 ( .A(u5__abc_54027_n1793), .B(u5__abc_54027_n1760), .Y(u5__abc_54027_n1794) );
  AND2X2 AND2X2_6599 ( .A(u5__abc_54027_n580), .B(u5__abc_54027_n406), .Y(u5__abc_54027_n1795) );
  AND2X2 AND2X2_66 ( .A(u0__abc_49347_n1100_1), .B(u0_lmr_req2), .Y(u0__abc_49347_n1118_1) );
  AND2X2 AND2X2_660 ( .A(u0__abc_49347_n2789), .B(u0__abc_49347_n2724_bF_buf3), .Y(u0__abc_49347_n2790) );
  AND2X2 AND2X2_6600 ( .A(u5__abc_54027_n1111), .B(u5__abc_54027_n1367), .Y(u5__abc_54027_n1796) );
  AND2X2 AND2X2_6601 ( .A(u5__abc_54027_n1795), .B(u5__abc_54027_n1796), .Y(u5__abc_54027_n1797) );
  AND2X2 AND2X2_6602 ( .A(u5__abc_54027_n1356), .B(u5__abc_54027_n509), .Y(u5__abc_54027_n1798) );
  AND2X2 AND2X2_6603 ( .A(u5__abc_54027_n1799), .B(u5__abc_54027_n1800), .Y(u5__abc_54027_n1801) );
  AND2X2 AND2X2_6604 ( .A(u5__abc_54027_n1797), .B(u5__abc_54027_n1801), .Y(u5__abc_54027_n1802) );
  AND2X2 AND2X2_6605 ( .A(u5__abc_54027_n1794), .B(u5__abc_54027_n1802), .Y(u5__abc_54027_n1803) );
  AND2X2 AND2X2_6606 ( .A(u5__abc_54027_n1702), .B(u5__abc_54027_n1429), .Y(u5__abc_54027_n1804) );
  AND2X2 AND2X2_6607 ( .A(u5__abc_54027_n1803), .B(u5__abc_54027_n1804), .Y(u5__abc_54027_n1805) );
  AND2X2 AND2X2_6608 ( .A(u5__abc_54027_n1805), .B(u5__abc_54027_n1769), .Y(u5__abc_54027_n1806) );
  AND2X2 AND2X2_6609 ( .A(u5__abc_54027_n1792), .B(u5__abc_54027_n1806), .Y(u5__abc_54027_n1807) );
  AND2X2 AND2X2_661 ( .A(u0_tms2_2_), .B(u0_cs2_bF_buf2), .Y(u0__abc_49347_n2791) );
  AND2X2 AND2X2_6610 ( .A(u5__abc_54027_n283), .B(u5__abc_54027_n290_1), .Y(u5__abc_54027_n1809) );
  AND2X2 AND2X2_6611 ( .A(u5__abc_54027_n1365), .B(u5__abc_54027_n1810), .Y(u5__abc_54027_n1811) );
  AND2X2 AND2X2_6612 ( .A(u5__abc_54027_n1482), .B(u5__abc_54027_n1811), .Y(u5__abc_54027_n1812) );
  AND2X2 AND2X2_6613 ( .A(u5__abc_54027_n1716), .B(u5__abc_54027_n1636), .Y(u5__abc_54027_n1813) );
  AND2X2 AND2X2_6614 ( .A(u5__abc_54027_n1813), .B(u5__abc_54027_n1812), .Y(u5__abc_54027_n1814) );
  AND2X2 AND2X2_6615 ( .A(u5__abc_54027_n1361), .B(u5__abc_54027_n1442), .Y(u5__abc_54027_n1815) );
  AND2X2 AND2X2_6616 ( .A(u5__abc_54027_n1699), .B(u5__abc_54027_n1801), .Y(u5__abc_54027_n1816) );
  AND2X2 AND2X2_6617 ( .A(u5__abc_54027_n1815), .B(u5__abc_54027_n1816), .Y(u5__abc_54027_n1817) );
  AND2X2 AND2X2_6618 ( .A(u5__abc_54027_n1817), .B(u5__abc_54027_n1814), .Y(u5__abc_54027_n1818) );
  AND2X2 AND2X2_6619 ( .A(u5__abc_54027_n1818), .B(u5__abc_54027_n1778), .Y(u5__abc_54027_n1819) );
  AND2X2 AND2X2_662 ( .A(u0__abc_49347_n2792), .B(u0__abc_49347_n2723_bF_buf3), .Y(u0__abc_49347_n2793) );
  AND2X2 AND2X2_6620 ( .A(u5__abc_54027_n1819), .B(u5__abc_54027_n1737), .Y(u5__abc_54027_n1820) );
  AND2X2 AND2X2_6621 ( .A(u5__abc_54027_n1792), .B(u5__abc_54027_n1820), .Y(u5__abc_54027_n1821) );
  AND2X2 AND2X2_6622 ( .A(u5__abc_54027_n1672), .B(u5__abc_54027_n1319), .Y(u5__abc_54027_n1823) );
  AND2X2 AND2X2_6623 ( .A(u5__abc_54027_n1823), .B(u5__abc_54027_n678), .Y(u5__abc_54027_n1824) );
  AND2X2 AND2X2_6624 ( .A(u5__abc_54027_n1649), .B(u5__abc_54027_n1321), .Y(u5__abc_54027_n1825) );
  AND2X2 AND2X2_6625 ( .A(u5__abc_54027_n1648), .B(u5__abc_54027_n1825), .Y(u5__abc_54027_n1826) );
  AND2X2 AND2X2_6626 ( .A(u5__abc_54027_n1827), .B(u5_ap_en), .Y(u5__abc_54027_n1828) );
  AND2X2 AND2X2_6627 ( .A(u5__abc_54027_n420), .B(u5__abc_54027_n1676), .Y(u5__abc_54027_n1830) );
  AND2X2 AND2X2_6628 ( .A(u5__abc_54027_n1829), .B(u5__abc_54027_n1830), .Y(u5__abc_54027_n1831) );
  AND2X2 AND2X2_6629 ( .A(u5__abc_54027_n1831), .B(u5__abc_54027_n1675), .Y(u5__abc_54027_n1832) );
  AND2X2 AND2X2_663 ( .A(u0_tms1_2_), .B(u0_cs1_bF_buf2), .Y(u0__abc_49347_n2794) );
  AND2X2 AND2X2_6630 ( .A(u5__abc_54027_n1647), .B(u5__abc_54027_n680), .Y(u5__abc_54027_n1833) );
  AND2X2 AND2X2_6631 ( .A(u5__abc_54027_n573), .B(u5_cmd_asserted_bF_buf3), .Y(u5__abc_54027_n1834) );
  AND2X2 AND2X2_6632 ( .A(u5__abc_54027_n1553), .B(u5__abc_54027_n630_1), .Y(u5__abc_54027_n1835) );
  AND2X2 AND2X2_6633 ( .A(u5__abc_54027_n1660), .B(u5__abc_54027_n1835), .Y(u5__abc_54027_n1836) );
  AND2X2 AND2X2_6634 ( .A(u5__abc_54027_n873), .B(u5__abc_54027_n1358), .Y(u5__abc_54027_n1838) );
  AND2X2 AND2X2_6635 ( .A(u5__abc_54027_n359), .B(u5__abc_54027_n350), .Y(u5__abc_54027_n1839) );
  AND2X2 AND2X2_6636 ( .A(u5__abc_54027_n1839), .B(u5__abc_54027_n1383_1), .Y(u5__abc_54027_n1840) );
  AND2X2 AND2X2_6637 ( .A(u5__abc_54027_n857), .B(u5_cmd_asserted_bF_buf2), .Y(u5__abc_54027_n1845) );
  AND2X2 AND2X2_6638 ( .A(u5__abc_54027_n1318), .B(u5__abc_54027_n1316), .Y(u5__abc_54027_n1846) );
  AND2X2 AND2X2_6639 ( .A(u5__abc_54027_n387_1), .B(u5__abc_54027_n1347), .Y(u5__abc_54027_n1853) );
  AND2X2 AND2X2_664 ( .A(u0__abc_49347_n1175_bF_buf3), .B(u0__abc_49347_n2797), .Y(u0__abc_49347_n2798) );
  AND2X2 AND2X2_6640 ( .A(u5__abc_54027_n1326), .B(u5__abc_54027_n315), .Y(u5__abc_54027_n1855) );
  AND2X2 AND2X2_6641 ( .A(u5__abc_54027_n1858), .B(u5__abc_54027_n422), .Y(u5__abc_54027_n1859) );
  AND2X2 AND2X2_6642 ( .A(u5__abc_54027_n1859), .B(u5__abc_54027_n1857), .Y(u5__abc_54027_n1860) );
  AND2X2 AND2X2_6643 ( .A(u5__abc_54027_n424), .B(u5__abc_54027_n456), .Y(u5__abc_54027_n1861) );
  AND2X2 AND2X2_6644 ( .A(u5__abc_54027_n420), .B(u5__abc_54027_n480), .Y(u5__abc_54027_n1862) );
  AND2X2 AND2X2_6645 ( .A(u5__abc_54027_n619), .B(u5__abc_54027_n598), .Y(u5__abc_54027_n1869) );
  AND2X2 AND2X2_6646 ( .A(u5__abc_54027_n1876), .B(u5__abc_54027_n1877), .Y(u5__abc_54027_n1878) );
  AND2X2 AND2X2_6647 ( .A(u5_no_wb_cycle_FF_INPUT), .B(u5__abc_54027_n1878), .Y(u5__abc_54027_n1879) );
  AND2X2 AND2X2_6648 ( .A(u5__abc_54027_n1879), .B(u5__abc_54027_n513_1), .Y(u5__abc_54027_n1880) );
  AND2X2 AND2X2_6649 ( .A(u5__abc_54027_n1880), .B(u5__abc_54027_n873), .Y(u5__abc_54027_n1881) );
  AND2X2 AND2X2_665 ( .A(u0__abc_49347_n2796), .B(u0__abc_49347_n2798), .Y(u0__abc_49347_n2799) );
  AND2X2 AND2X2_6650 ( .A(u5__abc_54027_n1563), .B(u5__abc_54027_n596), .Y(u5__abc_54027_n1884) );
  AND2X2 AND2X2_6651 ( .A(u5__abc_54027_n1885), .B(u5__abc_54027_n511), .Y(u5__abc_54027_n1886) );
  AND2X2 AND2X2_6652 ( .A(u5__abc_54027_n1887), .B(u5__abc_54027_n351_bF_buf0), .Y(u5__abc_54027_n1888) );
  AND2X2 AND2X2_6653 ( .A(u5__abc_54027_n477), .B(u5_tmr_done), .Y(u5__abc_54027_n1889) );
  AND2X2 AND2X2_6654 ( .A(u5__abc_54027_n1523), .B(u5__abc_54027_n503), .Y(u5__abc_54027_n1890) );
  AND2X2 AND2X2_6655 ( .A(u5__abc_54027_n1839), .B(u5_wb_cycle), .Y(u5__abc_54027_n1891) );
  AND2X2 AND2X2_6656 ( .A(u5__abc_54027_n1892), .B(u5__abc_54027_n1889), .Y(u5__abc_54027_n1893) );
  AND2X2 AND2X2_6657 ( .A(u5__abc_54027_n1474), .B(u5__abc_54027_n1471), .Y(u5__abc_54027_n1894) );
  AND2X2 AND2X2_6658 ( .A(u5__abc_54027_n1895), .B(u5_wb_cycle), .Y(u5__abc_54027_n1896) );
  AND2X2 AND2X2_6659 ( .A(u5__abc_54027_n1904), .B(u5__abc_54027_n971), .Y(u5__abc_54027_n1905) );
  AND2X2 AND2X2_666 ( .A(u0__abc_49347_n1176_1_bF_buf3), .B(tms_3_), .Y(u0__abc_49347_n2801) );
  AND2X2 AND2X2_6660 ( .A(u5__abc_54027_n1361), .B(u5__abc_54027_n1905), .Y(u5__abc_54027_n1906) );
  AND2X2 AND2X2_6661 ( .A(u5__abc_54027_n347), .B(u5__abc_54027_n561), .Y(u5__abc_54027_n1911) );
  AND2X2 AND2X2_6662 ( .A(u5__abc_54027_n377), .B(u5__abc_54027_n1346), .Y(u5__abc_54027_n1914) );
  AND2X2 AND2X2_6663 ( .A(u5__abc_54027_n1915), .B(u5_tmr2_done), .Y(next_adr) );
  AND2X2 AND2X2_6664 ( .A(u5__abc_54027_n473), .B(u5__abc_54027_n519), .Y(u5__abc_54027_n1918) );
  AND2X2 AND2X2_6665 ( .A(u5__abc_54027_n1918), .B(u5__abc_54027_n648), .Y(u5__abc_54027_n1919) );
  AND2X2 AND2X2_6666 ( .A(u5__abc_54027_n424), .B(u5__abc_54027_n1921), .Y(u5__abc_54027_n1922) );
  AND2X2 AND2X2_6667 ( .A(u5__abc_54027_n1922), .B(u5__abc_54027_n454), .Y(u5__abc_54027_n1923) );
  AND2X2 AND2X2_6668 ( .A(u5__abc_54027_n1923), .B(u5__abc_54027_n1920), .Y(u5__abc_54027_n1924) );
  AND2X2 AND2X2_6669 ( .A(u5__abc_54027_n1926), .B(u5_cmd_a10_r), .Y(u5__abc_54027_n1927) );
  AND2X2 AND2X2_667 ( .A(u0_tms5_3_), .B(u0_cs5_bF_buf1), .Y(u0__abc_49347_n2802) );
  AND2X2 AND2X2_6670 ( .A(u5__abc_54027_n617), .B(u5__abc_54027_n1928), .Y(u5__abc_54027_n1929) );
  AND2X2 AND2X2_6671 ( .A(u5__abc_54027_n401), .B(u5__abc_54027_n1296), .Y(u5__abc_54027_n1934) );
  AND2X2 AND2X2_6672 ( .A(u5__abc_54027_n1934), .B(u5__abc_54027_n393), .Y(u5__abc_54027_n1935) );
  AND2X2 AND2X2_6673 ( .A(u5__abc_54027_n1935), .B(u5__abc_54027_n381), .Y(u5__abc_54027_n1936) );
  AND2X2 AND2X2_6674 ( .A(u5__abc_54027_n588), .B(u5__abc_54027_n599), .Y(u5__abc_54027_n1937) );
  AND2X2 AND2X2_6675 ( .A(u5__abc_54027_n1936), .B(u5__abc_54027_n1938), .Y(u5__abc_54027_n1939) );
  AND2X2 AND2X2_6676 ( .A(u5__abc_54027_n1933), .B(u5__abc_54027_n1939), .Y(u5_oe__FF_INPUT) );
  AND2X2 AND2X2_6677 ( .A(u5__abc_54027_n659), .B(u5__abc_54027_n434), .Y(u5__abc_54027_n1941) );
  AND2X2 AND2X2_6678 ( .A(u5__abc_54027_n1461), .B(u5__abc_54027_n1297), .Y(u5__abc_54027_n1942) );
  AND2X2 AND2X2_6679 ( .A(u5__abc_54027_n1941), .B(u5__abc_54027_n1942), .Y(u5__abc_54027_n1943) );
  AND2X2 AND2X2_668 ( .A(u0__abc_49347_n2804), .B(u0__abc_49347_n2730_bF_buf2), .Y(u0__abc_49347_n2805) );
  AND2X2 AND2X2_6680 ( .A(u5__abc_54027_n364), .B(u5__abc_54027_n458), .Y(u5__abc_54027_n1944) );
  AND2X2 AND2X2_6681 ( .A(u5__abc_54027_n368), .B(u5__abc_54027_n418), .Y(u5__abc_54027_n1945) );
  AND2X2 AND2X2_6682 ( .A(u5__abc_54027_n1945), .B(u5__abc_54027_n1944), .Y(u5__abc_54027_n1946) );
  AND2X2 AND2X2_6683 ( .A(u5__abc_54027_n1943), .B(u5__abc_54027_n1946), .Y(u5__abc_54027_n1947) );
  AND2X2 AND2X2_6684 ( .A(u5__abc_54027_n1559), .B(u5__abc_54027_n1401), .Y(u5__abc_54027_n1948) );
  AND2X2 AND2X2_6685 ( .A(u5__abc_54027_n1904), .B(u5__abc_54027_n1948), .Y(u5__abc_54027_n1949) );
  AND2X2 AND2X2_6686 ( .A(u5__abc_54027_n1949), .B(u5__abc_54027_n454), .Y(u5__abc_54027_n1950) );
  AND2X2 AND2X2_6687 ( .A(u5__abc_54027_n396), .B(u5__abc_54027_n400), .Y(u5__abc_54027_n1951) );
  AND2X2 AND2X2_6688 ( .A(u5__abc_54027_n1951), .B(u5__abc_54027_n1492), .Y(u5__abc_54027_n1952) );
  AND2X2 AND2X2_6689 ( .A(u5__abc_54027_n1954), .B(u5__abc_54027_n1953), .Y(u5__abc_54027_n1955) );
  AND2X2 AND2X2_669 ( .A(u0__abc_49347_n2805), .B(u0__abc_49347_n2803), .Y(u0__abc_49347_n2806) );
  AND2X2 AND2X2_6690 ( .A(u5__abc_54027_n1955), .B(u5__abc_54027_n1952), .Y(u5__abc_54027_n1956) );
  AND2X2 AND2X2_6691 ( .A(u5__abc_54027_n1956), .B(u5__abc_54027_n1950), .Y(u5__abc_54027_n1957) );
  AND2X2 AND2X2_6692 ( .A(u5__abc_54027_n1957), .B(u5__abc_54027_n1947), .Y(u5__abc_54027_n1958) );
  AND2X2 AND2X2_6693 ( .A(u5__abc_54027_n1530), .B(u5__abc_54027_n1750), .Y(u5__abc_54027_n1959) );
  AND2X2 AND2X2_6694 ( .A(u5__abc_54027_n1960), .B(u5__abc_54027_n1961), .Y(u5__abc_54027_n1962) );
  AND2X2 AND2X2_6695 ( .A(u5__abc_54027_n1962), .B(u5__abc_54027_n1959), .Y(u5__abc_54027_n1963) );
  AND2X2 AND2X2_6696 ( .A(u5__abc_54027_n308), .B(u5__abc_54027_n1963), .Y(u5__abc_54027_n1964) );
  AND2X2 AND2X2_6697 ( .A(u5__abc_54027_n393), .B(u5__abc_54027_n1047), .Y(u5__abc_54027_n1965) );
  AND2X2 AND2X2_6698 ( .A(u5__abc_54027_n1964), .B(u5__abc_54027_n1965), .Y(u5__abc_54027_n1966) );
  AND2X2 AND2X2_6699 ( .A(u5__abc_54027_n398), .B(u5__abc_54027_n378), .Y(u5__abc_54027_n1967) );
  AND2X2 AND2X2_67 ( .A(init_req), .B(u0_init_req2), .Y(u0__abc_49347_n1119) );
  AND2X2 AND2X2_670 ( .A(u0__abc_49347_n2807), .B(u0__abc_49347_n2726_bF_buf2), .Y(u0__abc_49347_n2808) );
  AND2X2 AND2X2_6700 ( .A(u5__abc_54027_n373), .B(u5__abc_54027_n1967), .Y(u5__abc_54027_n1968) );
  AND2X2 AND2X2_6701 ( .A(u5__abc_54027_n653), .B(u5__abc_54027_n444), .Y(u5__abc_54027_n1969) );
  AND2X2 AND2X2_6702 ( .A(u5__abc_54027_n1306), .B(u5__abc_54027_n1970), .Y(u5__abc_54027_n1971) );
  AND2X2 AND2X2_6703 ( .A(u5__abc_54027_n1969), .B(u5__abc_54027_n1971), .Y(u5__abc_54027_n1972) );
  AND2X2 AND2X2_6704 ( .A(u5__abc_54027_n1968), .B(u5__abc_54027_n1972), .Y(u5__abc_54027_n1973) );
  AND2X2 AND2X2_6705 ( .A(u5__abc_54027_n853), .B(u5__abc_54027_n1974), .Y(u5__abc_54027_n1975) );
  AND2X2 AND2X2_6706 ( .A(u5__abc_54027_n1976), .B(u5__abc_54027_n1977), .Y(u5__abc_54027_n1978) );
  AND2X2 AND2X2_6707 ( .A(u5__abc_54027_n1975), .B(u5__abc_54027_n1978), .Y(u5__abc_54027_n1979) );
  AND2X2 AND2X2_6708 ( .A(u5__abc_54027_n1980), .B(u5__abc_54027_n406), .Y(u5__abc_54027_n1981) );
  AND2X2 AND2X2_6709 ( .A(u5__abc_54027_n448), .B(u5__abc_54027_n429_1), .Y(u5__abc_54027_n1982) );
  AND2X2 AND2X2_671 ( .A(u0_tms4_3_), .B(u0_cs4_bF_buf1), .Y(u0__abc_49347_n2809) );
  AND2X2 AND2X2_6710 ( .A(u5__abc_54027_n1981), .B(u5__abc_54027_n1982), .Y(u5__abc_54027_n1983) );
  AND2X2 AND2X2_6711 ( .A(u5__abc_54027_n1983), .B(u5__abc_54027_n1979), .Y(u5__abc_54027_n1984) );
  AND2X2 AND2X2_6712 ( .A(u5__abc_54027_n1973), .B(u5__abc_54027_n1984), .Y(u5__abc_54027_n1985) );
  AND2X2 AND2X2_6713 ( .A(u5__abc_54027_n1966), .B(u5__abc_54027_n1985), .Y(u5__abc_54027_n1986) );
  AND2X2 AND2X2_6714 ( .A(u5__abc_54027_n1986), .B(u5__abc_54027_n1958), .Y(u5_suspended_d) );
  AND2X2 AND2X2_6715 ( .A(u5__abc_54027_n870), .B(u5_cke_r), .Y(u5__abc_54027_n1988) );
  AND2X2 AND2X2_6716 ( .A(u5_cnt), .B(u5_wb_cycle), .Y(u5__abc_54027_n1989) );
  AND2X2 AND2X2_6717 ( .A(u5__abc_54027_n1326), .B(u5__abc_54027_n1989), .Y(u5__abc_54027_n1990) );
  AND2X2 AND2X2_6718 ( .A(u5__abc_54027_n1990), .B(u5__abc_54027_n477), .Y(u5__abc_54027_n1991) );
  AND2X2 AND2X2_6719 ( .A(u5__abc_54027_n1992), .B(_auto_iopadmap_cc_313_execute_56251), .Y(u5__abc_54027_n1993) );
  AND2X2 AND2X2_672 ( .A(u0__abc_49347_n2810), .B(u0__abc_49347_n2725_bF_buf2), .Y(u0__abc_49347_n2811) );
  AND2X2 AND2X2_6720 ( .A(u5__abc_54027_n1995), .B(u5__abc_54027_n1988), .Y(u5_cke__FF_INPUT) );
  AND2X2 AND2X2_6721 ( .A(wb_stb_i_bF_buf4), .B(wb_cyc_i), .Y(u5__abc_54027_n1997) );
  AND2X2 AND2X2_6722 ( .A(u5__abc_54027_n1997), .B(cs_le_bF_buf2), .Y(u5_lookup_ready1_FF_INPUT) );
  AND2X2 AND2X2_6723 ( .A(u5__abc_54027_n1997), .B(u5_lookup_ready1), .Y(u5_lookup_ready2_FF_INPUT) );
  AND2X2 AND2X2_6724 ( .A(u5__abc_54027_n1107), .B(u5__abc_54027_n1142), .Y(u5__abc_54027_n2001) );
  AND2X2 AND2X2_6725 ( .A(u5__abc_54027_n2001), .B(u5__abc_54027_n1112), .Y(u5__abc_54027_n2002) );
  AND2X2 AND2X2_6726 ( .A(u5__abc_54027_n2000), .B(u5__abc_54027_n2002), .Y(u5_tmr2_done_FF_INPUT) );
  AND2X2 AND2X2_6727 ( .A(u5__abc_54027_n387_1), .B(u5__abc_54027_n2004), .Y(u5_pack_le2_d) );
  AND2X2 AND2X2_6728 ( .A(u5__abc_54027_n2006), .B(u5__abc_54027_n314), .Y(u5_cnt_next) );
  AND2X2 AND2X2_6729 ( .A(u5__abc_54027_n646), .B(u5_kro), .Y(bank_set) );
  AND2X2 AND2X2_673 ( .A(u0_tms3_3_), .B(u0_cs3_bF_buf1), .Y(u0__abc_49347_n2812) );
  AND2X2 AND2X2_6730 ( .A(u5__abc_54027_n2009), .B(susp_sel), .Y(u5__abc_54027_n2010) );
  AND2X2 AND2X2_6731 ( .A(u5_wb_cycle), .B(wb_cyc_i), .Y(u5__abc_54027_n2013) );
  AND2X2 AND2X2_6732 ( .A(u5__abc_54027_n2013), .B(u5__abc_54027_n2012), .Y(u5__abc_54027_n2014) );
  AND2X2 AND2X2_6733 ( .A(u5__abc_54027_n414), .B(u1_wr_cycle), .Y(u5__abc_54027_n2016) );
  AND2X2 AND2X2_6734 ( .A(u5__abc_54027_n1725), .B(u5__abc_54027_n1563), .Y(u5__abc_54027_n2019) );
  AND2X2 AND2X2_6735 ( .A(u5__abc_54027_n2020), .B(u5__abc_54027_n2017), .Y(u5__abc_54027_n2021) );
  AND2X2 AND2X2_6736 ( .A(wb_cyc_i), .B(wb_stb_i_bF_buf3), .Y(u6__abc_56056_n132) );
  AND2X2 AND2X2_6737 ( .A(u6__abc_56056_n135_1), .B(u6__abc_56056_n136), .Y(u6__abc_56056_n137) );
  AND2X2 AND2X2_6738 ( .A(u6__abc_56056_n137), .B(u6__abc_56056_n134), .Y(u6__abc_56056_n138_1) );
  AND2X2 AND2X2_6739 ( .A(u6__abc_56056_n141_1), .B(u6__abc_56056_n142_1), .Y(u6__abc_56056_n143) );
  AND2X2 AND2X2_674 ( .A(u0__abc_49347_n2813), .B(u0__abc_49347_n2724_bF_buf2), .Y(u0__abc_49347_n2814) );
  AND2X2 AND2X2_6740 ( .A(u6__abc_56056_n143), .B(u6__abc_56056_n140_1), .Y(u6__abc_56056_n144) );
  AND2X2 AND2X2_6741 ( .A(u6__abc_56056_n144_bF_buf5), .B(mem_ack), .Y(u6__abc_56056_n145_1) );
  AND2X2 AND2X2_6742 ( .A(u6__abc_56056_n139_1), .B(u6__abc_56056_n145_1), .Y(u6__abc_56056_n146_1) );
  AND2X2 AND2X2_6743 ( .A(u6__abc_56056_n140_1), .B(\wb_addr_i[29] ), .Y(u6__abc_56056_n147) );
  AND2X2 AND2X2_6744 ( .A(u6__abc_56056_n148_1), .B(\wb_addr_i[30] ), .Y(u6__abc_56056_n149_1) );
  AND2X2 AND2X2_6745 ( .A(u6__abc_56056_n149_1), .B(u6__abc_56056_n132), .Y(u6__abc_56056_n150_1) );
  AND2X2 AND2X2_6746 ( .A(u6__abc_56056_n150_1), .B(u6__abc_56056_n147), .Y(u6__abc_56056_n151) );
  AND2X2 AND2X2_6747 ( .A(u6__abc_56056_n155_1), .B(u6__abc_56056_n153), .Y(u6_wb_data_o_0__FF_INPUT) );
  AND2X2 AND2X2_6748 ( .A(u6__abc_56056_n158), .B(u6__abc_56056_n157_1), .Y(u6_wb_data_o_1__FF_INPUT) );
  AND2X2 AND2X2_6749 ( .A(u6__abc_56056_n161), .B(u6__abc_56056_n160), .Y(u6_wb_data_o_2__FF_INPUT) );
  AND2X2 AND2X2_675 ( .A(u0_tms2_3_), .B(u0_cs2_bF_buf1), .Y(u0__abc_49347_n2815) );
  AND2X2 AND2X2_6750 ( .A(u6__abc_56056_n164), .B(u6__abc_56056_n163_1), .Y(u6_wb_data_o_3__FF_INPUT) );
  AND2X2 AND2X2_6751 ( .A(u6__abc_56056_n167_1), .B(u6__abc_56056_n166_1), .Y(u6_wb_data_o_4__FF_INPUT) );
  AND2X2 AND2X2_6752 ( .A(u6__abc_56056_n170), .B(u6__abc_56056_n169), .Y(u6_wb_data_o_5__FF_INPUT) );
  AND2X2 AND2X2_6753 ( .A(u6__abc_56056_n173), .B(u6__abc_56056_n172), .Y(u6_wb_data_o_6__FF_INPUT) );
  AND2X2 AND2X2_6754 ( .A(u6__abc_56056_n176), .B(u6__abc_56056_n175), .Y(u6_wb_data_o_7__FF_INPUT) );
  AND2X2 AND2X2_6755 ( .A(u6__abc_56056_n179), .B(u6__abc_56056_n178), .Y(u6_wb_data_o_8__FF_INPUT) );
  AND2X2 AND2X2_6756 ( .A(u6__abc_56056_n182), .B(u6__abc_56056_n181), .Y(u6_wb_data_o_9__FF_INPUT) );
  AND2X2 AND2X2_6757 ( .A(u6__abc_56056_n185), .B(u6__abc_56056_n184), .Y(u6_wb_data_o_10__FF_INPUT) );
  AND2X2 AND2X2_6758 ( .A(u6__abc_56056_n188), .B(u6__abc_56056_n187), .Y(u6_wb_data_o_11__FF_INPUT) );
  AND2X2 AND2X2_6759 ( .A(u6__abc_56056_n191), .B(u6__abc_56056_n190), .Y(u6_wb_data_o_12__FF_INPUT) );
  AND2X2 AND2X2_676 ( .A(u0__abc_49347_n2816_1), .B(u0__abc_49347_n2723_bF_buf2), .Y(u0__abc_49347_n2817) );
  AND2X2 AND2X2_6760 ( .A(u6__abc_56056_n194), .B(u6__abc_56056_n193), .Y(u6_wb_data_o_13__FF_INPUT) );
  AND2X2 AND2X2_6761 ( .A(u6__abc_56056_n197), .B(u6__abc_56056_n196), .Y(u6_wb_data_o_14__FF_INPUT) );
  AND2X2 AND2X2_6762 ( .A(u6__abc_56056_n200), .B(u6__abc_56056_n199), .Y(u6_wb_data_o_15__FF_INPUT) );
  AND2X2 AND2X2_6763 ( .A(u6__abc_56056_n203), .B(u6__abc_56056_n202), .Y(u6_wb_data_o_16__FF_INPUT) );
  AND2X2 AND2X2_6764 ( .A(u6__abc_56056_n206), .B(u6__abc_56056_n205), .Y(u6_wb_data_o_17__FF_INPUT) );
  AND2X2 AND2X2_6765 ( .A(u6__abc_56056_n209), .B(u6__abc_56056_n208), .Y(u6_wb_data_o_18__FF_INPUT) );
  AND2X2 AND2X2_6766 ( .A(u6__abc_56056_n212), .B(u6__abc_56056_n211), .Y(u6_wb_data_o_19__FF_INPUT) );
  AND2X2 AND2X2_6767 ( .A(u6__abc_56056_n215), .B(u6__abc_56056_n214), .Y(u6_wb_data_o_20__FF_INPUT) );
  AND2X2 AND2X2_6768 ( .A(u6__abc_56056_n218), .B(u6__abc_56056_n217), .Y(u6_wb_data_o_21__FF_INPUT) );
  AND2X2 AND2X2_6769 ( .A(u6__abc_56056_n221), .B(u6__abc_56056_n220), .Y(u6_wb_data_o_22__FF_INPUT) );
  AND2X2 AND2X2_677 ( .A(u0_tms1_3_), .B(u0_cs1_bF_buf1), .Y(u0__abc_49347_n2818) );
  AND2X2 AND2X2_6770 ( .A(u6__abc_56056_n224), .B(u6__abc_56056_n223), .Y(u6_wb_data_o_23__FF_INPUT) );
  AND2X2 AND2X2_6771 ( .A(u6__abc_56056_n227), .B(u6__abc_56056_n226), .Y(u6_wb_data_o_24__FF_INPUT) );
  AND2X2 AND2X2_6772 ( .A(u6__abc_56056_n230), .B(u6__abc_56056_n229), .Y(u6_wb_data_o_25__FF_INPUT) );
  AND2X2 AND2X2_6773 ( .A(u6__abc_56056_n233), .B(u6__abc_56056_n232), .Y(u6_wb_data_o_26__FF_INPUT) );
  AND2X2 AND2X2_6774 ( .A(u6__abc_56056_n236), .B(u6__abc_56056_n235), .Y(u6_wb_data_o_27__FF_INPUT) );
  AND2X2 AND2X2_6775 ( .A(u6__abc_56056_n239), .B(u6__abc_56056_n238), .Y(u6_wb_data_o_28__FF_INPUT) );
  AND2X2 AND2X2_6776 ( .A(u6__abc_56056_n242), .B(u6__abc_56056_n241), .Y(u6_wb_data_o_29__FF_INPUT) );
  AND2X2 AND2X2_6777 ( .A(u6__abc_56056_n245), .B(u6__abc_56056_n244), .Y(u6_wb_data_o_30__FF_INPUT) );
  AND2X2 AND2X2_6778 ( .A(u6__abc_56056_n248), .B(u6__abc_56056_n247), .Y(u6_wb_data_o_31__FF_INPUT) );
  AND2X2 AND2X2_6779 ( .A(u6__abc_56056_n132), .B(wb_we_i), .Y(u6__abc_56056_n250) );
  AND2X2 AND2X2_678 ( .A(u0__abc_49347_n1175_bF_buf2), .B(u0__abc_49347_n2821), .Y(u0__abc_49347_n2822) );
  AND2X2 AND2X2_6780 ( .A(u6__abc_56056_n133), .B(u1_wr_hold), .Y(u6__abc_56056_n251) );
  AND2X2 AND2X2_6781 ( .A(u6__abc_56056_n253), .B(u6_rmw_en), .Y(u6__abc_56056_n254) );
  AND2X2 AND2X2_6782 ( .A(u6__abc_56056_n250), .B(u6__abc_56056_n254), .Y(u6_rmw_r_FF_INPUT) );
  AND2X2 AND2X2_6783 ( .A(u6__abc_56056_n144_bF_buf1), .B(wb_stb_i_bF_buf2), .Y(u6__abc_56056_n257) );
  AND2X2 AND2X2_6784 ( .A(u6__abc_56056_n257), .B(u6__abc_56056_n256), .Y(u6__abc_56056_n258) );
  AND2X2 AND2X2_6785 ( .A(u6__abc_56056_n261), .B(u6__abc_56056_n260), .Y(u6__abc_56056_n262) );
  AND2X2 AND2X2_6786 ( .A(u6__abc_56056_n262), .B(wb_cyc_i), .Y(u6__abc_56056_n263) );
  AND2X2 AND2X2_6787 ( .A(u6__abc_56056_n259), .B(u6__abc_56056_n263), .Y(u6_read_go_r1_FF_INPUT) );
  AND2X2 AND2X2_6788 ( .A(wb_cyc_i), .B(u6_read_go_r1), .Y(u6_read_go_r_FF_INPUT) );
  AND2X2 AND2X2_6789 ( .A(u6__abc_56056_n262), .B(u6_read_go_r_FF_INPUT), .Y(u3_wb_read_go) );
  AND2X2 AND2X2_679 ( .A(u0__abc_49347_n2820), .B(u0__abc_49347_n2822), .Y(u0__abc_49347_n2823) );
  AND2X2 AND2X2_6790 ( .A(u6__abc_56056_n257), .B(wb_we_i), .Y(u6__abc_56056_n267) );
  AND2X2 AND2X2_6791 ( .A(u6__abc_56056_n268), .B(wb_cyc_i), .Y(u6_write_go_r1_FF_INPUT) );
  AND2X2 AND2X2_6792 ( .A(wb_cyc_i), .B(u6_write_go_r1), .Y(u6__abc_56056_n272) );
  AND2X2 AND2X2_6793 ( .A(u6__abc_56056_n271), .B(u6__abc_56056_n272), .Y(u6_write_go_r_FF_INPUT) );
  AND2X2 AND2X2_6794 ( .A(u6__abc_56056_n262), .B(u6_write_go_r_FF_INPUT), .Y(u1_wb_write_go) );
  AND2X2 AND2X2_6795 ( .A(u6__abc_56056_n275), .B(u6__abc_56056_n276), .Y(u6__abc_56056_n277) );
  AND2X2 AND2X2_6796 ( .A(u6__abc_56056_n277), .B(u6__abc_56056_n132), .Y(u6__abc_56056_n278) );
  AND2X2 AND2X2_6797 ( .A(u6__abc_56056_n144_bF_buf0), .B(u6__abc_56056_n278), .Y(u6__abc_56056_n279) );
  AND2X2 AND2X2_6798 ( .A(u6__abc_56056_n148_1), .B(u6_wb_first_r), .Y(u6__abc_56056_n281) );
  AND2X2 AND2X2_6799 ( .A(u6__abc_56056_n281), .B(u6__abc_56056_n280), .Y(u6__abc_56056_n282) );
  AND2X2 AND2X2_68 ( .A(u0__abc_49347_n1117_1), .B(u0__abc_49347_n1120_1), .Y(u0__abc_49347_n1121) );
  AND2X2 AND2X2_680 ( .A(u0__abc_49347_n1176_1_bF_buf2), .B(tms_4_), .Y(u0__abc_49347_n2825) );
  AND2X2 AND2X2_6800 ( .A(u6__abc_56056_n144_bF_buf5), .B(u6__abc_56056_n280), .Y(u6__abc_56056_n285) );
  AND2X2 AND2X2_6801 ( .A(u6__abc_56056_n284), .B(u6__abc_56056_n285), .Y(u6_wb_err_FF_INPUT) );
  AND2X2 AND2X2_6802 ( .A(u6__abc_56056_n270), .B(wb_cyc_i), .Y(u6__abc_56056_n288) );
  AND2X2 AND2X2_6803 ( .A(u6__abc_56056_n287), .B(u6__abc_56056_n288), .Y(u5_wb_wait) );
  AND2X2 AND2X2_6804 ( .A(wb_cyc_i), .B(u6_rmw_en), .Y(u6__abc_56056_n290) );
  AND2X2 AND2X2_6805 ( .A(u7__abc_47535_n75_1), .B(data_oe), .Y(u7__abc_47535_n76) );
  AND2X2 AND2X2_6806 ( .A(u7__abc_47535_n79_1), .B(u7__abc_47535_n77_1), .Y(u7__abc_47535_n80_1) );
  AND2X2 AND2X2_6807 ( .A(u7__abc_47535_n83_1), .B(data_oe), .Y(u7__abc_47535_n84) );
  AND2X2 AND2X2_6808 ( .A(u7__abc_47535_n86_1), .B(data_oe), .Y(u7__abc_47535_n87_1) );
  AND2X2 AND2X2_6809 ( .A(u7__abc_47535_n89_1), .B(data_oe), .Y(u7__abc_47535_n90_1) );
  AND2X2 AND2X2_681 ( .A(u0_tms5_4_), .B(u0_cs5_bF_buf0), .Y(u0__abc_49347_n2826) );
  AND2X2 AND2X2_6810 ( .A(wb_stb_i_bF_buf0), .B(wb_cyc_i), .Y(u7__abc_47535_n92_1) );
  AND2X2 AND2X2_6811 ( .A(u7__abc_47535_n92_1), .B(\wb_sel_i[0] ), .Y(u7__abc_47535_n93) );
  AND2X2 AND2X2_6812 ( .A(u7__abc_47535_n94_1), .B(u7_mc_dqm_r_0_), .Y(u7__abc_47535_n95_1) );
  AND2X2 AND2X2_6813 ( .A(u7__abc_47535_n92_1), .B(\wb_sel_i[1] ), .Y(u7__abc_47535_n97_1) );
  AND2X2 AND2X2_6814 ( .A(u7__abc_47535_n94_1), .B(u7_mc_dqm_r_1_), .Y(u7__abc_47535_n98_1) );
  AND2X2 AND2X2_6815 ( .A(u7__abc_47535_n92_1), .B(\wb_sel_i[2] ), .Y(u7__abc_47535_n100) );
  AND2X2 AND2X2_6816 ( .A(u7__abc_47535_n94_1), .B(u7_mc_dqm_r_2_), .Y(u7__abc_47535_n101) );
  AND2X2 AND2X2_6817 ( .A(u7__abc_47535_n92_1), .B(\wb_sel_i[3] ), .Y(u7__abc_47535_n103) );
  AND2X2 AND2X2_6818 ( .A(u7__abc_47535_n94_1), .B(u7_mc_dqm_r_3_), .Y(u7__abc_47535_n104) );
  AND2X2 AND2X2_6819 ( .A(spec_req_cs_0_bF_buf5), .B(lmr_sel_bF_buf1), .Y(u7__abc_47535_n110) );
  AND2X2 AND2X2_682 ( .A(u0__abc_49347_n2828), .B(u0__abc_49347_n2730_bF_buf1), .Y(u0__abc_49347_n2829) );
  AND2X2 AND2X2_6820 ( .A(u7__abc_47535_n109), .B(u7__abc_47535_n111), .Y(u7__abc_47535_n112) );
  AND2X2 AND2X2_6821 ( .A(u7__abc_47535_n112), .B(u7__abc_47535_n107), .Y(u7__abc_47535_n113) );
  AND2X2 AND2X2_6822 ( .A(u7__abc_47535_n106), .B(u7__abc_47535_n115), .Y(u7__abc_47535_n116) );
  AND2X2 AND2X2_6823 ( .A(lmr_sel_bF_buf6), .B(spec_req_cs_1_bF_buf5), .Y(u7__abc_47535_n121) );
  AND2X2 AND2X2_6824 ( .A(u7__abc_47535_n120), .B(u7__abc_47535_n122), .Y(u7__abc_47535_n123) );
  AND2X2 AND2X2_6825 ( .A(u7__abc_47535_n123), .B(u7__abc_47535_n107), .Y(u7__abc_47535_n124) );
  AND2X2 AND2X2_6826 ( .A(u7__abc_47535_n106), .B(u7__abc_47535_n125), .Y(u7__abc_47535_n126) );
  AND2X2 AND2X2_6827 ( .A(lmr_sel_bF_buf4), .B(spec_req_cs_2_bF_buf5), .Y(u7__abc_47535_n131) );
  AND2X2 AND2X2_6828 ( .A(u7__abc_47535_n130), .B(u7__abc_47535_n132), .Y(u7__abc_47535_n133) );
  AND2X2 AND2X2_6829 ( .A(u7__abc_47535_n133), .B(u7__abc_47535_n107), .Y(u7__abc_47535_n134) );
  AND2X2 AND2X2_683 ( .A(u0__abc_49347_n2829), .B(u0__abc_49347_n2827), .Y(u0__abc_49347_n2830) );
  AND2X2 AND2X2_6830 ( .A(u7__abc_47535_n106), .B(u7__abc_47535_n135), .Y(u7__abc_47535_n136) );
  AND2X2 AND2X2_6831 ( .A(lmr_sel_bF_buf2), .B(spec_req_cs_3_bF_buf5), .Y(u7__abc_47535_n141) );
  AND2X2 AND2X2_6832 ( .A(u7__abc_47535_n140), .B(u7__abc_47535_n142), .Y(u7__abc_47535_n143) );
  AND2X2 AND2X2_6833 ( .A(u7__abc_47535_n143), .B(u7__abc_47535_n107), .Y(u7__abc_47535_n144) );
  AND2X2 AND2X2_6834 ( .A(u7__abc_47535_n106), .B(u7__abc_47535_n145), .Y(u7__abc_47535_n146) );
  AND2X2 AND2X2_6835 ( .A(lmr_sel_bF_buf0), .B(spec_req_cs_4_bF_buf5), .Y(u7__abc_47535_n151) );
  AND2X2 AND2X2_6836 ( .A(u7__abc_47535_n150), .B(u7__abc_47535_n152), .Y(u7__abc_47535_n153) );
  AND2X2 AND2X2_6837 ( .A(u7__abc_47535_n153), .B(u7__abc_47535_n107), .Y(u7__abc_47535_n154) );
  AND2X2 AND2X2_6838 ( .A(u7__abc_47535_n106), .B(u7__abc_47535_n155), .Y(u7__abc_47535_n156) );
  AND2X2 AND2X2_6839 ( .A(lmr_sel_bF_buf5), .B(spec_req_cs_5_bF_buf5), .Y(u7__abc_47535_n161) );
  AND2X2 AND2X2_684 ( .A(u0__abc_49347_n2831), .B(u0__abc_49347_n2726_bF_buf1), .Y(u0__abc_49347_n2832) );
  AND2X2 AND2X2_6840 ( .A(u7__abc_47535_n160), .B(u7__abc_47535_n162), .Y(u7__abc_47535_n163) );
  AND2X2 AND2X2_6841 ( .A(u7__abc_47535_n163), .B(u7__abc_47535_n107), .Y(u7__abc_47535_n164) );
  AND2X2 AND2X2_6842 ( .A(u7__abc_47535_n106), .B(u7__abc_47535_n165), .Y(u7__abc_47535_n166) );
  AND2X2 AND2X2_6843 ( .A(lmr_sel_bF_buf3), .B(spec_req_cs_6_bF_buf1), .Y(u7__abc_47535_n171) );
  AND2X2 AND2X2_6844 ( .A(u7__abc_47535_n170), .B(u7__abc_47535_n172), .Y(u7__abc_47535_n173) );
  AND2X2 AND2X2_6845 ( .A(u7__abc_47535_n173), .B(u7__abc_47535_n107), .Y(u7__abc_47535_n174) );
  AND2X2 AND2X2_6846 ( .A(u7__abc_47535_n106), .B(u7__abc_47535_n175), .Y(u7__abc_47535_n176) );
  AND2X2 AND2X2_6847 ( .A(lmr_sel_bF_buf1), .B(spec_req_cs_7_), .Y(u7__abc_47535_n181) );
  AND2X2 AND2X2_6848 ( .A(u7__abc_47535_n180), .B(u7__abc_47535_n182), .Y(u7__abc_47535_n183) );
  AND2X2 AND2X2_6849 ( .A(u7__abc_47535_n183), .B(u7__abc_47535_n107), .Y(u7__abc_47535_n184) );
  AND2X2 AND2X2_685 ( .A(u0_tms4_4_), .B(u0_cs4_bF_buf0), .Y(u0__abc_49347_n2833) );
  AND2X2 AND2X2_6850 ( .A(u7__abc_47535_n106), .B(u7__abc_47535_n185), .Y(u7__abc_47535_n186) );
  AND2X2 AND2X2_6851 ( .A(u7__abc_47535_n191), .B(u7__abc_47535_n192), .Y(u7_mc_rp_FF_INPUT) );
  AND2X2 AND2X2_6852 ( .A(data_oe), .B(mc_c_oe_d), .Y(u7__abc_47535_n195) );
  AND2X2 AND2X2_6853 ( .A(u7__abc_47535_n195), .B(u7__abc_47535_n194), .Y(u7_mc_data_oe_FF_INPUT) );
  AND2X2 AND2X2_686 ( .A(u0__abc_49347_n2834), .B(u0__abc_49347_n2725_bF_buf1), .Y(u0__abc_49347_n2835) );
  AND2X2 AND2X2_687 ( .A(u0_tms3_4_), .B(u0_cs3_bF_buf0), .Y(u0__abc_49347_n2836) );
  AND2X2 AND2X2_688 ( .A(u0__abc_49347_n2837), .B(u0__abc_49347_n2724_bF_buf1), .Y(u0__abc_49347_n2838) );
  AND2X2 AND2X2_689 ( .A(u0_tms2_4_), .B(u0_cs2_bF_buf0), .Y(u0__abc_49347_n2839) );
  AND2X2 AND2X2_69 ( .A(u0__abc_49347_n1105_1), .B(u0__abc_49347_n1121), .Y(u0__abc_49347_n1122_1) );
  AND2X2 AND2X2_690 ( .A(u0__abc_49347_n2840), .B(u0__abc_49347_n2723_bF_buf1), .Y(u0__abc_49347_n2841) );
  AND2X2 AND2X2_691 ( .A(u0_tms1_4_), .B(u0_cs1_bF_buf0), .Y(u0__abc_49347_n2842) );
  AND2X2 AND2X2_692 ( .A(u0__abc_49347_n1175_bF_buf1), .B(u0__abc_49347_n2845), .Y(u0__abc_49347_n2846) );
  AND2X2 AND2X2_693 ( .A(u0__abc_49347_n2844), .B(u0__abc_49347_n2846), .Y(u0__abc_49347_n2847) );
  AND2X2 AND2X2_694 ( .A(u0__abc_49347_n1176_1_bF_buf1), .B(tms_5_), .Y(u0__abc_49347_n2849) );
  AND2X2 AND2X2_695 ( .A(u0_tms5_5_), .B(u0_cs5_bF_buf5), .Y(u0__abc_49347_n2850) );
  AND2X2 AND2X2_696 ( .A(u0__abc_49347_n2852), .B(u0__abc_49347_n2730_bF_buf0), .Y(u0__abc_49347_n2853) );
  AND2X2 AND2X2_697 ( .A(u0__abc_49347_n2853), .B(u0__abc_49347_n2851), .Y(u0__abc_49347_n2854) );
  AND2X2 AND2X2_698 ( .A(u0__abc_49347_n2855), .B(u0__abc_49347_n2726_bF_buf0), .Y(u0__abc_49347_n2856) );
  AND2X2 AND2X2_699 ( .A(u0_tms4_5_), .B(u0_cs4_bF_buf5), .Y(u0__abc_49347_n2857) );
  AND2X2 AND2X2_7 ( .A(_abc_55805_n257), .B(_abc_55805_n258), .Y(obct_cs_2_) );
  AND2X2 AND2X2_70 ( .A(u0__abc_49347_n1113_1), .B(spec_req_cs_3_bF_buf4), .Y(u0__abc_49347_n1124_1) );
  AND2X2 AND2X2_700 ( .A(u0__abc_49347_n2858), .B(u0__abc_49347_n2725_bF_buf0), .Y(u0__abc_49347_n2859) );
  AND2X2 AND2X2_701 ( .A(u0_tms3_5_), .B(u0_cs3_bF_buf5), .Y(u0__abc_49347_n2860) );
  AND2X2 AND2X2_702 ( .A(u0__abc_49347_n2861), .B(u0__abc_49347_n2724_bF_buf0), .Y(u0__abc_49347_n2862) );
  AND2X2 AND2X2_703 ( .A(u0_tms2_5_), .B(u0_cs2_bF_buf5), .Y(u0__abc_49347_n2863) );
  AND2X2 AND2X2_704 ( .A(u0__abc_49347_n2864), .B(u0__abc_49347_n2723_bF_buf0), .Y(u0__abc_49347_n2865) );
  AND2X2 AND2X2_705 ( .A(u0_tms1_5_), .B(u0_cs1_bF_buf5), .Y(u0__abc_49347_n2866) );
  AND2X2 AND2X2_706 ( .A(u0__abc_49347_n1175_bF_buf0), .B(u0__abc_49347_n2869), .Y(u0__abc_49347_n2870) );
  AND2X2 AND2X2_707 ( .A(u0__abc_49347_n2868), .B(u0__abc_49347_n2870), .Y(u0__abc_49347_n2871) );
  AND2X2 AND2X2_708 ( .A(u0__abc_49347_n1176_1_bF_buf0), .B(tms_6_), .Y(u0__abc_49347_n2873) );
  AND2X2 AND2X2_709 ( .A(u0_tms5_6_), .B(u0_cs5_bF_buf4), .Y(u0__abc_49347_n2874) );
  AND2X2 AND2X2_71 ( .A(u0__abc_49347_n1117_1), .B(u0__abc_49347_n1125), .Y(u0__abc_49347_n1126_1) );
  AND2X2 AND2X2_710 ( .A(u0__abc_49347_n2876), .B(u0__abc_49347_n2730_bF_buf5), .Y(u0__abc_49347_n2877) );
  AND2X2 AND2X2_711 ( .A(u0__abc_49347_n2877), .B(u0__abc_49347_n2875), .Y(u0__abc_49347_n2878) );
  AND2X2 AND2X2_712 ( .A(u0__abc_49347_n2879), .B(u0__abc_49347_n2726_bF_buf5), .Y(u0__abc_49347_n2880) );
  AND2X2 AND2X2_713 ( .A(u0_tms4_6_), .B(u0_cs4_bF_buf4), .Y(u0__abc_49347_n2881_1) );
  AND2X2 AND2X2_714 ( .A(u0__abc_49347_n2882), .B(u0__abc_49347_n2725_bF_buf5), .Y(u0__abc_49347_n2883) );
  AND2X2 AND2X2_715 ( .A(u0_tms3_6_), .B(u0_cs3_bF_buf4), .Y(u0__abc_49347_n2884) );
  AND2X2 AND2X2_716 ( .A(u0__abc_49347_n2885), .B(u0__abc_49347_n2724_bF_buf5), .Y(u0__abc_49347_n2886) );
  AND2X2 AND2X2_717 ( .A(u0_tms2_6_), .B(u0_cs2_bF_buf4), .Y(u0__abc_49347_n2887) );
  AND2X2 AND2X2_718 ( .A(u0__abc_49347_n2888), .B(u0__abc_49347_n2723_bF_buf5), .Y(u0__abc_49347_n2889) );
  AND2X2 AND2X2_719 ( .A(u0_tms1_6_), .B(u0_cs1_bF_buf4), .Y(u0__abc_49347_n2890) );
  AND2X2 AND2X2_72 ( .A(u0__abc_49347_n1100_1), .B(u0_lmr_req3), .Y(u0__abc_49347_n1127) );
  AND2X2 AND2X2_720 ( .A(u0__abc_49347_n1175_bF_buf6), .B(u0__abc_49347_n2893), .Y(u0__abc_49347_n2894) );
  AND2X2 AND2X2_721 ( .A(u0__abc_49347_n2892), .B(u0__abc_49347_n2894), .Y(u0__abc_49347_n2895) );
  AND2X2 AND2X2_722 ( .A(u0__abc_49347_n1176_1_bF_buf6), .B(tms_7_), .Y(u0__abc_49347_n2897) );
  AND2X2 AND2X2_723 ( .A(u0_tms5_7_), .B(u0_cs5_bF_buf3), .Y(u0__abc_49347_n2898) );
  AND2X2 AND2X2_724 ( .A(u0__abc_49347_n2900), .B(u0__abc_49347_n2730_bF_buf4), .Y(u0__abc_49347_n2901) );
  AND2X2 AND2X2_725 ( .A(u0__abc_49347_n2901), .B(u0__abc_49347_n2899), .Y(u0__abc_49347_n2902) );
  AND2X2 AND2X2_726 ( .A(u0__abc_49347_n2903), .B(u0__abc_49347_n2726_bF_buf4), .Y(u0__abc_49347_n2904) );
  AND2X2 AND2X2_727 ( .A(u0_tms4_7_), .B(u0_cs4_bF_buf3), .Y(u0__abc_49347_n2905) );
  AND2X2 AND2X2_728 ( .A(u0__abc_49347_n2906), .B(u0__abc_49347_n2725_bF_buf4), .Y(u0__abc_49347_n2907) );
  AND2X2 AND2X2_729 ( .A(u0_tms3_7_), .B(u0_cs3_bF_buf3), .Y(u0__abc_49347_n2908) );
  AND2X2 AND2X2_73 ( .A(init_req), .B(u0_init_req3), .Y(u0__abc_49347_n1128_1) );
  AND2X2 AND2X2_730 ( .A(u0__abc_49347_n2909), .B(u0__abc_49347_n2724_bF_buf4), .Y(u0__abc_49347_n2910) );
  AND2X2 AND2X2_731 ( .A(u0_tms2_7_), .B(u0_cs2_bF_buf3), .Y(u0__abc_49347_n2911) );
  AND2X2 AND2X2_732 ( .A(u0__abc_49347_n2912), .B(u0__abc_49347_n2723_bF_buf4), .Y(u0__abc_49347_n2913_1) );
  AND2X2 AND2X2_733 ( .A(u0_tms1_7_), .B(u0_cs1_bF_buf3), .Y(u0__abc_49347_n2914) );
  AND2X2 AND2X2_734 ( .A(u0__abc_49347_n1175_bF_buf5), .B(u0__abc_49347_n2917), .Y(u0__abc_49347_n2918) );
  AND2X2 AND2X2_735 ( .A(u0__abc_49347_n2916), .B(u0__abc_49347_n2918), .Y(u0__abc_49347_n2919) );
  AND2X2 AND2X2_736 ( .A(u0__abc_49347_n1176_1_bF_buf5), .B(tms_8_), .Y(u0__abc_49347_n2921) );
  AND2X2 AND2X2_737 ( .A(u0_tms5_8_), .B(u0_cs5_bF_buf2), .Y(u0__abc_49347_n2922) );
  AND2X2 AND2X2_738 ( .A(u0__abc_49347_n2924), .B(u0__abc_49347_n2730_bF_buf3), .Y(u0__abc_49347_n2925) );
  AND2X2 AND2X2_739 ( .A(u0__abc_49347_n2925), .B(u0__abc_49347_n2923), .Y(u0__abc_49347_n2926) );
  AND2X2 AND2X2_74 ( .A(u0__abc_49347_n1105_1), .B(u0__abc_49347_n1129), .Y(u0__abc_49347_n1130_1) );
  AND2X2 AND2X2_740 ( .A(u0__abc_49347_n2927), .B(u0__abc_49347_n2726_bF_buf3), .Y(u0__abc_49347_n2928) );
  AND2X2 AND2X2_741 ( .A(u0_tms4_8_), .B(u0_cs4_bF_buf2), .Y(u0__abc_49347_n2929) );
  AND2X2 AND2X2_742 ( .A(u0__abc_49347_n2930), .B(u0__abc_49347_n2725_bF_buf3), .Y(u0__abc_49347_n2931) );
  AND2X2 AND2X2_743 ( .A(u0_tms3_8_), .B(u0_cs3_bF_buf2), .Y(u0__abc_49347_n2932) );
  AND2X2 AND2X2_744 ( .A(u0__abc_49347_n2933), .B(u0__abc_49347_n2724_bF_buf3), .Y(u0__abc_49347_n2934) );
  AND2X2 AND2X2_745 ( .A(u0_tms2_8_), .B(u0_cs2_bF_buf2), .Y(u0__abc_49347_n2935) );
  AND2X2 AND2X2_746 ( .A(u0__abc_49347_n2936), .B(u0__abc_49347_n2723_bF_buf3), .Y(u0__abc_49347_n2937) );
  AND2X2 AND2X2_747 ( .A(u0_tms1_8_), .B(u0_cs1_bF_buf2), .Y(u0__abc_49347_n2938) );
  AND2X2 AND2X2_748 ( .A(u0__abc_49347_n1175_bF_buf4), .B(u0__abc_49347_n2941), .Y(u0__abc_49347_n2942) );
  AND2X2 AND2X2_749 ( .A(u0__abc_49347_n2940), .B(u0__abc_49347_n2942), .Y(u0__abc_49347_n2943) );
  AND2X2 AND2X2_75 ( .A(u0__abc_49347_n1130_1), .B(u0__abc_49347_n1126_1), .Y(u0__abc_49347_n1131) );
  AND2X2 AND2X2_750 ( .A(u0__abc_49347_n1176_1_bF_buf4), .B(tms_9_), .Y(u0__abc_49347_n2945_1) );
  AND2X2 AND2X2_751 ( .A(u0_tms5_9_), .B(u0_cs5_bF_buf1), .Y(u0__abc_49347_n2946) );
  AND2X2 AND2X2_752 ( .A(u0__abc_49347_n2948), .B(u0__abc_49347_n2730_bF_buf2), .Y(u0__abc_49347_n2949) );
  AND2X2 AND2X2_753 ( .A(u0__abc_49347_n2949), .B(u0__abc_49347_n2947), .Y(u0__abc_49347_n2950) );
  AND2X2 AND2X2_754 ( .A(u0__abc_49347_n2951), .B(u0__abc_49347_n2726_bF_buf2), .Y(u0__abc_49347_n2952) );
  AND2X2 AND2X2_755 ( .A(u0_tms4_9_), .B(u0_cs4_bF_buf1), .Y(u0__abc_49347_n2953) );
  AND2X2 AND2X2_756 ( .A(u0__abc_49347_n2954), .B(u0__abc_49347_n2725_bF_buf2), .Y(u0__abc_49347_n2955) );
  AND2X2 AND2X2_757 ( .A(u0_tms3_9_), .B(u0_cs3_bF_buf1), .Y(u0__abc_49347_n2956) );
  AND2X2 AND2X2_758 ( .A(u0__abc_49347_n2957), .B(u0__abc_49347_n2724_bF_buf2), .Y(u0__abc_49347_n2958) );
  AND2X2 AND2X2_759 ( .A(u0_tms2_9_), .B(u0_cs2_bF_buf1), .Y(u0__abc_49347_n2959) );
  AND2X2 AND2X2_76 ( .A(u0__abc_49347_n1113_1), .B(spec_req_cs_4_bF_buf4), .Y(u0__abc_49347_n1133_1) );
  AND2X2 AND2X2_760 ( .A(u0__abc_49347_n2960), .B(u0__abc_49347_n2723_bF_buf2), .Y(u0__abc_49347_n2961) );
  AND2X2 AND2X2_761 ( .A(u0_tms1_9_), .B(u0_cs1_bF_buf1), .Y(u0__abc_49347_n2962) );
  AND2X2 AND2X2_762 ( .A(u0__abc_49347_n1175_bF_buf3), .B(u0__abc_49347_n2965), .Y(u0__abc_49347_n2966) );
  AND2X2 AND2X2_763 ( .A(u0__abc_49347_n2964), .B(u0__abc_49347_n2966), .Y(u0__abc_49347_n2967) );
  AND2X2 AND2X2_764 ( .A(u0__abc_49347_n1176_1_bF_buf3), .B(tms_10_), .Y(u0__abc_49347_n2969) );
  AND2X2 AND2X2_765 ( .A(u0_tms5_10_), .B(u0_cs5_bF_buf0), .Y(u0__abc_49347_n2970) );
  AND2X2 AND2X2_766 ( .A(u0__abc_49347_n2972), .B(u0__abc_49347_n2730_bF_buf1), .Y(u0__abc_49347_n2973) );
  AND2X2 AND2X2_767 ( .A(u0__abc_49347_n2973), .B(u0__abc_49347_n2971), .Y(u0__abc_49347_n2974) );
  AND2X2 AND2X2_768 ( .A(u0__abc_49347_n2975), .B(u0__abc_49347_n2726_bF_buf1), .Y(u0__abc_49347_n2976) );
  AND2X2 AND2X2_769 ( .A(u0_tms4_10_), .B(u0_cs4_bF_buf0), .Y(u0__abc_49347_n2977_1) );
  AND2X2 AND2X2_77 ( .A(u0__abc_49347_n1126_1), .B(u0__abc_49347_n1104), .Y(u0__abc_49347_n1135_1) );
  AND2X2 AND2X2_770 ( .A(u0__abc_49347_n2978), .B(u0__abc_49347_n2725_bF_buf1), .Y(u0__abc_49347_n2979) );
  AND2X2 AND2X2_771 ( .A(u0_tms3_10_), .B(u0_cs3_bF_buf0), .Y(u0__abc_49347_n2980) );
  AND2X2 AND2X2_772 ( .A(u0__abc_49347_n2981), .B(u0__abc_49347_n2724_bF_buf1), .Y(u0__abc_49347_n2982) );
  AND2X2 AND2X2_773 ( .A(u0_tms2_10_), .B(u0_cs2_bF_buf0), .Y(u0__abc_49347_n2983) );
  AND2X2 AND2X2_774 ( .A(u0__abc_49347_n2984), .B(u0__abc_49347_n2723_bF_buf1), .Y(u0__abc_49347_n2985) );
  AND2X2 AND2X2_775 ( .A(u0_tms1_10_), .B(u0_cs1_bF_buf0), .Y(u0__abc_49347_n2986) );
  AND2X2 AND2X2_776 ( .A(u0__abc_49347_n1175_bF_buf2), .B(u0__abc_49347_n2989), .Y(u0__abc_49347_n2990) );
  AND2X2 AND2X2_777 ( .A(u0__abc_49347_n2988), .B(u0__abc_49347_n2990), .Y(u0__abc_49347_n2991) );
  AND2X2 AND2X2_778 ( .A(u0__abc_49347_n1176_1_bF_buf2), .B(tms_11_), .Y(u0__abc_49347_n2993) );
  AND2X2 AND2X2_779 ( .A(u0_tms5_11_), .B(u0_cs5_bF_buf5), .Y(u0__abc_49347_n2994) );
  AND2X2 AND2X2_78 ( .A(u0__abc_49347_n1135_1), .B(u0__abc_49347_n1134_1), .Y(u0__abc_49347_n1136) );
  AND2X2 AND2X2_780 ( .A(u0__abc_49347_n2996), .B(u0__abc_49347_n2730_bF_buf0), .Y(u0__abc_49347_n2997) );
  AND2X2 AND2X2_781 ( .A(u0__abc_49347_n2997), .B(u0__abc_49347_n2995), .Y(u0__abc_49347_n2998) );
  AND2X2 AND2X2_782 ( .A(u0__abc_49347_n2999), .B(u0__abc_49347_n2726_bF_buf0), .Y(u0__abc_49347_n3000) );
  AND2X2 AND2X2_783 ( .A(u0_tms4_11_), .B(u0_cs4_bF_buf5), .Y(u0__abc_49347_n3001) );
  AND2X2 AND2X2_784 ( .A(u0__abc_49347_n3002), .B(u0__abc_49347_n2725_bF_buf0), .Y(u0__abc_49347_n3003) );
  AND2X2 AND2X2_785 ( .A(u0_tms3_11_), .B(u0_cs3_bF_buf5), .Y(u0__abc_49347_n3004) );
  AND2X2 AND2X2_786 ( .A(u0__abc_49347_n3005), .B(u0__abc_49347_n2724_bF_buf0), .Y(u0__abc_49347_n3006) );
  AND2X2 AND2X2_787 ( .A(u0_tms2_11_), .B(u0_cs2_bF_buf5), .Y(u0__abc_49347_n3007) );
  AND2X2 AND2X2_788 ( .A(u0__abc_49347_n3008), .B(u0__abc_49347_n2723_bF_buf0), .Y(u0__abc_49347_n3009_1) );
  AND2X2 AND2X2_789 ( .A(u0_tms1_11_), .B(u0_cs1_bF_buf5), .Y(u0__abc_49347_n3010) );
  AND2X2 AND2X2_79 ( .A(u0__abc_49347_n1100_1), .B(u0_lmr_req4), .Y(u0__abc_49347_n1137_1) );
  AND2X2 AND2X2_790 ( .A(u0__abc_49347_n1175_bF_buf1), .B(u0__abc_49347_n3013), .Y(u0__abc_49347_n3014) );
  AND2X2 AND2X2_791 ( .A(u0__abc_49347_n3012), .B(u0__abc_49347_n3014), .Y(u0__abc_49347_n3015) );
  AND2X2 AND2X2_792 ( .A(u0__abc_49347_n1176_1_bF_buf1), .B(tms_12_), .Y(u0__abc_49347_n3017) );
  AND2X2 AND2X2_793 ( .A(u0_tms5_12_), .B(u0_cs5_bF_buf4), .Y(u0__abc_49347_n3018) );
  AND2X2 AND2X2_794 ( .A(u0__abc_49347_n3020), .B(u0__abc_49347_n2730_bF_buf5), .Y(u0__abc_49347_n3021) );
  AND2X2 AND2X2_795 ( .A(u0__abc_49347_n3021), .B(u0__abc_49347_n3019), .Y(u0__abc_49347_n3022) );
  AND2X2 AND2X2_796 ( .A(u0__abc_49347_n3023), .B(u0__abc_49347_n2726_bF_buf5), .Y(u0__abc_49347_n3024) );
  AND2X2 AND2X2_797 ( .A(u0_tms4_12_), .B(u0_cs4_bF_buf4), .Y(u0__abc_49347_n3025) );
  AND2X2 AND2X2_798 ( .A(u0__abc_49347_n3026), .B(u0__abc_49347_n2725_bF_buf5), .Y(u0__abc_49347_n3027) );
  AND2X2 AND2X2_799 ( .A(u0_tms3_12_), .B(u0_cs3_bF_buf4), .Y(u0__abc_49347_n3028) );
  AND2X2 AND2X2_8 ( .A(_abc_55805_n260), .B(_abc_55805_n261), .Y(_abc_55805_n262) );
  AND2X2 AND2X2_80 ( .A(init_req), .B(u0_init_req4), .Y(u0__abc_49347_n1138) );
  AND2X2 AND2X2_800 ( .A(u0__abc_49347_n3029), .B(u0__abc_49347_n2724_bF_buf5), .Y(u0__abc_49347_n3030) );
  AND2X2 AND2X2_801 ( .A(u0_tms2_12_), .B(u0_cs2_bF_buf4), .Y(u0__abc_49347_n3031) );
  AND2X2 AND2X2_802 ( .A(u0__abc_49347_n3032), .B(u0__abc_49347_n2723_bF_buf5), .Y(u0__abc_49347_n3033) );
  AND2X2 AND2X2_803 ( .A(u0_tms1_12_), .B(u0_cs1_bF_buf4), .Y(u0__abc_49347_n3034) );
  AND2X2 AND2X2_804 ( .A(u0__abc_49347_n1175_bF_buf0), .B(u0__abc_49347_n3037), .Y(u0__abc_49347_n3038) );
  AND2X2 AND2X2_805 ( .A(u0__abc_49347_n3036), .B(u0__abc_49347_n3038), .Y(u0__abc_49347_n3039) );
  AND2X2 AND2X2_806 ( .A(u0__abc_49347_n1176_1_bF_buf0), .B(tms_13_), .Y(u0__abc_49347_n3041_1) );
  AND2X2 AND2X2_807 ( .A(u0_tms5_13_), .B(u0_cs5_bF_buf3), .Y(u0__abc_49347_n3042) );
  AND2X2 AND2X2_808 ( .A(u0__abc_49347_n3044), .B(u0__abc_49347_n2730_bF_buf4), .Y(u0__abc_49347_n3045) );
  AND2X2 AND2X2_809 ( .A(u0__abc_49347_n3045), .B(u0__abc_49347_n3043), .Y(u0__abc_49347_n3046) );
  AND2X2 AND2X2_81 ( .A(u0__abc_49347_n1139_1), .B(u0_sreq_cs_le), .Y(u0__abc_49347_n1140) );
  AND2X2 AND2X2_810 ( .A(u0__abc_49347_n3047), .B(u0__abc_49347_n2726_bF_buf4), .Y(u0__abc_49347_n3048) );
  AND2X2 AND2X2_811 ( .A(u0_tms4_13_), .B(u0_cs4_bF_buf3), .Y(u0__abc_49347_n3049) );
  AND2X2 AND2X2_812 ( .A(u0__abc_49347_n3050), .B(u0__abc_49347_n2725_bF_buf4), .Y(u0__abc_49347_n3051) );
  AND2X2 AND2X2_813 ( .A(u0_tms3_13_), .B(u0_cs3_bF_buf3), .Y(u0__abc_49347_n3052) );
  AND2X2 AND2X2_814 ( .A(u0__abc_49347_n3053), .B(u0__abc_49347_n2724_bF_buf4), .Y(u0__abc_49347_n3054) );
  AND2X2 AND2X2_815 ( .A(u0_tms2_13_), .B(u0_cs2_bF_buf3), .Y(u0__abc_49347_n3055) );
  AND2X2 AND2X2_816 ( .A(u0__abc_49347_n3056), .B(u0__abc_49347_n2723_bF_buf4), .Y(u0__abc_49347_n3057) );
  AND2X2 AND2X2_817 ( .A(u0_tms1_13_), .B(u0_cs1_bF_buf3), .Y(u0__abc_49347_n3058) );
  AND2X2 AND2X2_818 ( .A(u0__abc_49347_n1175_bF_buf6), .B(u0__abc_49347_n3061), .Y(u0__abc_49347_n3062) );
  AND2X2 AND2X2_819 ( .A(u0__abc_49347_n3060), .B(u0__abc_49347_n3062), .Y(u0__abc_49347_n3063) );
  AND2X2 AND2X2_82 ( .A(u0__abc_49347_n1136), .B(u0__abc_49347_n1140), .Y(u0__abc_49347_n1141_1) );
  AND2X2 AND2X2_820 ( .A(u0__abc_49347_n1176_1_bF_buf6), .B(tms_14_), .Y(u0__abc_49347_n3065) );
  AND2X2 AND2X2_821 ( .A(u0_tms5_14_), .B(u0_cs5_bF_buf2), .Y(u0__abc_49347_n3066) );
  AND2X2 AND2X2_822 ( .A(u0__abc_49347_n3068), .B(u0__abc_49347_n2730_bF_buf3), .Y(u0__abc_49347_n3069) );
  AND2X2 AND2X2_823 ( .A(u0__abc_49347_n3069), .B(u0__abc_49347_n3067), .Y(u0__abc_49347_n3070) );
  AND2X2 AND2X2_824 ( .A(u0__abc_49347_n3071), .B(u0__abc_49347_n2726_bF_buf3), .Y(u0__abc_49347_n3072) );
  AND2X2 AND2X2_825 ( .A(u0_tms4_14_), .B(u0_cs4_bF_buf2), .Y(u0__abc_49347_n3073_1) );
  AND2X2 AND2X2_826 ( .A(u0__abc_49347_n3074), .B(u0__abc_49347_n2725_bF_buf3), .Y(u0__abc_49347_n3075) );
  AND2X2 AND2X2_827 ( .A(u0_tms3_14_), .B(u0_cs3_bF_buf2), .Y(u0__abc_49347_n3076) );
  AND2X2 AND2X2_828 ( .A(u0__abc_49347_n3077), .B(u0__abc_49347_n2724_bF_buf3), .Y(u0__abc_49347_n3078) );
  AND2X2 AND2X2_829 ( .A(u0_tms2_14_), .B(u0_cs2_bF_buf2), .Y(u0__abc_49347_n3079) );
  AND2X2 AND2X2_83 ( .A(u0__abc_49347_n1113_1), .B(spec_req_cs_5_bF_buf4), .Y(u0__abc_49347_n1143_1) );
  AND2X2 AND2X2_830 ( .A(u0__abc_49347_n3080), .B(u0__abc_49347_n2723_bF_buf3), .Y(u0__abc_49347_n3081) );
  AND2X2 AND2X2_831 ( .A(u0_tms1_14_), .B(u0_cs1_bF_buf2), .Y(u0__abc_49347_n3082) );
  AND2X2 AND2X2_832 ( .A(u0__abc_49347_n1175_bF_buf5), .B(u0__abc_49347_n3085), .Y(u0__abc_49347_n3086) );
  AND2X2 AND2X2_833 ( .A(u0__abc_49347_n3084), .B(u0__abc_49347_n3086), .Y(u0__abc_49347_n3087) );
  AND2X2 AND2X2_834 ( .A(u0__abc_49347_n1176_1_bF_buf5), .B(tms_15_), .Y(u0__abc_49347_n3089) );
  AND2X2 AND2X2_835 ( .A(u0_tms5_15_), .B(u0_cs5_bF_buf1), .Y(u0__abc_49347_n3090) );
  AND2X2 AND2X2_836 ( .A(u0__abc_49347_n3092), .B(u0__abc_49347_n2730_bF_buf2), .Y(u0__abc_49347_n3093) );
  AND2X2 AND2X2_837 ( .A(u0__abc_49347_n3093), .B(u0__abc_49347_n3091), .Y(u0__abc_49347_n3094) );
  AND2X2 AND2X2_838 ( .A(u0__abc_49347_n3095), .B(u0__abc_49347_n2726_bF_buf2), .Y(u0__abc_49347_n3096) );
  AND2X2 AND2X2_839 ( .A(u0_tms4_15_), .B(u0_cs4_bF_buf1), .Y(u0__abc_49347_n3097) );
  AND2X2 AND2X2_84 ( .A(u0__abc_49347_n1100_1), .B(u0_lmr_req5), .Y(u0__abc_49347_n1144) );
  AND2X2 AND2X2_840 ( .A(u0__abc_49347_n3098), .B(u0__abc_49347_n2725_bF_buf2), .Y(u0__abc_49347_n3099) );
  AND2X2 AND2X2_841 ( .A(u0_tms3_15_), .B(u0_cs3_bF_buf1), .Y(u0__abc_49347_n3100) );
  AND2X2 AND2X2_842 ( .A(u0__abc_49347_n3101), .B(u0__abc_49347_n2724_bF_buf2), .Y(u0__abc_49347_n3102) );
  AND2X2 AND2X2_843 ( .A(u0_tms2_15_), .B(u0_cs2_bF_buf1), .Y(u0__abc_49347_n3103) );
  AND2X2 AND2X2_844 ( .A(u0__abc_49347_n3104), .B(u0__abc_49347_n2723_bF_buf2), .Y(u0__abc_49347_n3105_1) );
  AND2X2 AND2X2_845 ( .A(u0_tms1_15_), .B(u0_cs1_bF_buf1), .Y(u0__abc_49347_n3106_1) );
  AND2X2 AND2X2_846 ( .A(u0__abc_49347_n1175_bF_buf4), .B(u0__abc_49347_n3109), .Y(u0__abc_49347_n3110_1) );
  AND2X2 AND2X2_847 ( .A(u0__abc_49347_n3108_1), .B(u0__abc_49347_n3110_1), .Y(u0__abc_49347_n3111) );
  AND2X2 AND2X2_848 ( .A(u0__abc_49347_n1176_1_bF_buf4), .B(tms_16_), .Y(u0__abc_49347_n3113) );
  AND2X2 AND2X2_849 ( .A(u0_tms5_16_), .B(u0_cs5_bF_buf0), .Y(u0__abc_49347_n3114) );
  AND2X2 AND2X2_85 ( .A(init_req), .B(u0_init_req5), .Y(u0__abc_49347_n1145_1) );
  AND2X2 AND2X2_850 ( .A(u0__abc_49347_n3116_1), .B(u0__abc_49347_n2730_bF_buf1), .Y(u0__abc_49347_n3117) );
  AND2X2 AND2X2_851 ( .A(u0__abc_49347_n3117), .B(u0__abc_49347_n3115_1), .Y(u0__abc_49347_n3118) );
  AND2X2 AND2X2_852 ( .A(u0__abc_49347_n3119), .B(u0__abc_49347_n2726_bF_buf1), .Y(u0__abc_49347_n3120_1) );
  AND2X2 AND2X2_853 ( .A(u0_tms4_16_), .B(u0_cs4_bF_buf0), .Y(u0__abc_49347_n3121) );
  AND2X2 AND2X2_854 ( .A(u0__abc_49347_n3122), .B(u0__abc_49347_n2725_bF_buf1), .Y(u0__abc_49347_n3123_1) );
  AND2X2 AND2X2_855 ( .A(u0_tms3_16_), .B(u0_cs3_bF_buf0), .Y(u0__abc_49347_n3124) );
  AND2X2 AND2X2_856 ( .A(u0__abc_49347_n3125), .B(u0__abc_49347_n2724_bF_buf1), .Y(u0__abc_49347_n3126_1) );
  AND2X2 AND2X2_857 ( .A(u0_tms2_16_), .B(u0_cs2_bF_buf0), .Y(u0__abc_49347_n3127) );
  AND2X2 AND2X2_858 ( .A(u0__abc_49347_n3128), .B(u0__abc_49347_n2723_bF_buf1), .Y(u0__abc_49347_n3129_1) );
  AND2X2 AND2X2_859 ( .A(u0_tms1_16_), .B(u0_cs1_bF_buf0), .Y(u0__abc_49347_n3130) );
  AND2X2 AND2X2_86 ( .A(u0__abc_49347_n1105_1), .B(u0__abc_49347_n1146), .Y(u0__abc_49347_n1147_1) );
  AND2X2 AND2X2_860 ( .A(u0__abc_49347_n1175_bF_buf3), .B(u0__abc_49347_n3133), .Y(u0__abc_49347_n3134) );
  AND2X2 AND2X2_861 ( .A(u0__abc_49347_n3132_1), .B(u0__abc_49347_n3134), .Y(u0__abc_49347_n3135_1) );
  AND2X2 AND2X2_862 ( .A(u0__abc_49347_n1176_1_bF_buf3), .B(tms_17_), .Y(u0__abc_49347_n3137) );
  AND2X2 AND2X2_863 ( .A(u0_tms5_17_), .B(u0_cs5_bF_buf5), .Y(u0__abc_49347_n3138_1) );
  AND2X2 AND2X2_864 ( .A(u0__abc_49347_n3140), .B(u0__abc_49347_n2730_bF_buf0), .Y(u0__abc_49347_n3141_1) );
  AND2X2 AND2X2_865 ( .A(u0__abc_49347_n3141_1), .B(u0__abc_49347_n3139), .Y(u0__abc_49347_n3142) );
  AND2X2 AND2X2_866 ( .A(u0__abc_49347_n3143), .B(u0__abc_49347_n2726_bF_buf0), .Y(u0__abc_49347_n3144_1) );
  AND2X2 AND2X2_867 ( .A(u0_tms4_17_), .B(u0_cs4_bF_buf5), .Y(u0__abc_49347_n3145_1) );
  AND2X2 AND2X2_868 ( .A(u0__abc_49347_n3146), .B(u0__abc_49347_n2725_bF_buf0), .Y(u0__abc_49347_n3147_1) );
  AND2X2 AND2X2_869 ( .A(u0_tms3_17_), .B(u0_cs3_bF_buf5), .Y(u0__abc_49347_n3148) );
  AND2X2 AND2X2_87 ( .A(u0__abc_49347_n1134_1), .B(u0__abc_49347_n1148), .Y(u0__abc_49347_n1149_1) );
  AND2X2 AND2X2_870 ( .A(u0__abc_49347_n3149_1), .B(u0__abc_49347_n2724_bF_buf0), .Y(u0__abc_49347_n3150) );
  AND2X2 AND2X2_871 ( .A(u0_tms2_17_), .B(u0_cs2_bF_buf5), .Y(u0__abc_49347_n3151_1) );
  AND2X2 AND2X2_872 ( .A(u0__abc_49347_n3152), .B(u0__abc_49347_n2723_bF_buf0), .Y(u0__abc_49347_n3153_1) );
  AND2X2 AND2X2_873 ( .A(u0_tms1_17_), .B(u0_cs1_bF_buf5), .Y(u0__abc_49347_n3154) );
  AND2X2 AND2X2_874 ( .A(u0__abc_49347_n1175_bF_buf2), .B(u0__abc_49347_n3157), .Y(u0__abc_49347_n3158) );
  AND2X2 AND2X2_875 ( .A(u0__abc_49347_n3156_1), .B(u0__abc_49347_n3158), .Y(u0__abc_49347_n3159) );
  AND2X2 AND2X2_876 ( .A(u0__abc_49347_n1176_1_bF_buf2), .B(tms_18_), .Y(u0__abc_49347_n3161) );
  AND2X2 AND2X2_877 ( .A(u0_tms5_18_), .B(u0_cs5_bF_buf4), .Y(u0__abc_49347_n3162) );
  AND2X2 AND2X2_878 ( .A(u0__abc_49347_n3164), .B(u0__abc_49347_n2730_bF_buf5), .Y(u0__abc_49347_n3165) );
  AND2X2 AND2X2_879 ( .A(u0__abc_49347_n3165), .B(u0__abc_49347_n3163_1), .Y(u0__abc_49347_n3166) );
  AND2X2 AND2X2_88 ( .A(u0__abc_49347_n1126_1), .B(u0__abc_49347_n1149_1), .Y(u0__abc_49347_n1150_1) );
  AND2X2 AND2X2_880 ( .A(u0__abc_49347_n3167), .B(u0__abc_49347_n2726_bF_buf5), .Y(u0__abc_49347_n3168) );
  AND2X2 AND2X2_881 ( .A(u0_tms4_18_), .B(u0_cs4_bF_buf4), .Y(u0__abc_49347_n3169) );
  AND2X2 AND2X2_882 ( .A(u0__abc_49347_n3170_1), .B(u0__abc_49347_n2725_bF_buf5), .Y(u0__abc_49347_n3171_1) );
  AND2X2 AND2X2_883 ( .A(u0_tms3_18_), .B(u0_cs3_bF_buf4), .Y(u0__abc_49347_n3172_1) );
  AND2X2 AND2X2_884 ( .A(u0__abc_49347_n3173_1), .B(u0__abc_49347_n2724_bF_buf5), .Y(u0__abc_49347_n3174_1) );
  AND2X2 AND2X2_885 ( .A(u0_tms2_18_), .B(u0_cs2_bF_buf4), .Y(u0__abc_49347_n3175_1) );
  AND2X2 AND2X2_886 ( .A(u0__abc_49347_n3176_1), .B(u0__abc_49347_n2723_bF_buf5), .Y(u0__abc_49347_n3177_1) );
  AND2X2 AND2X2_887 ( .A(u0_tms1_18_), .B(u0_cs1_bF_buf4), .Y(u0__abc_49347_n3178_1) );
  AND2X2 AND2X2_888 ( .A(u0__abc_49347_n1175_bF_buf1), .B(u0__abc_49347_n3181_1), .Y(u0__abc_49347_n3182_1) );
  AND2X2 AND2X2_889 ( .A(u0__abc_49347_n3180_1), .B(u0__abc_49347_n3182_1), .Y(u0__abc_49347_n3183_1) );
  AND2X2 AND2X2_89 ( .A(u0__abc_49347_n1150_1), .B(u0__abc_49347_n1147_1), .Y(u0__abc_49347_n1151_1) );
  AND2X2 AND2X2_890 ( .A(u0__abc_49347_n1176_1_bF_buf1), .B(tms_19_), .Y(u0__abc_49347_n3185_1) );
  AND2X2 AND2X2_891 ( .A(u0_tms5_19_), .B(u0_cs5_bF_buf3), .Y(u0__abc_49347_n3186_1) );
  AND2X2 AND2X2_892 ( .A(u0__abc_49347_n3188_1), .B(u0__abc_49347_n2730_bF_buf4), .Y(u0__abc_49347_n3189) );
  AND2X2 AND2X2_893 ( .A(u0__abc_49347_n3189), .B(u0__abc_49347_n3187_1), .Y(u0__abc_49347_n3190) );
  AND2X2 AND2X2_894 ( .A(u0__abc_49347_n3191), .B(u0__abc_49347_n2726_bF_buf4), .Y(u0__abc_49347_n3192) );
  AND2X2 AND2X2_895 ( .A(u0_tms4_19_), .B(u0_cs4_bF_buf3), .Y(u0__abc_49347_n3193) );
  AND2X2 AND2X2_896 ( .A(u0__abc_49347_n3194), .B(u0__abc_49347_n2725_bF_buf4), .Y(u0__abc_49347_n3195) );
  AND2X2 AND2X2_897 ( .A(u0_tms3_19_), .B(u0_cs3_bF_buf3), .Y(u0__abc_49347_n3196) );
  AND2X2 AND2X2_898 ( .A(u0__abc_49347_n3197), .B(u0__abc_49347_n2724_bF_buf4), .Y(u0__abc_49347_n3198) );
  AND2X2 AND2X2_899 ( .A(u0_tms2_19_), .B(u0_cs2_bF_buf3), .Y(u0__abc_49347_n3199) );
  AND2X2 AND2X2_9 ( .A(_abc_55805_n263), .B(_abc_55805_n264), .Y(obct_cs_3_) );
  AND2X2 AND2X2_90 ( .A(u0__abc_49347_n1153), .B(u0_sreq_cs_le), .Y(u0__abc_49347_n1154_1) );
  AND2X2 AND2X2_900 ( .A(u0__abc_49347_n3200), .B(u0__abc_49347_n2723_bF_buf4), .Y(u0__abc_49347_n3201) );
  AND2X2 AND2X2_901 ( .A(u0_tms1_19_), .B(u0_cs1_bF_buf3), .Y(u0__abc_49347_n3202) );
  AND2X2 AND2X2_902 ( .A(u0__abc_49347_n1175_bF_buf0), .B(u0__abc_49347_n3205), .Y(u0__abc_49347_n3206) );
  AND2X2 AND2X2_903 ( .A(u0__abc_49347_n3204), .B(u0__abc_49347_n3206), .Y(u0__abc_49347_n3207) );
  AND2X2 AND2X2_904 ( .A(u0__abc_49347_n1176_1_bF_buf0), .B(tms_20_), .Y(u0__abc_49347_n3209) );
  AND2X2 AND2X2_905 ( .A(u0_tms5_20_), .B(u0_cs5_bF_buf2), .Y(u0__abc_49347_n3210) );
  AND2X2 AND2X2_906 ( .A(u0__abc_49347_n3212), .B(u0__abc_49347_n2730_bF_buf3), .Y(u0__abc_49347_n3213) );
  AND2X2 AND2X2_907 ( .A(u0__abc_49347_n3213), .B(u0__abc_49347_n3211), .Y(u0__abc_49347_n3214) );
  AND2X2 AND2X2_908 ( .A(u0__abc_49347_n3215), .B(u0__abc_49347_n2726_bF_buf3), .Y(u0__abc_49347_n3216) );
  AND2X2 AND2X2_909 ( .A(u0_tms4_20_), .B(u0_cs4_bF_buf2), .Y(u0__abc_49347_n3217) );
  AND2X2 AND2X2_91 ( .A(u0__abc_49347_n1100_1), .B(1'b0), .Y(u0__abc_49347_n1155) );
  AND2X2 AND2X2_910 ( .A(u0__abc_49347_n3218), .B(u0__abc_49347_n2725_bF_buf3), .Y(u0__abc_49347_n3219) );
  AND2X2 AND2X2_911 ( .A(u0_tms3_20_), .B(u0_cs3_bF_buf2), .Y(u0__abc_49347_n3220) );
  AND2X2 AND2X2_912 ( .A(u0__abc_49347_n3221), .B(u0__abc_49347_n2724_bF_buf3), .Y(u0__abc_49347_n3222) );
  AND2X2 AND2X2_913 ( .A(u0_tms2_20_), .B(u0_cs2_bF_buf2), .Y(u0__abc_49347_n3223) );
  AND2X2 AND2X2_914 ( .A(u0__abc_49347_n3224), .B(u0__abc_49347_n2723_bF_buf3), .Y(u0__abc_49347_n3225) );
  AND2X2 AND2X2_915 ( .A(u0_tms1_20_), .B(u0_cs1_bF_buf2), .Y(u0__abc_49347_n3226) );
  AND2X2 AND2X2_916 ( .A(u0__abc_49347_n1175_bF_buf6), .B(u0__abc_49347_n3229), .Y(u0__abc_49347_n3230) );
  AND2X2 AND2X2_917 ( .A(u0__abc_49347_n3228), .B(u0__abc_49347_n3230), .Y(u0__abc_49347_n3231) );
  AND2X2 AND2X2_918 ( .A(u0__abc_49347_n1176_1_bF_buf6), .B(tms_21_), .Y(u0__abc_49347_n3233) );
  AND2X2 AND2X2_919 ( .A(u0_tms5_21_), .B(u0_cs5_bF_buf1), .Y(u0__abc_49347_n3234) );
  AND2X2 AND2X2_92 ( .A(init_req), .B(1'b0), .Y(u0__abc_49347_n1156_1) );
  AND2X2 AND2X2_920 ( .A(u0__abc_49347_n3236), .B(u0__abc_49347_n2730_bF_buf2), .Y(u0__abc_49347_n3237) );
  AND2X2 AND2X2_921 ( .A(u0__abc_49347_n3237), .B(u0__abc_49347_n3235), .Y(u0__abc_49347_n3238) );
  AND2X2 AND2X2_922 ( .A(u0__abc_49347_n3239), .B(u0__abc_49347_n2726_bF_buf2), .Y(u0__abc_49347_n3240) );
  AND2X2 AND2X2_923 ( .A(u0_tms4_21_), .B(u0_cs4_bF_buf1), .Y(u0__abc_49347_n3241) );
  AND2X2 AND2X2_924 ( .A(u0__abc_49347_n3242), .B(u0__abc_49347_n2725_bF_buf2), .Y(u0__abc_49347_n3243) );
  AND2X2 AND2X2_925 ( .A(u0_tms3_21_), .B(u0_cs3_bF_buf1), .Y(u0__abc_49347_n3244) );
  AND2X2 AND2X2_926 ( .A(u0__abc_49347_n3245), .B(u0__abc_49347_n2724_bF_buf2), .Y(u0__abc_49347_n3246) );
  AND2X2 AND2X2_927 ( .A(u0_tms2_21_), .B(u0_cs2_bF_buf1), .Y(u0__abc_49347_n3247) );
  AND2X2 AND2X2_928 ( .A(u0__abc_49347_n3248), .B(u0__abc_49347_n2723_bF_buf2), .Y(u0__abc_49347_n3249) );
  AND2X2 AND2X2_929 ( .A(u0_tms1_21_), .B(u0_cs1_bF_buf1), .Y(u0__abc_49347_n3250) );
  AND2X2 AND2X2_93 ( .A(u0__abc_49347_n1148), .B(u0__abc_49347_n1157), .Y(u0__abc_49347_n1158_1) );
  AND2X2 AND2X2_930 ( .A(u0__abc_49347_n1175_bF_buf5), .B(u0__abc_49347_n3253), .Y(u0__abc_49347_n3254) );
  AND2X2 AND2X2_931 ( .A(u0__abc_49347_n3252), .B(u0__abc_49347_n3254), .Y(u0__abc_49347_n3255) );
  AND2X2 AND2X2_932 ( .A(u0__abc_49347_n1176_1_bF_buf5), .B(tms_22_), .Y(u0__abc_49347_n3257) );
  AND2X2 AND2X2_933 ( .A(u0_tms5_22_), .B(u0_cs5_bF_buf0), .Y(u0__abc_49347_n3258) );
  AND2X2 AND2X2_934 ( .A(u0__abc_49347_n3260), .B(u0__abc_49347_n2730_bF_buf1), .Y(u0__abc_49347_n3261) );
  AND2X2 AND2X2_935 ( .A(u0__abc_49347_n3261), .B(u0__abc_49347_n3259), .Y(u0__abc_49347_n3262) );
  AND2X2 AND2X2_936 ( .A(u0__abc_49347_n3263), .B(u0__abc_49347_n2726_bF_buf1), .Y(u0__abc_49347_n3264) );
  AND2X2 AND2X2_937 ( .A(u0_tms4_22_), .B(u0_cs4_bF_buf0), .Y(u0__abc_49347_n3265) );
  AND2X2 AND2X2_938 ( .A(u0__abc_49347_n3266), .B(u0__abc_49347_n2725_bF_buf1), .Y(u0__abc_49347_n3267) );
  AND2X2 AND2X2_939 ( .A(u0_tms3_22_), .B(u0_cs3_bF_buf0), .Y(u0__abc_49347_n3268) );
  AND2X2 AND2X2_94 ( .A(u0__abc_49347_n1158_1), .B(u0__abc_49347_n1154_1), .Y(u0__abc_49347_n1159) );
  AND2X2 AND2X2_940 ( .A(u0__abc_49347_n3269), .B(u0__abc_49347_n2724_bF_buf1), .Y(u0__abc_49347_n3270) );
  AND2X2 AND2X2_941 ( .A(u0_tms2_22_), .B(u0_cs2_bF_buf0), .Y(u0__abc_49347_n3271) );
  AND2X2 AND2X2_942 ( .A(u0__abc_49347_n3272), .B(u0__abc_49347_n2723_bF_buf1), .Y(u0__abc_49347_n3273) );
  AND2X2 AND2X2_943 ( .A(u0_tms1_22_), .B(u0_cs1_bF_buf0), .Y(u0__abc_49347_n3274) );
  AND2X2 AND2X2_944 ( .A(u0__abc_49347_n1175_bF_buf4), .B(u0__abc_49347_n3277), .Y(u0__abc_49347_n3278) );
  AND2X2 AND2X2_945 ( .A(u0__abc_49347_n3276), .B(u0__abc_49347_n3278), .Y(u0__abc_49347_n3279) );
  AND2X2 AND2X2_946 ( .A(u0__abc_49347_n1176_1_bF_buf4), .B(tms_23_), .Y(u0__abc_49347_n3281) );
  AND2X2 AND2X2_947 ( .A(u0_tms5_23_), .B(u0_cs5_bF_buf5), .Y(u0__abc_49347_n3282) );
  AND2X2 AND2X2_948 ( .A(u0__abc_49347_n3284), .B(u0__abc_49347_n2730_bF_buf0), .Y(u0__abc_49347_n3285) );
  AND2X2 AND2X2_949 ( .A(u0__abc_49347_n3285), .B(u0__abc_49347_n3283), .Y(u0__abc_49347_n3286) );
  AND2X2 AND2X2_95 ( .A(u0__abc_49347_n1136), .B(u0__abc_49347_n1159), .Y(u0__abc_49347_n1160_1) );
  AND2X2 AND2X2_950 ( .A(u0__abc_49347_n3287), .B(u0__abc_49347_n2726_bF_buf0), .Y(u0__abc_49347_n3288) );
  AND2X2 AND2X2_951 ( .A(u0_tms4_23_), .B(u0_cs4_bF_buf5), .Y(u0__abc_49347_n3289) );
  AND2X2 AND2X2_952 ( .A(u0__abc_49347_n3290), .B(u0__abc_49347_n2725_bF_buf0), .Y(u0__abc_49347_n3291) );
  AND2X2 AND2X2_953 ( .A(u0_tms3_23_), .B(u0_cs3_bF_buf5), .Y(u0__abc_49347_n3292) );
  AND2X2 AND2X2_954 ( .A(u0__abc_49347_n3293), .B(u0__abc_49347_n2724_bF_buf0), .Y(u0__abc_49347_n3294) );
  AND2X2 AND2X2_955 ( .A(u0_tms2_23_), .B(u0_cs2_bF_buf5), .Y(u0__abc_49347_n3295) );
  AND2X2 AND2X2_956 ( .A(u0__abc_49347_n3296), .B(u0__abc_49347_n2723_bF_buf0), .Y(u0__abc_49347_n3297) );
  AND2X2 AND2X2_957 ( .A(u0_tms1_23_), .B(u0_cs1_bF_buf5), .Y(u0__abc_49347_n3298) );
  AND2X2 AND2X2_958 ( .A(u0__abc_49347_n1175_bF_buf3), .B(u0__abc_49347_n3301), .Y(u0__abc_49347_n3302) );
  AND2X2 AND2X2_959 ( .A(u0__abc_49347_n3300), .B(u0__abc_49347_n3302), .Y(u0__abc_49347_n3303) );
  AND2X2 AND2X2_96 ( .A(u0__abc_49347_n1113_1), .B(spec_req_cs_6_bF_buf4), .Y(u0__abc_49347_n1161) );
  AND2X2 AND2X2_960 ( .A(u0__abc_49347_n1176_1_bF_buf3), .B(tms_24_), .Y(u0__abc_49347_n3305) );
  AND2X2 AND2X2_961 ( .A(u0_tms5_24_), .B(u0_cs5_bF_buf4), .Y(u0__abc_49347_n3306) );
  AND2X2 AND2X2_962 ( .A(u0__abc_49347_n3308), .B(u0__abc_49347_n2730_bF_buf5), .Y(u0__abc_49347_n3309) );
  AND2X2 AND2X2_963 ( .A(u0__abc_49347_n3309), .B(u0__abc_49347_n3307), .Y(u0__abc_49347_n3310) );
  AND2X2 AND2X2_964 ( .A(u0__abc_49347_n3311), .B(u0__abc_49347_n2726_bF_buf5), .Y(u0__abc_49347_n3312) );
  AND2X2 AND2X2_965 ( .A(u0_tms4_24_), .B(u0_cs4_bF_buf4), .Y(u0__abc_49347_n3313) );
  AND2X2 AND2X2_966 ( .A(u0__abc_49347_n3314), .B(u0__abc_49347_n2725_bF_buf5), .Y(u0__abc_49347_n3315) );
  AND2X2 AND2X2_967 ( .A(u0_tms3_24_), .B(u0_cs3_bF_buf4), .Y(u0__abc_49347_n3316) );
  AND2X2 AND2X2_968 ( .A(u0__abc_49347_n3317), .B(u0__abc_49347_n2724_bF_buf5), .Y(u0__abc_49347_n3318) );
  AND2X2 AND2X2_969 ( .A(u0_tms2_24_), .B(u0_cs2_bF_buf4), .Y(u0__abc_49347_n3319) );
  AND2X2 AND2X2_97 ( .A(u0__abc_49347_n1113_1), .B(spec_req_cs_7_), .Y(u0__abc_49347_n1163) );
  AND2X2 AND2X2_970 ( .A(u0__abc_49347_n3320), .B(u0__abc_49347_n2723_bF_buf5), .Y(u0__abc_49347_n3321) );
  AND2X2 AND2X2_971 ( .A(u0_tms1_24_), .B(u0_cs1_bF_buf4), .Y(u0__abc_49347_n3322) );
  AND2X2 AND2X2_972 ( .A(u0__abc_49347_n1175_bF_buf2), .B(u0__abc_49347_n3325), .Y(u0__abc_49347_n3326) );
  AND2X2 AND2X2_973 ( .A(u0__abc_49347_n3324), .B(u0__abc_49347_n3326), .Y(u0__abc_49347_n3327) );
  AND2X2 AND2X2_974 ( .A(u0__abc_49347_n1176_1_bF_buf2), .B(tms_25_), .Y(u0__abc_49347_n3329) );
  AND2X2 AND2X2_975 ( .A(u0_tms5_25_), .B(u0_cs5_bF_buf3), .Y(u0__abc_49347_n3330) );
  AND2X2 AND2X2_976 ( .A(u0__abc_49347_n3332), .B(u0__abc_49347_n2730_bF_buf4), .Y(u0__abc_49347_n3333) );
  AND2X2 AND2X2_977 ( .A(u0__abc_49347_n3333), .B(u0__abc_49347_n3331), .Y(u0__abc_49347_n3334) );
  AND2X2 AND2X2_978 ( .A(u0__abc_49347_n3335), .B(u0__abc_49347_n2726_bF_buf4), .Y(u0__abc_49347_n3336) );
  AND2X2 AND2X2_979 ( .A(u0_tms4_25_), .B(u0_cs4_bF_buf3), .Y(u0__abc_49347_n3337) );
  AND2X2 AND2X2_98 ( .A(u0__abc_49347_n1165), .B(u0__abc_49347_n1166_1), .Y(u0__abc_49347_n1167_1) );
  AND2X2 AND2X2_980 ( .A(u0__abc_49347_n3338), .B(u0__abc_49347_n2725_bF_buf4), .Y(u0__abc_49347_n3339) );
  AND2X2 AND2X2_981 ( .A(u0_tms3_25_), .B(u0_cs3_bF_buf3), .Y(u0__abc_49347_n3340) );
  AND2X2 AND2X2_982 ( .A(u0__abc_49347_n3341), .B(u0__abc_49347_n2724_bF_buf4), .Y(u0__abc_49347_n3342) );
  AND2X2 AND2X2_983 ( .A(u0_tms2_25_), .B(u0_cs2_bF_buf3), .Y(u0__abc_49347_n3343) );
  AND2X2 AND2X2_984 ( .A(u0__abc_49347_n3344), .B(u0__abc_49347_n2723_bF_buf4), .Y(u0__abc_49347_n3345) );
  AND2X2 AND2X2_985 ( .A(u0_tms1_25_), .B(u0_cs1_bF_buf3), .Y(u0__abc_49347_n3346) );
  AND2X2 AND2X2_986 ( .A(u0__abc_49347_n1175_bF_buf1), .B(u0__abc_49347_n3349), .Y(u0__abc_49347_n3350) );
  AND2X2 AND2X2_987 ( .A(u0__abc_49347_n3348), .B(u0__abc_49347_n3350), .Y(u0__abc_49347_n3351) );
  AND2X2 AND2X2_988 ( .A(u0__abc_49347_n1176_1_bF_buf1), .B(tms_26_), .Y(u0__abc_49347_n3353) );
  AND2X2 AND2X2_989 ( .A(u0_tms5_26_), .B(u0_cs5_bF_buf2), .Y(u0__abc_49347_n3354) );
  AND2X2 AND2X2_99 ( .A(u0__abc_49347_n1164_1), .B(u0__abc_49347_n1167_1), .Y(u0__abc_49347_n1168_1) );
  AND2X2 AND2X2_990 ( .A(u0__abc_49347_n3356), .B(u0__abc_49347_n2730_bF_buf3), .Y(u0__abc_49347_n3357) );
  AND2X2 AND2X2_991 ( .A(u0__abc_49347_n3357), .B(u0__abc_49347_n3355), .Y(u0__abc_49347_n3358) );
  AND2X2 AND2X2_992 ( .A(u0__abc_49347_n3359), .B(u0__abc_49347_n2726_bF_buf3), .Y(u0__abc_49347_n3360) );
  AND2X2 AND2X2_993 ( .A(u0_tms4_26_), .B(u0_cs4_bF_buf2), .Y(u0__abc_49347_n3361) );
  AND2X2 AND2X2_994 ( .A(u0__abc_49347_n3362), .B(u0__abc_49347_n2725_bF_buf3), .Y(u0__abc_49347_n3363) );
  AND2X2 AND2X2_995 ( .A(u0_tms3_26_), .B(u0_cs3_bF_buf2), .Y(u0__abc_49347_n3364) );
  AND2X2 AND2X2_996 ( .A(u0__abc_49347_n3365), .B(u0__abc_49347_n2724_bF_buf3), .Y(u0__abc_49347_n3366) );
  AND2X2 AND2X2_997 ( .A(u0_tms2_26_), .B(u0_cs2_bF_buf2), .Y(u0__abc_49347_n3367) );
  AND2X2 AND2X2_998 ( .A(u0__abc_49347_n3368), .B(u0__abc_49347_n2723_bF_buf3), .Y(u0__abc_49347_n3369) );
  AND2X2 AND2X2_999 ( .A(u0_tms1_26_), .B(u0_cs1_bF_buf2), .Y(u0__abc_49347_n3370) );
  BUFX2 BUFX2_1 ( .A(clk_i), .Y(clk_i_hier0_bF_buf10) );
  BUFX2 BUFX2_10 ( .A(clk_i), .Y(clk_i_hier0_bF_buf1) );
  BUFX2 BUFX2_100 ( .A(u2_u5__abc_47660_n137), .Y(u2_u5__abc_47660_n137_bF_buf0) );
  BUFX2 BUFX2_1000 ( .A(_auto_iopadmap_cc_313_execute_56255_0_), .Y(\mc_cs_pad_o_[0] ) );
  BUFX2 BUFX2_1001 ( .A(_auto_iopadmap_cc_313_execute_56255_1_), .Y(\mc_cs_pad_o_[1] ) );
  BUFX2 BUFX2_1002 ( .A(_auto_iopadmap_cc_313_execute_56255_2_), .Y(\mc_cs_pad_o_[2] ) );
  BUFX2 BUFX2_1003 ( .A(_auto_iopadmap_cc_313_execute_56255_3_), .Y(\mc_cs_pad_o_[3] ) );
  BUFX2 BUFX2_1004 ( .A(_auto_iopadmap_cc_313_execute_56255_4_), .Y(\mc_cs_pad_o_[4] ) );
  BUFX2 BUFX2_1005 ( .A(_auto_iopadmap_cc_313_execute_56255_5_), .Y(\mc_cs_pad_o_[5] ) );
  BUFX2 BUFX2_1006 ( .A(_auto_iopadmap_cc_313_execute_56255_6_), .Y(\mc_cs_pad_o_[6] ) );
  BUFX2 BUFX2_1007 ( .A(_auto_iopadmap_cc_313_execute_56255_7_), .Y(\mc_cs_pad_o_[7] ) );
  BUFX2 BUFX2_1008 ( .A(_auto_iopadmap_cc_313_execute_56264_0_), .Y(\mc_data_pad_o[0] ) );
  BUFX2 BUFX2_1009 ( .A(_auto_iopadmap_cc_313_execute_56264_1_), .Y(\mc_data_pad_o[1] ) );
  BUFX2 BUFX2_101 ( .A(clk_i_hier0_bF_buf10), .Y(clk_i_bF_buf125) );
  BUFX2 BUFX2_1010 ( .A(_auto_iopadmap_cc_313_execute_56264_2_), .Y(\mc_data_pad_o[2] ) );
  BUFX2 BUFX2_1011 ( .A(_auto_iopadmap_cc_313_execute_56264_3_), .Y(\mc_data_pad_o[3] ) );
  BUFX2 BUFX2_1012 ( .A(_auto_iopadmap_cc_313_execute_56264_4_), .Y(\mc_data_pad_o[4] ) );
  BUFX2 BUFX2_1013 ( .A(_auto_iopadmap_cc_313_execute_56264_5_), .Y(\mc_data_pad_o[5] ) );
  BUFX2 BUFX2_1014 ( .A(_auto_iopadmap_cc_313_execute_56264_6_), .Y(\mc_data_pad_o[6] ) );
  BUFX2 BUFX2_1015 ( .A(_auto_iopadmap_cc_313_execute_56264_7_), .Y(\mc_data_pad_o[7] ) );
  BUFX2 BUFX2_1016 ( .A(_auto_iopadmap_cc_313_execute_56264_8_), .Y(\mc_data_pad_o[8] ) );
  BUFX2 BUFX2_1017 ( .A(_auto_iopadmap_cc_313_execute_56264_9_), .Y(\mc_data_pad_o[9] ) );
  BUFX2 BUFX2_1018 ( .A(_auto_iopadmap_cc_313_execute_56264_10_), .Y(\mc_data_pad_o[10] ) );
  BUFX2 BUFX2_1019 ( .A(_auto_iopadmap_cc_313_execute_56264_11_), .Y(\mc_data_pad_o[11] ) );
  BUFX2 BUFX2_102 ( .A(clk_i_hier0_bF_buf9), .Y(clk_i_bF_buf124) );
  BUFX2 BUFX2_1020 ( .A(_auto_iopadmap_cc_313_execute_56264_12_), .Y(\mc_data_pad_o[12] ) );
  BUFX2 BUFX2_1021 ( .A(_auto_iopadmap_cc_313_execute_56264_13_), .Y(\mc_data_pad_o[13] ) );
  BUFX2 BUFX2_1022 ( .A(_auto_iopadmap_cc_313_execute_56264_14_), .Y(\mc_data_pad_o[14] ) );
  BUFX2 BUFX2_1023 ( .A(_auto_iopadmap_cc_313_execute_56264_15_), .Y(\mc_data_pad_o[15] ) );
  BUFX2 BUFX2_1024 ( .A(_auto_iopadmap_cc_313_execute_56264_16_), .Y(\mc_data_pad_o[16] ) );
  BUFX2 BUFX2_1025 ( .A(_auto_iopadmap_cc_313_execute_56264_17_), .Y(\mc_data_pad_o[17] ) );
  BUFX2 BUFX2_1026 ( .A(_auto_iopadmap_cc_313_execute_56264_18_), .Y(\mc_data_pad_o[18] ) );
  BUFX2 BUFX2_1027 ( .A(_auto_iopadmap_cc_313_execute_56264_19_), .Y(\mc_data_pad_o[19] ) );
  BUFX2 BUFX2_1028 ( .A(_auto_iopadmap_cc_313_execute_56264_20_), .Y(\mc_data_pad_o[20] ) );
  BUFX2 BUFX2_1029 ( .A(_auto_iopadmap_cc_313_execute_56264_21_), .Y(\mc_data_pad_o[21] ) );
  BUFX2 BUFX2_103 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf123) );
  BUFX2 BUFX2_1030 ( .A(_auto_iopadmap_cc_313_execute_56264_22_), .Y(\mc_data_pad_o[22] ) );
  BUFX2 BUFX2_1031 ( .A(_auto_iopadmap_cc_313_execute_56264_23_), .Y(\mc_data_pad_o[23] ) );
  BUFX2 BUFX2_1032 ( .A(_auto_iopadmap_cc_313_execute_56264_24_), .Y(\mc_data_pad_o[24] ) );
  BUFX2 BUFX2_1033 ( .A(_auto_iopadmap_cc_313_execute_56264_25_), .Y(\mc_data_pad_o[25] ) );
  BUFX2 BUFX2_1034 ( .A(_auto_iopadmap_cc_313_execute_56264_26_), .Y(\mc_data_pad_o[26] ) );
  BUFX2 BUFX2_1035 ( .A(_auto_iopadmap_cc_313_execute_56264_27_), .Y(\mc_data_pad_o[27] ) );
  BUFX2 BUFX2_1036 ( .A(_auto_iopadmap_cc_313_execute_56264_28_), .Y(\mc_data_pad_o[28] ) );
  BUFX2 BUFX2_1037 ( .A(_auto_iopadmap_cc_313_execute_56264_29_), .Y(\mc_data_pad_o[29] ) );
  BUFX2 BUFX2_1038 ( .A(_auto_iopadmap_cc_313_execute_56264_30_), .Y(\mc_data_pad_o[30] ) );
  BUFX2 BUFX2_1039 ( .A(_auto_iopadmap_cc_313_execute_56264_31_), .Y(\mc_data_pad_o[31] ) );
  BUFX2 BUFX2_104 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf122) );
  BUFX2 BUFX2_1040 ( .A(_auto_iopadmap_cc_313_execute_56297), .Y(mc_doe_pad_doe_o) );
  BUFX2 BUFX2_1041 ( .A(_auto_iopadmap_cc_313_execute_56299_0_), .Y(\mc_dp_pad_o[0] ) );
  BUFX2 BUFX2_1042 ( .A(_auto_iopadmap_cc_313_execute_56299_1_), .Y(\mc_dp_pad_o[1] ) );
  BUFX2 BUFX2_1043 ( .A(_auto_iopadmap_cc_313_execute_56299_2_), .Y(\mc_dp_pad_o[2] ) );
  BUFX2 BUFX2_1044 ( .A(_auto_iopadmap_cc_313_execute_56299_3_), .Y(\mc_dp_pad_o[3] ) );
  BUFX2 BUFX2_1045 ( .A(_auto_iopadmap_cc_313_execute_56304_0_), .Y(\mc_dqm_pad_o[0] ) );
  BUFX2 BUFX2_1046 ( .A(_auto_iopadmap_cc_313_execute_56304_1_), .Y(\mc_dqm_pad_o[1] ) );
  BUFX2 BUFX2_1047 ( .A(_auto_iopadmap_cc_313_execute_56304_2_), .Y(\mc_dqm_pad_o[2] ) );
  BUFX2 BUFX2_1048 ( .A(_auto_iopadmap_cc_313_execute_56304_3_), .Y(\mc_dqm_pad_o[3] ) );
  BUFX2 BUFX2_1049 ( .A(_auto_iopadmap_cc_313_execute_56309), .Y(mc_oe_pad_o_) );
  BUFX2 BUFX2_105 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf121) );
  BUFX2 BUFX2_1050 ( .A(_auto_iopadmap_cc_313_execute_56311), .Y(mc_ras_pad_o_) );
  BUFX2 BUFX2_1051 ( .A(_auto_iopadmap_cc_313_execute_56313), .Y(mc_rp_pad_o_) );
  BUFX2 BUFX2_1052 ( .A(_auto_iopadmap_cc_313_execute_56315), .Y(mc_vpen_pad_o) );
  BUFX2 BUFX2_1053 ( .A(_auto_iopadmap_cc_313_execute_56317), .Y(mc_we_pad_o_) );
  BUFX2 BUFX2_1054 ( .A(_auto_iopadmap_cc_313_execute_56319), .Y(mc_zz_pad_o) );
  BUFX2 BUFX2_1055 ( .A(_auto_iopadmap_cc_313_execute_56321_0_), .Y(\poc_o[0] ) );
  BUFX2 BUFX2_1056 ( .A(_auto_iopadmap_cc_313_execute_56321_1_), .Y(\poc_o[1] ) );
  BUFX2 BUFX2_1057 ( .A(_auto_iopadmap_cc_313_execute_56321_2_), .Y(\poc_o[2] ) );
  BUFX2 BUFX2_1058 ( .A(_auto_iopadmap_cc_313_execute_56321_3_), .Y(\poc_o[3] ) );
  BUFX2 BUFX2_1059 ( .A(_auto_iopadmap_cc_313_execute_56321_4_), .Y(\poc_o[4] ) );
  BUFX2 BUFX2_106 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf120) );
  BUFX2 BUFX2_1060 ( .A(_auto_iopadmap_cc_313_execute_56321_5_), .Y(\poc_o[5] ) );
  BUFX2 BUFX2_1061 ( .A(_auto_iopadmap_cc_313_execute_56321_6_), .Y(\poc_o[6] ) );
  BUFX2 BUFX2_1062 ( .A(_auto_iopadmap_cc_313_execute_56321_7_), .Y(\poc_o[7] ) );
  BUFX2 BUFX2_1063 ( .A(_auto_iopadmap_cc_313_execute_56321_8_), .Y(\poc_o[8] ) );
  BUFX2 BUFX2_1064 ( .A(_auto_iopadmap_cc_313_execute_56321_9_), .Y(\poc_o[9] ) );
  BUFX2 BUFX2_1065 ( .A(_auto_iopadmap_cc_313_execute_56321_10_), .Y(\poc_o[10] ) );
  BUFX2 BUFX2_1066 ( .A(_auto_iopadmap_cc_313_execute_56321_11_), .Y(\poc_o[11] ) );
  BUFX2 BUFX2_1067 ( .A(_auto_iopadmap_cc_313_execute_56321_12_), .Y(\poc_o[12] ) );
  BUFX2 BUFX2_1068 ( .A(_auto_iopadmap_cc_313_execute_56321_13_), .Y(\poc_o[13] ) );
  BUFX2 BUFX2_1069 ( .A(_auto_iopadmap_cc_313_execute_56321_14_), .Y(\poc_o[14] ) );
  BUFX2 BUFX2_107 ( .A(clk_i_hier0_bF_buf4), .Y(clk_i_bF_buf119) );
  BUFX2 BUFX2_1070 ( .A(_auto_iopadmap_cc_313_execute_56321_15_), .Y(\poc_o[15] ) );
  BUFX2 BUFX2_1071 ( .A(_auto_iopadmap_cc_313_execute_56321_16_), .Y(\poc_o[16] ) );
  BUFX2 BUFX2_1072 ( .A(_auto_iopadmap_cc_313_execute_56321_17_), .Y(\poc_o[17] ) );
  BUFX2 BUFX2_1073 ( .A(_auto_iopadmap_cc_313_execute_56321_18_), .Y(\poc_o[18] ) );
  BUFX2 BUFX2_1074 ( .A(_auto_iopadmap_cc_313_execute_56321_19_), .Y(\poc_o[19] ) );
  BUFX2 BUFX2_1075 ( .A(_auto_iopadmap_cc_313_execute_56321_20_), .Y(\poc_o[20] ) );
  BUFX2 BUFX2_1076 ( .A(_auto_iopadmap_cc_313_execute_56321_21_), .Y(\poc_o[21] ) );
  BUFX2 BUFX2_1077 ( .A(_auto_iopadmap_cc_313_execute_56321_22_), .Y(\poc_o[22] ) );
  BUFX2 BUFX2_1078 ( .A(_auto_iopadmap_cc_313_execute_56321_23_), .Y(\poc_o[23] ) );
  BUFX2 BUFX2_1079 ( .A(_auto_iopadmap_cc_313_execute_56321_24_), .Y(\poc_o[24] ) );
  BUFX2 BUFX2_108 ( .A(clk_i_hier0_bF_buf3), .Y(clk_i_bF_buf118) );
  BUFX2 BUFX2_1080 ( .A(_auto_iopadmap_cc_313_execute_56321_25_), .Y(\poc_o[25] ) );
  BUFX2 BUFX2_1081 ( .A(_auto_iopadmap_cc_313_execute_56321_26_), .Y(\poc_o[26] ) );
  BUFX2 BUFX2_1082 ( .A(_auto_iopadmap_cc_313_execute_56321_27_), .Y(\poc_o[27] ) );
  BUFX2 BUFX2_1083 ( .A(_auto_iopadmap_cc_313_execute_56321_28_), .Y(\poc_o[28] ) );
  BUFX2 BUFX2_1084 ( .A(_auto_iopadmap_cc_313_execute_56321_29_), .Y(\poc_o[29] ) );
  BUFX2 BUFX2_1085 ( .A(_auto_iopadmap_cc_313_execute_56321_30_), .Y(\poc_o[30] ) );
  BUFX2 BUFX2_1086 ( .A(_auto_iopadmap_cc_313_execute_56321_31_), .Y(\poc_o[31] ) );
  BUFX2 BUFX2_1087 ( .A(_auto_iopadmap_cc_313_execute_56354), .Y(suspended_o) );
  BUFX2 BUFX2_1088 ( .A(_auto_iopadmap_cc_313_execute_56356), .Y(wb_ack_o) );
  BUFX2 BUFX2_1089 ( .A(_auto_iopadmap_cc_313_execute_56358_0_), .Y(\wb_data_o[0] ) );
  BUFX2 BUFX2_109 ( .A(clk_i_hier0_bF_buf2), .Y(clk_i_bF_buf117) );
  BUFX2 BUFX2_1090 ( .A(_auto_iopadmap_cc_313_execute_56358_1_), .Y(\wb_data_o[1] ) );
  BUFX2 BUFX2_1091 ( .A(_auto_iopadmap_cc_313_execute_56358_2_), .Y(\wb_data_o[2] ) );
  BUFX2 BUFX2_1092 ( .A(_auto_iopadmap_cc_313_execute_56358_3_), .Y(\wb_data_o[3] ) );
  BUFX2 BUFX2_1093 ( .A(_auto_iopadmap_cc_313_execute_56358_4_), .Y(\wb_data_o[4] ) );
  BUFX2 BUFX2_1094 ( .A(_auto_iopadmap_cc_313_execute_56358_5_), .Y(\wb_data_o[5] ) );
  BUFX2 BUFX2_1095 ( .A(_auto_iopadmap_cc_313_execute_56358_6_), .Y(\wb_data_o[6] ) );
  BUFX2 BUFX2_1096 ( .A(_auto_iopadmap_cc_313_execute_56358_7_), .Y(\wb_data_o[7] ) );
  BUFX2 BUFX2_1097 ( .A(_auto_iopadmap_cc_313_execute_56358_8_), .Y(\wb_data_o[8] ) );
  BUFX2 BUFX2_1098 ( .A(_auto_iopadmap_cc_313_execute_56358_9_), .Y(\wb_data_o[9] ) );
  BUFX2 BUFX2_1099 ( .A(_auto_iopadmap_cc_313_execute_56358_10_), .Y(\wb_data_o[10] ) );
  BUFX2 BUFX2_11 ( .A(clk_i), .Y(clk_i_hier0_bF_buf0) );
  BUFX2 BUFX2_110 ( .A(clk_i_hier0_bF_buf1), .Y(clk_i_bF_buf116) );
  BUFX2 BUFX2_1100 ( .A(_auto_iopadmap_cc_313_execute_56358_11_), .Y(\wb_data_o[11] ) );
  BUFX2 BUFX2_1101 ( .A(_auto_iopadmap_cc_313_execute_56358_12_), .Y(\wb_data_o[12] ) );
  BUFX2 BUFX2_1102 ( .A(_auto_iopadmap_cc_313_execute_56358_13_), .Y(\wb_data_o[13] ) );
  BUFX2 BUFX2_1103 ( .A(_auto_iopadmap_cc_313_execute_56358_14_), .Y(\wb_data_o[14] ) );
  BUFX2 BUFX2_1104 ( .A(_auto_iopadmap_cc_313_execute_56358_15_), .Y(\wb_data_o[15] ) );
  BUFX2 BUFX2_1105 ( .A(_auto_iopadmap_cc_313_execute_56358_16_), .Y(\wb_data_o[16] ) );
  BUFX2 BUFX2_1106 ( .A(_auto_iopadmap_cc_313_execute_56358_17_), .Y(\wb_data_o[17] ) );
  BUFX2 BUFX2_1107 ( .A(_auto_iopadmap_cc_313_execute_56358_18_), .Y(\wb_data_o[18] ) );
  BUFX2 BUFX2_1108 ( .A(_auto_iopadmap_cc_313_execute_56358_19_), .Y(\wb_data_o[19] ) );
  BUFX2 BUFX2_1109 ( .A(_auto_iopadmap_cc_313_execute_56358_20_), .Y(\wb_data_o[20] ) );
  BUFX2 BUFX2_111 ( .A(clk_i_hier0_bF_buf0), .Y(clk_i_bF_buf115) );
  BUFX2 BUFX2_1110 ( .A(_auto_iopadmap_cc_313_execute_56358_21_), .Y(\wb_data_o[21] ) );
  BUFX2 BUFX2_1111 ( .A(_auto_iopadmap_cc_313_execute_56358_22_), .Y(\wb_data_o[22] ) );
  BUFX2 BUFX2_1112 ( .A(_auto_iopadmap_cc_313_execute_56358_23_), .Y(\wb_data_o[23] ) );
  BUFX2 BUFX2_1113 ( .A(_auto_iopadmap_cc_313_execute_56358_24_), .Y(\wb_data_o[24] ) );
  BUFX2 BUFX2_1114 ( .A(_auto_iopadmap_cc_313_execute_56358_25_), .Y(\wb_data_o[25] ) );
  BUFX2 BUFX2_1115 ( .A(_auto_iopadmap_cc_313_execute_56358_26_), .Y(\wb_data_o[26] ) );
  BUFX2 BUFX2_1116 ( .A(_auto_iopadmap_cc_313_execute_56358_27_), .Y(\wb_data_o[27] ) );
  BUFX2 BUFX2_1117 ( .A(_auto_iopadmap_cc_313_execute_56358_28_), .Y(\wb_data_o[28] ) );
  BUFX2 BUFX2_1118 ( .A(_auto_iopadmap_cc_313_execute_56358_29_), .Y(\wb_data_o[29] ) );
  BUFX2 BUFX2_1119 ( .A(_auto_iopadmap_cc_313_execute_56358_30_), .Y(\wb_data_o[30] ) );
  BUFX2 BUFX2_112 ( .A(clk_i_hier0_bF_buf10), .Y(clk_i_bF_buf114) );
  BUFX2 BUFX2_1120 ( .A(_auto_iopadmap_cc_313_execute_56358_31_), .Y(\wb_data_o[31] ) );
  BUFX2 BUFX2_1121 ( .A(_auto_iopadmap_cc_313_execute_56391), .Y(wb_err_o) );
  BUFX2 BUFX2_113 ( .A(clk_i_hier0_bF_buf9), .Y(clk_i_bF_buf113) );
  BUFX2 BUFX2_114 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf112) );
  BUFX2 BUFX2_115 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf111) );
  BUFX2 BUFX2_116 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf110) );
  BUFX2 BUFX2_117 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf109) );
  BUFX2 BUFX2_118 ( .A(clk_i_hier0_bF_buf4), .Y(clk_i_bF_buf108) );
  BUFX2 BUFX2_119 ( .A(clk_i_hier0_bF_buf3), .Y(clk_i_bF_buf107) );
  BUFX2 BUFX2_12 ( .A(u0_u3__abc_44466_n239_1), .Y(u0_u3__abc_44466_n239_1_bF_buf4) );
  BUFX2 BUFX2_120 ( .A(clk_i_hier0_bF_buf2), .Y(clk_i_bF_buf106) );
  BUFX2 BUFX2_121 ( .A(clk_i_hier0_bF_buf1), .Y(clk_i_bF_buf105) );
  BUFX2 BUFX2_122 ( .A(clk_i_hier0_bF_buf0), .Y(clk_i_bF_buf104) );
  BUFX2 BUFX2_123 ( .A(clk_i_hier0_bF_buf10), .Y(clk_i_bF_buf103) );
  BUFX2 BUFX2_124 ( .A(clk_i_hier0_bF_buf9), .Y(clk_i_bF_buf102) );
  BUFX2 BUFX2_125 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf101) );
  BUFX2 BUFX2_126 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf100) );
  BUFX2 BUFX2_127 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf99) );
  BUFX2 BUFX2_128 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf98) );
  BUFX2 BUFX2_129 ( .A(clk_i_hier0_bF_buf4), .Y(clk_i_bF_buf97) );
  BUFX2 BUFX2_13 ( .A(u0_u3__abc_44466_n239_1), .Y(u0_u3__abc_44466_n239_1_bF_buf3) );
  BUFX2 BUFX2_130 ( .A(clk_i_hier0_bF_buf3), .Y(clk_i_bF_buf96) );
  BUFX2 BUFX2_131 ( .A(clk_i_hier0_bF_buf2), .Y(clk_i_bF_buf95) );
  BUFX2 BUFX2_132 ( .A(clk_i_hier0_bF_buf1), .Y(clk_i_bF_buf94) );
  BUFX2 BUFX2_133 ( .A(clk_i_hier0_bF_buf0), .Y(clk_i_bF_buf93) );
  BUFX2 BUFX2_134 ( .A(clk_i_hier0_bF_buf10), .Y(clk_i_bF_buf92) );
  BUFX2 BUFX2_135 ( .A(clk_i_hier0_bF_buf9), .Y(clk_i_bF_buf91) );
  BUFX2 BUFX2_136 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf90) );
  BUFX2 BUFX2_137 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf89) );
  BUFX2 BUFX2_138 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf88) );
  BUFX2 BUFX2_139 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf87) );
  BUFX2 BUFX2_14 ( .A(u0_u3__abc_44466_n239_1), .Y(u0_u3__abc_44466_n239_1_bF_buf2) );
  BUFX2 BUFX2_140 ( .A(clk_i_hier0_bF_buf4), .Y(clk_i_bF_buf86) );
  BUFX2 BUFX2_141 ( .A(clk_i_hier0_bF_buf3), .Y(clk_i_bF_buf85) );
  BUFX2 BUFX2_142 ( .A(clk_i_hier0_bF_buf2), .Y(clk_i_bF_buf84) );
  BUFX2 BUFX2_143 ( .A(clk_i_hier0_bF_buf1), .Y(clk_i_bF_buf83) );
  BUFX2 BUFX2_144 ( .A(clk_i_hier0_bF_buf0), .Y(clk_i_bF_buf82) );
  BUFX2 BUFX2_145 ( .A(clk_i_hier0_bF_buf10), .Y(clk_i_bF_buf81) );
  BUFX2 BUFX2_146 ( .A(clk_i_hier0_bF_buf9), .Y(clk_i_bF_buf80) );
  BUFX2 BUFX2_147 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf79) );
  BUFX2 BUFX2_148 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf78) );
  BUFX2 BUFX2_149 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf77) );
  BUFX2 BUFX2_15 ( .A(u0_u3__abc_44466_n239_1), .Y(u0_u3__abc_44466_n239_1_bF_buf1) );
  BUFX2 BUFX2_150 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf76) );
  BUFX2 BUFX2_151 ( .A(clk_i_hier0_bF_buf4), .Y(clk_i_bF_buf75) );
  BUFX2 BUFX2_152 ( .A(clk_i_hier0_bF_buf3), .Y(clk_i_bF_buf74) );
  BUFX2 BUFX2_153 ( .A(clk_i_hier0_bF_buf2), .Y(clk_i_bF_buf73) );
  BUFX2 BUFX2_154 ( .A(clk_i_hier0_bF_buf1), .Y(clk_i_bF_buf72) );
  BUFX2 BUFX2_155 ( .A(clk_i_hier0_bF_buf0), .Y(clk_i_bF_buf71) );
  BUFX2 BUFX2_156 ( .A(clk_i_hier0_bF_buf10), .Y(clk_i_bF_buf70) );
  BUFX2 BUFX2_157 ( .A(clk_i_hier0_bF_buf9), .Y(clk_i_bF_buf69) );
  BUFX2 BUFX2_158 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf68) );
  BUFX2 BUFX2_159 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf67) );
  BUFX2 BUFX2_16 ( .A(u0_u3__abc_44466_n239_1), .Y(u0_u3__abc_44466_n239_1_bF_buf0) );
  BUFX2 BUFX2_160 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf66) );
  BUFX2 BUFX2_161 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf65) );
  BUFX2 BUFX2_162 ( .A(clk_i_hier0_bF_buf4), .Y(clk_i_bF_buf64) );
  BUFX2 BUFX2_163 ( .A(clk_i_hier0_bF_buf3), .Y(clk_i_bF_buf63) );
  BUFX2 BUFX2_164 ( .A(clk_i_hier0_bF_buf2), .Y(clk_i_bF_buf62) );
  BUFX2 BUFX2_165 ( .A(clk_i_hier0_bF_buf1), .Y(clk_i_bF_buf61) );
  BUFX2 BUFX2_166 ( .A(clk_i_hier0_bF_buf0), .Y(clk_i_bF_buf60) );
  BUFX2 BUFX2_167 ( .A(clk_i_hier0_bF_buf10), .Y(clk_i_bF_buf59) );
  BUFX2 BUFX2_168 ( .A(clk_i_hier0_bF_buf9), .Y(clk_i_bF_buf58) );
  BUFX2 BUFX2_169 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf57) );
  BUFX2 BUFX2_17 ( .A(u0_u3_rst_r2), .Y(u0_u3_rst_r2_bF_buf5) );
  BUFX2 BUFX2_170 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf56) );
  BUFX2 BUFX2_171 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf55) );
  BUFX2 BUFX2_172 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf54) );
  BUFX2 BUFX2_173 ( .A(clk_i_hier0_bF_buf4), .Y(clk_i_bF_buf53) );
  BUFX2 BUFX2_174 ( .A(clk_i_hier0_bF_buf3), .Y(clk_i_bF_buf52) );
  BUFX2 BUFX2_175 ( .A(clk_i_hier0_bF_buf2), .Y(clk_i_bF_buf51) );
  BUFX2 BUFX2_176 ( .A(clk_i_hier0_bF_buf1), .Y(clk_i_bF_buf50) );
  BUFX2 BUFX2_177 ( .A(clk_i_hier0_bF_buf0), .Y(clk_i_bF_buf49) );
  BUFX2 BUFX2_178 ( .A(clk_i_hier0_bF_buf10), .Y(clk_i_bF_buf48) );
  BUFX2 BUFX2_179 ( .A(clk_i_hier0_bF_buf9), .Y(clk_i_bF_buf47) );
  BUFX2 BUFX2_18 ( .A(u0_u3_rst_r2), .Y(u0_u3_rst_r2_bF_buf4) );
  BUFX2 BUFX2_180 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf46) );
  BUFX2 BUFX2_181 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf45) );
  BUFX2 BUFX2_182 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf44) );
  BUFX2 BUFX2_183 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf43) );
  BUFX2 BUFX2_184 ( .A(clk_i_hier0_bF_buf4), .Y(clk_i_bF_buf42) );
  BUFX2 BUFX2_185 ( .A(clk_i_hier0_bF_buf3), .Y(clk_i_bF_buf41) );
  BUFX2 BUFX2_186 ( .A(clk_i_hier0_bF_buf2), .Y(clk_i_bF_buf40) );
  BUFX2 BUFX2_187 ( .A(clk_i_hier0_bF_buf1), .Y(clk_i_bF_buf39) );
  BUFX2 BUFX2_188 ( .A(clk_i_hier0_bF_buf0), .Y(clk_i_bF_buf38) );
  BUFX2 BUFX2_189 ( .A(clk_i_hier0_bF_buf10), .Y(clk_i_bF_buf37) );
  BUFX2 BUFX2_19 ( .A(u0_u3_rst_r2), .Y(u0_u3_rst_r2_bF_buf3) );
  BUFX2 BUFX2_190 ( .A(clk_i_hier0_bF_buf9), .Y(clk_i_bF_buf36) );
  BUFX2 BUFX2_191 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf35) );
  BUFX2 BUFX2_192 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf34) );
  BUFX2 BUFX2_193 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf33) );
  BUFX2 BUFX2_194 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf32) );
  BUFX2 BUFX2_195 ( .A(clk_i_hier0_bF_buf4), .Y(clk_i_bF_buf31) );
  BUFX2 BUFX2_196 ( .A(clk_i_hier0_bF_buf3), .Y(clk_i_bF_buf30) );
  BUFX2 BUFX2_197 ( .A(clk_i_hier0_bF_buf2), .Y(clk_i_bF_buf29) );
  BUFX2 BUFX2_198 ( .A(clk_i_hier0_bF_buf1), .Y(clk_i_bF_buf28) );
  BUFX2 BUFX2_199 ( .A(clk_i_hier0_bF_buf0), .Y(clk_i_bF_buf27) );
  BUFX2 BUFX2_2 ( .A(clk_i), .Y(clk_i_hier0_bF_buf9) );
  BUFX2 BUFX2_20 ( .A(u0_u3_rst_r2), .Y(u0_u3_rst_r2_bF_buf2) );
  BUFX2 BUFX2_200 ( .A(clk_i_hier0_bF_buf10), .Y(clk_i_bF_buf26) );
  BUFX2 BUFX2_201 ( .A(clk_i_hier0_bF_buf9), .Y(clk_i_bF_buf25) );
  BUFX2 BUFX2_202 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf24) );
  BUFX2 BUFX2_203 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf23) );
  BUFX2 BUFX2_204 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf22) );
  BUFX2 BUFX2_205 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf21) );
  BUFX2 BUFX2_206 ( .A(clk_i_hier0_bF_buf4), .Y(clk_i_bF_buf20) );
  BUFX2 BUFX2_207 ( .A(clk_i_hier0_bF_buf3), .Y(clk_i_bF_buf19) );
  BUFX2 BUFX2_208 ( .A(clk_i_hier0_bF_buf2), .Y(clk_i_bF_buf18) );
  BUFX2 BUFX2_209 ( .A(clk_i_hier0_bF_buf1), .Y(clk_i_bF_buf17) );
  BUFX2 BUFX2_21 ( .A(u0_u3_rst_r2), .Y(u0_u3_rst_r2_bF_buf1) );
  BUFX2 BUFX2_210 ( .A(clk_i_hier0_bF_buf0), .Y(clk_i_bF_buf16) );
  BUFX2 BUFX2_211 ( .A(clk_i_hier0_bF_buf10), .Y(clk_i_bF_buf15) );
  BUFX2 BUFX2_212 ( .A(clk_i_hier0_bF_buf9), .Y(clk_i_bF_buf14) );
  BUFX2 BUFX2_213 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf13) );
  BUFX2 BUFX2_214 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf12) );
  BUFX2 BUFX2_215 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf11) );
  BUFX2 BUFX2_216 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf10) );
  BUFX2 BUFX2_217 ( .A(clk_i_hier0_bF_buf4), .Y(clk_i_bF_buf9) );
  BUFX2 BUFX2_218 ( .A(clk_i_hier0_bF_buf3), .Y(clk_i_bF_buf8) );
  BUFX2 BUFX2_219 ( .A(clk_i_hier0_bF_buf2), .Y(clk_i_bF_buf7) );
  BUFX2 BUFX2_22 ( .A(u0_u3_rst_r2), .Y(u0_u3_rst_r2_bF_buf0) );
  BUFX2 BUFX2_220 ( .A(clk_i_hier0_bF_buf1), .Y(clk_i_bF_buf6) );
  BUFX2 BUFX2_221 ( .A(clk_i_hier0_bF_buf0), .Y(clk_i_bF_buf5) );
  BUFX2 BUFX2_222 ( .A(clk_i_hier0_bF_buf10), .Y(clk_i_bF_buf4) );
  BUFX2 BUFX2_223 ( .A(clk_i_hier0_bF_buf9), .Y(clk_i_bF_buf3) );
  BUFX2 BUFX2_224 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf2) );
  BUFX2 BUFX2_225 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf1) );
  BUFX2 BUFX2_226 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf0) );
  BUFX2 BUFX2_227 ( .A(u0__abc_49347_n2723), .Y(u0__abc_49347_n2723_bF_buf5) );
  BUFX2 BUFX2_228 ( .A(u0__abc_49347_n2723), .Y(u0__abc_49347_n2723_bF_buf4) );
  BUFX2 BUFX2_229 ( .A(u0__abc_49347_n2723), .Y(u0__abc_49347_n2723_bF_buf3) );
  BUFX2 BUFX2_23 ( .A(u3_u0__abc_48231_n382), .Y(u3_u0__abc_48231_n382_bF_buf7) );
  BUFX2 BUFX2_230 ( .A(u0__abc_49347_n2723), .Y(u0__abc_49347_n2723_bF_buf2) );
  BUFX2 BUFX2_231 ( .A(u0__abc_49347_n2723), .Y(u0__abc_49347_n2723_bF_buf1) );
  BUFX2 BUFX2_232 ( .A(u0__abc_49347_n2723), .Y(u0__abc_49347_n2723_bF_buf0) );
  BUFX2 BUFX2_233 ( .A(u0__abc_49347_n2724), .Y(u0__abc_49347_n2724_bF_buf5) );
  BUFX2 BUFX2_234 ( .A(u0__abc_49347_n2724), .Y(u0__abc_49347_n2724_bF_buf4) );
  BUFX2 BUFX2_235 ( .A(u0__abc_49347_n2724), .Y(u0__abc_49347_n2724_bF_buf3) );
  BUFX2 BUFX2_236 ( .A(u0__abc_49347_n2724), .Y(u0__abc_49347_n2724_bF_buf2) );
  BUFX2 BUFX2_237 ( .A(u0__abc_49347_n2724), .Y(u0__abc_49347_n2724_bF_buf1) );
  BUFX2 BUFX2_238 ( .A(u0__abc_49347_n2724), .Y(u0__abc_49347_n2724_bF_buf0) );
  BUFX2 BUFX2_239 ( .A(u0__abc_49347_n2725), .Y(u0__abc_49347_n2725_bF_buf5) );
  BUFX2 BUFX2_24 ( .A(u3_u0__abc_48231_n382), .Y(u3_u0__abc_48231_n382_bF_buf6) );
  BUFX2 BUFX2_240 ( .A(u0__abc_49347_n2725), .Y(u0__abc_49347_n2725_bF_buf4) );
  BUFX2 BUFX2_241 ( .A(u0__abc_49347_n2725), .Y(u0__abc_49347_n2725_bF_buf3) );
  BUFX2 BUFX2_242 ( .A(u0__abc_49347_n2725), .Y(u0__abc_49347_n2725_bF_buf2) );
  BUFX2 BUFX2_243 ( .A(u0__abc_49347_n2725), .Y(u0__abc_49347_n2725_bF_buf1) );
  BUFX2 BUFX2_244 ( .A(u0__abc_49347_n2725), .Y(u0__abc_49347_n2725_bF_buf0) );
  BUFX2 BUFX2_245 ( .A(u0__abc_49347_n2726), .Y(u0__abc_49347_n2726_bF_buf5) );
  BUFX2 BUFX2_246 ( .A(u0__abc_49347_n2726), .Y(u0__abc_49347_n2726_bF_buf4) );
  BUFX2 BUFX2_247 ( .A(u0__abc_49347_n2726), .Y(u0__abc_49347_n2726_bF_buf3) );
  BUFX2 BUFX2_248 ( .A(u0__abc_49347_n2726), .Y(u0__abc_49347_n2726_bF_buf2) );
  BUFX2 BUFX2_249 ( .A(u0__abc_49347_n2726), .Y(u0__abc_49347_n2726_bF_buf1) );
  BUFX2 BUFX2_25 ( .A(u3_u0__abc_48231_n382), .Y(u3_u0__abc_48231_n382_bF_buf5) );
  BUFX2 BUFX2_250 ( .A(u0__abc_49347_n2726), .Y(u0__abc_49347_n2726_bF_buf0) );
  BUFX2 BUFX2_251 ( .A(u0__abc_49347_n2728), .Y(u0__abc_49347_n2728_bF_buf5) );
  BUFX2 BUFX2_252 ( .A(u0__abc_49347_n2728), .Y(u0__abc_49347_n2728_bF_buf4) );
  BUFX2 BUFX2_253 ( .A(u0__abc_49347_n2728), .Y(u0__abc_49347_n2728_bF_buf3) );
  BUFX2 BUFX2_254 ( .A(u0__abc_49347_n2728), .Y(u0__abc_49347_n2728_bF_buf2) );
  BUFX2 BUFX2_255 ( .A(u0__abc_49347_n2728), .Y(u0__abc_49347_n2728_bF_buf1) );
  BUFX2 BUFX2_256 ( .A(u0__abc_49347_n2728), .Y(u0__abc_49347_n2728_bF_buf0) );
  BUFX2 BUFX2_257 ( .A(bank_adr_1_), .Y(bank_adr_1_bF_buf3) );
  BUFX2 BUFX2_258 ( .A(bank_adr_1_), .Y(bank_adr_1_bF_buf2) );
  BUFX2 BUFX2_259 ( .A(bank_adr_1_), .Y(bank_adr_1_bF_buf1) );
  BUFX2 BUFX2_26 ( .A(u3_u0__abc_48231_n382), .Y(u3_u0__abc_48231_n382_bF_buf4) );
  BUFX2 BUFX2_260 ( .A(bank_adr_1_), .Y(bank_adr_1_bF_buf0) );
  BUFX2 BUFX2_261 ( .A(u0__abc_49347_n1953_1), .Y(u0__abc_49347_n1953_1_bF_buf3) );
  BUFX2 BUFX2_262 ( .A(u0__abc_49347_n1953_1), .Y(u0__abc_49347_n1953_1_bF_buf2) );
  BUFX2 BUFX2_263 ( .A(u0__abc_49347_n1953_1), .Y(u0__abc_49347_n1953_1_bF_buf1) );
  BUFX2 BUFX2_264 ( .A(u0__abc_49347_n1953_1), .Y(u0__abc_49347_n1953_1_bF_buf0) );
  BUFX2 BUFX2_265 ( .A(u0__abc_49347_n4571), .Y(u0__abc_49347_n4571_bF_buf4) );
  BUFX2 BUFX2_266 ( .A(u0__abc_49347_n4571), .Y(u0__abc_49347_n4571_bF_buf3) );
  BUFX2 BUFX2_267 ( .A(u0__abc_49347_n4571), .Y(u0__abc_49347_n4571_bF_buf2) );
  BUFX2 BUFX2_268 ( .A(u0__abc_49347_n4571), .Y(u0__abc_49347_n4571_bF_buf1) );
  BUFX2 BUFX2_269 ( .A(u0__abc_49347_n4571), .Y(u0__abc_49347_n4571_bF_buf0) );
  BUFX2 BUFX2_27 ( .A(u3_u0__abc_48231_n382), .Y(u3_u0__abc_48231_n382_bF_buf3) );
  BUFX2 BUFX2_270 ( .A(u2_u3__abc_47660_n137), .Y(u2_u3__abc_47660_n137_bF_buf4) );
  BUFX2 BUFX2_271 ( .A(u2_u3__abc_47660_n137), .Y(u2_u3__abc_47660_n137_bF_buf3) );
  BUFX2 BUFX2_272 ( .A(u2_u3__abc_47660_n137), .Y(u2_u3__abc_47660_n137_bF_buf2) );
  BUFX2 BUFX2_273 ( .A(u2_u3__abc_47660_n137), .Y(u2_u3__abc_47660_n137_bF_buf1) );
  BUFX2 BUFX2_274 ( .A(u2_u3__abc_47660_n137), .Y(u2_u3__abc_47660_n137_bF_buf0) );
  BUFX2 BUFX2_275 ( .A(u3_u0__abc_48231_n1034), .Y(u3_u0__abc_48231_n1034_bF_buf5) );
  BUFX2 BUFX2_276 ( .A(u3_u0__abc_48231_n1034), .Y(u3_u0__abc_48231_n1034_bF_buf4) );
  BUFX2 BUFX2_277 ( .A(u3_u0__abc_48231_n1034), .Y(u3_u0__abc_48231_n1034_bF_buf3) );
  BUFX2 BUFX2_278 ( .A(u3_u0__abc_48231_n1034), .Y(u3_u0__abc_48231_n1034_bF_buf2) );
  BUFX2 BUFX2_279 ( .A(u3_u0__abc_48231_n1034), .Y(u3_u0__abc_48231_n1034_bF_buf1) );
  BUFX2 BUFX2_28 ( .A(u3_u0__abc_48231_n382), .Y(u3_u0__abc_48231_n382_bF_buf2) );
  BUFX2 BUFX2_280 ( .A(u3_u0__abc_48231_n1034), .Y(u3_u0__abc_48231_n1034_bF_buf0) );
  BUFX2 BUFX2_281 ( .A(spec_req_cs_5_), .Y(spec_req_cs_5_bF_buf5) );
  BUFX2 BUFX2_282 ( .A(spec_req_cs_5_), .Y(spec_req_cs_5_bF_buf4) );
  BUFX2 BUFX2_283 ( .A(spec_req_cs_5_), .Y(spec_req_cs_5_bF_buf3) );
  BUFX2 BUFX2_284 ( .A(spec_req_cs_5_), .Y(spec_req_cs_5_bF_buf2) );
  BUFX2 BUFX2_285 ( .A(spec_req_cs_5_), .Y(spec_req_cs_5_bF_buf1) );
  BUFX2 BUFX2_286 ( .A(spec_req_cs_5_), .Y(spec_req_cs_5_bF_buf0) );
  BUFX2 BUFX2_287 ( .A(row_adr_10_), .Y(row_adr_10_bF_buf6) );
  BUFX2 BUFX2_288 ( .A(row_adr_10_), .Y(row_adr_10_bF_buf5) );
  BUFX2 BUFX2_289 ( .A(row_adr_10_), .Y(row_adr_10_bF_buf4) );
  BUFX2 BUFX2_29 ( .A(u3_u0__abc_48231_n382), .Y(u3_u0__abc_48231_n382_bF_buf1) );
  BUFX2 BUFX2_290 ( .A(row_adr_10_), .Y(row_adr_10_bF_buf3) );
  BUFX2 BUFX2_291 ( .A(row_adr_10_), .Y(row_adr_10_bF_buf2) );
  BUFX2 BUFX2_292 ( .A(row_adr_10_), .Y(row_adr_10_bF_buf1) );
  BUFX2 BUFX2_293 ( .A(row_adr_10_), .Y(row_adr_10_bF_buf0) );
  BUFX2 BUFX2_294 ( .A(u0__abc_49347_n4511), .Y(u0__abc_49347_n4511_bF_buf4) );
  BUFX2 BUFX2_295 ( .A(u0__abc_49347_n4511), .Y(u0__abc_49347_n4511_bF_buf3) );
  BUFX2 BUFX2_296 ( .A(u0__abc_49347_n4511), .Y(u0__abc_49347_n4511_bF_buf2) );
  BUFX2 BUFX2_297 ( .A(u0__abc_49347_n4511), .Y(u0__abc_49347_n4511_bF_buf1) );
  BUFX2 BUFX2_298 ( .A(u0__abc_49347_n4511), .Y(u0__abc_49347_n4511_bF_buf0) );
  BUFX2 BUFX2_299 ( .A(u0__abc_49347_n4516), .Y(u0__abc_49347_n4516_bF_buf4) );
  BUFX2 BUFX2_3 ( .A(clk_i), .Y(clk_i_hier0_bF_buf8) );
  BUFX2 BUFX2_30 ( .A(u3_u0__abc_48231_n382), .Y(u3_u0__abc_48231_n382_bF_buf0) );
  BUFX2 BUFX2_300 ( .A(u0__abc_49347_n4516), .Y(u0__abc_49347_n4516_bF_buf3) );
  BUFX2 BUFX2_301 ( .A(u0__abc_49347_n4516), .Y(u0__abc_49347_n4516_bF_buf2) );
  BUFX2 BUFX2_302 ( .A(u0__abc_49347_n4516), .Y(u0__abc_49347_n4516_bF_buf1) );
  BUFX2 BUFX2_303 ( .A(u0__abc_49347_n4516), .Y(u0__abc_49347_n4516_bF_buf0) );
  BUFX2 BUFX2_304 ( .A(u0__abc_49347_n4519), .Y(u0__abc_49347_n4519_bF_buf4) );
  BUFX2 BUFX2_305 ( .A(u0__abc_49347_n4519), .Y(u0__abc_49347_n4519_bF_buf3) );
  BUFX2 BUFX2_306 ( .A(u0__abc_49347_n4519), .Y(u0__abc_49347_n4519_bF_buf2) );
  BUFX2 BUFX2_307 ( .A(u0__abc_49347_n4519), .Y(u0__abc_49347_n4519_bF_buf1) );
  BUFX2 BUFX2_308 ( .A(u0__abc_49347_n4519), .Y(u0__abc_49347_n4519_bF_buf0) );
  BUFX2 BUFX2_309 ( .A(spec_req_cs_2_), .Y(spec_req_cs_2_bF_buf5) );
  BUFX2 BUFX2_31 ( .A(u0_u1_lmr_req_we_FF_INPUT), .Y(u0_u1_lmr_req_we_FF_INPUT_bF_buf7) );
  BUFX2 BUFX2_310 ( .A(spec_req_cs_2_), .Y(spec_req_cs_2_bF_buf4) );
  BUFX2 BUFX2_311 ( .A(spec_req_cs_2_), .Y(spec_req_cs_2_bF_buf3) );
  BUFX2 BUFX2_312 ( .A(spec_req_cs_2_), .Y(spec_req_cs_2_bF_buf2) );
  BUFX2 BUFX2_313 ( .A(spec_req_cs_2_), .Y(spec_req_cs_2_bF_buf1) );
  BUFX2 BUFX2_314 ( .A(spec_req_cs_2_), .Y(spec_req_cs_2_bF_buf0) );
  BUFX2 BUFX2_315 ( .A(csc_5_), .Y(csc_5_bF_buf4) );
  BUFX2 BUFX2_316 ( .A(csc_5_), .Y(csc_5_bF_buf3) );
  BUFX2 BUFX2_317 ( .A(csc_5_), .Y(csc_5_bF_buf2) );
  BUFX2 BUFX2_318 ( .A(csc_5_), .Y(csc_5_bF_buf1) );
  BUFX2 BUFX2_319 ( .A(csc_5_), .Y(csc_5_bF_buf0) );
  BUFX2 BUFX2_32 ( .A(u0_u1_lmr_req_we_FF_INPUT), .Y(u0_u1_lmr_req_we_FF_INPUT_bF_buf6) );
  BUFX2 BUFX2_320 ( .A(u2_u1__abc_47660_n137), .Y(u2_u1__abc_47660_n137_bF_buf4) );
  BUFX2 BUFX2_321 ( .A(u2_u1__abc_47660_n137), .Y(u2_u1__abc_47660_n137_bF_buf3) );
  BUFX2 BUFX2_322 ( .A(u2_u1__abc_47660_n137), .Y(u2_u1__abc_47660_n137_bF_buf2) );
  BUFX2 BUFX2_323 ( .A(u2_u1__abc_47660_n137), .Y(u2_u1__abc_47660_n137_bF_buf1) );
  BUFX2 BUFX2_324 ( .A(u2_u1__abc_47660_n137), .Y(u2_u1__abc_47660_n137_bF_buf0) );
  BUFX2 BUFX2_325 ( .A(u1__abc_45852_n893), .Y(u1__abc_45852_n893_bF_buf4) );
  BUFX2 BUFX2_326 ( .A(u1__abc_45852_n893), .Y(u1__abc_45852_n893_bF_buf3) );
  BUFX2 BUFX2_327 ( .A(u1__abc_45852_n893), .Y(u1__abc_45852_n893_bF_buf2) );
  BUFX2 BUFX2_328 ( .A(u1__abc_45852_n893), .Y(u1__abc_45852_n893_bF_buf1) );
  BUFX2 BUFX2_329 ( .A(u1__abc_45852_n893), .Y(u1__abc_45852_n893_bF_buf0) );
  BUFX2 BUFX2_33 ( .A(u0_u1_lmr_req_we_FF_INPUT), .Y(u0_u1_lmr_req_we_FF_INPUT_bF_buf5) );
  BUFX2 BUFX2_330 ( .A(u1__abc_45852_n897), .Y(u1__abc_45852_n897_bF_buf3) );
  BUFX2 BUFX2_331 ( .A(u1__abc_45852_n897), .Y(u1__abc_45852_n897_bF_buf2) );
  BUFX2 BUFX2_332 ( .A(u1__abc_45852_n897), .Y(u1__abc_45852_n897_bF_buf1) );
  BUFX2 BUFX2_333 ( .A(u1__abc_45852_n897), .Y(u1__abc_45852_n897_bF_buf0) );
  BUFX2 BUFX2_334 ( .A(u5__abc_54027_n1575), .Y(u5__abc_54027_n1575_bF_buf6) );
  BUFX2 BUFX2_335 ( .A(u5__abc_54027_n1575), .Y(u5__abc_54027_n1575_bF_buf5) );
  BUFX2 BUFX2_336 ( .A(u5__abc_54027_n1575), .Y(u5__abc_54027_n1575_bF_buf4) );
  BUFX2 BUFX2_337 ( .A(u5__abc_54027_n1575), .Y(u5__abc_54027_n1575_bF_buf3) );
  BUFX2 BUFX2_338 ( .A(u5__abc_54027_n1575), .Y(u5__abc_54027_n1575_bF_buf2) );
  BUFX2 BUFX2_339 ( .A(u5__abc_54027_n1575), .Y(u5__abc_54027_n1575_bF_buf1) );
  BUFX2 BUFX2_34 ( .A(u0_u1_lmr_req_we_FF_INPUT), .Y(u0_u1_lmr_req_we_FF_INPUT_bF_buf4) );
  BUFX2 BUFX2_340 ( .A(u5__abc_54027_n1575), .Y(u5__abc_54027_n1575_bF_buf0) );
  BUFX2 BUFX2_341 ( .A(u0_u3_init_req_we_FF_INPUT), .Y(u0_u3_init_req_we_FF_INPUT_bF_buf5) );
  BUFX2 BUFX2_342 ( .A(u0_u3_init_req_we_FF_INPUT), .Y(u0_u3_init_req_we_FF_INPUT_bF_buf4) );
  BUFX2 BUFX2_343 ( .A(u0_u3_init_req_we_FF_INPUT), .Y(u0_u3_init_req_we_FF_INPUT_bF_buf3) );
  BUFX2 BUFX2_344 ( .A(u0_u3_init_req_we_FF_INPUT), .Y(u0_u3_init_req_we_FF_INPUT_bF_buf2) );
  BUFX2 BUFX2_345 ( .A(u0_u3_init_req_we_FF_INPUT), .Y(u0_u3_init_req_we_FF_INPUT_bF_buf1) );
  BUFX2 BUFX2_346 ( .A(u0_u3_init_req_we_FF_INPUT), .Y(u0_u3_init_req_we_FF_INPUT_bF_buf0) );
  BUFX2 BUFX2_347 ( .A(page_size_10_), .Y(page_size_10_bF_buf3) );
  BUFX2 BUFX2_348 ( .A(page_size_10_), .Y(page_size_10_bF_buf2) );
  BUFX2 BUFX2_349 ( .A(page_size_10_), .Y(page_size_10_bF_buf1) );
  BUFX2 BUFX2_35 ( .A(u0_u1_lmr_req_we_FF_INPUT), .Y(u0_u1_lmr_req_we_FF_INPUT_bF_buf3) );
  BUFX2 BUFX2_350 ( .A(page_size_10_), .Y(page_size_10_bF_buf0) );
  BUFX2 BUFX2_351 ( .A(u0_u5_lmr_req_we_FF_INPUT), .Y(u0_u5_lmr_req_we_FF_INPUT_bF_buf7) );
  BUFX2 BUFX2_352 ( .A(u0_u5_lmr_req_we_FF_INPUT), .Y(u0_u5_lmr_req_we_FF_INPUT_bF_buf6) );
  BUFX2 BUFX2_353 ( .A(u0_u5_lmr_req_we_FF_INPUT), .Y(u0_u5_lmr_req_we_FF_INPUT_bF_buf5) );
  BUFX2 BUFX2_354 ( .A(u0_u5_lmr_req_we_FF_INPUT), .Y(u0_u5_lmr_req_we_FF_INPUT_bF_buf4) );
  BUFX2 BUFX2_355 ( .A(u0_u5_lmr_req_we_FF_INPUT), .Y(u0_u5_lmr_req_we_FF_INPUT_bF_buf3) );
  BUFX2 BUFX2_356 ( .A(u0_u5_lmr_req_we_FF_INPUT), .Y(u0_u5_lmr_req_we_FF_INPUT_bF_buf2) );
  BUFX2 BUFX2_357 ( .A(u0_u5_lmr_req_we_FF_INPUT), .Y(u0_u5_lmr_req_we_FF_INPUT_bF_buf1) );
  BUFX2 BUFX2_358 ( .A(u0_u5_lmr_req_we_FF_INPUT), .Y(u0_u5_lmr_req_we_FF_INPUT_bF_buf0) );
  BUFX2 BUFX2_359 ( .A(lmr_sel), .Y(lmr_sel_bF_buf6) );
  BUFX2 BUFX2_36 ( .A(u0_u1_lmr_req_we_FF_INPUT), .Y(u0_u1_lmr_req_we_FF_INPUT_bF_buf2) );
  BUFX2 BUFX2_360 ( .A(lmr_sel), .Y(lmr_sel_bF_buf5) );
  BUFX2 BUFX2_361 ( .A(lmr_sel), .Y(lmr_sel_bF_buf4) );
  BUFX2 BUFX2_362 ( .A(lmr_sel), .Y(lmr_sel_bF_buf3) );
  BUFX2 BUFX2_363 ( .A(lmr_sel), .Y(lmr_sel_bF_buf2) );
  BUFX2 BUFX2_364 ( .A(lmr_sel), .Y(lmr_sel_bF_buf1) );
  BUFX2 BUFX2_365 ( .A(lmr_sel), .Y(lmr_sel_bF_buf0) );
  BUFX2 BUFX2_366 ( .A(u0_u5__abc_45296_n218), .Y(u0_u5__abc_45296_n218_bF_buf7) );
  BUFX2 BUFX2_367 ( .A(u0_u5__abc_45296_n218), .Y(u0_u5__abc_45296_n218_bF_buf6) );
  BUFX2 BUFX2_368 ( .A(u0_u5__abc_45296_n218), .Y(u0_u5__abc_45296_n218_bF_buf5) );
  BUFX2 BUFX2_369 ( .A(u0_u5__abc_45296_n218), .Y(u0_u5__abc_45296_n218_bF_buf4) );
  BUFX2 BUFX2_37 ( .A(u0_u1_lmr_req_we_FF_INPUT), .Y(u0_u1_lmr_req_we_FF_INPUT_bF_buf1) );
  BUFX2 BUFX2_370 ( .A(u0_u5__abc_45296_n218), .Y(u0_u5__abc_45296_n218_bF_buf3) );
  BUFX2 BUFX2_371 ( .A(u0_u5__abc_45296_n218), .Y(u0_u5__abc_45296_n218_bF_buf2) );
  BUFX2 BUFX2_372 ( .A(u0_u5__abc_45296_n218), .Y(u0_u5__abc_45296_n218_bF_buf1) );
  BUFX2 BUFX2_373 ( .A(u0_u5__abc_45296_n218), .Y(u0_u5__abc_45296_n218_bF_buf0) );
  BUFX2 BUFX2_374 ( .A(row_adr_9_), .Y(row_adr_9_bF_buf6) );
  BUFX2 BUFX2_375 ( .A(row_adr_9_), .Y(row_adr_9_bF_buf5) );
  BUFX2 BUFX2_376 ( .A(row_adr_9_), .Y(row_adr_9_bF_buf4) );
  BUFX2 BUFX2_377 ( .A(row_adr_9_), .Y(row_adr_9_bF_buf3) );
  BUFX2 BUFX2_378 ( .A(row_adr_9_), .Y(row_adr_9_bF_buf2) );
  BUFX2 BUFX2_379 ( .A(row_adr_9_), .Y(row_adr_9_bF_buf1) );
  BUFX2 BUFX2_38 ( .A(u0_u1_lmr_req_we_FF_INPUT), .Y(u0_u1_lmr_req_we_FF_INPUT_bF_buf0) );
  BUFX2 BUFX2_380 ( .A(row_adr_9_), .Y(row_adr_9_bF_buf0) );
  BUFX2 BUFX2_381 ( .A(u0_u0__abc_43300_n219_1), .Y(u0_u0__abc_43300_n219_1_bF_buf4) );
  BUFX2 BUFX2_382 ( .A(u0_u0__abc_43300_n219_1), .Y(u0_u0__abc_43300_n219_1_bF_buf3) );
  BUFX2 BUFX2_383 ( .A(u0_u0__abc_43300_n219_1), .Y(u0_u0__abc_43300_n219_1_bF_buf2) );
  BUFX2 BUFX2_384 ( .A(u0_u0__abc_43300_n219_1), .Y(u0_u0__abc_43300_n219_1_bF_buf1) );
  BUFX2 BUFX2_385 ( .A(u0_u0__abc_43300_n219_1), .Y(u0_u0__abc_43300_n219_1_bF_buf0) );
  BUFX2 BUFX2_386 ( .A(row_adr_6_), .Y(row_adr_6_bF_buf6) );
  BUFX2 BUFX2_387 ( .A(row_adr_6_), .Y(row_adr_6_bF_buf5) );
  BUFX2 BUFX2_388 ( .A(row_adr_6_), .Y(row_adr_6_bF_buf4) );
  BUFX2 BUFX2_389 ( .A(row_adr_6_), .Y(row_adr_6_bF_buf3) );
  BUFX2 BUFX2_39 ( .A(rst_i), .Y(rst_i_bF_buf3) );
  BUFX2 BUFX2_390 ( .A(row_adr_6_), .Y(row_adr_6_bF_buf2) );
  BUFX2 BUFX2_391 ( .A(row_adr_6_), .Y(row_adr_6_bF_buf1) );
  BUFX2 BUFX2_392 ( .A(row_adr_6_), .Y(row_adr_6_bF_buf0) );
  BUFX2 BUFX2_393 ( .A(u3__abc_46775_n450), .Y(u3__abc_46775_n450_bF_buf3) );
  BUFX2 BUFX2_394 ( .A(u3__abc_46775_n450), .Y(u3__abc_46775_n450_bF_buf2) );
  BUFX2 BUFX2_395 ( .A(u3__abc_46775_n450), .Y(u3__abc_46775_n450_bF_buf1) );
  BUFX2 BUFX2_396 ( .A(u3__abc_46775_n450), .Y(u3__abc_46775_n450_bF_buf0) );
  BUFX2 BUFX2_397 ( .A(u3__abc_46775_n452), .Y(u3__abc_46775_n452_bF_buf3) );
  BUFX2 BUFX2_398 ( .A(u3__abc_46775_n452), .Y(u3__abc_46775_n452_bF_buf2) );
  BUFX2 BUFX2_399 ( .A(u3__abc_46775_n452), .Y(u3__abc_46775_n452_bF_buf1) );
  BUFX2 BUFX2_4 ( .A(clk_i), .Y(clk_i_hier0_bF_buf7) );
  BUFX2 BUFX2_40 ( .A(rst_i), .Y(rst_i_bF_buf2) );
  BUFX2 BUFX2_400 ( .A(u3__abc_46775_n452), .Y(u3__abc_46775_n452_bF_buf0) );
  BUFX2 BUFX2_401 ( .A(u0__abc_49347_n4304), .Y(u0__abc_49347_n4304_bF_buf4) );
  BUFX2 BUFX2_402 ( .A(u0__abc_49347_n4304), .Y(u0__abc_49347_n4304_bF_buf3) );
  BUFX2 BUFX2_403 ( .A(u0__abc_49347_n4304), .Y(u0__abc_49347_n4304_bF_buf2) );
  BUFX2 BUFX2_404 ( .A(u0__abc_49347_n4304), .Y(u0__abc_49347_n4304_bF_buf1) );
  BUFX2 BUFX2_405 ( .A(u0__abc_49347_n4304), .Y(u0__abc_49347_n4304_bF_buf0) );
  BUFX2 BUFX2_406 ( .A(u0__abc_49347_n1176_1), .Y(u0__abc_49347_n1176_1_bF_buf6) );
  BUFX2 BUFX2_407 ( .A(u0__abc_49347_n1176_1), .Y(u0__abc_49347_n1176_1_bF_buf5) );
  BUFX2 BUFX2_408 ( .A(u0__abc_49347_n1176_1), .Y(u0__abc_49347_n1176_1_bF_buf4) );
  BUFX2 BUFX2_409 ( .A(u0__abc_49347_n1176_1), .Y(u0__abc_49347_n1176_1_bF_buf3) );
  BUFX2 BUFX2_41 ( .A(rst_i), .Y(rst_i_bF_buf1) );
  BUFX2 BUFX2_410 ( .A(u0__abc_49347_n1176_1), .Y(u0__abc_49347_n1176_1_bF_buf2) );
  BUFX2 BUFX2_411 ( .A(u0__abc_49347_n1176_1), .Y(u0__abc_49347_n1176_1_bF_buf1) );
  BUFX2 BUFX2_412 ( .A(u0__abc_49347_n1176_1), .Y(u0__abc_49347_n1176_1_bF_buf0) );
  BUFX2 BUFX2_413 ( .A(u0_u0__abc_43300_n218), .Y(u0_u0__abc_43300_n218_bF_buf7) );
  BUFX2 BUFX2_414 ( .A(u0_u0__abc_43300_n218), .Y(u0_u0__abc_43300_n218_bF_buf6) );
  BUFX2 BUFX2_415 ( .A(u0_u0__abc_43300_n218), .Y(u0_u0__abc_43300_n218_bF_buf5) );
  BUFX2 BUFX2_416 ( .A(u0_u0__abc_43300_n218), .Y(u0_u0__abc_43300_n218_bF_buf4) );
  BUFX2 BUFX2_417 ( .A(u0_u0__abc_43300_n218), .Y(u0_u0__abc_43300_n218_bF_buf3) );
  BUFX2 BUFX2_418 ( .A(u0_u0__abc_43300_n218), .Y(u0_u0__abc_43300_n218_bF_buf2) );
  BUFX2 BUFX2_419 ( .A(u0_u0__abc_43300_n218), .Y(u0_u0__abc_43300_n218_bF_buf1) );
  BUFX2 BUFX2_42 ( .A(rst_i), .Y(rst_i_bF_buf0) );
  BUFX2 BUFX2_420 ( .A(u0_u0__abc_43300_n218), .Y(u0_u0__abc_43300_n218_bF_buf0) );
  BUFX2 BUFX2_421 ( .A(row_adr_3_), .Y(row_adr_3_bF_buf6) );
  BUFX2 BUFX2_422 ( .A(row_adr_3_), .Y(row_adr_3_bF_buf5) );
  BUFX2 BUFX2_423 ( .A(row_adr_3_), .Y(row_adr_3_bF_buf4) );
  BUFX2 BUFX2_424 ( .A(row_adr_3_), .Y(row_adr_3_bF_buf3) );
  BUFX2 BUFX2_425 ( .A(row_adr_3_), .Y(row_adr_3_bF_buf2) );
  BUFX2 BUFX2_426 ( .A(row_adr_3_), .Y(row_adr_3_bF_buf1) );
  BUFX2 BUFX2_427 ( .A(row_adr_3_), .Y(row_adr_3_bF_buf0) );
  BUFX2 BUFX2_428 ( .A(cs_le), .Y(cs_le_bF_buf4) );
  BUFX2 BUFX2_429 ( .A(cs_le), .Y(cs_le_bF_buf3) );
  BUFX2 BUFX2_43 ( .A(u0_u1__abc_43657_n219_1), .Y(u0_u1__abc_43657_n219_1_bF_buf7) );
  BUFX2 BUFX2_430 ( .A(cs_le), .Y(cs_le_bF_buf2) );
  BUFX2 BUFX2_431 ( .A(cs_le), .Y(cs_le_bF_buf1) );
  BUFX2 BUFX2_432 ( .A(cs_le), .Y(cs_le_bF_buf0) );
  BUFX2 BUFX2_433 ( .A(u0__abc_49347_n2748), .Y(u0__abc_49347_n2748_bF_buf5) );
  BUFX2 BUFX2_434 ( .A(u0__abc_49347_n2748), .Y(u0__abc_49347_n2748_bF_buf4) );
  BUFX2 BUFX2_435 ( .A(u0__abc_49347_n2748), .Y(u0__abc_49347_n2748_bF_buf3) );
  BUFX2 BUFX2_436 ( .A(u0__abc_49347_n2748), .Y(u0__abc_49347_n2748_bF_buf2) );
  BUFX2 BUFX2_437 ( .A(u0__abc_49347_n2748), .Y(u0__abc_49347_n2748_bF_buf1) );
  BUFX2 BUFX2_438 ( .A(u0__abc_49347_n2748), .Y(u0__abc_49347_n2748_bF_buf0) );
  BUFX2 BUFX2_439 ( .A(csc_s_5_), .Y(csc_s_5_bF_buf4) );
  BUFX2 BUFX2_44 ( .A(u0_u1__abc_43657_n219_1), .Y(u0_u1__abc_43657_n219_1_bF_buf6) );
  BUFX2 BUFX2_440 ( .A(csc_s_5_), .Y(csc_s_5_bF_buf3) );
  BUFX2 BUFX2_441 ( .A(csc_s_5_), .Y(csc_s_5_bF_buf2) );
  BUFX2 BUFX2_442 ( .A(csc_s_5_), .Y(csc_s_5_bF_buf1) );
  BUFX2 BUFX2_443 ( .A(csc_s_5_), .Y(csc_s_5_bF_buf0) );
  BUFX2 BUFX2_444 ( .A(row_adr_0_), .Y(row_adr_0_bF_buf6) );
  BUFX2 BUFX2_445 ( .A(row_adr_0_), .Y(row_adr_0_bF_buf5) );
  BUFX2 BUFX2_446 ( .A(row_adr_0_), .Y(row_adr_0_bF_buf4) );
  BUFX2 BUFX2_447 ( .A(row_adr_0_), .Y(row_adr_0_bF_buf3) );
  BUFX2 BUFX2_448 ( .A(row_adr_0_), .Y(row_adr_0_bF_buf2) );
  BUFX2 BUFX2_449 ( .A(row_adr_0_), .Y(row_adr_0_bF_buf1) );
  BUFX2 BUFX2_45 ( .A(u0_u1__abc_43657_n219_1), .Y(u0_u1__abc_43657_n219_1_bF_buf5) );
  BUFX2 BUFX2_450 ( .A(row_adr_0_), .Y(row_adr_0_bF_buf0) );
  BUFX2 BUFX2_451 ( .A(next_adr), .Y(next_adr_bF_buf4) );
  BUFX2 BUFX2_452 ( .A(next_adr), .Y(next_adr_bF_buf3) );
  BUFX2 BUFX2_453 ( .A(next_adr), .Y(next_adr_bF_buf2) );
  BUFX2 BUFX2_454 ( .A(next_adr), .Y(next_adr_bF_buf1) );
  BUFX2 BUFX2_455 ( .A(next_adr), .Y(next_adr_bF_buf0) );
  BUFX2 BUFX2_456 ( .A(u5__abc_54027_n565), .Y(u5__abc_54027_n565_bF_buf4) );
  BUFX2 BUFX2_457 ( .A(u5__abc_54027_n565), .Y(u5__abc_54027_n565_bF_buf3) );
  BUFX2 BUFX2_458 ( .A(u5__abc_54027_n565), .Y(u5__abc_54027_n565_bF_buf2) );
  BUFX2 BUFX2_459 ( .A(u5__abc_54027_n565), .Y(u5__abc_54027_n565_bF_buf1) );
  BUFX2 BUFX2_46 ( .A(u0_u1__abc_43657_n219_1), .Y(u0_u1__abc_43657_n219_1_bF_buf4) );
  BUFX2 BUFX2_460 ( .A(u5__abc_54027_n565), .Y(u5__abc_54027_n565_bF_buf0) );
  BUFX2 BUFX2_461 ( .A(u4__abc_49152_n191), .Y(u4__abc_49152_n191_bF_buf3) );
  BUFX2 BUFX2_462 ( .A(u4__abc_49152_n191), .Y(u4__abc_49152_n191_bF_buf2) );
  BUFX2 BUFX2_463 ( .A(u4__abc_49152_n191), .Y(u4__abc_49152_n191_bF_buf1) );
  BUFX2 BUFX2_464 ( .A(u4__abc_49152_n191), .Y(u4__abc_49152_n191_bF_buf0) );
  BUFX2 BUFX2_465 ( .A(bank_adr_0_), .Y(bank_adr_0_bF_buf3) );
  BUFX2 BUFX2_466 ( .A(bank_adr_0_), .Y(bank_adr_0_bF_buf2) );
  BUFX2 BUFX2_467 ( .A(bank_adr_0_), .Y(bank_adr_0_bF_buf1) );
  BUFX2 BUFX2_468 ( .A(bank_adr_0_), .Y(bank_adr_0_bF_buf0) );
  BUFX2 BUFX2_469 ( .A(\wb_addr_i[23] ), .Y(wb_addr_i_23_bF_buf3) );
  BUFX2 BUFX2_47 ( .A(u0_u1__abc_43657_n219_1), .Y(u0_u1__abc_43657_n219_1_bF_buf3) );
  BUFX2 BUFX2_470 ( .A(\wb_addr_i[23] ), .Y(wb_addr_i_23_bF_buf2) );
  BUFX2 BUFX2_471 ( .A(\wb_addr_i[23] ), .Y(wb_addr_i_23_bF_buf1) );
  BUFX2 BUFX2_472 ( .A(\wb_addr_i[23] ), .Y(wb_addr_i_23_bF_buf0) );
  BUFX2 BUFX2_473 ( .A(csc_s_2_), .Y(csc_s_2_bF_buf4) );
  BUFX2 BUFX2_474 ( .A(csc_s_2_), .Y(csc_s_2_bF_buf3) );
  BUFX2 BUFX2_475 ( .A(csc_s_2_), .Y(csc_s_2_bF_buf2) );
  BUFX2 BUFX2_476 ( .A(csc_s_2_), .Y(csc_s_2_bF_buf1) );
  BUFX2 BUFX2_477 ( .A(csc_s_2_), .Y(csc_s_2_bF_buf0) );
  BUFX2 BUFX2_478 ( .A(u1__abc_45852_n276), .Y(u1__abc_45852_n276_bF_buf4) );
  BUFX2 BUFX2_479 ( .A(u1__abc_45852_n276), .Y(u1__abc_45852_n276_bF_buf3) );
  BUFX2 BUFX2_48 ( .A(u0_u1__abc_43657_n219_1), .Y(u0_u1__abc_43657_n219_1_bF_buf2) );
  BUFX2 BUFX2_480 ( .A(u1__abc_45852_n276), .Y(u1__abc_45852_n276_bF_buf2) );
  BUFX2 BUFX2_481 ( .A(u1__abc_45852_n276), .Y(u1__abc_45852_n276_bF_buf1) );
  BUFX2 BUFX2_482 ( .A(u1__abc_45852_n276), .Y(u1__abc_45852_n276_bF_buf0) );
  BUFX2 BUFX2_483 ( .A(u2_u4__abc_47660_n137), .Y(u2_u4__abc_47660_n137_bF_buf4) );
  BUFX2 BUFX2_484 ( .A(u2_u4__abc_47660_n137), .Y(u2_u4__abc_47660_n137_bF_buf3) );
  BUFX2 BUFX2_485 ( .A(u2_u4__abc_47660_n137), .Y(u2_u4__abc_47660_n137_bF_buf2) );
  BUFX2 BUFX2_486 ( .A(u2_u4__abc_47660_n137), .Y(u2_u4__abc_47660_n137_bF_buf1) );
  BUFX2 BUFX2_487 ( .A(u2_u4__abc_47660_n137), .Y(u2_u4__abc_47660_n137_bF_buf0) );
  BUFX2 BUFX2_488 ( .A(u0_u2__abc_44109_n209), .Y(u0_u2__abc_44109_n209_bF_buf7) );
  BUFX2 BUFX2_489 ( .A(u0_u2__abc_44109_n209), .Y(u0_u2__abc_44109_n209_bF_buf6) );
  BUFX2 BUFX2_49 ( .A(u0_u1__abc_43657_n219_1), .Y(u0_u1__abc_43657_n219_1_bF_buf1) );
  BUFX2 BUFX2_490 ( .A(u0_u2__abc_44109_n209), .Y(u0_u2__abc_44109_n209_bF_buf5) );
  BUFX2 BUFX2_491 ( .A(u0_u2__abc_44109_n209), .Y(u0_u2__abc_44109_n209_bF_buf4) );
  BUFX2 BUFX2_492 ( .A(u0_u2__abc_44109_n209), .Y(u0_u2__abc_44109_n209_bF_buf3) );
  BUFX2 BUFX2_493 ( .A(u0_u2__abc_44109_n209), .Y(u0_u2__abc_44109_n209_bF_buf2) );
  BUFX2 BUFX2_494 ( .A(u0_u2__abc_44109_n209), .Y(u0_u2__abc_44109_n209_bF_buf1) );
  BUFX2 BUFX2_495 ( .A(u0_u2__abc_44109_n209), .Y(u0_u2__abc_44109_n209_bF_buf0) );
  BUFX2 BUFX2_496 ( .A(u0__abc_49347_n4560), .Y(u0__abc_49347_n4560_bF_buf4) );
  BUFX2 BUFX2_497 ( .A(u0__abc_49347_n4560), .Y(u0__abc_49347_n4560_bF_buf3) );
  BUFX2 BUFX2_498 ( .A(u0__abc_49347_n4560), .Y(u0__abc_49347_n4560_bF_buf2) );
  BUFX2 BUFX2_499 ( .A(u0__abc_49347_n4560), .Y(u0__abc_49347_n4560_bF_buf1) );
  BUFX2 BUFX2_5 ( .A(clk_i), .Y(clk_i_hier0_bF_buf6) );
  BUFX2 BUFX2_50 ( .A(u0_u1__abc_43657_n219_1), .Y(u0_u1__abc_43657_n219_1_bF_buf0) );
  BUFX2 BUFX2_500 ( .A(u0__abc_49347_n4560), .Y(u0__abc_49347_n4560_bF_buf0) );
  BUFX2 BUFX2_501 ( .A(u0__abc_49347_n4562), .Y(u0__abc_49347_n4562_bF_buf4) );
  BUFX2 BUFX2_502 ( .A(u0__abc_49347_n4562), .Y(u0__abc_49347_n4562_bF_buf3) );
  BUFX2 BUFX2_503 ( .A(u0__abc_49347_n4562), .Y(u0__abc_49347_n4562_bF_buf2) );
  BUFX2 BUFX2_504 ( .A(u0__abc_49347_n4562), .Y(u0__abc_49347_n4562_bF_buf1) );
  BUFX2 BUFX2_505 ( .A(u0__abc_49347_n4562), .Y(u0__abc_49347_n4562_bF_buf0) );
  BUFX2 BUFX2_506 ( .A(u0__abc_49347_n4567), .Y(u0__abc_49347_n4567_bF_buf4) );
  BUFX2 BUFX2_507 ( .A(u0__abc_49347_n4567), .Y(u0__abc_49347_n4567_bF_buf3) );
  BUFX2 BUFX2_508 ( .A(u0__abc_49347_n4567), .Y(u0__abc_49347_n4567_bF_buf2) );
  BUFX2 BUFX2_509 ( .A(u0__abc_49347_n4567), .Y(u0__abc_49347_n4567_bF_buf1) );
  BUFX2 BUFX2_51 ( .A(row_adr_7_), .Y(row_adr_7_bF_buf6) );
  BUFX2 BUFX2_510 ( .A(u0__abc_49347_n4567), .Y(u0__abc_49347_n4567_bF_buf0) );
  BUFX2 BUFX2_511 ( .A(u3_u0__abc_48231_n1050), .Y(u3_u0__abc_48231_n1050_bF_buf5) );
  BUFX2 BUFX2_512 ( .A(u3_u0__abc_48231_n1050), .Y(u3_u0__abc_48231_n1050_bF_buf4) );
  BUFX2 BUFX2_513 ( .A(u3_u0__abc_48231_n1050), .Y(u3_u0__abc_48231_n1050_bF_buf3) );
  BUFX2 BUFX2_514 ( .A(u3_u0__abc_48231_n1050), .Y(u3_u0__abc_48231_n1050_bF_buf2) );
  BUFX2 BUFX2_515 ( .A(u3_u0__abc_48231_n1050), .Y(u3_u0__abc_48231_n1050_bF_buf1) );
  BUFX2 BUFX2_516 ( .A(u3_u0__abc_48231_n1050), .Y(u3_u0__abc_48231_n1050_bF_buf0) );
  BUFX2 BUFX2_517 ( .A(u0_cs0), .Y(u0_cs0_bF_buf5) );
  BUFX2 BUFX2_518 ( .A(u0_cs0), .Y(u0_cs0_bF_buf4) );
  BUFX2 BUFX2_519 ( .A(u0_cs0), .Y(u0_cs0_bF_buf3) );
  BUFX2 BUFX2_52 ( .A(row_adr_7_), .Y(row_adr_7_bF_buf5) );
  BUFX2 BUFX2_520 ( .A(u0_cs0), .Y(u0_cs0_bF_buf2) );
  BUFX2 BUFX2_521 ( .A(u0_cs0), .Y(u0_cs0_bF_buf1) );
  BUFX2 BUFX2_522 ( .A(u0_cs0), .Y(u0_cs0_bF_buf0) );
  BUFX2 BUFX2_523 ( .A(u0_cs1), .Y(u0_cs1_bF_buf5) );
  BUFX2 BUFX2_524 ( .A(u0_cs1), .Y(u0_cs1_bF_buf4) );
  BUFX2 BUFX2_525 ( .A(u0_cs1), .Y(u0_cs1_bF_buf3) );
  BUFX2 BUFX2_526 ( .A(u0_cs1), .Y(u0_cs1_bF_buf2) );
  BUFX2 BUFX2_527 ( .A(u0_cs1), .Y(u0_cs1_bF_buf1) );
  BUFX2 BUFX2_528 ( .A(u0_cs1), .Y(u0_cs1_bF_buf0) );
  BUFX2 BUFX2_529 ( .A(u0_cs2), .Y(u0_cs2_bF_buf5) );
  BUFX2 BUFX2_53 ( .A(row_adr_7_), .Y(row_adr_7_bF_buf4) );
  BUFX2 BUFX2_530 ( .A(u0_cs2), .Y(u0_cs2_bF_buf4) );
  BUFX2 BUFX2_531 ( .A(u0_cs2), .Y(u0_cs2_bF_buf3) );
  BUFX2 BUFX2_532 ( .A(u0_cs2), .Y(u0_cs2_bF_buf2) );
  BUFX2 BUFX2_533 ( .A(u0_cs2), .Y(u0_cs2_bF_buf1) );
  BUFX2 BUFX2_534 ( .A(u0_cs2), .Y(u0_cs2_bF_buf0) );
  BUFX2 BUFX2_535 ( .A(u0_cs3), .Y(u0_cs3_bF_buf5) );
  BUFX2 BUFX2_536 ( .A(u0_cs3), .Y(u0_cs3_bF_buf4) );
  BUFX2 BUFX2_537 ( .A(u0_cs3), .Y(u0_cs3_bF_buf3) );
  BUFX2 BUFX2_538 ( .A(u0_cs3), .Y(u0_cs3_bF_buf2) );
  BUFX2 BUFX2_539 ( .A(u0_cs3), .Y(u0_cs3_bF_buf1) );
  BUFX2 BUFX2_54 ( .A(row_adr_7_), .Y(row_adr_7_bF_buf3) );
  BUFX2 BUFX2_540 ( .A(u0_cs3), .Y(u0_cs3_bF_buf0) );
  BUFX2 BUFX2_541 ( .A(u0_cs4), .Y(u0_cs4_bF_buf5) );
  BUFX2 BUFX2_542 ( .A(u0_cs4), .Y(u0_cs4_bF_buf4) );
  BUFX2 BUFX2_543 ( .A(u0_cs4), .Y(u0_cs4_bF_buf3) );
  BUFX2 BUFX2_544 ( .A(u0_cs4), .Y(u0_cs4_bF_buf2) );
  BUFX2 BUFX2_545 ( .A(u0_cs4), .Y(u0_cs4_bF_buf1) );
  BUFX2 BUFX2_546 ( .A(u0_cs4), .Y(u0_cs4_bF_buf0) );
  BUFX2 BUFX2_547 ( .A(u0_cs5), .Y(u0_cs5_bF_buf5) );
  BUFX2 BUFX2_548 ( .A(u0_cs5), .Y(u0_cs5_bF_buf4) );
  BUFX2 BUFX2_549 ( .A(u0_cs5), .Y(u0_cs5_bF_buf3) );
  BUFX2 BUFX2_55 ( .A(row_adr_7_), .Y(row_adr_7_bF_buf2) );
  BUFX2 BUFX2_550 ( .A(u0_cs5), .Y(u0_cs5_bF_buf2) );
  BUFX2 BUFX2_551 ( .A(u0_cs5), .Y(u0_cs5_bF_buf1) );
  BUFX2 BUFX2_552 ( .A(u0_cs5), .Y(u0_cs5_bF_buf0) );
  BUFX2 BUFX2_553 ( .A(row_adr_12_), .Y(row_adr_12_bF_buf6) );
  BUFX2 BUFX2_554 ( .A(row_adr_12_), .Y(row_adr_12_bF_buf5) );
  BUFX2 BUFX2_555 ( .A(row_adr_12_), .Y(row_adr_12_bF_buf4) );
  BUFX2 BUFX2_556 ( .A(row_adr_12_), .Y(row_adr_12_bF_buf3) );
  BUFX2 BUFX2_557 ( .A(row_adr_12_), .Y(row_adr_12_bF_buf2) );
  BUFX2 BUFX2_558 ( .A(row_adr_12_), .Y(row_adr_12_bF_buf1) );
  BUFX2 BUFX2_559 ( .A(row_adr_12_), .Y(row_adr_12_bF_buf0) );
  BUFX2 BUFX2_56 ( .A(row_adr_7_), .Y(row_adr_7_bF_buf1) );
  BUFX2 BUFX2_560 ( .A(u0__abc_49347_n4531), .Y(u0__abc_49347_n4531_bF_buf4) );
  BUFX2 BUFX2_561 ( .A(u0__abc_49347_n4531), .Y(u0__abc_49347_n4531_bF_buf3) );
  BUFX2 BUFX2_562 ( .A(u0__abc_49347_n4531), .Y(u0__abc_49347_n4531_bF_buf2) );
  BUFX2 BUFX2_563 ( .A(u0__abc_49347_n4531), .Y(u0__abc_49347_n4531_bF_buf1) );
  BUFX2 BUFX2_564 ( .A(u0__abc_49347_n4531), .Y(u0__abc_49347_n4531_bF_buf0) );
  BUFX2 BUFX2_565 ( .A(u0__abc_49347_n4535), .Y(u0__abc_49347_n4535_bF_buf4) );
  BUFX2 BUFX2_566 ( .A(u0__abc_49347_n4535), .Y(u0__abc_49347_n4535_bF_buf3) );
  BUFX2 BUFX2_567 ( .A(u0__abc_49347_n4535), .Y(u0__abc_49347_n4535_bF_buf2) );
  BUFX2 BUFX2_568 ( .A(u0__abc_49347_n4535), .Y(u0__abc_49347_n4535_bF_buf1) );
  BUFX2 BUFX2_569 ( .A(u0__abc_49347_n4535), .Y(u0__abc_49347_n4535_bF_buf0) );
  BUFX2 BUFX2_57 ( .A(row_adr_7_), .Y(row_adr_7_bF_buf0) );
  BUFX2 BUFX2_570 ( .A(u0__abc_49347_n4537), .Y(u0__abc_49347_n4537_bF_buf4) );
  BUFX2 BUFX2_571 ( .A(u0__abc_49347_n4537), .Y(u0__abc_49347_n4537_bF_buf3) );
  BUFX2 BUFX2_572 ( .A(u0__abc_49347_n4537), .Y(u0__abc_49347_n4537_bF_buf2) );
  BUFX2 BUFX2_573 ( .A(u0__abc_49347_n4537), .Y(u0__abc_49347_n4537_bF_buf1) );
  BUFX2 BUFX2_574 ( .A(u0__abc_49347_n4537), .Y(u0__abc_49347_n4537_bF_buf0) );
  BUFX2 BUFX2_575 ( .A(u0__abc_49347_n4539), .Y(u0__abc_49347_n4539_bF_buf4) );
  BUFX2 BUFX2_576 ( .A(u0__abc_49347_n4539), .Y(u0__abc_49347_n4539_bF_buf3) );
  BUFX2 BUFX2_577 ( .A(u0__abc_49347_n4539), .Y(u0__abc_49347_n4539_bF_buf2) );
  BUFX2 BUFX2_578 ( .A(u0__abc_49347_n4539), .Y(u0__abc_49347_n4539_bF_buf1) );
  BUFX2 BUFX2_579 ( .A(u0__abc_49347_n4539), .Y(u0__abc_49347_n4539_bF_buf0) );
  BUFX2 BUFX2_58 ( .A(u0_u0_lmr_req_we_FF_INPUT), .Y(u0_u0_lmr_req_we_FF_INPUT_bF_buf4) );
  BUFX2 BUFX2_580 ( .A(u0__abc_49347_n3188), .Y(u0__abc_49347_n3188_bF_buf10) );
  BUFX2 BUFX2_581 ( .A(u0__abc_49347_n3188), .Y(u0__abc_49347_n3188_bF_buf9) );
  BUFX2 BUFX2_582 ( .A(u0__abc_49347_n3188), .Y(u0__abc_49347_n3188_bF_buf8) );
  BUFX2 BUFX2_583 ( .A(u0__abc_49347_n3188), .Y(u0__abc_49347_n3188_bF_buf7) );
  BUFX2 BUFX2_584 ( .A(u0__abc_49347_n3188), .Y(u0__abc_49347_n3188_bF_buf6) );
  BUFX2 BUFX2_585 ( .A(u0__abc_49347_n3188), .Y(u0__abc_49347_n3188_bF_buf5) );
  BUFX2 BUFX2_586 ( .A(u0__abc_49347_n3188), .Y(u0__abc_49347_n3188_bF_buf4) );
  BUFX2 BUFX2_587 ( .A(u0__abc_49347_n3188), .Y(u0__abc_49347_n3188_bF_buf3) );
  BUFX2 BUFX2_588 ( .A(u0__abc_49347_n3188), .Y(u0__abc_49347_n3188_bF_buf2) );
  BUFX2 BUFX2_589 ( .A(u0__abc_49347_n3188), .Y(u0__abc_49347_n3188_bF_buf1) );
  BUFX2 BUFX2_59 ( .A(u0_u0_lmr_req_we_FF_INPUT), .Y(u0_u0_lmr_req_we_FF_INPUT_bF_buf3) );
  BUFX2 BUFX2_590 ( .A(u0__abc_49347_n3188), .Y(u0__abc_49347_n3188_bF_buf0) );
  BUFX2 BUFX2_591 ( .A(u0_u2__abc_44109_n210_1), .Y(u0_u2__abc_44109_n210_1_bF_buf4) );
  BUFX2 BUFX2_592 ( .A(u0_u2__abc_44109_n210_1), .Y(u0_u2__abc_44109_n210_1_bF_buf3) );
  BUFX2 BUFX2_593 ( .A(u0_u2__abc_44109_n210_1), .Y(u0_u2__abc_44109_n210_1_bF_buf2) );
  BUFX2 BUFX2_594 ( .A(u0_u2__abc_44109_n210_1), .Y(u0_u2__abc_44109_n210_1_bF_buf1) );
  BUFX2 BUFX2_595 ( .A(u0_u2__abc_44109_n210_1), .Y(u0_u2__abc_44109_n210_1_bF_buf0) );
  BUFX2 BUFX2_596 ( .A(spec_req_cs_4_), .Y(spec_req_cs_4_bF_buf5) );
  BUFX2 BUFX2_597 ( .A(spec_req_cs_4_), .Y(spec_req_cs_4_bF_buf4) );
  BUFX2 BUFX2_598 ( .A(spec_req_cs_4_), .Y(spec_req_cs_4_bF_buf3) );
  BUFX2 BUFX2_599 ( .A(spec_req_cs_4_), .Y(spec_req_cs_4_bF_buf2) );
  BUFX2 BUFX2_6 ( .A(clk_i), .Y(clk_i_hier0_bF_buf5) );
  BUFX2 BUFX2_60 ( .A(u0_u0_lmr_req_we_FF_INPUT), .Y(u0_u0_lmr_req_we_FF_INPUT_bF_buf2) );
  BUFX2 BUFX2_600 ( .A(spec_req_cs_4_), .Y(spec_req_cs_4_bF_buf1) );
  BUFX2 BUFX2_601 ( .A(spec_req_cs_4_), .Y(spec_req_cs_4_bF_buf0) );
  BUFX2 BUFX2_602 ( .A(u3__abc_46775_n275), .Y(u3__abc_46775_n275_bF_buf4) );
  BUFX2 BUFX2_603 ( .A(u3__abc_46775_n275), .Y(u3__abc_46775_n275_bF_buf3) );
  BUFX2 BUFX2_604 ( .A(u3__abc_46775_n275), .Y(u3__abc_46775_n275_bF_buf2) );
  BUFX2 BUFX2_605 ( .A(u3__abc_46775_n275), .Y(u3__abc_46775_n275_bF_buf1) );
  BUFX2 BUFX2_606 ( .A(u3__abc_46775_n275), .Y(u3__abc_46775_n275_bF_buf0) );
  BUFX2 BUFX2_607 ( .A(u3__abc_46775_n279), .Y(u3__abc_46775_n279_bF_buf5) );
  BUFX2 BUFX2_608 ( .A(u3__abc_46775_n279), .Y(u3__abc_46775_n279_bF_buf4) );
  BUFX2 BUFX2_609 ( .A(u3__abc_46775_n279), .Y(u3__abc_46775_n279_bF_buf3) );
  BUFX2 BUFX2_61 ( .A(u0_u0_lmr_req_we_FF_INPUT), .Y(u0_u0_lmr_req_we_FF_INPUT_bF_buf1) );
  BUFX2 BUFX2_610 ( .A(u3__abc_46775_n279), .Y(u3__abc_46775_n279_bF_buf2) );
  BUFX2 BUFX2_611 ( .A(u3__abc_46775_n279), .Y(u3__abc_46775_n279_bF_buf1) );
  BUFX2 BUFX2_612 ( .A(u3__abc_46775_n279), .Y(u3__abc_46775_n279_bF_buf0) );
  BUFX2 BUFX2_613 ( .A(u1__abc_45852_n562), .Y(u1__abc_45852_n562_bF_buf3) );
  BUFX2 BUFX2_614 ( .A(u1__abc_45852_n562), .Y(u1__abc_45852_n562_bF_buf2) );
  BUFX2 BUFX2_615 ( .A(u1__abc_45852_n562), .Y(u1__abc_45852_n562_bF_buf1) );
  BUFX2 BUFX2_616 ( .A(u1__abc_45852_n562), .Y(u1__abc_45852_n562_bF_buf0) );
  BUFX2 BUFX2_617 ( .A(u0_u4_init_req_we_FF_INPUT), .Y(u0_u4_init_req_we_FF_INPUT_bF_buf7) );
  BUFX2 BUFX2_618 ( .A(u0_u4_init_req_we_FF_INPUT), .Y(u0_u4_init_req_we_FF_INPUT_bF_buf6) );
  BUFX2 BUFX2_619 ( .A(u0_u4_init_req_we_FF_INPUT), .Y(u0_u4_init_req_we_FF_INPUT_bF_buf5) );
  BUFX2 BUFX2_62 ( .A(u0_u0_lmr_req_we_FF_INPUT), .Y(u0_u0_lmr_req_we_FF_INPUT_bF_buf0) );
  BUFX2 BUFX2_620 ( .A(u0_u4_init_req_we_FF_INPUT), .Y(u0_u4_init_req_we_FF_INPUT_bF_buf4) );
  BUFX2 BUFX2_621 ( .A(u0_u4_init_req_we_FF_INPUT), .Y(u0_u4_init_req_we_FF_INPUT_bF_buf3) );
  BUFX2 BUFX2_622 ( .A(u0_u4_init_req_we_FF_INPUT), .Y(u0_u4_init_req_we_FF_INPUT_bF_buf2) );
  BUFX2 BUFX2_623 ( .A(u0_u4_init_req_we_FF_INPUT), .Y(u0_u4_init_req_we_FF_INPUT_bF_buf1) );
  BUFX2 BUFX2_624 ( .A(u0_u4_init_req_we_FF_INPUT), .Y(u0_u4_init_req_we_FF_INPUT_bF_buf0) );
  BUFX2 BUFX2_625 ( .A(u2_u2__abc_47660_n137), .Y(u2_u2__abc_47660_n137_bF_buf4) );
  BUFX2 BUFX2_626 ( .A(u2_u2__abc_47660_n137), .Y(u2_u2__abc_47660_n137_bF_buf3) );
  BUFX2 BUFX2_627 ( .A(u2_u2__abc_47660_n137), .Y(u2_u2__abc_47660_n137_bF_buf2) );
  BUFX2 BUFX2_628 ( .A(u2_u2__abc_47660_n137), .Y(u2_u2__abc_47660_n137_bF_buf1) );
  BUFX2 BUFX2_629 ( .A(u2_u2__abc_47660_n137), .Y(u2_u2__abc_47660_n137_bF_buf0) );
  BUFX2 BUFX2_63 ( .A(u3_u0__abc_48231_n708), .Y(u3_u0__abc_48231_n708_bF_buf7) );
  BUFX2 BUFX2_630 ( .A(u0__abc_49347_n1952_1), .Y(u0__abc_49347_n1952_1_bF_buf3) );
  BUFX2 BUFX2_631 ( .A(u0__abc_49347_n1952_1), .Y(u0__abc_49347_n1952_1_bF_buf2) );
  BUFX2 BUFX2_632 ( .A(u0__abc_49347_n1952_1), .Y(u0__abc_49347_n1952_1_bF_buf1) );
  BUFX2 BUFX2_633 ( .A(u0__abc_49347_n1952_1), .Y(u0__abc_49347_n1952_1_bF_buf0) );
  BUFX2 BUFX2_634 ( .A(u0__abc_49347_n4507), .Y(u0__abc_49347_n4507_bF_buf3) );
  BUFX2 BUFX2_635 ( .A(u0__abc_49347_n4507), .Y(u0__abc_49347_n4507_bF_buf2) );
  BUFX2 BUFX2_636 ( .A(u0__abc_49347_n4507), .Y(u0__abc_49347_n4507_bF_buf1) );
  BUFX2 BUFX2_637 ( .A(u0__abc_49347_n4507), .Y(u0__abc_49347_n4507_bF_buf0) );
  BUFX2 BUFX2_638 ( .A(u0__abc_49347_n1178_1), .Y(u0__abc_49347_n1178_1_bF_buf5) );
  BUFX2 BUFX2_639 ( .A(u0__abc_49347_n1178_1), .Y(u0__abc_49347_n1178_1_bF_buf4) );
  BUFX2 BUFX2_64 ( .A(u3_u0__abc_48231_n708), .Y(u3_u0__abc_48231_n708_bF_buf6) );
  BUFX2 BUFX2_640 ( .A(u0__abc_49347_n1178_1), .Y(u0__abc_49347_n1178_1_bF_buf3) );
  BUFX2 BUFX2_641 ( .A(u0__abc_49347_n1178_1), .Y(u0__abc_49347_n1178_1_bF_buf2) );
  BUFX2 BUFX2_642 ( .A(u0__abc_49347_n1178_1), .Y(u0__abc_49347_n1178_1_bF_buf1) );
  BUFX2 BUFX2_643 ( .A(u0__abc_49347_n1178_1), .Y(u0__abc_49347_n1178_1_bF_buf0) );
  BUFX2 BUFX2_644 ( .A(u0_u4__abc_44844_n209_1), .Y(u0_u4__abc_44844_n209_1_bF_buf7) );
  BUFX2 BUFX2_645 ( .A(u0_u4__abc_44844_n209_1), .Y(u0_u4__abc_44844_n209_1_bF_buf6) );
  BUFX2 BUFX2_646 ( .A(u0_u4__abc_44844_n209_1), .Y(u0_u4__abc_44844_n209_1_bF_buf5) );
  BUFX2 BUFX2_647 ( .A(u0_u4__abc_44844_n209_1), .Y(u0_u4__abc_44844_n209_1_bF_buf4) );
  BUFX2 BUFX2_648 ( .A(u0_u4__abc_44844_n209_1), .Y(u0_u4__abc_44844_n209_1_bF_buf3) );
  BUFX2 BUFX2_649 ( .A(u0_u4__abc_44844_n209_1), .Y(u0_u4__abc_44844_n209_1_bF_buf2) );
  BUFX2 BUFX2_65 ( .A(u3_u0__abc_48231_n708), .Y(u3_u0__abc_48231_n708_bF_buf5) );
  BUFX2 BUFX2_650 ( .A(u0_u4__abc_44844_n209_1), .Y(u0_u4__abc_44844_n209_1_bF_buf1) );
  BUFX2 BUFX2_651 ( .A(u0_u4__abc_44844_n209_1), .Y(u0_u4__abc_44844_n209_1_bF_buf0) );
  BUFX2 BUFX2_652 ( .A(u0_u0_init_req_we_FF_INPUT), .Y(u0_u0_init_req_we_FF_INPUT_bF_buf4) );
  BUFX2 BUFX2_653 ( .A(u0_u0_init_req_we_FF_INPUT), .Y(u0_u0_init_req_we_FF_INPUT_bF_buf3) );
  BUFX2 BUFX2_654 ( .A(u0_u0_init_req_we_FF_INPUT), .Y(u0_u0_init_req_we_FF_INPUT_bF_buf2) );
  BUFX2 BUFX2_655 ( .A(u0_u0_init_req_we_FF_INPUT), .Y(u0_u0_init_req_we_FF_INPUT_bF_buf1) );
  BUFX2 BUFX2_656 ( .A(u0_u0_init_req_we_FF_INPUT), .Y(u0_u0_init_req_we_FF_INPUT_bF_buf0) );
  BUFX2 BUFX2_657 ( .A(spec_req_cs_1_), .Y(spec_req_cs_1_bF_buf5) );
  BUFX2 BUFX2_658 ( .A(spec_req_cs_1_), .Y(spec_req_cs_1_bF_buf4) );
  BUFX2 BUFX2_659 ( .A(spec_req_cs_1_), .Y(spec_req_cs_1_bF_buf3) );
  BUFX2 BUFX2_66 ( .A(u3_u0__abc_48231_n708), .Y(u3_u0__abc_48231_n708_bF_buf4) );
  BUFX2 BUFX2_660 ( .A(spec_req_cs_1_), .Y(spec_req_cs_1_bF_buf2) );
  BUFX2 BUFX2_661 ( .A(spec_req_cs_1_), .Y(spec_req_cs_1_bF_buf1) );
  BUFX2 BUFX2_662 ( .A(spec_req_cs_1_), .Y(spec_req_cs_1_bF_buf0) );
  BUFX2 BUFX2_663 ( .A(u3__abc_46775_n625), .Y(u3__abc_46775_n625_bF_buf4) );
  BUFX2 BUFX2_664 ( .A(u3__abc_46775_n625), .Y(u3__abc_46775_n625_bF_buf3) );
  BUFX2 BUFX2_665 ( .A(u3__abc_46775_n625), .Y(u3__abc_46775_n625_bF_buf2) );
  BUFX2 BUFX2_666 ( .A(u3__abc_46775_n625), .Y(u3__abc_46775_n625_bF_buf1) );
  BUFX2 BUFX2_667 ( .A(u3__abc_46775_n625), .Y(u3__abc_46775_n625_bF_buf0) );
  BUFX2 BUFX2_668 ( .A(u0__abc_49347_n4443), .Y(u0__abc_49347_n4443_bF_buf3) );
  BUFX2 BUFX2_669 ( .A(u0__abc_49347_n4443), .Y(u0__abc_49347_n4443_bF_buf2) );
  BUFX2 BUFX2_67 ( .A(u3_u0__abc_48231_n708), .Y(u3_u0__abc_48231_n708_bF_buf3) );
  BUFX2 BUFX2_670 ( .A(u0__abc_49347_n4443), .Y(u0__abc_49347_n4443_bF_buf1) );
  BUFX2 BUFX2_671 ( .A(u0__abc_49347_n4443), .Y(u0__abc_49347_n4443_bF_buf0) );
  BUFX2 BUFX2_672 ( .A(u0__abc_49347_n4444), .Y(u0__abc_49347_n4444_bF_buf3) );
  BUFX2 BUFX2_673 ( .A(u0__abc_49347_n4444), .Y(u0__abc_49347_n4444_bF_buf2) );
  BUFX2 BUFX2_674 ( .A(u0__abc_49347_n4444), .Y(u0__abc_49347_n4444_bF_buf1) );
  BUFX2 BUFX2_675 ( .A(u0__abc_49347_n4444), .Y(u0__abc_49347_n4444_bF_buf0) );
  BUFX2 BUFX2_676 ( .A(u0__abc_49347_n1181), .Y(u0__abc_49347_n1181_bF_buf5) );
  BUFX2 BUFX2_677 ( .A(u0__abc_49347_n1181), .Y(u0__abc_49347_n1181_bF_buf4) );
  BUFX2 BUFX2_678 ( .A(u0__abc_49347_n1181), .Y(u0__abc_49347_n1181_bF_buf3) );
  BUFX2 BUFX2_679 ( .A(u0__abc_49347_n1181), .Y(u0__abc_49347_n1181_bF_buf2) );
  BUFX2 BUFX2_68 ( .A(u3_u0__abc_48231_n708), .Y(u3_u0__abc_48231_n708_bF_buf2) );
  BUFX2 BUFX2_680 ( .A(u0__abc_49347_n1181), .Y(u0__abc_49347_n1181_bF_buf1) );
  BUFX2 BUFX2_681 ( .A(u0__abc_49347_n1181), .Y(u0__abc_49347_n1181_bF_buf0) );
  BUFX2 BUFX2_682 ( .A(u0__abc_49347_n1185), .Y(u0__abc_49347_n1185_bF_buf5) );
  BUFX2 BUFX2_683 ( .A(u0__abc_49347_n1185), .Y(u0__abc_49347_n1185_bF_buf4) );
  BUFX2 BUFX2_684 ( .A(u0__abc_49347_n1185), .Y(u0__abc_49347_n1185_bF_buf3) );
  BUFX2 BUFX2_685 ( .A(u0__abc_49347_n1185), .Y(u0__abc_49347_n1185_bF_buf2) );
  BUFX2 BUFX2_686 ( .A(u0__abc_49347_n1185), .Y(u0__abc_49347_n1185_bF_buf1) );
  BUFX2 BUFX2_687 ( .A(u0__abc_49347_n1185), .Y(u0__abc_49347_n1185_bF_buf0) );
  BUFX2 BUFX2_688 ( .A(u0_u0__abc_43300_n350), .Y(u0_u0__abc_43300_n350_bF_buf4) );
  BUFX2 BUFX2_689 ( .A(u0_u0__abc_43300_n350), .Y(u0_u0__abc_43300_n350_bF_buf3) );
  BUFX2 BUFX2_69 ( .A(u3_u0__abc_48231_n708), .Y(u3_u0__abc_48231_n708_bF_buf1) );
  BUFX2 BUFX2_690 ( .A(u0_u0__abc_43300_n350), .Y(u0_u0__abc_43300_n350_bF_buf2) );
  BUFX2 BUFX2_691 ( .A(u0_u0__abc_43300_n350), .Y(u0_u0__abc_43300_n350_bF_buf1) );
  BUFX2 BUFX2_692 ( .A(u0_u0__abc_43300_n350), .Y(u0_u0__abc_43300_n350_bF_buf0) );
  BUFX2 BUFX2_693 ( .A(u0__abc_49347_n1183_1), .Y(u0__abc_49347_n1183_1_bF_buf5) );
  BUFX2 BUFX2_694 ( .A(u0__abc_49347_n1183_1), .Y(u0__abc_49347_n1183_1_bF_buf4) );
  BUFX2 BUFX2_695 ( .A(u0__abc_49347_n1183_1), .Y(u0__abc_49347_n1183_1_bF_buf3) );
  BUFX2 BUFX2_696 ( .A(u0__abc_49347_n1183_1), .Y(u0__abc_49347_n1183_1_bF_buf2) );
  BUFX2 BUFX2_697 ( .A(u0__abc_49347_n1183_1), .Y(u0__abc_49347_n1183_1_bF_buf1) );
  BUFX2 BUFX2_698 ( .A(u0__abc_49347_n1183_1), .Y(u0__abc_49347_n1183_1_bF_buf0) );
  BUFX2 BUFX2_699 ( .A(u5_cmd_asserted), .Y(u5_cmd_asserted_bF_buf3) );
  BUFX2 BUFX2_7 ( .A(clk_i), .Y(clk_i_hier0_bF_buf4) );
  BUFX2 BUFX2_70 ( .A(u3_u0__abc_48231_n708), .Y(u3_u0__abc_48231_n708_bF_buf0) );
  BUFX2 BUFX2_700 ( .A(u5_cmd_asserted), .Y(u5_cmd_asserted_bF_buf2) );
  BUFX2 BUFX2_701 ( .A(u5_cmd_asserted), .Y(u5_cmd_asserted_bF_buf1) );
  BUFX2 BUFX2_702 ( .A(u5_cmd_asserted), .Y(u5_cmd_asserted_bF_buf0) );
  BUFX2 BUFX2_703 ( .A(u2_u0__abc_47660_n137), .Y(u2_u0__abc_47660_n137_bF_buf4) );
  BUFX2 BUFX2_704 ( .A(u2_u0__abc_47660_n137), .Y(u2_u0__abc_47660_n137_bF_buf3) );
  BUFX2 BUFX2_705 ( .A(u2_u0__abc_47660_n137), .Y(u2_u0__abc_47660_n137_bF_buf2) );
  BUFX2 BUFX2_706 ( .A(u2_u0__abc_47660_n137), .Y(u2_u0__abc_47660_n137_bF_buf1) );
  BUFX2 BUFX2_707 ( .A(u2_u0__abc_47660_n137), .Y(u2_u0__abc_47660_n137_bF_buf0) );
  BUFX2 BUFX2_708 ( .A(u5__abc_54027_n351), .Y(u5__abc_54027_n351_bF_buf3) );
  BUFX2 BUFX2_709 ( .A(u5__abc_54027_n351), .Y(u5__abc_54027_n351_bF_buf2) );
  BUFX2 BUFX2_71 ( .A(u0_u2_init_req_we_FF_INPUT), .Y(u0_u2_init_req_we_FF_INPUT_bF_buf4) );
  BUFX2 BUFX2_710 ( .A(u5__abc_54027_n351), .Y(u5__abc_54027_n351_bF_buf1) );
  BUFX2 BUFX2_711 ( .A(u5__abc_54027_n351), .Y(u5__abc_54027_n351_bF_buf0) );
  BUFX2 BUFX2_712 ( .A(u0_u4_lmr_req_we_FF_INPUT), .Y(u0_u4_lmr_req_we_FF_INPUT_bF_buf7) );
  BUFX2 BUFX2_713 ( .A(u0_u4_lmr_req_we_FF_INPUT), .Y(u0_u4_lmr_req_we_FF_INPUT_bF_buf6) );
  BUFX2 BUFX2_714 ( .A(u0_u4_lmr_req_we_FF_INPUT), .Y(u0_u4_lmr_req_we_FF_INPUT_bF_buf5) );
  BUFX2 BUFX2_715 ( .A(u0_u4_lmr_req_we_FF_INPUT), .Y(u0_u4_lmr_req_we_FF_INPUT_bF_buf4) );
  BUFX2 BUFX2_716 ( .A(u0_u4_lmr_req_we_FF_INPUT), .Y(u0_u4_lmr_req_we_FF_INPUT_bF_buf3) );
  BUFX2 BUFX2_717 ( .A(u0_u4_lmr_req_we_FF_INPUT), .Y(u0_u4_lmr_req_we_FF_INPUT_bF_buf2) );
  BUFX2 BUFX2_718 ( .A(u0_u4_lmr_req_we_FF_INPUT), .Y(u0_u4_lmr_req_we_FF_INPUT_bF_buf1) );
  BUFX2 BUFX2_719 ( .A(u0_u4_lmr_req_we_FF_INPUT), .Y(u0_u4_lmr_req_we_FF_INPUT_bF_buf0) );
  BUFX2 BUFX2_72 ( .A(u0_u2_init_req_we_FF_INPUT), .Y(u0_u2_init_req_we_FF_INPUT_bF_buf3) );
  BUFX2 BUFX2_720 ( .A(u1__abc_45852_n821), .Y(u1__abc_45852_n821_bF_buf3) );
  BUFX2 BUFX2_721 ( .A(u1__abc_45852_n821), .Y(u1__abc_45852_n821_bF_buf2) );
  BUFX2 BUFX2_722 ( .A(u1__abc_45852_n821), .Y(u1__abc_45852_n821_bF_buf1) );
  BUFX2 BUFX2_723 ( .A(u1__abc_45852_n821), .Y(u1__abc_45852_n821_bF_buf0) );
  BUFX2 BUFX2_724 ( .A(u0_u3_lmr_req_we_FF_INPUT), .Y(u0_u3_lmr_req_we_FF_INPUT_bF_buf4) );
  BUFX2 BUFX2_725 ( .A(u0_u3_lmr_req_we_FF_INPUT), .Y(u0_u3_lmr_req_we_FF_INPUT_bF_buf3) );
  BUFX2 BUFX2_726 ( .A(u0_u3_lmr_req_we_FF_INPUT), .Y(u0_u3_lmr_req_we_FF_INPUT_bF_buf2) );
  BUFX2 BUFX2_727 ( .A(u0_u3_lmr_req_we_FF_INPUT), .Y(u0_u3_lmr_req_we_FF_INPUT_bF_buf1) );
  BUFX2 BUFX2_728 ( .A(u0_u3_lmr_req_we_FF_INPUT), .Y(u0_u3_lmr_req_we_FF_INPUT_bF_buf0) );
  BUFX2 BUFX2_729 ( .A(wb_stb_i), .Y(wb_stb_i_bF_buf5) );
  BUFX2 BUFX2_73 ( .A(u0_u2_init_req_we_FF_INPUT), .Y(u0_u2_init_req_we_FF_INPUT_bF_buf2) );
  BUFX2 BUFX2_730 ( .A(wb_stb_i), .Y(wb_stb_i_bF_buf4) );
  BUFX2 BUFX2_731 ( .A(wb_stb_i), .Y(wb_stb_i_bF_buf3) );
  BUFX2 BUFX2_732 ( .A(wb_stb_i), .Y(wb_stb_i_bF_buf2) );
  BUFX2 BUFX2_733 ( .A(wb_stb_i), .Y(wb_stb_i_bF_buf1) );
  BUFX2 BUFX2_734 ( .A(wb_stb_i), .Y(wb_stb_i_bF_buf0) );
  BUFX2 BUFX2_735 ( .A(u0_u2__abc_44109_n340), .Y(u0_u2__abc_44109_n340_bF_buf4) );
  BUFX2 BUFX2_736 ( .A(u0_u2__abc_44109_n340), .Y(u0_u2__abc_44109_n340_bF_buf3) );
  BUFX2 BUFX2_737 ( .A(u0_u2__abc_44109_n340), .Y(u0_u2__abc_44109_n340_bF_buf2) );
  BUFX2 BUFX2_738 ( .A(u0_u2__abc_44109_n340), .Y(u0_u2__abc_44109_n340_bF_buf1) );
  BUFX2 BUFX2_739 ( .A(u0_u2__abc_44109_n340), .Y(u0_u2__abc_44109_n340_bF_buf0) );
  BUFX2 BUFX2_74 ( .A(u0_u2_init_req_we_FF_INPUT), .Y(u0_u2_init_req_we_FF_INPUT_bF_buf1) );
  BUFX2 BUFX2_740 ( .A(row_adr_8_), .Y(row_adr_8_bF_buf6) );
  BUFX2 BUFX2_741 ( .A(row_adr_8_), .Y(row_adr_8_bF_buf5) );
  BUFX2 BUFX2_742 ( .A(row_adr_8_), .Y(row_adr_8_bF_buf4) );
  BUFX2 BUFX2_743 ( .A(row_adr_8_), .Y(row_adr_8_bF_buf3) );
  BUFX2 BUFX2_744 ( .A(row_adr_8_), .Y(row_adr_8_bF_buf2) );
  BUFX2 BUFX2_745 ( .A(row_adr_8_), .Y(row_adr_8_bF_buf1) );
  BUFX2 BUFX2_746 ( .A(row_adr_8_), .Y(row_adr_8_bF_buf0) );
  BUFX2 BUFX2_747 ( .A(u0_u2_lmr_req_we_FF_INPUT), .Y(u0_u2_lmr_req_we_FF_INPUT_bF_buf4) );
  BUFX2 BUFX2_748 ( .A(u0_u2_lmr_req_we_FF_INPUT), .Y(u0_u2_lmr_req_we_FF_INPUT_bF_buf3) );
  BUFX2 BUFX2_749 ( .A(u0_u2_lmr_req_we_FF_INPUT), .Y(u0_u2_lmr_req_we_FF_INPUT_bF_buf2) );
  BUFX2 BUFX2_75 ( .A(u0_u2_init_req_we_FF_INPUT), .Y(u0_u2_init_req_we_FF_INPUT_bF_buf0) );
  BUFX2 BUFX2_750 ( .A(u0_u2_lmr_req_we_FF_INPUT), .Y(u0_u2_lmr_req_we_FF_INPUT_bF_buf1) );
  BUFX2 BUFX2_751 ( .A(u0_u2_lmr_req_we_FF_INPUT), .Y(u0_u2_lmr_req_we_FF_INPUT_bF_buf0) );
  BUFX2 BUFX2_752 ( .A(row_adr_5_), .Y(row_adr_5_bF_buf6) );
  BUFX2 BUFX2_753 ( .A(row_adr_5_), .Y(row_adr_5_bF_buf5) );
  BUFX2 BUFX2_754 ( .A(row_adr_5_), .Y(row_adr_5_bF_buf4) );
  BUFX2 BUFX2_755 ( .A(row_adr_5_), .Y(row_adr_5_bF_buf3) );
  BUFX2 BUFX2_756 ( .A(row_adr_5_), .Y(row_adr_5_bF_buf2) );
  BUFX2 BUFX2_757 ( .A(row_adr_5_), .Y(row_adr_5_bF_buf1) );
  BUFX2 BUFX2_758 ( .A(row_adr_5_), .Y(row_adr_5_bF_buf0) );
  BUFX2 BUFX2_759 ( .A(u6__abc_56056_n154), .Y(u6__abc_56056_n154_bF_buf4) );
  BUFX2 BUFX2_76 ( .A(row_adr_4_), .Y(row_adr_4_bF_buf6) );
  BUFX2 BUFX2_760 ( .A(u6__abc_56056_n154), .Y(u6__abc_56056_n154_bF_buf3) );
  BUFX2 BUFX2_761 ( .A(u6__abc_56056_n154), .Y(u6__abc_56056_n154_bF_buf2) );
  BUFX2 BUFX2_762 ( .A(u6__abc_56056_n154), .Y(u6__abc_56056_n154_bF_buf1) );
  BUFX2 BUFX2_763 ( .A(u6__abc_56056_n154), .Y(u6__abc_56056_n154_bF_buf0) );
  BUFX2 BUFX2_764 ( .A(u1__abc_45852_n554_1), .Y(u1__abc_45852_n554_1_bF_buf4) );
  BUFX2 BUFX2_765 ( .A(u1__abc_45852_n554_1), .Y(u1__abc_45852_n554_1_bF_buf3) );
  BUFX2 BUFX2_766 ( .A(u1__abc_45852_n554_1), .Y(u1__abc_45852_n554_1_bF_buf2) );
  BUFX2 BUFX2_767 ( .A(u1__abc_45852_n554_1), .Y(u1__abc_45852_n554_1_bF_buf1) );
  BUFX2 BUFX2_768 ( .A(u1__abc_45852_n554_1), .Y(u1__abc_45852_n554_1_bF_buf0) );
  BUFX2 BUFX2_769 ( .A(u3__abc_46775_n448), .Y(u3__abc_46775_n448_bF_buf3) );
  BUFX2 BUFX2_77 ( .A(row_adr_4_), .Y(row_adr_4_bF_buf5) );
  BUFX2 BUFX2_770 ( .A(u3__abc_46775_n448), .Y(u3__abc_46775_n448_bF_buf2) );
  BUFX2 BUFX2_771 ( .A(u3__abc_46775_n448), .Y(u3__abc_46775_n448_bF_buf1) );
  BUFX2 BUFX2_772 ( .A(u3__abc_46775_n448), .Y(u3__abc_46775_n448_bF_buf0) );
  BUFX2 BUFX2_773 ( .A(row_adr_2_), .Y(row_adr_2_bF_buf6) );
  BUFX2 BUFX2_774 ( .A(row_adr_2_), .Y(row_adr_2_bF_buf5) );
  BUFX2 BUFX2_775 ( .A(row_adr_2_), .Y(row_adr_2_bF_buf4) );
  BUFX2 BUFX2_776 ( .A(row_adr_2_), .Y(row_adr_2_bF_buf3) );
  BUFX2 BUFX2_777 ( .A(row_adr_2_), .Y(row_adr_2_bF_buf2) );
  BUFX2 BUFX2_778 ( .A(row_adr_2_), .Y(row_adr_2_bF_buf1) );
  BUFX2 BUFX2_779 ( .A(row_adr_2_), .Y(row_adr_2_bF_buf0) );
  BUFX2 BUFX2_78 ( .A(row_adr_4_), .Y(row_adr_4_bF_buf4) );
  BUFX2 BUFX2_780 ( .A(u0_u3__abc_44466_n364), .Y(u0_u3__abc_44466_n364_bF_buf4) );
  BUFX2 BUFX2_781 ( .A(u0_u3__abc_44466_n364), .Y(u0_u3__abc_44466_n364_bF_buf3) );
  BUFX2 BUFX2_782 ( .A(u0_u3__abc_44466_n364), .Y(u0_u3__abc_44466_n364_bF_buf2) );
  BUFX2 BUFX2_783 ( .A(u0_u3__abc_44466_n364), .Y(u0_u3__abc_44466_n364_bF_buf1) );
  BUFX2 BUFX2_784 ( .A(u0_u3__abc_44466_n364), .Y(u0_u3__abc_44466_n364_bF_buf0) );
  BUFX2 BUFX2_785 ( .A(u0__abc_49347_n2730), .Y(u0__abc_49347_n2730_bF_buf5) );
  BUFX2 BUFX2_786 ( .A(u0__abc_49347_n2730), .Y(u0__abc_49347_n2730_bF_buf4) );
  BUFX2 BUFX2_787 ( .A(u0__abc_49347_n2730), .Y(u0__abc_49347_n2730_bF_buf3) );
  BUFX2 BUFX2_788 ( .A(u0__abc_49347_n2730), .Y(u0__abc_49347_n2730_bF_buf2) );
  BUFX2 BUFX2_789 ( .A(u0__abc_49347_n2730), .Y(u0__abc_49347_n2730_bF_buf1) );
  BUFX2 BUFX2_79 ( .A(row_adr_4_), .Y(row_adr_4_bF_buf3) );
  BUFX2 BUFX2_790 ( .A(u0__abc_49347_n2730), .Y(u0__abc_49347_n2730_bF_buf0) );
  BUFX2 BUFX2_791 ( .A(u0_u3__abc_44466_n205_1), .Y(u0_u3__abc_44466_n205_1_bF_buf4) );
  BUFX2 BUFX2_792 ( .A(u0_u3__abc_44466_n205_1), .Y(u0_u3__abc_44466_n205_1_bF_buf3) );
  BUFX2 BUFX2_793 ( .A(u0_u3__abc_44466_n205_1), .Y(u0_u3__abc_44466_n205_1_bF_buf2) );
  BUFX2 BUFX2_794 ( .A(u0_u3__abc_44466_n205_1), .Y(u0_u3__abc_44466_n205_1_bF_buf1) );
  BUFX2 BUFX2_795 ( .A(u0_u3__abc_44466_n205_1), .Y(u0_u3__abc_44466_n205_1_bF_buf0) );
  BUFX2 BUFX2_796 ( .A(\wb_addr_i[25] ), .Y(wb_addr_i_25_bF_buf3) );
  BUFX2 BUFX2_797 ( .A(\wb_addr_i[25] ), .Y(wb_addr_i_25_bF_buf2) );
  BUFX2 BUFX2_798 ( .A(\wb_addr_i[25] ), .Y(wb_addr_i_25_bF_buf1) );
  BUFX2 BUFX2_799 ( .A(\wb_addr_i[25] ), .Y(wb_addr_i_25_bF_buf0) );
  BUFX2 BUFX2_8 ( .A(clk_i), .Y(clk_i_hier0_bF_buf3) );
  BUFX2 BUFX2_80 ( .A(row_adr_4_), .Y(row_adr_4_bF_buf2) );
  BUFX2 BUFX2_800 ( .A(u3__abc_46775_n277_1), .Y(u3__abc_46775_n277_1_bF_buf5) );
  BUFX2 BUFX2_801 ( .A(u3__abc_46775_n277_1), .Y(u3__abc_46775_n277_1_bF_buf4) );
  BUFX2 BUFX2_802 ( .A(u3__abc_46775_n277_1), .Y(u3__abc_46775_n277_1_bF_buf3) );
  BUFX2 BUFX2_803 ( .A(u3__abc_46775_n277_1), .Y(u3__abc_46775_n277_1_bF_buf2) );
  BUFX2 BUFX2_804 ( .A(u3__abc_46775_n277_1), .Y(u3__abc_46775_n277_1_bF_buf1) );
  BUFX2 BUFX2_805 ( .A(u3__abc_46775_n277_1), .Y(u3__abc_46775_n277_1_bF_buf0) );
  BUFX2 BUFX2_806 ( .A(u0_u5_init_req_we_FF_INPUT), .Y(u0_u5_init_req_we_FF_INPUT_bF_buf7) );
  BUFX2 BUFX2_807 ( .A(u0_u5_init_req_we_FF_INPUT), .Y(u0_u5_init_req_we_FF_INPUT_bF_buf6) );
  BUFX2 BUFX2_808 ( .A(u0_u5_init_req_we_FF_INPUT), .Y(u0_u5_init_req_we_FF_INPUT_bF_buf5) );
  BUFX2 BUFX2_809 ( .A(u0_u5_init_req_we_FF_INPUT), .Y(u0_u5_init_req_we_FF_INPUT_bF_buf4) );
  BUFX2 BUFX2_81 ( .A(row_adr_4_), .Y(row_adr_4_bF_buf1) );
  BUFX2 BUFX2_810 ( .A(u0_u5_init_req_we_FF_INPUT), .Y(u0_u5_init_req_we_FF_INPUT_bF_buf3) );
  BUFX2 BUFX2_811 ( .A(u0_u5_init_req_we_FF_INPUT), .Y(u0_u5_init_req_we_FF_INPUT_bF_buf2) );
  BUFX2 BUFX2_812 ( .A(u0_u5_init_req_we_FF_INPUT), .Y(u0_u5_init_req_we_FF_INPUT_bF_buf1) );
  BUFX2 BUFX2_813 ( .A(u0_u5_init_req_we_FF_INPUT), .Y(u0_u5_init_req_we_FF_INPUT_bF_buf0) );
  BUFX2 BUFX2_814 ( .A(u0__abc_49347_n4582), .Y(u0__abc_49347_n4582_bF_buf4) );
  BUFX2 BUFX2_815 ( .A(u0__abc_49347_n4582), .Y(u0__abc_49347_n4582_bF_buf3) );
  BUFX2 BUFX2_816 ( .A(u0__abc_49347_n4582), .Y(u0__abc_49347_n4582_bF_buf2) );
  BUFX2 BUFX2_817 ( .A(u0__abc_49347_n4582), .Y(u0__abc_49347_n4582_bF_buf1) );
  BUFX2 BUFX2_818 ( .A(u0__abc_49347_n4582), .Y(u0__abc_49347_n4582_bF_buf0) );
  BUFX2 BUFX2_819 ( .A(u0__abc_49347_n4584), .Y(u0__abc_49347_n4584_bF_buf4) );
  BUFX2 BUFX2_82 ( .A(row_adr_4_), .Y(row_adr_4_bF_buf0) );
  BUFX2 BUFX2_820 ( .A(u0__abc_49347_n4584), .Y(u0__abc_49347_n4584_bF_buf3) );
  BUFX2 BUFX2_821 ( .A(u0__abc_49347_n4584), .Y(u0__abc_49347_n4584_bF_buf2) );
  BUFX2 BUFX2_822 ( .A(u0__abc_49347_n4584), .Y(u0__abc_49347_n4584_bF_buf1) );
  BUFX2 BUFX2_823 ( .A(u0__abc_49347_n4584), .Y(u0__abc_49347_n4584_bF_buf0) );
  BUFX2 BUFX2_824 ( .A(u0__abc_49347_n4586), .Y(u0__abc_49347_n4586_bF_buf4) );
  BUFX2 BUFX2_825 ( .A(u0__abc_49347_n4586), .Y(u0__abc_49347_n4586_bF_buf3) );
  BUFX2 BUFX2_826 ( .A(u0__abc_49347_n4586), .Y(u0__abc_49347_n4586_bF_buf2) );
  BUFX2 BUFX2_827 ( .A(u0__abc_49347_n4586), .Y(u0__abc_49347_n4586_bF_buf1) );
  BUFX2 BUFX2_828 ( .A(u0__abc_49347_n4586), .Y(u0__abc_49347_n4586_bF_buf0) );
  BUFX2 BUFX2_829 ( .A(u0__abc_49347_n4589), .Y(u0__abc_49347_n4589_bF_buf4) );
  BUFX2 BUFX2_83 ( .A(u6__abc_56056_n144), .Y(u6__abc_56056_n144_bF_buf5) );
  BUFX2 BUFX2_830 ( .A(u0__abc_49347_n4589), .Y(u0__abc_49347_n4589_bF_buf3) );
  BUFX2 BUFX2_831 ( .A(u0__abc_49347_n4589), .Y(u0__abc_49347_n4589_bF_buf2) );
  BUFX2 BUFX2_832 ( .A(u0__abc_49347_n4589), .Y(u0__abc_49347_n4589_bF_buf1) );
  BUFX2 BUFX2_833 ( .A(u0__abc_49347_n4589), .Y(u0__abc_49347_n4589_bF_buf0) );
  BUFX2 BUFX2_834 ( .A(u1__abc_45852_n261), .Y(u1__abc_45852_n261_bF_buf4) );
  BUFX2 BUFX2_835 ( .A(u1__abc_45852_n261), .Y(u1__abc_45852_n261_bF_buf3) );
  BUFX2 BUFX2_836 ( .A(u1__abc_45852_n261), .Y(u1__abc_45852_n261_bF_buf2) );
  BUFX2 BUFX2_837 ( .A(u1__abc_45852_n261), .Y(u1__abc_45852_n261_bF_buf1) );
  BUFX2 BUFX2_838 ( .A(u1__abc_45852_n261), .Y(u1__abc_45852_n261_bF_buf0) );
  BUFX2 BUFX2_839 ( .A(u0_u1_init_req_we_FF_INPUT), .Y(u0_u1_init_req_we_FF_INPUT_bF_buf7) );
  BUFX2 BUFX2_84 ( .A(u6__abc_56056_n144), .Y(u6__abc_56056_n144_bF_buf4) );
  BUFX2 BUFX2_840 ( .A(u0_u1_init_req_we_FF_INPUT), .Y(u0_u1_init_req_we_FF_INPUT_bF_buf6) );
  BUFX2 BUFX2_841 ( .A(u0_u1_init_req_we_FF_INPUT), .Y(u0_u1_init_req_we_FF_INPUT_bF_buf5) );
  BUFX2 BUFX2_842 ( .A(u0_u1_init_req_we_FF_INPUT), .Y(u0_u1_init_req_we_FF_INPUT_bF_buf4) );
  BUFX2 BUFX2_843 ( .A(u0_u1_init_req_we_FF_INPUT), .Y(u0_u1_init_req_we_FF_INPUT_bF_buf3) );
  BUFX2 BUFX2_844 ( .A(u0_u1_init_req_we_FF_INPUT), .Y(u0_u1_init_req_we_FF_INPUT_bF_buf2) );
  BUFX2 BUFX2_845 ( .A(u0_u1_init_req_we_FF_INPUT), .Y(u0_u1_init_req_we_FF_INPUT_bF_buf1) );
  BUFX2 BUFX2_846 ( .A(u0_u1_init_req_we_FF_INPUT), .Y(u0_u1_init_req_we_FF_INPUT_bF_buf0) );
  BUFX2 BUFX2_847 ( .A(u3_u0__abc_48231_n563), .Y(u3_u0__abc_48231_n563_bF_buf7) );
  BUFX2 BUFX2_848 ( .A(u3_u0__abc_48231_n563), .Y(u3_u0__abc_48231_n563_bF_buf6) );
  BUFX2 BUFX2_849 ( .A(u3_u0__abc_48231_n563), .Y(u3_u0__abc_48231_n563_bF_buf5) );
  BUFX2 BUFX2_85 ( .A(u6__abc_56056_n144), .Y(u6__abc_56056_n144_bF_buf3) );
  BUFX2 BUFX2_850 ( .A(u3_u0__abc_48231_n563), .Y(u3_u0__abc_48231_n563_bF_buf4) );
  BUFX2 BUFX2_851 ( .A(u3_u0__abc_48231_n563), .Y(u3_u0__abc_48231_n563_bF_buf3) );
  BUFX2 BUFX2_852 ( .A(u3_u0__abc_48231_n563), .Y(u3_u0__abc_48231_n563_bF_buf2) );
  BUFX2 BUFX2_853 ( .A(u3_u0__abc_48231_n563), .Y(u3_u0__abc_48231_n563_bF_buf1) );
  BUFX2 BUFX2_854 ( .A(u3_u0__abc_48231_n563), .Y(u3_u0__abc_48231_n563_bF_buf0) );
  BUFX2 BUFX2_855 ( .A(_abc_55805_n240), .Y(_abc_55805_n240_bF_buf5) );
  BUFX2 BUFX2_856 ( .A(_abc_55805_n240), .Y(_abc_55805_n240_bF_buf4) );
  BUFX2 BUFX2_857 ( .A(_abc_55805_n240), .Y(_abc_55805_n240_bF_buf3) );
  BUFX2 BUFX2_858 ( .A(_abc_55805_n240), .Y(_abc_55805_n240_bF_buf2) );
  BUFX2 BUFX2_859 ( .A(_abc_55805_n240), .Y(_abc_55805_n240_bF_buf1) );
  BUFX2 BUFX2_86 ( .A(u6__abc_56056_n144), .Y(u6__abc_56056_n144_bF_buf2) );
  BUFX2 BUFX2_860 ( .A(_abc_55805_n240), .Y(_abc_55805_n240_bF_buf0) );
  BUFX2 BUFX2_861 ( .A(u3_u0__abc_48231_n1042), .Y(u3_u0__abc_48231_n1042_bF_buf5) );
  BUFX2 BUFX2_862 ( .A(u3_u0__abc_48231_n1042), .Y(u3_u0__abc_48231_n1042_bF_buf4) );
  BUFX2 BUFX2_863 ( .A(u3_u0__abc_48231_n1042), .Y(u3_u0__abc_48231_n1042_bF_buf3) );
  BUFX2 BUFX2_864 ( .A(u3_u0__abc_48231_n1042), .Y(u3_u0__abc_48231_n1042_bF_buf2) );
  BUFX2 BUFX2_865 ( .A(u3_u0__abc_48231_n1042), .Y(u3_u0__abc_48231_n1042_bF_buf1) );
  BUFX2 BUFX2_866 ( .A(u3_u0__abc_48231_n1042), .Y(u3_u0__abc_48231_n1042_bF_buf0) );
  BUFX2 BUFX2_867 ( .A(u0_rst_r3), .Y(u0_rst_r3_bF_buf4) );
  BUFX2 BUFX2_868 ( .A(u0_rst_r3), .Y(u0_rst_r3_bF_buf3) );
  BUFX2 BUFX2_869 ( .A(u0_rst_r3), .Y(u0_rst_r3_bF_buf2) );
  BUFX2 BUFX2_87 ( .A(u6__abc_56056_n144), .Y(u6__abc_56056_n144_bF_buf1) );
  BUFX2 BUFX2_870 ( .A(u0_rst_r3), .Y(u0_rst_r3_bF_buf1) );
  BUFX2 BUFX2_871 ( .A(u0_rst_r3), .Y(u0_rst_r3_bF_buf0) );
  BUFX2 BUFX2_872 ( .A(u3_u0__abc_48231_n1047), .Y(u3_u0__abc_48231_n1047_bF_buf5) );
  BUFX2 BUFX2_873 ( .A(u3_u0__abc_48231_n1047), .Y(u3_u0__abc_48231_n1047_bF_buf4) );
  BUFX2 BUFX2_874 ( .A(u3_u0__abc_48231_n1047), .Y(u3_u0__abc_48231_n1047_bF_buf3) );
  BUFX2 BUFX2_875 ( .A(u3_u0__abc_48231_n1047), .Y(u3_u0__abc_48231_n1047_bF_buf2) );
  BUFX2 BUFX2_876 ( .A(u3_u0__abc_48231_n1047), .Y(u3_u0__abc_48231_n1047_bF_buf1) );
  BUFX2 BUFX2_877 ( .A(u3_u0__abc_48231_n1047), .Y(u3_u0__abc_48231_n1047_bF_buf0) );
  BUFX2 BUFX2_878 ( .A(spec_req_cs_6_), .Y(spec_req_cs_6_bF_buf5) );
  BUFX2 BUFX2_879 ( .A(spec_req_cs_6_), .Y(spec_req_cs_6_bF_buf4) );
  BUFX2 BUFX2_88 ( .A(u6__abc_56056_n144), .Y(u6__abc_56056_n144_bF_buf0) );
  BUFX2 BUFX2_880 ( .A(spec_req_cs_6_), .Y(spec_req_cs_6_bF_buf3) );
  BUFX2 BUFX2_881 ( .A(spec_req_cs_6_), .Y(spec_req_cs_6_bF_buf2) );
  BUFX2 BUFX2_882 ( .A(spec_req_cs_6_), .Y(spec_req_cs_6_bF_buf1) );
  BUFX2 BUFX2_883 ( .A(spec_req_cs_6_), .Y(spec_req_cs_6_bF_buf0) );
  BUFX2 BUFX2_884 ( .A(row_adr_11_), .Y(row_adr_11_bF_buf6) );
  BUFX2 BUFX2_885 ( .A(row_adr_11_), .Y(row_adr_11_bF_buf5) );
  BUFX2 BUFX2_886 ( .A(row_adr_11_), .Y(row_adr_11_bF_buf4) );
  BUFX2 BUFX2_887 ( .A(row_adr_11_), .Y(row_adr_11_bF_buf3) );
  BUFX2 BUFX2_888 ( .A(row_adr_11_), .Y(row_adr_11_bF_buf2) );
  BUFX2 BUFX2_889 ( .A(row_adr_11_), .Y(row_adr_11_bF_buf1) );
  BUFX2 BUFX2_89 ( .A(row_adr_1_), .Y(row_adr_1_bF_buf6) );
  BUFX2 BUFX2_890 ( .A(row_adr_11_), .Y(row_adr_11_bF_buf0) );
  BUFX2 BUFX2_891 ( .A(u0__abc_49347_n4526), .Y(u0__abc_49347_n4526_bF_buf4) );
  BUFX2 BUFX2_892 ( .A(u0__abc_49347_n4526), .Y(u0__abc_49347_n4526_bF_buf3) );
  BUFX2 BUFX2_893 ( .A(u0__abc_49347_n4526), .Y(u0__abc_49347_n4526_bF_buf2) );
  BUFX2 BUFX2_894 ( .A(u0__abc_49347_n4526), .Y(u0__abc_49347_n4526_bF_buf1) );
  BUFX2 BUFX2_895 ( .A(u0__abc_49347_n4526), .Y(u0__abc_49347_n4526_bF_buf0) );
  BUFX2 BUFX2_896 ( .A(u0__abc_49347_n4528), .Y(u0__abc_49347_n4528_bF_buf4) );
  BUFX2 BUFX2_897 ( .A(u0__abc_49347_n4528), .Y(u0__abc_49347_n4528_bF_buf3) );
  BUFX2 BUFX2_898 ( .A(u0__abc_49347_n4528), .Y(u0__abc_49347_n4528_bF_buf2) );
  BUFX2 BUFX2_899 ( .A(u0__abc_49347_n4528), .Y(u0__abc_49347_n4528_bF_buf1) );
  BUFX2 BUFX2_9 ( .A(clk_i), .Y(clk_i_hier0_bF_buf2) );
  BUFX2 BUFX2_90 ( .A(row_adr_1_), .Y(row_adr_1_bF_buf5) );
  BUFX2 BUFX2_900 ( .A(u0__abc_49347_n4528), .Y(u0__abc_49347_n4528_bF_buf0) );
  BUFX2 BUFX2_901 ( .A(u0__abc_49347_n1180_1), .Y(u0__abc_49347_n1180_1_bF_buf5) );
  BUFX2 BUFX2_902 ( .A(u0__abc_49347_n1180_1), .Y(u0__abc_49347_n1180_1_bF_buf4) );
  BUFX2 BUFX2_903 ( .A(u0__abc_49347_n1180_1), .Y(u0__abc_49347_n1180_1_bF_buf3) );
  BUFX2 BUFX2_904 ( .A(u0__abc_49347_n1180_1), .Y(u0__abc_49347_n1180_1_bF_buf2) );
  BUFX2 BUFX2_905 ( .A(u0__abc_49347_n1180_1), .Y(u0__abc_49347_n1180_1_bF_buf1) );
  BUFX2 BUFX2_906 ( .A(u0__abc_49347_n1180_1), .Y(u0__abc_49347_n1180_1_bF_buf0) );
  BUFX2 BUFX2_907 ( .A(spec_req_cs_3_), .Y(spec_req_cs_3_bF_buf5) );
  BUFX2 BUFX2_908 ( .A(spec_req_cs_3_), .Y(spec_req_cs_3_bF_buf4) );
  BUFX2 BUFX2_909 ( .A(spec_req_cs_3_), .Y(spec_req_cs_3_bF_buf3) );
  BUFX2 BUFX2_91 ( .A(row_adr_1_), .Y(row_adr_1_bF_buf4) );
  BUFX2 BUFX2_910 ( .A(spec_req_cs_3_), .Y(spec_req_cs_3_bF_buf2) );
  BUFX2 BUFX2_911 ( .A(spec_req_cs_3_), .Y(spec_req_cs_3_bF_buf1) );
  BUFX2 BUFX2_912 ( .A(spec_req_cs_3_), .Y(spec_req_cs_3_bF_buf0) );
  BUFX2 BUFX2_913 ( .A(u1__abc_45852_n556), .Y(u1__abc_45852_n556_bF_buf3) );
  BUFX2 BUFX2_914 ( .A(u1__abc_45852_n556), .Y(u1__abc_45852_n556_bF_buf2) );
  BUFX2 BUFX2_915 ( .A(u1__abc_45852_n556), .Y(u1__abc_45852_n556_bF_buf1) );
  BUFX2 BUFX2_916 ( .A(u1__abc_45852_n556), .Y(u1__abc_45852_n556_bF_buf0) );
  BUFX2 BUFX2_917 ( .A(u3_u0__abc_48231_n853), .Y(u3_u0__abc_48231_n853_bF_buf7) );
  BUFX2 BUFX2_918 ( .A(u3_u0__abc_48231_n853), .Y(u3_u0__abc_48231_n853_bF_buf6) );
  BUFX2 BUFX2_919 ( .A(u3_u0__abc_48231_n853), .Y(u3_u0__abc_48231_n853_bF_buf5) );
  BUFX2 BUFX2_92 ( .A(row_adr_1_), .Y(row_adr_1_bF_buf3) );
  BUFX2 BUFX2_920 ( .A(u3_u0__abc_48231_n853), .Y(u3_u0__abc_48231_n853_bF_buf4) );
  BUFX2 BUFX2_921 ( .A(u3_u0__abc_48231_n853), .Y(u3_u0__abc_48231_n853_bF_buf3) );
  BUFX2 BUFX2_922 ( .A(u3_u0__abc_48231_n853), .Y(u3_u0__abc_48231_n853_bF_buf2) );
  BUFX2 BUFX2_923 ( .A(u3_u0__abc_48231_n853), .Y(u3_u0__abc_48231_n853_bF_buf1) );
  BUFX2 BUFX2_924 ( .A(u3_u0__abc_48231_n853), .Y(u3_u0__abc_48231_n853_bF_buf0) );
  BUFX2 BUFX2_925 ( .A(spec_req_cs_0_), .Y(spec_req_cs_0_bF_buf5) );
  BUFX2 BUFX2_926 ( .A(spec_req_cs_0_), .Y(spec_req_cs_0_bF_buf4) );
  BUFX2 BUFX2_927 ( .A(spec_req_cs_0_), .Y(spec_req_cs_0_bF_buf3) );
  BUFX2 BUFX2_928 ( .A(spec_req_cs_0_), .Y(spec_req_cs_0_bF_buf2) );
  BUFX2 BUFX2_929 ( .A(spec_req_cs_0_), .Y(spec_req_cs_0_bF_buf1) );
  BUFX2 BUFX2_93 ( .A(row_adr_1_), .Y(row_adr_1_bF_buf2) );
  BUFX2 BUFX2_930 ( .A(spec_req_cs_0_), .Y(spec_req_cs_0_bF_buf0) );
  BUFX2 BUFX2_931 ( .A(u1__abc_45852_n901), .Y(u1__abc_45852_n901_bF_buf4) );
  BUFX2 BUFX2_932 ( .A(u1__abc_45852_n901), .Y(u1__abc_45852_n901_bF_buf3) );
  BUFX2 BUFX2_933 ( .A(u1__abc_45852_n901), .Y(u1__abc_45852_n901_bF_buf2) );
  BUFX2 BUFX2_934 ( .A(u1__abc_45852_n901), .Y(u1__abc_45852_n901_bF_buf1) );
  BUFX2 BUFX2_935 ( .A(u1__abc_45852_n901), .Y(u1__abc_45852_n901_bF_buf0) );
  BUFX2 BUFX2_936 ( .A(u1__abc_45852_n903), .Y(u1__abc_45852_n903_bF_buf3) );
  BUFX2 BUFX2_937 ( .A(u1__abc_45852_n903), .Y(u1__abc_45852_n903_bF_buf2) );
  BUFX2 BUFX2_938 ( .A(u1__abc_45852_n903), .Y(u1__abc_45852_n903_bF_buf1) );
  BUFX2 BUFX2_939 ( .A(u1__abc_45852_n903), .Y(u1__abc_45852_n903_bF_buf0) );
  BUFX2 BUFX2_94 ( .A(row_adr_1_), .Y(row_adr_1_bF_buf1) );
  BUFX2 BUFX2_940 ( .A(u0__abc_49347_n1203), .Y(u0__abc_49347_n1203_bF_buf5) );
  BUFX2 BUFX2_941 ( .A(u0__abc_49347_n1203), .Y(u0__abc_49347_n1203_bF_buf4) );
  BUFX2 BUFX2_942 ( .A(u0__abc_49347_n1203), .Y(u0__abc_49347_n1203_bF_buf3) );
  BUFX2 BUFX2_943 ( .A(u0__abc_49347_n1203), .Y(u0__abc_49347_n1203_bF_buf2) );
  BUFX2 BUFX2_944 ( .A(u0__abc_49347_n1203), .Y(u0__abc_49347_n1203_bF_buf1) );
  BUFX2 BUFX2_945 ( .A(u0__abc_49347_n1203), .Y(u0__abc_49347_n1203_bF_buf0) );
  BUFX2 BUFX2_946 ( .A(mc_clk_i), .Y(mc_clk_i_bF_buf10) );
  BUFX2 BUFX2_947 ( .A(mc_clk_i), .Y(mc_clk_i_bF_buf9) );
  BUFX2 BUFX2_948 ( .A(mc_clk_i), .Y(mc_clk_i_bF_buf8) );
  BUFX2 BUFX2_949 ( .A(mc_clk_i), .Y(mc_clk_i_bF_buf7) );
  BUFX2 BUFX2_95 ( .A(row_adr_1_), .Y(row_adr_1_bF_buf0) );
  BUFX2 BUFX2_950 ( .A(mc_clk_i), .Y(mc_clk_i_bF_buf6) );
  BUFX2 BUFX2_951 ( .A(mc_clk_i), .Y(mc_clk_i_bF_buf5) );
  BUFX2 BUFX2_952 ( .A(mc_clk_i), .Y(mc_clk_i_bF_buf4) );
  BUFX2 BUFX2_953 ( .A(mc_clk_i), .Y(mc_clk_i_bF_buf3) );
  BUFX2 BUFX2_954 ( .A(mc_clk_i), .Y(mc_clk_i_bF_buf2) );
  BUFX2 BUFX2_955 ( .A(mc_clk_i), .Y(mc_clk_i_bF_buf1) );
  BUFX2 BUFX2_956 ( .A(mc_clk_i), .Y(mc_clk_i_bF_buf0) );
  BUFX2 BUFX2_957 ( .A(u0__abc_49347_n1175), .Y(u0__abc_49347_n1175_bF_buf6) );
  BUFX2 BUFX2_958 ( .A(u0__abc_49347_n1175), .Y(u0__abc_49347_n1175_bF_buf5) );
  BUFX2 BUFX2_959 ( .A(u0__abc_49347_n1175), .Y(u0__abc_49347_n1175_bF_buf4) );
  BUFX2 BUFX2_96 ( .A(u2_u5__abc_47660_n137), .Y(u2_u5__abc_47660_n137_bF_buf4) );
  BUFX2 BUFX2_960 ( .A(u0__abc_49347_n1175), .Y(u0__abc_49347_n1175_bF_buf3) );
  BUFX2 BUFX2_961 ( .A(u0__abc_49347_n1175), .Y(u0__abc_49347_n1175_bF_buf2) );
  BUFX2 BUFX2_962 ( .A(u0__abc_49347_n1175), .Y(u0__abc_49347_n1175_bF_buf1) );
  BUFX2 BUFX2_963 ( .A(u0__abc_49347_n1175), .Y(u0__abc_49347_n1175_bF_buf0) );
  BUFX2 BUFX2_964 ( .A(u0__abc_49347_n1179), .Y(u0__abc_49347_n1179_bF_buf5) );
  BUFX2 BUFX2_965 ( .A(u0__abc_49347_n1179), .Y(u0__abc_49347_n1179_bF_buf4) );
  BUFX2 BUFX2_966 ( .A(u0__abc_49347_n1179), .Y(u0__abc_49347_n1179_bF_buf3) );
  BUFX2 BUFX2_967 ( .A(u0__abc_49347_n1179), .Y(u0__abc_49347_n1179_bF_buf2) );
  BUFX2 BUFX2_968 ( .A(u0__abc_49347_n1179), .Y(u0__abc_49347_n1179_bF_buf1) );
  BUFX2 BUFX2_969 ( .A(u0__abc_49347_n1179), .Y(u0__abc_49347_n1179_bF_buf0) );
  BUFX2 BUFX2_97 ( .A(u2_u5__abc_47660_n137), .Y(u2_u5__abc_47660_n137_bF_buf3) );
  BUFX2 BUFX2_970 ( .A(_auto_iopadmap_cc_313_execute_56218_0_), .Y(\mc_addr_pad_o[0] ) );
  BUFX2 BUFX2_971 ( .A(_auto_iopadmap_cc_313_execute_56218_1_), .Y(\mc_addr_pad_o[1] ) );
  BUFX2 BUFX2_972 ( .A(_auto_iopadmap_cc_313_execute_56218_2_), .Y(\mc_addr_pad_o[2] ) );
  BUFX2 BUFX2_973 ( .A(_auto_iopadmap_cc_313_execute_56218_3_), .Y(\mc_addr_pad_o[3] ) );
  BUFX2 BUFX2_974 ( .A(_auto_iopadmap_cc_313_execute_56218_4_), .Y(\mc_addr_pad_o[4] ) );
  BUFX2 BUFX2_975 ( .A(_auto_iopadmap_cc_313_execute_56218_5_), .Y(\mc_addr_pad_o[5] ) );
  BUFX2 BUFX2_976 ( .A(_auto_iopadmap_cc_313_execute_56218_6_), .Y(\mc_addr_pad_o[6] ) );
  BUFX2 BUFX2_977 ( .A(_auto_iopadmap_cc_313_execute_56218_7_), .Y(\mc_addr_pad_o[7] ) );
  BUFX2 BUFX2_978 ( .A(_auto_iopadmap_cc_313_execute_56218_8_), .Y(\mc_addr_pad_o[8] ) );
  BUFX2 BUFX2_979 ( .A(_auto_iopadmap_cc_313_execute_56218_9_), .Y(\mc_addr_pad_o[9] ) );
  BUFX2 BUFX2_98 ( .A(u2_u5__abc_47660_n137), .Y(u2_u5__abc_47660_n137_bF_buf2) );
  BUFX2 BUFX2_980 ( .A(_auto_iopadmap_cc_313_execute_56218_10_), .Y(\mc_addr_pad_o[10] ) );
  BUFX2 BUFX2_981 ( .A(_auto_iopadmap_cc_313_execute_56218_11_), .Y(\mc_addr_pad_o[11] ) );
  BUFX2 BUFX2_982 ( .A(_auto_iopadmap_cc_313_execute_56218_12_), .Y(\mc_addr_pad_o[12] ) );
  BUFX2 BUFX2_983 ( .A(_auto_iopadmap_cc_313_execute_56218_13_), .Y(\mc_addr_pad_o[13] ) );
  BUFX2 BUFX2_984 ( .A(_auto_iopadmap_cc_313_execute_56218_14_), .Y(\mc_addr_pad_o[14] ) );
  BUFX2 BUFX2_985 ( .A(_auto_iopadmap_cc_313_execute_56218_15_), .Y(\mc_addr_pad_o[15] ) );
  BUFX2 BUFX2_986 ( .A(_auto_iopadmap_cc_313_execute_56218_16_), .Y(\mc_addr_pad_o[16] ) );
  BUFX2 BUFX2_987 ( .A(_auto_iopadmap_cc_313_execute_56218_17_), .Y(\mc_addr_pad_o[17] ) );
  BUFX2 BUFX2_988 ( .A(_auto_iopadmap_cc_313_execute_56218_18_), .Y(\mc_addr_pad_o[18] ) );
  BUFX2 BUFX2_989 ( .A(_auto_iopadmap_cc_313_execute_56218_19_), .Y(\mc_addr_pad_o[19] ) );
  BUFX2 BUFX2_99 ( .A(u2_u5__abc_47660_n137), .Y(u2_u5__abc_47660_n137_bF_buf1) );
  BUFX2 BUFX2_990 ( .A(_auto_iopadmap_cc_313_execute_56218_20_), .Y(\mc_addr_pad_o[20] ) );
  BUFX2 BUFX2_991 ( .A(_auto_iopadmap_cc_313_execute_56218_21_), .Y(\mc_addr_pad_o[21] ) );
  BUFX2 BUFX2_992 ( .A(_auto_iopadmap_cc_313_execute_56218_22_), .Y(\mc_addr_pad_o[22] ) );
  BUFX2 BUFX2_993 ( .A(_auto_iopadmap_cc_313_execute_56218_23_), .Y(\mc_addr_pad_o[23] ) );
  BUFX2 BUFX2_994 ( .A(_auto_iopadmap_cc_313_execute_56243), .Y(mc_adsc_pad_o_) );
  BUFX2 BUFX2_995 ( .A(_auto_iopadmap_cc_313_execute_56245), .Y(mc_adv_pad_o_) );
  BUFX2 BUFX2_996 ( .A(_auto_iopadmap_cc_313_execute_56247), .Y(mc_bg_pad_o) );
  BUFX2 BUFX2_997 ( .A(_auto_iopadmap_cc_313_execute_56249), .Y(mc_cas_pad_o_) );
  BUFX2 BUFX2_998 ( .A(_auto_iopadmap_cc_313_execute_56251), .Y(mc_cke_pad_o_) );
  BUFX2 BUFX2_999 ( .A(_auto_iopadmap_cc_313_execute_56253), .Y(mc_coe_pad_coe_o) );
  DFFPOSX1 DFFPOSX1_1 ( .CLK(clk_i_bF_buf125), .D(mem_ack), .Q(mem_ack_r) );
  DFFPOSX1 DFFPOSX1_10 ( .CLK(clk_i_bF_buf116), .D(u0_poc_6__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56321_6_) );
  DFFPOSX1 DFFPOSX1_100 ( .CLK(clk_i_bF_buf24), .D(u0_u0_csc_26__FF_INPUT), .Q(u0_csc0_26_) );
  DFFPOSX1 DFFPOSX1_1000 ( .CLK(clk_i_bF_buf66), .D(u3_u0_r1_12__FF_INPUT), .Q(u3_u0_r1_12_) );
  DFFPOSX1 DFFPOSX1_1001 ( .CLK(clk_i_bF_buf65), .D(u3_u0_r1_13__FF_INPUT), .Q(u3_u0_r1_13_) );
  DFFPOSX1 DFFPOSX1_1002 ( .CLK(clk_i_bF_buf64), .D(u3_u0_r1_14__FF_INPUT), .Q(u3_u0_r1_14_) );
  DFFPOSX1 DFFPOSX1_1003 ( .CLK(clk_i_bF_buf63), .D(u3_u0_r1_15__FF_INPUT), .Q(u3_u0_r1_15_) );
  DFFPOSX1 DFFPOSX1_1004 ( .CLK(clk_i_bF_buf62), .D(u3_u0_r1_16__FF_INPUT), .Q(u3_u0_r1_16_) );
  DFFPOSX1 DFFPOSX1_1005 ( .CLK(clk_i_bF_buf61), .D(u3_u0_r1_17__FF_INPUT), .Q(u3_u0_r1_17_) );
  DFFPOSX1 DFFPOSX1_1006 ( .CLK(clk_i_bF_buf60), .D(u3_u0_r1_18__FF_INPUT), .Q(u3_u0_r1_18_) );
  DFFPOSX1 DFFPOSX1_1007 ( .CLK(clk_i_bF_buf59), .D(u3_u0_r1_19__FF_INPUT), .Q(u3_u0_r1_19_) );
  DFFPOSX1 DFFPOSX1_1008 ( .CLK(clk_i_bF_buf58), .D(u3_u0_r1_20__FF_INPUT), .Q(u3_u0_r1_20_) );
  DFFPOSX1 DFFPOSX1_1009 ( .CLK(clk_i_bF_buf57), .D(u3_u0_r1_21__FF_INPUT), .Q(u3_u0_r1_21_) );
  DFFPOSX1 DFFPOSX1_101 ( .CLK(clk_i_bF_buf23), .D(u0_u0_csc_27__FF_INPUT), .Q(u0_csc0_27_) );
  DFFPOSX1 DFFPOSX1_1010 ( .CLK(clk_i_bF_buf56), .D(u3_u0_r1_22__FF_INPUT), .Q(u3_u0_r1_22_) );
  DFFPOSX1 DFFPOSX1_1011 ( .CLK(clk_i_bF_buf55), .D(u3_u0_r1_23__FF_INPUT), .Q(u3_u0_r1_23_) );
  DFFPOSX1 DFFPOSX1_1012 ( .CLK(clk_i_bF_buf54), .D(u3_u0_r1_24__FF_INPUT), .Q(u3_u0_r1_24_) );
  DFFPOSX1 DFFPOSX1_1013 ( .CLK(clk_i_bF_buf53), .D(u3_u0_r1_25__FF_INPUT), .Q(u3_u0_r1_25_) );
  DFFPOSX1 DFFPOSX1_1014 ( .CLK(clk_i_bF_buf52), .D(u3_u0_r1_26__FF_INPUT), .Q(u3_u0_r1_26_) );
  DFFPOSX1 DFFPOSX1_1015 ( .CLK(clk_i_bF_buf51), .D(u3_u0_r1_27__FF_INPUT), .Q(u3_u0_r1_27_) );
  DFFPOSX1 DFFPOSX1_1016 ( .CLK(clk_i_bF_buf50), .D(u3_u0_r1_28__FF_INPUT), .Q(u3_u0_r1_28_) );
  DFFPOSX1 DFFPOSX1_1017 ( .CLK(clk_i_bF_buf49), .D(u3_u0_r1_29__FF_INPUT), .Q(u3_u0_r1_29_) );
  DFFPOSX1 DFFPOSX1_1018 ( .CLK(clk_i_bF_buf48), .D(u3_u0_r1_30__FF_INPUT), .Q(u3_u0_r1_30_) );
  DFFPOSX1 DFFPOSX1_1019 ( .CLK(clk_i_bF_buf47), .D(u3_u0_r1_31__FF_INPUT), .Q(u3_u0_r1_31_) );
  DFFPOSX1 DFFPOSX1_102 ( .CLK(clk_i_bF_buf22), .D(u0_u0_csc_28__FF_INPUT), .Q(u0_csc0_28_) );
  DFFPOSX1 DFFPOSX1_1020 ( .CLK(clk_i_bF_buf46), .D(u3_u0_r1_32__FF_INPUT), .Q(u3_u0_r1_32_) );
  DFFPOSX1 DFFPOSX1_1021 ( .CLK(clk_i_bF_buf45), .D(u3_u0_r1_33__FF_INPUT), .Q(u3_u0_r1_33_) );
  DFFPOSX1 DFFPOSX1_1022 ( .CLK(clk_i_bF_buf44), .D(u3_u0_r1_34__FF_INPUT), .Q(u3_u0_r1_34_) );
  DFFPOSX1 DFFPOSX1_1023 ( .CLK(clk_i_bF_buf43), .D(u3_u0_r1_35__FF_INPUT), .Q(u3_u0_r1_35_) );
  DFFPOSX1 DFFPOSX1_1024 ( .CLK(clk_i_bF_buf42), .D(u3_u0_r0_0__FF_INPUT), .Q(u3_u0_r0_0_) );
  DFFPOSX1 DFFPOSX1_1025 ( .CLK(clk_i_bF_buf41), .D(u3_u0_r0_1__FF_INPUT), .Q(u3_u0_r0_1_) );
  DFFPOSX1 DFFPOSX1_1026 ( .CLK(clk_i_bF_buf40), .D(u3_u0_r0_2__FF_INPUT), .Q(u3_u0_r0_2_) );
  DFFPOSX1 DFFPOSX1_1027 ( .CLK(clk_i_bF_buf39), .D(u3_u0_r0_3__FF_INPUT), .Q(u3_u0_r0_3_) );
  DFFPOSX1 DFFPOSX1_1028 ( .CLK(clk_i_bF_buf38), .D(u3_u0_r0_4__FF_INPUT), .Q(u3_u0_r0_4_) );
  DFFPOSX1 DFFPOSX1_1029 ( .CLK(clk_i_bF_buf37), .D(u3_u0_r0_5__FF_INPUT), .Q(u3_u0_r0_5_) );
  DFFPOSX1 DFFPOSX1_103 ( .CLK(clk_i_bF_buf21), .D(u0_u0_csc_29__FF_INPUT), .Q(u0_csc0_29_) );
  DFFPOSX1 DFFPOSX1_1030 ( .CLK(clk_i_bF_buf36), .D(u3_u0_r0_6__FF_INPUT), .Q(u3_u0_r0_6_) );
  DFFPOSX1 DFFPOSX1_1031 ( .CLK(clk_i_bF_buf35), .D(u3_u0_r0_7__FF_INPUT), .Q(u3_u0_r0_7_) );
  DFFPOSX1 DFFPOSX1_1032 ( .CLK(clk_i_bF_buf34), .D(u3_u0_r0_8__FF_INPUT), .Q(u3_u0_r0_8_) );
  DFFPOSX1 DFFPOSX1_1033 ( .CLK(clk_i_bF_buf33), .D(u3_u0_r0_9__FF_INPUT), .Q(u3_u0_r0_9_) );
  DFFPOSX1 DFFPOSX1_1034 ( .CLK(clk_i_bF_buf32), .D(u3_u0_r0_10__FF_INPUT), .Q(u3_u0_r0_10_) );
  DFFPOSX1 DFFPOSX1_1035 ( .CLK(clk_i_bF_buf31), .D(u3_u0_r0_11__FF_INPUT), .Q(u3_u0_r0_11_) );
  DFFPOSX1 DFFPOSX1_1036 ( .CLK(clk_i_bF_buf30), .D(u3_u0_r0_12__FF_INPUT), .Q(u3_u0_r0_12_) );
  DFFPOSX1 DFFPOSX1_1037 ( .CLK(clk_i_bF_buf29), .D(u3_u0_r0_13__FF_INPUT), .Q(u3_u0_r0_13_) );
  DFFPOSX1 DFFPOSX1_1038 ( .CLK(clk_i_bF_buf28), .D(u3_u0_r0_14__FF_INPUT), .Q(u3_u0_r0_14_) );
  DFFPOSX1 DFFPOSX1_1039 ( .CLK(clk_i_bF_buf27), .D(u3_u0_r0_15__FF_INPUT), .Q(u3_u0_r0_15_) );
  DFFPOSX1 DFFPOSX1_104 ( .CLK(clk_i_bF_buf20), .D(u0_u0_csc_30__FF_INPUT), .Q(u0_csc0_30_) );
  DFFPOSX1 DFFPOSX1_1040 ( .CLK(clk_i_bF_buf26), .D(u3_u0_r0_16__FF_INPUT), .Q(u3_u0_r0_16_) );
  DFFPOSX1 DFFPOSX1_1041 ( .CLK(clk_i_bF_buf25), .D(u3_u0_r0_17__FF_INPUT), .Q(u3_u0_r0_17_) );
  DFFPOSX1 DFFPOSX1_1042 ( .CLK(clk_i_bF_buf24), .D(u3_u0_r0_18__FF_INPUT), .Q(u3_u0_r0_18_) );
  DFFPOSX1 DFFPOSX1_1043 ( .CLK(clk_i_bF_buf23), .D(u3_u0_r0_19__FF_INPUT), .Q(u3_u0_r0_19_) );
  DFFPOSX1 DFFPOSX1_1044 ( .CLK(clk_i_bF_buf22), .D(u3_u0_r0_20__FF_INPUT), .Q(u3_u0_r0_20_) );
  DFFPOSX1 DFFPOSX1_1045 ( .CLK(clk_i_bF_buf21), .D(u3_u0_r0_21__FF_INPUT), .Q(u3_u0_r0_21_) );
  DFFPOSX1 DFFPOSX1_1046 ( .CLK(clk_i_bF_buf20), .D(u3_u0_r0_22__FF_INPUT), .Q(u3_u0_r0_22_) );
  DFFPOSX1 DFFPOSX1_1047 ( .CLK(clk_i_bF_buf19), .D(u3_u0_r0_23__FF_INPUT), .Q(u3_u0_r0_23_) );
  DFFPOSX1 DFFPOSX1_1048 ( .CLK(clk_i_bF_buf18), .D(u3_u0_r0_24__FF_INPUT), .Q(u3_u0_r0_24_) );
  DFFPOSX1 DFFPOSX1_1049 ( .CLK(clk_i_bF_buf17), .D(u3_u0_r0_25__FF_INPUT), .Q(u3_u0_r0_25_) );
  DFFPOSX1 DFFPOSX1_105 ( .CLK(clk_i_bF_buf19), .D(u0_u0_csc_31__FF_INPUT), .Q(u0_csc0_31_) );
  DFFPOSX1 DFFPOSX1_1050 ( .CLK(clk_i_bF_buf16), .D(u3_u0_r0_26__FF_INPUT), .Q(u3_u0_r0_26_) );
  DFFPOSX1 DFFPOSX1_1051 ( .CLK(clk_i_bF_buf15), .D(u3_u0_r0_27__FF_INPUT), .Q(u3_u0_r0_27_) );
  DFFPOSX1 DFFPOSX1_1052 ( .CLK(clk_i_bF_buf14), .D(u3_u0_r0_28__FF_INPUT), .Q(u3_u0_r0_28_) );
  DFFPOSX1 DFFPOSX1_1053 ( .CLK(clk_i_bF_buf13), .D(u3_u0_r0_29__FF_INPUT), .Q(u3_u0_r0_29_) );
  DFFPOSX1 DFFPOSX1_1054 ( .CLK(clk_i_bF_buf12), .D(u3_u0_r0_30__FF_INPUT), .Q(u3_u0_r0_30_) );
  DFFPOSX1 DFFPOSX1_1055 ( .CLK(clk_i_bF_buf11), .D(u3_u0_r0_31__FF_INPUT), .Q(u3_u0_r0_31_) );
  DFFPOSX1 DFFPOSX1_1056 ( .CLK(clk_i_bF_buf10), .D(u3_u0_r0_32__FF_INPUT), .Q(u3_u0_r0_32_) );
  DFFPOSX1 DFFPOSX1_1057 ( .CLK(clk_i_bF_buf9), .D(u3_u0_r0_33__FF_INPUT), .Q(u3_u0_r0_33_) );
  DFFPOSX1 DFFPOSX1_1058 ( .CLK(clk_i_bF_buf8), .D(u3_u0_r0_34__FF_INPUT), .Q(u3_u0_r0_34_) );
  DFFPOSX1 DFFPOSX1_1059 ( .CLK(clk_i_bF_buf7), .D(u3_u0_r0_35__FF_INPUT), .Q(u3_u0_r0_35_) );
  DFFPOSX1 DFFPOSX1_106 ( .CLK(clk_i_bF_buf18), .D(\wb_addr_i[2] ), .Q(u0_u0_addr_r_2_) );
  DFFPOSX1 DFFPOSX1_1060 ( .CLK(clk_i_bF_buf124), .D(u4_rfr_clr_FF_INPUT), .Q(u4_rfr_clr) );
  DFFPOSX1 DFFPOSX1_1061 ( .CLK(clk_i_bF_buf103), .D(u1_wb_write_go), .Q(u5_wb_write_go_r) );
  DFFPOSX1 DFFPOSX1_1062 ( .CLK(clk_i_bF_buf102), .D(cmd_a10), .Q(u5_cmd_a10_r) );
  DFFPOSX1 DFFPOSX1_1063 ( .CLK(clk_i_bF_buf101), .D(u5_burst_act_rd_FF_INPUT), .Q(u5_burst_act_rd) );
  DFFPOSX1 DFFPOSX1_1064 ( .CLK(clk_i_bF_buf100), .D(u5_burst_cnt_0__FF_INPUT), .Q(u5_burst_cnt_0_) );
  DFFPOSX1 DFFPOSX1_1065 ( .CLK(clk_i_bF_buf99), .D(u5_burst_cnt_1__FF_INPUT), .Q(u5_burst_cnt_1_) );
  DFFPOSX1 DFFPOSX1_1066 ( .CLK(clk_i_bF_buf98), .D(u5_burst_cnt_2__FF_INPUT), .Q(u5_burst_cnt_2_) );
  DFFPOSX1 DFFPOSX1_1067 ( .CLK(clk_i_bF_buf97), .D(u5_burst_cnt_3__FF_INPUT), .Q(u5_burst_cnt_3_) );
  DFFPOSX1 DFFPOSX1_1068 ( .CLK(clk_i_bF_buf96), .D(u5_burst_cnt_4__FF_INPUT), .Q(u5_burst_cnt_4_) );
  DFFPOSX1 DFFPOSX1_1069 ( .CLK(clk_i_bF_buf95), .D(u5_burst_cnt_5__FF_INPUT), .Q(u5_burst_cnt_5_) );
  DFFPOSX1 DFFPOSX1_107 ( .CLK(clk_i_bF_buf17), .D(\wb_addr_i[3] ), .Q(u0_u0_addr_r_3_) );
  DFFPOSX1 DFFPOSX1_1070 ( .CLK(clk_i_bF_buf94), .D(u5_burst_cnt_6__FF_INPUT), .Q(u5_burst_cnt_6_) );
  DFFPOSX1 DFFPOSX1_1071 ( .CLK(clk_i_bF_buf93), .D(u5_burst_cnt_7__FF_INPUT), .Q(u5_burst_cnt_7_) );
  DFFPOSX1 DFFPOSX1_1072 ( .CLK(clk_i_bF_buf92), .D(u5_burst_cnt_8__FF_INPUT), .Q(u5_burst_cnt_8_) );
  DFFPOSX1 DFFPOSX1_1073 ( .CLK(clk_i_bF_buf91), .D(u5_burst_cnt_9__FF_INPUT), .Q(u5_burst_cnt_9_) );
  DFFPOSX1 DFFPOSX1_1074 ( .CLK(clk_i_bF_buf90), .D(u5_burst_cnt_10__FF_INPUT), .Q(u5_burst_cnt_10_) );
  DFFPOSX1 DFFPOSX1_1075 ( .CLK(clk_i_bF_buf89), .D(u5_ir_cnt_done_FF_INPUT), .Q(u5_ir_cnt_done) );
  DFFPOSX1 DFFPOSX1_1076 ( .CLK(clk_i_bF_buf88), .D(u5_ir_cnt_0__FF_INPUT), .Q(u5_ir_cnt_0_) );
  DFFPOSX1 DFFPOSX1_1077 ( .CLK(clk_i_bF_buf87), .D(u5_ir_cnt_1__FF_INPUT), .Q(u5_ir_cnt_1_) );
  DFFPOSX1 DFFPOSX1_1078 ( .CLK(clk_i_bF_buf86), .D(u5_ir_cnt_2__FF_INPUT), .Q(u5_ir_cnt_2_) );
  DFFPOSX1 DFFPOSX1_1079 ( .CLK(clk_i_bF_buf85), .D(u5_ir_cnt_3__FF_INPUT), .Q(u5_ir_cnt_3_) );
  DFFPOSX1 DFFPOSX1_108 ( .CLK(clk_i_bF_buf16), .D(\wb_addr_i[4] ), .Q(u0_u0_addr_r_4_) );
  DFFPOSX1 DFFPOSX1_1080 ( .CLK(clk_i_bF_buf84), .D(u5_timer2_0__FF_INPUT), .Q(u5_timer2_0_) );
  DFFPOSX1 DFFPOSX1_1081 ( .CLK(clk_i_bF_buf83), .D(u5_timer2_1__FF_INPUT), .Q(u5_timer2_1_) );
  DFFPOSX1 DFFPOSX1_1082 ( .CLK(clk_i_bF_buf82), .D(u5_timer2_2__FF_INPUT), .Q(u5_timer2_2_) );
  DFFPOSX1 DFFPOSX1_1083 ( .CLK(clk_i_bF_buf81), .D(u5_timer2_3__FF_INPUT), .Q(u5_timer2_3_) );
  DFFPOSX1 DFFPOSX1_1084 ( .CLK(clk_i_bF_buf80), .D(u5_timer2_4__FF_INPUT), .Q(u5_timer2_4_) );
  DFFPOSX1 DFFPOSX1_1085 ( .CLK(clk_i_bF_buf79), .D(u5_timer2_5__FF_INPUT), .Q(u5_timer2_5_) );
  DFFPOSX1 DFFPOSX1_1086 ( .CLK(clk_i_bF_buf78), .D(u5_timer2_6__FF_INPUT), .Q(u5_timer2_6_) );
  DFFPOSX1 DFFPOSX1_1087 ( .CLK(clk_i_bF_buf77), .D(u5_timer2_7__FF_INPUT), .Q(u5_timer2_7_) );
  DFFPOSX1 DFFPOSX1_1088 ( .CLK(clk_i_bF_buf76), .D(u5_timer2_8__FF_INPUT), .Q(u5_timer2_8_) );
  DFFPOSX1 DFFPOSX1_1089 ( .CLK(clk_i_bF_buf75), .D(u5_cnt_next), .Q(u5_cnt) );
  DFFPOSX1 DFFPOSX1_109 ( .CLK(clk_i_bF_buf15), .D(\wb_addr_i[5] ), .Q(u0_u0_addr_r_5_) );
  DFFPOSX1 DFFPOSX1_1090 ( .CLK(clk_i_bF_buf74), .D(u5_wb_wait_r2), .Q(u5_wb_wait_r) );
  DFFPOSX1 DFFPOSX1_1091 ( .CLK(clk_i_bF_buf73), .D(u5_wb_wait), .Q(u5_wb_wait_r2) );
  DFFPOSX1 DFFPOSX1_1092 ( .CLK(clk_i_bF_buf72), .D(u5_cke_o_r2), .Q(u5_cke_o_del) );
  DFFPOSX1 DFFPOSX1_1093 ( .CLK(clk_i_bF_buf71), .D(u5_cke_o_r1), .Q(u5_cke_o_r2) );
  DFFPOSX1 DFFPOSX1_1094 ( .CLK(clk_i_bF_buf70), .D(_auto_iopadmap_cc_313_execute_56251), .Q(u5_cke_o_r1) );
  DFFPOSX1 DFFPOSX1_1095 ( .CLK(clk_i_bF_buf69), .D(u5_cke__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56251) );
  DFFPOSX1 DFFPOSX1_1096 ( .CLK(clk_i_bF_buf68), .D(u5_cke_d), .Q(u5_cke_r) );
  DFFPOSX1 DFFPOSX1_1097 ( .CLK(clk_i_bF_buf67), .D(u5_pack_le2_d), .Q(pack_le2) );
  DFFPOSX1 DFFPOSX1_1098 ( .CLK(clk_i_bF_buf66), .D(u5_pack_le1_d), .Q(pack_le1) );
  DFFPOSX1 DFFPOSX1_1099 ( .CLK(clk_i_bF_buf65), .D(u5_pack_le0_d), .Q(pack_le0) );
  DFFPOSX1 DFFPOSX1_11 ( .CLK(clk_i_bF_buf115), .D(u0_poc_7__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56321_7_) );
  DFFPOSX1 DFFPOSX1_110 ( .CLK(clk_i_bF_buf14), .D(\wb_addr_i[6] ), .Q(u0_u0_addr_r_6_) );
  DFFPOSX1 DFFPOSX1_1100 ( .CLK(clk_i_bF_buf64), .D(cs_le_d), .Q(cs_le) );
  DFFPOSX1 DFFPOSX1_1101 ( .CLK(clk_i_bF_buf63), .D(cs_le_bF_buf1), .Q(u5_cs_le_r1) );
  DFFPOSX1 DFFPOSX1_1102 ( .CLK(clk_i_bF_buf62), .D(u5_cs_le_r1), .Q(u5_cs_le_r) );
  DFFPOSX1 DFFPOSX1_1103 ( .CLK(clk_i_bF_buf61), .D(u5_lmr_ack_d), .Q(lmr_ack) );
  DFFPOSX1 DFFPOSX1_1104 ( .CLK(clk_i_bF_buf6), .D(u6_wb_data_o_0__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56358_0_) );
  DFFPOSX1 DFFPOSX1_1105 ( .CLK(clk_i_bF_buf5), .D(u6_wb_data_o_1__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56358_1_) );
  DFFPOSX1 DFFPOSX1_1106 ( .CLK(clk_i_bF_buf4), .D(u6_wb_data_o_2__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56358_2_) );
  DFFPOSX1 DFFPOSX1_1107 ( .CLK(clk_i_bF_buf3), .D(u6_wb_data_o_3__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56358_3_) );
  DFFPOSX1 DFFPOSX1_1108 ( .CLK(clk_i_bF_buf2), .D(u6_wb_data_o_4__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56358_4_) );
  DFFPOSX1 DFFPOSX1_1109 ( .CLK(clk_i_bF_buf1), .D(u6_wb_data_o_5__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56358_5_) );
  DFFPOSX1 DFFPOSX1_111 ( .CLK(clk_i_bF_buf6), .D(u0_u1_tms_0__FF_INPUT), .Q(u0_tms1_0_) );
  DFFPOSX1 DFFPOSX1_1110 ( .CLK(clk_i_bF_buf0), .D(u6_wb_data_o_6__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56358_6_) );
  DFFPOSX1 DFFPOSX1_1111 ( .CLK(clk_i_bF_buf125), .D(u6_wb_data_o_7__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56358_7_) );
  DFFPOSX1 DFFPOSX1_1112 ( .CLK(clk_i_bF_buf124), .D(u6_wb_data_o_8__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56358_8_) );
  DFFPOSX1 DFFPOSX1_1113 ( .CLK(clk_i_bF_buf123), .D(u6_wb_data_o_9__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56358_9_) );
  DFFPOSX1 DFFPOSX1_1114 ( .CLK(clk_i_bF_buf122), .D(u6_wb_data_o_10__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56358_10_) );
  DFFPOSX1 DFFPOSX1_1115 ( .CLK(clk_i_bF_buf121), .D(u6_wb_data_o_11__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56358_11_) );
  DFFPOSX1 DFFPOSX1_1116 ( .CLK(clk_i_bF_buf120), .D(u6_wb_data_o_12__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56358_12_) );
  DFFPOSX1 DFFPOSX1_1117 ( .CLK(clk_i_bF_buf119), .D(u6_wb_data_o_13__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56358_13_) );
  DFFPOSX1 DFFPOSX1_1118 ( .CLK(clk_i_bF_buf118), .D(u6_wb_data_o_14__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56358_14_) );
  DFFPOSX1 DFFPOSX1_1119 ( .CLK(clk_i_bF_buf117), .D(u6_wb_data_o_15__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56358_15_) );
  DFFPOSX1 DFFPOSX1_112 ( .CLK(clk_i_bF_buf5), .D(u0_u1_tms_1__FF_INPUT), .Q(u0_tms1_1_) );
  DFFPOSX1 DFFPOSX1_1120 ( .CLK(clk_i_bF_buf116), .D(u6_wb_data_o_16__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56358_16_) );
  DFFPOSX1 DFFPOSX1_1121 ( .CLK(clk_i_bF_buf115), .D(u6_wb_data_o_17__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56358_17_) );
  DFFPOSX1 DFFPOSX1_1122 ( .CLK(clk_i_bF_buf114), .D(u6_wb_data_o_18__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56358_18_) );
  DFFPOSX1 DFFPOSX1_1123 ( .CLK(clk_i_bF_buf113), .D(u6_wb_data_o_19__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56358_19_) );
  DFFPOSX1 DFFPOSX1_1124 ( .CLK(clk_i_bF_buf112), .D(u6_wb_data_o_20__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56358_20_) );
  DFFPOSX1 DFFPOSX1_1125 ( .CLK(clk_i_bF_buf111), .D(u6_wb_data_o_21__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56358_21_) );
  DFFPOSX1 DFFPOSX1_1126 ( .CLK(clk_i_bF_buf110), .D(u6_wb_data_o_22__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56358_22_) );
  DFFPOSX1 DFFPOSX1_1127 ( .CLK(clk_i_bF_buf109), .D(u6_wb_data_o_23__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56358_23_) );
  DFFPOSX1 DFFPOSX1_1128 ( .CLK(clk_i_bF_buf108), .D(u6_wb_data_o_24__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56358_24_) );
  DFFPOSX1 DFFPOSX1_1129 ( .CLK(clk_i_bF_buf107), .D(u6_wb_data_o_25__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56358_25_) );
  DFFPOSX1 DFFPOSX1_113 ( .CLK(clk_i_bF_buf4), .D(u0_u1_tms_2__FF_INPUT), .Q(u0_tms1_2_) );
  DFFPOSX1 DFFPOSX1_1130 ( .CLK(clk_i_bF_buf106), .D(u6_wb_data_o_26__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56358_26_) );
  DFFPOSX1 DFFPOSX1_1131 ( .CLK(clk_i_bF_buf105), .D(u6_wb_data_o_27__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56358_27_) );
  DFFPOSX1 DFFPOSX1_1132 ( .CLK(clk_i_bF_buf104), .D(u6_wb_data_o_28__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56358_28_) );
  DFFPOSX1 DFFPOSX1_1133 ( .CLK(clk_i_bF_buf103), .D(u6_wb_data_o_29__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56358_29_) );
  DFFPOSX1 DFFPOSX1_1134 ( .CLK(clk_i_bF_buf102), .D(u6_wb_data_o_30__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56358_30_) );
  DFFPOSX1 DFFPOSX1_1135 ( .CLK(clk_i_bF_buf101), .D(u6_wb_data_o_31__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56358_31_) );
  DFFPOSX1 DFFPOSX1_1136 ( .CLK(mc_clk_i_bF_buf9), .D(u7_mc_adv__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56245) );
  DFFPOSX1 DFFPOSX1_1137 ( .CLK(mc_clk_i_bF_buf8), .D(u7_mc_adsc__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56243) );
  DFFPOSX1 DFFPOSX1_1138 ( .CLK(mc_clk_i_bF_buf7), .D(ras_), .Q(_auto_iopadmap_cc_313_execute_56311) );
  DFFPOSX1 DFFPOSX1_1139 ( .CLK(mc_clk_i_bF_buf6), .D(cas_), .Q(_auto_iopadmap_cc_313_execute_56249) );
  DFFPOSX1 DFFPOSX1_114 ( .CLK(clk_i_bF_buf3), .D(u0_u1_tms_3__FF_INPUT), .Q(u0_tms1_3_) );
  DFFPOSX1 DFFPOSX1_1140 ( .CLK(mc_clk_i_bF_buf5), .D(u5_we_), .Q(_auto_iopadmap_cc_313_execute_56317) );
  DFFPOSX1 DFFPOSX1_1141 ( .CLK(mc_clk_i_bF_buf4), .D(u7_mc_dqm_0__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56304_0_) );
  DFFPOSX1 DFFPOSX1_1142 ( .CLK(mc_clk_i_bF_buf3), .D(u7_mc_dqm_1__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56304_1_) );
  DFFPOSX1 DFFPOSX1_1143 ( .CLK(mc_clk_i_bF_buf2), .D(u7_mc_dqm_2__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56304_2_) );
  DFFPOSX1 DFFPOSX1_1144 ( .CLK(mc_clk_i_bF_buf1), .D(u7_mc_dqm_3__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56304_3_) );
  DFFPOSX1 DFFPOSX1_1145 ( .CLK(clk_i_bF_buf90), .D(u7_mc_dqm_r_0_), .Q(u7_mc_dqm_r2_0_) );
  DFFPOSX1 DFFPOSX1_1146 ( .CLK(clk_i_bF_buf89), .D(u7_mc_dqm_r_1_), .Q(u7_mc_dqm_r2_1_) );
  DFFPOSX1 DFFPOSX1_1147 ( .CLK(clk_i_bF_buf88), .D(u7_mc_dqm_r_2_), .Q(u7_mc_dqm_r2_2_) );
  DFFPOSX1 DFFPOSX1_1148 ( .CLK(clk_i_bF_buf87), .D(u7_mc_dqm_r_3_), .Q(u7_mc_dqm_r2_3_) );
  DFFPOSX1 DFFPOSX1_1149 ( .CLK(clk_i_bF_buf86), .D(u7_mc_dqm_r_0__FF_INPUT), .Q(u7_mc_dqm_r_0_) );
  DFFPOSX1 DFFPOSX1_115 ( .CLK(clk_i_bF_buf2), .D(u0_u1_tms_4__FF_INPUT), .Q(u0_tms1_4_) );
  DFFPOSX1 DFFPOSX1_1150 ( .CLK(clk_i_bF_buf85), .D(u7_mc_dqm_r_1__FF_INPUT), .Q(u7_mc_dqm_r_1_) );
  DFFPOSX1 DFFPOSX1_1151 ( .CLK(clk_i_bF_buf84), .D(u7_mc_dqm_r_2__FF_INPUT), .Q(u7_mc_dqm_r_2_) );
  DFFPOSX1 DFFPOSX1_1152 ( .CLK(clk_i_bF_buf83), .D(u7_mc_dqm_r_3__FF_INPUT), .Q(u7_mc_dqm_r_3_) );
  DFFPOSX1 DFFPOSX1_1153 ( .CLK(mc_clk_i_bF_buf0), .D(mc_addr_d_0_), .Q(_auto_iopadmap_cc_313_execute_56218_0_) );
  DFFPOSX1 DFFPOSX1_1154 ( .CLK(mc_clk_i_bF_buf10), .D(mc_addr_d_1_), .Q(_auto_iopadmap_cc_313_execute_56218_1_) );
  DFFPOSX1 DFFPOSX1_1155 ( .CLK(mc_clk_i_bF_buf9), .D(mc_addr_d_2_), .Q(_auto_iopadmap_cc_313_execute_56218_2_) );
  DFFPOSX1 DFFPOSX1_1156 ( .CLK(mc_clk_i_bF_buf8), .D(mc_addr_d_3_), .Q(_auto_iopadmap_cc_313_execute_56218_3_) );
  DFFPOSX1 DFFPOSX1_1157 ( .CLK(mc_clk_i_bF_buf7), .D(mc_addr_d_4_), .Q(_auto_iopadmap_cc_313_execute_56218_4_) );
  DFFPOSX1 DFFPOSX1_1158 ( .CLK(mc_clk_i_bF_buf6), .D(mc_addr_d_5_), .Q(_auto_iopadmap_cc_313_execute_56218_5_) );
  DFFPOSX1 DFFPOSX1_1159 ( .CLK(mc_clk_i_bF_buf5), .D(mc_addr_d_6_), .Q(_auto_iopadmap_cc_313_execute_56218_6_) );
  DFFPOSX1 DFFPOSX1_116 ( .CLK(clk_i_bF_buf1), .D(u0_u1_tms_5__FF_INPUT), .Q(u0_tms1_5_) );
  DFFPOSX1 DFFPOSX1_1160 ( .CLK(mc_clk_i_bF_buf4), .D(mc_addr_d_7_), .Q(_auto_iopadmap_cc_313_execute_56218_7_) );
  DFFPOSX1 DFFPOSX1_1161 ( .CLK(mc_clk_i_bF_buf3), .D(mc_addr_d_8_), .Q(_auto_iopadmap_cc_313_execute_56218_8_) );
  DFFPOSX1 DFFPOSX1_1162 ( .CLK(mc_clk_i_bF_buf2), .D(mc_addr_d_9_), .Q(_auto_iopadmap_cc_313_execute_56218_9_) );
  DFFPOSX1 DFFPOSX1_1163 ( .CLK(mc_clk_i_bF_buf1), .D(mc_addr_d_10_), .Q(_auto_iopadmap_cc_313_execute_56218_10_) );
  DFFPOSX1 DFFPOSX1_1164 ( .CLK(mc_clk_i_bF_buf0), .D(mc_addr_d_11_), .Q(_auto_iopadmap_cc_313_execute_56218_11_) );
  DFFPOSX1 DFFPOSX1_1165 ( .CLK(mc_clk_i_bF_buf10), .D(mc_addr_d_12_), .Q(_auto_iopadmap_cc_313_execute_56218_12_) );
  DFFPOSX1 DFFPOSX1_1166 ( .CLK(mc_clk_i_bF_buf9), .D(mc_addr_d_13_), .Q(_auto_iopadmap_cc_313_execute_56218_13_) );
  DFFPOSX1 DFFPOSX1_1167 ( .CLK(mc_clk_i_bF_buf8), .D(mc_addr_d_14_), .Q(_auto_iopadmap_cc_313_execute_56218_14_) );
  DFFPOSX1 DFFPOSX1_1168 ( .CLK(mc_clk_i_bF_buf7), .D(mc_addr_d_15_), .Q(_auto_iopadmap_cc_313_execute_56218_15_) );
  DFFPOSX1 DFFPOSX1_1169 ( .CLK(mc_clk_i_bF_buf6), .D(mc_addr_d_16_), .Q(_auto_iopadmap_cc_313_execute_56218_16_) );
  DFFPOSX1 DFFPOSX1_117 ( .CLK(clk_i_bF_buf0), .D(u0_u1_tms_6__FF_INPUT), .Q(u0_tms1_6_) );
  DFFPOSX1 DFFPOSX1_1170 ( .CLK(mc_clk_i_bF_buf5), .D(mc_addr_d_17_), .Q(_auto_iopadmap_cc_313_execute_56218_17_) );
  DFFPOSX1 DFFPOSX1_1171 ( .CLK(mc_clk_i_bF_buf4), .D(mc_addr_d_18_), .Q(_auto_iopadmap_cc_313_execute_56218_18_) );
  DFFPOSX1 DFFPOSX1_1172 ( .CLK(mc_clk_i_bF_buf3), .D(mc_addr_d_19_), .Q(_auto_iopadmap_cc_313_execute_56218_19_) );
  DFFPOSX1 DFFPOSX1_1173 ( .CLK(mc_clk_i_bF_buf2), .D(mc_addr_d_20_), .Q(_auto_iopadmap_cc_313_execute_56218_20_) );
  DFFPOSX1 DFFPOSX1_1174 ( .CLK(mc_clk_i_bF_buf1), .D(mc_addr_d_21_), .Q(_auto_iopadmap_cc_313_execute_56218_21_) );
  DFFPOSX1 DFFPOSX1_1175 ( .CLK(mc_clk_i_bF_buf0), .D(mc_addr_d_22_), .Q(_auto_iopadmap_cc_313_execute_56218_22_) );
  DFFPOSX1 DFFPOSX1_1176 ( .CLK(mc_clk_i_bF_buf10), .D(mc_addr_d_23_), .Q(_auto_iopadmap_cc_313_execute_56218_23_) );
  DFFPOSX1 DFFPOSX1_1177 ( .CLK(mc_clk_i_bF_buf9), .D(mc_dp_od_0_), .Q(_auto_iopadmap_cc_313_execute_56299_0_) );
  DFFPOSX1 DFFPOSX1_1178 ( .CLK(mc_clk_i_bF_buf8), .D(mc_dp_od_1_), .Q(_auto_iopadmap_cc_313_execute_56299_1_) );
  DFFPOSX1 DFFPOSX1_1179 ( .CLK(mc_clk_i_bF_buf7), .D(mc_dp_od_2_), .Q(_auto_iopadmap_cc_313_execute_56299_2_) );
  DFFPOSX1 DFFPOSX1_118 ( .CLK(clk_i_bF_buf125), .D(u0_u1_tms_7__FF_INPUT), .Q(u0_tms1_7_) );
  DFFPOSX1 DFFPOSX1_1180 ( .CLK(mc_clk_i_bF_buf6), .D(mc_dp_od_3_), .Q(_auto_iopadmap_cc_313_execute_56299_3_) );
  DFFPOSX1 DFFPOSX1_1181 ( .CLK(mc_clk_i_bF_buf5), .D(mc_data_od_0_), .Q(_auto_iopadmap_cc_313_execute_56264_0_) );
  DFFPOSX1 DFFPOSX1_1182 ( .CLK(mc_clk_i_bF_buf4), .D(mc_data_od_1_), .Q(_auto_iopadmap_cc_313_execute_56264_1_) );
  DFFPOSX1 DFFPOSX1_1183 ( .CLK(mc_clk_i_bF_buf3), .D(mc_data_od_2_), .Q(_auto_iopadmap_cc_313_execute_56264_2_) );
  DFFPOSX1 DFFPOSX1_1184 ( .CLK(mc_clk_i_bF_buf2), .D(mc_data_od_3_), .Q(_auto_iopadmap_cc_313_execute_56264_3_) );
  DFFPOSX1 DFFPOSX1_1185 ( .CLK(mc_clk_i_bF_buf1), .D(mc_data_od_4_), .Q(_auto_iopadmap_cc_313_execute_56264_4_) );
  DFFPOSX1 DFFPOSX1_1186 ( .CLK(mc_clk_i_bF_buf0), .D(mc_data_od_5_), .Q(_auto_iopadmap_cc_313_execute_56264_5_) );
  DFFPOSX1 DFFPOSX1_1187 ( .CLK(mc_clk_i_bF_buf10), .D(mc_data_od_6_), .Q(_auto_iopadmap_cc_313_execute_56264_6_) );
  DFFPOSX1 DFFPOSX1_1188 ( .CLK(mc_clk_i_bF_buf9), .D(mc_data_od_7_), .Q(_auto_iopadmap_cc_313_execute_56264_7_) );
  DFFPOSX1 DFFPOSX1_1189 ( .CLK(mc_clk_i_bF_buf8), .D(mc_data_od_8_), .Q(_auto_iopadmap_cc_313_execute_56264_8_) );
  DFFPOSX1 DFFPOSX1_119 ( .CLK(clk_i_bF_buf124), .D(u0_u1_tms_8__FF_INPUT), .Q(u0_tms1_8_) );
  DFFPOSX1 DFFPOSX1_1190 ( .CLK(mc_clk_i_bF_buf7), .D(mc_data_od_9_), .Q(_auto_iopadmap_cc_313_execute_56264_9_) );
  DFFPOSX1 DFFPOSX1_1191 ( .CLK(mc_clk_i_bF_buf6), .D(mc_data_od_10_), .Q(_auto_iopadmap_cc_313_execute_56264_10_) );
  DFFPOSX1 DFFPOSX1_1192 ( .CLK(mc_clk_i_bF_buf5), .D(mc_data_od_11_), .Q(_auto_iopadmap_cc_313_execute_56264_11_) );
  DFFPOSX1 DFFPOSX1_1193 ( .CLK(mc_clk_i_bF_buf4), .D(mc_data_od_12_), .Q(_auto_iopadmap_cc_313_execute_56264_12_) );
  DFFPOSX1 DFFPOSX1_1194 ( .CLK(mc_clk_i_bF_buf3), .D(mc_data_od_13_), .Q(_auto_iopadmap_cc_313_execute_56264_13_) );
  DFFPOSX1 DFFPOSX1_1195 ( .CLK(mc_clk_i_bF_buf2), .D(mc_data_od_14_), .Q(_auto_iopadmap_cc_313_execute_56264_14_) );
  DFFPOSX1 DFFPOSX1_1196 ( .CLK(mc_clk_i_bF_buf1), .D(mc_data_od_15_), .Q(_auto_iopadmap_cc_313_execute_56264_15_) );
  DFFPOSX1 DFFPOSX1_1197 ( .CLK(mc_clk_i_bF_buf0), .D(mc_data_od_16_), .Q(_auto_iopadmap_cc_313_execute_56264_16_) );
  DFFPOSX1 DFFPOSX1_1198 ( .CLK(mc_clk_i_bF_buf10), .D(mc_data_od_17_), .Q(_auto_iopadmap_cc_313_execute_56264_17_) );
  DFFPOSX1 DFFPOSX1_1199 ( .CLK(mc_clk_i_bF_buf9), .D(mc_data_od_18_), .Q(_auto_iopadmap_cc_313_execute_56264_18_) );
  DFFPOSX1 DFFPOSX1_12 ( .CLK(clk_i_bF_buf114), .D(u0_poc_8__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56321_8_) );
  DFFPOSX1 DFFPOSX1_120 ( .CLK(clk_i_bF_buf123), .D(u0_u1_tms_9__FF_INPUT), .Q(u0_tms1_9_) );
  DFFPOSX1 DFFPOSX1_1200 ( .CLK(mc_clk_i_bF_buf8), .D(mc_data_od_19_), .Q(_auto_iopadmap_cc_313_execute_56264_19_) );
  DFFPOSX1 DFFPOSX1_1201 ( .CLK(mc_clk_i_bF_buf7), .D(mc_data_od_20_), .Q(_auto_iopadmap_cc_313_execute_56264_20_) );
  DFFPOSX1 DFFPOSX1_1202 ( .CLK(mc_clk_i_bF_buf6), .D(mc_data_od_21_), .Q(_auto_iopadmap_cc_313_execute_56264_21_) );
  DFFPOSX1 DFFPOSX1_1203 ( .CLK(mc_clk_i_bF_buf5), .D(mc_data_od_22_), .Q(_auto_iopadmap_cc_313_execute_56264_22_) );
  DFFPOSX1 DFFPOSX1_1204 ( .CLK(mc_clk_i_bF_buf4), .D(mc_data_od_23_), .Q(_auto_iopadmap_cc_313_execute_56264_23_) );
  DFFPOSX1 DFFPOSX1_1205 ( .CLK(mc_clk_i_bF_buf3), .D(mc_data_od_24_), .Q(_auto_iopadmap_cc_313_execute_56264_24_) );
  DFFPOSX1 DFFPOSX1_1206 ( .CLK(mc_clk_i_bF_buf2), .D(mc_data_od_25_), .Q(_auto_iopadmap_cc_313_execute_56264_25_) );
  DFFPOSX1 DFFPOSX1_1207 ( .CLK(mc_clk_i_bF_buf1), .D(mc_data_od_26_), .Q(_auto_iopadmap_cc_313_execute_56264_26_) );
  DFFPOSX1 DFFPOSX1_1208 ( .CLK(mc_clk_i_bF_buf0), .D(mc_data_od_27_), .Q(_auto_iopadmap_cc_313_execute_56264_27_) );
  DFFPOSX1 DFFPOSX1_1209 ( .CLK(mc_clk_i_bF_buf10), .D(mc_data_od_28_), .Q(_auto_iopadmap_cc_313_execute_56264_28_) );
  DFFPOSX1 DFFPOSX1_121 ( .CLK(clk_i_bF_buf122), .D(u0_u1_tms_10__FF_INPUT), .Q(u0_tms1_10_) );
  DFFPOSX1 DFFPOSX1_1210 ( .CLK(mc_clk_i_bF_buf9), .D(mc_data_od_29_), .Q(_auto_iopadmap_cc_313_execute_56264_29_) );
  DFFPOSX1 DFFPOSX1_1211 ( .CLK(mc_clk_i_bF_buf8), .D(mc_data_od_30_), .Q(_auto_iopadmap_cc_313_execute_56264_30_) );
  DFFPOSX1 DFFPOSX1_1212 ( .CLK(mc_clk_i_bF_buf7), .D(mc_data_od_31_), .Q(_auto_iopadmap_cc_313_execute_56264_31_) );
  DFFPOSX1 DFFPOSX1_1213 ( .CLK(mc_clk_i_bF_buf6), .D(mc_bg_d), .Q(_auto_iopadmap_cc_313_execute_56247) );
  DFFPOSX1 DFFPOSX1_1214 ( .CLK(mc_clk_i_bF_buf5), .D(mc_ack_pad_i), .Q(mc_ack_r) );
  DFFPOSX1 DFFPOSX1_1215 ( .CLK(mc_clk_i_bF_buf4), .D(mc_br_pad_i), .Q(mc_br_r) );
  DFFPOSX1 DFFPOSX1_1216 ( .CLK(mc_clk_i_bF_buf3), .D(u7_mc_rp_FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56313) );
  DFFPOSX1 DFFPOSX1_1217 ( .CLK(mc_clk_i_bF_buf2), .D(mc_c_oe_d), .Q(_auto_iopadmap_cc_313_execute_56253) );
  DFFPOSX1 DFFPOSX1_1218 ( .CLK(mc_clk_i_bF_buf1), .D(\mc_data_pad_i[0] ), .Q(mc_data_ir_0_) );
  DFFPOSX1 DFFPOSX1_1219 ( .CLK(mc_clk_i_bF_buf0), .D(\mc_data_pad_i[1] ), .Q(mc_data_ir_1_) );
  DFFPOSX1 DFFPOSX1_122 ( .CLK(clk_i_bF_buf121), .D(u0_u1_tms_11__FF_INPUT), .Q(u0_tms1_11_) );
  DFFPOSX1 DFFPOSX1_1220 ( .CLK(mc_clk_i_bF_buf10), .D(\mc_data_pad_i[2] ), .Q(mc_data_ir_2_) );
  DFFPOSX1 DFFPOSX1_1221 ( .CLK(mc_clk_i_bF_buf9), .D(\mc_data_pad_i[3] ), .Q(mc_data_ir_3_) );
  DFFPOSX1 DFFPOSX1_1222 ( .CLK(mc_clk_i_bF_buf8), .D(\mc_data_pad_i[4] ), .Q(mc_data_ir_4_) );
  DFFPOSX1 DFFPOSX1_1223 ( .CLK(mc_clk_i_bF_buf7), .D(\mc_data_pad_i[5] ), .Q(mc_data_ir_5_) );
  DFFPOSX1 DFFPOSX1_1224 ( .CLK(mc_clk_i_bF_buf6), .D(\mc_data_pad_i[6] ), .Q(mc_data_ir_6_) );
  DFFPOSX1 DFFPOSX1_1225 ( .CLK(mc_clk_i_bF_buf5), .D(\mc_data_pad_i[7] ), .Q(mc_data_ir_7_) );
  DFFPOSX1 DFFPOSX1_1226 ( .CLK(mc_clk_i_bF_buf4), .D(\mc_data_pad_i[8] ), .Q(mc_data_ir_8_) );
  DFFPOSX1 DFFPOSX1_1227 ( .CLK(mc_clk_i_bF_buf3), .D(\mc_data_pad_i[9] ), .Q(mc_data_ir_9_) );
  DFFPOSX1 DFFPOSX1_1228 ( .CLK(mc_clk_i_bF_buf2), .D(\mc_data_pad_i[10] ), .Q(mc_data_ir_10_) );
  DFFPOSX1 DFFPOSX1_1229 ( .CLK(mc_clk_i_bF_buf1), .D(\mc_data_pad_i[11] ), .Q(mc_data_ir_11_) );
  DFFPOSX1 DFFPOSX1_123 ( .CLK(clk_i_bF_buf120), .D(u0_u1_tms_12__FF_INPUT), .Q(u0_tms1_12_) );
  DFFPOSX1 DFFPOSX1_1230 ( .CLK(mc_clk_i_bF_buf0), .D(\mc_data_pad_i[12] ), .Q(mc_data_ir_12_) );
  DFFPOSX1 DFFPOSX1_1231 ( .CLK(mc_clk_i_bF_buf10), .D(\mc_data_pad_i[13] ), .Q(mc_data_ir_13_) );
  DFFPOSX1 DFFPOSX1_1232 ( .CLK(mc_clk_i_bF_buf9), .D(\mc_data_pad_i[14] ), .Q(mc_data_ir_14_) );
  DFFPOSX1 DFFPOSX1_1233 ( .CLK(mc_clk_i_bF_buf8), .D(\mc_data_pad_i[15] ), .Q(mc_data_ir_15_) );
  DFFPOSX1 DFFPOSX1_1234 ( .CLK(mc_clk_i_bF_buf7), .D(\mc_data_pad_i[16] ), .Q(mc_data_ir_16_) );
  DFFPOSX1 DFFPOSX1_1235 ( .CLK(mc_clk_i_bF_buf6), .D(\mc_data_pad_i[17] ), .Q(mc_data_ir_17_) );
  DFFPOSX1 DFFPOSX1_1236 ( .CLK(mc_clk_i_bF_buf5), .D(\mc_data_pad_i[18] ), .Q(mc_data_ir_18_) );
  DFFPOSX1 DFFPOSX1_1237 ( .CLK(mc_clk_i_bF_buf4), .D(\mc_data_pad_i[19] ), .Q(mc_data_ir_19_) );
  DFFPOSX1 DFFPOSX1_1238 ( .CLK(mc_clk_i_bF_buf3), .D(\mc_data_pad_i[20] ), .Q(mc_data_ir_20_) );
  DFFPOSX1 DFFPOSX1_1239 ( .CLK(mc_clk_i_bF_buf2), .D(\mc_data_pad_i[21] ), .Q(mc_data_ir_21_) );
  DFFPOSX1 DFFPOSX1_124 ( .CLK(clk_i_bF_buf119), .D(u0_u1_tms_13__FF_INPUT), .Q(u0_tms1_13_) );
  DFFPOSX1 DFFPOSX1_1240 ( .CLK(mc_clk_i_bF_buf1), .D(\mc_data_pad_i[22] ), .Q(mc_data_ir_22_) );
  DFFPOSX1 DFFPOSX1_1241 ( .CLK(mc_clk_i_bF_buf0), .D(\mc_data_pad_i[23] ), .Q(mc_data_ir_23_) );
  DFFPOSX1 DFFPOSX1_1242 ( .CLK(mc_clk_i_bF_buf10), .D(\mc_data_pad_i[24] ), .Q(mc_data_ir_24_) );
  DFFPOSX1 DFFPOSX1_1243 ( .CLK(mc_clk_i_bF_buf9), .D(\mc_data_pad_i[25] ), .Q(mc_data_ir_25_) );
  DFFPOSX1 DFFPOSX1_1244 ( .CLK(mc_clk_i_bF_buf8), .D(\mc_data_pad_i[26] ), .Q(mc_data_ir_26_) );
  DFFPOSX1 DFFPOSX1_1245 ( .CLK(mc_clk_i_bF_buf7), .D(\mc_data_pad_i[27] ), .Q(mc_data_ir_27_) );
  DFFPOSX1 DFFPOSX1_1246 ( .CLK(mc_clk_i_bF_buf6), .D(\mc_data_pad_i[28] ), .Q(mc_data_ir_28_) );
  DFFPOSX1 DFFPOSX1_1247 ( .CLK(mc_clk_i_bF_buf5), .D(\mc_data_pad_i[29] ), .Q(mc_data_ir_29_) );
  DFFPOSX1 DFFPOSX1_1248 ( .CLK(mc_clk_i_bF_buf4), .D(\mc_data_pad_i[30] ), .Q(mc_data_ir_30_) );
  DFFPOSX1 DFFPOSX1_1249 ( .CLK(mc_clk_i_bF_buf3), .D(\mc_data_pad_i[31] ), .Q(mc_data_ir_31_) );
  DFFPOSX1 DFFPOSX1_125 ( .CLK(clk_i_bF_buf118), .D(u0_u1_tms_14__FF_INPUT), .Q(u0_tms1_14_) );
  DFFPOSX1 DFFPOSX1_1250 ( .CLK(mc_clk_i_bF_buf2), .D(\mc_dp_pad_i[0] ), .Q(mc_data_ir_32_) );
  DFFPOSX1 DFFPOSX1_1251 ( .CLK(mc_clk_i_bF_buf1), .D(\mc_dp_pad_i[1] ), .Q(mc_data_ir_33_) );
  DFFPOSX1 DFFPOSX1_1252 ( .CLK(mc_clk_i_bF_buf0), .D(\mc_dp_pad_i[2] ), .Q(mc_data_ir_34_) );
  DFFPOSX1 DFFPOSX1_1253 ( .CLK(mc_clk_i_bF_buf10), .D(\mc_dp_pad_i[3] ), .Q(mc_data_ir_35_) );
  DFFPOSX1 DFFPOSX1_1254 ( .CLK(mc_clk_i_bF_buf9), .D(mc_sts_pad_i), .Q(mc_sts_ir) );
  DFFPOSX1 DFFPOSX1_1255 ( .CLK(mc_clk_i_bF_buf8), .D(_auto_iopadmap_cc_313_execute_56354), .Q(_auto_iopadmap_cc_313_execute_56319) );
  DFFPOSX1 DFFPOSX1_126 ( .CLK(clk_i_bF_buf117), .D(u0_u1_tms_15__FF_INPUT), .Q(u0_tms1_15_) );
  DFFPOSX1 DFFPOSX1_127 ( .CLK(clk_i_bF_buf116), .D(u0_u1_tms_16__FF_INPUT), .Q(u0_tms1_16_) );
  DFFPOSX1 DFFPOSX1_128 ( .CLK(clk_i_bF_buf115), .D(u0_u1_tms_17__FF_INPUT), .Q(u0_tms1_17_) );
  DFFPOSX1 DFFPOSX1_129 ( .CLK(clk_i_bF_buf114), .D(u0_u1_tms_18__FF_INPUT), .Q(u0_tms1_18_) );
  DFFPOSX1 DFFPOSX1_13 ( .CLK(clk_i_bF_buf113), .D(u0_poc_9__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56321_9_) );
  DFFPOSX1 DFFPOSX1_130 ( .CLK(clk_i_bF_buf113), .D(u0_u1_tms_19__FF_INPUT), .Q(u0_tms1_19_) );
  DFFPOSX1 DFFPOSX1_131 ( .CLK(clk_i_bF_buf112), .D(u0_u1_tms_20__FF_INPUT), .Q(u0_tms1_20_) );
  DFFPOSX1 DFFPOSX1_132 ( .CLK(clk_i_bF_buf111), .D(u0_u1_tms_21__FF_INPUT), .Q(u0_tms1_21_) );
  DFFPOSX1 DFFPOSX1_133 ( .CLK(clk_i_bF_buf110), .D(u0_u1_tms_22__FF_INPUT), .Q(u0_tms1_22_) );
  DFFPOSX1 DFFPOSX1_134 ( .CLK(clk_i_bF_buf109), .D(u0_u1_tms_23__FF_INPUT), .Q(u0_tms1_23_) );
  DFFPOSX1 DFFPOSX1_135 ( .CLK(clk_i_bF_buf108), .D(u0_u1_tms_24__FF_INPUT), .Q(u0_tms1_24_) );
  DFFPOSX1 DFFPOSX1_136 ( .CLK(clk_i_bF_buf107), .D(u0_u1_tms_25__FF_INPUT), .Q(u0_tms1_25_) );
  DFFPOSX1 DFFPOSX1_137 ( .CLK(clk_i_bF_buf106), .D(u0_u1_tms_26__FF_INPUT), .Q(u0_tms1_26_) );
  DFFPOSX1 DFFPOSX1_138 ( .CLK(clk_i_bF_buf105), .D(u0_u1_tms_27__FF_INPUT), .Q(u0_tms1_27_) );
  DFFPOSX1 DFFPOSX1_139 ( .CLK(clk_i_bF_buf104), .D(u0_u1_tms_28__FF_INPUT), .Q(u0_tms1_28_) );
  DFFPOSX1 DFFPOSX1_14 ( .CLK(clk_i_bF_buf112), .D(u0_poc_10__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56321_10_) );
  DFFPOSX1 DFFPOSX1_140 ( .CLK(clk_i_bF_buf103), .D(u0_u1_tms_29__FF_INPUT), .Q(u0_tms1_29_) );
  DFFPOSX1 DFFPOSX1_141 ( .CLK(clk_i_bF_buf102), .D(u0_u1_tms_30__FF_INPUT), .Q(u0_tms1_30_) );
  DFFPOSX1 DFFPOSX1_142 ( .CLK(clk_i_bF_buf101), .D(u0_u1_tms_31__FF_INPUT), .Q(u0_tms1_31_) );
  DFFPOSX1 DFFPOSX1_143 ( .CLK(clk_i_bF_buf100), .D(u0_u1_csc_0__FF_INPUT), .Q(u0_csc1_0_) );
  DFFPOSX1 DFFPOSX1_144 ( .CLK(clk_i_bF_buf99), .D(u0_u1_csc_1__FF_INPUT), .Q(u0_csc1_1_) );
  DFFPOSX1 DFFPOSX1_145 ( .CLK(clk_i_bF_buf98), .D(u0_u1_csc_2__FF_INPUT), .Q(u0_csc1_2_) );
  DFFPOSX1 DFFPOSX1_146 ( .CLK(clk_i_bF_buf97), .D(u0_u1_csc_3__FF_INPUT), .Q(u0_csc1_3_) );
  DFFPOSX1 DFFPOSX1_147 ( .CLK(clk_i_bF_buf96), .D(u0_u1_csc_4__FF_INPUT), .Q(u0_csc1_4_) );
  DFFPOSX1 DFFPOSX1_148 ( .CLK(clk_i_bF_buf95), .D(u0_u1_csc_5__FF_INPUT), .Q(u0_csc1_5_) );
  DFFPOSX1 DFFPOSX1_149 ( .CLK(clk_i_bF_buf94), .D(u0_u1_csc_6__FF_INPUT), .Q(u0_csc1_6_) );
  DFFPOSX1 DFFPOSX1_15 ( .CLK(clk_i_bF_buf111), .D(u0_poc_11__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56321_11_) );
  DFFPOSX1 DFFPOSX1_150 ( .CLK(clk_i_bF_buf93), .D(u0_u1_csc_7__FF_INPUT), .Q(u0_csc1_7_) );
  DFFPOSX1 DFFPOSX1_151 ( .CLK(clk_i_bF_buf92), .D(u0_u1_csc_8__FF_INPUT), .Q(u0_csc1_8_) );
  DFFPOSX1 DFFPOSX1_152 ( .CLK(clk_i_bF_buf91), .D(u0_u1_csc_9__FF_INPUT), .Q(u0_csc1_9_) );
  DFFPOSX1 DFFPOSX1_153 ( .CLK(clk_i_bF_buf90), .D(u0_u1_csc_10__FF_INPUT), .Q(u0_csc1_10_) );
  DFFPOSX1 DFFPOSX1_154 ( .CLK(clk_i_bF_buf89), .D(u0_u1_csc_11__FF_INPUT), .Q(u0_csc1_11_) );
  DFFPOSX1 DFFPOSX1_155 ( .CLK(clk_i_bF_buf88), .D(u0_u1_csc_12__FF_INPUT), .Q(u0_csc1_12_) );
  DFFPOSX1 DFFPOSX1_156 ( .CLK(clk_i_bF_buf87), .D(u0_u1_csc_13__FF_INPUT), .Q(u0_csc1_13_) );
  DFFPOSX1 DFFPOSX1_157 ( .CLK(clk_i_bF_buf86), .D(u0_u1_csc_14__FF_INPUT), .Q(u0_csc1_14_) );
  DFFPOSX1 DFFPOSX1_158 ( .CLK(clk_i_bF_buf85), .D(u0_u1_csc_15__FF_INPUT), .Q(u0_csc1_15_) );
  DFFPOSX1 DFFPOSX1_159 ( .CLK(clk_i_bF_buf84), .D(u0_u1_csc_16__FF_INPUT), .Q(u0_csc1_16_) );
  DFFPOSX1 DFFPOSX1_16 ( .CLK(clk_i_bF_buf110), .D(u0_poc_12__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56321_12_) );
  DFFPOSX1 DFFPOSX1_160 ( .CLK(clk_i_bF_buf83), .D(u0_u1_csc_17__FF_INPUT), .Q(u0_csc1_17_) );
  DFFPOSX1 DFFPOSX1_161 ( .CLK(clk_i_bF_buf82), .D(u0_u1_csc_18__FF_INPUT), .Q(u0_csc1_18_) );
  DFFPOSX1 DFFPOSX1_162 ( .CLK(clk_i_bF_buf81), .D(u0_u1_csc_19__FF_INPUT), .Q(u0_csc1_19_) );
  DFFPOSX1 DFFPOSX1_163 ( .CLK(clk_i_bF_buf80), .D(u0_u1_csc_20__FF_INPUT), .Q(u0_csc1_20_) );
  DFFPOSX1 DFFPOSX1_164 ( .CLK(clk_i_bF_buf79), .D(u0_u1_csc_21__FF_INPUT), .Q(u0_csc1_21_) );
  DFFPOSX1 DFFPOSX1_165 ( .CLK(clk_i_bF_buf78), .D(u0_u1_csc_22__FF_INPUT), .Q(u0_csc1_22_) );
  DFFPOSX1 DFFPOSX1_166 ( .CLK(clk_i_bF_buf77), .D(u0_u1_csc_23__FF_INPUT), .Q(u0_csc1_23_) );
  DFFPOSX1 DFFPOSX1_167 ( .CLK(clk_i_bF_buf76), .D(u0_u1_csc_24__FF_INPUT), .Q(u0_csc1_24_) );
  DFFPOSX1 DFFPOSX1_168 ( .CLK(clk_i_bF_buf75), .D(u0_u1_csc_25__FF_INPUT), .Q(u0_csc1_25_) );
  DFFPOSX1 DFFPOSX1_169 ( .CLK(clk_i_bF_buf74), .D(u0_u1_csc_26__FF_INPUT), .Q(u0_csc1_26_) );
  DFFPOSX1 DFFPOSX1_17 ( .CLK(clk_i_bF_buf109), .D(u0_poc_13__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56321_13_) );
  DFFPOSX1 DFFPOSX1_170 ( .CLK(clk_i_bF_buf73), .D(u0_u1_csc_27__FF_INPUT), .Q(u0_csc1_27_) );
  DFFPOSX1 DFFPOSX1_171 ( .CLK(clk_i_bF_buf72), .D(u0_u1_csc_28__FF_INPUT), .Q(u0_csc1_28_) );
  DFFPOSX1 DFFPOSX1_172 ( .CLK(clk_i_bF_buf71), .D(u0_u1_csc_29__FF_INPUT), .Q(u0_csc1_29_) );
  DFFPOSX1 DFFPOSX1_173 ( .CLK(clk_i_bF_buf70), .D(u0_u1_csc_30__FF_INPUT), .Q(u0_csc1_30_) );
  DFFPOSX1 DFFPOSX1_174 ( .CLK(clk_i_bF_buf69), .D(u0_u1_csc_31__FF_INPUT), .Q(u0_csc1_31_) );
  DFFPOSX1 DFFPOSX1_175 ( .CLK(clk_i_bF_buf68), .D(\wb_addr_i[2] ), .Q(u0_u1_addr_r_2_) );
  DFFPOSX1 DFFPOSX1_176 ( .CLK(clk_i_bF_buf67), .D(\wb_addr_i[3] ), .Q(u0_u1_addr_r_3_) );
  DFFPOSX1 DFFPOSX1_177 ( .CLK(clk_i_bF_buf66), .D(\wb_addr_i[4] ), .Q(u0_u1_addr_r_4_) );
  DFFPOSX1 DFFPOSX1_178 ( .CLK(clk_i_bF_buf65), .D(\wb_addr_i[5] ), .Q(u0_u1_addr_r_5_) );
  DFFPOSX1 DFFPOSX1_179 ( .CLK(clk_i_bF_buf64), .D(\wb_addr_i[6] ), .Q(u0_u1_addr_r_6_) );
  DFFPOSX1 DFFPOSX1_18 ( .CLK(clk_i_bF_buf108), .D(u0_poc_14__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56321_14_) );
  DFFPOSX1 DFFPOSX1_180 ( .CLK(clk_i_bF_buf56), .D(u0_u2_tms_0__FF_INPUT), .Q(u0_tms2_0_) );
  DFFPOSX1 DFFPOSX1_181 ( .CLK(clk_i_bF_buf55), .D(u0_u2_tms_1__FF_INPUT), .Q(u0_tms2_1_) );
  DFFPOSX1 DFFPOSX1_182 ( .CLK(clk_i_bF_buf54), .D(u0_u2_tms_2__FF_INPUT), .Q(u0_tms2_2_) );
  DFFPOSX1 DFFPOSX1_183 ( .CLK(clk_i_bF_buf53), .D(u0_u2_tms_3__FF_INPUT), .Q(u0_tms2_3_) );
  DFFPOSX1 DFFPOSX1_184 ( .CLK(clk_i_bF_buf52), .D(u0_u2_tms_4__FF_INPUT), .Q(u0_tms2_4_) );
  DFFPOSX1 DFFPOSX1_185 ( .CLK(clk_i_bF_buf51), .D(u0_u2_tms_5__FF_INPUT), .Q(u0_tms2_5_) );
  DFFPOSX1 DFFPOSX1_186 ( .CLK(clk_i_bF_buf50), .D(u0_u2_tms_6__FF_INPUT), .Q(u0_tms2_6_) );
  DFFPOSX1 DFFPOSX1_187 ( .CLK(clk_i_bF_buf49), .D(u0_u2_tms_7__FF_INPUT), .Q(u0_tms2_7_) );
  DFFPOSX1 DFFPOSX1_188 ( .CLK(clk_i_bF_buf48), .D(u0_u2_tms_8__FF_INPUT), .Q(u0_tms2_8_) );
  DFFPOSX1 DFFPOSX1_189 ( .CLK(clk_i_bF_buf47), .D(u0_u2_tms_9__FF_INPUT), .Q(u0_tms2_9_) );
  DFFPOSX1 DFFPOSX1_19 ( .CLK(clk_i_bF_buf107), .D(u0_poc_15__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56321_15_) );
  DFFPOSX1 DFFPOSX1_190 ( .CLK(clk_i_bF_buf46), .D(u0_u2_tms_10__FF_INPUT), .Q(u0_tms2_10_) );
  DFFPOSX1 DFFPOSX1_191 ( .CLK(clk_i_bF_buf45), .D(u0_u2_tms_11__FF_INPUT), .Q(u0_tms2_11_) );
  DFFPOSX1 DFFPOSX1_192 ( .CLK(clk_i_bF_buf44), .D(u0_u2_tms_12__FF_INPUT), .Q(u0_tms2_12_) );
  DFFPOSX1 DFFPOSX1_193 ( .CLK(clk_i_bF_buf43), .D(u0_u2_tms_13__FF_INPUT), .Q(u0_tms2_13_) );
  DFFPOSX1 DFFPOSX1_194 ( .CLK(clk_i_bF_buf42), .D(u0_u2_tms_14__FF_INPUT), .Q(u0_tms2_14_) );
  DFFPOSX1 DFFPOSX1_195 ( .CLK(clk_i_bF_buf41), .D(u0_u2_tms_15__FF_INPUT), .Q(u0_tms2_15_) );
  DFFPOSX1 DFFPOSX1_196 ( .CLK(clk_i_bF_buf40), .D(u0_u2_tms_16__FF_INPUT), .Q(u0_tms2_16_) );
  DFFPOSX1 DFFPOSX1_197 ( .CLK(clk_i_bF_buf39), .D(u0_u2_tms_17__FF_INPUT), .Q(u0_tms2_17_) );
  DFFPOSX1 DFFPOSX1_198 ( .CLK(clk_i_bF_buf38), .D(u0_u2_tms_18__FF_INPUT), .Q(u0_tms2_18_) );
  DFFPOSX1 DFFPOSX1_199 ( .CLK(clk_i_bF_buf37), .D(u0_u2_tms_19__FF_INPUT), .Q(u0_tms2_19_) );
  DFFPOSX1 DFFPOSX1_2 ( .CLK(clk_i_bF_buf124), .D(lmr_ack), .Q(u0_lmr_ack_r) );
  DFFPOSX1 DFFPOSX1_20 ( .CLK(clk_i_bF_buf106), .D(u0_poc_16__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56321_16_) );
  DFFPOSX1 DFFPOSX1_200 ( .CLK(clk_i_bF_buf36), .D(u0_u2_tms_20__FF_INPUT), .Q(u0_tms2_20_) );
  DFFPOSX1 DFFPOSX1_201 ( .CLK(clk_i_bF_buf35), .D(u0_u2_tms_21__FF_INPUT), .Q(u0_tms2_21_) );
  DFFPOSX1 DFFPOSX1_202 ( .CLK(clk_i_bF_buf34), .D(u0_u2_tms_22__FF_INPUT), .Q(u0_tms2_22_) );
  DFFPOSX1 DFFPOSX1_203 ( .CLK(clk_i_bF_buf33), .D(u0_u2_tms_23__FF_INPUT), .Q(u0_tms2_23_) );
  DFFPOSX1 DFFPOSX1_204 ( .CLK(clk_i_bF_buf32), .D(u0_u2_tms_24__FF_INPUT), .Q(u0_tms2_24_) );
  DFFPOSX1 DFFPOSX1_205 ( .CLK(clk_i_bF_buf31), .D(u0_u2_tms_25__FF_INPUT), .Q(u0_tms2_25_) );
  DFFPOSX1 DFFPOSX1_206 ( .CLK(clk_i_bF_buf30), .D(u0_u2_tms_26__FF_INPUT), .Q(u0_tms2_26_) );
  DFFPOSX1 DFFPOSX1_207 ( .CLK(clk_i_bF_buf29), .D(u0_u2_tms_27__FF_INPUT), .Q(u0_tms2_27_) );
  DFFPOSX1 DFFPOSX1_208 ( .CLK(clk_i_bF_buf28), .D(u0_u2_tms_28__FF_INPUT), .Q(u0_tms2_28_) );
  DFFPOSX1 DFFPOSX1_209 ( .CLK(clk_i_bF_buf27), .D(u0_u2_tms_29__FF_INPUT), .Q(u0_tms2_29_) );
  DFFPOSX1 DFFPOSX1_21 ( .CLK(clk_i_bF_buf105), .D(u0_poc_17__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56321_17_) );
  DFFPOSX1 DFFPOSX1_210 ( .CLK(clk_i_bF_buf26), .D(u0_u2_tms_30__FF_INPUT), .Q(u0_tms2_30_) );
  DFFPOSX1 DFFPOSX1_211 ( .CLK(clk_i_bF_buf25), .D(u0_u2_tms_31__FF_INPUT), .Q(u0_tms2_31_) );
  DFFPOSX1 DFFPOSX1_212 ( .CLK(clk_i_bF_buf24), .D(u0_u2_csc_0__FF_INPUT), .Q(u0_csc2_0_) );
  DFFPOSX1 DFFPOSX1_213 ( .CLK(clk_i_bF_buf23), .D(u0_u2_csc_1__FF_INPUT), .Q(u0_csc2_1_) );
  DFFPOSX1 DFFPOSX1_214 ( .CLK(clk_i_bF_buf22), .D(u0_u2_csc_2__FF_INPUT), .Q(u0_csc2_2_) );
  DFFPOSX1 DFFPOSX1_215 ( .CLK(clk_i_bF_buf21), .D(u0_u2_csc_3__FF_INPUT), .Q(u0_csc2_3_) );
  DFFPOSX1 DFFPOSX1_216 ( .CLK(clk_i_bF_buf20), .D(u0_u2_csc_4__FF_INPUT), .Q(u0_csc2_4_) );
  DFFPOSX1 DFFPOSX1_217 ( .CLK(clk_i_bF_buf19), .D(u0_u2_csc_5__FF_INPUT), .Q(u0_csc2_5_) );
  DFFPOSX1 DFFPOSX1_218 ( .CLK(clk_i_bF_buf18), .D(u0_u2_csc_6__FF_INPUT), .Q(u0_csc2_6_) );
  DFFPOSX1 DFFPOSX1_219 ( .CLK(clk_i_bF_buf17), .D(u0_u2_csc_7__FF_INPUT), .Q(u0_csc2_7_) );
  DFFPOSX1 DFFPOSX1_22 ( .CLK(clk_i_bF_buf104), .D(u0_poc_18__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56321_18_) );
  DFFPOSX1 DFFPOSX1_220 ( .CLK(clk_i_bF_buf16), .D(u0_u2_csc_8__FF_INPUT), .Q(u0_csc2_8_) );
  DFFPOSX1 DFFPOSX1_221 ( .CLK(clk_i_bF_buf15), .D(u0_u2_csc_9__FF_INPUT), .Q(u0_csc2_9_) );
  DFFPOSX1 DFFPOSX1_222 ( .CLK(clk_i_bF_buf14), .D(u0_u2_csc_10__FF_INPUT), .Q(u0_csc2_10_) );
  DFFPOSX1 DFFPOSX1_223 ( .CLK(clk_i_bF_buf13), .D(u0_u2_csc_11__FF_INPUT), .Q(u0_csc2_11_) );
  DFFPOSX1 DFFPOSX1_224 ( .CLK(clk_i_bF_buf12), .D(u0_u2_csc_12__FF_INPUT), .Q(u0_csc2_12_) );
  DFFPOSX1 DFFPOSX1_225 ( .CLK(clk_i_bF_buf11), .D(u0_u2_csc_13__FF_INPUT), .Q(u0_csc2_13_) );
  DFFPOSX1 DFFPOSX1_226 ( .CLK(clk_i_bF_buf10), .D(u0_u2_csc_14__FF_INPUT), .Q(u0_csc2_14_) );
  DFFPOSX1 DFFPOSX1_227 ( .CLK(clk_i_bF_buf9), .D(u0_u2_csc_15__FF_INPUT), .Q(u0_csc2_15_) );
  DFFPOSX1 DFFPOSX1_228 ( .CLK(clk_i_bF_buf8), .D(u0_u2_csc_16__FF_INPUT), .Q(u0_csc2_16_) );
  DFFPOSX1 DFFPOSX1_229 ( .CLK(clk_i_bF_buf7), .D(u0_u2_csc_17__FF_INPUT), .Q(u0_csc2_17_) );
  DFFPOSX1 DFFPOSX1_23 ( .CLK(clk_i_bF_buf103), .D(u0_poc_19__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56321_19_) );
  DFFPOSX1 DFFPOSX1_230 ( .CLK(clk_i_bF_buf6), .D(u0_u2_csc_18__FF_INPUT), .Q(u0_csc2_18_) );
  DFFPOSX1 DFFPOSX1_231 ( .CLK(clk_i_bF_buf5), .D(u0_u2_csc_19__FF_INPUT), .Q(u0_csc2_19_) );
  DFFPOSX1 DFFPOSX1_232 ( .CLK(clk_i_bF_buf4), .D(u0_u2_csc_20__FF_INPUT), .Q(u0_csc2_20_) );
  DFFPOSX1 DFFPOSX1_233 ( .CLK(clk_i_bF_buf3), .D(u0_u2_csc_21__FF_INPUT), .Q(u0_csc2_21_) );
  DFFPOSX1 DFFPOSX1_234 ( .CLK(clk_i_bF_buf2), .D(u0_u2_csc_22__FF_INPUT), .Q(u0_csc2_22_) );
  DFFPOSX1 DFFPOSX1_235 ( .CLK(clk_i_bF_buf1), .D(u0_u2_csc_23__FF_INPUT), .Q(u0_csc2_23_) );
  DFFPOSX1 DFFPOSX1_236 ( .CLK(clk_i_bF_buf0), .D(u0_u2_csc_24__FF_INPUT), .Q(u0_csc2_24_) );
  DFFPOSX1 DFFPOSX1_237 ( .CLK(clk_i_bF_buf125), .D(u0_u2_csc_25__FF_INPUT), .Q(u0_csc2_25_) );
  DFFPOSX1 DFFPOSX1_238 ( .CLK(clk_i_bF_buf124), .D(u0_u2_csc_26__FF_INPUT), .Q(u0_csc2_26_) );
  DFFPOSX1 DFFPOSX1_239 ( .CLK(clk_i_bF_buf123), .D(u0_u2_csc_27__FF_INPUT), .Q(u0_csc2_27_) );
  DFFPOSX1 DFFPOSX1_24 ( .CLK(clk_i_bF_buf102), .D(u0_poc_20__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56321_20_) );
  DFFPOSX1 DFFPOSX1_240 ( .CLK(clk_i_bF_buf122), .D(u0_u2_csc_28__FF_INPUT), .Q(u0_csc2_28_) );
  DFFPOSX1 DFFPOSX1_241 ( .CLK(clk_i_bF_buf121), .D(u0_u2_csc_29__FF_INPUT), .Q(u0_csc2_29_) );
  DFFPOSX1 DFFPOSX1_242 ( .CLK(clk_i_bF_buf120), .D(u0_u2_csc_30__FF_INPUT), .Q(u0_csc2_30_) );
  DFFPOSX1 DFFPOSX1_243 ( .CLK(clk_i_bF_buf119), .D(u0_u2_csc_31__FF_INPUT), .Q(u0_csc2_31_) );
  DFFPOSX1 DFFPOSX1_244 ( .CLK(clk_i_bF_buf118), .D(\wb_addr_i[2] ), .Q(u0_u2_addr_r_2_) );
  DFFPOSX1 DFFPOSX1_245 ( .CLK(clk_i_bF_buf117), .D(\wb_addr_i[3] ), .Q(u0_u2_addr_r_3_) );
  DFFPOSX1 DFFPOSX1_246 ( .CLK(clk_i_bF_buf116), .D(\wb_addr_i[4] ), .Q(u0_u2_addr_r_4_) );
  DFFPOSX1 DFFPOSX1_247 ( .CLK(clk_i_bF_buf115), .D(\wb_addr_i[5] ), .Q(u0_u2_addr_r_5_) );
  DFFPOSX1 DFFPOSX1_248 ( .CLK(clk_i_bF_buf114), .D(\wb_addr_i[6] ), .Q(u0_u2_addr_r_6_) );
  DFFPOSX1 DFFPOSX1_249 ( .CLK(clk_i_bF_buf106), .D(u0_u3_tms_0__FF_INPUT), .Q(u0_tms3_0_) );
  DFFPOSX1 DFFPOSX1_25 ( .CLK(clk_i_bF_buf101), .D(u0_poc_21__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56321_21_) );
  DFFPOSX1 DFFPOSX1_250 ( .CLK(clk_i_bF_buf105), .D(u0_u3_tms_1__FF_INPUT), .Q(u0_tms3_1_) );
  DFFPOSX1 DFFPOSX1_251 ( .CLK(clk_i_bF_buf104), .D(u0_u3_tms_2__FF_INPUT), .Q(u0_tms3_2_) );
  DFFPOSX1 DFFPOSX1_252 ( .CLK(clk_i_bF_buf103), .D(u0_u3_tms_3__FF_INPUT), .Q(u0_tms3_3_) );
  DFFPOSX1 DFFPOSX1_253 ( .CLK(clk_i_bF_buf102), .D(u0_u3_tms_4__FF_INPUT), .Q(u0_tms3_4_) );
  DFFPOSX1 DFFPOSX1_254 ( .CLK(clk_i_bF_buf101), .D(u0_u3_tms_5__FF_INPUT), .Q(u0_tms3_5_) );
  DFFPOSX1 DFFPOSX1_255 ( .CLK(clk_i_bF_buf100), .D(u0_u3_tms_6__FF_INPUT), .Q(u0_tms3_6_) );
  DFFPOSX1 DFFPOSX1_256 ( .CLK(clk_i_bF_buf99), .D(u0_u3_tms_7__FF_INPUT), .Q(u0_tms3_7_) );
  DFFPOSX1 DFFPOSX1_257 ( .CLK(clk_i_bF_buf98), .D(u0_u3_tms_8__FF_INPUT), .Q(u0_tms3_8_) );
  DFFPOSX1 DFFPOSX1_258 ( .CLK(clk_i_bF_buf97), .D(u0_u3_tms_9__FF_INPUT), .Q(u0_tms3_9_) );
  DFFPOSX1 DFFPOSX1_259 ( .CLK(clk_i_bF_buf96), .D(u0_u3_tms_10__FF_INPUT), .Q(u0_tms3_10_) );
  DFFPOSX1 DFFPOSX1_26 ( .CLK(clk_i_bF_buf100), .D(u0_poc_22__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56321_22_) );
  DFFPOSX1 DFFPOSX1_260 ( .CLK(clk_i_bF_buf95), .D(u0_u3_tms_11__FF_INPUT), .Q(u0_tms3_11_) );
  DFFPOSX1 DFFPOSX1_261 ( .CLK(clk_i_bF_buf94), .D(u0_u3_tms_12__FF_INPUT), .Q(u0_tms3_12_) );
  DFFPOSX1 DFFPOSX1_262 ( .CLK(clk_i_bF_buf93), .D(u0_u3_tms_13__FF_INPUT), .Q(u0_tms3_13_) );
  DFFPOSX1 DFFPOSX1_263 ( .CLK(clk_i_bF_buf92), .D(u0_u3_tms_14__FF_INPUT), .Q(u0_tms3_14_) );
  DFFPOSX1 DFFPOSX1_264 ( .CLK(clk_i_bF_buf91), .D(u0_u3_tms_15__FF_INPUT), .Q(u0_tms3_15_) );
  DFFPOSX1 DFFPOSX1_265 ( .CLK(clk_i_bF_buf90), .D(u0_u3_tms_16__FF_INPUT), .Q(u0_tms3_16_) );
  DFFPOSX1 DFFPOSX1_266 ( .CLK(clk_i_bF_buf89), .D(u0_u3_tms_17__FF_INPUT), .Q(u0_tms3_17_) );
  DFFPOSX1 DFFPOSX1_267 ( .CLK(clk_i_bF_buf88), .D(u0_u3_tms_18__FF_INPUT), .Q(u0_tms3_18_) );
  DFFPOSX1 DFFPOSX1_268 ( .CLK(clk_i_bF_buf87), .D(u0_u3_tms_19__FF_INPUT), .Q(u0_tms3_19_) );
  DFFPOSX1 DFFPOSX1_269 ( .CLK(clk_i_bF_buf86), .D(u0_u3_tms_20__FF_INPUT), .Q(u0_tms3_20_) );
  DFFPOSX1 DFFPOSX1_27 ( .CLK(clk_i_bF_buf99), .D(u0_poc_23__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56321_23_) );
  DFFPOSX1 DFFPOSX1_270 ( .CLK(clk_i_bF_buf85), .D(u0_u3_tms_21__FF_INPUT), .Q(u0_tms3_21_) );
  DFFPOSX1 DFFPOSX1_271 ( .CLK(clk_i_bF_buf84), .D(u0_u3_tms_22__FF_INPUT), .Q(u0_tms3_22_) );
  DFFPOSX1 DFFPOSX1_272 ( .CLK(clk_i_bF_buf83), .D(u0_u3_tms_23__FF_INPUT), .Q(u0_tms3_23_) );
  DFFPOSX1 DFFPOSX1_273 ( .CLK(clk_i_bF_buf82), .D(u0_u3_tms_24__FF_INPUT), .Q(u0_tms3_24_) );
  DFFPOSX1 DFFPOSX1_274 ( .CLK(clk_i_bF_buf81), .D(u0_u3_tms_25__FF_INPUT), .Q(u0_tms3_25_) );
  DFFPOSX1 DFFPOSX1_275 ( .CLK(clk_i_bF_buf80), .D(u0_u3_tms_26__FF_INPUT), .Q(u0_tms3_26_) );
  DFFPOSX1 DFFPOSX1_276 ( .CLK(clk_i_bF_buf79), .D(u0_u3_tms_27__FF_INPUT), .Q(u0_tms3_27_) );
  DFFPOSX1 DFFPOSX1_277 ( .CLK(clk_i_bF_buf78), .D(u0_u3_tms_28__FF_INPUT), .Q(u0_tms3_28_) );
  DFFPOSX1 DFFPOSX1_278 ( .CLK(clk_i_bF_buf77), .D(u0_u3_tms_29__FF_INPUT), .Q(u0_tms3_29_) );
  DFFPOSX1 DFFPOSX1_279 ( .CLK(clk_i_bF_buf76), .D(u0_u3_tms_30__FF_INPUT), .Q(u0_tms3_30_) );
  DFFPOSX1 DFFPOSX1_28 ( .CLK(clk_i_bF_buf98), .D(u0_poc_24__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56321_24_) );
  DFFPOSX1 DFFPOSX1_280 ( .CLK(clk_i_bF_buf75), .D(u0_u3_tms_31__FF_INPUT), .Q(u0_tms3_31_) );
  DFFPOSX1 DFFPOSX1_281 ( .CLK(clk_i_bF_buf74), .D(u0_u3_csc_0__FF_INPUT), .Q(u0_csc3_0_) );
  DFFPOSX1 DFFPOSX1_282 ( .CLK(clk_i_bF_buf73), .D(u0_u3_csc_1__FF_INPUT), .Q(u0_csc3_1_) );
  DFFPOSX1 DFFPOSX1_283 ( .CLK(clk_i_bF_buf72), .D(u0_u3_csc_2__FF_INPUT), .Q(u0_csc3_2_) );
  DFFPOSX1 DFFPOSX1_284 ( .CLK(clk_i_bF_buf71), .D(u0_u3_csc_3__FF_INPUT), .Q(u0_csc3_3_) );
  DFFPOSX1 DFFPOSX1_285 ( .CLK(clk_i_bF_buf70), .D(u0_u3_csc_4__FF_INPUT), .Q(u0_csc3_4_) );
  DFFPOSX1 DFFPOSX1_286 ( .CLK(clk_i_bF_buf69), .D(u0_u3_csc_5__FF_INPUT), .Q(u0_csc3_5_) );
  DFFPOSX1 DFFPOSX1_287 ( .CLK(clk_i_bF_buf68), .D(u0_u3_csc_6__FF_INPUT), .Q(u0_csc3_6_) );
  DFFPOSX1 DFFPOSX1_288 ( .CLK(clk_i_bF_buf67), .D(u0_u3_csc_7__FF_INPUT), .Q(u0_csc3_7_) );
  DFFPOSX1 DFFPOSX1_289 ( .CLK(clk_i_bF_buf66), .D(u0_u3_csc_8__FF_INPUT), .Q(u0_csc3_8_) );
  DFFPOSX1 DFFPOSX1_29 ( .CLK(clk_i_bF_buf97), .D(u0_poc_25__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56321_25_) );
  DFFPOSX1 DFFPOSX1_290 ( .CLK(clk_i_bF_buf65), .D(u0_u3_csc_9__FF_INPUT), .Q(u0_csc3_9_) );
  DFFPOSX1 DFFPOSX1_291 ( .CLK(clk_i_bF_buf64), .D(u0_u3_csc_10__FF_INPUT), .Q(u0_csc3_10_) );
  DFFPOSX1 DFFPOSX1_292 ( .CLK(clk_i_bF_buf63), .D(u0_u3_csc_11__FF_INPUT), .Q(u0_csc3_11_) );
  DFFPOSX1 DFFPOSX1_293 ( .CLK(clk_i_bF_buf62), .D(u0_u3_csc_12__FF_INPUT), .Q(u0_csc3_12_) );
  DFFPOSX1 DFFPOSX1_294 ( .CLK(clk_i_bF_buf61), .D(u0_u3_csc_13__FF_INPUT), .Q(u0_csc3_13_) );
  DFFPOSX1 DFFPOSX1_295 ( .CLK(clk_i_bF_buf60), .D(u0_u3_csc_14__FF_INPUT), .Q(u0_csc3_14_) );
  DFFPOSX1 DFFPOSX1_296 ( .CLK(clk_i_bF_buf59), .D(u0_u3_csc_15__FF_INPUT), .Q(u0_csc3_15_) );
  DFFPOSX1 DFFPOSX1_297 ( .CLK(clk_i_bF_buf58), .D(u0_u3_csc_16__FF_INPUT), .Q(u0_csc3_16_) );
  DFFPOSX1 DFFPOSX1_298 ( .CLK(clk_i_bF_buf57), .D(u0_u3_csc_17__FF_INPUT), .Q(u0_csc3_17_) );
  DFFPOSX1 DFFPOSX1_299 ( .CLK(clk_i_bF_buf56), .D(u0_u3_csc_18__FF_INPUT), .Q(u0_csc3_18_) );
  DFFPOSX1 DFFPOSX1_3 ( .CLK(clk_i_bF_buf123), .D(init_ack), .Q(u0_init_ack_r) );
  DFFPOSX1 DFFPOSX1_30 ( .CLK(clk_i_bF_buf96), .D(u0_poc_26__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56321_26_) );
  DFFPOSX1 DFFPOSX1_300 ( .CLK(clk_i_bF_buf55), .D(u0_u3_csc_19__FF_INPUT), .Q(u0_csc3_19_) );
  DFFPOSX1 DFFPOSX1_301 ( .CLK(clk_i_bF_buf54), .D(u0_u3_csc_20__FF_INPUT), .Q(u0_csc3_20_) );
  DFFPOSX1 DFFPOSX1_302 ( .CLK(clk_i_bF_buf53), .D(u0_u3_csc_21__FF_INPUT), .Q(u0_csc3_21_) );
  DFFPOSX1 DFFPOSX1_303 ( .CLK(clk_i_bF_buf52), .D(u0_u3_csc_22__FF_INPUT), .Q(u0_csc3_22_) );
  DFFPOSX1 DFFPOSX1_304 ( .CLK(clk_i_bF_buf51), .D(u0_u3_csc_23__FF_INPUT), .Q(u0_csc3_23_) );
  DFFPOSX1 DFFPOSX1_305 ( .CLK(clk_i_bF_buf50), .D(u0_u3_csc_24__FF_INPUT), .Q(u0_csc3_24_) );
  DFFPOSX1 DFFPOSX1_306 ( .CLK(clk_i_bF_buf49), .D(u0_u3_csc_25__FF_INPUT), .Q(u0_csc3_25_) );
  DFFPOSX1 DFFPOSX1_307 ( .CLK(clk_i_bF_buf48), .D(u0_u3_csc_26__FF_INPUT), .Q(u0_csc3_26_) );
  DFFPOSX1 DFFPOSX1_308 ( .CLK(clk_i_bF_buf47), .D(u0_u3_csc_27__FF_INPUT), .Q(u0_csc3_27_) );
  DFFPOSX1 DFFPOSX1_309 ( .CLK(clk_i_bF_buf46), .D(u0_u3_csc_28__FF_INPUT), .Q(u0_csc3_28_) );
  DFFPOSX1 DFFPOSX1_31 ( .CLK(clk_i_bF_buf95), .D(u0_poc_27__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56321_27_) );
  DFFPOSX1 DFFPOSX1_310 ( .CLK(clk_i_bF_buf45), .D(u0_u3_csc_29__FF_INPUT), .Q(u0_csc3_29_) );
  DFFPOSX1 DFFPOSX1_311 ( .CLK(clk_i_bF_buf44), .D(u0_u3_csc_30__FF_INPUT), .Q(u0_csc3_30_) );
  DFFPOSX1 DFFPOSX1_312 ( .CLK(clk_i_bF_buf43), .D(u0_u3_csc_31__FF_INPUT), .Q(u0_csc3_31_) );
  DFFPOSX1 DFFPOSX1_313 ( .CLK(clk_i_bF_buf42), .D(\wb_addr_i[2] ), .Q(u0_u3_addr_r_2_) );
  DFFPOSX1 DFFPOSX1_314 ( .CLK(clk_i_bF_buf41), .D(\wb_addr_i[3] ), .Q(u0_u3_addr_r_3_) );
  DFFPOSX1 DFFPOSX1_315 ( .CLK(clk_i_bF_buf40), .D(\wb_addr_i[4] ), .Q(u0_u3_addr_r_4_) );
  DFFPOSX1 DFFPOSX1_316 ( .CLK(clk_i_bF_buf39), .D(\wb_addr_i[5] ), .Q(u0_u3_addr_r_5_) );
  DFFPOSX1 DFFPOSX1_317 ( .CLK(clk_i_bF_buf38), .D(\wb_addr_i[6] ), .Q(u0_u3_addr_r_6_) );
  DFFPOSX1 DFFPOSX1_318 ( .CLK(clk_i_bF_buf30), .D(u0_u4_tms_0__FF_INPUT), .Q(u0_tms4_0_) );
  DFFPOSX1 DFFPOSX1_319 ( .CLK(clk_i_bF_buf29), .D(u0_u4_tms_1__FF_INPUT), .Q(u0_tms4_1_) );
  DFFPOSX1 DFFPOSX1_32 ( .CLK(clk_i_bF_buf94), .D(u0_poc_28__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56321_28_) );
  DFFPOSX1 DFFPOSX1_320 ( .CLK(clk_i_bF_buf28), .D(u0_u4_tms_2__FF_INPUT), .Q(u0_tms4_2_) );
  DFFPOSX1 DFFPOSX1_321 ( .CLK(clk_i_bF_buf27), .D(u0_u4_tms_3__FF_INPUT), .Q(u0_tms4_3_) );
  DFFPOSX1 DFFPOSX1_322 ( .CLK(clk_i_bF_buf26), .D(u0_u4_tms_4__FF_INPUT), .Q(u0_tms4_4_) );
  DFFPOSX1 DFFPOSX1_323 ( .CLK(clk_i_bF_buf25), .D(u0_u4_tms_5__FF_INPUT), .Q(u0_tms4_5_) );
  DFFPOSX1 DFFPOSX1_324 ( .CLK(clk_i_bF_buf24), .D(u0_u4_tms_6__FF_INPUT), .Q(u0_tms4_6_) );
  DFFPOSX1 DFFPOSX1_325 ( .CLK(clk_i_bF_buf23), .D(u0_u4_tms_7__FF_INPUT), .Q(u0_tms4_7_) );
  DFFPOSX1 DFFPOSX1_326 ( .CLK(clk_i_bF_buf22), .D(u0_u4_tms_8__FF_INPUT), .Q(u0_tms4_8_) );
  DFFPOSX1 DFFPOSX1_327 ( .CLK(clk_i_bF_buf21), .D(u0_u4_tms_9__FF_INPUT), .Q(u0_tms4_9_) );
  DFFPOSX1 DFFPOSX1_328 ( .CLK(clk_i_bF_buf20), .D(u0_u4_tms_10__FF_INPUT), .Q(u0_tms4_10_) );
  DFFPOSX1 DFFPOSX1_329 ( .CLK(clk_i_bF_buf19), .D(u0_u4_tms_11__FF_INPUT), .Q(u0_tms4_11_) );
  DFFPOSX1 DFFPOSX1_33 ( .CLK(clk_i_bF_buf93), .D(u0_poc_29__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56321_29_) );
  DFFPOSX1 DFFPOSX1_330 ( .CLK(clk_i_bF_buf18), .D(u0_u4_tms_12__FF_INPUT), .Q(u0_tms4_12_) );
  DFFPOSX1 DFFPOSX1_331 ( .CLK(clk_i_bF_buf17), .D(u0_u4_tms_13__FF_INPUT), .Q(u0_tms4_13_) );
  DFFPOSX1 DFFPOSX1_332 ( .CLK(clk_i_bF_buf16), .D(u0_u4_tms_14__FF_INPUT), .Q(u0_tms4_14_) );
  DFFPOSX1 DFFPOSX1_333 ( .CLK(clk_i_bF_buf15), .D(u0_u4_tms_15__FF_INPUT), .Q(u0_tms4_15_) );
  DFFPOSX1 DFFPOSX1_334 ( .CLK(clk_i_bF_buf14), .D(u0_u4_tms_16__FF_INPUT), .Q(u0_tms4_16_) );
  DFFPOSX1 DFFPOSX1_335 ( .CLK(clk_i_bF_buf13), .D(u0_u4_tms_17__FF_INPUT), .Q(u0_tms4_17_) );
  DFFPOSX1 DFFPOSX1_336 ( .CLK(clk_i_bF_buf12), .D(u0_u4_tms_18__FF_INPUT), .Q(u0_tms4_18_) );
  DFFPOSX1 DFFPOSX1_337 ( .CLK(clk_i_bF_buf11), .D(u0_u4_tms_19__FF_INPUT), .Q(u0_tms4_19_) );
  DFFPOSX1 DFFPOSX1_338 ( .CLK(clk_i_bF_buf10), .D(u0_u4_tms_20__FF_INPUT), .Q(u0_tms4_20_) );
  DFFPOSX1 DFFPOSX1_339 ( .CLK(clk_i_bF_buf9), .D(u0_u4_tms_21__FF_INPUT), .Q(u0_tms4_21_) );
  DFFPOSX1 DFFPOSX1_34 ( .CLK(clk_i_bF_buf92), .D(u0_poc_30__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56321_30_) );
  DFFPOSX1 DFFPOSX1_340 ( .CLK(clk_i_bF_buf8), .D(u0_u4_tms_22__FF_INPUT), .Q(u0_tms4_22_) );
  DFFPOSX1 DFFPOSX1_341 ( .CLK(clk_i_bF_buf7), .D(u0_u4_tms_23__FF_INPUT), .Q(u0_tms4_23_) );
  DFFPOSX1 DFFPOSX1_342 ( .CLK(clk_i_bF_buf6), .D(u0_u4_tms_24__FF_INPUT), .Q(u0_tms4_24_) );
  DFFPOSX1 DFFPOSX1_343 ( .CLK(clk_i_bF_buf5), .D(u0_u4_tms_25__FF_INPUT), .Q(u0_tms4_25_) );
  DFFPOSX1 DFFPOSX1_344 ( .CLK(clk_i_bF_buf4), .D(u0_u4_tms_26__FF_INPUT), .Q(u0_tms4_26_) );
  DFFPOSX1 DFFPOSX1_345 ( .CLK(clk_i_bF_buf3), .D(u0_u4_tms_27__FF_INPUT), .Q(u0_tms4_27_) );
  DFFPOSX1 DFFPOSX1_346 ( .CLK(clk_i_bF_buf2), .D(u0_u4_tms_28__FF_INPUT), .Q(u0_tms4_28_) );
  DFFPOSX1 DFFPOSX1_347 ( .CLK(clk_i_bF_buf1), .D(u0_u4_tms_29__FF_INPUT), .Q(u0_tms4_29_) );
  DFFPOSX1 DFFPOSX1_348 ( .CLK(clk_i_bF_buf0), .D(u0_u4_tms_30__FF_INPUT), .Q(u0_tms4_30_) );
  DFFPOSX1 DFFPOSX1_349 ( .CLK(clk_i_bF_buf125), .D(u0_u4_tms_31__FF_INPUT), .Q(u0_tms4_31_) );
  DFFPOSX1 DFFPOSX1_35 ( .CLK(clk_i_bF_buf91), .D(u0_poc_31__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56321_31_) );
  DFFPOSX1 DFFPOSX1_350 ( .CLK(clk_i_bF_buf124), .D(u0_u4_csc_0__FF_INPUT), .Q(u0_csc4_0_) );
  DFFPOSX1 DFFPOSX1_351 ( .CLK(clk_i_bF_buf123), .D(u0_u4_csc_1__FF_INPUT), .Q(u0_csc4_1_) );
  DFFPOSX1 DFFPOSX1_352 ( .CLK(clk_i_bF_buf122), .D(u0_u4_csc_2__FF_INPUT), .Q(u0_csc4_2_) );
  DFFPOSX1 DFFPOSX1_353 ( .CLK(clk_i_bF_buf121), .D(u0_u4_csc_3__FF_INPUT), .Q(u0_csc4_3_) );
  DFFPOSX1 DFFPOSX1_354 ( .CLK(clk_i_bF_buf120), .D(u0_u4_csc_4__FF_INPUT), .Q(u0_csc4_4_) );
  DFFPOSX1 DFFPOSX1_355 ( .CLK(clk_i_bF_buf119), .D(u0_u4_csc_5__FF_INPUT), .Q(u0_csc4_5_) );
  DFFPOSX1 DFFPOSX1_356 ( .CLK(clk_i_bF_buf118), .D(u0_u4_csc_6__FF_INPUT), .Q(u0_csc4_6_) );
  DFFPOSX1 DFFPOSX1_357 ( .CLK(clk_i_bF_buf117), .D(u0_u4_csc_7__FF_INPUT), .Q(u0_csc4_7_) );
  DFFPOSX1 DFFPOSX1_358 ( .CLK(clk_i_bF_buf116), .D(u0_u4_csc_8__FF_INPUT), .Q(u0_csc4_8_) );
  DFFPOSX1 DFFPOSX1_359 ( .CLK(clk_i_bF_buf115), .D(u0_u4_csc_9__FF_INPUT), .Q(u0_csc4_9_) );
  DFFPOSX1 DFFPOSX1_36 ( .CLK(clk_i_bF_buf90), .D(mc_sts_ir), .Q(u0_csr_0_) );
  DFFPOSX1 DFFPOSX1_360 ( .CLK(clk_i_bF_buf114), .D(u0_u4_csc_10__FF_INPUT), .Q(u0_csc4_10_) );
  DFFPOSX1 DFFPOSX1_361 ( .CLK(clk_i_bF_buf113), .D(u0_u4_csc_11__FF_INPUT), .Q(u0_csc4_11_) );
  DFFPOSX1 DFFPOSX1_362 ( .CLK(clk_i_bF_buf112), .D(u0_u4_csc_12__FF_INPUT), .Q(u0_csc4_12_) );
  DFFPOSX1 DFFPOSX1_363 ( .CLK(clk_i_bF_buf111), .D(u0_u4_csc_13__FF_INPUT), .Q(u0_csc4_13_) );
  DFFPOSX1 DFFPOSX1_364 ( .CLK(clk_i_bF_buf110), .D(u0_u4_csc_14__FF_INPUT), .Q(u0_csc4_14_) );
  DFFPOSX1 DFFPOSX1_365 ( .CLK(clk_i_bF_buf109), .D(u0_u4_csc_15__FF_INPUT), .Q(u0_csc4_15_) );
  DFFPOSX1 DFFPOSX1_366 ( .CLK(clk_i_bF_buf108), .D(u0_u4_csc_16__FF_INPUT), .Q(u0_csc4_16_) );
  DFFPOSX1 DFFPOSX1_367 ( .CLK(clk_i_bF_buf107), .D(u0_u4_csc_17__FF_INPUT), .Q(u0_csc4_17_) );
  DFFPOSX1 DFFPOSX1_368 ( .CLK(clk_i_bF_buf106), .D(u0_u4_csc_18__FF_INPUT), .Q(u0_csc4_18_) );
  DFFPOSX1 DFFPOSX1_369 ( .CLK(clk_i_bF_buf105), .D(u0_u4_csc_19__FF_INPUT), .Q(u0_csc4_19_) );
  DFFPOSX1 DFFPOSX1_37 ( .CLK(clk_i_bF_buf89), .D(\wb_addr_i[2] ), .Q(u0_wb_addr_r_2_) );
  DFFPOSX1 DFFPOSX1_370 ( .CLK(clk_i_bF_buf104), .D(u0_u4_csc_20__FF_INPUT), .Q(u0_csc4_20_) );
  DFFPOSX1 DFFPOSX1_371 ( .CLK(clk_i_bF_buf103), .D(u0_u4_csc_21__FF_INPUT), .Q(u0_csc4_21_) );
  DFFPOSX1 DFFPOSX1_372 ( .CLK(clk_i_bF_buf102), .D(u0_u4_csc_22__FF_INPUT), .Q(u0_csc4_22_) );
  DFFPOSX1 DFFPOSX1_373 ( .CLK(clk_i_bF_buf101), .D(u0_u4_csc_23__FF_INPUT), .Q(u0_csc4_23_) );
  DFFPOSX1 DFFPOSX1_374 ( .CLK(clk_i_bF_buf100), .D(u0_u4_csc_24__FF_INPUT), .Q(u0_csc4_24_) );
  DFFPOSX1 DFFPOSX1_375 ( .CLK(clk_i_bF_buf99), .D(u0_u4_csc_25__FF_INPUT), .Q(u0_csc4_25_) );
  DFFPOSX1 DFFPOSX1_376 ( .CLK(clk_i_bF_buf98), .D(u0_u4_csc_26__FF_INPUT), .Q(u0_csc4_26_) );
  DFFPOSX1 DFFPOSX1_377 ( .CLK(clk_i_bF_buf97), .D(u0_u4_csc_27__FF_INPUT), .Q(u0_csc4_27_) );
  DFFPOSX1 DFFPOSX1_378 ( .CLK(clk_i_bF_buf96), .D(u0_u4_csc_28__FF_INPUT), .Q(u0_csc4_28_) );
  DFFPOSX1 DFFPOSX1_379 ( .CLK(clk_i_bF_buf95), .D(u0_u4_csc_29__FF_INPUT), .Q(u0_csc4_29_) );
  DFFPOSX1 DFFPOSX1_38 ( .CLK(clk_i_bF_buf88), .D(\wb_addr_i[3] ), .Q(u0_wb_addr_r_3_) );
  DFFPOSX1 DFFPOSX1_380 ( .CLK(clk_i_bF_buf94), .D(u0_u4_csc_30__FF_INPUT), .Q(u0_csc4_30_) );
  DFFPOSX1 DFFPOSX1_381 ( .CLK(clk_i_bF_buf93), .D(u0_u4_csc_31__FF_INPUT), .Q(u0_csc4_31_) );
  DFFPOSX1 DFFPOSX1_382 ( .CLK(clk_i_bF_buf92), .D(\wb_addr_i[2] ), .Q(u0_u4_addr_r_2_) );
  DFFPOSX1 DFFPOSX1_383 ( .CLK(clk_i_bF_buf91), .D(\wb_addr_i[3] ), .Q(u0_u4_addr_r_3_) );
  DFFPOSX1 DFFPOSX1_384 ( .CLK(clk_i_bF_buf90), .D(\wb_addr_i[4] ), .Q(u0_u4_addr_r_4_) );
  DFFPOSX1 DFFPOSX1_385 ( .CLK(clk_i_bF_buf89), .D(\wb_addr_i[5] ), .Q(u0_u4_addr_r_5_) );
  DFFPOSX1 DFFPOSX1_386 ( .CLK(clk_i_bF_buf88), .D(\wb_addr_i[6] ), .Q(u0_u4_addr_r_6_) );
  DFFPOSX1 DFFPOSX1_387 ( .CLK(clk_i_bF_buf80), .D(u0_u5_tms_0__FF_INPUT), .Q(u0_tms5_0_) );
  DFFPOSX1 DFFPOSX1_388 ( .CLK(clk_i_bF_buf79), .D(u0_u5_tms_1__FF_INPUT), .Q(u0_tms5_1_) );
  DFFPOSX1 DFFPOSX1_389 ( .CLK(clk_i_bF_buf78), .D(u0_u5_tms_2__FF_INPUT), .Q(u0_tms5_2_) );
  DFFPOSX1 DFFPOSX1_39 ( .CLK(clk_i_bF_buf87), .D(\wb_addr_i[4] ), .Q(u0_wb_addr_r_4_) );
  DFFPOSX1 DFFPOSX1_390 ( .CLK(clk_i_bF_buf77), .D(u0_u5_tms_3__FF_INPUT), .Q(u0_tms5_3_) );
  DFFPOSX1 DFFPOSX1_391 ( .CLK(clk_i_bF_buf76), .D(u0_u5_tms_4__FF_INPUT), .Q(u0_tms5_4_) );
  DFFPOSX1 DFFPOSX1_392 ( .CLK(clk_i_bF_buf75), .D(u0_u5_tms_5__FF_INPUT), .Q(u0_tms5_5_) );
  DFFPOSX1 DFFPOSX1_393 ( .CLK(clk_i_bF_buf74), .D(u0_u5_tms_6__FF_INPUT), .Q(u0_tms5_6_) );
  DFFPOSX1 DFFPOSX1_394 ( .CLK(clk_i_bF_buf73), .D(u0_u5_tms_7__FF_INPUT), .Q(u0_tms5_7_) );
  DFFPOSX1 DFFPOSX1_395 ( .CLK(clk_i_bF_buf72), .D(u0_u5_tms_8__FF_INPUT), .Q(u0_tms5_8_) );
  DFFPOSX1 DFFPOSX1_396 ( .CLK(clk_i_bF_buf71), .D(u0_u5_tms_9__FF_INPUT), .Q(u0_tms5_9_) );
  DFFPOSX1 DFFPOSX1_397 ( .CLK(clk_i_bF_buf70), .D(u0_u5_tms_10__FF_INPUT), .Q(u0_tms5_10_) );
  DFFPOSX1 DFFPOSX1_398 ( .CLK(clk_i_bF_buf69), .D(u0_u5_tms_11__FF_INPUT), .Q(u0_tms5_11_) );
  DFFPOSX1 DFFPOSX1_399 ( .CLK(clk_i_bF_buf68), .D(u0_u5_tms_12__FF_INPUT), .Q(u0_tms5_12_) );
  DFFPOSX1 DFFPOSX1_4 ( .CLK(clk_i_bF_buf122), .D(u0_poc_0__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56321_0_) );
  DFFPOSX1 DFFPOSX1_40 ( .CLK(clk_i_bF_buf86), .D(\wb_addr_i[5] ), .Q(u0_wb_addr_r_5_) );
  DFFPOSX1 DFFPOSX1_400 ( .CLK(clk_i_bF_buf67), .D(u0_u5_tms_13__FF_INPUT), .Q(u0_tms5_13_) );
  DFFPOSX1 DFFPOSX1_401 ( .CLK(clk_i_bF_buf66), .D(u0_u5_tms_14__FF_INPUT), .Q(u0_tms5_14_) );
  DFFPOSX1 DFFPOSX1_402 ( .CLK(clk_i_bF_buf65), .D(u0_u5_tms_15__FF_INPUT), .Q(u0_tms5_15_) );
  DFFPOSX1 DFFPOSX1_403 ( .CLK(clk_i_bF_buf64), .D(u0_u5_tms_16__FF_INPUT), .Q(u0_tms5_16_) );
  DFFPOSX1 DFFPOSX1_404 ( .CLK(clk_i_bF_buf63), .D(u0_u5_tms_17__FF_INPUT), .Q(u0_tms5_17_) );
  DFFPOSX1 DFFPOSX1_405 ( .CLK(clk_i_bF_buf62), .D(u0_u5_tms_18__FF_INPUT), .Q(u0_tms5_18_) );
  DFFPOSX1 DFFPOSX1_406 ( .CLK(clk_i_bF_buf61), .D(u0_u5_tms_19__FF_INPUT), .Q(u0_tms5_19_) );
  DFFPOSX1 DFFPOSX1_407 ( .CLK(clk_i_bF_buf60), .D(u0_u5_tms_20__FF_INPUT), .Q(u0_tms5_20_) );
  DFFPOSX1 DFFPOSX1_408 ( .CLK(clk_i_bF_buf59), .D(u0_u5_tms_21__FF_INPUT), .Q(u0_tms5_21_) );
  DFFPOSX1 DFFPOSX1_409 ( .CLK(clk_i_bF_buf58), .D(u0_u5_tms_22__FF_INPUT), .Q(u0_tms5_22_) );
  DFFPOSX1 DFFPOSX1_41 ( .CLK(clk_i_bF_buf85), .D(\wb_addr_i[6] ), .Q(u0_wb_addr_r_6_) );
  DFFPOSX1 DFFPOSX1_410 ( .CLK(clk_i_bF_buf57), .D(u0_u5_tms_23__FF_INPUT), .Q(u0_tms5_23_) );
  DFFPOSX1 DFFPOSX1_411 ( .CLK(clk_i_bF_buf56), .D(u0_u5_tms_24__FF_INPUT), .Q(u0_tms5_24_) );
  DFFPOSX1 DFFPOSX1_412 ( .CLK(clk_i_bF_buf55), .D(u0_u5_tms_25__FF_INPUT), .Q(u0_tms5_25_) );
  DFFPOSX1 DFFPOSX1_413 ( .CLK(clk_i_bF_buf54), .D(u0_u5_tms_26__FF_INPUT), .Q(u0_tms5_26_) );
  DFFPOSX1 DFFPOSX1_414 ( .CLK(clk_i_bF_buf53), .D(u0_u5_tms_27__FF_INPUT), .Q(u0_tms5_27_) );
  DFFPOSX1 DFFPOSX1_415 ( .CLK(clk_i_bF_buf52), .D(u0_u5_tms_28__FF_INPUT), .Q(u0_tms5_28_) );
  DFFPOSX1 DFFPOSX1_416 ( .CLK(clk_i_bF_buf51), .D(u0_u5_tms_29__FF_INPUT), .Q(u0_tms5_29_) );
  DFFPOSX1 DFFPOSX1_417 ( .CLK(clk_i_bF_buf50), .D(u0_u5_tms_30__FF_INPUT), .Q(u0_tms5_30_) );
  DFFPOSX1 DFFPOSX1_418 ( .CLK(clk_i_bF_buf49), .D(u0_u5_tms_31__FF_INPUT), .Q(u0_tms5_31_) );
  DFFPOSX1 DFFPOSX1_419 ( .CLK(clk_i_bF_buf48), .D(u0_u5_csc_0__FF_INPUT), .Q(u0_csc5_0_) );
  DFFPOSX1 DFFPOSX1_42 ( .CLK(clk_i_bF_buf82), .D(u0_u0_tms_0__FF_INPUT), .Q(u0_tms0_0_) );
  DFFPOSX1 DFFPOSX1_420 ( .CLK(clk_i_bF_buf47), .D(u0_u5_csc_1__FF_INPUT), .Q(u0_csc5_1_) );
  DFFPOSX1 DFFPOSX1_421 ( .CLK(clk_i_bF_buf46), .D(u0_u5_csc_2__FF_INPUT), .Q(u0_csc5_2_) );
  DFFPOSX1 DFFPOSX1_422 ( .CLK(clk_i_bF_buf45), .D(u0_u5_csc_3__FF_INPUT), .Q(u0_csc5_3_) );
  DFFPOSX1 DFFPOSX1_423 ( .CLK(clk_i_bF_buf44), .D(u0_u5_csc_4__FF_INPUT), .Q(u0_csc5_4_) );
  DFFPOSX1 DFFPOSX1_424 ( .CLK(clk_i_bF_buf43), .D(u0_u5_csc_5__FF_INPUT), .Q(u0_csc5_5_) );
  DFFPOSX1 DFFPOSX1_425 ( .CLK(clk_i_bF_buf42), .D(u0_u5_csc_6__FF_INPUT), .Q(u0_csc5_6_) );
  DFFPOSX1 DFFPOSX1_426 ( .CLK(clk_i_bF_buf41), .D(u0_u5_csc_7__FF_INPUT), .Q(u0_csc5_7_) );
  DFFPOSX1 DFFPOSX1_427 ( .CLK(clk_i_bF_buf40), .D(u0_u5_csc_8__FF_INPUT), .Q(u0_csc5_8_) );
  DFFPOSX1 DFFPOSX1_428 ( .CLK(clk_i_bF_buf39), .D(u0_u5_csc_9__FF_INPUT), .Q(u0_csc5_9_) );
  DFFPOSX1 DFFPOSX1_429 ( .CLK(clk_i_bF_buf38), .D(u0_u5_csc_10__FF_INPUT), .Q(u0_csc5_10_) );
  DFFPOSX1 DFFPOSX1_43 ( .CLK(clk_i_bF_buf81), .D(u0_u0_tms_1__FF_INPUT), .Q(u0_tms0_1_) );
  DFFPOSX1 DFFPOSX1_430 ( .CLK(clk_i_bF_buf37), .D(u0_u5_csc_11__FF_INPUT), .Q(u0_csc5_11_) );
  DFFPOSX1 DFFPOSX1_431 ( .CLK(clk_i_bF_buf36), .D(u0_u5_csc_12__FF_INPUT), .Q(u0_csc5_12_) );
  DFFPOSX1 DFFPOSX1_432 ( .CLK(clk_i_bF_buf35), .D(u0_u5_csc_13__FF_INPUT), .Q(u0_csc5_13_) );
  DFFPOSX1 DFFPOSX1_433 ( .CLK(clk_i_bF_buf34), .D(u0_u5_csc_14__FF_INPUT), .Q(u0_csc5_14_) );
  DFFPOSX1 DFFPOSX1_434 ( .CLK(clk_i_bF_buf33), .D(u0_u5_csc_15__FF_INPUT), .Q(u0_csc5_15_) );
  DFFPOSX1 DFFPOSX1_435 ( .CLK(clk_i_bF_buf32), .D(u0_u5_csc_16__FF_INPUT), .Q(u0_csc5_16_) );
  DFFPOSX1 DFFPOSX1_436 ( .CLK(clk_i_bF_buf31), .D(u0_u5_csc_17__FF_INPUT), .Q(u0_csc5_17_) );
  DFFPOSX1 DFFPOSX1_437 ( .CLK(clk_i_bF_buf30), .D(u0_u5_csc_18__FF_INPUT), .Q(u0_csc5_18_) );
  DFFPOSX1 DFFPOSX1_438 ( .CLK(clk_i_bF_buf29), .D(u0_u5_csc_19__FF_INPUT), .Q(u0_csc5_19_) );
  DFFPOSX1 DFFPOSX1_439 ( .CLK(clk_i_bF_buf28), .D(u0_u5_csc_20__FF_INPUT), .Q(u0_csc5_20_) );
  DFFPOSX1 DFFPOSX1_44 ( .CLK(clk_i_bF_buf80), .D(u0_u0_tms_2__FF_INPUT), .Q(u0_tms0_2_) );
  DFFPOSX1 DFFPOSX1_440 ( .CLK(clk_i_bF_buf27), .D(u0_u5_csc_21__FF_INPUT), .Q(u0_csc5_21_) );
  DFFPOSX1 DFFPOSX1_441 ( .CLK(clk_i_bF_buf26), .D(u0_u5_csc_22__FF_INPUT), .Q(u0_csc5_22_) );
  DFFPOSX1 DFFPOSX1_442 ( .CLK(clk_i_bF_buf25), .D(u0_u5_csc_23__FF_INPUT), .Q(u0_csc5_23_) );
  DFFPOSX1 DFFPOSX1_443 ( .CLK(clk_i_bF_buf24), .D(u0_u5_csc_24__FF_INPUT), .Q(u0_csc5_24_) );
  DFFPOSX1 DFFPOSX1_444 ( .CLK(clk_i_bF_buf23), .D(u0_u5_csc_25__FF_INPUT), .Q(u0_csc5_25_) );
  DFFPOSX1 DFFPOSX1_445 ( .CLK(clk_i_bF_buf22), .D(u0_u5_csc_26__FF_INPUT), .Q(u0_csc5_26_) );
  DFFPOSX1 DFFPOSX1_446 ( .CLK(clk_i_bF_buf21), .D(u0_u5_csc_27__FF_INPUT), .Q(u0_csc5_27_) );
  DFFPOSX1 DFFPOSX1_447 ( .CLK(clk_i_bF_buf20), .D(u0_u5_csc_28__FF_INPUT), .Q(u0_csc5_28_) );
  DFFPOSX1 DFFPOSX1_448 ( .CLK(clk_i_bF_buf19), .D(u0_u5_csc_29__FF_INPUT), .Q(u0_csc5_29_) );
  DFFPOSX1 DFFPOSX1_449 ( .CLK(clk_i_bF_buf18), .D(u0_u5_csc_30__FF_INPUT), .Q(u0_csc5_30_) );
  DFFPOSX1 DFFPOSX1_45 ( .CLK(clk_i_bF_buf79), .D(u0_u0_tms_3__FF_INPUT), .Q(u0_tms0_3_) );
  DFFPOSX1 DFFPOSX1_450 ( .CLK(clk_i_bF_buf17), .D(u0_u5_csc_31__FF_INPUT), .Q(u0_csc5_31_) );
  DFFPOSX1 DFFPOSX1_451 ( .CLK(clk_i_bF_buf16), .D(\wb_addr_i[2] ), .Q(u0_u5_addr_r_2_) );
  DFFPOSX1 DFFPOSX1_452 ( .CLK(clk_i_bF_buf15), .D(\wb_addr_i[3] ), .Q(u0_u5_addr_r_3_) );
  DFFPOSX1 DFFPOSX1_453 ( .CLK(clk_i_bF_buf14), .D(\wb_addr_i[4] ), .Q(u0_u5_addr_r_4_) );
  DFFPOSX1 DFFPOSX1_454 ( .CLK(clk_i_bF_buf13), .D(\wb_addr_i[5] ), .Q(u0_u5_addr_r_5_) );
  DFFPOSX1 DFFPOSX1_455 ( .CLK(clk_i_bF_buf12), .D(\wb_addr_i[6] ), .Q(u0_u5_addr_r_6_) );
  DFFPOSX1 DFFPOSX1_456 ( .CLK(clk_i_bF_buf4), .D(u1_bank_adr_0__FF_INPUT), .Q(bank_adr_0_) );
  DFFPOSX1 DFFPOSX1_457 ( .CLK(clk_i_bF_buf3), .D(u1_bank_adr_1__FF_INPUT), .Q(bank_adr_1_) );
  DFFPOSX1 DFFPOSX1_458 ( .CLK(clk_i_bF_buf2), .D(u1_row_adr_0__FF_INPUT), .Q(row_adr_0_) );
  DFFPOSX1 DFFPOSX1_459 ( .CLK(clk_i_bF_buf1), .D(u1_row_adr_1__FF_INPUT), .Q(row_adr_1_) );
  DFFPOSX1 DFFPOSX1_46 ( .CLK(clk_i_bF_buf78), .D(u0_u0_tms_4__FF_INPUT), .Q(u0_tms0_4_) );
  DFFPOSX1 DFFPOSX1_460 ( .CLK(clk_i_bF_buf0), .D(u1_row_adr_2__FF_INPUT), .Q(row_adr_2_) );
  DFFPOSX1 DFFPOSX1_461 ( .CLK(clk_i_bF_buf125), .D(u1_row_adr_3__FF_INPUT), .Q(row_adr_3_) );
  DFFPOSX1 DFFPOSX1_462 ( .CLK(clk_i_bF_buf124), .D(u1_row_adr_4__FF_INPUT), .Q(row_adr_4_) );
  DFFPOSX1 DFFPOSX1_463 ( .CLK(clk_i_bF_buf123), .D(u1_row_adr_5__FF_INPUT), .Q(row_adr_5_) );
  DFFPOSX1 DFFPOSX1_464 ( .CLK(clk_i_bF_buf122), .D(u1_row_adr_6__FF_INPUT), .Q(row_adr_6_) );
  DFFPOSX1 DFFPOSX1_465 ( .CLK(clk_i_bF_buf121), .D(u1_row_adr_7__FF_INPUT), .Q(row_adr_7_) );
  DFFPOSX1 DFFPOSX1_466 ( .CLK(clk_i_bF_buf120), .D(u1_row_adr_8__FF_INPUT), .Q(row_adr_8_) );
  DFFPOSX1 DFFPOSX1_467 ( .CLK(clk_i_bF_buf119), .D(u1_row_adr_9__FF_INPUT), .Q(row_adr_9_) );
  DFFPOSX1 DFFPOSX1_468 ( .CLK(clk_i_bF_buf118), .D(u1_row_adr_10__FF_INPUT), .Q(row_adr_10_) );
  DFFPOSX1 DFFPOSX1_469 ( .CLK(clk_i_bF_buf117), .D(u1_row_adr_11__FF_INPUT), .Q(row_adr_11_) );
  DFFPOSX1 DFFPOSX1_47 ( .CLK(clk_i_bF_buf77), .D(u0_u0_tms_5__FF_INPUT), .Q(u0_tms0_5_) );
  DFFPOSX1 DFFPOSX1_470 ( .CLK(clk_i_bF_buf116), .D(u1_row_adr_12__FF_INPUT), .Q(row_adr_12_) );
  DFFPOSX1 DFFPOSX1_471 ( .CLK(clk_i_bF_buf115), .D(u1_col_adr_0__FF_INPUT), .Q(u1_col_adr_0_) );
  DFFPOSX1 DFFPOSX1_472 ( .CLK(clk_i_bF_buf114), .D(u1_col_adr_1__FF_INPUT), .Q(u1_col_adr_1_) );
  DFFPOSX1 DFFPOSX1_473 ( .CLK(clk_i_bF_buf113), .D(u1_col_adr_2__FF_INPUT), .Q(u1_col_adr_2_) );
  DFFPOSX1 DFFPOSX1_474 ( .CLK(clk_i_bF_buf112), .D(u1_col_adr_3__FF_INPUT), .Q(u1_col_adr_3_) );
  DFFPOSX1 DFFPOSX1_475 ( .CLK(clk_i_bF_buf111), .D(u1_col_adr_4__FF_INPUT), .Q(u1_col_adr_4_) );
  DFFPOSX1 DFFPOSX1_476 ( .CLK(clk_i_bF_buf110), .D(u1_col_adr_5__FF_INPUT), .Q(u1_col_adr_5_) );
  DFFPOSX1 DFFPOSX1_477 ( .CLK(clk_i_bF_buf109), .D(u1_col_adr_6__FF_INPUT), .Q(u1_col_adr_6_) );
  DFFPOSX1 DFFPOSX1_478 ( .CLK(clk_i_bF_buf108), .D(u1_col_adr_7__FF_INPUT), .Q(u1_col_adr_7_) );
  DFFPOSX1 DFFPOSX1_479 ( .CLK(clk_i_bF_buf107), .D(u1_col_adr_8__FF_INPUT), .Q(u1_col_adr_8_) );
  DFFPOSX1 DFFPOSX1_48 ( .CLK(clk_i_bF_buf76), .D(u0_u0_tms_6__FF_INPUT), .Q(u0_tms0_6_) );
  DFFPOSX1 DFFPOSX1_480 ( .CLK(clk_i_bF_buf106), .D(u1_col_adr_9__FF_INPUT), .Q(u1_col_adr_9_) );
  DFFPOSX1 DFFPOSX1_481 ( .CLK(clk_i_bF_buf105), .D(u1_acs_addr_0__FF_INPUT), .Q(u1_acs_addr_0_) );
  DFFPOSX1 DFFPOSX1_482 ( .CLK(clk_i_bF_buf104), .D(u1_acs_addr_1__FF_INPUT), .Q(u1_acs_addr_1_) );
  DFFPOSX1 DFFPOSX1_483 ( .CLK(clk_i_bF_buf103), .D(u1_acs_addr_2__FF_INPUT), .Q(u1_acs_addr_2_) );
  DFFPOSX1 DFFPOSX1_484 ( .CLK(clk_i_bF_buf102), .D(u1_acs_addr_3__FF_INPUT), .Q(u1_acs_addr_3_) );
  DFFPOSX1 DFFPOSX1_485 ( .CLK(clk_i_bF_buf101), .D(u1_acs_addr_4__FF_INPUT), .Q(u1_acs_addr_4_) );
  DFFPOSX1 DFFPOSX1_486 ( .CLK(clk_i_bF_buf100), .D(u1_acs_addr_5__FF_INPUT), .Q(u1_acs_addr_5_) );
  DFFPOSX1 DFFPOSX1_487 ( .CLK(clk_i_bF_buf99), .D(u1_acs_addr_6__FF_INPUT), .Q(u1_acs_addr_6_) );
  DFFPOSX1 DFFPOSX1_488 ( .CLK(clk_i_bF_buf98), .D(u1_acs_addr_7__FF_INPUT), .Q(u1_acs_addr_7_) );
  DFFPOSX1 DFFPOSX1_489 ( .CLK(clk_i_bF_buf97), .D(u1_acs_addr_8__FF_INPUT), .Q(u1_acs_addr_8_) );
  DFFPOSX1 DFFPOSX1_49 ( .CLK(clk_i_bF_buf75), .D(u0_u0_tms_7__FF_INPUT), .Q(u0_tms0_7_) );
  DFFPOSX1 DFFPOSX1_490 ( .CLK(clk_i_bF_buf96), .D(u1_acs_addr_9__FF_INPUT), .Q(u1_acs_addr_9_) );
  DFFPOSX1 DFFPOSX1_491 ( .CLK(clk_i_bF_buf95), .D(u1_acs_addr_10__FF_INPUT), .Q(u1_acs_addr_10_) );
  DFFPOSX1 DFFPOSX1_492 ( .CLK(clk_i_bF_buf94), .D(u1_acs_addr_11__FF_INPUT), .Q(u1_acs_addr_11_) );
  DFFPOSX1 DFFPOSX1_493 ( .CLK(clk_i_bF_buf93), .D(u1_acs_addr_12__FF_INPUT), .Q(u1_acs_addr_12_) );
  DFFPOSX1 DFFPOSX1_494 ( .CLK(clk_i_bF_buf92), .D(u1_acs_addr_13__FF_INPUT), .Q(u1_acs_addr_13_) );
  DFFPOSX1 DFFPOSX1_495 ( .CLK(clk_i_bF_buf91), .D(u1_acs_addr_14__FF_INPUT), .Q(u1_acs_addr_14_) );
  DFFPOSX1 DFFPOSX1_496 ( .CLK(clk_i_bF_buf90), .D(u1_acs_addr_15__FF_INPUT), .Q(u1_acs_addr_15_) );
  DFFPOSX1 DFFPOSX1_497 ( .CLK(clk_i_bF_buf89), .D(u1_acs_addr_16__FF_INPUT), .Q(u1_acs_addr_16_) );
  DFFPOSX1 DFFPOSX1_498 ( .CLK(clk_i_bF_buf88), .D(u1_acs_addr_17__FF_INPUT), .Q(u1_acs_addr_17_) );
  DFFPOSX1 DFFPOSX1_499 ( .CLK(clk_i_bF_buf87), .D(u1_acs_addr_18__FF_INPUT), .Q(u1_acs_addr_18_) );
  DFFPOSX1 DFFPOSX1_5 ( .CLK(clk_i_bF_buf121), .D(u0_poc_1__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56321_1_) );
  DFFPOSX1 DFFPOSX1_50 ( .CLK(clk_i_bF_buf74), .D(u0_u0_tms_8__FF_INPUT), .Q(u0_tms0_8_) );
  DFFPOSX1 DFFPOSX1_500 ( .CLK(clk_i_bF_buf86), .D(u1_acs_addr_19__FF_INPUT), .Q(u1_acs_addr_19_) );
  DFFPOSX1 DFFPOSX1_501 ( .CLK(clk_i_bF_buf85), .D(u1_acs_addr_20__FF_INPUT), .Q(u1_acs_addr_20_) );
  DFFPOSX1 DFFPOSX1_502 ( .CLK(clk_i_bF_buf84), .D(u1_acs_addr_21__FF_INPUT), .Q(u1_acs_addr_21_) );
  DFFPOSX1 DFFPOSX1_503 ( .CLK(clk_i_bF_buf83), .D(u1_acs_addr_22__FF_INPUT), .Q(u1_acs_addr_22_) );
  DFFPOSX1 DFFPOSX1_504 ( .CLK(clk_i_bF_buf82), .D(u1_acs_addr_23__FF_INPUT), .Q(u1_acs_addr_23_) );
  DFFPOSX1 DFFPOSX1_505 ( .CLK(clk_i_bF_buf81), .D(u1_sram_addr_0__FF_INPUT), .Q(u1_sram_addr_0_) );
  DFFPOSX1 DFFPOSX1_506 ( .CLK(clk_i_bF_buf80), .D(u1_sram_addr_1__FF_INPUT), .Q(u1_sram_addr_1_) );
  DFFPOSX1 DFFPOSX1_507 ( .CLK(clk_i_bF_buf79), .D(u1_sram_addr_2__FF_INPUT), .Q(u1_sram_addr_2_) );
  DFFPOSX1 DFFPOSX1_508 ( .CLK(clk_i_bF_buf78), .D(u1_sram_addr_3__FF_INPUT), .Q(u1_sram_addr_3_) );
  DFFPOSX1 DFFPOSX1_509 ( .CLK(clk_i_bF_buf77), .D(u1_sram_addr_4__FF_INPUT), .Q(u1_sram_addr_4_) );
  DFFPOSX1 DFFPOSX1_51 ( .CLK(clk_i_bF_buf73), .D(u0_u0_tms_9__FF_INPUT), .Q(u0_tms0_9_) );
  DFFPOSX1 DFFPOSX1_510 ( .CLK(clk_i_bF_buf76), .D(u1_sram_addr_5__FF_INPUT), .Q(u1_sram_addr_5_) );
  DFFPOSX1 DFFPOSX1_511 ( .CLK(clk_i_bF_buf75), .D(u1_sram_addr_6__FF_INPUT), .Q(u1_sram_addr_6_) );
  DFFPOSX1 DFFPOSX1_512 ( .CLK(clk_i_bF_buf74), .D(u1_sram_addr_7__FF_INPUT), .Q(u1_sram_addr_7_) );
  DFFPOSX1 DFFPOSX1_513 ( .CLK(clk_i_bF_buf73), .D(u1_sram_addr_8__FF_INPUT), .Q(u1_sram_addr_8_) );
  DFFPOSX1 DFFPOSX1_514 ( .CLK(clk_i_bF_buf72), .D(u1_sram_addr_9__FF_INPUT), .Q(u1_sram_addr_9_) );
  DFFPOSX1 DFFPOSX1_515 ( .CLK(clk_i_bF_buf71), .D(u1_sram_addr_10__FF_INPUT), .Q(u1_sram_addr_10_) );
  DFFPOSX1 DFFPOSX1_516 ( .CLK(clk_i_bF_buf70), .D(u1_sram_addr_11__FF_INPUT), .Q(u1_sram_addr_11_) );
  DFFPOSX1 DFFPOSX1_517 ( .CLK(clk_i_bF_buf69), .D(u1_sram_addr_12__FF_INPUT), .Q(u1_sram_addr_12_) );
  DFFPOSX1 DFFPOSX1_518 ( .CLK(clk_i_bF_buf68), .D(u1_sram_addr_13__FF_INPUT), .Q(u1_sram_addr_13_) );
  DFFPOSX1 DFFPOSX1_519 ( .CLK(clk_i_bF_buf67), .D(u1_sram_addr_14__FF_INPUT), .Q(u1_sram_addr_14_) );
  DFFPOSX1 DFFPOSX1_52 ( .CLK(clk_i_bF_buf72), .D(u0_u0_tms_10__FF_INPUT), .Q(u0_tms0_10_) );
  DFFPOSX1 DFFPOSX1_520 ( .CLK(clk_i_bF_buf66), .D(u1_sram_addr_15__FF_INPUT), .Q(u1_sram_addr_15_) );
  DFFPOSX1 DFFPOSX1_521 ( .CLK(clk_i_bF_buf65), .D(u1_sram_addr_16__FF_INPUT), .Q(u1_sram_addr_16_) );
  DFFPOSX1 DFFPOSX1_522 ( .CLK(clk_i_bF_buf64), .D(u1_sram_addr_17__FF_INPUT), .Q(u1_sram_addr_17_) );
  DFFPOSX1 DFFPOSX1_523 ( .CLK(clk_i_bF_buf63), .D(u1_sram_addr_18__FF_INPUT), .Q(u1_sram_addr_18_) );
  DFFPOSX1 DFFPOSX1_524 ( .CLK(clk_i_bF_buf62), .D(u1_sram_addr_19__FF_INPUT), .Q(u1_sram_addr_19_) );
  DFFPOSX1 DFFPOSX1_525 ( .CLK(clk_i_bF_buf61), .D(u1_sram_addr_20__FF_INPUT), .Q(u1_sram_addr_20_) );
  DFFPOSX1 DFFPOSX1_526 ( .CLK(clk_i_bF_buf60), .D(u1_sram_addr_21__FF_INPUT), .Q(u1_sram_addr_21_) );
  DFFPOSX1 DFFPOSX1_527 ( .CLK(clk_i_bF_buf59), .D(u1_sram_addr_22__FF_INPUT), .Q(u1_sram_addr_22_) );
  DFFPOSX1 DFFPOSX1_528 ( .CLK(clk_i_bF_buf58), .D(u1_sram_addr_23__FF_INPUT), .Q(u1_sram_addr_23_) );
  DFFPOSX1 DFFPOSX1_529 ( .CLK(clk_i_bF_buf57), .D(u1_u0_out_r_0__FF_INPUT), .Q(u1_acs_addr_pl1_0_) );
  DFFPOSX1 DFFPOSX1_53 ( .CLK(clk_i_bF_buf71), .D(u0_u0_tms_11__FF_INPUT), .Q(u0_tms0_11_) );
  DFFPOSX1 DFFPOSX1_530 ( .CLK(clk_i_bF_buf56), .D(u1_u0_out_r_1__FF_INPUT), .Q(u1_acs_addr_pl1_1_) );
  DFFPOSX1 DFFPOSX1_531 ( .CLK(clk_i_bF_buf55), .D(u1_u0_out_r_2__FF_INPUT), .Q(u1_acs_addr_pl1_2_) );
  DFFPOSX1 DFFPOSX1_532 ( .CLK(clk_i_bF_buf54), .D(u1_u0_out_r_3__FF_INPUT), .Q(u1_acs_addr_pl1_3_) );
  DFFPOSX1 DFFPOSX1_533 ( .CLK(clk_i_bF_buf53), .D(u1_u0_out_r_4__FF_INPUT), .Q(u1_acs_addr_pl1_4_) );
  DFFPOSX1 DFFPOSX1_534 ( .CLK(clk_i_bF_buf52), .D(u1_u0_out_r_5__FF_INPUT), .Q(u1_acs_addr_pl1_5_) );
  DFFPOSX1 DFFPOSX1_535 ( .CLK(clk_i_bF_buf51), .D(u1_u0_out_r_6__FF_INPUT), .Q(u1_acs_addr_pl1_6_) );
  DFFPOSX1 DFFPOSX1_536 ( .CLK(clk_i_bF_buf50), .D(u1_u0_out_r_7__FF_INPUT), .Q(u1_acs_addr_pl1_7_) );
  DFFPOSX1 DFFPOSX1_537 ( .CLK(clk_i_bF_buf49), .D(u1_u0_out_r_8__FF_INPUT), .Q(u1_acs_addr_pl1_8_) );
  DFFPOSX1 DFFPOSX1_538 ( .CLK(clk_i_bF_buf48), .D(u1_u0_out_r_9__FF_INPUT), .Q(u1_acs_addr_pl1_9_) );
  DFFPOSX1 DFFPOSX1_539 ( .CLK(clk_i_bF_buf47), .D(u1_u0_out_r_10__FF_INPUT), .Q(u1_acs_addr_pl1_10_) );
  DFFPOSX1 DFFPOSX1_54 ( .CLK(clk_i_bF_buf70), .D(u0_u0_tms_12__FF_INPUT), .Q(u0_tms0_12_) );
  DFFPOSX1 DFFPOSX1_540 ( .CLK(clk_i_bF_buf46), .D(u1_u0_out_r_11__FF_INPUT), .Q(u1_acs_addr_pl1_11_) );
  DFFPOSX1 DFFPOSX1_541 ( .CLK(clk_i_bF_buf45), .D(u1_u0_out_r_12__FF_INPUT), .Q(u1_u0_inc_next) );
  DFFPOSX1 DFFPOSX1_542 ( .CLK(clk_i_bF_buf44), .D(u2_row_same_FF_INPUT), .Q(row_same) );
  DFFPOSX1 DFFPOSX1_543 ( .CLK(clk_i_bF_buf43), .D(u2_bank_open_FF_INPUT), .Q(bank_open) );
  DFFPOSX1 DFFPOSX1_544 ( .CLK(clk_i_bF_buf42), .D(u2_u0_b3_last_row_0__FF_INPUT), .Q(u2_u0_b3_last_row_0_) );
  DFFPOSX1 DFFPOSX1_545 ( .CLK(clk_i_bF_buf41), .D(u2_u0_b3_last_row_1__FF_INPUT), .Q(u2_u0_b3_last_row_1_) );
  DFFPOSX1 DFFPOSX1_546 ( .CLK(clk_i_bF_buf40), .D(u2_u0_b3_last_row_2__FF_INPUT), .Q(u2_u0_b3_last_row_2_) );
  DFFPOSX1 DFFPOSX1_547 ( .CLK(clk_i_bF_buf39), .D(u2_u0_b3_last_row_3__FF_INPUT), .Q(u2_u0_b3_last_row_3_) );
  DFFPOSX1 DFFPOSX1_548 ( .CLK(clk_i_bF_buf38), .D(u2_u0_b3_last_row_4__FF_INPUT), .Q(u2_u0_b3_last_row_4_) );
  DFFPOSX1 DFFPOSX1_549 ( .CLK(clk_i_bF_buf37), .D(u2_u0_b3_last_row_5__FF_INPUT), .Q(u2_u0_b3_last_row_5_) );
  DFFPOSX1 DFFPOSX1_55 ( .CLK(clk_i_bF_buf69), .D(u0_u0_tms_13__FF_INPUT), .Q(u0_tms0_13_) );
  DFFPOSX1 DFFPOSX1_550 ( .CLK(clk_i_bF_buf36), .D(u2_u0_b3_last_row_6__FF_INPUT), .Q(u2_u0_b3_last_row_6_) );
  DFFPOSX1 DFFPOSX1_551 ( .CLK(clk_i_bF_buf35), .D(u2_u0_b3_last_row_7__FF_INPUT), .Q(u2_u0_b3_last_row_7_) );
  DFFPOSX1 DFFPOSX1_552 ( .CLK(clk_i_bF_buf34), .D(u2_u0_b3_last_row_8__FF_INPUT), .Q(u2_u0_b3_last_row_8_) );
  DFFPOSX1 DFFPOSX1_553 ( .CLK(clk_i_bF_buf33), .D(u2_u0_b3_last_row_9__FF_INPUT), .Q(u2_u0_b3_last_row_9_) );
  DFFPOSX1 DFFPOSX1_554 ( .CLK(clk_i_bF_buf32), .D(u2_u0_b3_last_row_10__FF_INPUT), .Q(u2_u0_b3_last_row_10_) );
  DFFPOSX1 DFFPOSX1_555 ( .CLK(clk_i_bF_buf31), .D(u2_u0_b3_last_row_11__FF_INPUT), .Q(u2_u0_b3_last_row_11_) );
  DFFPOSX1 DFFPOSX1_556 ( .CLK(clk_i_bF_buf30), .D(u2_u0_b3_last_row_12__FF_INPUT), .Q(u2_u0_b3_last_row_12_) );
  DFFPOSX1 DFFPOSX1_557 ( .CLK(clk_i_bF_buf29), .D(u2_u0_b2_last_row_0__FF_INPUT), .Q(u2_u0_b2_last_row_0_) );
  DFFPOSX1 DFFPOSX1_558 ( .CLK(clk_i_bF_buf28), .D(u2_u0_b2_last_row_1__FF_INPUT), .Q(u2_u0_b2_last_row_1_) );
  DFFPOSX1 DFFPOSX1_559 ( .CLK(clk_i_bF_buf27), .D(u2_u0_b2_last_row_2__FF_INPUT), .Q(u2_u0_b2_last_row_2_) );
  DFFPOSX1 DFFPOSX1_56 ( .CLK(clk_i_bF_buf68), .D(u0_u0_tms_14__FF_INPUT), .Q(u0_tms0_14_) );
  DFFPOSX1 DFFPOSX1_560 ( .CLK(clk_i_bF_buf26), .D(u2_u0_b2_last_row_3__FF_INPUT), .Q(u2_u0_b2_last_row_3_) );
  DFFPOSX1 DFFPOSX1_561 ( .CLK(clk_i_bF_buf25), .D(u2_u0_b2_last_row_4__FF_INPUT), .Q(u2_u0_b2_last_row_4_) );
  DFFPOSX1 DFFPOSX1_562 ( .CLK(clk_i_bF_buf24), .D(u2_u0_b2_last_row_5__FF_INPUT), .Q(u2_u0_b2_last_row_5_) );
  DFFPOSX1 DFFPOSX1_563 ( .CLK(clk_i_bF_buf23), .D(u2_u0_b2_last_row_6__FF_INPUT), .Q(u2_u0_b2_last_row_6_) );
  DFFPOSX1 DFFPOSX1_564 ( .CLK(clk_i_bF_buf22), .D(u2_u0_b2_last_row_7__FF_INPUT), .Q(u2_u0_b2_last_row_7_) );
  DFFPOSX1 DFFPOSX1_565 ( .CLK(clk_i_bF_buf21), .D(u2_u0_b2_last_row_8__FF_INPUT), .Q(u2_u0_b2_last_row_8_) );
  DFFPOSX1 DFFPOSX1_566 ( .CLK(clk_i_bF_buf20), .D(u2_u0_b2_last_row_9__FF_INPUT), .Q(u2_u0_b2_last_row_9_) );
  DFFPOSX1 DFFPOSX1_567 ( .CLK(clk_i_bF_buf19), .D(u2_u0_b2_last_row_10__FF_INPUT), .Q(u2_u0_b2_last_row_10_) );
  DFFPOSX1 DFFPOSX1_568 ( .CLK(clk_i_bF_buf18), .D(u2_u0_b2_last_row_11__FF_INPUT), .Q(u2_u0_b2_last_row_11_) );
  DFFPOSX1 DFFPOSX1_569 ( .CLK(clk_i_bF_buf17), .D(u2_u0_b2_last_row_12__FF_INPUT), .Q(u2_u0_b2_last_row_12_) );
  DFFPOSX1 DFFPOSX1_57 ( .CLK(clk_i_bF_buf67), .D(u0_u0_tms_15__FF_INPUT), .Q(u0_tms0_15_) );
  DFFPOSX1 DFFPOSX1_570 ( .CLK(clk_i_bF_buf16), .D(u2_u0_b1_last_row_0__FF_INPUT), .Q(u2_u0_b1_last_row_0_) );
  DFFPOSX1 DFFPOSX1_571 ( .CLK(clk_i_bF_buf15), .D(u2_u0_b1_last_row_1__FF_INPUT), .Q(u2_u0_b1_last_row_1_) );
  DFFPOSX1 DFFPOSX1_572 ( .CLK(clk_i_bF_buf14), .D(u2_u0_b1_last_row_2__FF_INPUT), .Q(u2_u0_b1_last_row_2_) );
  DFFPOSX1 DFFPOSX1_573 ( .CLK(clk_i_bF_buf13), .D(u2_u0_b1_last_row_3__FF_INPUT), .Q(u2_u0_b1_last_row_3_) );
  DFFPOSX1 DFFPOSX1_574 ( .CLK(clk_i_bF_buf12), .D(u2_u0_b1_last_row_4__FF_INPUT), .Q(u2_u0_b1_last_row_4_) );
  DFFPOSX1 DFFPOSX1_575 ( .CLK(clk_i_bF_buf11), .D(u2_u0_b1_last_row_5__FF_INPUT), .Q(u2_u0_b1_last_row_5_) );
  DFFPOSX1 DFFPOSX1_576 ( .CLK(clk_i_bF_buf10), .D(u2_u0_b1_last_row_6__FF_INPUT), .Q(u2_u0_b1_last_row_6_) );
  DFFPOSX1 DFFPOSX1_577 ( .CLK(clk_i_bF_buf9), .D(u2_u0_b1_last_row_7__FF_INPUT), .Q(u2_u0_b1_last_row_7_) );
  DFFPOSX1 DFFPOSX1_578 ( .CLK(clk_i_bF_buf8), .D(u2_u0_b1_last_row_8__FF_INPUT), .Q(u2_u0_b1_last_row_8_) );
  DFFPOSX1 DFFPOSX1_579 ( .CLK(clk_i_bF_buf7), .D(u2_u0_b1_last_row_9__FF_INPUT), .Q(u2_u0_b1_last_row_9_) );
  DFFPOSX1 DFFPOSX1_58 ( .CLK(clk_i_bF_buf66), .D(u0_u0_tms_16__FF_INPUT), .Q(u0_tms0_16_) );
  DFFPOSX1 DFFPOSX1_580 ( .CLK(clk_i_bF_buf6), .D(u2_u0_b1_last_row_10__FF_INPUT), .Q(u2_u0_b1_last_row_10_) );
  DFFPOSX1 DFFPOSX1_581 ( .CLK(clk_i_bF_buf5), .D(u2_u0_b1_last_row_11__FF_INPUT), .Q(u2_u0_b1_last_row_11_) );
  DFFPOSX1 DFFPOSX1_582 ( .CLK(clk_i_bF_buf4), .D(u2_u0_b1_last_row_12__FF_INPUT), .Q(u2_u0_b1_last_row_12_) );
  DFFPOSX1 DFFPOSX1_583 ( .CLK(clk_i_bF_buf3), .D(u2_u0_b0_last_row_0__FF_INPUT), .Q(u2_u0_b0_last_row_0_) );
  DFFPOSX1 DFFPOSX1_584 ( .CLK(clk_i_bF_buf2), .D(u2_u0_b0_last_row_1__FF_INPUT), .Q(u2_u0_b0_last_row_1_) );
  DFFPOSX1 DFFPOSX1_585 ( .CLK(clk_i_bF_buf1), .D(u2_u0_b0_last_row_2__FF_INPUT), .Q(u2_u0_b0_last_row_2_) );
  DFFPOSX1 DFFPOSX1_586 ( .CLK(clk_i_bF_buf0), .D(u2_u0_b0_last_row_3__FF_INPUT), .Q(u2_u0_b0_last_row_3_) );
  DFFPOSX1 DFFPOSX1_587 ( .CLK(clk_i_bF_buf125), .D(u2_u0_b0_last_row_4__FF_INPUT), .Q(u2_u0_b0_last_row_4_) );
  DFFPOSX1 DFFPOSX1_588 ( .CLK(clk_i_bF_buf124), .D(u2_u0_b0_last_row_5__FF_INPUT), .Q(u2_u0_b0_last_row_5_) );
  DFFPOSX1 DFFPOSX1_589 ( .CLK(clk_i_bF_buf123), .D(u2_u0_b0_last_row_6__FF_INPUT), .Q(u2_u0_b0_last_row_6_) );
  DFFPOSX1 DFFPOSX1_59 ( .CLK(clk_i_bF_buf65), .D(u0_u0_tms_17__FF_INPUT), .Q(u0_tms0_17_) );
  DFFPOSX1 DFFPOSX1_590 ( .CLK(clk_i_bF_buf122), .D(u2_u0_b0_last_row_7__FF_INPUT), .Q(u2_u0_b0_last_row_7_) );
  DFFPOSX1 DFFPOSX1_591 ( .CLK(clk_i_bF_buf121), .D(u2_u0_b0_last_row_8__FF_INPUT), .Q(u2_u0_b0_last_row_8_) );
  DFFPOSX1 DFFPOSX1_592 ( .CLK(clk_i_bF_buf120), .D(u2_u0_b0_last_row_9__FF_INPUT), .Q(u2_u0_b0_last_row_9_) );
  DFFPOSX1 DFFPOSX1_593 ( .CLK(clk_i_bF_buf119), .D(u2_u0_b0_last_row_10__FF_INPUT), .Q(u2_u0_b0_last_row_10_) );
  DFFPOSX1 DFFPOSX1_594 ( .CLK(clk_i_bF_buf118), .D(u2_u0_b0_last_row_11__FF_INPUT), .Q(u2_u0_b0_last_row_11_) );
  DFFPOSX1 DFFPOSX1_595 ( .CLK(clk_i_bF_buf117), .D(u2_u0_b0_last_row_12__FF_INPUT), .Q(u2_u0_b0_last_row_12_) );
  DFFPOSX1 DFFPOSX1_596 ( .CLK(clk_i_bF_buf112), .D(u2_u1_b3_last_row_0__FF_INPUT), .Q(u2_u1_b3_last_row_0_) );
  DFFPOSX1 DFFPOSX1_597 ( .CLK(clk_i_bF_buf111), .D(u2_u1_b3_last_row_1__FF_INPUT), .Q(u2_u1_b3_last_row_1_) );
  DFFPOSX1 DFFPOSX1_598 ( .CLK(clk_i_bF_buf110), .D(u2_u1_b3_last_row_2__FF_INPUT), .Q(u2_u1_b3_last_row_2_) );
  DFFPOSX1 DFFPOSX1_599 ( .CLK(clk_i_bF_buf109), .D(u2_u1_b3_last_row_3__FF_INPUT), .Q(u2_u1_b3_last_row_3_) );
  DFFPOSX1 DFFPOSX1_6 ( .CLK(clk_i_bF_buf120), .D(u0_poc_2__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56321_2_) );
  DFFPOSX1 DFFPOSX1_60 ( .CLK(clk_i_bF_buf64), .D(u0_u0_tms_18__FF_INPUT), .Q(u0_tms0_18_) );
  DFFPOSX1 DFFPOSX1_600 ( .CLK(clk_i_bF_buf108), .D(u2_u1_b3_last_row_4__FF_INPUT), .Q(u2_u1_b3_last_row_4_) );
  DFFPOSX1 DFFPOSX1_601 ( .CLK(clk_i_bF_buf107), .D(u2_u1_b3_last_row_5__FF_INPUT), .Q(u2_u1_b3_last_row_5_) );
  DFFPOSX1 DFFPOSX1_602 ( .CLK(clk_i_bF_buf106), .D(u2_u1_b3_last_row_6__FF_INPUT), .Q(u2_u1_b3_last_row_6_) );
  DFFPOSX1 DFFPOSX1_603 ( .CLK(clk_i_bF_buf105), .D(u2_u1_b3_last_row_7__FF_INPUT), .Q(u2_u1_b3_last_row_7_) );
  DFFPOSX1 DFFPOSX1_604 ( .CLK(clk_i_bF_buf104), .D(u2_u1_b3_last_row_8__FF_INPUT), .Q(u2_u1_b3_last_row_8_) );
  DFFPOSX1 DFFPOSX1_605 ( .CLK(clk_i_bF_buf103), .D(u2_u1_b3_last_row_9__FF_INPUT), .Q(u2_u1_b3_last_row_9_) );
  DFFPOSX1 DFFPOSX1_606 ( .CLK(clk_i_bF_buf102), .D(u2_u1_b3_last_row_10__FF_INPUT), .Q(u2_u1_b3_last_row_10_) );
  DFFPOSX1 DFFPOSX1_607 ( .CLK(clk_i_bF_buf101), .D(u2_u1_b3_last_row_11__FF_INPUT), .Q(u2_u1_b3_last_row_11_) );
  DFFPOSX1 DFFPOSX1_608 ( .CLK(clk_i_bF_buf100), .D(u2_u1_b3_last_row_12__FF_INPUT), .Q(u2_u1_b3_last_row_12_) );
  DFFPOSX1 DFFPOSX1_609 ( .CLK(clk_i_bF_buf99), .D(u2_u1_b2_last_row_0__FF_INPUT), .Q(u2_u1_b2_last_row_0_) );
  DFFPOSX1 DFFPOSX1_61 ( .CLK(clk_i_bF_buf63), .D(u0_u0_tms_19__FF_INPUT), .Q(u0_tms0_19_) );
  DFFPOSX1 DFFPOSX1_610 ( .CLK(clk_i_bF_buf98), .D(u2_u1_b2_last_row_1__FF_INPUT), .Q(u2_u1_b2_last_row_1_) );
  DFFPOSX1 DFFPOSX1_611 ( .CLK(clk_i_bF_buf97), .D(u2_u1_b2_last_row_2__FF_INPUT), .Q(u2_u1_b2_last_row_2_) );
  DFFPOSX1 DFFPOSX1_612 ( .CLK(clk_i_bF_buf96), .D(u2_u1_b2_last_row_3__FF_INPUT), .Q(u2_u1_b2_last_row_3_) );
  DFFPOSX1 DFFPOSX1_613 ( .CLK(clk_i_bF_buf95), .D(u2_u1_b2_last_row_4__FF_INPUT), .Q(u2_u1_b2_last_row_4_) );
  DFFPOSX1 DFFPOSX1_614 ( .CLK(clk_i_bF_buf94), .D(u2_u1_b2_last_row_5__FF_INPUT), .Q(u2_u1_b2_last_row_5_) );
  DFFPOSX1 DFFPOSX1_615 ( .CLK(clk_i_bF_buf93), .D(u2_u1_b2_last_row_6__FF_INPUT), .Q(u2_u1_b2_last_row_6_) );
  DFFPOSX1 DFFPOSX1_616 ( .CLK(clk_i_bF_buf92), .D(u2_u1_b2_last_row_7__FF_INPUT), .Q(u2_u1_b2_last_row_7_) );
  DFFPOSX1 DFFPOSX1_617 ( .CLK(clk_i_bF_buf91), .D(u2_u1_b2_last_row_8__FF_INPUT), .Q(u2_u1_b2_last_row_8_) );
  DFFPOSX1 DFFPOSX1_618 ( .CLK(clk_i_bF_buf90), .D(u2_u1_b2_last_row_9__FF_INPUT), .Q(u2_u1_b2_last_row_9_) );
  DFFPOSX1 DFFPOSX1_619 ( .CLK(clk_i_bF_buf89), .D(u2_u1_b2_last_row_10__FF_INPUT), .Q(u2_u1_b2_last_row_10_) );
  DFFPOSX1 DFFPOSX1_62 ( .CLK(clk_i_bF_buf62), .D(u0_u0_tms_20__FF_INPUT), .Q(u0_tms0_20_) );
  DFFPOSX1 DFFPOSX1_620 ( .CLK(clk_i_bF_buf88), .D(u2_u1_b2_last_row_11__FF_INPUT), .Q(u2_u1_b2_last_row_11_) );
  DFFPOSX1 DFFPOSX1_621 ( .CLK(clk_i_bF_buf87), .D(u2_u1_b2_last_row_12__FF_INPUT), .Q(u2_u1_b2_last_row_12_) );
  DFFPOSX1 DFFPOSX1_622 ( .CLK(clk_i_bF_buf86), .D(u2_u1_b1_last_row_0__FF_INPUT), .Q(u2_u1_b1_last_row_0_) );
  DFFPOSX1 DFFPOSX1_623 ( .CLK(clk_i_bF_buf85), .D(u2_u1_b1_last_row_1__FF_INPUT), .Q(u2_u1_b1_last_row_1_) );
  DFFPOSX1 DFFPOSX1_624 ( .CLK(clk_i_bF_buf84), .D(u2_u1_b1_last_row_2__FF_INPUT), .Q(u2_u1_b1_last_row_2_) );
  DFFPOSX1 DFFPOSX1_625 ( .CLK(clk_i_bF_buf83), .D(u2_u1_b1_last_row_3__FF_INPUT), .Q(u2_u1_b1_last_row_3_) );
  DFFPOSX1 DFFPOSX1_626 ( .CLK(clk_i_bF_buf82), .D(u2_u1_b1_last_row_4__FF_INPUT), .Q(u2_u1_b1_last_row_4_) );
  DFFPOSX1 DFFPOSX1_627 ( .CLK(clk_i_bF_buf81), .D(u2_u1_b1_last_row_5__FF_INPUT), .Q(u2_u1_b1_last_row_5_) );
  DFFPOSX1 DFFPOSX1_628 ( .CLK(clk_i_bF_buf80), .D(u2_u1_b1_last_row_6__FF_INPUT), .Q(u2_u1_b1_last_row_6_) );
  DFFPOSX1 DFFPOSX1_629 ( .CLK(clk_i_bF_buf79), .D(u2_u1_b1_last_row_7__FF_INPUT), .Q(u2_u1_b1_last_row_7_) );
  DFFPOSX1 DFFPOSX1_63 ( .CLK(clk_i_bF_buf61), .D(u0_u0_tms_21__FF_INPUT), .Q(u0_tms0_21_) );
  DFFPOSX1 DFFPOSX1_630 ( .CLK(clk_i_bF_buf78), .D(u2_u1_b1_last_row_8__FF_INPUT), .Q(u2_u1_b1_last_row_8_) );
  DFFPOSX1 DFFPOSX1_631 ( .CLK(clk_i_bF_buf77), .D(u2_u1_b1_last_row_9__FF_INPUT), .Q(u2_u1_b1_last_row_9_) );
  DFFPOSX1 DFFPOSX1_632 ( .CLK(clk_i_bF_buf76), .D(u2_u1_b1_last_row_10__FF_INPUT), .Q(u2_u1_b1_last_row_10_) );
  DFFPOSX1 DFFPOSX1_633 ( .CLK(clk_i_bF_buf75), .D(u2_u1_b1_last_row_11__FF_INPUT), .Q(u2_u1_b1_last_row_11_) );
  DFFPOSX1 DFFPOSX1_634 ( .CLK(clk_i_bF_buf74), .D(u2_u1_b1_last_row_12__FF_INPUT), .Q(u2_u1_b1_last_row_12_) );
  DFFPOSX1 DFFPOSX1_635 ( .CLK(clk_i_bF_buf73), .D(u2_u1_b0_last_row_0__FF_INPUT), .Q(u2_u1_b0_last_row_0_) );
  DFFPOSX1 DFFPOSX1_636 ( .CLK(clk_i_bF_buf72), .D(u2_u1_b0_last_row_1__FF_INPUT), .Q(u2_u1_b0_last_row_1_) );
  DFFPOSX1 DFFPOSX1_637 ( .CLK(clk_i_bF_buf71), .D(u2_u1_b0_last_row_2__FF_INPUT), .Q(u2_u1_b0_last_row_2_) );
  DFFPOSX1 DFFPOSX1_638 ( .CLK(clk_i_bF_buf70), .D(u2_u1_b0_last_row_3__FF_INPUT), .Q(u2_u1_b0_last_row_3_) );
  DFFPOSX1 DFFPOSX1_639 ( .CLK(clk_i_bF_buf69), .D(u2_u1_b0_last_row_4__FF_INPUT), .Q(u2_u1_b0_last_row_4_) );
  DFFPOSX1 DFFPOSX1_64 ( .CLK(clk_i_bF_buf60), .D(u0_u0_tms_22__FF_INPUT), .Q(u0_tms0_22_) );
  DFFPOSX1 DFFPOSX1_640 ( .CLK(clk_i_bF_buf68), .D(u2_u1_b0_last_row_5__FF_INPUT), .Q(u2_u1_b0_last_row_5_) );
  DFFPOSX1 DFFPOSX1_641 ( .CLK(clk_i_bF_buf67), .D(u2_u1_b0_last_row_6__FF_INPUT), .Q(u2_u1_b0_last_row_6_) );
  DFFPOSX1 DFFPOSX1_642 ( .CLK(clk_i_bF_buf66), .D(u2_u1_b0_last_row_7__FF_INPUT), .Q(u2_u1_b0_last_row_7_) );
  DFFPOSX1 DFFPOSX1_643 ( .CLK(clk_i_bF_buf65), .D(u2_u1_b0_last_row_8__FF_INPUT), .Q(u2_u1_b0_last_row_8_) );
  DFFPOSX1 DFFPOSX1_644 ( .CLK(clk_i_bF_buf64), .D(u2_u1_b0_last_row_9__FF_INPUT), .Q(u2_u1_b0_last_row_9_) );
  DFFPOSX1 DFFPOSX1_645 ( .CLK(clk_i_bF_buf63), .D(u2_u1_b0_last_row_10__FF_INPUT), .Q(u2_u1_b0_last_row_10_) );
  DFFPOSX1 DFFPOSX1_646 ( .CLK(clk_i_bF_buf62), .D(u2_u1_b0_last_row_11__FF_INPUT), .Q(u2_u1_b0_last_row_11_) );
  DFFPOSX1 DFFPOSX1_647 ( .CLK(clk_i_bF_buf61), .D(u2_u1_b0_last_row_12__FF_INPUT), .Q(u2_u1_b0_last_row_12_) );
  DFFPOSX1 DFFPOSX1_648 ( .CLK(clk_i_bF_buf56), .D(u2_u2_b3_last_row_0__FF_INPUT), .Q(u2_u2_b3_last_row_0_) );
  DFFPOSX1 DFFPOSX1_649 ( .CLK(clk_i_bF_buf55), .D(u2_u2_b3_last_row_1__FF_INPUT), .Q(u2_u2_b3_last_row_1_) );
  DFFPOSX1 DFFPOSX1_65 ( .CLK(clk_i_bF_buf59), .D(u0_u0_tms_23__FF_INPUT), .Q(u0_tms0_23_) );
  DFFPOSX1 DFFPOSX1_650 ( .CLK(clk_i_bF_buf54), .D(u2_u2_b3_last_row_2__FF_INPUT), .Q(u2_u2_b3_last_row_2_) );
  DFFPOSX1 DFFPOSX1_651 ( .CLK(clk_i_bF_buf53), .D(u2_u2_b3_last_row_3__FF_INPUT), .Q(u2_u2_b3_last_row_3_) );
  DFFPOSX1 DFFPOSX1_652 ( .CLK(clk_i_bF_buf52), .D(u2_u2_b3_last_row_4__FF_INPUT), .Q(u2_u2_b3_last_row_4_) );
  DFFPOSX1 DFFPOSX1_653 ( .CLK(clk_i_bF_buf51), .D(u2_u2_b3_last_row_5__FF_INPUT), .Q(u2_u2_b3_last_row_5_) );
  DFFPOSX1 DFFPOSX1_654 ( .CLK(clk_i_bF_buf50), .D(u2_u2_b3_last_row_6__FF_INPUT), .Q(u2_u2_b3_last_row_6_) );
  DFFPOSX1 DFFPOSX1_655 ( .CLK(clk_i_bF_buf49), .D(u2_u2_b3_last_row_7__FF_INPUT), .Q(u2_u2_b3_last_row_7_) );
  DFFPOSX1 DFFPOSX1_656 ( .CLK(clk_i_bF_buf48), .D(u2_u2_b3_last_row_8__FF_INPUT), .Q(u2_u2_b3_last_row_8_) );
  DFFPOSX1 DFFPOSX1_657 ( .CLK(clk_i_bF_buf47), .D(u2_u2_b3_last_row_9__FF_INPUT), .Q(u2_u2_b3_last_row_9_) );
  DFFPOSX1 DFFPOSX1_658 ( .CLK(clk_i_bF_buf46), .D(u2_u2_b3_last_row_10__FF_INPUT), .Q(u2_u2_b3_last_row_10_) );
  DFFPOSX1 DFFPOSX1_659 ( .CLK(clk_i_bF_buf45), .D(u2_u2_b3_last_row_11__FF_INPUT), .Q(u2_u2_b3_last_row_11_) );
  DFFPOSX1 DFFPOSX1_66 ( .CLK(clk_i_bF_buf58), .D(u0_u0_tms_24__FF_INPUT), .Q(u0_tms0_24_) );
  DFFPOSX1 DFFPOSX1_660 ( .CLK(clk_i_bF_buf44), .D(u2_u2_b3_last_row_12__FF_INPUT), .Q(u2_u2_b3_last_row_12_) );
  DFFPOSX1 DFFPOSX1_661 ( .CLK(clk_i_bF_buf43), .D(u2_u2_b2_last_row_0__FF_INPUT), .Q(u2_u2_b2_last_row_0_) );
  DFFPOSX1 DFFPOSX1_662 ( .CLK(clk_i_bF_buf42), .D(u2_u2_b2_last_row_1__FF_INPUT), .Q(u2_u2_b2_last_row_1_) );
  DFFPOSX1 DFFPOSX1_663 ( .CLK(clk_i_bF_buf41), .D(u2_u2_b2_last_row_2__FF_INPUT), .Q(u2_u2_b2_last_row_2_) );
  DFFPOSX1 DFFPOSX1_664 ( .CLK(clk_i_bF_buf40), .D(u2_u2_b2_last_row_3__FF_INPUT), .Q(u2_u2_b2_last_row_3_) );
  DFFPOSX1 DFFPOSX1_665 ( .CLK(clk_i_bF_buf39), .D(u2_u2_b2_last_row_4__FF_INPUT), .Q(u2_u2_b2_last_row_4_) );
  DFFPOSX1 DFFPOSX1_666 ( .CLK(clk_i_bF_buf38), .D(u2_u2_b2_last_row_5__FF_INPUT), .Q(u2_u2_b2_last_row_5_) );
  DFFPOSX1 DFFPOSX1_667 ( .CLK(clk_i_bF_buf37), .D(u2_u2_b2_last_row_6__FF_INPUT), .Q(u2_u2_b2_last_row_6_) );
  DFFPOSX1 DFFPOSX1_668 ( .CLK(clk_i_bF_buf36), .D(u2_u2_b2_last_row_7__FF_INPUT), .Q(u2_u2_b2_last_row_7_) );
  DFFPOSX1 DFFPOSX1_669 ( .CLK(clk_i_bF_buf35), .D(u2_u2_b2_last_row_8__FF_INPUT), .Q(u2_u2_b2_last_row_8_) );
  DFFPOSX1 DFFPOSX1_67 ( .CLK(clk_i_bF_buf57), .D(u0_u0_tms_25__FF_INPUT), .Q(u0_tms0_25_) );
  DFFPOSX1 DFFPOSX1_670 ( .CLK(clk_i_bF_buf34), .D(u2_u2_b2_last_row_9__FF_INPUT), .Q(u2_u2_b2_last_row_9_) );
  DFFPOSX1 DFFPOSX1_671 ( .CLK(clk_i_bF_buf33), .D(u2_u2_b2_last_row_10__FF_INPUT), .Q(u2_u2_b2_last_row_10_) );
  DFFPOSX1 DFFPOSX1_672 ( .CLK(clk_i_bF_buf32), .D(u2_u2_b2_last_row_11__FF_INPUT), .Q(u2_u2_b2_last_row_11_) );
  DFFPOSX1 DFFPOSX1_673 ( .CLK(clk_i_bF_buf31), .D(u2_u2_b2_last_row_12__FF_INPUT), .Q(u2_u2_b2_last_row_12_) );
  DFFPOSX1 DFFPOSX1_674 ( .CLK(clk_i_bF_buf30), .D(u2_u2_b1_last_row_0__FF_INPUT), .Q(u2_u2_b1_last_row_0_) );
  DFFPOSX1 DFFPOSX1_675 ( .CLK(clk_i_bF_buf29), .D(u2_u2_b1_last_row_1__FF_INPUT), .Q(u2_u2_b1_last_row_1_) );
  DFFPOSX1 DFFPOSX1_676 ( .CLK(clk_i_bF_buf28), .D(u2_u2_b1_last_row_2__FF_INPUT), .Q(u2_u2_b1_last_row_2_) );
  DFFPOSX1 DFFPOSX1_677 ( .CLK(clk_i_bF_buf27), .D(u2_u2_b1_last_row_3__FF_INPUT), .Q(u2_u2_b1_last_row_3_) );
  DFFPOSX1 DFFPOSX1_678 ( .CLK(clk_i_bF_buf26), .D(u2_u2_b1_last_row_4__FF_INPUT), .Q(u2_u2_b1_last_row_4_) );
  DFFPOSX1 DFFPOSX1_679 ( .CLK(clk_i_bF_buf25), .D(u2_u2_b1_last_row_5__FF_INPUT), .Q(u2_u2_b1_last_row_5_) );
  DFFPOSX1 DFFPOSX1_68 ( .CLK(clk_i_bF_buf56), .D(u0_u0_tms_26__FF_INPUT), .Q(u0_tms0_26_) );
  DFFPOSX1 DFFPOSX1_680 ( .CLK(clk_i_bF_buf24), .D(u2_u2_b1_last_row_6__FF_INPUT), .Q(u2_u2_b1_last_row_6_) );
  DFFPOSX1 DFFPOSX1_681 ( .CLK(clk_i_bF_buf23), .D(u2_u2_b1_last_row_7__FF_INPUT), .Q(u2_u2_b1_last_row_7_) );
  DFFPOSX1 DFFPOSX1_682 ( .CLK(clk_i_bF_buf22), .D(u2_u2_b1_last_row_8__FF_INPUT), .Q(u2_u2_b1_last_row_8_) );
  DFFPOSX1 DFFPOSX1_683 ( .CLK(clk_i_bF_buf21), .D(u2_u2_b1_last_row_9__FF_INPUT), .Q(u2_u2_b1_last_row_9_) );
  DFFPOSX1 DFFPOSX1_684 ( .CLK(clk_i_bF_buf20), .D(u2_u2_b1_last_row_10__FF_INPUT), .Q(u2_u2_b1_last_row_10_) );
  DFFPOSX1 DFFPOSX1_685 ( .CLK(clk_i_bF_buf19), .D(u2_u2_b1_last_row_11__FF_INPUT), .Q(u2_u2_b1_last_row_11_) );
  DFFPOSX1 DFFPOSX1_686 ( .CLK(clk_i_bF_buf18), .D(u2_u2_b1_last_row_12__FF_INPUT), .Q(u2_u2_b1_last_row_12_) );
  DFFPOSX1 DFFPOSX1_687 ( .CLK(clk_i_bF_buf17), .D(u2_u2_b0_last_row_0__FF_INPUT), .Q(u2_u2_b0_last_row_0_) );
  DFFPOSX1 DFFPOSX1_688 ( .CLK(clk_i_bF_buf16), .D(u2_u2_b0_last_row_1__FF_INPUT), .Q(u2_u2_b0_last_row_1_) );
  DFFPOSX1 DFFPOSX1_689 ( .CLK(clk_i_bF_buf15), .D(u2_u2_b0_last_row_2__FF_INPUT), .Q(u2_u2_b0_last_row_2_) );
  DFFPOSX1 DFFPOSX1_69 ( .CLK(clk_i_bF_buf55), .D(u0_u0_tms_27__FF_INPUT), .Q(u0_tms0_27_) );
  DFFPOSX1 DFFPOSX1_690 ( .CLK(clk_i_bF_buf14), .D(u2_u2_b0_last_row_3__FF_INPUT), .Q(u2_u2_b0_last_row_3_) );
  DFFPOSX1 DFFPOSX1_691 ( .CLK(clk_i_bF_buf13), .D(u2_u2_b0_last_row_4__FF_INPUT), .Q(u2_u2_b0_last_row_4_) );
  DFFPOSX1 DFFPOSX1_692 ( .CLK(clk_i_bF_buf12), .D(u2_u2_b0_last_row_5__FF_INPUT), .Q(u2_u2_b0_last_row_5_) );
  DFFPOSX1 DFFPOSX1_693 ( .CLK(clk_i_bF_buf11), .D(u2_u2_b0_last_row_6__FF_INPUT), .Q(u2_u2_b0_last_row_6_) );
  DFFPOSX1 DFFPOSX1_694 ( .CLK(clk_i_bF_buf10), .D(u2_u2_b0_last_row_7__FF_INPUT), .Q(u2_u2_b0_last_row_7_) );
  DFFPOSX1 DFFPOSX1_695 ( .CLK(clk_i_bF_buf9), .D(u2_u2_b0_last_row_8__FF_INPUT), .Q(u2_u2_b0_last_row_8_) );
  DFFPOSX1 DFFPOSX1_696 ( .CLK(clk_i_bF_buf8), .D(u2_u2_b0_last_row_9__FF_INPUT), .Q(u2_u2_b0_last_row_9_) );
  DFFPOSX1 DFFPOSX1_697 ( .CLK(clk_i_bF_buf7), .D(u2_u2_b0_last_row_10__FF_INPUT), .Q(u2_u2_b0_last_row_10_) );
  DFFPOSX1 DFFPOSX1_698 ( .CLK(clk_i_bF_buf6), .D(u2_u2_b0_last_row_11__FF_INPUT), .Q(u2_u2_b0_last_row_11_) );
  DFFPOSX1 DFFPOSX1_699 ( .CLK(clk_i_bF_buf5), .D(u2_u2_b0_last_row_12__FF_INPUT), .Q(u2_u2_b0_last_row_12_) );
  DFFPOSX1 DFFPOSX1_7 ( .CLK(clk_i_bF_buf119), .D(u0_poc_3__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56321_3_) );
  DFFPOSX1 DFFPOSX1_70 ( .CLK(clk_i_bF_buf54), .D(u0_u0_tms_28__FF_INPUT), .Q(u0_tms0_28_) );
  DFFPOSX1 DFFPOSX1_700 ( .CLK(clk_i_bF_buf0), .D(u2_u3_b3_last_row_0__FF_INPUT), .Q(u2_u3_b3_last_row_0_) );
  DFFPOSX1 DFFPOSX1_701 ( .CLK(clk_i_bF_buf125), .D(u2_u3_b3_last_row_1__FF_INPUT), .Q(u2_u3_b3_last_row_1_) );
  DFFPOSX1 DFFPOSX1_702 ( .CLK(clk_i_bF_buf124), .D(u2_u3_b3_last_row_2__FF_INPUT), .Q(u2_u3_b3_last_row_2_) );
  DFFPOSX1 DFFPOSX1_703 ( .CLK(clk_i_bF_buf123), .D(u2_u3_b3_last_row_3__FF_INPUT), .Q(u2_u3_b3_last_row_3_) );
  DFFPOSX1 DFFPOSX1_704 ( .CLK(clk_i_bF_buf122), .D(u2_u3_b3_last_row_4__FF_INPUT), .Q(u2_u3_b3_last_row_4_) );
  DFFPOSX1 DFFPOSX1_705 ( .CLK(clk_i_bF_buf121), .D(u2_u3_b3_last_row_5__FF_INPUT), .Q(u2_u3_b3_last_row_5_) );
  DFFPOSX1 DFFPOSX1_706 ( .CLK(clk_i_bF_buf120), .D(u2_u3_b3_last_row_6__FF_INPUT), .Q(u2_u3_b3_last_row_6_) );
  DFFPOSX1 DFFPOSX1_707 ( .CLK(clk_i_bF_buf119), .D(u2_u3_b3_last_row_7__FF_INPUT), .Q(u2_u3_b3_last_row_7_) );
  DFFPOSX1 DFFPOSX1_708 ( .CLK(clk_i_bF_buf118), .D(u2_u3_b3_last_row_8__FF_INPUT), .Q(u2_u3_b3_last_row_8_) );
  DFFPOSX1 DFFPOSX1_709 ( .CLK(clk_i_bF_buf117), .D(u2_u3_b3_last_row_9__FF_INPUT), .Q(u2_u3_b3_last_row_9_) );
  DFFPOSX1 DFFPOSX1_71 ( .CLK(clk_i_bF_buf53), .D(u0_u0_tms_29__FF_INPUT), .Q(u0_tms0_29_) );
  DFFPOSX1 DFFPOSX1_710 ( .CLK(clk_i_bF_buf116), .D(u2_u3_b3_last_row_10__FF_INPUT), .Q(u2_u3_b3_last_row_10_) );
  DFFPOSX1 DFFPOSX1_711 ( .CLK(clk_i_bF_buf115), .D(u2_u3_b3_last_row_11__FF_INPUT), .Q(u2_u3_b3_last_row_11_) );
  DFFPOSX1 DFFPOSX1_712 ( .CLK(clk_i_bF_buf114), .D(u2_u3_b3_last_row_12__FF_INPUT), .Q(u2_u3_b3_last_row_12_) );
  DFFPOSX1 DFFPOSX1_713 ( .CLK(clk_i_bF_buf113), .D(u2_u3_b2_last_row_0__FF_INPUT), .Q(u2_u3_b2_last_row_0_) );
  DFFPOSX1 DFFPOSX1_714 ( .CLK(clk_i_bF_buf112), .D(u2_u3_b2_last_row_1__FF_INPUT), .Q(u2_u3_b2_last_row_1_) );
  DFFPOSX1 DFFPOSX1_715 ( .CLK(clk_i_bF_buf111), .D(u2_u3_b2_last_row_2__FF_INPUT), .Q(u2_u3_b2_last_row_2_) );
  DFFPOSX1 DFFPOSX1_716 ( .CLK(clk_i_bF_buf110), .D(u2_u3_b2_last_row_3__FF_INPUT), .Q(u2_u3_b2_last_row_3_) );
  DFFPOSX1 DFFPOSX1_717 ( .CLK(clk_i_bF_buf109), .D(u2_u3_b2_last_row_4__FF_INPUT), .Q(u2_u3_b2_last_row_4_) );
  DFFPOSX1 DFFPOSX1_718 ( .CLK(clk_i_bF_buf108), .D(u2_u3_b2_last_row_5__FF_INPUT), .Q(u2_u3_b2_last_row_5_) );
  DFFPOSX1 DFFPOSX1_719 ( .CLK(clk_i_bF_buf107), .D(u2_u3_b2_last_row_6__FF_INPUT), .Q(u2_u3_b2_last_row_6_) );
  DFFPOSX1 DFFPOSX1_72 ( .CLK(clk_i_bF_buf52), .D(u0_u0_tms_30__FF_INPUT), .Q(u0_tms0_30_) );
  DFFPOSX1 DFFPOSX1_720 ( .CLK(clk_i_bF_buf106), .D(u2_u3_b2_last_row_7__FF_INPUT), .Q(u2_u3_b2_last_row_7_) );
  DFFPOSX1 DFFPOSX1_721 ( .CLK(clk_i_bF_buf105), .D(u2_u3_b2_last_row_8__FF_INPUT), .Q(u2_u3_b2_last_row_8_) );
  DFFPOSX1 DFFPOSX1_722 ( .CLK(clk_i_bF_buf104), .D(u2_u3_b2_last_row_9__FF_INPUT), .Q(u2_u3_b2_last_row_9_) );
  DFFPOSX1 DFFPOSX1_723 ( .CLK(clk_i_bF_buf103), .D(u2_u3_b2_last_row_10__FF_INPUT), .Q(u2_u3_b2_last_row_10_) );
  DFFPOSX1 DFFPOSX1_724 ( .CLK(clk_i_bF_buf102), .D(u2_u3_b2_last_row_11__FF_INPUT), .Q(u2_u3_b2_last_row_11_) );
  DFFPOSX1 DFFPOSX1_725 ( .CLK(clk_i_bF_buf101), .D(u2_u3_b2_last_row_12__FF_INPUT), .Q(u2_u3_b2_last_row_12_) );
  DFFPOSX1 DFFPOSX1_726 ( .CLK(clk_i_bF_buf100), .D(u2_u3_b1_last_row_0__FF_INPUT), .Q(u2_u3_b1_last_row_0_) );
  DFFPOSX1 DFFPOSX1_727 ( .CLK(clk_i_bF_buf99), .D(u2_u3_b1_last_row_1__FF_INPUT), .Q(u2_u3_b1_last_row_1_) );
  DFFPOSX1 DFFPOSX1_728 ( .CLK(clk_i_bF_buf98), .D(u2_u3_b1_last_row_2__FF_INPUT), .Q(u2_u3_b1_last_row_2_) );
  DFFPOSX1 DFFPOSX1_729 ( .CLK(clk_i_bF_buf97), .D(u2_u3_b1_last_row_3__FF_INPUT), .Q(u2_u3_b1_last_row_3_) );
  DFFPOSX1 DFFPOSX1_73 ( .CLK(clk_i_bF_buf51), .D(u0_u0_tms_31__FF_INPUT), .Q(u0_tms0_31_) );
  DFFPOSX1 DFFPOSX1_730 ( .CLK(clk_i_bF_buf96), .D(u2_u3_b1_last_row_4__FF_INPUT), .Q(u2_u3_b1_last_row_4_) );
  DFFPOSX1 DFFPOSX1_731 ( .CLK(clk_i_bF_buf95), .D(u2_u3_b1_last_row_5__FF_INPUT), .Q(u2_u3_b1_last_row_5_) );
  DFFPOSX1 DFFPOSX1_732 ( .CLK(clk_i_bF_buf94), .D(u2_u3_b1_last_row_6__FF_INPUT), .Q(u2_u3_b1_last_row_6_) );
  DFFPOSX1 DFFPOSX1_733 ( .CLK(clk_i_bF_buf93), .D(u2_u3_b1_last_row_7__FF_INPUT), .Q(u2_u3_b1_last_row_7_) );
  DFFPOSX1 DFFPOSX1_734 ( .CLK(clk_i_bF_buf92), .D(u2_u3_b1_last_row_8__FF_INPUT), .Q(u2_u3_b1_last_row_8_) );
  DFFPOSX1 DFFPOSX1_735 ( .CLK(clk_i_bF_buf91), .D(u2_u3_b1_last_row_9__FF_INPUT), .Q(u2_u3_b1_last_row_9_) );
  DFFPOSX1 DFFPOSX1_736 ( .CLK(clk_i_bF_buf90), .D(u2_u3_b1_last_row_10__FF_INPUT), .Q(u2_u3_b1_last_row_10_) );
  DFFPOSX1 DFFPOSX1_737 ( .CLK(clk_i_bF_buf89), .D(u2_u3_b1_last_row_11__FF_INPUT), .Q(u2_u3_b1_last_row_11_) );
  DFFPOSX1 DFFPOSX1_738 ( .CLK(clk_i_bF_buf88), .D(u2_u3_b1_last_row_12__FF_INPUT), .Q(u2_u3_b1_last_row_12_) );
  DFFPOSX1 DFFPOSX1_739 ( .CLK(clk_i_bF_buf87), .D(u2_u3_b0_last_row_0__FF_INPUT), .Q(u2_u3_b0_last_row_0_) );
  DFFPOSX1 DFFPOSX1_74 ( .CLK(clk_i_bF_buf50), .D(u0_u0_csc_0__FF_INPUT), .Q(u0_csc0_0_) );
  DFFPOSX1 DFFPOSX1_740 ( .CLK(clk_i_bF_buf86), .D(u2_u3_b0_last_row_1__FF_INPUT), .Q(u2_u3_b0_last_row_1_) );
  DFFPOSX1 DFFPOSX1_741 ( .CLK(clk_i_bF_buf85), .D(u2_u3_b0_last_row_2__FF_INPUT), .Q(u2_u3_b0_last_row_2_) );
  DFFPOSX1 DFFPOSX1_742 ( .CLK(clk_i_bF_buf84), .D(u2_u3_b0_last_row_3__FF_INPUT), .Q(u2_u3_b0_last_row_3_) );
  DFFPOSX1 DFFPOSX1_743 ( .CLK(clk_i_bF_buf83), .D(u2_u3_b0_last_row_4__FF_INPUT), .Q(u2_u3_b0_last_row_4_) );
  DFFPOSX1 DFFPOSX1_744 ( .CLK(clk_i_bF_buf82), .D(u2_u3_b0_last_row_5__FF_INPUT), .Q(u2_u3_b0_last_row_5_) );
  DFFPOSX1 DFFPOSX1_745 ( .CLK(clk_i_bF_buf81), .D(u2_u3_b0_last_row_6__FF_INPUT), .Q(u2_u3_b0_last_row_6_) );
  DFFPOSX1 DFFPOSX1_746 ( .CLK(clk_i_bF_buf80), .D(u2_u3_b0_last_row_7__FF_INPUT), .Q(u2_u3_b0_last_row_7_) );
  DFFPOSX1 DFFPOSX1_747 ( .CLK(clk_i_bF_buf79), .D(u2_u3_b0_last_row_8__FF_INPUT), .Q(u2_u3_b0_last_row_8_) );
  DFFPOSX1 DFFPOSX1_748 ( .CLK(clk_i_bF_buf78), .D(u2_u3_b0_last_row_9__FF_INPUT), .Q(u2_u3_b0_last_row_9_) );
  DFFPOSX1 DFFPOSX1_749 ( .CLK(clk_i_bF_buf77), .D(u2_u3_b0_last_row_10__FF_INPUT), .Q(u2_u3_b0_last_row_10_) );
  DFFPOSX1 DFFPOSX1_75 ( .CLK(clk_i_bF_buf49), .D(u0_u0_csc_1__FF_INPUT), .Q(u0_csc0_1_) );
  DFFPOSX1 DFFPOSX1_750 ( .CLK(clk_i_bF_buf76), .D(u2_u3_b0_last_row_11__FF_INPUT), .Q(u2_u3_b0_last_row_11_) );
  DFFPOSX1 DFFPOSX1_751 ( .CLK(clk_i_bF_buf75), .D(u2_u3_b0_last_row_12__FF_INPUT), .Q(u2_u3_b0_last_row_12_) );
  DFFPOSX1 DFFPOSX1_752 ( .CLK(clk_i_bF_buf70), .D(u2_u4_b3_last_row_0__FF_INPUT), .Q(u2_u4_b3_last_row_0_) );
  DFFPOSX1 DFFPOSX1_753 ( .CLK(clk_i_bF_buf69), .D(u2_u4_b3_last_row_1__FF_INPUT), .Q(u2_u4_b3_last_row_1_) );
  DFFPOSX1 DFFPOSX1_754 ( .CLK(clk_i_bF_buf68), .D(u2_u4_b3_last_row_2__FF_INPUT), .Q(u2_u4_b3_last_row_2_) );
  DFFPOSX1 DFFPOSX1_755 ( .CLK(clk_i_bF_buf67), .D(u2_u4_b3_last_row_3__FF_INPUT), .Q(u2_u4_b3_last_row_3_) );
  DFFPOSX1 DFFPOSX1_756 ( .CLK(clk_i_bF_buf66), .D(u2_u4_b3_last_row_4__FF_INPUT), .Q(u2_u4_b3_last_row_4_) );
  DFFPOSX1 DFFPOSX1_757 ( .CLK(clk_i_bF_buf65), .D(u2_u4_b3_last_row_5__FF_INPUT), .Q(u2_u4_b3_last_row_5_) );
  DFFPOSX1 DFFPOSX1_758 ( .CLK(clk_i_bF_buf64), .D(u2_u4_b3_last_row_6__FF_INPUT), .Q(u2_u4_b3_last_row_6_) );
  DFFPOSX1 DFFPOSX1_759 ( .CLK(clk_i_bF_buf63), .D(u2_u4_b3_last_row_7__FF_INPUT), .Q(u2_u4_b3_last_row_7_) );
  DFFPOSX1 DFFPOSX1_76 ( .CLK(clk_i_bF_buf48), .D(u0_u0_csc_2__FF_INPUT), .Q(u0_csc0_2_) );
  DFFPOSX1 DFFPOSX1_760 ( .CLK(clk_i_bF_buf62), .D(u2_u4_b3_last_row_8__FF_INPUT), .Q(u2_u4_b3_last_row_8_) );
  DFFPOSX1 DFFPOSX1_761 ( .CLK(clk_i_bF_buf61), .D(u2_u4_b3_last_row_9__FF_INPUT), .Q(u2_u4_b3_last_row_9_) );
  DFFPOSX1 DFFPOSX1_762 ( .CLK(clk_i_bF_buf60), .D(u2_u4_b3_last_row_10__FF_INPUT), .Q(u2_u4_b3_last_row_10_) );
  DFFPOSX1 DFFPOSX1_763 ( .CLK(clk_i_bF_buf59), .D(u2_u4_b3_last_row_11__FF_INPUT), .Q(u2_u4_b3_last_row_11_) );
  DFFPOSX1 DFFPOSX1_764 ( .CLK(clk_i_bF_buf58), .D(u2_u4_b3_last_row_12__FF_INPUT), .Q(u2_u4_b3_last_row_12_) );
  DFFPOSX1 DFFPOSX1_765 ( .CLK(clk_i_bF_buf57), .D(u2_u4_b2_last_row_0__FF_INPUT), .Q(u2_u4_b2_last_row_0_) );
  DFFPOSX1 DFFPOSX1_766 ( .CLK(clk_i_bF_buf56), .D(u2_u4_b2_last_row_1__FF_INPUT), .Q(u2_u4_b2_last_row_1_) );
  DFFPOSX1 DFFPOSX1_767 ( .CLK(clk_i_bF_buf55), .D(u2_u4_b2_last_row_2__FF_INPUT), .Q(u2_u4_b2_last_row_2_) );
  DFFPOSX1 DFFPOSX1_768 ( .CLK(clk_i_bF_buf54), .D(u2_u4_b2_last_row_3__FF_INPUT), .Q(u2_u4_b2_last_row_3_) );
  DFFPOSX1 DFFPOSX1_769 ( .CLK(clk_i_bF_buf53), .D(u2_u4_b2_last_row_4__FF_INPUT), .Q(u2_u4_b2_last_row_4_) );
  DFFPOSX1 DFFPOSX1_77 ( .CLK(clk_i_bF_buf47), .D(u0_u0_csc_3__FF_INPUT), .Q(u0_csc0_3_) );
  DFFPOSX1 DFFPOSX1_770 ( .CLK(clk_i_bF_buf52), .D(u2_u4_b2_last_row_5__FF_INPUT), .Q(u2_u4_b2_last_row_5_) );
  DFFPOSX1 DFFPOSX1_771 ( .CLK(clk_i_bF_buf51), .D(u2_u4_b2_last_row_6__FF_INPUT), .Q(u2_u4_b2_last_row_6_) );
  DFFPOSX1 DFFPOSX1_772 ( .CLK(clk_i_bF_buf50), .D(u2_u4_b2_last_row_7__FF_INPUT), .Q(u2_u4_b2_last_row_7_) );
  DFFPOSX1 DFFPOSX1_773 ( .CLK(clk_i_bF_buf49), .D(u2_u4_b2_last_row_8__FF_INPUT), .Q(u2_u4_b2_last_row_8_) );
  DFFPOSX1 DFFPOSX1_774 ( .CLK(clk_i_bF_buf48), .D(u2_u4_b2_last_row_9__FF_INPUT), .Q(u2_u4_b2_last_row_9_) );
  DFFPOSX1 DFFPOSX1_775 ( .CLK(clk_i_bF_buf47), .D(u2_u4_b2_last_row_10__FF_INPUT), .Q(u2_u4_b2_last_row_10_) );
  DFFPOSX1 DFFPOSX1_776 ( .CLK(clk_i_bF_buf46), .D(u2_u4_b2_last_row_11__FF_INPUT), .Q(u2_u4_b2_last_row_11_) );
  DFFPOSX1 DFFPOSX1_777 ( .CLK(clk_i_bF_buf45), .D(u2_u4_b2_last_row_12__FF_INPUT), .Q(u2_u4_b2_last_row_12_) );
  DFFPOSX1 DFFPOSX1_778 ( .CLK(clk_i_bF_buf44), .D(u2_u4_b1_last_row_0__FF_INPUT), .Q(u2_u4_b1_last_row_0_) );
  DFFPOSX1 DFFPOSX1_779 ( .CLK(clk_i_bF_buf43), .D(u2_u4_b1_last_row_1__FF_INPUT), .Q(u2_u4_b1_last_row_1_) );
  DFFPOSX1 DFFPOSX1_78 ( .CLK(clk_i_bF_buf46), .D(u0_u0_csc_4__FF_INPUT), .Q(u0_csc0_4_) );
  DFFPOSX1 DFFPOSX1_780 ( .CLK(clk_i_bF_buf42), .D(u2_u4_b1_last_row_2__FF_INPUT), .Q(u2_u4_b1_last_row_2_) );
  DFFPOSX1 DFFPOSX1_781 ( .CLK(clk_i_bF_buf41), .D(u2_u4_b1_last_row_3__FF_INPUT), .Q(u2_u4_b1_last_row_3_) );
  DFFPOSX1 DFFPOSX1_782 ( .CLK(clk_i_bF_buf40), .D(u2_u4_b1_last_row_4__FF_INPUT), .Q(u2_u4_b1_last_row_4_) );
  DFFPOSX1 DFFPOSX1_783 ( .CLK(clk_i_bF_buf39), .D(u2_u4_b1_last_row_5__FF_INPUT), .Q(u2_u4_b1_last_row_5_) );
  DFFPOSX1 DFFPOSX1_784 ( .CLK(clk_i_bF_buf38), .D(u2_u4_b1_last_row_6__FF_INPUT), .Q(u2_u4_b1_last_row_6_) );
  DFFPOSX1 DFFPOSX1_785 ( .CLK(clk_i_bF_buf37), .D(u2_u4_b1_last_row_7__FF_INPUT), .Q(u2_u4_b1_last_row_7_) );
  DFFPOSX1 DFFPOSX1_786 ( .CLK(clk_i_bF_buf36), .D(u2_u4_b1_last_row_8__FF_INPUT), .Q(u2_u4_b1_last_row_8_) );
  DFFPOSX1 DFFPOSX1_787 ( .CLK(clk_i_bF_buf35), .D(u2_u4_b1_last_row_9__FF_INPUT), .Q(u2_u4_b1_last_row_9_) );
  DFFPOSX1 DFFPOSX1_788 ( .CLK(clk_i_bF_buf34), .D(u2_u4_b1_last_row_10__FF_INPUT), .Q(u2_u4_b1_last_row_10_) );
  DFFPOSX1 DFFPOSX1_789 ( .CLK(clk_i_bF_buf33), .D(u2_u4_b1_last_row_11__FF_INPUT), .Q(u2_u4_b1_last_row_11_) );
  DFFPOSX1 DFFPOSX1_79 ( .CLK(clk_i_bF_buf45), .D(u0_u0_csc_5__FF_INPUT), .Q(u0_csc0_5_) );
  DFFPOSX1 DFFPOSX1_790 ( .CLK(clk_i_bF_buf32), .D(u2_u4_b1_last_row_12__FF_INPUT), .Q(u2_u4_b1_last_row_12_) );
  DFFPOSX1 DFFPOSX1_791 ( .CLK(clk_i_bF_buf31), .D(u2_u4_b0_last_row_0__FF_INPUT), .Q(u2_u4_b0_last_row_0_) );
  DFFPOSX1 DFFPOSX1_792 ( .CLK(clk_i_bF_buf30), .D(u2_u4_b0_last_row_1__FF_INPUT), .Q(u2_u4_b0_last_row_1_) );
  DFFPOSX1 DFFPOSX1_793 ( .CLK(clk_i_bF_buf29), .D(u2_u4_b0_last_row_2__FF_INPUT), .Q(u2_u4_b0_last_row_2_) );
  DFFPOSX1 DFFPOSX1_794 ( .CLK(clk_i_bF_buf28), .D(u2_u4_b0_last_row_3__FF_INPUT), .Q(u2_u4_b0_last_row_3_) );
  DFFPOSX1 DFFPOSX1_795 ( .CLK(clk_i_bF_buf27), .D(u2_u4_b0_last_row_4__FF_INPUT), .Q(u2_u4_b0_last_row_4_) );
  DFFPOSX1 DFFPOSX1_796 ( .CLK(clk_i_bF_buf26), .D(u2_u4_b0_last_row_5__FF_INPUT), .Q(u2_u4_b0_last_row_5_) );
  DFFPOSX1 DFFPOSX1_797 ( .CLK(clk_i_bF_buf25), .D(u2_u4_b0_last_row_6__FF_INPUT), .Q(u2_u4_b0_last_row_6_) );
  DFFPOSX1 DFFPOSX1_798 ( .CLK(clk_i_bF_buf24), .D(u2_u4_b0_last_row_7__FF_INPUT), .Q(u2_u4_b0_last_row_7_) );
  DFFPOSX1 DFFPOSX1_799 ( .CLK(clk_i_bF_buf23), .D(u2_u4_b0_last_row_8__FF_INPUT), .Q(u2_u4_b0_last_row_8_) );
  DFFPOSX1 DFFPOSX1_8 ( .CLK(clk_i_bF_buf118), .D(u0_poc_4__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56321_4_) );
  DFFPOSX1 DFFPOSX1_80 ( .CLK(clk_i_bF_buf44), .D(u0_u0_csc_6__FF_INPUT), .Q(u0_csc0_6_) );
  DFFPOSX1 DFFPOSX1_800 ( .CLK(clk_i_bF_buf22), .D(u2_u4_b0_last_row_9__FF_INPUT), .Q(u2_u4_b0_last_row_9_) );
  DFFPOSX1 DFFPOSX1_801 ( .CLK(clk_i_bF_buf21), .D(u2_u4_b0_last_row_10__FF_INPUT), .Q(u2_u4_b0_last_row_10_) );
  DFFPOSX1 DFFPOSX1_802 ( .CLK(clk_i_bF_buf20), .D(u2_u4_b0_last_row_11__FF_INPUT), .Q(u2_u4_b0_last_row_11_) );
  DFFPOSX1 DFFPOSX1_803 ( .CLK(clk_i_bF_buf19), .D(u2_u4_b0_last_row_12__FF_INPUT), .Q(u2_u4_b0_last_row_12_) );
  DFFPOSX1 DFFPOSX1_804 ( .CLK(clk_i_bF_buf14), .D(u2_u5_b3_last_row_0__FF_INPUT), .Q(u2_u5_b3_last_row_0_) );
  DFFPOSX1 DFFPOSX1_805 ( .CLK(clk_i_bF_buf13), .D(u2_u5_b3_last_row_1__FF_INPUT), .Q(u2_u5_b3_last_row_1_) );
  DFFPOSX1 DFFPOSX1_806 ( .CLK(clk_i_bF_buf12), .D(u2_u5_b3_last_row_2__FF_INPUT), .Q(u2_u5_b3_last_row_2_) );
  DFFPOSX1 DFFPOSX1_807 ( .CLK(clk_i_bF_buf11), .D(u2_u5_b3_last_row_3__FF_INPUT), .Q(u2_u5_b3_last_row_3_) );
  DFFPOSX1 DFFPOSX1_808 ( .CLK(clk_i_bF_buf10), .D(u2_u5_b3_last_row_4__FF_INPUT), .Q(u2_u5_b3_last_row_4_) );
  DFFPOSX1 DFFPOSX1_809 ( .CLK(clk_i_bF_buf9), .D(u2_u5_b3_last_row_5__FF_INPUT), .Q(u2_u5_b3_last_row_5_) );
  DFFPOSX1 DFFPOSX1_81 ( .CLK(clk_i_bF_buf43), .D(u0_u0_csc_7__FF_INPUT), .Q(u0_csc0_7_) );
  DFFPOSX1 DFFPOSX1_810 ( .CLK(clk_i_bF_buf8), .D(u2_u5_b3_last_row_6__FF_INPUT), .Q(u2_u5_b3_last_row_6_) );
  DFFPOSX1 DFFPOSX1_811 ( .CLK(clk_i_bF_buf7), .D(u2_u5_b3_last_row_7__FF_INPUT), .Q(u2_u5_b3_last_row_7_) );
  DFFPOSX1 DFFPOSX1_812 ( .CLK(clk_i_bF_buf6), .D(u2_u5_b3_last_row_8__FF_INPUT), .Q(u2_u5_b3_last_row_8_) );
  DFFPOSX1 DFFPOSX1_813 ( .CLK(clk_i_bF_buf5), .D(u2_u5_b3_last_row_9__FF_INPUT), .Q(u2_u5_b3_last_row_9_) );
  DFFPOSX1 DFFPOSX1_814 ( .CLK(clk_i_bF_buf4), .D(u2_u5_b3_last_row_10__FF_INPUT), .Q(u2_u5_b3_last_row_10_) );
  DFFPOSX1 DFFPOSX1_815 ( .CLK(clk_i_bF_buf3), .D(u2_u5_b3_last_row_11__FF_INPUT), .Q(u2_u5_b3_last_row_11_) );
  DFFPOSX1 DFFPOSX1_816 ( .CLK(clk_i_bF_buf2), .D(u2_u5_b3_last_row_12__FF_INPUT), .Q(u2_u5_b3_last_row_12_) );
  DFFPOSX1 DFFPOSX1_817 ( .CLK(clk_i_bF_buf1), .D(u2_u5_b2_last_row_0__FF_INPUT), .Q(u2_u5_b2_last_row_0_) );
  DFFPOSX1 DFFPOSX1_818 ( .CLK(clk_i_bF_buf0), .D(u2_u5_b2_last_row_1__FF_INPUT), .Q(u2_u5_b2_last_row_1_) );
  DFFPOSX1 DFFPOSX1_819 ( .CLK(clk_i_bF_buf125), .D(u2_u5_b2_last_row_2__FF_INPUT), .Q(u2_u5_b2_last_row_2_) );
  DFFPOSX1 DFFPOSX1_82 ( .CLK(clk_i_bF_buf42), .D(u0_u0_csc_8__FF_INPUT), .Q(u0_csc0_8_) );
  DFFPOSX1 DFFPOSX1_820 ( .CLK(clk_i_bF_buf124), .D(u2_u5_b2_last_row_3__FF_INPUT), .Q(u2_u5_b2_last_row_3_) );
  DFFPOSX1 DFFPOSX1_821 ( .CLK(clk_i_bF_buf123), .D(u2_u5_b2_last_row_4__FF_INPUT), .Q(u2_u5_b2_last_row_4_) );
  DFFPOSX1 DFFPOSX1_822 ( .CLK(clk_i_bF_buf122), .D(u2_u5_b2_last_row_5__FF_INPUT), .Q(u2_u5_b2_last_row_5_) );
  DFFPOSX1 DFFPOSX1_823 ( .CLK(clk_i_bF_buf121), .D(u2_u5_b2_last_row_6__FF_INPUT), .Q(u2_u5_b2_last_row_6_) );
  DFFPOSX1 DFFPOSX1_824 ( .CLK(clk_i_bF_buf120), .D(u2_u5_b2_last_row_7__FF_INPUT), .Q(u2_u5_b2_last_row_7_) );
  DFFPOSX1 DFFPOSX1_825 ( .CLK(clk_i_bF_buf119), .D(u2_u5_b2_last_row_8__FF_INPUT), .Q(u2_u5_b2_last_row_8_) );
  DFFPOSX1 DFFPOSX1_826 ( .CLK(clk_i_bF_buf118), .D(u2_u5_b2_last_row_9__FF_INPUT), .Q(u2_u5_b2_last_row_9_) );
  DFFPOSX1 DFFPOSX1_827 ( .CLK(clk_i_bF_buf117), .D(u2_u5_b2_last_row_10__FF_INPUT), .Q(u2_u5_b2_last_row_10_) );
  DFFPOSX1 DFFPOSX1_828 ( .CLK(clk_i_bF_buf116), .D(u2_u5_b2_last_row_11__FF_INPUT), .Q(u2_u5_b2_last_row_11_) );
  DFFPOSX1 DFFPOSX1_829 ( .CLK(clk_i_bF_buf115), .D(u2_u5_b2_last_row_12__FF_INPUT), .Q(u2_u5_b2_last_row_12_) );
  DFFPOSX1 DFFPOSX1_83 ( .CLK(clk_i_bF_buf41), .D(u0_u0_csc_9__FF_INPUT), .Q(u0_csc0_9_) );
  DFFPOSX1 DFFPOSX1_830 ( .CLK(clk_i_bF_buf114), .D(u2_u5_b1_last_row_0__FF_INPUT), .Q(u2_u5_b1_last_row_0_) );
  DFFPOSX1 DFFPOSX1_831 ( .CLK(clk_i_bF_buf113), .D(u2_u5_b1_last_row_1__FF_INPUT), .Q(u2_u5_b1_last_row_1_) );
  DFFPOSX1 DFFPOSX1_832 ( .CLK(clk_i_bF_buf112), .D(u2_u5_b1_last_row_2__FF_INPUT), .Q(u2_u5_b1_last_row_2_) );
  DFFPOSX1 DFFPOSX1_833 ( .CLK(clk_i_bF_buf111), .D(u2_u5_b1_last_row_3__FF_INPUT), .Q(u2_u5_b1_last_row_3_) );
  DFFPOSX1 DFFPOSX1_834 ( .CLK(clk_i_bF_buf110), .D(u2_u5_b1_last_row_4__FF_INPUT), .Q(u2_u5_b1_last_row_4_) );
  DFFPOSX1 DFFPOSX1_835 ( .CLK(clk_i_bF_buf109), .D(u2_u5_b1_last_row_5__FF_INPUT), .Q(u2_u5_b1_last_row_5_) );
  DFFPOSX1 DFFPOSX1_836 ( .CLK(clk_i_bF_buf108), .D(u2_u5_b1_last_row_6__FF_INPUT), .Q(u2_u5_b1_last_row_6_) );
  DFFPOSX1 DFFPOSX1_837 ( .CLK(clk_i_bF_buf107), .D(u2_u5_b1_last_row_7__FF_INPUT), .Q(u2_u5_b1_last_row_7_) );
  DFFPOSX1 DFFPOSX1_838 ( .CLK(clk_i_bF_buf106), .D(u2_u5_b1_last_row_8__FF_INPUT), .Q(u2_u5_b1_last_row_8_) );
  DFFPOSX1 DFFPOSX1_839 ( .CLK(clk_i_bF_buf105), .D(u2_u5_b1_last_row_9__FF_INPUT), .Q(u2_u5_b1_last_row_9_) );
  DFFPOSX1 DFFPOSX1_84 ( .CLK(clk_i_bF_buf40), .D(u0_u0_csc_10__FF_INPUT), .Q(u0_csc0_10_) );
  DFFPOSX1 DFFPOSX1_840 ( .CLK(clk_i_bF_buf104), .D(u2_u5_b1_last_row_10__FF_INPUT), .Q(u2_u5_b1_last_row_10_) );
  DFFPOSX1 DFFPOSX1_841 ( .CLK(clk_i_bF_buf103), .D(u2_u5_b1_last_row_11__FF_INPUT), .Q(u2_u5_b1_last_row_11_) );
  DFFPOSX1 DFFPOSX1_842 ( .CLK(clk_i_bF_buf102), .D(u2_u5_b1_last_row_12__FF_INPUT), .Q(u2_u5_b1_last_row_12_) );
  DFFPOSX1 DFFPOSX1_843 ( .CLK(clk_i_bF_buf101), .D(u2_u5_b0_last_row_0__FF_INPUT), .Q(u2_u5_b0_last_row_0_) );
  DFFPOSX1 DFFPOSX1_844 ( .CLK(clk_i_bF_buf100), .D(u2_u5_b0_last_row_1__FF_INPUT), .Q(u2_u5_b0_last_row_1_) );
  DFFPOSX1 DFFPOSX1_845 ( .CLK(clk_i_bF_buf99), .D(u2_u5_b0_last_row_2__FF_INPUT), .Q(u2_u5_b0_last_row_2_) );
  DFFPOSX1 DFFPOSX1_846 ( .CLK(clk_i_bF_buf98), .D(u2_u5_b0_last_row_3__FF_INPUT), .Q(u2_u5_b0_last_row_3_) );
  DFFPOSX1 DFFPOSX1_847 ( .CLK(clk_i_bF_buf97), .D(u2_u5_b0_last_row_4__FF_INPUT), .Q(u2_u5_b0_last_row_4_) );
  DFFPOSX1 DFFPOSX1_848 ( .CLK(clk_i_bF_buf96), .D(u2_u5_b0_last_row_5__FF_INPUT), .Q(u2_u5_b0_last_row_5_) );
  DFFPOSX1 DFFPOSX1_849 ( .CLK(clk_i_bF_buf95), .D(u2_u5_b0_last_row_6__FF_INPUT), .Q(u2_u5_b0_last_row_6_) );
  DFFPOSX1 DFFPOSX1_85 ( .CLK(clk_i_bF_buf39), .D(u0_u0_csc_11__FF_INPUT), .Q(u0_csc0_11_) );
  DFFPOSX1 DFFPOSX1_850 ( .CLK(clk_i_bF_buf94), .D(u2_u5_b0_last_row_7__FF_INPUT), .Q(u2_u5_b0_last_row_7_) );
  DFFPOSX1 DFFPOSX1_851 ( .CLK(clk_i_bF_buf93), .D(u2_u5_b0_last_row_8__FF_INPUT), .Q(u2_u5_b0_last_row_8_) );
  DFFPOSX1 DFFPOSX1_852 ( .CLK(clk_i_bF_buf92), .D(u2_u5_b0_last_row_9__FF_INPUT), .Q(u2_u5_b0_last_row_9_) );
  DFFPOSX1 DFFPOSX1_853 ( .CLK(clk_i_bF_buf91), .D(u2_u5_b0_last_row_10__FF_INPUT), .Q(u2_u5_b0_last_row_10_) );
  DFFPOSX1 DFFPOSX1_854 ( .CLK(clk_i_bF_buf90), .D(u2_u5_b0_last_row_11__FF_INPUT), .Q(u2_u5_b0_last_row_11_) );
  DFFPOSX1 DFFPOSX1_855 ( .CLK(clk_i_bF_buf89), .D(u2_u5_b0_last_row_12__FF_INPUT), .Q(u2_u5_b0_last_row_12_) );
  DFFPOSX1 DFFPOSX1_856 ( .CLK(clk_i_bF_buf84), .D(u3_mc_dp_o_0__FF_INPUT), .Q(mc_dp_od_0_) );
  DFFPOSX1 DFFPOSX1_857 ( .CLK(clk_i_bF_buf83), .D(u3_mc_dp_o_1__FF_INPUT), .Q(mc_dp_od_1_) );
  DFFPOSX1 DFFPOSX1_858 ( .CLK(clk_i_bF_buf82), .D(u3_mc_dp_o_2__FF_INPUT), .Q(mc_dp_od_2_) );
  DFFPOSX1 DFFPOSX1_859 ( .CLK(clk_i_bF_buf81), .D(u3_mc_dp_o_3__FF_INPUT), .Q(mc_dp_od_3_) );
  DFFPOSX1 DFFPOSX1_86 ( .CLK(clk_i_bF_buf38), .D(u0_u0_csc_12__FF_INPUT), .Q(u0_csc0_12_) );
  DFFPOSX1 DFFPOSX1_860 ( .CLK(clk_i_bF_buf80), .D(u3_byte2_0__FF_INPUT), .Q(u3_byte2_0_) );
  DFFPOSX1 DFFPOSX1_861 ( .CLK(clk_i_bF_buf79), .D(u3_byte2_1__FF_INPUT), .Q(u3_byte2_1_) );
  DFFPOSX1 DFFPOSX1_862 ( .CLK(clk_i_bF_buf78), .D(u3_byte2_2__FF_INPUT), .Q(u3_byte2_2_) );
  DFFPOSX1 DFFPOSX1_863 ( .CLK(clk_i_bF_buf77), .D(u3_byte2_3__FF_INPUT), .Q(u3_byte2_3_) );
  DFFPOSX1 DFFPOSX1_864 ( .CLK(clk_i_bF_buf76), .D(u3_byte2_4__FF_INPUT), .Q(u3_byte2_4_) );
  DFFPOSX1 DFFPOSX1_865 ( .CLK(clk_i_bF_buf75), .D(u3_byte2_5__FF_INPUT), .Q(u3_byte2_5_) );
  DFFPOSX1 DFFPOSX1_866 ( .CLK(clk_i_bF_buf74), .D(u3_byte2_6__FF_INPUT), .Q(u3_byte2_6_) );
  DFFPOSX1 DFFPOSX1_867 ( .CLK(clk_i_bF_buf73), .D(u3_byte2_7__FF_INPUT), .Q(u3_byte2_7_) );
  DFFPOSX1 DFFPOSX1_868 ( .CLK(clk_i_bF_buf72), .D(u3_byte1_0__FF_INPUT), .Q(u3_byte1_0_) );
  DFFPOSX1 DFFPOSX1_869 ( .CLK(clk_i_bF_buf71), .D(u3_byte1_1__FF_INPUT), .Q(u3_byte1_1_) );
  DFFPOSX1 DFFPOSX1_87 ( .CLK(clk_i_bF_buf37), .D(u0_u0_csc_13__FF_INPUT), .Q(u0_csc0_13_) );
  DFFPOSX1 DFFPOSX1_870 ( .CLK(clk_i_bF_buf70), .D(u3_byte1_2__FF_INPUT), .Q(u3_byte1_2_) );
  DFFPOSX1 DFFPOSX1_871 ( .CLK(clk_i_bF_buf69), .D(u3_byte1_3__FF_INPUT), .Q(u3_byte1_3_) );
  DFFPOSX1 DFFPOSX1_872 ( .CLK(clk_i_bF_buf68), .D(u3_byte1_4__FF_INPUT), .Q(u3_byte1_4_) );
  DFFPOSX1 DFFPOSX1_873 ( .CLK(clk_i_bF_buf67), .D(u3_byte1_5__FF_INPUT), .Q(u3_byte1_5_) );
  DFFPOSX1 DFFPOSX1_874 ( .CLK(clk_i_bF_buf66), .D(u3_byte1_6__FF_INPUT), .Q(u3_byte1_6_) );
  DFFPOSX1 DFFPOSX1_875 ( .CLK(clk_i_bF_buf65), .D(u3_byte1_7__FF_INPUT), .Q(u3_byte1_7_) );
  DFFPOSX1 DFFPOSX1_876 ( .CLK(clk_i_bF_buf64), .D(u3_byte0_0__FF_INPUT), .Q(u3_byte0_0_) );
  DFFPOSX1 DFFPOSX1_877 ( .CLK(clk_i_bF_buf63), .D(u3_byte0_1__FF_INPUT), .Q(u3_byte0_1_) );
  DFFPOSX1 DFFPOSX1_878 ( .CLK(clk_i_bF_buf62), .D(u3_byte0_2__FF_INPUT), .Q(u3_byte0_2_) );
  DFFPOSX1 DFFPOSX1_879 ( .CLK(clk_i_bF_buf61), .D(u3_byte0_3__FF_INPUT), .Q(u3_byte0_3_) );
  DFFPOSX1 DFFPOSX1_88 ( .CLK(clk_i_bF_buf36), .D(u0_u0_csc_14__FF_INPUT), .Q(u0_csc0_14_) );
  DFFPOSX1 DFFPOSX1_880 ( .CLK(clk_i_bF_buf60), .D(u3_byte0_4__FF_INPUT), .Q(u3_byte0_4_) );
  DFFPOSX1 DFFPOSX1_881 ( .CLK(clk_i_bF_buf59), .D(u3_byte0_5__FF_INPUT), .Q(u3_byte0_5_) );
  DFFPOSX1 DFFPOSX1_882 ( .CLK(clk_i_bF_buf58), .D(u3_byte0_6__FF_INPUT), .Q(u3_byte0_6_) );
  DFFPOSX1 DFFPOSX1_883 ( .CLK(clk_i_bF_buf57), .D(u3_byte0_7__FF_INPUT), .Q(u3_byte0_7_) );
  DFFPOSX1 DFFPOSX1_884 ( .CLK(clk_i_bF_buf56), .D(u3_mc_data_o_0__FF_INPUT), .Q(mc_data_od_0_) );
  DFFPOSX1 DFFPOSX1_885 ( .CLK(clk_i_bF_buf55), .D(u3_mc_data_o_1__FF_INPUT), .Q(mc_data_od_1_) );
  DFFPOSX1 DFFPOSX1_886 ( .CLK(clk_i_bF_buf54), .D(u3_mc_data_o_2__FF_INPUT), .Q(mc_data_od_2_) );
  DFFPOSX1 DFFPOSX1_887 ( .CLK(clk_i_bF_buf53), .D(u3_mc_data_o_3__FF_INPUT), .Q(mc_data_od_3_) );
  DFFPOSX1 DFFPOSX1_888 ( .CLK(clk_i_bF_buf52), .D(u3_mc_data_o_4__FF_INPUT), .Q(mc_data_od_4_) );
  DFFPOSX1 DFFPOSX1_889 ( .CLK(clk_i_bF_buf51), .D(u3_mc_data_o_5__FF_INPUT), .Q(mc_data_od_5_) );
  DFFPOSX1 DFFPOSX1_89 ( .CLK(clk_i_bF_buf35), .D(u0_u0_csc_15__FF_INPUT), .Q(u0_csc0_15_) );
  DFFPOSX1 DFFPOSX1_890 ( .CLK(clk_i_bF_buf50), .D(u3_mc_data_o_6__FF_INPUT), .Q(mc_data_od_6_) );
  DFFPOSX1 DFFPOSX1_891 ( .CLK(clk_i_bF_buf49), .D(u3_mc_data_o_7__FF_INPUT), .Q(mc_data_od_7_) );
  DFFPOSX1 DFFPOSX1_892 ( .CLK(clk_i_bF_buf48), .D(u3_mc_data_o_8__FF_INPUT), .Q(mc_data_od_8_) );
  DFFPOSX1 DFFPOSX1_893 ( .CLK(clk_i_bF_buf47), .D(u3_mc_data_o_9__FF_INPUT), .Q(mc_data_od_9_) );
  DFFPOSX1 DFFPOSX1_894 ( .CLK(clk_i_bF_buf46), .D(u3_mc_data_o_10__FF_INPUT), .Q(mc_data_od_10_) );
  DFFPOSX1 DFFPOSX1_895 ( .CLK(clk_i_bF_buf45), .D(u3_mc_data_o_11__FF_INPUT), .Q(mc_data_od_11_) );
  DFFPOSX1 DFFPOSX1_896 ( .CLK(clk_i_bF_buf44), .D(u3_mc_data_o_12__FF_INPUT), .Q(mc_data_od_12_) );
  DFFPOSX1 DFFPOSX1_897 ( .CLK(clk_i_bF_buf43), .D(u3_mc_data_o_13__FF_INPUT), .Q(mc_data_od_13_) );
  DFFPOSX1 DFFPOSX1_898 ( .CLK(clk_i_bF_buf42), .D(u3_mc_data_o_14__FF_INPUT), .Q(mc_data_od_14_) );
  DFFPOSX1 DFFPOSX1_899 ( .CLK(clk_i_bF_buf41), .D(u3_mc_data_o_15__FF_INPUT), .Q(mc_data_od_15_) );
  DFFPOSX1 DFFPOSX1_9 ( .CLK(clk_i_bF_buf117), .D(u0_poc_5__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56321_5_) );
  DFFPOSX1 DFFPOSX1_90 ( .CLK(clk_i_bF_buf34), .D(u0_u0_csc_16__FF_INPUT), .Q(u0_csc0_16_) );
  DFFPOSX1 DFFPOSX1_900 ( .CLK(clk_i_bF_buf40), .D(u3_mc_data_o_16__FF_INPUT), .Q(mc_data_od_16_) );
  DFFPOSX1 DFFPOSX1_901 ( .CLK(clk_i_bF_buf39), .D(u3_mc_data_o_17__FF_INPUT), .Q(mc_data_od_17_) );
  DFFPOSX1 DFFPOSX1_902 ( .CLK(clk_i_bF_buf38), .D(u3_mc_data_o_18__FF_INPUT), .Q(mc_data_od_18_) );
  DFFPOSX1 DFFPOSX1_903 ( .CLK(clk_i_bF_buf37), .D(u3_mc_data_o_19__FF_INPUT), .Q(mc_data_od_19_) );
  DFFPOSX1 DFFPOSX1_904 ( .CLK(clk_i_bF_buf36), .D(u3_mc_data_o_20__FF_INPUT), .Q(mc_data_od_20_) );
  DFFPOSX1 DFFPOSX1_905 ( .CLK(clk_i_bF_buf35), .D(u3_mc_data_o_21__FF_INPUT), .Q(mc_data_od_21_) );
  DFFPOSX1 DFFPOSX1_906 ( .CLK(clk_i_bF_buf34), .D(u3_mc_data_o_22__FF_INPUT), .Q(mc_data_od_22_) );
  DFFPOSX1 DFFPOSX1_907 ( .CLK(clk_i_bF_buf33), .D(u3_mc_data_o_23__FF_INPUT), .Q(mc_data_od_23_) );
  DFFPOSX1 DFFPOSX1_908 ( .CLK(clk_i_bF_buf32), .D(u3_mc_data_o_24__FF_INPUT), .Q(mc_data_od_24_) );
  DFFPOSX1 DFFPOSX1_909 ( .CLK(clk_i_bF_buf31), .D(u3_mc_data_o_25__FF_INPUT), .Q(mc_data_od_25_) );
  DFFPOSX1 DFFPOSX1_91 ( .CLK(clk_i_bF_buf33), .D(u0_u0_csc_17__FF_INPUT), .Q(u0_csc0_17_) );
  DFFPOSX1 DFFPOSX1_910 ( .CLK(clk_i_bF_buf30), .D(u3_mc_data_o_26__FF_INPUT), .Q(mc_data_od_26_) );
  DFFPOSX1 DFFPOSX1_911 ( .CLK(clk_i_bF_buf29), .D(u3_mc_data_o_27__FF_INPUT), .Q(mc_data_od_27_) );
  DFFPOSX1 DFFPOSX1_912 ( .CLK(clk_i_bF_buf28), .D(u3_mc_data_o_28__FF_INPUT), .Q(mc_data_od_28_) );
  DFFPOSX1 DFFPOSX1_913 ( .CLK(clk_i_bF_buf27), .D(u3_mc_data_o_29__FF_INPUT), .Q(mc_data_od_29_) );
  DFFPOSX1 DFFPOSX1_914 ( .CLK(clk_i_bF_buf26), .D(u3_mc_data_o_30__FF_INPUT), .Q(mc_data_od_30_) );
  DFFPOSX1 DFFPOSX1_915 ( .CLK(clk_i_bF_buf25), .D(u3_mc_data_o_31__FF_INPUT), .Q(mc_data_od_31_) );
  DFFPOSX1 DFFPOSX1_916 ( .CLK(clk_i_bF_buf24), .D(u3_u0_r3_0__FF_INPUT), .Q(u3_u0_r3_0_) );
  DFFPOSX1 DFFPOSX1_917 ( .CLK(clk_i_bF_buf23), .D(u3_u0_r3_1__FF_INPUT), .Q(u3_u0_r3_1_) );
  DFFPOSX1 DFFPOSX1_918 ( .CLK(clk_i_bF_buf22), .D(u3_u0_r3_2__FF_INPUT), .Q(u3_u0_r3_2_) );
  DFFPOSX1 DFFPOSX1_919 ( .CLK(clk_i_bF_buf21), .D(u3_u0_r3_3__FF_INPUT), .Q(u3_u0_r3_3_) );
  DFFPOSX1 DFFPOSX1_92 ( .CLK(clk_i_bF_buf32), .D(u0_u0_csc_18__FF_INPUT), .Q(u0_csc0_18_) );
  DFFPOSX1 DFFPOSX1_920 ( .CLK(clk_i_bF_buf20), .D(u3_u0_r3_4__FF_INPUT), .Q(u3_u0_r3_4_) );
  DFFPOSX1 DFFPOSX1_921 ( .CLK(clk_i_bF_buf19), .D(u3_u0_r3_5__FF_INPUT), .Q(u3_u0_r3_5_) );
  DFFPOSX1 DFFPOSX1_922 ( .CLK(clk_i_bF_buf18), .D(u3_u0_r3_6__FF_INPUT), .Q(u3_u0_r3_6_) );
  DFFPOSX1 DFFPOSX1_923 ( .CLK(clk_i_bF_buf17), .D(u3_u0_r3_7__FF_INPUT), .Q(u3_u0_r3_7_) );
  DFFPOSX1 DFFPOSX1_924 ( .CLK(clk_i_bF_buf16), .D(u3_u0_r3_8__FF_INPUT), .Q(u3_u0_r3_8_) );
  DFFPOSX1 DFFPOSX1_925 ( .CLK(clk_i_bF_buf15), .D(u3_u0_r3_9__FF_INPUT), .Q(u3_u0_r3_9_) );
  DFFPOSX1 DFFPOSX1_926 ( .CLK(clk_i_bF_buf14), .D(u3_u0_r3_10__FF_INPUT), .Q(u3_u0_r3_10_) );
  DFFPOSX1 DFFPOSX1_927 ( .CLK(clk_i_bF_buf13), .D(u3_u0_r3_11__FF_INPUT), .Q(u3_u0_r3_11_) );
  DFFPOSX1 DFFPOSX1_928 ( .CLK(clk_i_bF_buf12), .D(u3_u0_r3_12__FF_INPUT), .Q(u3_u0_r3_12_) );
  DFFPOSX1 DFFPOSX1_929 ( .CLK(clk_i_bF_buf11), .D(u3_u0_r3_13__FF_INPUT), .Q(u3_u0_r3_13_) );
  DFFPOSX1 DFFPOSX1_93 ( .CLK(clk_i_bF_buf31), .D(u0_u0_csc_19__FF_INPUT), .Q(u0_csc0_19_) );
  DFFPOSX1 DFFPOSX1_930 ( .CLK(clk_i_bF_buf10), .D(u3_u0_r3_14__FF_INPUT), .Q(u3_u0_r3_14_) );
  DFFPOSX1 DFFPOSX1_931 ( .CLK(clk_i_bF_buf9), .D(u3_u0_r3_15__FF_INPUT), .Q(u3_u0_r3_15_) );
  DFFPOSX1 DFFPOSX1_932 ( .CLK(clk_i_bF_buf8), .D(u3_u0_r3_16__FF_INPUT), .Q(u3_u0_r3_16_) );
  DFFPOSX1 DFFPOSX1_933 ( .CLK(clk_i_bF_buf7), .D(u3_u0_r3_17__FF_INPUT), .Q(u3_u0_r3_17_) );
  DFFPOSX1 DFFPOSX1_934 ( .CLK(clk_i_bF_buf6), .D(u3_u0_r3_18__FF_INPUT), .Q(u3_u0_r3_18_) );
  DFFPOSX1 DFFPOSX1_935 ( .CLK(clk_i_bF_buf5), .D(u3_u0_r3_19__FF_INPUT), .Q(u3_u0_r3_19_) );
  DFFPOSX1 DFFPOSX1_936 ( .CLK(clk_i_bF_buf4), .D(u3_u0_r3_20__FF_INPUT), .Q(u3_u0_r3_20_) );
  DFFPOSX1 DFFPOSX1_937 ( .CLK(clk_i_bF_buf3), .D(u3_u0_r3_21__FF_INPUT), .Q(u3_u0_r3_21_) );
  DFFPOSX1 DFFPOSX1_938 ( .CLK(clk_i_bF_buf2), .D(u3_u0_r3_22__FF_INPUT), .Q(u3_u0_r3_22_) );
  DFFPOSX1 DFFPOSX1_939 ( .CLK(clk_i_bF_buf1), .D(u3_u0_r3_23__FF_INPUT), .Q(u3_u0_r3_23_) );
  DFFPOSX1 DFFPOSX1_94 ( .CLK(clk_i_bF_buf30), .D(u0_u0_csc_20__FF_INPUT), .Q(u0_csc0_20_) );
  DFFPOSX1 DFFPOSX1_940 ( .CLK(clk_i_bF_buf0), .D(u3_u0_r3_24__FF_INPUT), .Q(u3_u0_r3_24_) );
  DFFPOSX1 DFFPOSX1_941 ( .CLK(clk_i_bF_buf125), .D(u3_u0_r3_25__FF_INPUT), .Q(u3_u0_r3_25_) );
  DFFPOSX1 DFFPOSX1_942 ( .CLK(clk_i_bF_buf124), .D(u3_u0_r3_26__FF_INPUT), .Q(u3_u0_r3_26_) );
  DFFPOSX1 DFFPOSX1_943 ( .CLK(clk_i_bF_buf123), .D(u3_u0_r3_27__FF_INPUT), .Q(u3_u0_r3_27_) );
  DFFPOSX1 DFFPOSX1_944 ( .CLK(clk_i_bF_buf122), .D(u3_u0_r3_28__FF_INPUT), .Q(u3_u0_r3_28_) );
  DFFPOSX1 DFFPOSX1_945 ( .CLK(clk_i_bF_buf121), .D(u3_u0_r3_29__FF_INPUT), .Q(u3_u0_r3_29_) );
  DFFPOSX1 DFFPOSX1_946 ( .CLK(clk_i_bF_buf120), .D(u3_u0_r3_30__FF_INPUT), .Q(u3_u0_r3_30_) );
  DFFPOSX1 DFFPOSX1_947 ( .CLK(clk_i_bF_buf119), .D(u3_u0_r3_31__FF_INPUT), .Q(u3_u0_r3_31_) );
  DFFPOSX1 DFFPOSX1_948 ( .CLK(clk_i_bF_buf118), .D(u3_u0_r3_32__FF_INPUT), .Q(u3_u0_r3_32_) );
  DFFPOSX1 DFFPOSX1_949 ( .CLK(clk_i_bF_buf117), .D(u3_u0_r3_33__FF_INPUT), .Q(u3_u0_r3_33_) );
  DFFPOSX1 DFFPOSX1_95 ( .CLK(clk_i_bF_buf29), .D(u0_u0_csc_21__FF_INPUT), .Q(u0_csc0_21_) );
  DFFPOSX1 DFFPOSX1_950 ( .CLK(clk_i_bF_buf116), .D(u3_u0_r3_34__FF_INPUT), .Q(u3_u0_r3_34_) );
  DFFPOSX1 DFFPOSX1_951 ( .CLK(clk_i_bF_buf115), .D(u3_u0_r3_35__FF_INPUT), .Q(u3_u0_r3_35_) );
  DFFPOSX1 DFFPOSX1_952 ( .CLK(clk_i_bF_buf114), .D(u3_u0_r2_0__FF_INPUT), .Q(u3_u0_r2_0_) );
  DFFPOSX1 DFFPOSX1_953 ( .CLK(clk_i_bF_buf113), .D(u3_u0_r2_1__FF_INPUT), .Q(u3_u0_r2_1_) );
  DFFPOSX1 DFFPOSX1_954 ( .CLK(clk_i_bF_buf112), .D(u3_u0_r2_2__FF_INPUT), .Q(u3_u0_r2_2_) );
  DFFPOSX1 DFFPOSX1_955 ( .CLK(clk_i_bF_buf111), .D(u3_u0_r2_3__FF_INPUT), .Q(u3_u0_r2_3_) );
  DFFPOSX1 DFFPOSX1_956 ( .CLK(clk_i_bF_buf110), .D(u3_u0_r2_4__FF_INPUT), .Q(u3_u0_r2_4_) );
  DFFPOSX1 DFFPOSX1_957 ( .CLK(clk_i_bF_buf109), .D(u3_u0_r2_5__FF_INPUT), .Q(u3_u0_r2_5_) );
  DFFPOSX1 DFFPOSX1_958 ( .CLK(clk_i_bF_buf108), .D(u3_u0_r2_6__FF_INPUT), .Q(u3_u0_r2_6_) );
  DFFPOSX1 DFFPOSX1_959 ( .CLK(clk_i_bF_buf107), .D(u3_u0_r2_7__FF_INPUT), .Q(u3_u0_r2_7_) );
  DFFPOSX1 DFFPOSX1_96 ( .CLK(clk_i_bF_buf28), .D(u0_u0_csc_22__FF_INPUT), .Q(u0_csc0_22_) );
  DFFPOSX1 DFFPOSX1_960 ( .CLK(clk_i_bF_buf106), .D(u3_u0_r2_8__FF_INPUT), .Q(u3_u0_r2_8_) );
  DFFPOSX1 DFFPOSX1_961 ( .CLK(clk_i_bF_buf105), .D(u3_u0_r2_9__FF_INPUT), .Q(u3_u0_r2_9_) );
  DFFPOSX1 DFFPOSX1_962 ( .CLK(clk_i_bF_buf104), .D(u3_u0_r2_10__FF_INPUT), .Q(u3_u0_r2_10_) );
  DFFPOSX1 DFFPOSX1_963 ( .CLK(clk_i_bF_buf103), .D(u3_u0_r2_11__FF_INPUT), .Q(u3_u0_r2_11_) );
  DFFPOSX1 DFFPOSX1_964 ( .CLK(clk_i_bF_buf102), .D(u3_u0_r2_12__FF_INPUT), .Q(u3_u0_r2_12_) );
  DFFPOSX1 DFFPOSX1_965 ( .CLK(clk_i_bF_buf101), .D(u3_u0_r2_13__FF_INPUT), .Q(u3_u0_r2_13_) );
  DFFPOSX1 DFFPOSX1_966 ( .CLK(clk_i_bF_buf100), .D(u3_u0_r2_14__FF_INPUT), .Q(u3_u0_r2_14_) );
  DFFPOSX1 DFFPOSX1_967 ( .CLK(clk_i_bF_buf99), .D(u3_u0_r2_15__FF_INPUT), .Q(u3_u0_r2_15_) );
  DFFPOSX1 DFFPOSX1_968 ( .CLK(clk_i_bF_buf98), .D(u3_u0_r2_16__FF_INPUT), .Q(u3_u0_r2_16_) );
  DFFPOSX1 DFFPOSX1_969 ( .CLK(clk_i_bF_buf97), .D(u3_u0_r2_17__FF_INPUT), .Q(u3_u0_r2_17_) );
  DFFPOSX1 DFFPOSX1_97 ( .CLK(clk_i_bF_buf27), .D(u0_u0_csc_23__FF_INPUT), .Q(u0_csc0_23_) );
  DFFPOSX1 DFFPOSX1_970 ( .CLK(clk_i_bF_buf96), .D(u3_u0_r2_18__FF_INPUT), .Q(u3_u0_r2_18_) );
  DFFPOSX1 DFFPOSX1_971 ( .CLK(clk_i_bF_buf95), .D(u3_u0_r2_19__FF_INPUT), .Q(u3_u0_r2_19_) );
  DFFPOSX1 DFFPOSX1_972 ( .CLK(clk_i_bF_buf94), .D(u3_u0_r2_20__FF_INPUT), .Q(u3_u0_r2_20_) );
  DFFPOSX1 DFFPOSX1_973 ( .CLK(clk_i_bF_buf93), .D(u3_u0_r2_21__FF_INPUT), .Q(u3_u0_r2_21_) );
  DFFPOSX1 DFFPOSX1_974 ( .CLK(clk_i_bF_buf92), .D(u3_u0_r2_22__FF_INPUT), .Q(u3_u0_r2_22_) );
  DFFPOSX1 DFFPOSX1_975 ( .CLK(clk_i_bF_buf91), .D(u3_u0_r2_23__FF_INPUT), .Q(u3_u0_r2_23_) );
  DFFPOSX1 DFFPOSX1_976 ( .CLK(clk_i_bF_buf90), .D(u3_u0_r2_24__FF_INPUT), .Q(u3_u0_r2_24_) );
  DFFPOSX1 DFFPOSX1_977 ( .CLK(clk_i_bF_buf89), .D(u3_u0_r2_25__FF_INPUT), .Q(u3_u0_r2_25_) );
  DFFPOSX1 DFFPOSX1_978 ( .CLK(clk_i_bF_buf88), .D(u3_u0_r2_26__FF_INPUT), .Q(u3_u0_r2_26_) );
  DFFPOSX1 DFFPOSX1_979 ( .CLK(clk_i_bF_buf87), .D(u3_u0_r2_27__FF_INPUT), .Q(u3_u0_r2_27_) );
  DFFPOSX1 DFFPOSX1_98 ( .CLK(clk_i_bF_buf26), .D(u0_u0_csc_24__FF_INPUT), .Q(u0_csc0_24_) );
  DFFPOSX1 DFFPOSX1_980 ( .CLK(clk_i_bF_buf86), .D(u3_u0_r2_28__FF_INPUT), .Q(u3_u0_r2_28_) );
  DFFPOSX1 DFFPOSX1_981 ( .CLK(clk_i_bF_buf85), .D(u3_u0_r2_29__FF_INPUT), .Q(u3_u0_r2_29_) );
  DFFPOSX1 DFFPOSX1_982 ( .CLK(clk_i_bF_buf84), .D(u3_u0_r2_30__FF_INPUT), .Q(u3_u0_r2_30_) );
  DFFPOSX1 DFFPOSX1_983 ( .CLK(clk_i_bF_buf83), .D(u3_u0_r2_31__FF_INPUT), .Q(u3_u0_r2_31_) );
  DFFPOSX1 DFFPOSX1_984 ( .CLK(clk_i_bF_buf82), .D(u3_u0_r2_32__FF_INPUT), .Q(u3_u0_r2_32_) );
  DFFPOSX1 DFFPOSX1_985 ( .CLK(clk_i_bF_buf81), .D(u3_u0_r2_33__FF_INPUT), .Q(u3_u0_r2_33_) );
  DFFPOSX1 DFFPOSX1_986 ( .CLK(clk_i_bF_buf80), .D(u3_u0_r2_34__FF_INPUT), .Q(u3_u0_r2_34_) );
  DFFPOSX1 DFFPOSX1_987 ( .CLK(clk_i_bF_buf79), .D(u3_u0_r2_35__FF_INPUT), .Q(u3_u0_r2_35_) );
  DFFPOSX1 DFFPOSX1_988 ( .CLK(clk_i_bF_buf78), .D(u3_u0_r1_0__FF_INPUT), .Q(u3_u0_r1_0_) );
  DFFPOSX1 DFFPOSX1_989 ( .CLK(clk_i_bF_buf77), .D(u3_u0_r1_1__FF_INPUT), .Q(u3_u0_r1_1_) );
  DFFPOSX1 DFFPOSX1_99 ( .CLK(clk_i_bF_buf25), .D(u0_u0_csc_25__FF_INPUT), .Q(u0_csc0_25_) );
  DFFPOSX1 DFFPOSX1_990 ( .CLK(clk_i_bF_buf76), .D(u3_u0_r1_2__FF_INPUT), .Q(u3_u0_r1_2_) );
  DFFPOSX1 DFFPOSX1_991 ( .CLK(clk_i_bF_buf75), .D(u3_u0_r1_3__FF_INPUT), .Q(u3_u0_r1_3_) );
  DFFPOSX1 DFFPOSX1_992 ( .CLK(clk_i_bF_buf74), .D(u3_u0_r1_4__FF_INPUT), .Q(u3_u0_r1_4_) );
  DFFPOSX1 DFFPOSX1_993 ( .CLK(clk_i_bF_buf73), .D(u3_u0_r1_5__FF_INPUT), .Q(u3_u0_r1_5_) );
  DFFPOSX1 DFFPOSX1_994 ( .CLK(clk_i_bF_buf72), .D(u3_u0_r1_6__FF_INPUT), .Q(u3_u0_r1_6_) );
  DFFPOSX1 DFFPOSX1_995 ( .CLK(clk_i_bF_buf71), .D(u3_u0_r1_7__FF_INPUT), .Q(u3_u0_r1_7_) );
  DFFPOSX1 DFFPOSX1_996 ( .CLK(clk_i_bF_buf70), .D(u3_u0_r1_8__FF_INPUT), .Q(u3_u0_r1_8_) );
  DFFPOSX1 DFFPOSX1_997 ( .CLK(clk_i_bF_buf69), .D(u3_u0_r1_9__FF_INPUT), .Q(u3_u0_r1_9_) );
  DFFPOSX1 DFFPOSX1_998 ( .CLK(clk_i_bF_buf68), .D(u3_u0_r1_10__FF_INPUT), .Q(u3_u0_r1_10_) );
  DFFPOSX1 DFFPOSX1_999 ( .CLK(clk_i_bF_buf67), .D(u3_u0_r1_11__FF_INPUT), .Q(u3_u0_r1_11_) );
  DFFSR DFFSR_1 ( .CLK(clk_i_bF_buf84), .D(u0_lmr_req_FF_INPUT), .Q(lmr_req), .R(u0__abc_49347_n3188_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_10 ( .CLK(clk_i_bF_buf75), .D(u0_spec_req_cs_6__FF_INPUT), .Q(spec_req_cs_6_), .R(u0__abc_49347_n3188_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_100 ( .CLK(clk_i_bF_buf111), .D(u0_csc_mask_r_1__FF_INPUT), .Q(u0_csc_mask_1_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf10) );
  DFFSR DFFSR_101 ( .CLK(clk_i_bF_buf110), .D(u0_csc_mask_r_2__FF_INPUT), .Q(u0_csc_mask_2_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf9) );
  DFFSR DFFSR_102 ( .CLK(clk_i_bF_buf109), .D(u0_csc_mask_r_3__FF_INPUT), .Q(u0_csc_mask_3_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf8) );
  DFFSR DFFSR_103 ( .CLK(clk_i_bF_buf108), .D(u0_csc_mask_r_4__FF_INPUT), .Q(u0_csc_mask_4_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf7) );
  DFFSR DFFSR_104 ( .CLK(clk_i_bF_buf107), .D(u0_csc_mask_r_5__FF_INPUT), .Q(u0_csc_mask_5_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf6) );
  DFFSR DFFSR_105 ( .CLK(clk_i_bF_buf106), .D(u0_csc_mask_r_6__FF_INPUT), .Q(u0_csc_mask_6_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf5) );
  DFFSR DFFSR_106 ( .CLK(clk_i_bF_buf105), .D(u0_csc_mask_r_7__FF_INPUT), .Q(u0_csc_mask_7_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf4) );
  DFFSR DFFSR_107 ( .CLK(clk_i_bF_buf104), .D(u0_csc_mask_r_8__FF_INPUT), .Q(u0_csc_mask_8_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf3) );
  DFFSR DFFSR_108 ( .CLK(clk_i_bF_buf103), .D(u0_csc_mask_r_9__FF_INPUT), .Q(u0_csc_mask_9_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf2) );
  DFFSR DFFSR_109 ( .CLK(clk_i_bF_buf102), .D(u0_csc_mask_r_10__FF_INPUT), .Q(u0_csc_mask_10_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf1) );
  DFFSR DFFSR_11 ( .CLK(clk_i_bF_buf74), .D(u0_spec_req_cs_7__FF_INPUT), .Q(spec_req_cs_7_), .R(u0__abc_49347_n3188_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_110 ( .CLK(clk_i_bF_buf101), .D(u0_csr_r_0__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56315), .R(u0__abc_49347_n3188_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_111 ( .CLK(clk_i_bF_buf100), .D(u0_csr_r_1__FF_INPUT), .Q(fs), .R(u0__abc_49347_n3188_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_112 ( .CLK(clk_i_bF_buf99), .D(u0_csr_r_2__FF_INPUT), .Q(u0_csr_3_), .R(u0__abc_49347_n3188_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_113 ( .CLK(clk_i_bF_buf98), .D(u0_csr_r_3__FF_INPUT), .Q(u0_csr_4_), .R(u0__abc_49347_n3188_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_114 ( .CLK(clk_i_bF_buf97), .D(u0_csr_r_4__FF_INPUT), .Q(u0_csr_5_), .R(u0__abc_49347_n3188_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_115 ( .CLK(clk_i_bF_buf96), .D(u0_csr_r_5__FF_INPUT), .Q(u0_csr_6_), .R(u0__abc_49347_n3188_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_116 ( .CLK(clk_i_bF_buf95), .D(u0_csr_r_6__FF_INPUT), .Q(u0_csr_7_), .R(u0__abc_49347_n3188_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_117 ( .CLK(clk_i_bF_buf94), .D(u0_csr_r_7__FF_INPUT), .Q(ref_int_0_), .R(u0__abc_49347_n3188_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_118 ( .CLK(clk_i_bF_buf93), .D(u0_csr_r_8__FF_INPUT), .Q(ref_int_1_), .R(u0__abc_49347_n3188_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_119 ( .CLK(clk_i_bF_buf92), .D(u0_csr_r_9__FF_INPUT), .Q(ref_int_2_), .R(u0__abc_49347_n3188_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_12 ( .CLK(clk_i_bF_buf73), .D(u0_sp_tms_0__FF_INPUT), .Q(sp_tms_0_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf10) );
  DFFSR DFFSR_120 ( .CLK(clk_i_bF_buf91), .D(u0_csr_r2_0__FF_INPUT), .Q(rfr_ps_val_0_), .R(u0__abc_49347_n3188_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_121 ( .CLK(clk_i_bF_buf90), .D(u0_csr_r2_1__FF_INPUT), .Q(rfr_ps_val_1_), .R(u0__abc_49347_n3188_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_122 ( .CLK(clk_i_bF_buf89), .D(u0_csr_r2_2__FF_INPUT), .Q(rfr_ps_val_2_), .R(u0__abc_49347_n3188_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_123 ( .CLK(clk_i_bF_buf88), .D(u0_csr_r2_3__FF_INPUT), .Q(rfr_ps_val_3_), .R(u0__abc_49347_n3188_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_124 ( .CLK(clk_i_bF_buf87), .D(u0_csr_r2_4__FF_INPUT), .Q(rfr_ps_val_4_), .R(u0__abc_49347_n3188_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_125 ( .CLK(clk_i_bF_buf86), .D(u0_csr_r2_5__FF_INPUT), .Q(rfr_ps_val_5_), .R(u0__abc_49347_n3188_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_126 ( .CLK(clk_i_bF_buf85), .D(u0_csr_r2_6__FF_INPUT), .Q(rfr_ps_val_6_), .R(u0__abc_49347_n3188_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_127 ( .CLK(clk_i_bF_buf84), .D(u0_csr_r2_7__FF_INPUT), .Q(rfr_ps_val_7_), .R(u0__abc_49347_n3188_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_128 ( .CLK(clk_i_bF_buf83), .D(u0_rf_we_FF_INPUT), .Q(u0_rf_we), .R(u0__abc_49347_n3188_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_129 ( .CLK(clk_i_bF_buf13), .D(u0_u0_inited_FF_INPUT), .Q(u0_u0_inited), .R(u0_u0__abc_43300_n325), .S(1'b1) );
  DFFSR DFFSR_13 ( .CLK(clk_i_bF_buf72), .D(u0_sp_tms_1__FF_INPUT), .Q(sp_tms_1_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf9) );
  DFFSR DFFSR_130 ( .CLK(clk_i_bF_buf12), .D(u0_u0_init_req_FF_INPUT), .Q(u0_init_req0), .R(u0_u0__abc_43300_n325), .S(1'b1) );
  DFFSR DFFSR_131 ( .CLK(clk_i_bF_buf11), .D(u0_u0_init_req_we_FF_INPUT_bF_buf1), .Q(u0_u0_init_req_we), .R(u0_u0__abc_43300_n325), .S(1'b1) );
  DFFSR DFFSR_132 ( .CLK(clk_i_bF_buf10), .D(u0_u0_lmr_req_FF_INPUT), .Q(u0_lmr_req0), .R(u0_u0__abc_43300_n325), .S(1'b1) );
  DFFSR DFFSR_133 ( .CLK(clk_i_bF_buf9), .D(u0_u0_lmr_req_we_FF_INPUT_bF_buf1), .Q(u0_u0_lmr_req_we), .R(u0_u0__abc_43300_n325), .S(1'b1) );
  DFFSR DFFSR_134 ( .CLK(clk_i_bF_buf8), .D(u0_u0_rst_r1), .Q(u0_u0_rst_r2), .R(1'b1), .S(u0_u0__abc_43300_n325) );
  DFFSR DFFSR_135 ( .CLK(clk_i_bF_buf7), .D(1'b0), .Q(u0_u0_rst_r1), .R(1'b1), .S(u0_u0__abc_43300_n325) );
  DFFSR DFFSR_136 ( .CLK(clk_i_bF_buf63), .D(u0_u1_inited_FF_INPUT), .Q(u0_u1_inited), .R(u0_u1__abc_43657_n324), .S(1'b1) );
  DFFSR DFFSR_137 ( .CLK(clk_i_bF_buf62), .D(u0_u1_init_req_FF_INPUT), .Q(u0_init_req1), .R(u0_u1__abc_43657_n324), .S(1'b1) );
  DFFSR DFFSR_138 ( .CLK(clk_i_bF_buf61), .D(u0_u1_init_req_we_FF_INPUT_bF_buf7), .Q(u0_u1_init_req_we), .R(u0_u1__abc_43657_n324), .S(1'b1) );
  DFFSR DFFSR_139 ( .CLK(clk_i_bF_buf60), .D(u0_u1_lmr_req_FF_INPUT), .Q(u0_lmr_req1), .R(u0_u1__abc_43657_n324), .S(1'b1) );
  DFFSR DFFSR_14 ( .CLK(clk_i_bF_buf71), .D(u0_sp_tms_2__FF_INPUT), .Q(sp_tms_2_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf8) );
  DFFSR DFFSR_140 ( .CLK(clk_i_bF_buf59), .D(u0_u1_lmr_req_we_FF_INPUT_bF_buf7), .Q(u0_u1_lmr_req_we), .R(u0_u1__abc_43657_n324), .S(1'b1) );
  DFFSR DFFSR_141 ( .CLK(clk_i_bF_buf58), .D(u0_u1_rst_r1), .Q(u0_u1_rst_r2), .R(1'b1), .S(u0_u1__abc_43657_n324) );
  DFFSR DFFSR_142 ( .CLK(clk_i_bF_buf57), .D(1'b0), .Q(u0_u1_rst_r1), .R(1'b1), .S(u0_u1__abc_43657_n324) );
  DFFSR DFFSR_143 ( .CLK(clk_i_bF_buf113), .D(u0_u2_inited_FF_INPUT), .Q(u0_u2_inited), .R(u0_u2__abc_44109_n324), .S(1'b1) );
  DFFSR DFFSR_144 ( .CLK(clk_i_bF_buf112), .D(u0_u2_init_req_FF_INPUT), .Q(u0_init_req2), .R(u0_u2__abc_44109_n324), .S(1'b1) );
  DFFSR DFFSR_145 ( .CLK(clk_i_bF_buf111), .D(u0_u2_init_req_we_FF_INPUT_bF_buf1), .Q(u0_u2_init_req_we), .R(u0_u2__abc_44109_n324), .S(1'b1) );
  DFFSR DFFSR_146 ( .CLK(clk_i_bF_buf110), .D(u0_u2_lmr_req_FF_INPUT), .Q(u0_lmr_req2), .R(u0_u2__abc_44109_n324), .S(1'b1) );
  DFFSR DFFSR_147 ( .CLK(clk_i_bF_buf109), .D(u0_u2_lmr_req_we_FF_INPUT_bF_buf1), .Q(u0_u2_lmr_req_we), .R(u0_u2__abc_44109_n324), .S(1'b1) );
  DFFSR DFFSR_148 ( .CLK(clk_i_bF_buf108), .D(u0_u2_rst_r1), .Q(u0_u2_rst_r2), .R(1'b1), .S(u0_u2__abc_44109_n324) );
  DFFSR DFFSR_149 ( .CLK(clk_i_bF_buf107), .D(1'b0), .Q(u0_u2_rst_r1), .R(1'b1), .S(u0_u2__abc_44109_n324) );
  DFFSR DFFSR_15 ( .CLK(clk_i_bF_buf70), .D(u0_sp_tms_3__FF_INPUT), .Q(sp_tms_3_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf7) );
  DFFSR DFFSR_150 ( .CLK(clk_i_bF_buf37), .D(u0_u3_inited_FF_INPUT), .Q(u0_u3_inited), .R(u0_u3__abc_44466_n328), .S(1'b1) );
  DFFSR DFFSR_151 ( .CLK(clk_i_bF_buf36), .D(u0_u3_init_req_FF_INPUT), .Q(u0_init_req3), .R(u0_u3__abc_44466_n328), .S(1'b1) );
  DFFSR DFFSR_152 ( .CLK(clk_i_bF_buf35), .D(u0_u3_init_req_we_FF_INPUT_bF_buf3), .Q(u0_u3_init_req_we), .R(u0_u3__abc_44466_n328), .S(1'b1) );
  DFFSR DFFSR_153 ( .CLK(clk_i_bF_buf34), .D(u0_u3_lmr_req_FF_INPUT), .Q(u0_lmr_req3), .R(u0_u3__abc_44466_n328), .S(1'b1) );
  DFFSR DFFSR_154 ( .CLK(clk_i_bF_buf33), .D(u0_u3_lmr_req_we_FF_INPUT_bF_buf1), .Q(u0_u3_lmr_req_we), .R(u0_u3__abc_44466_n328), .S(1'b1) );
  DFFSR DFFSR_155 ( .CLK(clk_i_bF_buf32), .D(u0_u3_rst_r1), .Q(u0_u3_rst_r2), .R(1'b1), .S(u0_u3__abc_44466_n328) );
  DFFSR DFFSR_156 ( .CLK(clk_i_bF_buf31), .D(1'b0), .Q(u0_u3_rst_r1), .R(1'b1), .S(u0_u3__abc_44466_n328) );
  DFFSR DFFSR_157 ( .CLK(clk_i_bF_buf87), .D(u0_u4_inited_FF_INPUT), .Q(u0_u4_inited), .R(u0_u4__abc_44844_n324), .S(1'b1) );
  DFFSR DFFSR_158 ( .CLK(clk_i_bF_buf86), .D(u0_u4_init_req_FF_INPUT), .Q(u0_init_req4), .R(u0_u4__abc_44844_n324), .S(1'b1) );
  DFFSR DFFSR_159 ( .CLK(clk_i_bF_buf85), .D(u0_u4_init_req_we_FF_INPUT_bF_buf7), .Q(u0_u4_init_req_we), .R(u0_u4__abc_44844_n324), .S(1'b1) );
  DFFSR DFFSR_16 ( .CLK(clk_i_bF_buf69), .D(u0_sp_tms_4__FF_INPUT), .Q(sp_tms_4_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf6) );
  DFFSR DFFSR_160 ( .CLK(clk_i_bF_buf84), .D(u0_u4_lmr_req_FF_INPUT), .Q(u0_lmr_req4), .R(u0_u4__abc_44844_n324), .S(1'b1) );
  DFFSR DFFSR_161 ( .CLK(clk_i_bF_buf83), .D(u0_u4_lmr_req_we_FF_INPUT_bF_buf7), .Q(u0_u4_lmr_req_we), .R(u0_u4__abc_44844_n324), .S(1'b1) );
  DFFSR DFFSR_162 ( .CLK(clk_i_bF_buf82), .D(u0_u4_rst_r1), .Q(u0_u4_rst_r2), .R(1'b1), .S(u0_u4__abc_44844_n324) );
  DFFSR DFFSR_163 ( .CLK(clk_i_bF_buf81), .D(1'b0), .Q(u0_u4_rst_r1), .R(1'b1), .S(u0_u4__abc_44844_n324) );
  DFFSR DFFSR_164 ( .CLK(clk_i_bF_buf11), .D(u0_u5_inited_FF_INPUT), .Q(u0_u5_inited), .R(u0_u5__abc_45296_n325), .S(1'b1) );
  DFFSR DFFSR_165 ( .CLK(clk_i_bF_buf10), .D(u0_u5_init_req_FF_INPUT), .Q(u0_init_req5), .R(u0_u5__abc_45296_n325), .S(1'b1) );
  DFFSR DFFSR_166 ( .CLK(clk_i_bF_buf9), .D(u0_u5_init_req_we_FF_INPUT_bF_buf7), .Q(u0_u5_init_req_we), .R(u0_u5__abc_45296_n325), .S(1'b1) );
  DFFSR DFFSR_167 ( .CLK(clk_i_bF_buf8), .D(u0_u5_lmr_req_FF_INPUT), .Q(u0_lmr_req5), .R(u0_u5__abc_45296_n325), .S(1'b1) );
  DFFSR DFFSR_168 ( .CLK(clk_i_bF_buf7), .D(u0_u5_lmr_req_we_FF_INPUT_bF_buf7), .Q(u0_u5_lmr_req_we), .R(u0_u5__abc_45296_n325), .S(1'b1) );
  DFFSR DFFSR_169 ( .CLK(clk_i_bF_buf6), .D(u0_u5_rst_r1), .Q(u0_u5_rst_r2), .R(1'b1), .S(u0_u5__abc_45296_n325) );
  DFFSR DFFSR_17 ( .CLK(clk_i_bF_buf68), .D(u0_sp_tms_5__FF_INPUT), .Q(sp_tms_5_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf5) );
  DFFSR DFFSR_170 ( .CLK(clk_i_bF_buf5), .D(1'b0), .Q(u0_u5_rst_r1), .R(1'b1), .S(u0_u5__abc_45296_n325) );
  DFFSR DFFSR_171 ( .CLK(clk_i_bF_buf116), .D(u2_u0_bank3_open_FF_INPUT), .Q(u2_u0_bank3_open), .R(u2_u0__abc_47660_n305), .S(1'b1) );
  DFFSR DFFSR_172 ( .CLK(clk_i_bF_buf115), .D(u2_u0_bank2_open_FF_INPUT), .Q(u2_u0_bank2_open), .R(u2_u0__abc_47660_n305), .S(1'b1) );
  DFFSR DFFSR_173 ( .CLK(clk_i_bF_buf114), .D(u2_u0_bank1_open_FF_INPUT), .Q(u2_u0_bank1_open), .R(u2_u0__abc_47660_n305), .S(1'b1) );
  DFFSR DFFSR_174 ( .CLK(clk_i_bF_buf113), .D(u2_u0_bank0_open_FF_INPUT), .Q(u2_u0_bank0_open), .R(u2_u0__abc_47660_n305), .S(1'b1) );
  DFFSR DFFSR_175 ( .CLK(clk_i_bF_buf60), .D(u2_u1_bank3_open_FF_INPUT), .Q(u2_u1_bank3_open), .R(u2_u1__abc_47660_n305), .S(1'b1) );
  DFFSR DFFSR_176 ( .CLK(clk_i_bF_buf59), .D(u2_u1_bank2_open_FF_INPUT), .Q(u2_u1_bank2_open), .R(u2_u1__abc_47660_n305), .S(1'b1) );
  DFFSR DFFSR_177 ( .CLK(clk_i_bF_buf58), .D(u2_u1_bank1_open_FF_INPUT), .Q(u2_u1_bank1_open), .R(u2_u1__abc_47660_n305), .S(1'b1) );
  DFFSR DFFSR_178 ( .CLK(clk_i_bF_buf57), .D(u2_u1_bank0_open_FF_INPUT), .Q(u2_u1_bank0_open), .R(u2_u1__abc_47660_n305), .S(1'b1) );
  DFFSR DFFSR_179 ( .CLK(clk_i_bF_buf4), .D(u2_u2_bank3_open_FF_INPUT), .Q(u2_u2_bank3_open), .R(u2_u2__abc_47660_n305), .S(1'b1) );
  DFFSR DFFSR_18 ( .CLK(clk_i_bF_buf67), .D(u0_sp_tms_6__FF_INPUT), .Q(sp_tms_6_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf4) );
  DFFSR DFFSR_180 ( .CLK(clk_i_bF_buf3), .D(u2_u2_bank2_open_FF_INPUT), .Q(u2_u2_bank2_open), .R(u2_u2__abc_47660_n305), .S(1'b1) );
  DFFSR DFFSR_181 ( .CLK(clk_i_bF_buf2), .D(u2_u2_bank1_open_FF_INPUT), .Q(u2_u2_bank1_open), .R(u2_u2__abc_47660_n305), .S(1'b1) );
  DFFSR DFFSR_182 ( .CLK(clk_i_bF_buf1), .D(u2_u2_bank0_open_FF_INPUT), .Q(u2_u2_bank0_open), .R(u2_u2__abc_47660_n305), .S(1'b1) );
  DFFSR DFFSR_183 ( .CLK(clk_i_bF_buf74), .D(u2_u3_bank3_open_FF_INPUT), .Q(u2_u3_bank3_open), .R(u2_u3__abc_47660_n305), .S(1'b1) );
  DFFSR DFFSR_184 ( .CLK(clk_i_bF_buf73), .D(u2_u3_bank2_open_FF_INPUT), .Q(u2_u3_bank2_open), .R(u2_u3__abc_47660_n305), .S(1'b1) );
  DFFSR DFFSR_185 ( .CLK(clk_i_bF_buf72), .D(u2_u3_bank1_open_FF_INPUT), .Q(u2_u3_bank1_open), .R(u2_u3__abc_47660_n305), .S(1'b1) );
  DFFSR DFFSR_186 ( .CLK(clk_i_bF_buf71), .D(u2_u3_bank0_open_FF_INPUT), .Q(u2_u3_bank0_open), .R(u2_u3__abc_47660_n305), .S(1'b1) );
  DFFSR DFFSR_187 ( .CLK(clk_i_bF_buf18), .D(u2_u4_bank3_open_FF_INPUT), .Q(u2_u4_bank3_open), .R(u2_u4__abc_47660_n305), .S(1'b1) );
  DFFSR DFFSR_188 ( .CLK(clk_i_bF_buf17), .D(u2_u4_bank2_open_FF_INPUT), .Q(u2_u4_bank2_open), .R(u2_u4__abc_47660_n305), .S(1'b1) );
  DFFSR DFFSR_189 ( .CLK(clk_i_bF_buf16), .D(u2_u4_bank1_open_FF_INPUT), .Q(u2_u4_bank1_open), .R(u2_u4__abc_47660_n305), .S(1'b1) );
  DFFSR DFFSR_19 ( .CLK(clk_i_bF_buf66), .D(u0_sp_tms_7__FF_INPUT), .Q(sp_tms_7_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf3) );
  DFFSR DFFSR_190 ( .CLK(clk_i_bF_buf15), .D(u2_u4_bank0_open_FF_INPUT), .Q(u2_u4_bank0_open), .R(u2_u4__abc_47660_n305), .S(1'b1) );
  DFFSR DFFSR_191 ( .CLK(clk_i_bF_buf88), .D(u2_u5_bank3_open_FF_INPUT), .Q(u2_u5_bank3_open), .R(u2_u5__abc_47660_n305), .S(1'b1) );
  DFFSR DFFSR_192 ( .CLK(clk_i_bF_buf87), .D(u2_u5_bank2_open_FF_INPUT), .Q(u2_u5_bank2_open), .R(u2_u5__abc_47660_n305), .S(1'b1) );
  DFFSR DFFSR_193 ( .CLK(clk_i_bF_buf86), .D(u2_u5_bank1_open_FF_INPUT), .Q(u2_u5_bank1_open), .R(u2_u5__abc_47660_n305), .S(1'b1) );
  DFFSR DFFSR_194 ( .CLK(clk_i_bF_buf85), .D(u2_u5_bank0_open_FF_INPUT), .Q(u2_u5_bank0_open), .R(u2_u5__abc_47660_n305), .S(1'b1) );
  DFFSR DFFSR_195 ( .CLK(clk_i_bF_buf6), .D(u3_u0_wr_adr_0__FF_INPUT), .Q(u3_u0_wr_adr_0_), .R(1'b1), .S(u3_u0__abc_48231_n514) );
  DFFSR DFFSR_196 ( .CLK(clk_i_bF_buf5), .D(u3_u0_wr_adr_1__FF_INPUT), .Q(u3_u0_wr_adr_1_), .R(u3_u0__abc_48231_n514), .S(1'b1) );
  DFFSR DFFSR_197 ( .CLK(clk_i_bF_buf4), .D(u3_u0_wr_adr_2__FF_INPUT), .Q(u3_u0_wr_adr_2_), .R(u3_u0__abc_48231_n514), .S(1'b1) );
  DFFSR DFFSR_198 ( .CLK(clk_i_bF_buf3), .D(u3_u0_wr_adr_3__FF_INPUT), .Q(u3_u0_wr_adr_3_), .R(u3_u0__abc_48231_n514), .S(1'b1) );
  DFFSR DFFSR_199 ( .CLK(clk_i_bF_buf2), .D(u3_u0_rd_adr_0__FF_INPUT), .Q(u3_u0_rd_adr_0_), .R(1'b1), .S(u3_u0__abc_48231_n514) );
  DFFSR DFFSR_2 ( .CLK(clk_i_bF_buf83), .D(u0_init_req_FF_INPUT), .Q(init_req), .R(u0__abc_49347_n3188_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_20 ( .CLK(clk_i_bF_buf65), .D(u0_sp_tms_8__FF_INPUT), .Q(sp_tms_8_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf2) );
  DFFSR DFFSR_200 ( .CLK(clk_i_bF_buf1), .D(u3_u0_rd_adr_1__FF_INPUT), .Q(u3_u0_rd_adr_1_), .R(u3_u0__abc_48231_n514), .S(1'b1) );
  DFFSR DFFSR_201 ( .CLK(clk_i_bF_buf0), .D(u3_u0_rd_adr_2__FF_INPUT), .Q(u3_u0_rd_adr_2_), .R(u3_u0__abc_48231_n514), .S(1'b1) );
  DFFSR DFFSR_202 ( .CLK(clk_i_bF_buf125), .D(u3_u0_rd_adr_3__FF_INPUT), .Q(u3_u0_rd_adr_3_), .R(u3_u0__abc_48231_n514), .S(1'b1) );
  DFFSR DFFSR_203 ( .CLK(clk_i_bF_buf123), .D(u4_rfr_req_FF_INPUT), .Q(rfr_req), .R(u4__abc_49152_n191_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_204 ( .CLK(clk_i_bF_buf122), .D(u4_rfr_cnt_0__FF_INPUT), .Q(u4_rfr_cnt_0_), .R(u4__abc_49152_n191_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_205 ( .CLK(clk_i_bF_buf121), .D(u4_rfr_cnt_1__FF_INPUT), .Q(u4_rfr_cnt_1_), .R(u4__abc_49152_n191_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_206 ( .CLK(clk_i_bF_buf120), .D(u4_rfr_cnt_2__FF_INPUT), .Q(u4_rfr_cnt_2_), .R(u4__abc_49152_n191_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_207 ( .CLK(clk_i_bF_buf119), .D(u4_rfr_cnt_3__FF_INPUT), .Q(u4_rfr_cnt_3_), .R(u4__abc_49152_n191_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_208 ( .CLK(clk_i_bF_buf118), .D(u4_rfr_cnt_4__FF_INPUT), .Q(u4_rfr_cnt_4_), .R(u4__abc_49152_n191_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_209 ( .CLK(clk_i_bF_buf117), .D(u4_rfr_cnt_5__FF_INPUT), .Q(u4_rfr_cnt_5_), .R(u4__abc_49152_n191_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_21 ( .CLK(clk_i_bF_buf64), .D(u0_sp_tms_9__FF_INPUT), .Q(sp_tms_9_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf1) );
  DFFSR DFFSR_210 ( .CLK(clk_i_bF_buf116), .D(u4_rfr_cnt_6__FF_INPUT), .Q(u4_rfr_cnt_6_), .R(u4__abc_49152_n191_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_211 ( .CLK(clk_i_bF_buf115), .D(u4_rfr_cnt_7__FF_INPUT), .Q(u4_rfr_cnt_7_), .R(u4__abc_49152_n191_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_212 ( .CLK(clk_i_bF_buf114), .D(u4_ps_cnt_clr), .Q(u4_rfr_ce), .R(u4__abc_49152_n191_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_213 ( .CLK(clk_i_bF_buf113), .D(u4_rfr_early_FF_INPUT), .Q(u4_rfr_early), .R(u4__abc_49152_n191_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_214 ( .CLK(clk_i_bF_buf112), .D(u4_ps_cnt_0__FF_INPUT), .Q(u4_ps_cnt_0_), .R(u4__abc_49152_n191_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_215 ( .CLK(clk_i_bF_buf111), .D(u4_ps_cnt_1__FF_INPUT), .Q(u4_ps_cnt_1_), .R(u4__abc_49152_n191_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_216 ( .CLK(clk_i_bF_buf110), .D(u4_ps_cnt_2__FF_INPUT), .Q(u4_ps_cnt_2_), .R(u4__abc_49152_n191_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_217 ( .CLK(clk_i_bF_buf109), .D(u4_ps_cnt_3__FF_INPUT), .Q(u4_ps_cnt_3_), .R(u4__abc_49152_n191_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_218 ( .CLK(clk_i_bF_buf108), .D(u4_ps_cnt_4__FF_INPUT), .Q(u4_ps_cnt_4_), .R(u4__abc_49152_n191_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_219 ( .CLK(clk_i_bF_buf107), .D(u4_ps_cnt_5__FF_INPUT), .Q(u4_ps_cnt_5_), .R(u4__abc_49152_n191_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_22 ( .CLK(clk_i_bF_buf63), .D(u0_sp_tms_10__FF_INPUT), .Q(sp_tms_10_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf0) );
  DFFSR DFFSR_220 ( .CLK(clk_i_bF_buf106), .D(u4_ps_cnt_6__FF_INPUT), .Q(u4_ps_cnt_6_), .R(u4__abc_49152_n191_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_221 ( .CLK(clk_i_bF_buf105), .D(u4_ps_cnt_7__FF_INPUT), .Q(u4_ps_cnt_7_), .R(u4__abc_49152_n191_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_222 ( .CLK(clk_i_bF_buf104), .D(u4_rfr_en_FF_INPUT), .Q(u4_rfr_en), .R(u4__abc_49152_n191_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_223 ( .CLK(clk_i_bF_buf60), .D(u5__abc_41027_n1845), .Q(u5_state_0_), .R(u5__abc_54027_n1575_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_224 ( .CLK(clk_i_bF_buf59), .D(u5__abc_41027_n1846), .Q(u5_state_1_), .R(u5__abc_54027_n1575_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_225 ( .CLK(clk_i_bF_buf58), .D(u5__abc_41027_n1847), .Q(u5_state_2_), .R(u5__abc_54027_n1575_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_226 ( .CLK(clk_i_bF_buf57), .D(u5__abc_41027_n1848), .Q(u5_state_3_), .R(u5__abc_54027_n1575_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_227 ( .CLK(clk_i_bF_buf56), .D(u5__abc_41027_n1849), .Q(u5_state_4_), .R(u5__abc_54027_n1575_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_228 ( .CLK(clk_i_bF_buf55), .D(u5__abc_41027_n1850), .Q(u5_state_5_), .R(u5__abc_54027_n1575_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_229 ( .CLK(clk_i_bF_buf54), .D(u5__abc_41027_n1851), .Q(u5_state_6_), .R(u5__abc_54027_n1575_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_23 ( .CLK(clk_i_bF_buf62), .D(u0_sp_tms_11__FF_INPUT), .Q(sp_tms_11_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf10) );
  DFFSR DFFSR_230 ( .CLK(clk_i_bF_buf53), .D(u5_wb_stb_first_FF_INPUT), .Q(u5_wb_stb_first), .R(u5__abc_54027_n1575_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_231 ( .CLK(clk_i_bF_buf52), .D(dv), .Q(u5_dv_r), .R(u5__abc_54027_n1575_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_232 ( .CLK(clk_i_bF_buf51), .D(u5_ap_en_FF_INPUT), .Q(u5_ap_en), .R(u5__abc_54027_n1575_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_233 ( .CLK(clk_i_bF_buf50), .D(u5_timer_is_zero), .Q(u5_tmr_done), .R(u5__abc_54027_n1575_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_234 ( .CLK(clk_i_bF_buf49), .D(u5_timer_0__FF_INPUT), .Q(u5_timer_0_), .R(u5__abc_54027_n1575_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_235 ( .CLK(clk_i_bF_buf48), .D(u5_timer_1__FF_INPUT), .Q(u5_timer_1_), .R(1'b1), .S(u5__abc_54027_n1575_bF_buf1) );
  DFFSR DFFSR_236 ( .CLK(clk_i_bF_buf47), .D(u5_timer_2__FF_INPUT), .Q(u5_timer_2_), .R(u5__abc_54027_n1575_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_237 ( .CLK(clk_i_bF_buf46), .D(u5_timer_3__FF_INPUT), .Q(u5_timer_3_), .R(1'b1), .S(u5__abc_54027_n1575_bF_buf6) );
  DFFSR DFFSR_238 ( .CLK(clk_i_bF_buf45), .D(u5_timer_4__FF_INPUT), .Q(u5_timer_4_), .R(1'b1), .S(u5__abc_54027_n1575_bF_buf5) );
  DFFSR DFFSR_239 ( .CLK(clk_i_bF_buf44), .D(u5_timer_5__FF_INPUT), .Q(u5_timer_5_), .R(1'b1), .S(u5__abc_54027_n1575_bF_buf4) );
  DFFSR DFFSR_24 ( .CLK(clk_i_bF_buf61), .D(u0_sp_tms_12__FF_INPUT), .Q(sp_tms_12_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf9) );
  DFFSR DFFSR_240 ( .CLK(clk_i_bF_buf43), .D(u5_timer_6__FF_INPUT), .Q(u5_timer_6_), .R(1'b1), .S(u5__abc_54027_n1575_bF_buf3) );
  DFFSR DFFSR_241 ( .CLK(clk_i_bF_buf42), .D(u5_timer_7__FF_INPUT), .Q(u5_timer_7_), .R(1'b1), .S(u5__abc_54027_n1575_bF_buf2) );
  DFFSR DFFSR_242 ( .CLK(clk_i_bF_buf41), .D(u5_tmr2_done_FF_INPUT), .Q(u5_tmr2_done), .R(u5__abc_54027_n1575_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_243 ( .CLK(clk_i_bF_buf40), .D(u5_susp_sel_r_FF_INPUT), .Q(susp_sel), .R(u5__abc_54027_n1575_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_244 ( .CLK(clk_i_bF_buf39), .D(u5_rfr_ack_d), .Q(rfr_ack), .R(u5__abc_54027_n1575_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_245 ( .CLK(clk_i_bF_buf38), .D(u5_suspended_d), .Q(_auto_iopadmap_cc_313_execute_56354), .R(u5__abc_54027_n1575_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_246 ( .CLK(clk_i_bF_buf37), .D(resume_req_i), .Q(u5_resume_req_r), .R(u5__abc_54027_n1575_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_247 ( .CLK(clk_i_bF_buf36), .D(susp_req_i), .Q(u5_susp_req_r), .R(u5__abc_54027_n1575_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_248 ( .CLK(clk_i_bF_buf35), .D(u5_ack_cnt_0__FF_INPUT), .Q(u5_ack_cnt_0_), .R(u5__abc_54027_n1575_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_249 ( .CLK(clk_i_bF_buf34), .D(u5_ack_cnt_1__FF_INPUT), .Q(u5_ack_cnt_1_), .R(u5__abc_54027_n1575_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_25 ( .CLK(clk_i_bF_buf60), .D(u0_sp_tms_13__FF_INPUT), .Q(sp_tms_13_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf8) );
  DFFSR DFFSR_250 ( .CLK(clk_i_bF_buf33), .D(u5_ack_cnt_2__FF_INPUT), .Q(u5_ack_cnt_2_), .R(u5__abc_54027_n1575_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_251 ( .CLK(clk_i_bF_buf32), .D(u5_ack_cnt_3__FF_INPUT), .Q(u5_ack_cnt_3_), .R(u5__abc_54027_n1575_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_252 ( .CLK(clk_i_bF_buf31), .D(u5_no_wb_cycle_FF_INPUT), .Q(u5_no_wb_cycle), .R(u5__abc_54027_n1575_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_253 ( .CLK(clk_i_bF_buf30), .D(u5_wb_cycle_FF_INPUT), .Q(u5_wb_cycle), .R(u5__abc_54027_n1575_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_254 ( .CLK(clk_i_bF_buf29), .D(u5_wr_cycle_FF_INPUT), .Q(u1_wr_cycle), .R(u5__abc_54027_n1575_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_255 ( .CLK(clk_i_bF_buf28), .D(u5_lookup_ready2_FF_INPUT), .Q(u5_lookup_ready2), .R(u5__abc_54027_n1575_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_256 ( .CLK(clk_i_bF_buf27), .D(u5_lookup_ready1_FF_INPUT), .Q(u5_lookup_ready1), .R(u5__abc_54027_n1575_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_257 ( .CLK(clk_i_bF_buf26), .D(u5_data_oe_FF_INPUT), .Q(data_oe), .R(u5__abc_54027_n1575_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_258 ( .CLK(clk_i_bF_buf25), .D(u5_data_oe_r), .Q(u5_data_oe_r2), .R(u5__abc_54027_n1575_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_259 ( .CLK(clk_i_bF_buf24), .D(u5_data_oe_d), .Q(u5_data_oe_r), .R(u5__abc_54027_n1575_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_26 ( .CLK(clk_i_bF_buf59), .D(u0_sp_tms_14__FF_INPUT), .Q(sp_tms_14_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf7) );
  DFFSR DFFSR_260 ( .CLK(clk_i_bF_buf23), .D(u5_oe__FF_INPUT), .Q(oe_), .R(1'b1), .S(u5__abc_54027_n1575_bF_buf4) );
  DFFSR DFFSR_261 ( .CLK(clk_i_bF_buf22), .D(u5_cmd_asserted2_FF_INPUT), .Q(u5_cmd_asserted2), .R(u5__abc_54027_n1575_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_262 ( .CLK(clk_i_bF_buf21), .D(u5_cmd_asserted_FF_INPUT), .Q(u5_cmd_asserted), .R(u5__abc_54027_n1575_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_263 ( .CLK(clk_i_bF_buf20), .D(u5_cmd_r_0_), .Q(u5_cmd_del_0_), .R(1'b1), .S(u5__abc_54027_n1575_bF_buf1) );
  DFFSR DFFSR_264 ( .CLK(clk_i_bF_buf19), .D(u5_cmd_r_1_), .Q(u5_cmd_del_1_), .R(1'b1), .S(u5__abc_54027_n1575_bF_buf0) );
  DFFSR DFFSR_265 ( .CLK(clk_i_bF_buf18), .D(u5_cmd_r_2_), .Q(u5_cmd_del_2_), .R(1'b1), .S(u5__abc_54027_n1575_bF_buf6) );
  DFFSR DFFSR_266 ( .CLK(clk_i_bF_buf17), .D(u5_cmd_r_3_), .Q(u5_cmd_del_3_), .R(u5__abc_54027_n1575_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_267 ( .CLK(clk_i_bF_buf16), .D(u5_cmd_0_), .Q(u5_cmd_r_0_), .R(1'b1), .S(u5__abc_54027_n1575_bF_buf4) );
  DFFSR DFFSR_268 ( .CLK(clk_i_bF_buf15), .D(u5_cmd_1_), .Q(u5_cmd_r_1_), .R(1'b1), .S(u5__abc_54027_n1575_bF_buf3) );
  DFFSR DFFSR_269 ( .CLK(clk_i_bF_buf14), .D(u5_cmd_2_), .Q(u5_cmd_r_2_), .R(1'b1), .S(u5__abc_54027_n1575_bF_buf2) );
  DFFSR DFFSR_27 ( .CLK(clk_i_bF_buf58), .D(u0_sp_tms_15__FF_INPUT), .Q(sp_tms_15_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf6) );
  DFFSR DFFSR_270 ( .CLK(clk_i_bF_buf13), .D(u5_cmd_3_), .Q(u5_cmd_r_3_), .R(u5__abc_54027_n1575_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_271 ( .CLK(clk_i_bF_buf12), .D(mem_ack), .Q(u5_mem_ack_r), .R(u5__abc_54027_n1575_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_272 ( .CLK(clk_i_bF_buf11), .D(u5_mc_adv_r_FF_INPUT), .Q(u5_mc_adv_r), .R(u5__abc_54027_n1575_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_273 ( .CLK(clk_i_bF_buf10), .D(u5_mc_adv_r1_FF_INPUT), .Q(u5_mc_adv_r1), .R(u5__abc_54027_n1575_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_274 ( .CLK(clk_i_bF_buf9), .D(u5_mc_le_FF_INPUT), .Q(u5_mc_le), .R(u5__abc_54027_n1573), .S(1'b1) );
  DFFSR DFFSR_275 ( .CLK(clk_i_bF_buf8), .D(u5_mc_c_oe_d), .Q(mc_c_oe_d), .R(u5__abc_54027_n1575_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_276 ( .CLK(clk_i_bF_buf7), .D(u5_rsts1), .Q(u5_rsts), .R(1'b1), .S(u5__abc_54027_n1575_bF_buf3) );
  DFFSR DFFSR_277 ( .CLK(mc_clk_i_bF_buf10), .D(1'b0), .Q(u5_rsts1), .R(1'b1), .S(u5__abc_54027_n1575_bF_buf2) );
  DFFSR DFFSR_278 ( .CLK(clk_i_bF_buf100), .D(u6_wb_err_FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56391), .R(u6__abc_56056_n167), .S(1'b1) );
  DFFSR DFFSR_279 ( .CLK(clk_i_bF_buf99), .D(u6_wb_ack_o_FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56356), .R(u6__abc_56056_n167), .S(1'b1) );
  DFFSR DFFSR_28 ( .CLK(clk_i_bF_buf57), .D(u0_sp_tms_16__FF_INPUT), .Q(sp_tms_16_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf5) );
  DFFSR DFFSR_280 ( .CLK(clk_i_bF_buf98), .D(u6_wr_hold_FF_INPUT), .Q(u1_wr_hold), .R(u6__abc_56056_n167), .S(1'b1) );
  DFFSR DFFSR_281 ( .CLK(clk_i_bF_buf97), .D(u5_wb_first), .Q(u6_wb_first_r), .R(u6__abc_56056_n167), .S(1'b1) );
  DFFSR DFFSR_282 ( .CLK(clk_i_bF_buf96), .D(u6_write_go_r_FF_INPUT), .Q(u6_write_go_r), .R(u6__abc_56056_n167), .S(1'b1) );
  DFFSR DFFSR_283 ( .CLK(clk_i_bF_buf95), .D(u6_write_go_r1_FF_INPUT), .Q(u6_write_go_r1), .R(u6__abc_56056_n167), .S(1'b1) );
  DFFSR DFFSR_284 ( .CLK(clk_i_bF_buf94), .D(u6_read_go_r_FF_INPUT), .Q(u6_read_go_r), .R(u6__abc_56056_n167), .S(1'b1) );
  DFFSR DFFSR_285 ( .CLK(clk_i_bF_buf93), .D(u6_read_go_r1_FF_INPUT), .Q(u6_read_go_r1), .R(u6__abc_56056_n167), .S(1'b1) );
  DFFSR DFFSR_286 ( .CLK(clk_i_bF_buf92), .D(u6_rmw_r_FF_INPUT), .Q(u6_rmw_r), .R(u6__abc_56056_n167), .S(1'b1) );
  DFFSR DFFSR_287 ( .CLK(clk_i_bF_buf91), .D(u6_rmw_en_FF_INPUT), .Q(u6_rmw_en), .R(u6__abc_56056_n167), .S(1'b1) );
  DFFSR DFFSR_288 ( .CLK(mc_clk_i_bF_buf7), .D(u7_mc_cs__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56255_7_), .R(1'b1), .S(u7__abc_47535_n99) );
  DFFSR DFFSR_289 ( .CLK(mc_clk_i_bF_buf6), .D(u7_mc_cs__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56255_6_), .R(1'b1), .S(u7__abc_47535_n99) );
  DFFSR DFFSR_29 ( .CLK(clk_i_bF_buf56), .D(u0_sp_tms_17__FF_INPUT), .Q(sp_tms_17_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf4) );
  DFFSR DFFSR_290 ( .CLK(mc_clk_i_bF_buf5), .D(u7_mc_cs__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56255_5_), .R(1'b1), .S(u7__abc_47535_n99) );
  DFFSR DFFSR_291 ( .CLK(mc_clk_i_bF_buf4), .D(u7_mc_cs__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56255_4_), .R(1'b1), .S(u7__abc_47535_n99) );
  DFFSR DFFSR_292 ( .CLK(mc_clk_i_bF_buf3), .D(u7_mc_cs__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56255_3_), .R(1'b1), .S(u7__abc_47535_n99) );
  DFFSR DFFSR_293 ( .CLK(mc_clk_i_bF_buf2), .D(u7_mc_cs__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56255_2_), .R(1'b1), .S(u7__abc_47535_n99) );
  DFFSR DFFSR_294 ( .CLK(mc_clk_i_bF_buf1), .D(u7_mc_cs__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56255_1_), .R(1'b1), .S(u7__abc_47535_n99) );
  DFFSR DFFSR_295 ( .CLK(mc_clk_i_bF_buf0), .D(u7_mc_cs__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56255_0_), .R(1'b1), .S(u7__abc_47535_n99) );
  DFFSR DFFSR_296 ( .CLK(mc_clk_i_bF_buf10), .D(u7_mc_oe__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56309), .R(1'b1), .S(u7__abc_47535_n99) );
  DFFSR DFFSR_297 ( .CLK(mc_clk_i_bF_buf9), .D(u7_mc_data_oe_FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_56297), .R(u7__abc_47535_n99), .S(1'b1) );
  DFFSR DFFSR_3 ( .CLK(clk_i_bF_buf82), .D(u0_sreq_cs_le_FF_INPUT), .Q(u0_sreq_cs_le), .R(u0__abc_49347_n3188_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_30 ( .CLK(clk_i_bF_buf55), .D(u0_sp_tms_18__FF_INPUT), .Q(sp_tms_18_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf3) );
  DFFSR DFFSR_31 ( .CLK(clk_i_bF_buf54), .D(u0_sp_tms_19__FF_INPUT), .Q(sp_tms_19_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf2) );
  DFFSR DFFSR_32 ( .CLK(clk_i_bF_buf53), .D(u0_sp_tms_20__FF_INPUT), .Q(sp_tms_20_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf1) );
  DFFSR DFFSR_33 ( .CLK(clk_i_bF_buf52), .D(u0_sp_tms_21__FF_INPUT), .Q(sp_tms_21_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf0) );
  DFFSR DFFSR_34 ( .CLK(clk_i_bF_buf51), .D(u0_sp_tms_22__FF_INPUT), .Q(sp_tms_22_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf10) );
  DFFSR DFFSR_35 ( .CLK(clk_i_bF_buf50), .D(u0_sp_tms_23__FF_INPUT), .Q(sp_tms_23_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf9) );
  DFFSR DFFSR_36 ( .CLK(clk_i_bF_buf49), .D(u0_sp_tms_24__FF_INPUT), .Q(sp_tms_24_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf8) );
  DFFSR DFFSR_37 ( .CLK(clk_i_bF_buf48), .D(u0_sp_tms_25__FF_INPUT), .Q(sp_tms_25_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf7) );
  DFFSR DFFSR_38 ( .CLK(clk_i_bF_buf47), .D(u0_sp_tms_26__FF_INPUT), .Q(sp_tms_26_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf6) );
  DFFSR DFFSR_39 ( .CLK(clk_i_bF_buf46), .D(u0_sp_tms_27__FF_INPUT), .Q(sp_tms_27_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf5) );
  DFFSR DFFSR_4 ( .CLK(clk_i_bF_buf81), .D(u0_spec_req_cs_0__FF_INPUT), .Q(spec_req_cs_0_), .R(u0__abc_49347_n3188_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_40 ( .CLK(clk_i_bF_buf45), .D(u0_sp_csc_1__FF_INPUT), .Q(sp_csc_1_), .R(u0__abc_49347_n3188_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_41 ( .CLK(clk_i_bF_buf44), .D(u0_sp_csc_2__FF_INPUT), .Q(sp_csc_2_), .R(u0__abc_49347_n3188_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_42 ( .CLK(clk_i_bF_buf43), .D(u0_sp_csc_3__FF_INPUT), .Q(sp_csc_3_), .R(u0__abc_49347_n3188_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_43 ( .CLK(clk_i_bF_buf42), .D(u0_sp_csc_4__FF_INPUT), .Q(sp_csc_4_), .R(u0__abc_49347_n3188_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_44 ( .CLK(clk_i_bF_buf41), .D(u0_sp_csc_5__FF_INPUT), .Q(sp_csc_5_), .R(u0__abc_49347_n3188_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_45 ( .CLK(clk_i_bF_buf40), .D(u0_sp_csc_6__FF_INPUT), .Q(sp_csc_6_), .R(u0__abc_49347_n3188_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_46 ( .CLK(clk_i_bF_buf39), .D(u0_sp_csc_7__FF_INPUT), .Q(sp_csc_7_), .R(u0__abc_49347_n3188_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_47 ( .CLK(clk_i_bF_buf38), .D(u0_sp_csc_9__FF_INPUT), .Q(sp_csc_9_), .R(u0__abc_49347_n3188_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_48 ( .CLK(clk_i_bF_buf37), .D(u0_sp_csc_10__FF_INPUT), .Q(sp_csc_10_), .R(u0__abc_49347_n3188_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_49 ( .CLK(clk_i_bF_buf36), .D(u0_tms_0__FF_INPUT), .Q(tms_0_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf6) );
  DFFSR DFFSR_5 ( .CLK(clk_i_bF_buf80), .D(u0_spec_req_cs_1__FF_INPUT), .Q(spec_req_cs_1_), .R(u0__abc_49347_n3188_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_50 ( .CLK(clk_i_bF_buf35), .D(u0_tms_1__FF_INPUT), .Q(tms_1_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf5) );
  DFFSR DFFSR_51 ( .CLK(clk_i_bF_buf34), .D(u0_tms_2__FF_INPUT), .Q(tms_2_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf4) );
  DFFSR DFFSR_52 ( .CLK(clk_i_bF_buf33), .D(u0_tms_3__FF_INPUT), .Q(tms_3_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf3) );
  DFFSR DFFSR_53 ( .CLK(clk_i_bF_buf32), .D(u0_tms_4__FF_INPUT), .Q(tms_4_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf2) );
  DFFSR DFFSR_54 ( .CLK(clk_i_bF_buf31), .D(u0_tms_5__FF_INPUT), .Q(tms_5_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf1) );
  DFFSR DFFSR_55 ( .CLK(clk_i_bF_buf30), .D(u0_tms_6__FF_INPUT), .Q(tms_6_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf0) );
  DFFSR DFFSR_56 ( .CLK(clk_i_bF_buf29), .D(u0_tms_7__FF_INPUT), .Q(tms_7_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf10) );
  DFFSR DFFSR_57 ( .CLK(clk_i_bF_buf28), .D(u0_tms_8__FF_INPUT), .Q(tms_8_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf9) );
  DFFSR DFFSR_58 ( .CLK(clk_i_bF_buf27), .D(u0_tms_9__FF_INPUT), .Q(tms_9_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf8) );
  DFFSR DFFSR_59 ( .CLK(clk_i_bF_buf26), .D(u0_tms_10__FF_INPUT), .Q(tms_10_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf7) );
  DFFSR DFFSR_6 ( .CLK(clk_i_bF_buf79), .D(u0_spec_req_cs_2__FF_INPUT), .Q(spec_req_cs_2_), .R(u0__abc_49347_n3188_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_60 ( .CLK(clk_i_bF_buf25), .D(u0_tms_11__FF_INPUT), .Q(tms_11_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf6) );
  DFFSR DFFSR_61 ( .CLK(clk_i_bF_buf24), .D(u0_tms_12__FF_INPUT), .Q(tms_12_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf5) );
  DFFSR DFFSR_62 ( .CLK(clk_i_bF_buf23), .D(u0_tms_13__FF_INPUT), .Q(tms_13_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf4) );
  DFFSR DFFSR_63 ( .CLK(clk_i_bF_buf22), .D(u0_tms_14__FF_INPUT), .Q(tms_14_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf3) );
  DFFSR DFFSR_64 ( .CLK(clk_i_bF_buf21), .D(u0_tms_15__FF_INPUT), .Q(tms_15_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf2) );
  DFFSR DFFSR_65 ( .CLK(clk_i_bF_buf20), .D(u0_tms_16__FF_INPUT), .Q(tms_16_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf1) );
  DFFSR DFFSR_66 ( .CLK(clk_i_bF_buf19), .D(u0_tms_17__FF_INPUT), .Q(tms_17_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf0) );
  DFFSR DFFSR_67 ( .CLK(clk_i_bF_buf18), .D(u0_tms_18__FF_INPUT), .Q(tms_18_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf10) );
  DFFSR DFFSR_68 ( .CLK(clk_i_bF_buf17), .D(u0_tms_19__FF_INPUT), .Q(tms_19_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf9) );
  DFFSR DFFSR_69 ( .CLK(clk_i_bF_buf16), .D(u0_tms_20__FF_INPUT), .Q(tms_20_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf8) );
  DFFSR DFFSR_7 ( .CLK(clk_i_bF_buf78), .D(u0_spec_req_cs_3__FF_INPUT), .Q(spec_req_cs_3_), .R(u0__abc_49347_n3188_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_70 ( .CLK(clk_i_bF_buf15), .D(u0_tms_21__FF_INPUT), .Q(tms_21_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf7) );
  DFFSR DFFSR_71 ( .CLK(clk_i_bF_buf14), .D(u0_tms_22__FF_INPUT), .Q(tms_22_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf6) );
  DFFSR DFFSR_72 ( .CLK(clk_i_bF_buf13), .D(u0_tms_23__FF_INPUT), .Q(tms_23_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf5) );
  DFFSR DFFSR_73 ( .CLK(clk_i_bF_buf12), .D(u0_tms_24__FF_INPUT), .Q(tms_24_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf4) );
  DFFSR DFFSR_74 ( .CLK(clk_i_bF_buf11), .D(u0_tms_25__FF_INPUT), .Q(tms_25_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf3) );
  DFFSR DFFSR_75 ( .CLK(clk_i_bF_buf10), .D(u0_tms_26__FF_INPUT), .Q(tms_26_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf2) );
  DFFSR DFFSR_76 ( .CLK(clk_i_bF_buf9), .D(u0_tms_27__FF_INPUT), .Q(tms_27_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf1) );
  DFFSR DFFSR_77 ( .CLK(clk_i_bF_buf8), .D(u0_csc_1__FF_INPUT), .Q(csc_1_), .R(u0__abc_49347_n3188_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_78 ( .CLK(clk_i_bF_buf7), .D(u0_csc_2__FF_INPUT), .Q(csc_2_), .R(u0__abc_49347_n3188_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_79 ( .CLK(clk_i_bF_buf6), .D(u0_csc_3__FF_INPUT), .Q(csc_3_), .R(u0__abc_49347_n3188_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_8 ( .CLK(clk_i_bF_buf77), .D(u0_spec_req_cs_4__FF_INPUT), .Q(spec_req_cs_4_), .R(u0__abc_49347_n3188_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_80 ( .CLK(clk_i_bF_buf5), .D(u0_csc_4__FF_INPUT), .Q(csc_4_), .R(u0__abc_49347_n3188_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_81 ( .CLK(clk_i_bF_buf4), .D(u0_csc_5__FF_INPUT), .Q(csc_5_), .R(u0__abc_49347_n3188_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_82 ( .CLK(clk_i_bF_buf3), .D(u0_csc_6__FF_INPUT), .Q(csc_6_), .R(u0__abc_49347_n3188_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_83 ( .CLK(clk_i_bF_buf2), .D(u0_csc_7__FF_INPUT), .Q(csc_7_), .R(u0__abc_49347_n3188_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_84 ( .CLK(clk_i_bF_buf1), .D(u0_csc_9__FF_INPUT), .Q(csc_9_), .R(u0__abc_49347_n3188_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_85 ( .CLK(clk_i_bF_buf0), .D(u0_csc_10__FF_INPUT), .Q(csc_10_), .R(u0__abc_49347_n3188_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_86 ( .CLK(clk_i_bF_buf125), .D(u0_csc_11__FF_INPUT), .Q(u3_pen), .R(u0__abc_49347_n3188_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_87 ( .CLK(clk_i_bF_buf124), .D(u0_wp_err_FF_INPUT), .Q(u0_wp_err), .R(u0__abc_49347_n3188_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_88 ( .CLK(clk_i_bF_buf123), .D(u0_cs_0__FF_INPUT), .Q(cs_0_), .R(u0__abc_49347_n3188_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_89 ( .CLK(clk_i_bF_buf122), .D(u0_cs_1__FF_INPUT), .Q(cs_1_), .R(u0__abc_49347_n3188_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_9 ( .CLK(clk_i_bF_buf76), .D(u0_spec_req_cs_5__FF_INPUT), .Q(spec_req_cs_5_), .R(u0__abc_49347_n3188_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_90 ( .CLK(clk_i_bF_buf121), .D(u0_cs_2__FF_INPUT), .Q(cs_2_), .R(u0__abc_49347_n3188_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_91 ( .CLK(clk_i_bF_buf120), .D(u0_cs_3__FF_INPUT), .Q(cs_3_), .R(u0__abc_49347_n3188_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_92 ( .CLK(clk_i_bF_buf119), .D(u0_cs_4__FF_INPUT), .Q(cs_4_), .R(u0__abc_49347_n3188_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_93 ( .CLK(clk_i_bF_buf118), .D(u0_cs_5__FF_INPUT), .Q(cs_5_), .R(u0__abc_49347_n3188_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_94 ( .CLK(clk_i_bF_buf117), .D(u0_cs_6__FF_INPUT), .Q(cs_6_), .R(u0__abc_49347_n3188_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_95 ( .CLK(clk_i_bF_buf116), .D(u0_cs_7__FF_INPUT), .Q(cs_7_), .R(u0__abc_49347_n3188_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_96 ( .CLK(clk_i_bF_buf115), .D(u0_rst_r2), .Q(u0_rst_r3), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf3) );
  DFFSR DFFSR_97 ( .CLK(clk_i_bF_buf114), .D(u0_rst_r1), .Q(u0_rst_r2), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf2) );
  DFFSR DFFSR_98 ( .CLK(clk_i_bF_buf113), .D(1'b0), .Q(u0_rst_r1), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf1) );
  DFFSR DFFSR_99 ( .CLK(clk_i_bF_buf112), .D(u0_csc_mask_r_0__FF_INPUT), .Q(u0_csc_mask_0_), .R(1'b1), .S(u0__abc_49347_n3188_bF_buf0) );
  INVX1 INVX1_1 ( .A(init_ack), .Y(_abc_55805_n238_1) );
  INVX1 INVX1_10 ( .A(u0__abc_49347_n1157), .Y(u0__abc_49347_n1164_1) );
  INVX1 INVX1_100 ( .A(u0_u1__abc_43657_n233_1), .Y(u0_u1__abc_43657_n234_1) );
  INVX1 INVX1_1000 ( .A(\wb_data_i[1] ), .Y(u3__abc_46775_n285_1) );
  INVX1 INVX1_1001 ( .A(\wb_data_i[0] ), .Y(u3__abc_46775_n287_1) );
  INVX1 INVX1_1002 ( .A(u3__abc_46775_n290_1), .Y(u3__abc_46775_n291_1) );
  INVX1 INVX1_1003 ( .A(u3__abc_46775_n293), .Y(u3__abc_46775_n294) );
  INVX1 INVX1_1004 ( .A(u3__abc_46775_n296_1), .Y(u3__abc_46775_n297_1) );
  INVX1 INVX1_1005 ( .A(u3__abc_46775_n298), .Y(u3__abc_46775_n299) );
  INVX1 INVX1_1006 ( .A(\wb_data_i[5] ), .Y(u3__abc_46775_n300_1) );
  INVX1 INVX1_1007 ( .A(\wb_data_i[4] ), .Y(u3__abc_46775_n302_1) );
  INVX1 INVX1_1008 ( .A(u3__abc_46775_n304), .Y(u3__abc_46775_n305_1) );
  INVX1 INVX1_1009 ( .A(u3__abc_46775_n308), .Y(u3__abc_46775_n309) );
  INVX1 INVX1_101 ( .A(\wb_data_i[3] ), .Y(u0_u1__abc_43657_n238) );
  INVX1 INVX1_1010 ( .A(u3__abc_46775_n317_1), .Y(u3__abc_46775_n318) );
  INVX1 INVX1_1011 ( .A(\wb_data_i[9] ), .Y(u3__abc_46775_n320_1) );
  INVX1 INVX1_1012 ( .A(\wb_data_i[8] ), .Y(u3__abc_46775_n322_1) );
  INVX1 INVX1_1013 ( .A(u3__abc_46775_n324), .Y(u3__abc_46775_n325_1) );
  INVX1 INVX1_1014 ( .A(u3__abc_46775_n326_1), .Y(u3__abc_46775_n327_1) );
  INVX1 INVX1_1015 ( .A(u3__abc_46775_n329), .Y(u3__abc_46775_n330_1) );
  INVX1 INVX1_1016 ( .A(u3__abc_46775_n332_1), .Y(u3__abc_46775_n333) );
  INVX1 INVX1_1017 ( .A(u3__abc_46775_n334), .Y(u3__abc_46775_n335_1) );
  INVX1 INVX1_1018 ( .A(\wb_data_i[13] ), .Y(u3__abc_46775_n336_1) );
  INVX1 INVX1_1019 ( .A(\wb_data_i[12] ), .Y(u3__abc_46775_n338) );
  INVX1 INVX1_102 ( .A(u0_u1__abc_43657_n239_1), .Y(u0_u1__abc_43657_n240_1) );
  INVX1 INVX1_1020 ( .A(u3__abc_46775_n340_1), .Y(u3__abc_46775_n341_1) );
  INVX1 INVX1_1021 ( .A(u3__abc_46775_n344), .Y(u3__abc_46775_n345_1) );
  INVX1 INVX1_1022 ( .A(u3__abc_46775_n352_1), .Y(u3__abc_46775_n353) );
  INVX1 INVX1_1023 ( .A(\wb_data_i[17] ), .Y(u3__abc_46775_n355_1) );
  INVX1 INVX1_1024 ( .A(\wb_data_i[16] ), .Y(u3__abc_46775_n357_1) );
  INVX1 INVX1_1025 ( .A(u3__abc_46775_n359), .Y(u3__abc_46775_n360_1) );
  INVX1 INVX1_1026 ( .A(u3__abc_46775_n361_1), .Y(u3__abc_46775_n362_1) );
  INVX1 INVX1_1027 ( .A(u3__abc_46775_n366_1), .Y(u3__abc_46775_n367_1) );
  INVX1 INVX1_1028 ( .A(u3__abc_46775_n368_1), .Y(u3__abc_46775_n369) );
  INVX1 INVX1_1029 ( .A(\wb_data_i[21] ), .Y(u3__abc_46775_n370_1) );
  INVX1 INVX1_103 ( .A(\wb_data_i[4] ), .Y(u0_u1__abc_43657_n244) );
  INVX1 INVX1_1030 ( .A(\wb_data_i[20] ), .Y(u3__abc_46775_n372_1) );
  INVX1 INVX1_1031 ( .A(u3__abc_46775_n374), .Y(u3__abc_46775_n375) );
  INVX1 INVX1_1032 ( .A(u3__abc_46775_n378), .Y(u3__abc_46775_n379) );
  INVX1 INVX1_1033 ( .A(u3__abc_46775_n364), .Y(u3__abc_46775_n381_1) );
  INVX1 INVX1_1034 ( .A(u3__abc_46775_n388), .Y(u3__abc_46775_n389) );
  INVX1 INVX1_1035 ( .A(\wb_data_i[25] ), .Y(u3__abc_46775_n391) );
  INVX1 INVX1_1036 ( .A(\wb_data_i[24] ), .Y(u3__abc_46775_n393_1) );
  INVX1 INVX1_1037 ( .A(u3__abc_46775_n395), .Y(u3__abc_46775_n396) );
  INVX1 INVX1_1038 ( .A(u3__abc_46775_n397), .Y(u3__abc_46775_n398) );
  INVX1 INVX1_1039 ( .A(u3__abc_46775_n402_1), .Y(u3__abc_46775_n403) );
  INVX1 INVX1_104 ( .A(u0_u1__abc_43657_n245_1), .Y(u0_u1__abc_43657_n246_1) );
  INVX1 INVX1_1040 ( .A(u3__abc_46775_n404), .Y(u3__abc_46775_n405) );
  INVX1 INVX1_1041 ( .A(\wb_data_i[29] ), .Y(u3__abc_46775_n406) );
  INVX1 INVX1_1042 ( .A(\wb_data_i[28] ), .Y(u3__abc_46775_n408) );
  INVX1 INVX1_1043 ( .A(u3__abc_46775_n410), .Y(u3__abc_46775_n411_1) );
  INVX1 INVX1_1044 ( .A(u3__abc_46775_n414_1), .Y(u3__abc_46775_n415) );
  INVX1 INVX1_1045 ( .A(u3__abc_46775_n400), .Y(u3__abc_46775_n417) );
  INVX1 INVX1_1046 ( .A(csc_4_), .Y(u3__abc_46775_n449) );
  INVX1 INVX1_1047 ( .A(wb_cyc_i), .Y(u3__abc_46775_n850) );
  INVX1 INVX1_1048 ( .A(u3__abc_46775_n855), .Y(u3__abc_46775_n856) );
  INVX1 INVX1_1049 ( .A(u3__abc_46775_n857), .Y(u3__abc_46775_n858) );
  INVX1 INVX1_105 ( .A(\wb_data_i[5] ), .Y(u0_u1__abc_43657_n250) );
  INVX1 INVX1_1050 ( .A(u3_rd_fifo_out_33_), .Y(u3__abc_46775_n859) );
  INVX1 INVX1_1051 ( .A(u3_rd_fifo_out_9_), .Y(u3__abc_46775_n860) );
  INVX1 INVX1_1052 ( .A(u3_rd_fifo_out_8_), .Y(u3__abc_46775_n862) );
  INVX1 INVX1_1053 ( .A(u3__abc_46775_n876), .Y(u3__abc_46775_n877) );
  INVX1 INVX1_1054 ( .A(u3__abc_46775_n879), .Y(u3__abc_46775_n880) );
  INVX1 INVX1_1055 ( .A(u3__abc_46775_n881), .Y(u3__abc_46775_n882) );
  INVX1 INVX1_1056 ( .A(u3_rd_fifo_out_11_), .Y(u3__abc_46775_n883) );
  INVX1 INVX1_1057 ( .A(u3__abc_46775_n884), .Y(u3__abc_46775_n885) );
  INVX1 INVX1_1058 ( .A(u3__abc_46775_n887), .Y(u3__abc_46775_n888) );
  INVX1 INVX1_1059 ( .A(u3__abc_46775_n891), .Y(u3__abc_46775_n892) );
  INVX1 INVX1_106 ( .A(u0_u1__abc_43657_n251_1), .Y(u0_u1__abc_43657_n252_1) );
  INVX1 INVX1_1060 ( .A(u3__abc_46775_n898), .Y(u3__abc_46775_n899) );
  INVX1 INVX1_1061 ( .A(u3__abc_46775_n900), .Y(u3__abc_46775_n901) );
  INVX1 INVX1_1062 ( .A(u3_rd_fifo_out_34_), .Y(u3__abc_46775_n902) );
  INVX1 INVX1_1063 ( .A(u3__abc_46775_n904), .Y(u3__abc_46775_n905) );
  INVX1 INVX1_1064 ( .A(u3_rd_fifo_out_16_), .Y(u3__abc_46775_n908) );
  INVX1 INVX1_1065 ( .A(u3_rd_fifo_out_17_), .Y(u3__abc_46775_n909) );
  INVX1 INVX1_1066 ( .A(u3__abc_46775_n919), .Y(u3__abc_46775_n920) );
  INVX1 INVX1_1067 ( .A(u3__abc_46775_n922), .Y(u3__abc_46775_n923) );
  INVX1 INVX1_1068 ( .A(u3__abc_46775_n924), .Y(u3__abc_46775_n925) );
  INVX1 INVX1_1069 ( .A(u3_rd_fifo_out_19_), .Y(u3__abc_46775_n926) );
  INVX1 INVX1_107 ( .A(\wb_data_i[6] ), .Y(u0_u1__abc_43657_n256) );
  INVX1 INVX1_1070 ( .A(u3__abc_46775_n927), .Y(u3__abc_46775_n928) );
  INVX1 INVX1_1071 ( .A(u3__abc_46775_n930), .Y(u3__abc_46775_n931) );
  INVX1 INVX1_1072 ( .A(u3__abc_46775_n934), .Y(u3__abc_46775_n935) );
  INVX1 INVX1_1073 ( .A(u3__abc_46775_n942), .Y(u3__abc_46775_n943) );
  INVX1 INVX1_1074 ( .A(u3__abc_46775_n944), .Y(u3__abc_46775_n945) );
  INVX1 INVX1_1075 ( .A(u3_rd_fifo_out_32_), .Y(u3__abc_46775_n946) );
  INVX1 INVX1_1076 ( .A(u3__abc_46775_n948), .Y(u3__abc_46775_n949) );
  INVX1 INVX1_1077 ( .A(u3_rd_fifo_out_0_), .Y(u3__abc_46775_n952) );
  INVX1 INVX1_1078 ( .A(u3_rd_fifo_out_1_), .Y(u3__abc_46775_n953) );
  INVX1 INVX1_1079 ( .A(u3__abc_46775_n963), .Y(u3__abc_46775_n964) );
  INVX1 INVX1_108 ( .A(u0_u1__abc_43657_n257), .Y(u0_u1__abc_43657_n258) );
  INVX1 INVX1_1080 ( .A(u3__abc_46775_n966), .Y(u3__abc_46775_n967) );
  INVX1 INVX1_1081 ( .A(u3__abc_46775_n968), .Y(u3__abc_46775_n969) );
  INVX1 INVX1_1082 ( .A(u3_rd_fifo_out_3_), .Y(u3__abc_46775_n970) );
  INVX1 INVX1_1083 ( .A(u3__abc_46775_n971), .Y(u3__abc_46775_n972) );
  INVX1 INVX1_1084 ( .A(u3__abc_46775_n974), .Y(u3__abc_46775_n975) );
  INVX1 INVX1_1085 ( .A(u3__abc_46775_n978), .Y(u3__abc_46775_n979) );
  INVX1 INVX1_1086 ( .A(u3__abc_46775_n985), .Y(u3__abc_46775_n986) );
  INVX1 INVX1_1087 ( .A(u3__abc_46775_n987), .Y(u3__abc_46775_n988) );
  INVX1 INVX1_1088 ( .A(u3_rd_fifo_out_35_), .Y(u3__abc_46775_n989) );
  INVX1 INVX1_1089 ( .A(u3__abc_46775_n991), .Y(u3__abc_46775_n992) );
  INVX1 INVX1_109 ( .A(\wb_data_i[7] ), .Y(u0_u1__abc_43657_n262) );
  INVX1 INVX1_1090 ( .A(u3_rd_fifo_out_24_), .Y(u3__abc_46775_n995) );
  INVX1 INVX1_1091 ( .A(u3_rd_fifo_out_25_), .Y(u3__abc_46775_n997) );
  INVX1 INVX1_1092 ( .A(u3__abc_46775_n1007), .Y(u3__abc_46775_n1008) );
  INVX1 INVX1_1093 ( .A(u3__abc_46775_n1010), .Y(u3__abc_46775_n1011) );
  INVX1 INVX1_1094 ( .A(u3__abc_46775_n1012), .Y(u3__abc_46775_n1013) );
  INVX1 INVX1_1095 ( .A(u3_rd_fifo_out_27_), .Y(u3__abc_46775_n1014) );
  INVX1 INVX1_1096 ( .A(u3__abc_46775_n1015), .Y(u3__abc_46775_n1016) );
  INVX1 INVX1_1097 ( .A(u3__abc_46775_n1018), .Y(u3__abc_46775_n1019) );
  INVX1 INVX1_1098 ( .A(u3__abc_46775_n1022), .Y(u3__abc_46775_n1023) );
  INVX1 INVX1_1099 ( .A(wb_we_i), .Y(u3__abc_46775_n1030) );
  INVX1 INVX1_11 ( .A(u0__abc_49347_n4265), .Y(u0__abc_49347_n4274) );
  INVX1 INVX1_110 ( .A(u0_u1__abc_43657_n263), .Y(u0_u1__abc_43657_n264) );
  INVX1 INVX1_1100 ( .A(mc_data_ir_0_), .Y(u3_u0__abc_48231_n384_1) );
  INVX1 INVX1_1101 ( .A(u3_u0__abc_48231_n385), .Y(u3_u0__abc_48231_n386) );
  INVX1 INVX1_1102 ( .A(mc_data_ir_1_), .Y(u3_u0__abc_48231_n389) );
  INVX1 INVX1_1103 ( .A(u3_u0__abc_48231_n390), .Y(u3_u0__abc_48231_n391) );
  INVX1 INVX1_1104 ( .A(mc_data_ir_2_), .Y(u3_u0__abc_48231_n394) );
  INVX1 INVX1_1105 ( .A(u3_u0__abc_48231_n395), .Y(u3_u0__abc_48231_n396_1) );
  INVX1 INVX1_1106 ( .A(mc_data_ir_3_), .Y(u3_u0__abc_48231_n399) );
  INVX1 INVX1_1107 ( .A(u3_u0__abc_48231_n400_1), .Y(u3_u0__abc_48231_n401) );
  INVX1 INVX1_1108 ( .A(mc_data_ir_4_), .Y(u3_u0__abc_48231_n404_1) );
  INVX1 INVX1_1109 ( .A(u3_u0__abc_48231_n405), .Y(u3_u0__abc_48231_n406) );
  INVX1 INVX1_111 ( .A(\wb_data_i[8] ), .Y(u0_u1__abc_43657_n268) );
  INVX1 INVX1_1110 ( .A(mc_data_ir_5_), .Y(u3_u0__abc_48231_n409) );
  INVX1 INVX1_1111 ( .A(u3_u0__abc_48231_n410), .Y(u3_u0__abc_48231_n411) );
  INVX1 INVX1_1112 ( .A(mc_data_ir_6_), .Y(u3_u0__abc_48231_n414) );
  INVX1 INVX1_1113 ( .A(u3_u0__abc_48231_n415), .Y(u3_u0__abc_48231_n416_1) );
  INVX1 INVX1_1114 ( .A(mc_data_ir_7_), .Y(u3_u0__abc_48231_n419) );
  INVX1 INVX1_1115 ( .A(u3_u0__abc_48231_n420_1), .Y(u3_u0__abc_48231_n421) );
  INVX1 INVX1_1116 ( .A(mc_data_ir_8_), .Y(u3_u0__abc_48231_n424_1) );
  INVX1 INVX1_1117 ( .A(u3_u0__abc_48231_n425), .Y(u3_u0__abc_48231_n426) );
  INVX1 INVX1_1118 ( .A(mc_data_ir_9_), .Y(u3_u0__abc_48231_n429) );
  INVX1 INVX1_1119 ( .A(u3_u0__abc_48231_n430), .Y(u3_u0__abc_48231_n431) );
  INVX1 INVX1_112 ( .A(u0_u1__abc_43657_n269), .Y(u0_u1__abc_43657_n270) );
  INVX1 INVX1_1120 ( .A(mc_data_ir_10_), .Y(u3_u0__abc_48231_n434) );
  INVX1 INVX1_1121 ( .A(u3_u0__abc_48231_n435), .Y(u3_u0__abc_48231_n436_1) );
  INVX1 INVX1_1122 ( .A(mc_data_ir_11_), .Y(u3_u0__abc_48231_n439) );
  INVX1 INVX1_1123 ( .A(u3_u0__abc_48231_n440_1), .Y(u3_u0__abc_48231_n441) );
  INVX1 INVX1_1124 ( .A(mc_data_ir_12_), .Y(u3_u0__abc_48231_n444_1) );
  INVX1 INVX1_1125 ( .A(u3_u0__abc_48231_n445), .Y(u3_u0__abc_48231_n446) );
  INVX1 INVX1_1126 ( .A(mc_data_ir_13_), .Y(u3_u0__abc_48231_n449) );
  INVX1 INVX1_1127 ( .A(u3_u0__abc_48231_n450), .Y(u3_u0__abc_48231_n451) );
  INVX1 INVX1_1128 ( .A(mc_data_ir_14_), .Y(u3_u0__abc_48231_n454) );
  INVX1 INVX1_1129 ( .A(u3_u0__abc_48231_n455), .Y(u3_u0__abc_48231_n456_1) );
  INVX1 INVX1_113 ( .A(\wb_data_i[9] ), .Y(u0_u1__abc_43657_n274_1) );
  INVX1 INVX1_1130 ( .A(mc_data_ir_15_), .Y(u3_u0__abc_48231_n459) );
  INVX1 INVX1_1131 ( .A(u3_u0__abc_48231_n460_1), .Y(u3_u0__abc_48231_n461) );
  INVX1 INVX1_1132 ( .A(mc_data_ir_16_), .Y(u3_u0__abc_48231_n464_1) );
  INVX1 INVX1_1133 ( .A(u3_u0__abc_48231_n465), .Y(u3_u0__abc_48231_n466) );
  INVX1 INVX1_1134 ( .A(mc_data_ir_17_), .Y(u3_u0__abc_48231_n469) );
  INVX1 INVX1_1135 ( .A(u3_u0__abc_48231_n470), .Y(u3_u0__abc_48231_n471) );
  INVX1 INVX1_1136 ( .A(mc_data_ir_18_), .Y(u3_u0__abc_48231_n474) );
  INVX1 INVX1_1137 ( .A(u3_u0__abc_48231_n475), .Y(u3_u0__abc_48231_n476_1) );
  INVX1 INVX1_1138 ( .A(mc_data_ir_19_), .Y(u3_u0__abc_48231_n479) );
  INVX1 INVX1_1139 ( .A(u3_u0__abc_48231_n480_1), .Y(u3_u0__abc_48231_n481) );
  INVX1 INVX1_114 ( .A(u0_u1__abc_43657_n275), .Y(u0_u1__abc_43657_n276_1) );
  INVX1 INVX1_1140 ( .A(mc_data_ir_20_), .Y(u3_u0__abc_48231_n484_1) );
  INVX1 INVX1_1141 ( .A(u3_u0__abc_48231_n485), .Y(u3_u0__abc_48231_n486) );
  INVX1 INVX1_1142 ( .A(mc_data_ir_21_), .Y(u3_u0__abc_48231_n489) );
  INVX1 INVX1_1143 ( .A(u3_u0__abc_48231_n490), .Y(u3_u0__abc_48231_n491) );
  INVX1 INVX1_1144 ( .A(mc_data_ir_22_), .Y(u3_u0__abc_48231_n494) );
  INVX1 INVX1_1145 ( .A(u3_u0__abc_48231_n495), .Y(u3_u0__abc_48231_n496_1) );
  INVX1 INVX1_1146 ( .A(mc_data_ir_23_), .Y(u3_u0__abc_48231_n499) );
  INVX1 INVX1_1147 ( .A(u3_u0__abc_48231_n500_1), .Y(u3_u0__abc_48231_n501) );
  INVX1 INVX1_1148 ( .A(mc_data_ir_24_), .Y(u3_u0__abc_48231_n504_1) );
  INVX1 INVX1_1149 ( .A(u3_u0__abc_48231_n505), .Y(u3_u0__abc_48231_n506) );
  INVX1 INVX1_115 ( .A(\wb_data_i[10] ), .Y(u0_u1__abc_43657_n280) );
  INVX1 INVX1_1150 ( .A(mc_data_ir_25_), .Y(u3_u0__abc_48231_n509) );
  INVX1 INVX1_1151 ( .A(u3_u0__abc_48231_n510), .Y(u3_u0__abc_48231_n511) );
  INVX1 INVX1_1152 ( .A(mc_data_ir_26_), .Y(u3_u0__abc_48231_n514_1) );
  INVX1 INVX1_1153 ( .A(u3_u0__abc_48231_n515), .Y(u3_u0__abc_48231_n516) );
  INVX1 INVX1_1154 ( .A(mc_data_ir_27_), .Y(u3_u0__abc_48231_n519) );
  INVX1 INVX1_1155 ( .A(u3_u0__abc_48231_n520), .Y(u3_u0__abc_48231_n521) );
  INVX1 INVX1_1156 ( .A(mc_data_ir_28_), .Y(u3_u0__abc_48231_n524) );
  INVX1 INVX1_1157 ( .A(u3_u0__abc_48231_n525), .Y(u3_u0__abc_48231_n526) );
  INVX1 INVX1_1158 ( .A(mc_data_ir_29_), .Y(u3_u0__abc_48231_n529) );
  INVX1 INVX1_1159 ( .A(u3_u0__abc_48231_n530), .Y(u3_u0__abc_48231_n531) );
  INVX1 INVX1_116 ( .A(u0_u1__abc_43657_n281), .Y(u0_u1__abc_43657_n282_1) );
  INVX1 INVX1_1160 ( .A(mc_data_ir_30_), .Y(u3_u0__abc_48231_n534) );
  INVX1 INVX1_1161 ( .A(u3_u0__abc_48231_n535), .Y(u3_u0__abc_48231_n536) );
  INVX1 INVX1_1162 ( .A(mc_data_ir_31_), .Y(u3_u0__abc_48231_n539) );
  INVX1 INVX1_1163 ( .A(u3_u0__abc_48231_n540), .Y(u3_u0__abc_48231_n541) );
  INVX1 INVX1_1164 ( .A(mc_data_ir_32_), .Y(u3_u0__abc_48231_n544) );
  INVX1 INVX1_1165 ( .A(u3_u0__abc_48231_n545), .Y(u3_u0__abc_48231_n546) );
  INVX1 INVX1_1166 ( .A(mc_data_ir_33_), .Y(u3_u0__abc_48231_n549) );
  INVX1 INVX1_1167 ( .A(u3_u0__abc_48231_n550), .Y(u3_u0__abc_48231_n551) );
  INVX1 INVX1_1168 ( .A(mc_data_ir_34_), .Y(u3_u0__abc_48231_n554) );
  INVX1 INVX1_1169 ( .A(u3_u0__abc_48231_n555), .Y(u3_u0__abc_48231_n556) );
  INVX1 INVX1_117 ( .A(\wb_data_i[11] ), .Y(u0_u1__abc_43657_n286_1) );
  INVX1 INVX1_1170 ( .A(mc_data_ir_35_), .Y(u3_u0__abc_48231_n559) );
  INVX1 INVX1_1171 ( .A(u3_u0__abc_48231_n560), .Y(u3_u0__abc_48231_n561) );
  INVX1 INVX1_1172 ( .A(u3_u0__abc_48231_n565), .Y(u3_u0__abc_48231_n566) );
  INVX1 INVX1_1173 ( .A(u3_u0__abc_48231_n569), .Y(u3_u0__abc_48231_n570) );
  INVX1 INVX1_1174 ( .A(u3_u0__abc_48231_n573), .Y(u3_u0__abc_48231_n574) );
  INVX1 INVX1_1175 ( .A(u3_u0__abc_48231_n577), .Y(u3_u0__abc_48231_n578) );
  INVX1 INVX1_1176 ( .A(u3_u0__abc_48231_n581), .Y(u3_u0__abc_48231_n582) );
  INVX1 INVX1_1177 ( .A(u3_u0__abc_48231_n585), .Y(u3_u0__abc_48231_n586) );
  INVX1 INVX1_1178 ( .A(u3_u0__abc_48231_n589), .Y(u3_u0__abc_48231_n590) );
  INVX1 INVX1_1179 ( .A(u3_u0__abc_48231_n593), .Y(u3_u0__abc_48231_n594) );
  INVX1 INVX1_118 ( .A(u0_u1__abc_43657_n287), .Y(u0_u1__abc_43657_n288_1) );
  INVX1 INVX1_1180 ( .A(u3_u0__abc_48231_n597), .Y(u3_u0__abc_48231_n598) );
  INVX1 INVX1_1181 ( .A(u3_u0__abc_48231_n601), .Y(u3_u0__abc_48231_n602) );
  INVX1 INVX1_1182 ( .A(u3_u0__abc_48231_n605), .Y(u3_u0__abc_48231_n606) );
  INVX1 INVX1_1183 ( .A(u3_u0__abc_48231_n609), .Y(u3_u0__abc_48231_n610) );
  INVX1 INVX1_1184 ( .A(u3_u0__abc_48231_n613), .Y(u3_u0__abc_48231_n614) );
  INVX1 INVX1_1185 ( .A(u3_u0__abc_48231_n617), .Y(u3_u0__abc_48231_n618) );
  INVX1 INVX1_1186 ( .A(u3_u0__abc_48231_n621), .Y(u3_u0__abc_48231_n622) );
  INVX1 INVX1_1187 ( .A(u3_u0__abc_48231_n625), .Y(u3_u0__abc_48231_n626) );
  INVX1 INVX1_1188 ( .A(u3_u0__abc_48231_n629), .Y(u3_u0__abc_48231_n630) );
  INVX1 INVX1_1189 ( .A(u3_u0__abc_48231_n633), .Y(u3_u0__abc_48231_n634) );
  INVX1 INVX1_119 ( .A(\wb_data_i[12] ), .Y(u0_u1__abc_43657_n292) );
  INVX1 INVX1_1190 ( .A(u3_u0__abc_48231_n637), .Y(u3_u0__abc_48231_n638) );
  INVX1 INVX1_1191 ( .A(u3_u0__abc_48231_n641), .Y(u3_u0__abc_48231_n642) );
  INVX1 INVX1_1192 ( .A(u3_u0__abc_48231_n645), .Y(u3_u0__abc_48231_n646) );
  INVX1 INVX1_1193 ( .A(u3_u0__abc_48231_n649), .Y(u3_u0__abc_48231_n650) );
  INVX1 INVX1_1194 ( .A(u3_u0__abc_48231_n653), .Y(u3_u0__abc_48231_n654) );
  INVX1 INVX1_1195 ( .A(u3_u0__abc_48231_n657), .Y(u3_u0__abc_48231_n658) );
  INVX1 INVX1_1196 ( .A(u3_u0__abc_48231_n661), .Y(u3_u0__abc_48231_n662) );
  INVX1 INVX1_1197 ( .A(u3_u0__abc_48231_n665), .Y(u3_u0__abc_48231_n666) );
  INVX1 INVX1_1198 ( .A(u3_u0__abc_48231_n669), .Y(u3_u0__abc_48231_n670) );
  INVX1 INVX1_1199 ( .A(u3_u0__abc_48231_n673), .Y(u3_u0__abc_48231_n674) );
  INVX1 INVX1_12 ( .A(u0_rf_we), .Y(u0__abc_49347_n4400) );
  INVX1 INVX1_120 ( .A(u0_u1__abc_43657_n293), .Y(u0_u1__abc_43657_n294) );
  INVX1 INVX1_1200 ( .A(u3_u0__abc_48231_n677), .Y(u3_u0__abc_48231_n678) );
  INVX1 INVX1_1201 ( .A(u3_u0__abc_48231_n681), .Y(u3_u0__abc_48231_n682) );
  INVX1 INVX1_1202 ( .A(u3_u0__abc_48231_n685), .Y(u3_u0__abc_48231_n686) );
  INVX1 INVX1_1203 ( .A(u3_u0__abc_48231_n689), .Y(u3_u0__abc_48231_n690) );
  INVX1 INVX1_1204 ( .A(u3_u0__abc_48231_n693), .Y(u3_u0__abc_48231_n694) );
  INVX1 INVX1_1205 ( .A(u3_u0__abc_48231_n697), .Y(u3_u0__abc_48231_n698) );
  INVX1 INVX1_1206 ( .A(u3_u0__abc_48231_n701), .Y(u3_u0__abc_48231_n702) );
  INVX1 INVX1_1207 ( .A(u3_u0__abc_48231_n705), .Y(u3_u0__abc_48231_n706) );
  INVX1 INVX1_1208 ( .A(u3_u0__abc_48231_n710), .Y(u3_u0__abc_48231_n711) );
  INVX1 INVX1_1209 ( .A(u3_u0__abc_48231_n714), .Y(u3_u0__abc_48231_n715) );
  INVX1 INVX1_121 ( .A(\wb_data_i[13] ), .Y(u0_u1__abc_43657_n298) );
  INVX1 INVX1_1210 ( .A(u3_u0__abc_48231_n718), .Y(u3_u0__abc_48231_n719) );
  INVX1 INVX1_1211 ( .A(u3_u0__abc_48231_n722), .Y(u3_u0__abc_48231_n723) );
  INVX1 INVX1_1212 ( .A(u3_u0__abc_48231_n726), .Y(u3_u0__abc_48231_n727) );
  INVX1 INVX1_1213 ( .A(u3_u0__abc_48231_n730), .Y(u3_u0__abc_48231_n731) );
  INVX1 INVX1_1214 ( .A(u3_u0__abc_48231_n734), .Y(u3_u0__abc_48231_n735) );
  INVX1 INVX1_1215 ( .A(u3_u0__abc_48231_n738), .Y(u3_u0__abc_48231_n739) );
  INVX1 INVX1_1216 ( .A(u3_u0__abc_48231_n742), .Y(u3_u0__abc_48231_n743) );
  INVX1 INVX1_1217 ( .A(u3_u0__abc_48231_n746), .Y(u3_u0__abc_48231_n747) );
  INVX1 INVX1_1218 ( .A(u3_u0__abc_48231_n750), .Y(u3_u0__abc_48231_n751) );
  INVX1 INVX1_1219 ( .A(u3_u0__abc_48231_n754), .Y(u3_u0__abc_48231_n755) );
  INVX1 INVX1_122 ( .A(u0_u1__abc_43657_n299), .Y(u0_u1__abc_43657_n300) );
  INVX1 INVX1_1220 ( .A(u3_u0__abc_48231_n758), .Y(u3_u0__abc_48231_n759) );
  INVX1 INVX1_1221 ( .A(u3_u0__abc_48231_n762), .Y(u3_u0__abc_48231_n763) );
  INVX1 INVX1_1222 ( .A(u3_u0__abc_48231_n766), .Y(u3_u0__abc_48231_n767) );
  INVX1 INVX1_1223 ( .A(u3_u0__abc_48231_n770), .Y(u3_u0__abc_48231_n771) );
  INVX1 INVX1_1224 ( .A(u3_u0__abc_48231_n774), .Y(u3_u0__abc_48231_n775) );
  INVX1 INVX1_1225 ( .A(u3_u0__abc_48231_n778), .Y(u3_u0__abc_48231_n779) );
  INVX1 INVX1_1226 ( .A(u3_u0__abc_48231_n782), .Y(u3_u0__abc_48231_n783) );
  INVX1 INVX1_1227 ( .A(u3_u0__abc_48231_n786), .Y(u3_u0__abc_48231_n787) );
  INVX1 INVX1_1228 ( .A(u3_u0__abc_48231_n790), .Y(u3_u0__abc_48231_n791) );
  INVX1 INVX1_1229 ( .A(u3_u0__abc_48231_n794), .Y(u3_u0__abc_48231_n795) );
  INVX1 INVX1_123 ( .A(\wb_data_i[14] ), .Y(u0_u1__abc_43657_n304) );
  INVX1 INVX1_1230 ( .A(u3_u0__abc_48231_n798), .Y(u3_u0__abc_48231_n799) );
  INVX1 INVX1_1231 ( .A(u3_u0__abc_48231_n802), .Y(u3_u0__abc_48231_n803) );
  INVX1 INVX1_1232 ( .A(u3_u0__abc_48231_n806), .Y(u3_u0__abc_48231_n807) );
  INVX1 INVX1_1233 ( .A(u3_u0__abc_48231_n810), .Y(u3_u0__abc_48231_n811) );
  INVX1 INVX1_1234 ( .A(u3_u0__abc_48231_n814), .Y(u3_u0__abc_48231_n815) );
  INVX1 INVX1_1235 ( .A(u3_u0__abc_48231_n818), .Y(u3_u0__abc_48231_n819) );
  INVX1 INVX1_1236 ( .A(u3_u0__abc_48231_n822), .Y(u3_u0__abc_48231_n823) );
  INVX1 INVX1_1237 ( .A(u3_u0__abc_48231_n826), .Y(u3_u0__abc_48231_n827) );
  INVX1 INVX1_1238 ( .A(u3_u0__abc_48231_n830), .Y(u3_u0__abc_48231_n831) );
  INVX1 INVX1_1239 ( .A(u3_u0__abc_48231_n834), .Y(u3_u0__abc_48231_n835) );
  INVX1 INVX1_124 ( .A(u0_u1__abc_43657_n305), .Y(u0_u1__abc_43657_n306) );
  INVX1 INVX1_1240 ( .A(u3_u0__abc_48231_n838), .Y(u3_u0__abc_48231_n839) );
  INVX1 INVX1_1241 ( .A(u3_u0__abc_48231_n842), .Y(u3_u0__abc_48231_n843) );
  INVX1 INVX1_1242 ( .A(u3_u0__abc_48231_n846), .Y(u3_u0__abc_48231_n847) );
  INVX1 INVX1_1243 ( .A(u3_u0__abc_48231_n850), .Y(u3_u0__abc_48231_n851) );
  INVX1 INVX1_1244 ( .A(u3_u0__abc_48231_n855), .Y(u3_u0__abc_48231_n856) );
  INVX1 INVX1_1245 ( .A(u3_u0__abc_48231_n859), .Y(u3_u0__abc_48231_n860) );
  INVX1 INVX1_1246 ( .A(u3_u0__abc_48231_n863), .Y(u3_u0__abc_48231_n864) );
  INVX1 INVX1_1247 ( .A(u3_u0__abc_48231_n867), .Y(u3_u0__abc_48231_n868) );
  INVX1 INVX1_1248 ( .A(u3_u0__abc_48231_n871), .Y(u3_u0__abc_48231_n872) );
  INVX1 INVX1_1249 ( .A(u3_u0__abc_48231_n875), .Y(u3_u0__abc_48231_n876) );
  INVX1 INVX1_125 ( .A(\wb_data_i[15] ), .Y(u0_u1__abc_43657_n310) );
  INVX1 INVX1_1250 ( .A(u3_u0__abc_48231_n879), .Y(u3_u0__abc_48231_n880) );
  INVX1 INVX1_1251 ( .A(u3_u0__abc_48231_n883), .Y(u3_u0__abc_48231_n884) );
  INVX1 INVX1_1252 ( .A(u3_u0__abc_48231_n887), .Y(u3_u0__abc_48231_n888) );
  INVX1 INVX1_1253 ( .A(u3_u0__abc_48231_n891), .Y(u3_u0__abc_48231_n892) );
  INVX1 INVX1_1254 ( .A(u3_u0__abc_48231_n895), .Y(u3_u0__abc_48231_n896) );
  INVX1 INVX1_1255 ( .A(u3_u0__abc_48231_n899), .Y(u3_u0__abc_48231_n900) );
  INVX1 INVX1_1256 ( .A(u3_u0__abc_48231_n903), .Y(u3_u0__abc_48231_n904) );
  INVX1 INVX1_1257 ( .A(u3_u0__abc_48231_n907), .Y(u3_u0__abc_48231_n908) );
  INVX1 INVX1_1258 ( .A(u3_u0__abc_48231_n911), .Y(u3_u0__abc_48231_n912) );
  INVX1 INVX1_1259 ( .A(u3_u0__abc_48231_n915), .Y(u3_u0__abc_48231_n916) );
  INVX1 INVX1_126 ( .A(u0_u1__abc_43657_n311_1), .Y(u0_u1__abc_43657_n312) );
  INVX1 INVX1_1260 ( .A(u3_u0__abc_48231_n919), .Y(u3_u0__abc_48231_n920) );
  INVX1 INVX1_1261 ( .A(u3_u0__abc_48231_n923), .Y(u3_u0__abc_48231_n924) );
  INVX1 INVX1_1262 ( .A(u3_u0__abc_48231_n927), .Y(u3_u0__abc_48231_n928) );
  INVX1 INVX1_1263 ( .A(u3_u0__abc_48231_n931), .Y(u3_u0__abc_48231_n932) );
  INVX1 INVX1_1264 ( .A(u3_u0__abc_48231_n935), .Y(u3_u0__abc_48231_n936) );
  INVX1 INVX1_1265 ( .A(u3_u0__abc_48231_n939), .Y(u3_u0__abc_48231_n940) );
  INVX1 INVX1_1266 ( .A(u3_u0__abc_48231_n943), .Y(u3_u0__abc_48231_n944) );
  INVX1 INVX1_1267 ( .A(u3_u0__abc_48231_n947), .Y(u3_u0__abc_48231_n948) );
  INVX1 INVX1_1268 ( .A(u3_u0__abc_48231_n951), .Y(u3_u0__abc_48231_n952) );
  INVX1 INVX1_1269 ( .A(u3_u0__abc_48231_n955), .Y(u3_u0__abc_48231_n956) );
  INVX1 INVX1_127 ( .A(\wb_data_i[16] ), .Y(u0_u1__abc_43657_n316_1) );
  INVX1 INVX1_1270 ( .A(u3_u0__abc_48231_n959), .Y(u3_u0__abc_48231_n960) );
  INVX1 INVX1_1271 ( .A(u3_u0__abc_48231_n963), .Y(u3_u0__abc_48231_n964) );
  INVX1 INVX1_1272 ( .A(u3_u0__abc_48231_n967), .Y(u3_u0__abc_48231_n968) );
  INVX1 INVX1_1273 ( .A(u3_u0__abc_48231_n971), .Y(u3_u0__abc_48231_n972) );
  INVX1 INVX1_1274 ( .A(u3_u0__abc_48231_n975), .Y(u3_u0__abc_48231_n976) );
  INVX1 INVX1_1275 ( .A(u3_u0__abc_48231_n979), .Y(u3_u0__abc_48231_n980) );
  INVX1 INVX1_1276 ( .A(u3_u0__abc_48231_n983), .Y(u3_u0__abc_48231_n984) );
  INVX1 INVX1_1277 ( .A(u3_u0__abc_48231_n987), .Y(u3_u0__abc_48231_n988) );
  INVX1 INVX1_1278 ( .A(u3_u0__abc_48231_n991), .Y(u3_u0__abc_48231_n992) );
  INVX1 INVX1_1279 ( .A(u3_u0__abc_48231_n995), .Y(u3_u0__abc_48231_n996) );
  INVX1 INVX1_128 ( .A(u0_u1__abc_43657_n317), .Y(u0_u1__abc_43657_n318) );
  INVX1 INVX1_1280 ( .A(dv), .Y(u3_u0__abc_48231_n998) );
  INVX1 INVX1_1281 ( .A(u3_re), .Y(u3_u0__abc_48231_n1012) );
  INVX1 INVX1_1282 ( .A(u3_u0_rd_adr_3_), .Y(u3_u0__abc_48231_n1029) );
  INVX1 INVX1_1283 ( .A(u3_u0_rd_adr_2_), .Y(u3_u0__abc_48231_n1030) );
  INVX1 INVX1_1284 ( .A(u3_u0_rd_adr_0_), .Y(u3_u0__abc_48231_n1032) );
  INVX1 INVX1_1285 ( .A(u3_u0__abc_48231_n1034_bF_buf5), .Y(u3_u0__abc_48231_n1035) );
  INVX1 INVX1_1286 ( .A(u3_u0_rd_adr_1_), .Y(u3_u0__abc_48231_n1044) );
  INVX1 INVX1_1287 ( .A(rfr_ps_val_5_), .Y(u4__abc_49152_n72) );
  INVX1 INVX1_1288 ( .A(u4_ps_cnt_5_), .Y(u4__abc_49152_n74) );
  INVX1 INVX1_1289 ( .A(rfr_ps_val_4_), .Y(u4__abc_49152_n77) );
  INVX1 INVX1_129 ( .A(\wb_data_i[17] ), .Y(u0_u1__abc_43657_n322_1) );
  INVX1 INVX1_1290 ( .A(u4_ps_cnt_4_), .Y(u4__abc_49152_n79_1) );
  INVX1 INVX1_1291 ( .A(rfr_ps_val_6_), .Y(u4__abc_49152_n83) );
  INVX1 INVX1_1292 ( .A(u4_ps_cnt_6_), .Y(u4__abc_49152_n85_1) );
  INVX1 INVX1_1293 ( .A(rfr_ps_val_7_), .Y(u4__abc_49152_n88_1) );
  INVX1 INVX1_1294 ( .A(u4_ps_cnt_7_), .Y(u4__abc_49152_n90_1) );
  INVX1 INVX1_1295 ( .A(rfr_ps_val_0_), .Y(u4__abc_49152_n95) );
  INVX1 INVX1_1296 ( .A(u4_ps_cnt_0_), .Y(u4__abc_49152_n97) );
  INVX1 INVX1_1297 ( .A(rfr_ps_val_1_), .Y(u4__abc_49152_n100) );
  INVX1 INVX1_1298 ( .A(u4_ps_cnt_1_), .Y(u4__abc_49152_n102_1) );
  INVX1 INVX1_1299 ( .A(rfr_ps_val_2_), .Y(u4__abc_49152_n106) );
  INVX1 INVX1_13 ( .A(u0__abc_49347_n4402), .Y(u0__abc_49347_n4403) );
  INVX1 INVX1_130 ( .A(u0_u1__abc_43657_n323_1), .Y(u0_u1__abc_43657_n324_1) );
  INVX1 INVX1_1300 ( .A(u4_ps_cnt_2_), .Y(u4__abc_49152_n108_1) );
  INVX1 INVX1_1301 ( .A(u4__abc_49152_n112), .Y(u4__abc_49152_n113_1) );
  INVX1 INVX1_1302 ( .A(u4__abc_49152_n117), .Y(u4_rfr_early_FF_INPUT) );
  INVX1 INVX1_1303 ( .A(u4__abc_49152_n122), .Y(u4__abc_49152_n123) );
  INVX1 INVX1_1304 ( .A(u4__abc_49152_n128), .Y(u4__abc_49152_n129_1) );
  INVX1 INVX1_1305 ( .A(u4__abc_49152_n135), .Y(u4__abc_49152_n136) );
  INVX1 INVX1_1306 ( .A(u4__abc_49152_n140), .Y(u4__abc_49152_n141_1) );
  INVX1 INVX1_1307 ( .A(u4__abc_49152_n145), .Y(u4__abc_49152_n146) );
  INVX1 INVX1_1308 ( .A(u4__abc_49152_n152), .Y(u4__abc_49152_n153) );
  INVX1 INVX1_1309 ( .A(u4__abc_49152_n156), .Y(u4__abc_49152_n157) );
  INVX1 INVX1_131 ( .A(\wb_data_i[18] ), .Y(u0_u1__abc_43657_n328) );
  INVX1 INVX1_1310 ( .A(u4__abc_49152_n163), .Y(u4__abc_49152_n164) );
  INVX1 INVX1_1311 ( .A(rfr_ps_val_3_), .Y(u4__abc_49152_n170) );
  INVX1 INVX1_1312 ( .A(u4__abc_49152_n175), .Y(u4_ps_cnt_clr) );
  INVX1 INVX1_1313 ( .A(u4__abc_49152_n178), .Y(u4__abc_49152_n179) );
  INVX1 INVX1_1314 ( .A(u4__abc_49152_n183), .Y(u4__abc_49152_n184) );
  INVX1 INVX1_1315 ( .A(u4__abc_49152_n194), .Y(u4__abc_49152_n195) );
  INVX1 INVX1_1316 ( .A(u4__abc_49152_n200), .Y(u4__abc_49152_n201) );
  INVX1 INVX1_1317 ( .A(u4__abc_49152_n205), .Y(u4__abc_49152_n206) );
  INVX1 INVX1_1318 ( .A(u4__abc_49152_n215), .Y(u4__abc_49152_n216) );
  INVX1 INVX1_1319 ( .A(u4__abc_49152_n219), .Y(u4__abc_49152_n220) );
  INVX1 INVX1_132 ( .A(u0_u1__abc_43657_n329), .Y(u0_u1__abc_43657_n330) );
  INVX1 INVX1_1320 ( .A(ref_int_0_), .Y(u4__abc_49152_n228) );
  INVX1 INVX1_1321 ( .A(ref_int_1_), .Y(u4__abc_49152_n234) );
  INVX1 INVX1_1322 ( .A(ref_int_2_), .Y(u4__abc_49152_n246) );
  INVX1 INVX1_1323 ( .A(u5_burst_cnt_5_), .Y(u5__abc_54027_n248_1) );
  INVX1 INVX1_1324 ( .A(u5_burst_cnt_4_), .Y(u5__abc_54027_n249_1) );
  INVX1 INVX1_1325 ( .A(u5__abc_54027_n252_1), .Y(u5__abc_54027_n253_1) );
  INVX1 INVX1_1326 ( .A(u5_burst_cnt_10_), .Y(u5__abc_54027_n256_1) );
  INVX1 INVX1_1327 ( .A(u5_burst_cnt_9_), .Y(u5__abc_54027_n257) );
  INVX1 INVX1_1328 ( .A(u5_burst_cnt_8_), .Y(u5__abc_54027_n258) );
  INVX1 INVX1_1329 ( .A(u5_burst_cnt_6_), .Y(u5__abc_54027_n260_1) );
  INVX1 INVX1_133 ( .A(\wb_data_i[19] ), .Y(u0_u1__abc_43657_n334) );
  INVX1 INVX1_1330 ( .A(u5_burst_cnt_7_), .Y(u5__abc_54027_n261) );
  INVX1 INVX1_1331 ( .A(u5__abc_54027_n265), .Y(u5_burst_act_rd_FF_INPUT) );
  INVX1 INVX1_1332 ( .A(u5_state_5_), .Y(u5__abc_54027_n268_1) );
  INVX1 INVX1_1333 ( .A(u5_state_3_), .Y(u5__abc_54027_n271) );
  INVX1 INVX1_1334 ( .A(u5_state_4_), .Y(u5__abc_54027_n276) );
  INVX1 INVX1_1335 ( .A(u5_state_2_), .Y(u5__abc_54027_n279) );
  INVX1 INVX1_1336 ( .A(u5_state_1_), .Y(u5__abc_54027_n281) );
  INVX1 INVX1_1337 ( .A(u5_state_0_), .Y(u5__abc_54027_n286) );
  INVX1 INVX1_1338 ( .A(u5__abc_54027_n294), .Y(u5__abc_54027_n295) );
  INVX1 INVX1_1339 ( .A(u5__abc_54027_n297), .Y(u5__abc_54027_n298_1) );
  INVX1 INVX1_134 ( .A(u0_u1__abc_43657_n335), .Y(u0_u1__abc_43657_n336) );
  INVX1 INVX1_1340 ( .A(u5__abc_54027_n301_1), .Y(u5__abc_54027_n302) );
  INVX1 INVX1_1341 ( .A(u5__abc_54027_n304), .Y(u5__abc_54027_n305) );
  INVX1 INVX1_1342 ( .A(u5__abc_54027_n308), .Y(u5__abc_54027_n309) );
  INVX1 INVX1_1343 ( .A(u5_cnt), .Y(u5__abc_54027_n314) );
  INVX1 INVX1_1344 ( .A(u5_dv_r), .Y(u5__abc_54027_n320) );
  INVX1 INVX1_1345 ( .A(u5__abc_54027_n325), .Y(u5__abc_54027_n326) );
  INVX1 INVX1_1346 ( .A(u5_timer_5_), .Y(u5__abc_54027_n327) );
  INVX1 INVX1_1347 ( .A(u5_timer_4_), .Y(u5__abc_54027_n328_1) );
  INVX1 INVX1_1348 ( .A(u5__abc_54027_n333_1), .Y(u5__abc_54027_n334) );
  INVX1 INVX1_1349 ( .A(u5_ir_cnt_1_), .Y(u5__abc_54027_n336) );
  INVX1 INVX1_135 ( .A(\wb_data_i[20] ), .Y(u0_u1__abc_43657_n340) );
  INVX1 INVX1_1350 ( .A(u5_ir_cnt_0_), .Y(u5__abc_54027_n337) );
  INVX1 INVX1_1351 ( .A(u5_ir_cnt_3_), .Y(u5__abc_54027_n339) );
  INVX1 INVX1_1352 ( .A(u5_ir_cnt_2_), .Y(u5__abc_54027_n340) );
  INVX1 INVX1_1353 ( .A(u5__abc_54027_n360), .Y(u5__abc_54027_n361) );
  INVX1 INVX1_1354 ( .A(u5__abc_54027_n362), .Y(u5__abc_54027_n363) );
  INVX1 INVX1_1355 ( .A(u5_pack_le1_d), .Y(u5__abc_54027_n365_1) );
  INVX1 INVX1_1356 ( .A(u5__abc_54027_n366_1), .Y(u5__abc_54027_n367_1) );
  INVX1 INVX1_1357 ( .A(u5__abc_54027_n371), .Y(u5__abc_54027_n372) );
  INVX1 INVX1_1358 ( .A(u5__abc_54027_n375), .Y(u5__abc_54027_n376) );
  INVX1 INVX1_1359 ( .A(u5__abc_54027_n377), .Y(u5__abc_54027_n378) );
  INVX1 INVX1_136 ( .A(u0_u1__abc_43657_n341), .Y(u0_u1__abc_43657_n342) );
  INVX1 INVX1_1360 ( .A(u5__abc_54027_n382), .Y(u5__abc_54027_n383) );
  INVX1 INVX1_1361 ( .A(u5__abc_54027_n384), .Y(u5__abc_54027_n385) );
  INVX1 INVX1_1362 ( .A(u5__abc_54027_n387_1), .Y(u5__abc_54027_n388_1) );
  INVX1 INVX1_1363 ( .A(u5__abc_54027_n390_1), .Y(u5__abc_54027_n391) );
  INVX1 INVX1_1364 ( .A(u5__abc_54027_n270), .Y(u5__abc_54027_n394_1) );
  INVX1 INVX1_1365 ( .A(u5__abc_54027_n296), .Y(u5__abc_54027_n395) );
  INVX1 INVX1_1366 ( .A(u5__abc_54027_n397), .Y(u5__abc_54027_n398) );
  INVX1 INVX1_1367 ( .A(u5__abc_54027_n288_1), .Y(u5__abc_54027_n399) );
  INVX1 INVX1_1368 ( .A(u5__abc_54027_n405), .Y(u5__abc_54027_n406) );
  INVX1 INVX1_1369 ( .A(u5__abc_54027_n416), .Y(u5__abc_54027_n417) );
  INVX1 INVX1_137 ( .A(\wb_data_i[21] ), .Y(u0_u1__abc_43657_n346) );
  INVX1 INVX1_1370 ( .A(u5__abc_54027_n422), .Y(u5__abc_54027_n423) );
  INVX1 INVX1_1371 ( .A(u5__abc_54027_n428), .Y(u5__abc_54027_n429_1) );
  INVX1 INVX1_1372 ( .A(u5__abc_54027_n430_1), .Y(u5__abc_54027_n431) );
  INVX1 INVX1_1373 ( .A(u5__abc_54027_n432_1), .Y(u5__abc_54027_n433_1) );
  INVX1 INVX1_1374 ( .A(u5__abc_54027_n437_1), .Y(u5__abc_54027_n438_1) );
  INVX1 INVX1_1375 ( .A(u5__abc_54027_n445), .Y(u5__abc_54027_n446_1) );
  INVX1 INVX1_1376 ( .A(u5__abc_54027_n447_1), .Y(u5__abc_54027_n448) );
  INVX1 INVX1_1377 ( .A(u5__abc_54027_n347), .Y(u5__abc_54027_n451_1) );
  INVX1 INVX1_1378 ( .A(u5__abc_54027_n452_1), .Y(u5__abc_54027_n453) );
  INVX1 INVX1_1379 ( .A(u5__abc_54027_n354), .Y(u5__abc_54027_n456) );
  INVX1 INVX1_138 ( .A(u0_u1__abc_43657_n347), .Y(u0_u1__abc_43657_n348) );
  INVX1 INVX1_1380 ( .A(u5__abc_54027_n355), .Y(u5__abc_54027_n457) );
  INVX1 INVX1_1381 ( .A(u5__abc_54027_n461_1), .Y(u5__abc_54027_n462) );
  INVX1 INVX1_1382 ( .A(u5_wb_write_go_r), .Y(u5__abc_54027_n467) );
  INVX1 INVX1_1383 ( .A(tms_s_0_), .Y(u5__abc_54027_n468_1) );
  INVX1 INVX1_1384 ( .A(tms_s_2_), .Y(u5__abc_54027_n469) );
  INVX1 INVX1_1385 ( .A(tms_s_1_), .Y(u5__abc_54027_n470_1) );
  INVX1 INVX1_1386 ( .A(u5__abc_54027_n473), .Y(u5__abc_54027_n474) );
  INVX1 INVX1_1387 ( .A(csc_s_3_), .Y(u5__abc_54027_n488) );
  INVX1 INVX1_1388 ( .A(u3_wb_read_go), .Y(u5__abc_54027_n500) );
  INVX1 INVX1_1389 ( .A(u1_wb_write_go), .Y(u5__abc_54027_n501) );
  INVX1 INVX1_139 ( .A(\wb_data_i[22] ), .Y(u0_u1__abc_43657_n352) );
  INVX1 INVX1_1390 ( .A(u5_no_wb_cycle_FF_INPUT), .Y(u5__abc_54027_n503) );
  INVX1 INVX1_1391 ( .A(u5_wb_cycle), .Y(u5__abc_54027_n506) );
  INVX1 INVX1_1392 ( .A(u5__abc_54027_n507), .Y(u5__abc_54027_n508) );
  INVX1 INVX1_1393 ( .A(u5__abc_54027_n509), .Y(u5__abc_54027_n510) );
  INVX1 INVX1_1394 ( .A(rfr_req), .Y(u5__abc_54027_n511) );
  INVX1 INVX1_1395 ( .A(init_req), .Y(u5__abc_54027_n512_1) );
  INVX1 INVX1_1396 ( .A(u5__abc_54027_n522), .Y(u5__abc_54027_n523_1) );
  INVX1 INVX1_1397 ( .A(u5__abc_54027_n529), .Y(u5__abc_54027_n530) );
  INVX1 INVX1_1398 ( .A(u5__abc_54027_n538), .Y(u5__abc_54027_n539) );
  INVX1 INVX1_1399 ( .A(u5_wb_wait_r), .Y(u5__abc_54027_n545_1) );
  INVX1 INVX1_14 ( .A(u0__abc_49347_n4404), .Y(u0__abc_49347_n4405) );
  INVX1 INVX1_140 ( .A(u0_u1__abc_43657_n353), .Y(u0_u1__abc_43657_n354) );
  INVX1 INVX1_1400 ( .A(u5__abc_54027_n550), .Y(u5__abc_54027_n551) );
  INVX1 INVX1_1401 ( .A(u5__abc_54027_n484_1), .Y(u5__abc_54027_n556) );
  INVX1 INVX1_1402 ( .A(u5__abc_54027_n485), .Y(u5__abc_54027_n557) );
  INVX1 INVX1_1403 ( .A(susp_sel), .Y(u5__abc_54027_n560) );
  INVX1 INVX1_1404 ( .A(rfr_ack), .Y(u5__abc_54027_n561) );
  INVX1 INVX1_1405 ( .A(u5__abc_54027_n563_1), .Y(u5__abc_54027_n564) );
  INVX1 INVX1_1406 ( .A(u5__abc_54027_n570), .Y(u5__abc_54027_n571) );
  INVX1 INVX1_1407 ( .A(u5__abc_54027_n573), .Y(u5__abc_54027_n574) );
  INVX1 INVX1_1408 ( .A(csc_s_1_), .Y(u5__abc_54027_n590) );
  INVX1 INVX1_1409 ( .A(u5__abc_54027_n591), .Y(u5__abc_54027_n592_1) );
  INVX1 INVX1_141 ( .A(\wb_data_i[23] ), .Y(u0_u1__abc_43657_n358) );
  INVX1 INVX1_1410 ( .A(u5__abc_54027_n593), .Y(u5__abc_54027_n594) );
  INVX1 INVX1_1411 ( .A(u5__abc_54027_n601_1), .Y(u5__abc_54027_n602) );
  INVX1 INVX1_1412 ( .A(u5__abc_54027_n607), .Y(u5_cmd_3_) );
  INVX1 INVX1_1413 ( .A(u5__abc_54027_n440), .Y(u5__abc_54027_n618) );
  INVX1 INVX1_1414 ( .A(u5_mem_ack_r), .Y(u5__abc_54027_n629) );
  INVX1 INVX1_1415 ( .A(u5__abc_54027_n630_1), .Y(u5__abc_54027_n631) );
  INVX1 INVX1_1416 ( .A(u5_ack_cnt_2_), .Y(u5__abc_54027_n635) );
  INVX1 INVX1_1417 ( .A(u5_ack_cnt_1_), .Y(u5__abc_54027_n636) );
  INVX1 INVX1_1418 ( .A(u5_ack_cnt_0_), .Y(u5__abc_54027_n637) );
  INVX1 INVX1_1419 ( .A(u5__abc_54027_n639), .Y(u5__abc_54027_n640) );
  INVX1 INVX1_142 ( .A(u0_u1__abc_43657_n359), .Y(u0_u1__abc_43657_n360) );
  INVX1 INVX1_1420 ( .A(u5__abc_54027_n641), .Y(u5__abc_54027_n642) );
  INVX1 INVX1_1421 ( .A(u5__abc_54027_n651), .Y(u5__abc_54027_n652) );
  INVX1 INVX1_1422 ( .A(err), .Y(u5__abc_54027_n653) );
  INVX1 INVX1_1423 ( .A(u5__abc_54027_n661), .Y(u5__abc_54027_n662) );
  INVX1 INVX1_1424 ( .A(u5__abc_54027_n489), .Y(u5__abc_54027_n666_1) );
  INVX1 INVX1_1425 ( .A(u5__abc_54027_n667), .Y(u5__abc_54027_n668) );
  INVX1 INVX1_1426 ( .A(u5__abc_54027_n345), .Y(u5__abc_54027_n670) );
  INVX1 INVX1_1427 ( .A(u5__abc_54027_n348), .Y(u5__abc_54027_n671) );
  INVX1 INVX1_1428 ( .A(u5__abc_54027_n352), .Y(u5__abc_54027_n673) );
  INVX1 INVX1_1429 ( .A(u5__abc_54027_n684), .Y(u5__abc_54027_n685_1) );
  INVX1 INVX1_143 ( .A(\wb_data_i[24] ), .Y(u0_u1__abc_43657_n364) );
  INVX1 INVX1_1430 ( .A(u5__abc_54027_n689), .Y(mem_ack) );
  INVX1 INVX1_1431 ( .A(u5_burst_cnt_0_), .Y(u5__abc_54027_n698) );
  INVX1 INVX1_1432 ( .A(u5__abc_54027_n700), .Y(u5__abc_54027_n701) );
  INVX1 INVX1_1433 ( .A(u5__abc_54027_n704), .Y(u5__abc_54027_n715) );
  INVX1 INVX1_1434 ( .A(u5_burst_cnt_1_), .Y(u5__abc_54027_n717) );
  INVX1 INVX1_1435 ( .A(u5_burst_cnt_2_), .Y(u5__abc_54027_n728) );
  INVX1 INVX1_1436 ( .A(u5__abc_54027_n718), .Y(u5__abc_54027_n730) );
  INVX1 INVX1_1437 ( .A(u5__abc_54027_n754), .Y(u5__abc_54027_n761) );
  INVX1 INVX1_1438 ( .A(u5__abc_54027_n763_1), .Y(u5__abc_54027_n770) );
  INVX1 INVX1_1439 ( .A(u5__abc_54027_n772_1), .Y(u5__abc_54027_n779) );
  INVX1 INVX1_144 ( .A(u0_u1__abc_43657_n365), .Y(u0_u1__abc_43657_n366) );
  INVX1 INVX1_1440 ( .A(u5__abc_54027_n789), .Y(u5__abc_54027_n790) );
  INVX1 INVX1_1441 ( .A(u5__abc_54027_n799), .Y(u5__abc_54027_n801_1) );
  INVX1 INVX1_1442 ( .A(u5__abc_54027_n812), .Y(u5__abc_54027_n814) );
  INVX1 INVX1_1443 ( .A(u5__abc_54027_n825), .Y(u5__abc_54027_n826) );
  INVX1 INVX1_1444 ( .A(u5__abc_54027_n828), .Y(u5__abc_54027_n831) );
  INVX1 INVX1_1445 ( .A(u5__abc_54027_n833_1), .Y(u5__abc_54027_n836) );
  INVX1 INVX1_1446 ( .A(u5__abc_54027_n838), .Y(u5__abc_54027_n841) );
  INVX1 INVX1_1447 ( .A(u5__abc_54027_n848), .Y(u5__abc_54027_n849) );
  INVX1 INVX1_1448 ( .A(u5__abc_54027_n852), .Y(u5__abc_54027_n853) );
  INVX1 INVX1_1449 ( .A(u5__abc_54027_n858), .Y(u5__abc_54027_n859) );
  INVX1 INVX1_145 ( .A(\wb_data_i[25] ), .Y(u0_u1__abc_43657_n370) );
  INVX1 INVX1_1450 ( .A(u5__abc_54027_n863), .Y(u5__abc_54027_n864) );
  INVX1 INVX1_1451 ( .A(u5__abc_54027_n867), .Y(u5__abc_54027_n868_1) );
  INVX1 INVX1_1452 ( .A(u5__abc_54027_n869_1), .Y(u5__abc_54027_n870) );
  INVX1 INVX1_1453 ( .A(u5__abc_54027_n871), .Y(u5__abc_54027_n872) );
  INVX1 INVX1_1454 ( .A(u5__abc_54027_n882_1), .Y(u5__abc_54027_n883) );
  INVX1 INVX1_1455 ( .A(u5__abc_54027_n894), .Y(u5__abc_54027_n895_1) );
  INVX1 INVX1_1456 ( .A(u5__abc_54027_n903), .Y(u5__abc_54027_n904) );
  INVX1 INVX1_1457 ( .A(u5__abc_54027_n905_1), .Y(u5__abc_54027_n906_1) );
  INVX1 INVX1_1458 ( .A(u5__abc_54027_n854), .Y(u5__abc_54027_n907) );
  INVX1 INVX1_1459 ( .A(u5__abc_54027_n331), .Y(u5__abc_54027_n921) );
  INVX1 INVX1_146 ( .A(u0_u1__abc_43657_n371), .Y(u0_u1__abc_43657_n372) );
  INVX1 INVX1_1460 ( .A(u5__abc_54027_n862), .Y(u5__abc_54027_n922) );
  INVX1 INVX1_1461 ( .A(tms_s_21_), .Y(u5__abc_54027_n941) );
  INVX1 INVX1_1462 ( .A(tms_s_16_), .Y(u5__abc_54027_n942_1) );
  INVX1 INVX1_1463 ( .A(u5__abc_54027_n873), .Y(u5__abc_54027_n971) );
  INVX1 INVX1_1464 ( .A(u5__abc_54027_n923), .Y(u5__abc_54027_n973) );
  INVX1 INVX1_1465 ( .A(u5_timer_2_), .Y(u5__abc_54027_n975) );
  INVX1 INVX1_1466 ( .A(u5__abc_54027_n966), .Y(u5__abc_54027_n987) );
  INVX1 INVX1_1467 ( .A(u5__abc_54027_n1009), .Y(u5__abc_54027_n1010) );
  INVX1 INVX1_1468 ( .A(u5__abc_54027_n875), .Y(u5__abc_54027_n1017) );
  INVX1 INVX1_1469 ( .A(u5__abc_54027_n976), .Y(u5__abc_54027_n1019) );
  INVX1 INVX1_147 ( .A(\wb_data_i[26] ), .Y(u0_u1__abc_43657_n376) );
  INVX1 INVX1_1470 ( .A(u5__abc_54027_n1018), .Y(u5__abc_54027_n1043) );
  INVX1 INVX1_1471 ( .A(u5__abc_54027_n1042), .Y(u5__abc_54027_n1058_1) );
  INVX1 INVX1_1472 ( .A(u5__abc_54027_n1057), .Y(u5__abc_54027_n1067) );
  INVX1 INVX1_1473 ( .A(u5_timer_6_), .Y(u5__abc_54027_n1069) );
  INVX1 INVX1_1474 ( .A(u5__abc_54027_n1072), .Y(u5__abc_54027_n1079) );
  INVX1 INVX1_1475 ( .A(u5__abc_54027_n1092), .Y(u5__abc_54027_n1093) );
  INVX1 INVX1_1476 ( .A(u5_timer2_0_), .Y(u5__abc_54027_n1095) );
  INVX1 INVX1_1477 ( .A(u5__abc_54027_n1107), .Y(u5__abc_54027_n1108) );
  INVX1 INVX1_1478 ( .A(u5__abc_54027_n1096), .Y(u5__abc_54027_n1119) );
  INVX1 INVX1_1479 ( .A(u5__abc_54027_n1084), .Y(u5__abc_54027_n1142) );
  INVX1 INVX1_148 ( .A(u0_u1__abc_43657_n377), .Y(u0_u1__abc_43657_n378) );
  INVX1 INVX1_1480 ( .A(u5__abc_54027_n1097), .Y(u5__abc_54027_n1145) );
  INVX1 INVX1_1481 ( .A(u5__abc_54027_n1098), .Y(u5__abc_54027_n1165) );
  INVX1 INVX1_1482 ( .A(u5__abc_54027_n1099), .Y(u5__abc_54027_n1191) );
  INVX1 INVX1_1483 ( .A(u5__abc_54027_n1100), .Y(u5__abc_54027_n1209) );
  INVX1 INVX1_1484 ( .A(u5__abc_54027_n1101), .Y(u5__abc_54027_n1222) );
  INVX1 INVX1_1485 ( .A(u5__abc_54027_n1102), .Y(u5__abc_54027_n1234) );
  INVX1 INVX1_1486 ( .A(u5__abc_54027_n1250), .Y(u5__abc_54027_n1251) );
  INVX1 INVX1_1487 ( .A(u5__abc_54027_n1252), .Y(u5__abc_54027_n1253) );
  INVX1 INVX1_1488 ( .A(u5_no_wb_cycle), .Y(u5__abc_54027_n1255) );
  INVX1 INVX1_1489 ( .A(u5__abc_54027_n1261), .Y(u5__abc_54027_n1262) );
  INVX1 INVX1_149 ( .A(\wb_data_i[27] ), .Y(u0_u1__abc_43657_n382) );
  INVX1 INVX1_1490 ( .A(u5__abc_54027_n1270), .Y(u5__abc_54027_n1271) );
  INVX1 INVX1_1491 ( .A(u5__abc_54027_n1281), .Y(u5__abc_54027_n1282) );
  INVX1 INVX1_1492 ( .A(u5__abc_54027_n319), .Y(u5__abc_54027_n1294) );
  INVX1 INVX1_1493 ( .A(u5__abc_54027_n1295), .Y(u5__abc_54027_n1296) );
  INVX1 INVX1_1494 ( .A(u5__abc_54027_n1297), .Y(u5__abc_54027_n1298) );
  INVX1 INVX1_1495 ( .A(u5__abc_54027_n313_1), .Y(u5__abc_54027_n1306) );
  INVX1 INVX1_1496 ( .A(u5__abc_54027_n1308), .Y(u5__abc_54027_n1309) );
  INVX1 INVX1_1497 ( .A(u5__abc_54027_n1313), .Y(u5__abc_54027_n1314) );
  INVX1 INVX1_1498 ( .A(u5__abc_54027_n1316), .Y(u5__abc_54027_n1317) );
  INVX1 INVX1_1499 ( .A(u5__abc_54027_n1323), .Y(u5__abc_54027_n1324) );
  INVX1 INVX1_15 ( .A(\wb_addr_i[5] ), .Y(u0__abc_49347_n4499) );
  INVX1 INVX1_150 ( .A(u0_u1__abc_43657_n383), .Y(u0_u1__abc_43657_n384) );
  INVX1 INVX1_1500 ( .A(u5__abc_54027_n678), .Y(u5__abc_54027_n1326) );
  INVX1 INVX1_1501 ( .A(u5__abc_54027_n1327), .Y(u5__abc_54027_n1328) );
  INVX1 INVX1_1502 ( .A(u5__abc_54027_n1333), .Y(u5__abc_54027_n1334) );
  INVX1 INVX1_1503 ( .A(u5__abc_54027_n1336), .Y(u5__abc_54027_n1337) );
  INVX1 INVX1_1504 ( .A(u5__abc_54027_n1339), .Y(u5__abc_54027_n1340) );
  INVX1 INVX1_1505 ( .A(u5__abc_54027_n1344), .Y(u5__abc_54027_n1345) );
  INVX1 INVX1_1506 ( .A(csc_s_5_bF_buf1), .Y(u5__abc_54027_n1346) );
  INVX1 INVX1_1507 ( .A(u5__abc_54027_n1350), .Y(u5__abc_54027_n1351) );
  INVX1 INVX1_1508 ( .A(u5__abc_54027_n505_1), .Y(u5__abc_54027_n1352) );
  INVX1 INVX1_1509 ( .A(u5__abc_54027_n1354), .Y(u5__abc_54027_n1355) );
  INVX1 INVX1_151 ( .A(\wb_data_i[28] ), .Y(u0_u1__abc_43657_n388) );
  INVX1 INVX1_1510 ( .A(u5__abc_54027_n1356), .Y(u5__abc_54027_n1357) );
  INVX1 INVX1_1511 ( .A(mc_br_r), .Y(u5__abc_54027_n1358) );
  INVX1 INVX1_1512 ( .A(u5__abc_54027_n1364_1), .Y(u5__abc_54027_n1365) );
  INVX1 INVX1_1513 ( .A(u5__abc_54027_n1366), .Y(u5__abc_54027_n1367) );
  INVX1 INVX1_1514 ( .A(u5__abc_54027_n1370), .Y(u5__abc_54027_n1371) );
  INVX1 INVX1_1515 ( .A(u5__abc_54027_n1377), .Y(u5__abc_54027_n1378_1) );
  INVX1 INVX1_1516 ( .A(u5__abc_54027_n1381_1), .Y(u5__abc_54027_n1382) );
  INVX1 INVX1_1517 ( .A(u5__abc_54027_n1384), .Y(u5__abc_54027_n1385) );
  INVX1 INVX1_1518 ( .A(u5__abc_54027_n1387), .Y(u5__abc_54027_n1388) );
  INVX1 INVX1_1519 ( .A(u5__abc_54027_n1393), .Y(u5__abc_54027_n1394) );
  INVX1 INVX1_152 ( .A(u0_u1__abc_43657_n389), .Y(u0_u1__abc_43657_n390) );
  INVX1 INVX1_1520 ( .A(u5__abc_54027_n646), .Y(u5__abc_54027_n1401) );
  INVX1 INVX1_1521 ( .A(u5__abc_54027_n1407_1), .Y(u5__abc_54027_n1408) );
  INVX1 INVX1_1522 ( .A(u5__abc_54027_n1409), .Y(u5__abc_54027_n1410) );
  INVX1 INVX1_1523 ( .A(u5__abc_54027_n1416), .Y(u5__abc_54027_n1417) );
  INVX1 INVX1_1524 ( .A(u5__abc_54027_n1422), .Y(u5__abc_54027_n1423) );
  INVX1 INVX1_1525 ( .A(u5__abc_54027_n491), .Y(u5__abc_54027_n1424) );
  INVX1 INVX1_1526 ( .A(u5__abc_54027_n587), .Y(u5__abc_54027_n1425) );
  INVX1 INVX1_1527 ( .A(u5__abc_54027_n1427), .Y(u5__abc_54027_n1428) );
  INVX1 INVX1_1528 ( .A(mc_ack_r), .Y(u5__abc_54027_n1433) );
  INVX1 INVX1_1529 ( .A(u5__abc_54027_n1434), .Y(u5__abc_54027_n1435) );
  INVX1 INVX1_153 ( .A(\wb_data_i[29] ), .Y(u0_u1__abc_43657_n394) );
  INVX1 INVX1_1530 ( .A(u5__abc_54027_n1441), .Y(u5__abc_54027_n1442) );
  INVX1 INVX1_1531 ( .A(u5__abc_54027_n1445_1), .Y(u5__abc_54027_n1446) );
  INVX1 INVX1_1532 ( .A(u5__abc_54027_n1450_1), .Y(u5__abc_54027_n1451) );
  INVX1 INVX1_1533 ( .A(u5__abc_54027_n1453), .Y(u5__abc_54027_n1454_1) );
  INVX1 INVX1_1534 ( .A(u5__abc_54027_n1459), .Y(u5__abc_54027_n1460) );
  INVX1 INVX1_1535 ( .A(u5__abc_54027_n660), .Y(u5__abc_54027_n1467_1) );
  INVX1 INVX1_1536 ( .A(u5__abc_54027_n1470), .Y(u5__abc_54027_n1471) );
  INVX1 INVX1_1537 ( .A(u5__abc_54027_n1472), .Y(u5__abc_54027_n1473) );
  INVX1 INVX1_1538 ( .A(u5__abc_54027_n1476_1), .Y(u5__abc_54027_n1477) );
  INVX1 INVX1_1539 ( .A(u5__abc_54027_n1481), .Y(u5__abc_54027_n1482) );
  INVX1 INVX1_154 ( .A(u0_u1__abc_43657_n395), .Y(u0_u1__abc_43657_n396) );
  INVX1 INVX1_1540 ( .A(u5__abc_54027_n1484), .Y(u5__abc_54027_n1485) );
  INVX1 INVX1_1541 ( .A(u5__abc_54027_n1330), .Y(u5__abc_54027_n1489) );
  INVX1 INVX1_1542 ( .A(u5__abc_54027_n1490), .Y(u5__abc_54027_n1491_1) );
  INVX1 INVX1_1543 ( .A(u5__abc_54027_n598), .Y(u5__abc_54027_n1494) );
  INVX1 INVX1_1544 ( .A(u5__abc_54027_n1421), .Y(u5__abc_54027_n1495) );
  INVX1 INVX1_1545 ( .A(u5_lookup_ready2), .Y(u5__abc_54027_n1514) );
  INVX1 INVX1_1546 ( .A(u5__abc_54027_n1528), .Y(u5__abc_54027_n1529) );
  INVX1 INVX1_1547 ( .A(u5__abc_54027_n1518), .Y(u5__abc_54027_n1530) );
  INVX1 INVX1_1548 ( .A(u5__abc_54027_n1532), .Y(u5__abc_54027_n1533_1) );
  INVX1 INVX1_1549 ( .A(u5__abc_54027_n1535), .Y(u5__abc_54027_n1536) );
  INVX1 INVX1_155 ( .A(\wb_data_i[30] ), .Y(u0_u1__abc_43657_n400) );
  INVX1 INVX1_1550 ( .A(u5__abc_54027_n1545), .Y(u5__abc_41027_n1845) );
  INVX1 INVX1_1551 ( .A(u5__abc_54027_n1342), .Y(u5__abc_54027_n1547_1) );
  INVX1 INVX1_1552 ( .A(u5_ap_en), .Y(u5__abc_54027_n1551_1) );
  INVX1 INVX1_1553 ( .A(u5__abc_54027_n1552_1), .Y(u5__abc_54027_n1553) );
  INVX1 INVX1_1554 ( .A(u5__abc_54027_n615), .Y(u5__abc_54027_n1559) );
  INVX1 INVX1_1555 ( .A(u5__abc_54027_n1568), .Y(u5__abc_54027_n1569) );
  INVX1 INVX1_1556 ( .A(row_same), .Y(u5__abc_54027_n1573_1) );
  INVX1 INVX1_1557 ( .A(u5__abc_54027_n1577), .Y(u5__abc_54027_n1578) );
  INVX1 INVX1_1558 ( .A(u5__abc_54027_n1581), .Y(u5__abc_54027_n1582) );
  INVX1 INVX1_1559 ( .A(u5__abc_54027_n1585), .Y(u5__abc_54027_n1586) );
  INVX1 INVX1_156 ( .A(u0_u1__abc_43657_n401), .Y(u0_u1__abc_43657_n402) );
  INVX1 INVX1_1560 ( .A(u5__abc_54027_n1596), .Y(u5__abc_54027_n1597) );
  INVX1 INVX1_1561 ( .A(u5__abc_54027_n1600), .Y(u5__abc_54027_n1601) );
  INVX1 INVX1_1562 ( .A(u5__abc_54027_n1602), .Y(u5__abc_54027_n1603) );
  INVX1 INVX1_1563 ( .A(u5_ir_cnt_done), .Y(u5__abc_54027_n1604) );
  INVX1 INVX1_1564 ( .A(u5__abc_54027_n1605), .Y(u5__abc_54027_n1606) );
  INVX1 INVX1_1565 ( .A(u5__abc_54027_n1615), .Y(u5__abc_54027_n1616) );
  INVX1 INVX1_1566 ( .A(u5__abc_54027_n1630), .Y(u5__abc_54027_n1631) );
  INVX1 INVX1_1567 ( .A(u5__abc_54027_n1634), .Y(u5__abc_54027_n1635) );
  INVX1 INVX1_1568 ( .A(u5__abc_54027_n1643), .Y(u5__abc_54027_n1644) );
  INVX1 INVX1_1569 ( .A(u5__abc_54027_n1647), .Y(u5__abc_54027_n1648) );
  INVX1 INVX1_157 ( .A(\wb_data_i[31] ), .Y(u0_u1__abc_43657_n406) );
  INVX1 INVX1_1570 ( .A(u5__abc_54027_n475_1), .Y(u5__abc_54027_n1649) );
  INVX1 INVX1_1571 ( .A(u5__abc_54027_n1550), .Y(u5__abc_54027_n1659) );
  INVX1 INVX1_1572 ( .A(u5__abc_54027_n1662), .Y(u5__abc_54027_n1663) );
  INVX1 INVX1_1573 ( .A(u5__abc_54027_n1664), .Y(u5__abc_54027_n1665) );
  INVX1 INVX1_1574 ( .A(u5__abc_54027_n1667), .Y(u5__abc_54027_n1668) );
  INVX1 INVX1_1575 ( .A(u5__abc_54027_n1669), .Y(u5__abc_54027_n1670) );
  INVX1 INVX1_1576 ( .A(u5__abc_54027_n476), .Y(u5__abc_54027_n1672) );
  INVX1 INVX1_1577 ( .A(u5__abc_54027_n1678), .Y(u5__abc_54027_n1679) );
  INVX1 INVX1_1578 ( .A(u5__abc_54027_n1680), .Y(u5__abc_54027_n1681) );
  INVX1 INVX1_1579 ( .A(u5__abc_54027_n1683), .Y(u5__abc_54027_n1684) );
  INVX1 INVX1_158 ( .A(u0_u1__abc_43657_n407), .Y(u0_u1__abc_43657_n408) );
  INVX1 INVX1_1580 ( .A(u5__abc_54027_n1687), .Y(u5__abc_54027_n1688) );
  INVX1 INVX1_1581 ( .A(u5__abc_54027_n1704), .Y(u5__abc_54027_n1705) );
  INVX1 INVX1_1582 ( .A(u5__abc_54027_n1710), .Y(u5__abc_54027_n1711) );
  INVX1 INVX1_1583 ( .A(u5_resume_req_r), .Y(u5__abc_54027_n1712) );
  INVX1 INVX1_1584 ( .A(u5__abc_54027_n1715), .Y(u5__abc_54027_n1716) );
  INVX1 INVX1_1585 ( .A(u5__abc_54027_n1564), .Y(u5__abc_54027_n1726) );
  INVX1 INVX1_1586 ( .A(u5__abc_54027_n1729), .Y(u5__abc_54027_n1730) );
  INVX1 INVX1_1587 ( .A(u5__abc_54027_n1742), .Y(u5__abc_54027_n1743) );
  INVX1 INVX1_1588 ( .A(u5__abc_54027_n1335), .Y(u5__abc_54027_n1750) );
  INVX1 INVX1_1589 ( .A(u5__abc_54027_n1752), .Y(u5__abc_54027_n1753) );
  INVX1 INVX1_159 ( .A(u0_u1_addr_r_2_), .Y(u0_u1__abc_43657_n411) );
  INVX1 INVX1_1590 ( .A(u5__abc_54027_n620_1), .Y(u5__abc_54027_n1755) );
  INVX1 INVX1_1591 ( .A(u5__abc_54027_n1772), .Y(u5__abc_54027_n1773) );
  INVX1 INVX1_1592 ( .A(u5__abc_54027_n1782), .Y(u5__abc_54027_n1783) );
  INVX1 INVX1_1593 ( .A(u5__abc_54027_n1689), .Y(u5__abc_54027_n1786) );
  INVX1 INVX1_1594 ( .A(u5__abc_54027_n1798), .Y(u5__abc_54027_n1799) );
  INVX1 INVX1_1595 ( .A(u5__abc_54027_n1807), .Y(u5__abc_41027_n1849) );
  INVX1 INVX1_1596 ( .A(u5__abc_54027_n1809), .Y(u5__abc_54027_n1810) );
  INVX1 INVX1_1597 ( .A(u5__abc_54027_n1821), .Y(u5__abc_41027_n1850) );
  INVX1 INVX1_1598 ( .A(u5__abc_54027_n1653), .Y(u5__abc_54027_n1829) );
  INVX1 INVX1_1599 ( .A(u5__abc_54027_n1855), .Y(u5__abc_54027_n1856) );
  INVX1 INVX1_16 ( .A(\wb_addr_i[4] ), .Y(u0__abc_49347_n4500) );
  INVX1 INVX1_160 ( .A(u0_u1__abc_43657_n414), .Y(u0_u1__abc_43657_n415) );
  INVX1 INVX1_1600 ( .A(u5__abc_54027_n1493), .Y(u5__abc_54027_n1868) );
  INVX1 INVX1_1601 ( .A(lmr_req), .Y(u5__abc_54027_n1876) );
  INVX1 INVX1_1602 ( .A(u5_susp_req_r), .Y(u5__abc_54027_n1877) );
  INVX1 INVX1_1603 ( .A(u5__abc_54027_n1503), .Y(u5__abc_54027_n1883) );
  INVX1 INVX1_1604 ( .A(u5__abc_54027_n1875), .Y(u5__abc_54027_n1904) );
  INVX1 INVX1_1605 ( .A(u5__abc_54027_n450), .Y(u5__abc_54027_n1908) );
  INVX1 INVX1_1606 ( .A(u5__abc_54027_n386_1), .Y(u5__abc_54027_n1913) );
  INVX1 INVX1_1607 ( .A(u5__abc_54027_n1839), .Y(u5__abc_54027_n1921) );
  INVX1 INVX1_1608 ( .A(u5__abc_54027_n521), .Y(u5__abc_54027_n1925) );
  INVX1 INVX1_1609 ( .A(u5__abc_54027_n1690), .Y(u5__abc_54027_n1933) );
  INVX1 INVX1_161 ( .A(u0_u1__abc_43657_n419), .Y(u0_u1__abc_43657_n420) );
  INVX1 INVX1_1610 ( .A(u5__abc_54027_n1937), .Y(u5__abc_54027_n1938) );
  INVX1 INVX1_1611 ( .A(u5__abc_54027_n1865), .Y(u5__abc_54027_n1953) );
  INVX1 INVX1_1612 ( .A(u5__abc_54027_n1870), .Y(u5__abc_54027_n1954) );
  INVX1 INVX1_1613 ( .A(u5__abc_54027_n1549), .Y(u5__abc_54027_n1960) );
  INVX1 INVX1_1614 ( .A(u5__abc_54027_n1708), .Y(u5__abc_54027_n1961) );
  INVX1 INVX1_1615 ( .A(u5__abc_54027_n344_1), .Y(u5__abc_54027_n1970) );
  INVX1 INVX1_1616 ( .A(u5__abc_54027_n619), .Y(u5__abc_54027_n1974) );
  INVX1 INVX1_1617 ( .A(u5__abc_54027_n1456), .Y(u5__abc_54027_n1976) );
  INVX1 INVX1_1618 ( .A(u5__abc_54027_n1474), .Y(u5__abc_54027_n1977) );
  INVX1 INVX1_1619 ( .A(u5__abc_54027_n460), .Y(u5__abc_54027_n1980) );
  INVX1 INVX1_162 ( .A(u0_u1__abc_43657_n424), .Y(u0_u1__abc_43657_n425) );
  INVX1 INVX1_1620 ( .A(u5__abc_54027_n1990), .Y(u5__abc_54027_n1992) );
  INVX1 INVX1_1621 ( .A(u5__abc_54027_n1103), .Y(u5__abc_54027_n2000) );
  INVX1 INVX1_1622 ( .A(u5__abc_54027_n1369), .Y(u5__abc_54027_n2004) );
  INVX1 INVX1_1623 ( .A(not_mem_cyc), .Y(u5__abc_54027_n2012) );
  INVX1 INVX1_1624 ( .A(u5__abc_54027_n1948), .Y(u5__abc_54027_n2018) );
  INVX1 INVX1_1625 ( .A(u5_rsts), .Y(u5__abc_54027_n1573) );
  INVX1 INVX1_1626 ( .A(u6__abc_56056_n132), .Y(u6__abc_56056_n133) );
  INVX1 INVX1_1627 ( .A(par_err), .Y(u6__abc_56056_n134) );
  INVX1 INVX1_1628 ( .A(u0_wp_err), .Y(u6__abc_56056_n135_1) );
  INVX1 INVX1_1629 ( .A(err), .Y(u6__abc_56056_n136) );
  INVX1 INVX1_163 ( .A(u0_u1__abc_43657_n429), .Y(u0_u1__abc_43657_n430) );
  INVX1 INVX1_1630 ( .A(\wb_addr_i[31] ), .Y(u6__abc_56056_n140_1) );
  INVX1 INVX1_1631 ( .A(\wb_addr_i[30] ), .Y(u6__abc_56056_n141_1) );
  INVX1 INVX1_1632 ( .A(\wb_addr_i[29] ), .Y(u6__abc_56056_n142_1) );
  INVX1 INVX1_1633 ( .A(_auto_iopadmap_cc_313_execute_56356), .Y(u6__abc_56056_n148_1) );
  INVX1 INVX1_1634 ( .A(u1_wr_hold), .Y(u6__abc_56056_n253) );
  INVX1 INVX1_1635 ( .A(wb_we_i), .Y(u6__abc_56056_n256) );
  INVX1 INVX1_1636 ( .A(u6_rmw_r), .Y(u6__abc_56056_n260) );
  INVX1 INVX1_1637 ( .A(u6_rmw_r_FF_INPUT), .Y(u6__abc_56056_n261) );
  INVX1 INVX1_1638 ( .A(wb_stb_i_bF_buf1), .Y(u6__abc_56056_n270) );
  INVX1 INVX1_1639 ( .A(u6_read_go_r), .Y(u6__abc_56056_n275) );
  INVX1 INVX1_164 ( .A(u0_u1__abc_43657_n434), .Y(u0_u1__abc_43657_n435) );
  INVX1 INVX1_1640 ( .A(u6_write_go_r), .Y(u6__abc_56056_n276) );
  INVX1 INVX1_1641 ( .A(_auto_iopadmap_cc_313_execute_56391), .Y(u6__abc_56056_n280) );
  INVX1 INVX1_1642 ( .A(u6__abc_56056_n139_1), .Y(u6__abc_56056_n284) );
  INVX1 INVX1_1643 ( .A(u7_mc_dqm_r2_0_), .Y(u7__abc_47535_n75_1) );
  INVX1 INVX1_1644 ( .A(data_oe), .Y(u7__abc_47535_n77_1) );
  INVX1 INVX1_1645 ( .A(u5_wb_cycle), .Y(u7__abc_47535_n78) );
  INVX1 INVX1_1646 ( .A(u7_mc_dqm_r2_1_), .Y(u7__abc_47535_n83_1) );
  INVX1 INVX1_1647 ( .A(u7_mc_dqm_r2_2_), .Y(u7__abc_47535_n86_1) );
  INVX1 INVX1_1648 ( .A(u7_mc_dqm_r2_3_), .Y(u7__abc_47535_n89_1) );
  INVX1 INVX1_1649 ( .A(u7__abc_47535_n92_1), .Y(u7__abc_47535_n94_1) );
  INVX1 INVX1_165 ( .A(u0_u1__abc_43657_n439), .Y(u0_u1__abc_43657_n440) );
  INVX1 INVX1_1650 ( .A(cs_0_), .Y(u7__abc_47535_n108) );
  INVX1 INVX1_1651 ( .A(u7__abc_47535_n110), .Y(u7__abc_47535_n111) );
  INVX1 INVX1_1652 ( .A(cs_need_rfr_0_), .Y(u7__abc_47535_n115) );
  INVX1 INVX1_1653 ( .A(cs_1_), .Y(u7__abc_47535_n119) );
  INVX1 INVX1_1654 ( .A(u7__abc_47535_n121), .Y(u7__abc_47535_n122) );
  INVX1 INVX1_1655 ( .A(cs_need_rfr_1_), .Y(u7__abc_47535_n125) );
  INVX1 INVX1_1656 ( .A(cs_2_), .Y(u7__abc_47535_n129) );
  INVX1 INVX1_1657 ( .A(u7__abc_47535_n131), .Y(u7__abc_47535_n132) );
  INVX1 INVX1_1658 ( .A(cs_need_rfr_2_), .Y(u7__abc_47535_n135) );
  INVX1 INVX1_1659 ( .A(cs_3_), .Y(u7__abc_47535_n139) );
  INVX1 INVX1_166 ( .A(u0_u1__abc_43657_n444), .Y(u0_u1__abc_43657_n445) );
  INVX1 INVX1_1660 ( .A(u7__abc_47535_n141), .Y(u7__abc_47535_n142) );
  INVX1 INVX1_1661 ( .A(cs_need_rfr_3_), .Y(u7__abc_47535_n145) );
  INVX1 INVX1_1662 ( .A(cs_4_), .Y(u7__abc_47535_n149) );
  INVX1 INVX1_1663 ( .A(u7__abc_47535_n151), .Y(u7__abc_47535_n152) );
  INVX1 INVX1_1664 ( .A(cs_need_rfr_4_), .Y(u7__abc_47535_n155) );
  INVX1 INVX1_1665 ( .A(cs_5_), .Y(u7__abc_47535_n159) );
  INVX1 INVX1_1666 ( .A(u7__abc_47535_n161), .Y(u7__abc_47535_n162) );
  INVX1 INVX1_1667 ( .A(cs_need_rfr_5_), .Y(u7__abc_47535_n165) );
  INVX1 INVX1_1668 ( .A(cs_6_), .Y(u7__abc_47535_n169) );
  INVX1 INVX1_1669 ( .A(u7__abc_47535_n171), .Y(u7__abc_47535_n172) );
  INVX1 INVX1_167 ( .A(u0_u1__abc_43657_n449), .Y(u0_u1__abc_43657_n450) );
  INVX1 INVX1_1670 ( .A(cs_need_rfr_6_), .Y(u7__abc_47535_n175) );
  INVX1 INVX1_1671 ( .A(cs_7_), .Y(u7__abc_47535_n179) );
  INVX1 INVX1_1672 ( .A(u7__abc_47535_n181), .Y(u7__abc_47535_n182) );
  INVX1 INVX1_1673 ( .A(cs_need_rfr_7_), .Y(u7__abc_47535_n185) );
  INVX1 INVX1_1674 ( .A(mc_adsc_d), .Y(u7_mc_adsc__FF_INPUT) );
  INVX1 INVX1_1675 ( .A(mc_adv_d), .Y(u7_mc_adv__FF_INPUT) );
  INVX1 INVX1_1676 ( .A(fs), .Y(u7__abc_47535_n191) );
  INVX1 INVX1_1677 ( .A(_auto_iopadmap_cc_313_execute_56354), .Y(u7__abc_47535_n192) );
  INVX1 INVX1_1678 ( .A(susp_sel), .Y(u7__abc_47535_n194) );
  INVX1 INVX1_168 ( .A(u0_u1__abc_43657_n454), .Y(u0_u1__abc_43657_n455) );
  INVX1 INVX1_169 ( .A(u0_u1__abc_43657_n459), .Y(u0_u1__abc_43657_n460) );
  INVX1 INVX1_17 ( .A(\wb_addr_i[6] ), .Y(u0__abc_49347_n4502) );
  INVX1 INVX1_170 ( .A(u0_u1__abc_43657_n464), .Y(u0_u1__abc_43657_n465) );
  INVX1 INVX1_171 ( .A(u0_u1__abc_43657_n469), .Y(u0_u1__abc_43657_n470) );
  INVX1 INVX1_172 ( .A(u0_u1__abc_43657_n474), .Y(u0_u1__abc_43657_n475) );
  INVX1 INVX1_173 ( .A(u0_u1__abc_43657_n479), .Y(u0_u1__abc_43657_n480) );
  INVX1 INVX1_174 ( .A(u0_u1__abc_43657_n484), .Y(u0_u1__abc_43657_n485) );
  INVX1 INVX1_175 ( .A(u0_u1__abc_43657_n489), .Y(u0_u1__abc_43657_n490) );
  INVX1 INVX1_176 ( .A(u0_u1__abc_43657_n494), .Y(u0_u1__abc_43657_n495) );
  INVX1 INVX1_177 ( .A(u0_u1__abc_43657_n499), .Y(u0_u1__abc_43657_n500) );
  INVX1 INVX1_178 ( .A(u0_u1__abc_43657_n504), .Y(u0_u1__abc_43657_n505) );
  INVX1 INVX1_179 ( .A(u0_u1__abc_43657_n509), .Y(u0_u1__abc_43657_n510) );
  INVX1 INVX1_18 ( .A(\wb_addr_i[3] ), .Y(u0__abc_49347_n4503) );
  INVX1 INVX1_180 ( .A(u0_u1__abc_43657_n514), .Y(u0_u1__abc_43657_n515) );
  INVX1 INVX1_181 ( .A(u0_u1__abc_43657_n519), .Y(u0_u1__abc_43657_n520) );
  INVX1 INVX1_182 ( .A(u0_u1__abc_43657_n524), .Y(u0_u1__abc_43657_n525) );
  INVX1 INVX1_183 ( .A(u0_u1__abc_43657_n529), .Y(u0_u1__abc_43657_n530) );
  INVX1 INVX1_184 ( .A(u0_u1__abc_43657_n534), .Y(u0_u1__abc_43657_n535) );
  INVX1 INVX1_185 ( .A(u0_u1__abc_43657_n539), .Y(u0_u1__abc_43657_n540) );
  INVX1 INVX1_186 ( .A(u0_u1__abc_43657_n544), .Y(u0_u1__abc_43657_n545) );
  INVX1 INVX1_187 ( .A(u0_u1__abc_43657_n549), .Y(u0_u1__abc_43657_n550) );
  INVX1 INVX1_188 ( .A(u0_u1__abc_43657_n554), .Y(u0_u1__abc_43657_n555) );
  INVX1 INVX1_189 ( .A(u0_u1__abc_43657_n559), .Y(u0_u1__abc_43657_n560) );
  INVX1 INVX1_19 ( .A(\wb_addr_i[2] ), .Y(u0__abc_49347_n4504) );
  INVX1 INVX1_190 ( .A(u0_u1__abc_43657_n564), .Y(u0_u1__abc_43657_n565) );
  INVX1 INVX1_191 ( .A(u0_u1__abc_43657_n569), .Y(u0_u1__abc_43657_n570) );
  INVX1 INVX1_192 ( .A(u0_u1__abc_43657_n575), .Y(u0_u1__abc_43657_n576) );
  INVX1 INVX1_193 ( .A(u0_u1__abc_43657_n579), .Y(u0_u1__abc_43657_n580) );
  INVX1 INVX1_194 ( .A(wb_addr_i_23_bF_buf1), .Y(u0_u1__abc_43657_n583) );
  INVX1 INVX1_195 ( .A(u0_u1__abc_43657_n585), .Y(u0_u1__abc_43657_n586) );
  INVX1 INVX1_196 ( .A(u0_u1__abc_43657_n578), .Y(u0_u1__abc_43657_n587) );
  INVX1 INVX1_197 ( .A(u0_u1__abc_43657_n592), .Y(u0_u1__abc_43657_n593) );
  INVX1 INVX1_198 ( .A(u0_u1__abc_43657_n596), .Y(u0_u1__abc_43657_n597) );
  INVX1 INVX1_199 ( .A(wb_addr_i_25_bF_buf0), .Y(u0_u1__abc_43657_n600) );
  INVX1 INVX1_2 ( .A(lmr_ack), .Y(_abc_55805_n239_1) );
  INVX1 INVX1_20 ( .A(u0__abc_49347_n4511_bF_buf3), .Y(u0__abc_49347_n4545) );
  INVX1 INVX1_200 ( .A(u0_u1__abc_43657_n601), .Y(u0_u1__abc_43657_n602) );
  INVX1 INVX1_201 ( .A(u0_u1__abc_43657_n595), .Y(u0_u1__abc_43657_n603) );
  INVX1 INVX1_202 ( .A(u0_u1__abc_43657_n608), .Y(u0_u1__abc_43657_n609) );
  INVX1 INVX1_203 ( .A(u0_u1__abc_43657_n610), .Y(u0_u1__abc_43657_n611) );
  INVX1 INVX1_204 ( .A(u0_u1__abc_43657_n612), .Y(u0_u1__abc_43657_n615) );
  INVX1 INVX1_205 ( .A(u0_u1__abc_43657_n619), .Y(u0_u1__abc_43657_n620) );
  INVX1 INVX1_206 ( .A(u0_u1__abc_43657_n623), .Y(u0_u1__abc_43657_n624) );
  INVX1 INVX1_207 ( .A(u0_u1__abc_43657_n628), .Y(u0_u1__abc_43657_n629) );
  INVX1 INVX1_208 ( .A(u0_u1__abc_43657_n622), .Y(u0_u1__abc_43657_n631) );
  INVX1 INVX1_209 ( .A(u0_u1__abc_43657_n627), .Y(u0_u1__abc_43657_n635) );
  INVX1 INVX1_21 ( .A(u0__abc_49347_n4535_bF_buf3), .Y(u0__abc_49347_n4546) );
  INVX1 INVX1_210 ( .A(u0_u1__abc_43657_n573), .Y(u0_u1__abc_43657_n641) );
  INVX1 INVX1_211 ( .A(u0_init_ack1), .Y(u0_u1__abc_43657_n644) );
  INVX1 INVX1_212 ( .A(u0_u1_inited), .Y(u0_u1__abc_43657_n646) );
  INVX1 INVX1_213 ( .A(u0_u2_addr_r_2_), .Y(u0_u2__abc_44109_n201_1) );
  INVX1 INVX1_214 ( .A(u0_u2__abc_44109_n204_1), .Y(u0_u2__abc_44109_n205_1) );
  INVX1 INVX1_215 ( .A(u0_u2__abc_44109_n469), .Y(u0_u2__abc_44109_n470) );
  INVX1 INVX1_216 ( .A(u0_u2__abc_44109_n471), .Y(u0_u2__abc_44109_n473) );
  INVX1 INVX1_217 ( .A(u0_lmr_ack2), .Y(u0_u2__abc_44109_n474) );
  INVX1 INVX1_218 ( .A(u0_init_ack2), .Y(u0_u2__abc_44109_n478) );
  INVX1 INVX1_219 ( .A(u0_u2_inited), .Y(u0_u2__abc_44109_n480) );
  INVX1 INVX1_22 ( .A(u0__abc_49347_n4528_bF_buf3), .Y(u0__abc_49347_n4548) );
  INVX1 INVX1_220 ( .A(u0_u2__abc_44109_n488), .Y(u0_u2__abc_44109_n489) );
  INVX1 INVX1_221 ( .A(u0_u2__abc_44109_n492), .Y(u0_u2__abc_44109_n493) );
  INVX1 INVX1_222 ( .A(wb_addr_i_23_bF_buf3), .Y(u0_u2__abc_44109_n496) );
  INVX1 INVX1_223 ( .A(u0_u2__abc_44109_n498), .Y(u0_u2__abc_44109_n499) );
  INVX1 INVX1_224 ( .A(u0_u2__abc_44109_n491), .Y(u0_u2__abc_44109_n500) );
  INVX1 INVX1_225 ( .A(u0_u2__abc_44109_n505), .Y(u0_u2__abc_44109_n506) );
  INVX1 INVX1_226 ( .A(u0_u2__abc_44109_n509), .Y(u0_u2__abc_44109_n510) );
  INVX1 INVX1_227 ( .A(wb_addr_i_25_bF_buf2), .Y(u0_u2__abc_44109_n513) );
  INVX1 INVX1_228 ( .A(u0_u2__abc_44109_n514), .Y(u0_u2__abc_44109_n515) );
  INVX1 INVX1_229 ( .A(u0_u2__abc_44109_n508), .Y(u0_u2__abc_44109_n516) );
  INVX1 INVX1_23 ( .A(u0__abc_49347_n4537_bF_buf3), .Y(u0__abc_49347_n4549) );
  INVX1 INVX1_230 ( .A(u0_u2__abc_44109_n521), .Y(u0_u2__abc_44109_n522) );
  INVX1 INVX1_231 ( .A(u0_u2__abc_44109_n523), .Y(u0_u2__abc_44109_n524) );
  INVX1 INVX1_232 ( .A(u0_u2__abc_44109_n525), .Y(u0_u2__abc_44109_n528) );
  INVX1 INVX1_233 ( .A(u0_u2__abc_44109_n532), .Y(u0_u2__abc_44109_n533) );
  INVX1 INVX1_234 ( .A(u0_u2__abc_44109_n536), .Y(u0_u2__abc_44109_n537) );
  INVX1 INVX1_235 ( .A(u0_u2__abc_44109_n541), .Y(u0_u2__abc_44109_n542) );
  INVX1 INVX1_236 ( .A(u0_u2__abc_44109_n535), .Y(u0_u2__abc_44109_n544) );
  INVX1 INVX1_237 ( .A(u0_u2__abc_44109_n540), .Y(u0_u2__abc_44109_n548) );
  INVX1 INVX1_238 ( .A(u0_u2__abc_44109_n486), .Y(u0_u2__abc_44109_n554) );
  INVX1 INVX1_239 ( .A(u0_u3_addr_r_2_), .Y(u0_u3__abc_44466_n206_1) );
  INVX1 INVX1_24 ( .A(u0__abc_49347_n4507_bF_buf2), .Y(u0__abc_49347_n4552) );
  INVX1 INVX1_240 ( .A(u0_u3_addr_r_6_), .Y(u0_u3__abc_44466_n207) );
  INVX1 INVX1_241 ( .A(u0_u3_addr_r_4_), .Y(u0_u3__abc_44466_n208_1) );
  INVX1 INVX1_242 ( .A(\wb_data_i[0] ), .Y(u0_u3__abc_44466_n215_1) );
  INVX1 INVX1_243 ( .A(u0_u3__abc_44466_n216), .Y(u0_u3__abc_44466_n217_1) );
  INVX1 INVX1_244 ( .A(\wb_data_i[1] ), .Y(u0_u3__abc_44466_n225) );
  INVX1 INVX1_245 ( .A(u0_u3__abc_44466_n226_1), .Y(u0_u3__abc_44466_n227_1) );
  INVX1 INVX1_246 ( .A(\wb_data_i[2] ), .Y(u0_u3__abc_44466_n232_1) );
  INVX1 INVX1_247 ( .A(u0_u3__abc_44466_n233_1), .Y(u0_u3__abc_44466_n234) );
  INVX1 INVX1_248 ( .A(\wb_data_i[4] ), .Y(u0_u3__abc_44466_n244_1) );
  INVX1 INVX1_249 ( .A(u0_u3__abc_44466_n245_1), .Y(u0_u3__abc_44466_n246) );
  INVX1 INVX1_25 ( .A(u0__abc_49347_n4516_bF_buf3), .Y(u0__abc_49347_n4553) );
  INVX1 INVX1_250 ( .A(\wb_data_i[5] ), .Y(u0_u3__abc_44466_n252_1) );
  INVX1 INVX1_251 ( .A(u0_u3__abc_44466_n253), .Y(u0_u3__abc_44466_n254_1) );
  INVX1 INVX1_252 ( .A(u0_u3__abc_44466_n494), .Y(u0_u3__abc_44466_n495) );
  INVX1 INVX1_253 ( .A(u0_u3__abc_44466_n496), .Y(u0_u3__abc_44466_n498) );
  INVX1 INVX1_254 ( .A(u0_lmr_ack3), .Y(u0_u3__abc_44466_n499) );
  INVX1 INVX1_255 ( .A(u0_init_ack3), .Y(u0_u3__abc_44466_n503) );
  INVX1 INVX1_256 ( .A(u0_u3_inited), .Y(u0_u3__abc_44466_n505) );
  INVX1 INVX1_257 ( .A(u0_u3__abc_44466_n513), .Y(u0_u3__abc_44466_n514) );
  INVX1 INVX1_258 ( .A(u0_u3__abc_44466_n517), .Y(u0_u3__abc_44466_n518) );
  INVX1 INVX1_259 ( .A(wb_addr_i_23_bF_buf1), .Y(u0_u3__abc_44466_n521) );
  INVX1 INVX1_26 ( .A(u0__abc_49347_n4519_bF_buf3), .Y(u0__abc_49347_n4555) );
  INVX1 INVX1_260 ( .A(u0_u3__abc_44466_n523), .Y(u0_u3__abc_44466_n524) );
  INVX1 INVX1_261 ( .A(u0_u3__abc_44466_n516), .Y(u0_u3__abc_44466_n525) );
  INVX1 INVX1_262 ( .A(u0_u3__abc_44466_n530), .Y(u0_u3__abc_44466_n531) );
  INVX1 INVX1_263 ( .A(u0_u3__abc_44466_n534), .Y(u0_u3__abc_44466_n535) );
  INVX1 INVX1_264 ( .A(wb_addr_i_25_bF_buf0), .Y(u0_u3__abc_44466_n538) );
  INVX1 INVX1_265 ( .A(u0_u3__abc_44466_n539), .Y(u0_u3__abc_44466_n540) );
  INVX1 INVX1_266 ( .A(u0_u3__abc_44466_n533), .Y(u0_u3__abc_44466_n541) );
  INVX1 INVX1_267 ( .A(u0_u3__abc_44466_n546), .Y(u0_u3__abc_44466_n547) );
  INVX1 INVX1_268 ( .A(u0_u3__abc_44466_n548), .Y(u0_u3__abc_44466_n549) );
  INVX1 INVX1_269 ( .A(u0_u3__abc_44466_n550), .Y(u0_u3__abc_44466_n553) );
  INVX1 INVX1_27 ( .A(u0__abc_49347_n4526_bF_buf3), .Y(u0__abc_49347_n4556) );
  INVX1 INVX1_270 ( .A(u0_u3__abc_44466_n557), .Y(u0_u3__abc_44466_n558) );
  INVX1 INVX1_271 ( .A(u0_u3__abc_44466_n561), .Y(u0_u3__abc_44466_n562) );
  INVX1 INVX1_272 ( .A(u0_u3__abc_44466_n566), .Y(u0_u3__abc_44466_n567) );
  INVX1 INVX1_273 ( .A(u0_u3__abc_44466_n560), .Y(u0_u3__abc_44466_n569) );
  INVX1 INVX1_274 ( .A(u0_u3__abc_44466_n565), .Y(u0_u3__abc_44466_n573) );
  INVX1 INVX1_275 ( .A(u0_u3__abc_44466_n511), .Y(u0_u3__abc_44466_n579) );
  INVX1 INVX1_276 ( .A(u0_u4_addr_r_6_), .Y(u0_u4__abc_44844_n201_1) );
  INVX1 INVX1_277 ( .A(u0_u4_addr_r_3_), .Y(u0_u4__abc_44844_n202) );
  INVX1 INVX1_278 ( .A(\wb_data_i[0] ), .Y(u0_u4__abc_44844_n210_1) );
  INVX1 INVX1_279 ( .A(u0_u4__abc_44844_n211), .Y(u0_u4__abc_44844_n212_1) );
  INVX1 INVX1_28 ( .A(u0__abc_49347_n4560_bF_buf4), .Y(u0__abc_49347_n4561) );
  INVX1 INVX1_280 ( .A(\wb_data_i[1] ), .Y(u0_u4__abc_44844_n216_1) );
  INVX1 INVX1_281 ( .A(u0_u4__abc_44844_n217), .Y(u0_u4__abc_44844_n218_1) );
  INVX1 INVX1_282 ( .A(\wb_data_i[2] ), .Y(u0_u4__abc_44844_n222_1) );
  INVX1 INVX1_283 ( .A(u0_u4__abc_44844_n223), .Y(u0_u4__abc_44844_n224_1) );
  INVX1 INVX1_284 ( .A(\wb_data_i[3] ), .Y(u0_u4__abc_44844_n228_1) );
  INVX1 INVX1_285 ( .A(u0_u4__abc_44844_n229), .Y(u0_u4__abc_44844_n230_1) );
  INVX1 INVX1_286 ( .A(\wb_data_i[4] ), .Y(u0_u4__abc_44844_n234_1) );
  INVX1 INVX1_287 ( .A(u0_u4__abc_44844_n235), .Y(u0_u4__abc_44844_n236_1) );
  INVX1 INVX1_288 ( .A(\wb_data_i[5] ), .Y(u0_u4__abc_44844_n240_1) );
  INVX1 INVX1_289 ( .A(u0_u4__abc_44844_n241), .Y(u0_u4__abc_44844_n242_1) );
  INVX1 INVX1_29 ( .A(u0__abc_49347_n4562_bF_buf4), .Y(u0__abc_49347_n4563) );
  INVX1 INVX1_290 ( .A(\wb_data_i[6] ), .Y(u0_u4__abc_44844_n246_1) );
  INVX1 INVX1_291 ( .A(u0_u4__abc_44844_n247), .Y(u0_u4__abc_44844_n248_1) );
  INVX1 INVX1_292 ( .A(\wb_data_i[7] ), .Y(u0_u4__abc_44844_n252_1) );
  INVX1 INVX1_293 ( .A(u0_u4__abc_44844_n253), .Y(u0_u4__abc_44844_n254) );
  INVX1 INVX1_294 ( .A(\wb_data_i[8] ), .Y(u0_u4__abc_44844_n258_1) );
  INVX1 INVX1_295 ( .A(u0_u4__abc_44844_n259_1), .Y(u0_u4__abc_44844_n260_1) );
  INVX1 INVX1_296 ( .A(\wb_data_i[9] ), .Y(u0_u4__abc_44844_n264) );
  INVX1 INVX1_297 ( .A(u0_u4__abc_44844_n265), .Y(u0_u4__abc_44844_n266) );
  INVX1 INVX1_298 ( .A(\wb_data_i[10] ), .Y(u0_u4__abc_44844_n270_1) );
  INVX1 INVX1_299 ( .A(u0_u4__abc_44844_n271), .Y(u0_u4__abc_44844_n272) );
  INVX1 INVX1_3 ( .A(u0__abc_49347_n1103_1), .Y(u0__abc_49347_n1104) );
  INVX1 INVX1_30 ( .A(u0__abc_49347_n4565), .Y(u0__abc_49347_n4566) );
  INVX1 INVX1_300 ( .A(\wb_data_i[11] ), .Y(u0_u4__abc_44844_n276_1) );
  INVX1 INVX1_301 ( .A(u0_u4__abc_44844_n277), .Y(u0_u4__abc_44844_n278) );
  INVX1 INVX1_302 ( .A(\wb_data_i[12] ), .Y(u0_u4__abc_44844_n282) );
  INVX1 INVX1_303 ( .A(u0_u4__abc_44844_n283_1), .Y(u0_u4__abc_44844_n284) );
  INVX1 INVX1_304 ( .A(\wb_data_i[13] ), .Y(u0_u4__abc_44844_n288) );
  INVX1 INVX1_305 ( .A(u0_u4__abc_44844_n289), .Y(u0_u4__abc_44844_n290) );
  INVX1 INVX1_306 ( .A(\wb_data_i[14] ), .Y(u0_u4__abc_44844_n294) );
  INVX1 INVX1_307 ( .A(u0_u4__abc_44844_n295_1), .Y(u0_u4__abc_44844_n296) );
  INVX1 INVX1_308 ( .A(\wb_data_i[15] ), .Y(u0_u4__abc_44844_n300) );
  INVX1 INVX1_309 ( .A(u0_u4__abc_44844_n301), .Y(u0_u4__abc_44844_n302) );
  INVX1 INVX1_31 ( .A(u0__abc_49347_n4567_bF_buf4), .Y(u0__abc_49347_n4568) );
  INVX1 INVX1_310 ( .A(\wb_data_i[16] ), .Y(u0_u4__abc_44844_n306_1) );
  INVX1 INVX1_311 ( .A(u0_u4__abc_44844_n307), .Y(u0_u4__abc_44844_n308) );
  INVX1 INVX1_312 ( .A(\wb_data_i[17] ), .Y(u0_u4__abc_44844_n312) );
  INVX1 INVX1_313 ( .A(u0_u4__abc_44844_n313), .Y(u0_u4__abc_44844_n314) );
  INVX1 INVX1_314 ( .A(\wb_data_i[18] ), .Y(u0_u4__abc_44844_n318_1) );
  INVX1 INVX1_315 ( .A(u0_u4__abc_44844_n319), .Y(u0_u4__abc_44844_n320_1) );
  INVX1 INVX1_316 ( .A(\wb_data_i[19] ), .Y(u0_u4__abc_44844_n324_1) );
  INVX1 INVX1_317 ( .A(u0_u4__abc_44844_n325), .Y(u0_u4__abc_44844_n326) );
  INVX1 INVX1_318 ( .A(\wb_data_i[20] ), .Y(u0_u4__abc_44844_n330) );
  INVX1 INVX1_319 ( .A(u0_u4__abc_44844_n331), .Y(u0_u4__abc_44844_n332) );
  INVX1 INVX1_32 ( .A(u0__abc_49347_n4571_bF_buf4), .Y(u0__abc_49347_n4572) );
  INVX1 INVX1_320 ( .A(\wb_data_i[21] ), .Y(u0_u4__abc_44844_n336) );
  INVX1 INVX1_321 ( .A(u0_u4__abc_44844_n337), .Y(u0_u4__abc_44844_n338) );
  INVX1 INVX1_322 ( .A(\wb_data_i[22] ), .Y(u0_u4__abc_44844_n342) );
  INVX1 INVX1_323 ( .A(u0_u4__abc_44844_n343), .Y(u0_u4__abc_44844_n344) );
  INVX1 INVX1_324 ( .A(\wb_data_i[23] ), .Y(u0_u4__abc_44844_n348) );
  INVX1 INVX1_325 ( .A(u0_u4__abc_44844_n349), .Y(u0_u4__abc_44844_n350) );
  INVX1 INVX1_326 ( .A(\wb_data_i[24] ), .Y(u0_u4__abc_44844_n354) );
  INVX1 INVX1_327 ( .A(u0_u4__abc_44844_n355), .Y(u0_u4__abc_44844_n356) );
  INVX1 INVX1_328 ( .A(\wb_data_i[25] ), .Y(u0_u4__abc_44844_n360) );
  INVX1 INVX1_329 ( .A(u0_u4__abc_44844_n361), .Y(u0_u4__abc_44844_n362) );
  INVX1 INVX1_33 ( .A(u0__abc_49347_n4573), .Y(u0__abc_49347_n4574) );
  INVX1 INVX1_330 ( .A(\wb_data_i[26] ), .Y(u0_u4__abc_44844_n366) );
  INVX1 INVX1_331 ( .A(u0_u4__abc_44844_n367), .Y(u0_u4__abc_44844_n368) );
  INVX1 INVX1_332 ( .A(\wb_data_i[27] ), .Y(u0_u4__abc_44844_n372) );
  INVX1 INVX1_333 ( .A(u0_u4__abc_44844_n373), .Y(u0_u4__abc_44844_n374) );
  INVX1 INVX1_334 ( .A(\wb_data_i[28] ), .Y(u0_u4__abc_44844_n378) );
  INVX1 INVX1_335 ( .A(u0_u4__abc_44844_n379), .Y(u0_u4__abc_44844_n380) );
  INVX1 INVX1_336 ( .A(\wb_data_i[29] ), .Y(u0_u4__abc_44844_n384) );
  INVX1 INVX1_337 ( .A(u0_u4__abc_44844_n385), .Y(u0_u4__abc_44844_n386) );
  INVX1 INVX1_338 ( .A(\wb_data_i[30] ), .Y(u0_u4__abc_44844_n390) );
  INVX1 INVX1_339 ( .A(u0_u4__abc_44844_n391), .Y(u0_u4__abc_44844_n392) );
  INVX1 INVX1_34 ( .A(u0__abc_49347_n4531_bF_buf3), .Y(u0__abc_49347_n4577) );
  INVX1 INVX1_340 ( .A(\wb_data_i[31] ), .Y(u0_u4__abc_44844_n396) );
  INVX1 INVX1_341 ( .A(u0_u4__abc_44844_n397), .Y(u0_u4__abc_44844_n398) );
  INVX1 INVX1_342 ( .A(u0_u4__abc_44844_n402), .Y(u0_u4__abc_44844_n403) );
  INVX1 INVX1_343 ( .A(u0_u4__abc_44844_n404), .Y(u0_u4__abc_44844_n406) );
  INVX1 INVX1_344 ( .A(u0_lmr_ack4), .Y(u0_u4__abc_44844_n407) );
  INVX1 INVX1_345 ( .A(u0_u4_addr_r_2_), .Y(u0_u4__abc_44844_n411) );
  INVX1 INVX1_346 ( .A(u0_u4__abc_44844_n414), .Y(u0_u4__abc_44844_n415) );
  INVX1 INVX1_347 ( .A(u0_u4__abc_44844_n419), .Y(u0_u4__abc_44844_n420) );
  INVX1 INVX1_348 ( .A(u0_u4__abc_44844_n424), .Y(u0_u4__abc_44844_n425) );
  INVX1 INVX1_349 ( .A(u0_u4__abc_44844_n429), .Y(u0_u4__abc_44844_n430) );
  INVX1 INVX1_35 ( .A(u0__abc_49347_n4539_bF_buf3), .Y(u0__abc_49347_n4578) );
  INVX1 INVX1_350 ( .A(u0_u4__abc_44844_n434), .Y(u0_u4__abc_44844_n435) );
  INVX1 INVX1_351 ( .A(u0_u4__abc_44844_n439), .Y(u0_u4__abc_44844_n440) );
  INVX1 INVX1_352 ( .A(u0_u4__abc_44844_n444), .Y(u0_u4__abc_44844_n445) );
  INVX1 INVX1_353 ( .A(u0_u4__abc_44844_n449), .Y(u0_u4__abc_44844_n450) );
  INVX1 INVX1_354 ( .A(u0_u4__abc_44844_n454), .Y(u0_u4__abc_44844_n455) );
  INVX1 INVX1_355 ( .A(u0_u4__abc_44844_n459), .Y(u0_u4__abc_44844_n460) );
  INVX1 INVX1_356 ( .A(u0_u4__abc_44844_n464), .Y(u0_u4__abc_44844_n465) );
  INVX1 INVX1_357 ( .A(u0_u4__abc_44844_n469), .Y(u0_u4__abc_44844_n470) );
  INVX1 INVX1_358 ( .A(u0_u4__abc_44844_n474), .Y(u0_u4__abc_44844_n475) );
  INVX1 INVX1_359 ( .A(u0_u4__abc_44844_n479), .Y(u0_u4__abc_44844_n480) );
  INVX1 INVX1_36 ( .A(\wb_addr_i[31] ), .Y(u0__abc_49347_n5683) );
  INVX1 INVX1_360 ( .A(u0_u4__abc_44844_n484), .Y(u0_u4__abc_44844_n485) );
  INVX1 INVX1_361 ( .A(u0_u4__abc_44844_n489), .Y(u0_u4__abc_44844_n490) );
  INVX1 INVX1_362 ( .A(u0_u4__abc_44844_n494), .Y(u0_u4__abc_44844_n495) );
  INVX1 INVX1_363 ( .A(u0_u4__abc_44844_n499), .Y(u0_u4__abc_44844_n500) );
  INVX1 INVX1_364 ( .A(u0_u4__abc_44844_n504), .Y(u0_u4__abc_44844_n505) );
  INVX1 INVX1_365 ( .A(u0_u4__abc_44844_n509), .Y(u0_u4__abc_44844_n510) );
  INVX1 INVX1_366 ( .A(u0_u4__abc_44844_n514), .Y(u0_u4__abc_44844_n515) );
  INVX1 INVX1_367 ( .A(u0_u4__abc_44844_n519), .Y(u0_u4__abc_44844_n520) );
  INVX1 INVX1_368 ( .A(u0_u4__abc_44844_n524), .Y(u0_u4__abc_44844_n525) );
  INVX1 INVX1_369 ( .A(u0_u4__abc_44844_n529), .Y(u0_u4__abc_44844_n530) );
  INVX1 INVX1_37 ( .A(u0_csc0_1_), .Y(u0__abc_49347_n5692) );
  INVX1 INVX1_370 ( .A(u0_u4__abc_44844_n534), .Y(u0_u4__abc_44844_n535) );
  INVX1 INVX1_371 ( .A(u0_u4__abc_44844_n539), .Y(u0_u4__abc_44844_n540) );
  INVX1 INVX1_372 ( .A(u0_u4__abc_44844_n544), .Y(u0_u4__abc_44844_n545) );
  INVX1 INVX1_373 ( .A(u0_u4__abc_44844_n549), .Y(u0_u4__abc_44844_n550) );
  INVX1 INVX1_374 ( .A(u0_u4__abc_44844_n554), .Y(u0_u4__abc_44844_n555) );
  INVX1 INVX1_375 ( .A(u0_u4__abc_44844_n559), .Y(u0_u4__abc_44844_n560) );
  INVX1 INVX1_376 ( .A(u0_u4__abc_44844_n564), .Y(u0_u4__abc_44844_n565) );
  INVX1 INVX1_377 ( .A(u0_u4__abc_44844_n569), .Y(u0_u4__abc_44844_n570) );
  INVX1 INVX1_378 ( .A(u0_init_ack4), .Y(u0_u4__abc_44844_n573) );
  INVX1 INVX1_379 ( .A(u0_u4_inited), .Y(u0_u4__abc_44844_n575) );
  INVX1 INVX1_38 ( .A(u0_csc0_2_), .Y(u0__abc_49347_n5694) );
  INVX1 INVX1_380 ( .A(u0_u4__abc_44844_n583), .Y(u0_u4__abc_44844_n584) );
  INVX1 INVX1_381 ( .A(u0_u4__abc_44844_n587), .Y(u0_u4__abc_44844_n588) );
  INVX1 INVX1_382 ( .A(wb_addr_i_23_bF_buf3), .Y(u0_u4__abc_44844_n591) );
  INVX1 INVX1_383 ( .A(u0_u4__abc_44844_n593), .Y(u0_u4__abc_44844_n594) );
  INVX1 INVX1_384 ( .A(u0_u4__abc_44844_n586), .Y(u0_u4__abc_44844_n595) );
  INVX1 INVX1_385 ( .A(u0_u4__abc_44844_n600), .Y(u0_u4__abc_44844_n601) );
  INVX1 INVX1_386 ( .A(u0_u4__abc_44844_n604), .Y(u0_u4__abc_44844_n605) );
  INVX1 INVX1_387 ( .A(wb_addr_i_25_bF_buf2), .Y(u0_u4__abc_44844_n608) );
  INVX1 INVX1_388 ( .A(u0_u4__abc_44844_n609), .Y(u0_u4__abc_44844_n610) );
  INVX1 INVX1_389 ( .A(u0_u4__abc_44844_n603), .Y(u0_u4__abc_44844_n611) );
  INVX1 INVX1_39 ( .A(u0_csc0_3_), .Y(u0__abc_49347_n5695) );
  INVX1 INVX1_390 ( .A(u0_u4__abc_44844_n616), .Y(u0_u4__abc_44844_n617) );
  INVX1 INVX1_391 ( .A(u0_u4__abc_44844_n618), .Y(u0_u4__abc_44844_n619) );
  INVX1 INVX1_392 ( .A(u0_u4__abc_44844_n620), .Y(u0_u4__abc_44844_n623) );
  INVX1 INVX1_393 ( .A(u0_u4__abc_44844_n627), .Y(u0_u4__abc_44844_n628) );
  INVX1 INVX1_394 ( .A(u0_u4__abc_44844_n631), .Y(u0_u4__abc_44844_n632) );
  INVX1 INVX1_395 ( .A(u0_u4__abc_44844_n636), .Y(u0_u4__abc_44844_n637) );
  INVX1 INVX1_396 ( .A(u0_u4__abc_44844_n630), .Y(u0_u4__abc_44844_n639) );
  INVX1 INVX1_397 ( .A(u0_u4__abc_44844_n635), .Y(u0_u4__abc_44844_n643) );
  INVX1 INVX1_398 ( .A(u0_u4__abc_44844_n581), .Y(u0_u4__abc_44844_n649) );
  INVX1 INVX1_399 ( .A(u0_u5__abc_45296_n202_1), .Y(u0_u5__abc_45296_n203) );
  INVX1 INVX1_4 ( .A(u0__abc_49347_n1105_1), .Y(u0__abc_49347_n1106) );
  INVX1 INVX1_40 ( .A(u0_csc1_1_), .Y(u0__abc_49347_n5698) );
  INVX1 INVX1_400 ( .A(u0_u5__abc_45296_n204_1), .Y(u0_u5__abc_45296_n206) );
  INVX1 INVX1_401 ( .A(u0_lmr_ack5), .Y(u0_u5__abc_45296_n207_1) );
  INVX1 INVX1_402 ( .A(u0_u5_addr_r_6_), .Y(u0_u5__abc_45296_n211_1) );
  INVX1 INVX1_403 ( .A(\wb_data_i[0] ), .Y(u0_u5__abc_45296_n219_1) );
  INVX1 INVX1_404 ( .A(u0_u5__abc_45296_n220_1), .Y(u0_u5__abc_45296_n221) );
  INVX1 INVX1_405 ( .A(\wb_data_i[1] ), .Y(u0_u5__abc_45296_n225_1) );
  INVX1 INVX1_406 ( .A(u0_u5__abc_45296_n226_1), .Y(u0_u5__abc_45296_n227) );
  INVX1 INVX1_407 ( .A(\wb_data_i[2] ), .Y(u0_u5__abc_45296_n231_1) );
  INVX1 INVX1_408 ( .A(u0_u5__abc_45296_n232_1), .Y(u0_u5__abc_45296_n233) );
  INVX1 INVX1_409 ( .A(\wb_data_i[3] ), .Y(u0_u5__abc_45296_n237_1) );
  INVX1 INVX1_41 ( .A(u0_csc1_2_), .Y(u0__abc_49347_n5700) );
  INVX1 INVX1_410 ( .A(u0_u5__abc_45296_n238_1), .Y(u0_u5__abc_45296_n239) );
  INVX1 INVX1_411 ( .A(\wb_data_i[4] ), .Y(u0_u5__abc_45296_n243_1) );
  INVX1 INVX1_412 ( .A(u0_u5__abc_45296_n244_1), .Y(u0_u5__abc_45296_n245) );
  INVX1 INVX1_413 ( .A(\wb_data_i[5] ), .Y(u0_u5__abc_45296_n249_1) );
  INVX1 INVX1_414 ( .A(u0_u5__abc_45296_n250_1), .Y(u0_u5__abc_45296_n251) );
  INVX1 INVX1_415 ( .A(\wb_data_i[6] ), .Y(u0_u5__abc_45296_n255_1) );
  INVX1 INVX1_416 ( .A(u0_u5__abc_45296_n256), .Y(u0_u5__abc_45296_n257) );
  INVX1 INVX1_417 ( .A(\wb_data_i[7] ), .Y(u0_u5__abc_45296_n261) );
  INVX1 INVX1_418 ( .A(u0_u5__abc_45296_n262_1), .Y(u0_u5__abc_45296_n263) );
  INVX1 INVX1_419 ( .A(\wb_data_i[8] ), .Y(u0_u5__abc_45296_n267) );
  INVX1 INVX1_42 ( .A(u0_csc1_3_), .Y(u0__abc_49347_n5701) );
  INVX1 INVX1_420 ( .A(u0_u5__abc_45296_n268_1), .Y(u0_u5__abc_45296_n269) );
  INVX1 INVX1_421 ( .A(\wb_data_i[9] ), .Y(u0_u5__abc_45296_n273_1) );
  INVX1 INVX1_422 ( .A(u0_u5__abc_45296_n274), .Y(u0_u5__abc_45296_n275_1) );
  INVX1 INVX1_423 ( .A(\wb_data_i[10] ), .Y(u0_u5__abc_45296_n279_1) );
  INVX1 INVX1_424 ( .A(u0_u5__abc_45296_n280), .Y(u0_u5__abc_45296_n281) );
  INVX1 INVX1_425 ( .A(\wb_data_i[11] ), .Y(u0_u5__abc_45296_n285_1) );
  INVX1 INVX1_426 ( .A(u0_u5__abc_45296_n286), .Y(u0_u5__abc_45296_n287_1) );
  INVX1 INVX1_427 ( .A(\wb_data_i[12] ), .Y(u0_u5__abc_45296_n291) );
  INVX1 INVX1_428 ( .A(u0_u5__abc_45296_n292), .Y(u0_u5__abc_45296_n293) );
  INVX1 INVX1_429 ( .A(\wb_data_i[13] ), .Y(u0_u5__abc_45296_n297) );
  INVX1 INVX1_43 ( .A(u0_csc2_1_), .Y(u0__abc_49347_n5704) );
  INVX1 INVX1_430 ( .A(u0_u5__abc_45296_n298_1), .Y(u0_u5__abc_45296_n299) );
  INVX1 INVX1_431 ( .A(\wb_data_i[14] ), .Y(u0_u5__abc_45296_n303) );
  INVX1 INVX1_432 ( .A(u0_u5__abc_45296_n304), .Y(u0_u5__abc_45296_n305) );
  INVX1 INVX1_433 ( .A(\wb_data_i[15] ), .Y(u0_u5__abc_45296_n309) );
  INVX1 INVX1_434 ( .A(u0_u5__abc_45296_n310_1), .Y(u0_u5__abc_45296_n311) );
  INVX1 INVX1_435 ( .A(\wb_data_i[16] ), .Y(u0_u5__abc_45296_n315_1) );
  INVX1 INVX1_436 ( .A(u0_u5__abc_45296_n316_1), .Y(u0_u5__abc_45296_n317_1) );
  INVX1 INVX1_437 ( .A(\wb_data_i[17] ), .Y(u0_u5__abc_45296_n321_1) );
  INVX1 INVX1_438 ( .A(u0_u5__abc_45296_n322), .Y(u0_u5__abc_45296_n323_1) );
  INVX1 INVX1_439 ( .A(\wb_data_i[18] ), .Y(u0_u5__abc_45296_n327) );
  INVX1 INVX1_44 ( .A(u0_csc2_2_), .Y(u0__abc_49347_n5706) );
  INVX1 INVX1_440 ( .A(u0_u5__abc_45296_n328), .Y(u0_u5__abc_45296_n329) );
  INVX1 INVX1_441 ( .A(\wb_data_i[19] ), .Y(u0_u5__abc_45296_n333) );
  INVX1 INVX1_442 ( .A(u0_u5__abc_45296_n334), .Y(u0_u5__abc_45296_n335) );
  INVX1 INVX1_443 ( .A(\wb_data_i[20] ), .Y(u0_u5__abc_45296_n339) );
  INVX1 INVX1_444 ( .A(u0_u5__abc_45296_n340), .Y(u0_u5__abc_45296_n341) );
  INVX1 INVX1_445 ( .A(\wb_data_i[21] ), .Y(u0_u5__abc_45296_n345) );
  INVX1 INVX1_446 ( .A(u0_u5__abc_45296_n346), .Y(u0_u5__abc_45296_n347) );
  INVX1 INVX1_447 ( .A(\wb_data_i[22] ), .Y(u0_u5__abc_45296_n351) );
  INVX1 INVX1_448 ( .A(u0_u5__abc_45296_n352), .Y(u0_u5__abc_45296_n353) );
  INVX1 INVX1_449 ( .A(\wb_data_i[23] ), .Y(u0_u5__abc_45296_n357) );
  INVX1 INVX1_45 ( .A(u0_csc2_3_), .Y(u0__abc_49347_n5707) );
  INVX1 INVX1_450 ( .A(u0_u5__abc_45296_n358), .Y(u0_u5__abc_45296_n359) );
  INVX1 INVX1_451 ( .A(\wb_data_i[24] ), .Y(u0_u5__abc_45296_n363) );
  INVX1 INVX1_452 ( .A(u0_u5__abc_45296_n364), .Y(u0_u5__abc_45296_n365) );
  INVX1 INVX1_453 ( .A(\wb_data_i[25] ), .Y(u0_u5__abc_45296_n369) );
  INVX1 INVX1_454 ( .A(u0_u5__abc_45296_n370), .Y(u0_u5__abc_45296_n371) );
  INVX1 INVX1_455 ( .A(\wb_data_i[26] ), .Y(u0_u5__abc_45296_n375) );
  INVX1 INVX1_456 ( .A(u0_u5__abc_45296_n376), .Y(u0_u5__abc_45296_n377) );
  INVX1 INVX1_457 ( .A(\wb_data_i[27] ), .Y(u0_u5__abc_45296_n381) );
  INVX1 INVX1_458 ( .A(u0_u5__abc_45296_n382), .Y(u0_u5__abc_45296_n383) );
  INVX1 INVX1_459 ( .A(\wb_data_i[28] ), .Y(u0_u5__abc_45296_n387) );
  INVX1 INVX1_46 ( .A(u0_csc3_1_), .Y(u0__abc_49347_n5710) );
  INVX1 INVX1_460 ( .A(u0_u5__abc_45296_n388), .Y(u0_u5__abc_45296_n389) );
  INVX1 INVX1_461 ( .A(\wb_data_i[29] ), .Y(u0_u5__abc_45296_n393) );
  INVX1 INVX1_462 ( .A(u0_u5__abc_45296_n394), .Y(u0_u5__abc_45296_n395) );
  INVX1 INVX1_463 ( .A(\wb_data_i[30] ), .Y(u0_u5__abc_45296_n399) );
  INVX1 INVX1_464 ( .A(u0_u5__abc_45296_n400), .Y(u0_u5__abc_45296_n401) );
  INVX1 INVX1_465 ( .A(\wb_data_i[31] ), .Y(u0_u5__abc_45296_n405) );
  INVX1 INVX1_466 ( .A(u0_u5__abc_45296_n406), .Y(u0_u5__abc_45296_n407) );
  INVX1 INVX1_467 ( .A(u0_u5_addr_r_2_), .Y(u0_u5__abc_45296_n410) );
  INVX1 INVX1_468 ( .A(u0_u5__abc_45296_n413), .Y(u0_u5__abc_45296_n414) );
  INVX1 INVX1_469 ( .A(u0_u5__abc_45296_n418), .Y(u0_u5__abc_45296_n419) );
  INVX1 INVX1_47 ( .A(u0_csc3_2_), .Y(u0__abc_49347_n5712) );
  INVX1 INVX1_470 ( .A(u0_u5__abc_45296_n423), .Y(u0_u5__abc_45296_n424) );
  INVX1 INVX1_471 ( .A(u0_u5__abc_45296_n428), .Y(u0_u5__abc_45296_n429) );
  INVX1 INVX1_472 ( .A(u0_u5__abc_45296_n433), .Y(u0_u5__abc_45296_n434) );
  INVX1 INVX1_473 ( .A(u0_u5__abc_45296_n438), .Y(u0_u5__abc_45296_n439) );
  INVX1 INVX1_474 ( .A(u0_u5__abc_45296_n443), .Y(u0_u5__abc_45296_n444) );
  INVX1 INVX1_475 ( .A(u0_u5__abc_45296_n448), .Y(u0_u5__abc_45296_n449) );
  INVX1 INVX1_476 ( .A(u0_u5__abc_45296_n453), .Y(u0_u5__abc_45296_n454) );
  INVX1 INVX1_477 ( .A(u0_u5__abc_45296_n458), .Y(u0_u5__abc_45296_n459) );
  INVX1 INVX1_478 ( .A(u0_u5__abc_45296_n463), .Y(u0_u5__abc_45296_n464) );
  INVX1 INVX1_479 ( .A(u0_u5__abc_45296_n468), .Y(u0_u5__abc_45296_n469) );
  INVX1 INVX1_48 ( .A(u0_csc3_3_), .Y(u0__abc_49347_n5713) );
  INVX1 INVX1_480 ( .A(u0_u5__abc_45296_n473), .Y(u0_u5__abc_45296_n474) );
  INVX1 INVX1_481 ( .A(u0_u5__abc_45296_n478), .Y(u0_u5__abc_45296_n479) );
  INVX1 INVX1_482 ( .A(u0_u5__abc_45296_n483), .Y(u0_u5__abc_45296_n484) );
  INVX1 INVX1_483 ( .A(u0_u5__abc_45296_n488), .Y(u0_u5__abc_45296_n489) );
  INVX1 INVX1_484 ( .A(u0_u5__abc_45296_n493), .Y(u0_u5__abc_45296_n494) );
  INVX1 INVX1_485 ( .A(u0_u5__abc_45296_n498), .Y(u0_u5__abc_45296_n499) );
  INVX1 INVX1_486 ( .A(u0_u5__abc_45296_n503), .Y(u0_u5__abc_45296_n504) );
  INVX1 INVX1_487 ( .A(u0_u5__abc_45296_n508), .Y(u0_u5__abc_45296_n509) );
  INVX1 INVX1_488 ( .A(u0_u5__abc_45296_n513), .Y(u0_u5__abc_45296_n514) );
  INVX1 INVX1_489 ( .A(u0_u5__abc_45296_n518), .Y(u0_u5__abc_45296_n519) );
  INVX1 INVX1_49 ( .A(u0_csc4_1_), .Y(u0__abc_49347_n5716) );
  INVX1 INVX1_490 ( .A(u0_u5__abc_45296_n523), .Y(u0_u5__abc_45296_n524) );
  INVX1 INVX1_491 ( .A(u0_u5__abc_45296_n528), .Y(u0_u5__abc_45296_n529) );
  INVX1 INVX1_492 ( .A(u0_u5__abc_45296_n533), .Y(u0_u5__abc_45296_n534) );
  INVX1 INVX1_493 ( .A(u0_u5__abc_45296_n538), .Y(u0_u5__abc_45296_n539) );
  INVX1 INVX1_494 ( .A(u0_u5__abc_45296_n543), .Y(u0_u5__abc_45296_n544) );
  INVX1 INVX1_495 ( .A(u0_u5__abc_45296_n548), .Y(u0_u5__abc_45296_n549) );
  INVX1 INVX1_496 ( .A(u0_u5__abc_45296_n553), .Y(u0_u5__abc_45296_n554) );
  INVX1 INVX1_497 ( .A(u0_u5__abc_45296_n558), .Y(u0_u5__abc_45296_n559) );
  INVX1 INVX1_498 ( .A(u0_u5__abc_45296_n563), .Y(u0_u5__abc_45296_n564) );
  INVX1 INVX1_499 ( .A(u0_u5__abc_45296_n568), .Y(u0_u5__abc_45296_n569) );
  INVX1 INVX1_5 ( .A(u0__abc_49347_n1111_1), .Y(u0__abc_49347_n1117_1) );
  INVX1 INVX1_50 ( .A(u0_csc4_2_), .Y(u0__abc_49347_n5718) );
  INVX1 INVX1_500 ( .A(u0_u5__abc_45296_n574), .Y(u0_u5__abc_45296_n575) );
  INVX1 INVX1_501 ( .A(u0_u5__abc_45296_n578), .Y(u0_u5__abc_45296_n579) );
  INVX1 INVX1_502 ( .A(wb_addr_i_23_bF_buf1), .Y(u0_u5__abc_45296_n582) );
  INVX1 INVX1_503 ( .A(u0_u5__abc_45296_n584), .Y(u0_u5__abc_45296_n585) );
  INVX1 INVX1_504 ( .A(u0_u5__abc_45296_n577), .Y(u0_u5__abc_45296_n586) );
  INVX1 INVX1_505 ( .A(u0_u5__abc_45296_n591), .Y(u0_u5__abc_45296_n592) );
  INVX1 INVX1_506 ( .A(u0_u5__abc_45296_n595), .Y(u0_u5__abc_45296_n596) );
  INVX1 INVX1_507 ( .A(wb_addr_i_25_bF_buf0), .Y(u0_u5__abc_45296_n599) );
  INVX1 INVX1_508 ( .A(u0_u5__abc_45296_n600), .Y(u0_u5__abc_45296_n601) );
  INVX1 INVX1_509 ( .A(u0_u5__abc_45296_n594), .Y(u0_u5__abc_45296_n602) );
  INVX1 INVX1_51 ( .A(u0_csc4_3_), .Y(u0__abc_49347_n5719) );
  INVX1 INVX1_510 ( .A(u0_u5__abc_45296_n607), .Y(u0_u5__abc_45296_n608) );
  INVX1 INVX1_511 ( .A(u0_u5__abc_45296_n609), .Y(u0_u5__abc_45296_n610) );
  INVX1 INVX1_512 ( .A(u0_u5__abc_45296_n611), .Y(u0_u5__abc_45296_n614) );
  INVX1 INVX1_513 ( .A(u0_u5__abc_45296_n618), .Y(u0_u5__abc_45296_n619) );
  INVX1 INVX1_514 ( .A(u0_u5__abc_45296_n622), .Y(u0_u5__abc_45296_n623) );
  INVX1 INVX1_515 ( .A(u0_u5__abc_45296_n627), .Y(u0_u5__abc_45296_n628) );
  INVX1 INVX1_516 ( .A(u0_u5__abc_45296_n621), .Y(u0_u5__abc_45296_n630) );
  INVX1 INVX1_517 ( .A(u0_u5__abc_45296_n626), .Y(u0_u5__abc_45296_n634) );
  INVX1 INVX1_518 ( .A(u0_u5__abc_45296_n572), .Y(u0_u5__abc_45296_n640) );
  INVX1 INVX1_519 ( .A(u0_init_ack5), .Y(u0_u5__abc_45296_n643) );
  INVX1 INVX1_52 ( .A(u0_csc5_1_), .Y(u0__abc_49347_n5722) );
  INVX1 INVX1_520 ( .A(u0_u5_inited), .Y(u0_u5__abc_45296_n645) );
  INVX1 INVX1_521 ( .A(csc_s_7_), .Y(u1__abc_45852_n258_1) );
  INVX1 INVX1_522 ( .A(csc_s_6_), .Y(u1__abc_45852_n263) );
  INVX1 INVX1_523 ( .A(page_size_10_bF_buf3), .Y(u1__abc_45852_n267_1) );
  INVX1 INVX1_524 ( .A(csc_s_4_), .Y(u1__abc_45852_n269) );
  INVX1 INVX1_525 ( .A(csc_s_5_bF_buf2), .Y(u1__abc_45852_n275) );
  INVX1 INVX1_526 ( .A(u1__abc_45852_n277), .Y(u1__abc_45852_n278_1) );
  INVX1 INVX1_527 ( .A(u1__abc_45852_n272_1), .Y(u1__abc_45852_n291) );
  INVX1 INVX1_528 ( .A(u1__abc_45852_n297), .Y(u1__abc_45852_n298) );
  INVX1 INVX1_529 ( .A(u1__abc_45852_n273_1), .Y(u1__abc_45852_n362) );
  INVX1 INVX1_53 ( .A(u0_csc5_2_), .Y(u0__abc_49347_n5724) );
  INVX1 INVX1_530 ( .A(u1_wr_cycle), .Y(u1__abc_45852_n516) );
  INVX1 INVX1_531 ( .A(page_size_8_), .Y(u1__abc_45852_n546) );
  INVX1 INVX1_532 ( .A(u1__abc_45852_n893_bF_buf3), .Y(u1__abc_45852_n896) );
  INVX1 INVX1_533 ( .A(u1__abc_45852_n898), .Y(u1__abc_45852_n899) );
  INVX1 INVX1_534 ( .A(cas_), .Y(u1__abc_45852_n908) );
  INVX1 INVX1_535 ( .A(csc_s_2_bF_buf1), .Y(u1__abc_45852_n915) );
  INVX1 INVX1_536 ( .A(u1_u0__abc_45749_n52_1), .Y(u1_u0__abc_45749_n53_1) );
  INVX1 INVX1_537 ( .A(u1_u0__abc_45749_n56_1), .Y(u1_u0__abc_45749_n57) );
  INVX1 INVX1_538 ( .A(u1_u0__abc_45749_n62_1), .Y(u1_u0__abc_45749_n63_1) );
  INVX1 INVX1_539 ( .A(u1_u0__abc_45749_n65), .Y(u1_u0__abc_45749_n66) );
  INVX1 INVX1_54 ( .A(u0_csc5_3_), .Y(u0__abc_49347_n5725) );
  INVX1 INVX1_540 ( .A(u1_u0__abc_45749_n71_1), .Y(u1_u0__abc_45749_n72) );
  INVX1 INVX1_541 ( .A(u1_u0__abc_45749_n74_1), .Y(u1_u0__abc_45749_n75_1) );
  INVX1 INVX1_542 ( .A(u1_u0__abc_45749_n81), .Y(u1_u0__abc_45749_n82_1) );
  INVX1 INVX1_543 ( .A(u1_u0__abc_45749_n84), .Y(u1_u0__abc_45749_n85) );
  INVX1 INVX1_544 ( .A(u1_u0__abc_45749_n90), .Y(u1_u0__abc_45749_n91) );
  INVX1 INVX1_545 ( .A(u1_u0__abc_45749_n93), .Y(u1_u0__abc_45749_n94) );
  INVX1 INVX1_546 ( .A(u1_u0__abc_45749_n98), .Y(u1_u0__abc_45749_n99) );
  INVX1 INVX1_547 ( .A(u1_u0__abc_45749_n51), .Y(u1_u0__abc_45749_n101) );
  INVX1 INVX1_548 ( .A(u1_u0__abc_45749_n104), .Y(u1_u0__abc_45749_n105) );
  INVX1 INVX1_549 ( .A(u1_u0__abc_45749_n108), .Y(u1_u0__abc_45749_n109) );
  INVX1 INVX1_55 ( .A(1'b0), .Y(u0__abc_49347_n5728) );
  INVX1 INVX1_550 ( .A(u1_u0__abc_45749_n112), .Y(u1_u0__abc_45749_n113) );
  INVX1 INVX1_551 ( .A(u1_u0__abc_45749_n116), .Y(u1_u0__abc_45749_n117) );
  INVX1 INVX1_552 ( .A(u1_u0__abc_45749_n122), .Y(u1_u0__abc_45749_n123) );
  INVX1 INVX1_553 ( .A(u1_u0__abc_45749_n125), .Y(u1_u0__abc_45749_n126) );
  INVX1 INVX1_554 ( .A(u1_u0__abc_45749_n132), .Y(u1_u0__abc_45749_n133) );
  INVX1 INVX1_555 ( .A(u1_u0__abc_45749_n135), .Y(u1_u0__abc_45749_n136) );
  INVX1 INVX1_556 ( .A(u1_u0__abc_45749_n141), .Y(u1_u0__abc_45749_n142) );
  INVX1 INVX1_557 ( .A(u1_u0__abc_45749_n144), .Y(u1_u0__abc_45749_n145) );
  INVX1 INVX1_558 ( .A(u1_u0_out_r_12__FF_INPUT), .Y(u1_u0__abc_45749_n149) );
  INVX1 INVX1_559 ( .A(u1_acs_addr_0_), .Y(u1_u0_out_r_0__FF_INPUT) );
  INVX1 INVX1_56 ( .A(1'b0), .Y(u0__abc_49347_n5730) );
  INVX1 INVX1_560 ( .A(u2_u0__abc_47660_n140), .Y(u2_u0__abc_47660_n141) );
  INVX1 INVX1_561 ( .A(u2_u0__abc_47660_n145), .Y(u2_u0__abc_47660_n146) );
  INVX1 INVX1_562 ( .A(u2_u0__abc_47660_n150), .Y(u2_u0__abc_47660_n151) );
  INVX1 INVX1_563 ( .A(u2_u0__abc_47660_n155), .Y(u2_u0__abc_47660_n156) );
  INVX1 INVX1_564 ( .A(u2_u0__abc_47660_n160), .Y(u2_u0__abc_47660_n161) );
  INVX1 INVX1_565 ( .A(u2_u0__abc_47660_n165), .Y(u2_u0__abc_47660_n166) );
  INVX1 INVX1_566 ( .A(u2_u0__abc_47660_n170), .Y(u2_u0__abc_47660_n171) );
  INVX1 INVX1_567 ( .A(u2_u0__abc_47660_n175), .Y(u2_u0__abc_47660_n176) );
  INVX1 INVX1_568 ( .A(u2_u0__abc_47660_n180), .Y(u2_u0__abc_47660_n181) );
  INVX1 INVX1_569 ( .A(u2_u0__abc_47660_n185), .Y(u2_u0__abc_47660_n186) );
  INVX1 INVX1_57 ( .A(1'b0), .Y(u0__abc_49347_n5731) );
  INVX1 INVX1_570 ( .A(u2_u0__abc_47660_n190), .Y(u2_u0__abc_47660_n191) );
  INVX1 INVX1_571 ( .A(u2_u0__abc_47660_n195), .Y(u2_u0__abc_47660_n196) );
  INVX1 INVX1_572 ( .A(u2_u0__abc_47660_n200), .Y(u2_u0__abc_47660_n201) );
  INVX1 INVX1_573 ( .A(bank_adr_0_bF_buf0), .Y(u2_u0__abc_47660_n203) );
  INVX1 INVX1_574 ( .A(bank_adr_1_bF_buf3), .Y(u2_u0__abc_47660_n246) );
  INVX1 INVX1_575 ( .A(u2_u0_b0_last_row_12_), .Y(u2_u0__abc_47660_n331) );
  INVX1 INVX1_576 ( .A(u2_u0_b0_last_row_11_), .Y(u2_u0__abc_47660_n333) );
  INVX1 INVX1_577 ( .A(u2_u0_b0_last_row_9_), .Y(u2_u0__abc_47660_n339) );
  INVX1 INVX1_578 ( .A(u2_u0_b0_last_row_7_), .Y(u2_u0__abc_47660_n343) );
  INVX1 INVX1_579 ( .A(u2_u0_b0_last_row_4_), .Y(u2_u0__abc_47660_n351) );
  INVX1 INVX1_58 ( .A(1'b0), .Y(u0__abc_49347_n5734) );
  INVX1 INVX1_580 ( .A(u2_u0_b0_last_row_0_), .Y(u2_u0__abc_47660_n355) );
  INVX1 INVX1_581 ( .A(u2_u0_b0_last_row_5_), .Y(u2_u0__abc_47660_n360) );
  INVX1 INVX1_582 ( .A(u2_u0_b0_last_row_10_), .Y(u2_u0__abc_47660_n366) );
  INVX1 INVX1_583 ( .A(u2_u0_b0_last_row_8_), .Y(u2_u0__abc_47660_n371) );
  INVX1 INVX1_584 ( .A(u2_u0_b0_last_row_2_), .Y(u2_u0__abc_47660_n376) );
  INVX1 INVX1_585 ( .A(u2_u0_b0_last_row_1_), .Y(u2_u0__abc_47660_n379) );
  INVX1 INVX1_586 ( .A(u2_u0_b0_last_row_3_), .Y(u2_u0__abc_47660_n384) );
  INVX1 INVX1_587 ( .A(u2_u0_b0_last_row_6_), .Y(u2_u0__abc_47660_n389) );
  INVX1 INVX1_588 ( .A(u2_u0_b2_last_row_12_), .Y(u2_u0__abc_47660_n396) );
  INVX1 INVX1_589 ( .A(u2_u0_b2_last_row_11_), .Y(u2_u0__abc_47660_n398) );
  INVX1 INVX1_59 ( .A(1'b0), .Y(u0__abc_49347_n5736) );
  INVX1 INVX1_590 ( .A(u2_u0_b2_last_row_9_), .Y(u2_u0__abc_47660_n404) );
  INVX1 INVX1_591 ( .A(u2_u0_b2_last_row_7_), .Y(u2_u0__abc_47660_n408) );
  INVX1 INVX1_592 ( .A(u2_u0_b2_last_row_4_), .Y(u2_u0__abc_47660_n416) );
  INVX1 INVX1_593 ( .A(u2_u0_b2_last_row_0_), .Y(u2_u0__abc_47660_n420) );
  INVX1 INVX1_594 ( .A(u2_u0_b2_last_row_5_), .Y(u2_u0__abc_47660_n425) );
  INVX1 INVX1_595 ( .A(u2_u0_b2_last_row_10_), .Y(u2_u0__abc_47660_n431) );
  INVX1 INVX1_596 ( .A(u2_u0_b2_last_row_8_), .Y(u2_u0__abc_47660_n436) );
  INVX1 INVX1_597 ( .A(u2_u0_b2_last_row_2_), .Y(u2_u0__abc_47660_n441) );
  INVX1 INVX1_598 ( .A(u2_u0_b2_last_row_1_), .Y(u2_u0__abc_47660_n444) );
  INVX1 INVX1_599 ( .A(u2_u0_b2_last_row_3_), .Y(u2_u0__abc_47660_n449) );
  INVX1 INVX1_6 ( .A(u0__abc_49347_n1120_1), .Y(u0__abc_49347_n1125) );
  INVX1 INVX1_60 ( .A(1'b0), .Y(u0__abc_49347_n5737) );
  INVX1 INVX1_600 ( .A(u2_u0_b2_last_row_6_), .Y(u2_u0__abc_47660_n454) );
  INVX1 INVX1_601 ( .A(u2_u0_b1_last_row_12_), .Y(u2_u0__abc_47660_n462) );
  INVX1 INVX1_602 ( .A(u2_u0_b1_last_row_11_), .Y(u2_u0__abc_47660_n464) );
  INVX1 INVX1_603 ( .A(u2_u0_b1_last_row_9_), .Y(u2_u0__abc_47660_n470) );
  INVX1 INVX1_604 ( .A(u2_u0_b1_last_row_7_), .Y(u2_u0__abc_47660_n474) );
  INVX1 INVX1_605 ( .A(u2_u0_b1_last_row_4_), .Y(u2_u0__abc_47660_n482) );
  INVX1 INVX1_606 ( .A(u2_u0_b1_last_row_0_), .Y(u2_u0__abc_47660_n486) );
  INVX1 INVX1_607 ( .A(u2_u0_b1_last_row_5_), .Y(u2_u0__abc_47660_n491) );
  INVX1 INVX1_608 ( .A(u2_u0_b1_last_row_10_), .Y(u2_u0__abc_47660_n497) );
  INVX1 INVX1_609 ( .A(u2_u0_b1_last_row_8_), .Y(u2_u0__abc_47660_n502) );
  INVX1 INVX1_61 ( .A(lmr_req), .Y(u0__abc_49347_n5740) );
  INVX1 INVX1_610 ( .A(u2_u0_b1_last_row_2_), .Y(u2_u0__abc_47660_n507) );
  INVX1 INVX1_611 ( .A(u2_u0_b1_last_row_1_), .Y(u2_u0__abc_47660_n510) );
  INVX1 INVX1_612 ( .A(u2_u0_b1_last_row_3_), .Y(u2_u0__abc_47660_n515) );
  INVX1 INVX1_613 ( .A(u2_u0_b1_last_row_6_), .Y(u2_u0__abc_47660_n520) );
  INVX1 INVX1_614 ( .A(u2_u0_b3_last_row_9_), .Y(u2_u0__abc_47660_n527) );
  INVX1 INVX1_615 ( .A(u2_u0_b3_last_row_11_), .Y(u2_u0__abc_47660_n534) );
  INVX1 INVX1_616 ( .A(u2_u0_b3_last_row_8_), .Y(u2_u0__abc_47660_n538) );
  INVX1 INVX1_617 ( .A(u2_u0_b3_last_row_4_), .Y(u2_u0__abc_47660_n544) );
  INVX1 INVX1_618 ( .A(u2_u0_b3_last_row_3_), .Y(u2_u0__abc_47660_n547) );
  INVX1 INVX1_619 ( .A(u2_u0_b3_last_row_0_), .Y(u2_u0__abc_47660_n551) );
  INVX1 INVX1_62 ( .A(init_ack), .Y(u0__abc_49347_n5742) );
  INVX1 INVX1_620 ( .A(u2_u0_b3_last_row_2_), .Y(u2_u0__abc_47660_n555) );
  INVX1 INVX1_621 ( .A(u2_u0_b3_last_row_7_), .Y(u2_u0__abc_47660_n563) );
  INVX1 INVX1_622 ( .A(u2_u0_b3_last_row_10_), .Y(u2_u0__abc_47660_n566) );
  INVX1 INVX1_623 ( .A(u2_u0_b3_last_row_6_), .Y(u2_u0__abc_47660_n572) );
  INVX1 INVX1_624 ( .A(u2_u0_b3_last_row_5_), .Y(u2_u0__abc_47660_n575) );
  INVX1 INVX1_625 ( .A(u2_u0_b3_last_row_1_), .Y(u2_u0__abc_47660_n581) );
  INVX1 INVX1_626 ( .A(u2_u0_b3_last_row_12_), .Y(u2_u0__abc_47660_n585) );
  INVX1 INVX1_627 ( .A(u2_u0__abc_47660_n604), .Y(u2_u0__abc_47660_n605) );
  INVX1 INVX1_628 ( .A(u2_bank_clr_all_0), .Y(u2_u0__abc_47660_n606) );
  INVX1 INVX1_629 ( .A(u2_bank_clr_0), .Y(u2_u0__abc_47660_n610) );
  INVX1 INVX1_63 ( .A(lmr_ack), .Y(u0__abc_49347_n5744) );
  INVX1 INVX1_630 ( .A(u2_u0__abc_47660_n204), .Y(u2_u0__abc_47660_n611) );
  INVX1 INVX1_631 ( .A(u2_u0__abc_47660_n247), .Y(u2_u0__abc_47660_n616) );
  INVX1 INVX1_632 ( .A(u2_u0__abc_47660_n289), .Y(u2_u0__abc_47660_n621) );
  INVX1 INVX1_633 ( .A(u2_u1__abc_47660_n140), .Y(u2_u1__abc_47660_n141) );
  INVX1 INVX1_634 ( .A(u2_u1__abc_47660_n145), .Y(u2_u1__abc_47660_n146) );
  INVX1 INVX1_635 ( .A(u2_u1__abc_47660_n150), .Y(u2_u1__abc_47660_n151) );
  INVX1 INVX1_636 ( .A(u2_u1__abc_47660_n155), .Y(u2_u1__abc_47660_n156) );
  INVX1 INVX1_637 ( .A(u2_u1__abc_47660_n160), .Y(u2_u1__abc_47660_n161) );
  INVX1 INVX1_638 ( .A(u2_u1__abc_47660_n165), .Y(u2_u1__abc_47660_n166) );
  INVX1 INVX1_639 ( .A(u2_u1__abc_47660_n170), .Y(u2_u1__abc_47660_n171) );
  INVX1 INVX1_64 ( .A(u0_u0__abc_43300_n202_1), .Y(u0_u0__abc_43300_n203) );
  INVX1 INVX1_640 ( .A(u2_u1__abc_47660_n175), .Y(u2_u1__abc_47660_n176) );
  INVX1 INVX1_641 ( .A(u2_u1__abc_47660_n180), .Y(u2_u1__abc_47660_n181) );
  INVX1 INVX1_642 ( .A(u2_u1__abc_47660_n185), .Y(u2_u1__abc_47660_n186) );
  INVX1 INVX1_643 ( .A(u2_u1__abc_47660_n190), .Y(u2_u1__abc_47660_n191) );
  INVX1 INVX1_644 ( .A(u2_u1__abc_47660_n195), .Y(u2_u1__abc_47660_n196) );
  INVX1 INVX1_645 ( .A(u2_u1__abc_47660_n200), .Y(u2_u1__abc_47660_n201) );
  INVX1 INVX1_646 ( .A(bank_adr_0_bF_buf1), .Y(u2_u1__abc_47660_n203) );
  INVX1 INVX1_647 ( .A(bank_adr_1_bF_buf0), .Y(u2_u1__abc_47660_n246) );
  INVX1 INVX1_648 ( .A(u2_u1_b0_last_row_12_), .Y(u2_u1__abc_47660_n331) );
  INVX1 INVX1_649 ( .A(u2_u1_b0_last_row_11_), .Y(u2_u1__abc_47660_n333) );
  INVX1 INVX1_65 ( .A(u0_u0__abc_43300_n204_1), .Y(u0_u0__abc_43300_n206) );
  INVX1 INVX1_650 ( .A(u2_u1_b0_last_row_9_), .Y(u2_u1__abc_47660_n339) );
  INVX1 INVX1_651 ( .A(u2_u1_b0_last_row_7_), .Y(u2_u1__abc_47660_n343) );
  INVX1 INVX1_652 ( .A(u2_u1_b0_last_row_4_), .Y(u2_u1__abc_47660_n351) );
  INVX1 INVX1_653 ( .A(u2_u1_b0_last_row_0_), .Y(u2_u1__abc_47660_n355) );
  INVX1 INVX1_654 ( .A(u2_u1_b0_last_row_5_), .Y(u2_u1__abc_47660_n360) );
  INVX1 INVX1_655 ( .A(u2_u1_b0_last_row_10_), .Y(u2_u1__abc_47660_n366) );
  INVX1 INVX1_656 ( .A(u2_u1_b0_last_row_8_), .Y(u2_u1__abc_47660_n371) );
  INVX1 INVX1_657 ( .A(u2_u1_b0_last_row_2_), .Y(u2_u1__abc_47660_n376) );
  INVX1 INVX1_658 ( .A(u2_u1_b0_last_row_1_), .Y(u2_u1__abc_47660_n379) );
  INVX1 INVX1_659 ( .A(u2_u1_b0_last_row_3_), .Y(u2_u1__abc_47660_n384) );
  INVX1 INVX1_66 ( .A(u0_lmr_ack0), .Y(u0_u0__abc_43300_n207_1) );
  INVX1 INVX1_660 ( .A(u2_u1_b0_last_row_6_), .Y(u2_u1__abc_47660_n389) );
  INVX1 INVX1_661 ( .A(u2_u1_b2_last_row_12_), .Y(u2_u1__abc_47660_n396) );
  INVX1 INVX1_662 ( .A(u2_u1_b2_last_row_11_), .Y(u2_u1__abc_47660_n398) );
  INVX1 INVX1_663 ( .A(u2_u1_b2_last_row_9_), .Y(u2_u1__abc_47660_n404) );
  INVX1 INVX1_664 ( .A(u2_u1_b2_last_row_7_), .Y(u2_u1__abc_47660_n408) );
  INVX1 INVX1_665 ( .A(u2_u1_b2_last_row_4_), .Y(u2_u1__abc_47660_n416) );
  INVX1 INVX1_666 ( .A(u2_u1_b2_last_row_0_), .Y(u2_u1__abc_47660_n420) );
  INVX1 INVX1_667 ( .A(u2_u1_b2_last_row_5_), .Y(u2_u1__abc_47660_n425) );
  INVX1 INVX1_668 ( .A(u2_u1_b2_last_row_10_), .Y(u2_u1__abc_47660_n431) );
  INVX1 INVX1_669 ( .A(u2_u1_b2_last_row_8_), .Y(u2_u1__abc_47660_n436) );
  INVX1 INVX1_67 ( .A(u0_u0__abc_43300_n213_1), .Y(u0_u0__abc_43300_n214_1) );
  INVX1 INVX1_670 ( .A(u2_u1_b2_last_row_2_), .Y(u2_u1__abc_47660_n441) );
  INVX1 INVX1_671 ( .A(u2_u1_b2_last_row_1_), .Y(u2_u1__abc_47660_n444) );
  INVX1 INVX1_672 ( .A(u2_u1_b2_last_row_3_), .Y(u2_u1__abc_47660_n449) );
  INVX1 INVX1_673 ( .A(u2_u1_b2_last_row_6_), .Y(u2_u1__abc_47660_n454) );
  INVX1 INVX1_674 ( .A(u2_u1_b1_last_row_12_), .Y(u2_u1__abc_47660_n462) );
  INVX1 INVX1_675 ( .A(u2_u1_b1_last_row_11_), .Y(u2_u1__abc_47660_n464) );
  INVX1 INVX1_676 ( .A(u2_u1_b1_last_row_9_), .Y(u2_u1__abc_47660_n470) );
  INVX1 INVX1_677 ( .A(u2_u1_b1_last_row_7_), .Y(u2_u1__abc_47660_n474) );
  INVX1 INVX1_678 ( .A(u2_u1_b1_last_row_4_), .Y(u2_u1__abc_47660_n482) );
  INVX1 INVX1_679 ( .A(u2_u1_b1_last_row_0_), .Y(u2_u1__abc_47660_n486) );
  INVX1 INVX1_68 ( .A(u0_u0_addr_r_2_), .Y(u0_u0__abc_43300_n347) );
  INVX1 INVX1_680 ( .A(u2_u1_b1_last_row_5_), .Y(u2_u1__abc_47660_n491) );
  INVX1 INVX1_681 ( .A(u2_u1_b1_last_row_10_), .Y(u2_u1__abc_47660_n497) );
  INVX1 INVX1_682 ( .A(u2_u1_b1_last_row_8_), .Y(u2_u1__abc_47660_n502) );
  INVX1 INVX1_683 ( .A(u2_u1_b1_last_row_2_), .Y(u2_u1__abc_47660_n507) );
  INVX1 INVX1_684 ( .A(u2_u1_b1_last_row_1_), .Y(u2_u1__abc_47660_n510) );
  INVX1 INVX1_685 ( .A(u2_u1_b1_last_row_3_), .Y(u2_u1__abc_47660_n515) );
  INVX1 INVX1_686 ( .A(u2_u1_b1_last_row_6_), .Y(u2_u1__abc_47660_n520) );
  INVX1 INVX1_687 ( .A(u2_u1_b3_last_row_9_), .Y(u2_u1__abc_47660_n527) );
  INVX1 INVX1_688 ( .A(u2_u1_b3_last_row_11_), .Y(u2_u1__abc_47660_n534) );
  INVX1 INVX1_689 ( .A(u2_u1_b3_last_row_8_), .Y(u2_u1__abc_47660_n538) );
  INVX1 INVX1_69 ( .A(u0_u0__abc_43300_n480), .Y(u0_u0__abc_43300_n481) );
  INVX1 INVX1_690 ( .A(u2_u1_b3_last_row_4_), .Y(u2_u1__abc_47660_n544) );
  INVX1 INVX1_691 ( .A(u2_u1_b3_last_row_3_), .Y(u2_u1__abc_47660_n547) );
  INVX1 INVX1_692 ( .A(u2_u1_b3_last_row_0_), .Y(u2_u1__abc_47660_n551) );
  INVX1 INVX1_693 ( .A(u2_u1_b3_last_row_2_), .Y(u2_u1__abc_47660_n555) );
  INVX1 INVX1_694 ( .A(u2_u1_b3_last_row_7_), .Y(u2_u1__abc_47660_n563) );
  INVX1 INVX1_695 ( .A(u2_u1_b3_last_row_10_), .Y(u2_u1__abc_47660_n566) );
  INVX1 INVX1_696 ( .A(u2_u1_b3_last_row_6_), .Y(u2_u1__abc_47660_n572) );
  INVX1 INVX1_697 ( .A(u2_u1_b3_last_row_5_), .Y(u2_u1__abc_47660_n575) );
  INVX1 INVX1_698 ( .A(u2_u1_b3_last_row_1_), .Y(u2_u1__abc_47660_n581) );
  INVX1 INVX1_699 ( .A(u2_u1_b3_last_row_12_), .Y(u2_u1__abc_47660_n585) );
  INVX1 INVX1_7 ( .A(u0__abc_49347_n1129), .Y(u0__abc_49347_n1134_1) );
  INVX1 INVX1_70 ( .A(u0_u0__abc_43300_n484), .Y(u0_u0__abc_43300_n485) );
  INVX1 INVX1_700 ( .A(u2_u1__abc_47660_n604), .Y(u2_u1__abc_47660_n605) );
  INVX1 INVX1_701 ( .A(u2_bank_clr_all_1), .Y(u2_u1__abc_47660_n606) );
  INVX1 INVX1_702 ( .A(u2_bank_clr_1), .Y(u2_u1__abc_47660_n610) );
  INVX1 INVX1_703 ( .A(u2_u1__abc_47660_n204), .Y(u2_u1__abc_47660_n611) );
  INVX1 INVX1_704 ( .A(u2_u1__abc_47660_n247), .Y(u2_u1__abc_47660_n616) );
  INVX1 INVX1_705 ( .A(u2_u1__abc_47660_n289), .Y(u2_u1__abc_47660_n621) );
  INVX1 INVX1_706 ( .A(u2_u2__abc_47660_n140), .Y(u2_u2__abc_47660_n141) );
  INVX1 INVX1_707 ( .A(u2_u2__abc_47660_n145), .Y(u2_u2__abc_47660_n146) );
  INVX1 INVX1_708 ( .A(u2_u2__abc_47660_n150), .Y(u2_u2__abc_47660_n151) );
  INVX1 INVX1_709 ( .A(u2_u2__abc_47660_n155), .Y(u2_u2__abc_47660_n156) );
  INVX1 INVX1_71 ( .A(wb_addr_i_23_bF_buf3), .Y(u0_u0__abc_43300_n488) );
  INVX1 INVX1_710 ( .A(u2_u2__abc_47660_n160), .Y(u2_u2__abc_47660_n161) );
  INVX1 INVX1_711 ( .A(u2_u2__abc_47660_n165), .Y(u2_u2__abc_47660_n166) );
  INVX1 INVX1_712 ( .A(u2_u2__abc_47660_n170), .Y(u2_u2__abc_47660_n171) );
  INVX1 INVX1_713 ( .A(u2_u2__abc_47660_n175), .Y(u2_u2__abc_47660_n176) );
  INVX1 INVX1_714 ( .A(u2_u2__abc_47660_n180), .Y(u2_u2__abc_47660_n181) );
  INVX1 INVX1_715 ( .A(u2_u2__abc_47660_n185), .Y(u2_u2__abc_47660_n186) );
  INVX1 INVX1_716 ( .A(u2_u2__abc_47660_n190), .Y(u2_u2__abc_47660_n191) );
  INVX1 INVX1_717 ( .A(u2_u2__abc_47660_n195), .Y(u2_u2__abc_47660_n196) );
  INVX1 INVX1_718 ( .A(u2_u2__abc_47660_n200), .Y(u2_u2__abc_47660_n201) );
  INVX1 INVX1_719 ( .A(bank_adr_0_bF_buf2), .Y(u2_u2__abc_47660_n203) );
  INVX1 INVX1_72 ( .A(u0_u0__abc_43300_n490), .Y(u0_u0__abc_43300_n491) );
  INVX1 INVX1_720 ( .A(bank_adr_1_bF_buf1), .Y(u2_u2__abc_47660_n246) );
  INVX1 INVX1_721 ( .A(u2_u2_b0_last_row_12_), .Y(u2_u2__abc_47660_n331) );
  INVX1 INVX1_722 ( .A(u2_u2_b0_last_row_11_), .Y(u2_u2__abc_47660_n333) );
  INVX1 INVX1_723 ( .A(u2_u2_b0_last_row_9_), .Y(u2_u2__abc_47660_n339) );
  INVX1 INVX1_724 ( .A(u2_u2_b0_last_row_7_), .Y(u2_u2__abc_47660_n343) );
  INVX1 INVX1_725 ( .A(u2_u2_b0_last_row_4_), .Y(u2_u2__abc_47660_n351) );
  INVX1 INVX1_726 ( .A(u2_u2_b0_last_row_0_), .Y(u2_u2__abc_47660_n355) );
  INVX1 INVX1_727 ( .A(u2_u2_b0_last_row_5_), .Y(u2_u2__abc_47660_n360) );
  INVX1 INVX1_728 ( .A(u2_u2_b0_last_row_10_), .Y(u2_u2__abc_47660_n366) );
  INVX1 INVX1_729 ( .A(u2_u2_b0_last_row_8_), .Y(u2_u2__abc_47660_n371) );
  INVX1 INVX1_73 ( .A(u0_u0__abc_43300_n483), .Y(u0_u0__abc_43300_n492) );
  INVX1 INVX1_730 ( .A(u2_u2_b0_last_row_2_), .Y(u2_u2__abc_47660_n376) );
  INVX1 INVX1_731 ( .A(u2_u2_b0_last_row_1_), .Y(u2_u2__abc_47660_n379) );
  INVX1 INVX1_732 ( .A(u2_u2_b0_last_row_3_), .Y(u2_u2__abc_47660_n384) );
  INVX1 INVX1_733 ( .A(u2_u2_b0_last_row_6_), .Y(u2_u2__abc_47660_n389) );
  INVX1 INVX1_734 ( .A(u2_u2_b2_last_row_12_), .Y(u2_u2__abc_47660_n396) );
  INVX1 INVX1_735 ( .A(u2_u2_b2_last_row_11_), .Y(u2_u2__abc_47660_n398) );
  INVX1 INVX1_736 ( .A(u2_u2_b2_last_row_9_), .Y(u2_u2__abc_47660_n404) );
  INVX1 INVX1_737 ( .A(u2_u2_b2_last_row_7_), .Y(u2_u2__abc_47660_n408) );
  INVX1 INVX1_738 ( .A(u2_u2_b2_last_row_4_), .Y(u2_u2__abc_47660_n416) );
  INVX1 INVX1_739 ( .A(u2_u2_b2_last_row_0_), .Y(u2_u2__abc_47660_n420) );
  INVX1 INVX1_74 ( .A(u0_u0__abc_43300_n497), .Y(u0_u0__abc_43300_n498) );
  INVX1 INVX1_740 ( .A(u2_u2_b2_last_row_5_), .Y(u2_u2__abc_47660_n425) );
  INVX1 INVX1_741 ( .A(u2_u2_b2_last_row_10_), .Y(u2_u2__abc_47660_n431) );
  INVX1 INVX1_742 ( .A(u2_u2_b2_last_row_8_), .Y(u2_u2__abc_47660_n436) );
  INVX1 INVX1_743 ( .A(u2_u2_b2_last_row_2_), .Y(u2_u2__abc_47660_n441) );
  INVX1 INVX1_744 ( .A(u2_u2_b2_last_row_1_), .Y(u2_u2__abc_47660_n444) );
  INVX1 INVX1_745 ( .A(u2_u2_b2_last_row_3_), .Y(u2_u2__abc_47660_n449) );
  INVX1 INVX1_746 ( .A(u2_u2_b2_last_row_6_), .Y(u2_u2__abc_47660_n454) );
  INVX1 INVX1_747 ( .A(u2_u2_b1_last_row_12_), .Y(u2_u2__abc_47660_n462) );
  INVX1 INVX1_748 ( .A(u2_u2_b1_last_row_11_), .Y(u2_u2__abc_47660_n464) );
  INVX1 INVX1_749 ( .A(u2_u2_b1_last_row_9_), .Y(u2_u2__abc_47660_n470) );
  INVX1 INVX1_75 ( .A(u0_u0__abc_43300_n501), .Y(u0_u0__abc_43300_n502) );
  INVX1 INVX1_750 ( .A(u2_u2_b1_last_row_7_), .Y(u2_u2__abc_47660_n474) );
  INVX1 INVX1_751 ( .A(u2_u2_b1_last_row_4_), .Y(u2_u2__abc_47660_n482) );
  INVX1 INVX1_752 ( .A(u2_u2_b1_last_row_0_), .Y(u2_u2__abc_47660_n486) );
  INVX1 INVX1_753 ( .A(u2_u2_b1_last_row_5_), .Y(u2_u2__abc_47660_n491) );
  INVX1 INVX1_754 ( .A(u2_u2_b1_last_row_10_), .Y(u2_u2__abc_47660_n497) );
  INVX1 INVX1_755 ( .A(u2_u2_b1_last_row_8_), .Y(u2_u2__abc_47660_n502) );
  INVX1 INVX1_756 ( .A(u2_u2_b1_last_row_2_), .Y(u2_u2__abc_47660_n507) );
  INVX1 INVX1_757 ( .A(u2_u2_b1_last_row_1_), .Y(u2_u2__abc_47660_n510) );
  INVX1 INVX1_758 ( .A(u2_u2_b1_last_row_3_), .Y(u2_u2__abc_47660_n515) );
  INVX1 INVX1_759 ( .A(u2_u2_b1_last_row_6_), .Y(u2_u2__abc_47660_n520) );
  INVX1 INVX1_76 ( .A(wb_addr_i_25_bF_buf2), .Y(u0_u0__abc_43300_n505) );
  INVX1 INVX1_760 ( .A(u2_u2_b3_last_row_9_), .Y(u2_u2__abc_47660_n527) );
  INVX1 INVX1_761 ( .A(u2_u2_b3_last_row_11_), .Y(u2_u2__abc_47660_n534) );
  INVX1 INVX1_762 ( .A(u2_u2_b3_last_row_8_), .Y(u2_u2__abc_47660_n538) );
  INVX1 INVX1_763 ( .A(u2_u2_b3_last_row_4_), .Y(u2_u2__abc_47660_n544) );
  INVX1 INVX1_764 ( .A(u2_u2_b3_last_row_3_), .Y(u2_u2__abc_47660_n547) );
  INVX1 INVX1_765 ( .A(u2_u2_b3_last_row_0_), .Y(u2_u2__abc_47660_n551) );
  INVX1 INVX1_766 ( .A(u2_u2_b3_last_row_2_), .Y(u2_u2__abc_47660_n555) );
  INVX1 INVX1_767 ( .A(u2_u2_b3_last_row_7_), .Y(u2_u2__abc_47660_n563) );
  INVX1 INVX1_768 ( .A(u2_u2_b3_last_row_10_), .Y(u2_u2__abc_47660_n566) );
  INVX1 INVX1_769 ( .A(u2_u2_b3_last_row_6_), .Y(u2_u2__abc_47660_n572) );
  INVX1 INVX1_77 ( .A(u0_u0__abc_43300_n506), .Y(u0_u0__abc_43300_n507) );
  INVX1 INVX1_770 ( .A(u2_u2_b3_last_row_5_), .Y(u2_u2__abc_47660_n575) );
  INVX1 INVX1_771 ( .A(u2_u2_b3_last_row_1_), .Y(u2_u2__abc_47660_n581) );
  INVX1 INVX1_772 ( .A(u2_u2_b3_last_row_12_), .Y(u2_u2__abc_47660_n585) );
  INVX1 INVX1_773 ( .A(u2_u2__abc_47660_n604), .Y(u2_u2__abc_47660_n605) );
  INVX1 INVX1_774 ( .A(u2_bank_clr_all_2), .Y(u2_u2__abc_47660_n606) );
  INVX1 INVX1_775 ( .A(u2_bank_clr_2), .Y(u2_u2__abc_47660_n610) );
  INVX1 INVX1_776 ( .A(u2_u2__abc_47660_n204), .Y(u2_u2__abc_47660_n611) );
  INVX1 INVX1_777 ( .A(u2_u2__abc_47660_n247), .Y(u2_u2__abc_47660_n616) );
  INVX1 INVX1_778 ( .A(u2_u2__abc_47660_n289), .Y(u2_u2__abc_47660_n621) );
  INVX1 INVX1_779 ( .A(u2_u3__abc_47660_n140), .Y(u2_u3__abc_47660_n141) );
  INVX1 INVX1_78 ( .A(u0_u0__abc_43300_n500), .Y(u0_u0__abc_43300_n508) );
  INVX1 INVX1_780 ( .A(u2_u3__abc_47660_n145), .Y(u2_u3__abc_47660_n146) );
  INVX1 INVX1_781 ( .A(u2_u3__abc_47660_n150), .Y(u2_u3__abc_47660_n151) );
  INVX1 INVX1_782 ( .A(u2_u3__abc_47660_n155), .Y(u2_u3__abc_47660_n156) );
  INVX1 INVX1_783 ( .A(u2_u3__abc_47660_n160), .Y(u2_u3__abc_47660_n161) );
  INVX1 INVX1_784 ( .A(u2_u3__abc_47660_n165), .Y(u2_u3__abc_47660_n166) );
  INVX1 INVX1_785 ( .A(u2_u3__abc_47660_n170), .Y(u2_u3__abc_47660_n171) );
  INVX1 INVX1_786 ( .A(u2_u3__abc_47660_n175), .Y(u2_u3__abc_47660_n176) );
  INVX1 INVX1_787 ( .A(u2_u3__abc_47660_n180), .Y(u2_u3__abc_47660_n181) );
  INVX1 INVX1_788 ( .A(u2_u3__abc_47660_n185), .Y(u2_u3__abc_47660_n186) );
  INVX1 INVX1_789 ( .A(u2_u3__abc_47660_n190), .Y(u2_u3__abc_47660_n191) );
  INVX1 INVX1_79 ( .A(u0_u0__abc_43300_n513), .Y(u0_u0__abc_43300_n514) );
  INVX1 INVX1_790 ( .A(u2_u3__abc_47660_n195), .Y(u2_u3__abc_47660_n196) );
  INVX1 INVX1_791 ( .A(u2_u3__abc_47660_n200), .Y(u2_u3__abc_47660_n201) );
  INVX1 INVX1_792 ( .A(bank_adr_0_bF_buf3), .Y(u2_u3__abc_47660_n203) );
  INVX1 INVX1_793 ( .A(bank_adr_1_bF_buf2), .Y(u2_u3__abc_47660_n246) );
  INVX1 INVX1_794 ( .A(u2_u3_b0_last_row_12_), .Y(u2_u3__abc_47660_n331) );
  INVX1 INVX1_795 ( .A(u2_u3_b0_last_row_11_), .Y(u2_u3__abc_47660_n333) );
  INVX1 INVX1_796 ( .A(u2_u3_b0_last_row_9_), .Y(u2_u3__abc_47660_n339) );
  INVX1 INVX1_797 ( .A(u2_u3_b0_last_row_7_), .Y(u2_u3__abc_47660_n343) );
  INVX1 INVX1_798 ( .A(u2_u3_b0_last_row_4_), .Y(u2_u3__abc_47660_n351) );
  INVX1 INVX1_799 ( .A(u2_u3_b0_last_row_0_), .Y(u2_u3__abc_47660_n355) );
  INVX1 INVX1_8 ( .A(u0__abc_49347_n1139_1), .Y(u0__abc_49347_n1148) );
  INVX1 INVX1_80 ( .A(u0_u0__abc_43300_n515), .Y(u0_u0__abc_43300_n516) );
  INVX1 INVX1_800 ( .A(u2_u3_b0_last_row_5_), .Y(u2_u3__abc_47660_n360) );
  INVX1 INVX1_801 ( .A(u2_u3_b0_last_row_10_), .Y(u2_u3__abc_47660_n366) );
  INVX1 INVX1_802 ( .A(u2_u3_b0_last_row_8_), .Y(u2_u3__abc_47660_n371) );
  INVX1 INVX1_803 ( .A(u2_u3_b0_last_row_2_), .Y(u2_u3__abc_47660_n376) );
  INVX1 INVX1_804 ( .A(u2_u3_b0_last_row_1_), .Y(u2_u3__abc_47660_n379) );
  INVX1 INVX1_805 ( .A(u2_u3_b0_last_row_3_), .Y(u2_u3__abc_47660_n384) );
  INVX1 INVX1_806 ( .A(u2_u3_b0_last_row_6_), .Y(u2_u3__abc_47660_n389) );
  INVX1 INVX1_807 ( .A(u2_u3_b2_last_row_12_), .Y(u2_u3__abc_47660_n396) );
  INVX1 INVX1_808 ( .A(u2_u3_b2_last_row_11_), .Y(u2_u3__abc_47660_n398) );
  INVX1 INVX1_809 ( .A(u2_u3_b2_last_row_9_), .Y(u2_u3__abc_47660_n404) );
  INVX1 INVX1_81 ( .A(u0_u0__abc_43300_n517), .Y(u0_u0__abc_43300_n520) );
  INVX1 INVX1_810 ( .A(u2_u3_b2_last_row_7_), .Y(u2_u3__abc_47660_n408) );
  INVX1 INVX1_811 ( .A(u2_u3_b2_last_row_4_), .Y(u2_u3__abc_47660_n416) );
  INVX1 INVX1_812 ( .A(u2_u3_b2_last_row_0_), .Y(u2_u3__abc_47660_n420) );
  INVX1 INVX1_813 ( .A(u2_u3_b2_last_row_5_), .Y(u2_u3__abc_47660_n425) );
  INVX1 INVX1_814 ( .A(u2_u3_b2_last_row_10_), .Y(u2_u3__abc_47660_n431) );
  INVX1 INVX1_815 ( .A(u2_u3_b2_last_row_8_), .Y(u2_u3__abc_47660_n436) );
  INVX1 INVX1_816 ( .A(u2_u3_b2_last_row_2_), .Y(u2_u3__abc_47660_n441) );
  INVX1 INVX1_817 ( .A(u2_u3_b2_last_row_1_), .Y(u2_u3__abc_47660_n444) );
  INVX1 INVX1_818 ( .A(u2_u3_b2_last_row_3_), .Y(u2_u3__abc_47660_n449) );
  INVX1 INVX1_819 ( .A(u2_u3_b2_last_row_6_), .Y(u2_u3__abc_47660_n454) );
  INVX1 INVX1_82 ( .A(u0_u0__abc_43300_n524), .Y(u0_u0__abc_43300_n525) );
  INVX1 INVX1_820 ( .A(u2_u3_b1_last_row_12_), .Y(u2_u3__abc_47660_n462) );
  INVX1 INVX1_821 ( .A(u2_u3_b1_last_row_11_), .Y(u2_u3__abc_47660_n464) );
  INVX1 INVX1_822 ( .A(u2_u3_b1_last_row_9_), .Y(u2_u3__abc_47660_n470) );
  INVX1 INVX1_823 ( .A(u2_u3_b1_last_row_7_), .Y(u2_u3__abc_47660_n474) );
  INVX1 INVX1_824 ( .A(u2_u3_b1_last_row_4_), .Y(u2_u3__abc_47660_n482) );
  INVX1 INVX1_825 ( .A(u2_u3_b1_last_row_0_), .Y(u2_u3__abc_47660_n486) );
  INVX1 INVX1_826 ( .A(u2_u3_b1_last_row_5_), .Y(u2_u3__abc_47660_n491) );
  INVX1 INVX1_827 ( .A(u2_u3_b1_last_row_10_), .Y(u2_u3__abc_47660_n497) );
  INVX1 INVX1_828 ( .A(u2_u3_b1_last_row_8_), .Y(u2_u3__abc_47660_n502) );
  INVX1 INVX1_829 ( .A(u2_u3_b1_last_row_2_), .Y(u2_u3__abc_47660_n507) );
  INVX1 INVX1_83 ( .A(u0_u0__abc_43300_n528), .Y(u0_u0__abc_43300_n529) );
  INVX1 INVX1_830 ( .A(u2_u3_b1_last_row_1_), .Y(u2_u3__abc_47660_n510) );
  INVX1 INVX1_831 ( .A(u2_u3_b1_last_row_3_), .Y(u2_u3__abc_47660_n515) );
  INVX1 INVX1_832 ( .A(u2_u3_b1_last_row_6_), .Y(u2_u3__abc_47660_n520) );
  INVX1 INVX1_833 ( .A(u2_u3_b3_last_row_9_), .Y(u2_u3__abc_47660_n527) );
  INVX1 INVX1_834 ( .A(u2_u3_b3_last_row_11_), .Y(u2_u3__abc_47660_n534) );
  INVX1 INVX1_835 ( .A(u2_u3_b3_last_row_8_), .Y(u2_u3__abc_47660_n538) );
  INVX1 INVX1_836 ( .A(u2_u3_b3_last_row_4_), .Y(u2_u3__abc_47660_n544) );
  INVX1 INVX1_837 ( .A(u2_u3_b3_last_row_3_), .Y(u2_u3__abc_47660_n547) );
  INVX1 INVX1_838 ( .A(u2_u3_b3_last_row_0_), .Y(u2_u3__abc_47660_n551) );
  INVX1 INVX1_839 ( .A(u2_u3_b3_last_row_2_), .Y(u2_u3__abc_47660_n555) );
  INVX1 INVX1_84 ( .A(u0_u0__abc_43300_n533), .Y(u0_u0__abc_43300_n534) );
  INVX1 INVX1_840 ( .A(u2_u3_b3_last_row_7_), .Y(u2_u3__abc_47660_n563) );
  INVX1 INVX1_841 ( .A(u2_u3_b3_last_row_10_), .Y(u2_u3__abc_47660_n566) );
  INVX1 INVX1_842 ( .A(u2_u3_b3_last_row_6_), .Y(u2_u3__abc_47660_n572) );
  INVX1 INVX1_843 ( .A(u2_u3_b3_last_row_5_), .Y(u2_u3__abc_47660_n575) );
  INVX1 INVX1_844 ( .A(u2_u3_b3_last_row_1_), .Y(u2_u3__abc_47660_n581) );
  INVX1 INVX1_845 ( .A(u2_u3_b3_last_row_12_), .Y(u2_u3__abc_47660_n585) );
  INVX1 INVX1_846 ( .A(u2_u3__abc_47660_n604), .Y(u2_u3__abc_47660_n605) );
  INVX1 INVX1_847 ( .A(u2_bank_clr_all_3), .Y(u2_u3__abc_47660_n606) );
  INVX1 INVX1_848 ( .A(u2_bank_clr_3), .Y(u2_u3__abc_47660_n610) );
  INVX1 INVX1_849 ( .A(u2_u3__abc_47660_n204), .Y(u2_u3__abc_47660_n611) );
  INVX1 INVX1_85 ( .A(u0_u0__abc_43300_n527), .Y(u0_u0__abc_43300_n536) );
  INVX1 INVX1_850 ( .A(u2_u3__abc_47660_n247), .Y(u2_u3__abc_47660_n616) );
  INVX1 INVX1_851 ( .A(u2_u3__abc_47660_n289), .Y(u2_u3__abc_47660_n621) );
  INVX1 INVX1_852 ( .A(u2_u4__abc_47660_n140), .Y(u2_u4__abc_47660_n141) );
  INVX1 INVX1_853 ( .A(u2_u4__abc_47660_n145), .Y(u2_u4__abc_47660_n146) );
  INVX1 INVX1_854 ( .A(u2_u4__abc_47660_n150), .Y(u2_u4__abc_47660_n151) );
  INVX1 INVX1_855 ( .A(u2_u4__abc_47660_n155), .Y(u2_u4__abc_47660_n156) );
  INVX1 INVX1_856 ( .A(u2_u4__abc_47660_n160), .Y(u2_u4__abc_47660_n161) );
  INVX1 INVX1_857 ( .A(u2_u4__abc_47660_n165), .Y(u2_u4__abc_47660_n166) );
  INVX1 INVX1_858 ( .A(u2_u4__abc_47660_n170), .Y(u2_u4__abc_47660_n171) );
  INVX1 INVX1_859 ( .A(u2_u4__abc_47660_n175), .Y(u2_u4__abc_47660_n176) );
  INVX1 INVX1_86 ( .A(u0_u0__abc_43300_n532), .Y(u0_u0__abc_43300_n540) );
  INVX1 INVX1_860 ( .A(u2_u4__abc_47660_n180), .Y(u2_u4__abc_47660_n181) );
  INVX1 INVX1_861 ( .A(u2_u4__abc_47660_n185), .Y(u2_u4__abc_47660_n186) );
  INVX1 INVX1_862 ( .A(u2_u4__abc_47660_n190), .Y(u2_u4__abc_47660_n191) );
  INVX1 INVX1_863 ( .A(u2_u4__abc_47660_n195), .Y(u2_u4__abc_47660_n196) );
  INVX1 INVX1_864 ( .A(u2_u4__abc_47660_n200), .Y(u2_u4__abc_47660_n201) );
  INVX1 INVX1_865 ( .A(bank_adr_0_bF_buf0), .Y(u2_u4__abc_47660_n203) );
  INVX1 INVX1_866 ( .A(bank_adr_1_bF_buf3), .Y(u2_u4__abc_47660_n246) );
  INVX1 INVX1_867 ( .A(u2_u4_b0_last_row_12_), .Y(u2_u4__abc_47660_n331) );
  INVX1 INVX1_868 ( .A(u2_u4_b0_last_row_11_), .Y(u2_u4__abc_47660_n333) );
  INVX1 INVX1_869 ( .A(u2_u4_b0_last_row_9_), .Y(u2_u4__abc_47660_n339) );
  INVX1 INVX1_87 ( .A(u0_u0__abc_43300_n478), .Y(u0_u0__abc_43300_n546) );
  INVX1 INVX1_870 ( .A(u2_u4_b0_last_row_7_), .Y(u2_u4__abc_47660_n343) );
  INVX1 INVX1_871 ( .A(u2_u4_b0_last_row_4_), .Y(u2_u4__abc_47660_n351) );
  INVX1 INVX1_872 ( .A(u2_u4_b0_last_row_0_), .Y(u2_u4__abc_47660_n355) );
  INVX1 INVX1_873 ( .A(u2_u4_b0_last_row_5_), .Y(u2_u4__abc_47660_n360) );
  INVX1 INVX1_874 ( .A(u2_u4_b0_last_row_10_), .Y(u2_u4__abc_47660_n366) );
  INVX1 INVX1_875 ( .A(u2_u4_b0_last_row_8_), .Y(u2_u4__abc_47660_n371) );
  INVX1 INVX1_876 ( .A(u2_u4_b0_last_row_2_), .Y(u2_u4__abc_47660_n376) );
  INVX1 INVX1_877 ( .A(u2_u4_b0_last_row_1_), .Y(u2_u4__abc_47660_n379) );
  INVX1 INVX1_878 ( .A(u2_u4_b0_last_row_3_), .Y(u2_u4__abc_47660_n384) );
  INVX1 INVX1_879 ( .A(u2_u4_b0_last_row_6_), .Y(u2_u4__abc_47660_n389) );
  INVX1 INVX1_88 ( .A(u0_init_ack0), .Y(u0_u0__abc_43300_n549) );
  INVX1 INVX1_880 ( .A(u2_u4_b2_last_row_12_), .Y(u2_u4__abc_47660_n396) );
  INVX1 INVX1_881 ( .A(u2_u4_b2_last_row_11_), .Y(u2_u4__abc_47660_n398) );
  INVX1 INVX1_882 ( .A(u2_u4_b2_last_row_9_), .Y(u2_u4__abc_47660_n404) );
  INVX1 INVX1_883 ( .A(u2_u4_b2_last_row_7_), .Y(u2_u4__abc_47660_n408) );
  INVX1 INVX1_884 ( .A(u2_u4_b2_last_row_4_), .Y(u2_u4__abc_47660_n416) );
  INVX1 INVX1_885 ( .A(u2_u4_b2_last_row_0_), .Y(u2_u4__abc_47660_n420) );
  INVX1 INVX1_886 ( .A(u2_u4_b2_last_row_5_), .Y(u2_u4__abc_47660_n425) );
  INVX1 INVX1_887 ( .A(u2_u4_b2_last_row_10_), .Y(u2_u4__abc_47660_n431) );
  INVX1 INVX1_888 ( .A(u2_u4_b2_last_row_8_), .Y(u2_u4__abc_47660_n436) );
  INVX1 INVX1_889 ( .A(u2_u4_b2_last_row_2_), .Y(u2_u4__abc_47660_n441) );
  INVX1 INVX1_89 ( .A(u0_u0_inited), .Y(u0_u0__abc_43300_n551) );
  INVX1 INVX1_890 ( .A(u2_u4_b2_last_row_1_), .Y(u2_u4__abc_47660_n444) );
  INVX1 INVX1_891 ( .A(u2_u4_b2_last_row_3_), .Y(u2_u4__abc_47660_n449) );
  INVX1 INVX1_892 ( .A(u2_u4_b2_last_row_6_), .Y(u2_u4__abc_47660_n454) );
  INVX1 INVX1_893 ( .A(u2_u4_b1_last_row_12_), .Y(u2_u4__abc_47660_n462) );
  INVX1 INVX1_894 ( .A(u2_u4_b1_last_row_11_), .Y(u2_u4__abc_47660_n464) );
  INVX1 INVX1_895 ( .A(u2_u4_b1_last_row_9_), .Y(u2_u4__abc_47660_n470) );
  INVX1 INVX1_896 ( .A(u2_u4_b1_last_row_7_), .Y(u2_u4__abc_47660_n474) );
  INVX1 INVX1_897 ( .A(u2_u4_b1_last_row_4_), .Y(u2_u4__abc_47660_n482) );
  INVX1 INVX1_898 ( .A(u2_u4_b1_last_row_0_), .Y(u2_u4__abc_47660_n486) );
  INVX1 INVX1_899 ( .A(u2_u4_b1_last_row_5_), .Y(u2_u4__abc_47660_n491) );
  INVX1 INVX1_9 ( .A(u0__abc_49347_n1146), .Y(u0__abc_49347_n1153) );
  INVX1 INVX1_90 ( .A(u0_u1__abc_43657_n202), .Y(u0_u1__abc_43657_n203_1) );
  INVX1 INVX1_900 ( .A(u2_u4_b1_last_row_10_), .Y(u2_u4__abc_47660_n497) );
  INVX1 INVX1_901 ( .A(u2_u4_b1_last_row_8_), .Y(u2_u4__abc_47660_n502) );
  INVX1 INVX1_902 ( .A(u2_u4_b1_last_row_2_), .Y(u2_u4__abc_47660_n507) );
  INVX1 INVX1_903 ( .A(u2_u4_b1_last_row_1_), .Y(u2_u4__abc_47660_n510) );
  INVX1 INVX1_904 ( .A(u2_u4_b1_last_row_3_), .Y(u2_u4__abc_47660_n515) );
  INVX1 INVX1_905 ( .A(u2_u4_b1_last_row_6_), .Y(u2_u4__abc_47660_n520) );
  INVX1 INVX1_906 ( .A(u2_u4_b3_last_row_9_), .Y(u2_u4__abc_47660_n527) );
  INVX1 INVX1_907 ( .A(u2_u4_b3_last_row_11_), .Y(u2_u4__abc_47660_n534) );
  INVX1 INVX1_908 ( .A(u2_u4_b3_last_row_8_), .Y(u2_u4__abc_47660_n538) );
  INVX1 INVX1_909 ( .A(u2_u4_b3_last_row_4_), .Y(u2_u4__abc_47660_n544) );
  INVX1 INVX1_91 ( .A(u0_u1__abc_43657_n204_1), .Y(u0_u1__abc_43657_n206_1) );
  INVX1 INVX1_910 ( .A(u2_u4_b3_last_row_3_), .Y(u2_u4__abc_47660_n547) );
  INVX1 INVX1_911 ( .A(u2_u4_b3_last_row_0_), .Y(u2_u4__abc_47660_n551) );
  INVX1 INVX1_912 ( .A(u2_u4_b3_last_row_2_), .Y(u2_u4__abc_47660_n555) );
  INVX1 INVX1_913 ( .A(u2_u4_b3_last_row_7_), .Y(u2_u4__abc_47660_n563) );
  INVX1 INVX1_914 ( .A(u2_u4_b3_last_row_10_), .Y(u2_u4__abc_47660_n566) );
  INVX1 INVX1_915 ( .A(u2_u4_b3_last_row_6_), .Y(u2_u4__abc_47660_n572) );
  INVX1 INVX1_916 ( .A(u2_u4_b3_last_row_5_), .Y(u2_u4__abc_47660_n575) );
  INVX1 INVX1_917 ( .A(u2_u4_b3_last_row_1_), .Y(u2_u4__abc_47660_n581) );
  INVX1 INVX1_918 ( .A(u2_u4_b3_last_row_12_), .Y(u2_u4__abc_47660_n585) );
  INVX1 INVX1_919 ( .A(u2_u4__abc_47660_n604), .Y(u2_u4__abc_47660_n605) );
  INVX1 INVX1_92 ( .A(u0_lmr_ack1), .Y(u0_u1__abc_43657_n207_1) );
  INVX1 INVX1_920 ( .A(u2_bank_clr_all_4), .Y(u2_u4__abc_47660_n606) );
  INVX1 INVX1_921 ( .A(u2_bank_clr_4), .Y(u2_u4__abc_47660_n610) );
  INVX1 INVX1_922 ( .A(u2_u4__abc_47660_n204), .Y(u2_u4__abc_47660_n611) );
  INVX1 INVX1_923 ( .A(u2_u4__abc_47660_n247), .Y(u2_u4__abc_47660_n616) );
  INVX1 INVX1_924 ( .A(u2_u4__abc_47660_n289), .Y(u2_u4__abc_47660_n621) );
  INVX1 INVX1_925 ( .A(u2_u5__abc_47660_n140), .Y(u2_u5__abc_47660_n141) );
  INVX1 INVX1_926 ( .A(u2_u5__abc_47660_n145), .Y(u2_u5__abc_47660_n146) );
  INVX1 INVX1_927 ( .A(u2_u5__abc_47660_n150), .Y(u2_u5__abc_47660_n151) );
  INVX1 INVX1_928 ( .A(u2_u5__abc_47660_n155), .Y(u2_u5__abc_47660_n156) );
  INVX1 INVX1_929 ( .A(u2_u5__abc_47660_n160), .Y(u2_u5__abc_47660_n161) );
  INVX1 INVX1_93 ( .A(u0_u1_addr_r_6_), .Y(u0_u1__abc_43657_n211) );
  INVX1 INVX1_930 ( .A(u2_u5__abc_47660_n165), .Y(u2_u5__abc_47660_n166) );
  INVX1 INVX1_931 ( .A(u2_u5__abc_47660_n170), .Y(u2_u5__abc_47660_n171) );
  INVX1 INVX1_932 ( .A(u2_u5__abc_47660_n175), .Y(u2_u5__abc_47660_n176) );
  INVX1 INVX1_933 ( .A(u2_u5__abc_47660_n180), .Y(u2_u5__abc_47660_n181) );
  INVX1 INVX1_934 ( .A(u2_u5__abc_47660_n185), .Y(u2_u5__abc_47660_n186) );
  INVX1 INVX1_935 ( .A(u2_u5__abc_47660_n190), .Y(u2_u5__abc_47660_n191) );
  INVX1 INVX1_936 ( .A(u2_u5__abc_47660_n195), .Y(u2_u5__abc_47660_n196) );
  INVX1 INVX1_937 ( .A(u2_u5__abc_47660_n200), .Y(u2_u5__abc_47660_n201) );
  INVX1 INVX1_938 ( .A(bank_adr_0_bF_buf1), .Y(u2_u5__abc_47660_n203) );
  INVX1 INVX1_939 ( .A(bank_adr_1_bF_buf0), .Y(u2_u5__abc_47660_n246) );
  INVX1 INVX1_94 ( .A(u0_u1_addr_r_5_), .Y(u0_u1__abc_43657_n212_1) );
  INVX1 INVX1_940 ( .A(u2_u5_b0_last_row_12_), .Y(u2_u5__abc_47660_n331) );
  INVX1 INVX1_941 ( .A(u2_u5_b0_last_row_11_), .Y(u2_u5__abc_47660_n333) );
  INVX1 INVX1_942 ( .A(u2_u5_b0_last_row_9_), .Y(u2_u5__abc_47660_n339) );
  INVX1 INVX1_943 ( .A(u2_u5_b0_last_row_7_), .Y(u2_u5__abc_47660_n343) );
  INVX1 INVX1_944 ( .A(u2_u5_b0_last_row_4_), .Y(u2_u5__abc_47660_n351) );
  INVX1 INVX1_945 ( .A(u2_u5_b0_last_row_0_), .Y(u2_u5__abc_47660_n355) );
  INVX1 INVX1_946 ( .A(u2_u5_b0_last_row_5_), .Y(u2_u5__abc_47660_n360) );
  INVX1 INVX1_947 ( .A(u2_u5_b0_last_row_10_), .Y(u2_u5__abc_47660_n366) );
  INVX1 INVX1_948 ( .A(u2_u5_b0_last_row_8_), .Y(u2_u5__abc_47660_n371) );
  INVX1 INVX1_949 ( .A(u2_u5_b0_last_row_2_), .Y(u2_u5__abc_47660_n376) );
  INVX1 INVX1_95 ( .A(\wb_data_i[0] ), .Y(u0_u1__abc_43657_n220) );
  INVX1 INVX1_950 ( .A(u2_u5_b0_last_row_1_), .Y(u2_u5__abc_47660_n379) );
  INVX1 INVX1_951 ( .A(u2_u5_b0_last_row_3_), .Y(u2_u5__abc_47660_n384) );
  INVX1 INVX1_952 ( .A(u2_u5_b0_last_row_6_), .Y(u2_u5__abc_47660_n389) );
  INVX1 INVX1_953 ( .A(u2_u5_b2_last_row_12_), .Y(u2_u5__abc_47660_n396) );
  INVX1 INVX1_954 ( .A(u2_u5_b2_last_row_11_), .Y(u2_u5__abc_47660_n398) );
  INVX1 INVX1_955 ( .A(u2_u5_b2_last_row_9_), .Y(u2_u5__abc_47660_n404) );
  INVX1 INVX1_956 ( .A(u2_u5_b2_last_row_7_), .Y(u2_u5__abc_47660_n408) );
  INVX1 INVX1_957 ( .A(u2_u5_b2_last_row_4_), .Y(u2_u5__abc_47660_n416) );
  INVX1 INVX1_958 ( .A(u2_u5_b2_last_row_0_), .Y(u2_u5__abc_47660_n420) );
  INVX1 INVX1_959 ( .A(u2_u5_b2_last_row_5_), .Y(u2_u5__abc_47660_n425) );
  INVX1 INVX1_96 ( .A(u0_u1__abc_43657_n221_1), .Y(u0_u1__abc_43657_n222_1) );
  INVX1 INVX1_960 ( .A(u2_u5_b2_last_row_10_), .Y(u2_u5__abc_47660_n431) );
  INVX1 INVX1_961 ( .A(u2_u5_b2_last_row_8_), .Y(u2_u5__abc_47660_n436) );
  INVX1 INVX1_962 ( .A(u2_u5_b2_last_row_2_), .Y(u2_u5__abc_47660_n441) );
  INVX1 INVX1_963 ( .A(u2_u5_b2_last_row_1_), .Y(u2_u5__abc_47660_n444) );
  INVX1 INVX1_964 ( .A(u2_u5_b2_last_row_3_), .Y(u2_u5__abc_47660_n449) );
  INVX1 INVX1_965 ( .A(u2_u5_b2_last_row_6_), .Y(u2_u5__abc_47660_n454) );
  INVX1 INVX1_966 ( .A(u2_u5_b1_last_row_12_), .Y(u2_u5__abc_47660_n462) );
  INVX1 INVX1_967 ( .A(u2_u5_b1_last_row_11_), .Y(u2_u5__abc_47660_n464) );
  INVX1 INVX1_968 ( .A(u2_u5_b1_last_row_9_), .Y(u2_u5__abc_47660_n470) );
  INVX1 INVX1_969 ( .A(u2_u5_b1_last_row_7_), .Y(u2_u5__abc_47660_n474) );
  INVX1 INVX1_97 ( .A(\wb_data_i[1] ), .Y(u0_u1__abc_43657_n226) );
  INVX1 INVX1_970 ( .A(u2_u5_b1_last_row_4_), .Y(u2_u5__abc_47660_n482) );
  INVX1 INVX1_971 ( .A(u2_u5_b1_last_row_0_), .Y(u2_u5__abc_47660_n486) );
  INVX1 INVX1_972 ( .A(u2_u5_b1_last_row_5_), .Y(u2_u5__abc_47660_n491) );
  INVX1 INVX1_973 ( .A(u2_u5_b1_last_row_10_), .Y(u2_u5__abc_47660_n497) );
  INVX1 INVX1_974 ( .A(u2_u5_b1_last_row_8_), .Y(u2_u5__abc_47660_n502) );
  INVX1 INVX1_975 ( .A(u2_u5_b1_last_row_2_), .Y(u2_u5__abc_47660_n507) );
  INVX1 INVX1_976 ( .A(u2_u5_b1_last_row_1_), .Y(u2_u5__abc_47660_n510) );
  INVX1 INVX1_977 ( .A(u2_u5_b1_last_row_3_), .Y(u2_u5__abc_47660_n515) );
  INVX1 INVX1_978 ( .A(u2_u5_b1_last_row_6_), .Y(u2_u5__abc_47660_n520) );
  INVX1 INVX1_979 ( .A(u2_u5_b3_last_row_9_), .Y(u2_u5__abc_47660_n527) );
  INVX1 INVX1_98 ( .A(u0_u1__abc_43657_n227_1), .Y(u0_u1__abc_43657_n228_1) );
  INVX1 INVX1_980 ( .A(u2_u5_b3_last_row_11_), .Y(u2_u5__abc_47660_n534) );
  INVX1 INVX1_981 ( .A(u2_u5_b3_last_row_8_), .Y(u2_u5__abc_47660_n538) );
  INVX1 INVX1_982 ( .A(u2_u5_b3_last_row_4_), .Y(u2_u5__abc_47660_n544) );
  INVX1 INVX1_983 ( .A(u2_u5_b3_last_row_3_), .Y(u2_u5__abc_47660_n547) );
  INVX1 INVX1_984 ( .A(u2_u5_b3_last_row_0_), .Y(u2_u5__abc_47660_n551) );
  INVX1 INVX1_985 ( .A(u2_u5_b3_last_row_2_), .Y(u2_u5__abc_47660_n555) );
  INVX1 INVX1_986 ( .A(u2_u5_b3_last_row_7_), .Y(u2_u5__abc_47660_n563) );
  INVX1 INVX1_987 ( .A(u2_u5_b3_last_row_10_), .Y(u2_u5__abc_47660_n566) );
  INVX1 INVX1_988 ( .A(u2_u5_b3_last_row_6_), .Y(u2_u5__abc_47660_n572) );
  INVX1 INVX1_989 ( .A(u2_u5_b3_last_row_5_), .Y(u2_u5__abc_47660_n575) );
  INVX1 INVX1_99 ( .A(\wb_data_i[2] ), .Y(u0_u1__abc_43657_n232) );
  INVX1 INVX1_990 ( .A(u2_u5_b3_last_row_1_), .Y(u2_u5__abc_47660_n581) );
  INVX1 INVX1_991 ( .A(u2_u5_b3_last_row_12_), .Y(u2_u5__abc_47660_n585) );
  INVX1 INVX1_992 ( .A(u2_u5__abc_47660_n604), .Y(u2_u5__abc_47660_n605) );
  INVX1 INVX1_993 ( .A(u2_bank_clr_all_5), .Y(u2_u5__abc_47660_n606) );
  INVX1 INVX1_994 ( .A(u2_bank_clr_5), .Y(u2_u5__abc_47660_n610) );
  INVX1 INVX1_995 ( .A(u2_u5__abc_47660_n204), .Y(u2_u5__abc_47660_n611) );
  INVX1 INVX1_996 ( .A(u2_u5__abc_47660_n247), .Y(u2_u5__abc_47660_n616) );
  INVX1 INVX1_997 ( .A(u2_u5__abc_47660_n289), .Y(u2_u5__abc_47660_n621) );
  INVX1 INVX1_998 ( .A(u3__abc_46775_n281_1), .Y(u3__abc_46775_n282_1) );
  INVX1 INVX1_999 ( .A(u3__abc_46775_n283), .Y(u3__abc_46775_n284) );
  INVX2 INVX2_1 ( .A(init_req), .Y(u0__abc_49347_n1100_1) );
  INVX2 INVX2_10 ( .A(row_adr_7_bF_buf4), .Y(u2_u0__abc_47660_n174) );
  INVX2 INVX2_100 ( .A(u5__abc_54027_n654_1), .Y(u5__abc_54027_n655) );
  INVX2 INVX2_101 ( .A(u5__abc_54027_n657_1), .Y(u5__abc_54027_n658) );
  INVX2 INVX2_102 ( .A(u5__abc_54027_n702), .Y(u5__abc_54027_n703) );
  INVX2 INVX2_103 ( .A(u5__abc_54027_n850), .Y(u5__abc_54027_n892) );
  INVX2 INVX2_104 ( .A(u5__abc_54027_n1089), .Y(u5__abc_54027_n1090) );
  INVX2 INVX2_105 ( .A(u5__abc_54027_n1110), .Y(u5__abc_54027_n1111) );
  INVX2 INVX2_106 ( .A(u5__abc_54027_n1106), .Y(u5__abc_54027_n1124) );
  INVX2 INVX2_107 ( .A(u5_tmr2_done), .Y(u5__abc_54027_n1299) );
  INVX2 INVX2_108 ( .A(u7__abc_47535_n106), .Y(u7__abc_47535_n107) );
  INVX2 INVX2_109 ( .A(cs_en), .Y(u7__abc_47535_n114) );
  INVX2 INVX2_11 ( .A(row_adr_8_bF_buf4), .Y(u2_u0__abc_47660_n179) );
  INVX2 INVX2_12 ( .A(row_adr_9_bF_buf4), .Y(u2_u0__abc_47660_n184) );
  INVX2 INVX2_13 ( .A(row_adr_10_bF_buf4), .Y(u2_u0__abc_47660_n189) );
  INVX2 INVX2_14 ( .A(row_adr_11_bF_buf4), .Y(u2_u0__abc_47660_n194) );
  INVX2 INVX2_15 ( .A(row_adr_12_bF_buf4), .Y(u2_u0__abc_47660_n199) );
  INVX2 INVX2_16 ( .A(rst_i_bF_buf0), .Y(u2_u0__abc_47660_n305) );
  INVX2 INVX2_17 ( .A(row_adr_0_bF_buf3), .Y(u2_u1__abc_47660_n139) );
  INVX2 INVX2_18 ( .A(row_adr_1_bF_buf3), .Y(u2_u1__abc_47660_n144) );
  INVX2 INVX2_19 ( .A(row_adr_2_bF_buf3), .Y(u2_u1__abc_47660_n149) );
  INVX2 INVX2_2 ( .A(u0_sreq_cs_le), .Y(u0__abc_49347_n1113_1) );
  INVX2 INVX2_20 ( .A(row_adr_3_bF_buf3), .Y(u2_u1__abc_47660_n154) );
  INVX2 INVX2_21 ( .A(row_adr_4_bF_buf3), .Y(u2_u1__abc_47660_n159) );
  INVX2 INVX2_22 ( .A(row_adr_5_bF_buf3), .Y(u2_u1__abc_47660_n164) );
  INVX2 INVX2_23 ( .A(row_adr_6_bF_buf3), .Y(u2_u1__abc_47660_n169) );
  INVX2 INVX2_24 ( .A(row_adr_7_bF_buf3), .Y(u2_u1__abc_47660_n174) );
  INVX2 INVX2_25 ( .A(row_adr_8_bF_buf3), .Y(u2_u1__abc_47660_n179) );
  INVX2 INVX2_26 ( .A(row_adr_9_bF_buf3), .Y(u2_u1__abc_47660_n184) );
  INVX2 INVX2_27 ( .A(row_adr_10_bF_buf3), .Y(u2_u1__abc_47660_n189) );
  INVX2 INVX2_28 ( .A(row_adr_11_bF_buf3), .Y(u2_u1__abc_47660_n194) );
  INVX2 INVX2_29 ( .A(row_adr_12_bF_buf3), .Y(u2_u1__abc_47660_n199) );
  INVX2 INVX2_3 ( .A(row_adr_0_bF_buf4), .Y(u2_u0__abc_47660_n139) );
  INVX2 INVX2_30 ( .A(rst_i_bF_buf3), .Y(u2_u1__abc_47660_n305) );
  INVX2 INVX2_31 ( .A(row_adr_0_bF_buf2), .Y(u2_u2__abc_47660_n139) );
  INVX2 INVX2_32 ( .A(row_adr_1_bF_buf2), .Y(u2_u2__abc_47660_n144) );
  INVX2 INVX2_33 ( .A(row_adr_2_bF_buf2), .Y(u2_u2__abc_47660_n149) );
  INVX2 INVX2_34 ( .A(row_adr_3_bF_buf2), .Y(u2_u2__abc_47660_n154) );
  INVX2 INVX2_35 ( .A(row_adr_4_bF_buf2), .Y(u2_u2__abc_47660_n159) );
  INVX2 INVX2_36 ( .A(row_adr_5_bF_buf2), .Y(u2_u2__abc_47660_n164) );
  INVX2 INVX2_37 ( .A(row_adr_6_bF_buf2), .Y(u2_u2__abc_47660_n169) );
  INVX2 INVX2_38 ( .A(row_adr_7_bF_buf2), .Y(u2_u2__abc_47660_n174) );
  INVX2 INVX2_39 ( .A(row_adr_8_bF_buf2), .Y(u2_u2__abc_47660_n179) );
  INVX2 INVX2_4 ( .A(row_adr_1_bF_buf4), .Y(u2_u0__abc_47660_n144) );
  INVX2 INVX2_40 ( .A(row_adr_9_bF_buf2), .Y(u2_u2__abc_47660_n184) );
  INVX2 INVX2_41 ( .A(row_adr_10_bF_buf2), .Y(u2_u2__abc_47660_n189) );
  INVX2 INVX2_42 ( .A(row_adr_11_bF_buf2), .Y(u2_u2__abc_47660_n194) );
  INVX2 INVX2_43 ( .A(row_adr_12_bF_buf2), .Y(u2_u2__abc_47660_n199) );
  INVX2 INVX2_44 ( .A(rst_i_bF_buf2), .Y(u2_u2__abc_47660_n305) );
  INVX2 INVX2_45 ( .A(row_adr_0_bF_buf1), .Y(u2_u3__abc_47660_n139) );
  INVX2 INVX2_46 ( .A(row_adr_1_bF_buf1), .Y(u2_u3__abc_47660_n144) );
  INVX2 INVX2_47 ( .A(row_adr_2_bF_buf1), .Y(u2_u3__abc_47660_n149) );
  INVX2 INVX2_48 ( .A(row_adr_3_bF_buf1), .Y(u2_u3__abc_47660_n154) );
  INVX2 INVX2_49 ( .A(row_adr_4_bF_buf1), .Y(u2_u3__abc_47660_n159) );
  INVX2 INVX2_5 ( .A(row_adr_2_bF_buf4), .Y(u2_u0__abc_47660_n149) );
  INVX2 INVX2_50 ( .A(row_adr_5_bF_buf1), .Y(u2_u3__abc_47660_n164) );
  INVX2 INVX2_51 ( .A(row_adr_6_bF_buf1), .Y(u2_u3__abc_47660_n169) );
  INVX2 INVX2_52 ( .A(row_adr_7_bF_buf1), .Y(u2_u3__abc_47660_n174) );
  INVX2 INVX2_53 ( .A(row_adr_8_bF_buf1), .Y(u2_u3__abc_47660_n179) );
  INVX2 INVX2_54 ( .A(row_adr_9_bF_buf1), .Y(u2_u3__abc_47660_n184) );
  INVX2 INVX2_55 ( .A(row_adr_10_bF_buf1), .Y(u2_u3__abc_47660_n189) );
  INVX2 INVX2_56 ( .A(row_adr_11_bF_buf1), .Y(u2_u3__abc_47660_n194) );
  INVX2 INVX2_57 ( .A(row_adr_12_bF_buf1), .Y(u2_u3__abc_47660_n199) );
  INVX2 INVX2_58 ( .A(rst_i_bF_buf1), .Y(u2_u3__abc_47660_n305) );
  INVX2 INVX2_59 ( .A(row_adr_0_bF_buf0), .Y(u2_u4__abc_47660_n139) );
  INVX2 INVX2_6 ( .A(row_adr_3_bF_buf4), .Y(u2_u0__abc_47660_n154) );
  INVX2 INVX2_60 ( .A(row_adr_1_bF_buf0), .Y(u2_u4__abc_47660_n144) );
  INVX2 INVX2_61 ( .A(row_adr_2_bF_buf0), .Y(u2_u4__abc_47660_n149) );
  INVX2 INVX2_62 ( .A(row_adr_3_bF_buf0), .Y(u2_u4__abc_47660_n154) );
  INVX2 INVX2_63 ( .A(row_adr_4_bF_buf0), .Y(u2_u4__abc_47660_n159) );
  INVX2 INVX2_64 ( .A(row_adr_5_bF_buf0), .Y(u2_u4__abc_47660_n164) );
  INVX2 INVX2_65 ( .A(row_adr_6_bF_buf0), .Y(u2_u4__abc_47660_n169) );
  INVX2 INVX2_66 ( .A(row_adr_7_bF_buf0), .Y(u2_u4__abc_47660_n174) );
  INVX2 INVX2_67 ( .A(row_adr_8_bF_buf0), .Y(u2_u4__abc_47660_n179) );
  INVX2 INVX2_68 ( .A(row_adr_9_bF_buf0), .Y(u2_u4__abc_47660_n184) );
  INVX2 INVX2_69 ( .A(row_adr_10_bF_buf0), .Y(u2_u4__abc_47660_n189) );
  INVX2 INVX2_7 ( .A(row_adr_4_bF_buf4), .Y(u2_u0__abc_47660_n159) );
  INVX2 INVX2_70 ( .A(row_adr_11_bF_buf0), .Y(u2_u4__abc_47660_n194) );
  INVX2 INVX2_71 ( .A(row_adr_12_bF_buf0), .Y(u2_u4__abc_47660_n199) );
  INVX2 INVX2_72 ( .A(rst_i_bF_buf0), .Y(u2_u4__abc_47660_n305) );
  INVX2 INVX2_73 ( .A(row_adr_0_bF_buf6), .Y(u2_u5__abc_47660_n139) );
  INVX2 INVX2_74 ( .A(row_adr_1_bF_buf6), .Y(u2_u5__abc_47660_n144) );
  INVX2 INVX2_75 ( .A(row_adr_2_bF_buf6), .Y(u2_u5__abc_47660_n149) );
  INVX2 INVX2_76 ( .A(row_adr_3_bF_buf6), .Y(u2_u5__abc_47660_n154) );
  INVX2 INVX2_77 ( .A(row_adr_4_bF_buf6), .Y(u2_u5__abc_47660_n159) );
  INVX2 INVX2_78 ( .A(row_adr_5_bF_buf6), .Y(u2_u5__abc_47660_n164) );
  INVX2 INVX2_79 ( .A(row_adr_6_bF_buf6), .Y(u2_u5__abc_47660_n169) );
  INVX2 INVX2_8 ( .A(row_adr_5_bF_buf4), .Y(u2_u0__abc_47660_n164) );
  INVX2 INVX2_80 ( .A(row_adr_7_bF_buf6), .Y(u2_u5__abc_47660_n174) );
  INVX2 INVX2_81 ( .A(row_adr_8_bF_buf6), .Y(u2_u5__abc_47660_n179) );
  INVX2 INVX2_82 ( .A(row_adr_9_bF_buf6), .Y(u2_u5__abc_47660_n184) );
  INVX2 INVX2_83 ( .A(row_adr_10_bF_buf6), .Y(u2_u5__abc_47660_n189) );
  INVX2 INVX2_84 ( .A(row_adr_11_bF_buf6), .Y(u2_u5__abc_47660_n194) );
  INVX2 INVX2_85 ( .A(row_adr_12_bF_buf6), .Y(u2_u5__abc_47660_n199) );
  INVX2 INVX2_86 ( .A(rst_i_bF_buf3), .Y(u2_u5__abc_47660_n305) );
  INVX2 INVX2_87 ( .A(u3_rd_fifo_clr), .Y(u3_u0__abc_48231_n1002) );
  INVX2 INVX2_88 ( .A(rfr_ack), .Y(u4__abc_49152_n119) );
  INVX2 INVX2_89 ( .A(u5_state_6_), .Y(u5__abc_54027_n267) );
  INVX2 INVX2_9 ( .A(row_adr_6_bF_buf4), .Y(u2_u0__abc_47660_n169) );
  INVX2 INVX2_90 ( .A(u5_mc_le), .Y(u5_mc_le_FF_INPUT) );
  INVX2 INVX2_91 ( .A(u5__abc_54027_n420), .Y(u5__abc_54027_n421) );
  INVX2 INVX2_92 ( .A(u5__abc_54027_n425), .Y(u5__abc_54027_n426) );
  INVX2 INVX2_93 ( .A(u5__abc_54027_n435), .Y(u5__abc_54027_n436) );
  INVX2 INVX2_94 ( .A(u5__abc_54027_n291), .Y(u5__abc_54027_n444) );
  INVX2 INVX2_95 ( .A(u5_kro), .Y(u5__abc_54027_n519) );
  INVX2 INVX2_96 ( .A(u1_wr_cycle), .Y(u5__abc_54027_n533) );
  INVX2 INVX2_97 ( .A(u5__abc_54027_n582), .Y(u5__abc_54027_n583) );
  INVX2 INVX2_98 ( .A(u5__abc_54027_n595), .Y(u5__abc_54027_n596) );
  INVX2 INVX2_99 ( .A(u5__abc_54027_n424), .Y(u5__abc_54027_n614) );
  INVX4 INVX4_1 ( .A(_abc_55805_n237_1), .Y(_abc_55805_n245_1) );
  INVX4 INVX4_10 ( .A(rst_i_bF_buf1), .Y(u0_u5__abc_45296_n325) );
  INVX4 INVX4_11 ( .A(cs_le_bF_buf4), .Y(u1__abc_45852_n281) );
  INVX4 INVX4_12 ( .A(u1__abc_45852_n279_1), .Y(page_size_9_) );
  INVX4 INVX4_13 ( .A(u1_bas), .Y(u1__abc_45852_n290) );
  INVX4 INVX4_14 ( .A(u1__abc_45852_n519), .Y(u1__abc_45852_n520_1) );
  INVX4 INVX4_15 ( .A(row_sel), .Y(u1__abc_45852_n910) );
  INVX4 INVX4_16 ( .A(u1__abc_45852_n909), .Y(u1__abc_45852_n917) );
  INVX4 INVX4_17 ( .A(u2_u0__abc_47660_n205), .Y(u2_u0__abc_47660_n207) );
  INVX4 INVX4_18 ( .A(u2_u0__abc_47660_n248), .Y(u2_u0__abc_47660_n250) );
  INVX4 INVX4_19 ( .A(u2_u0__abc_47660_n290_1), .Y(u2_u0__abc_47660_n292_1) );
  INVX4 INVX4_2 ( .A(u0__abc_49347_n1952_1_bF_buf3), .Y(u0__abc_49347_n1953_1) );
  INVX4 INVX4_20 ( .A(u2_u1__abc_47660_n205), .Y(u2_u1__abc_47660_n207) );
  INVX4 INVX4_21 ( .A(u2_u1__abc_47660_n248), .Y(u2_u1__abc_47660_n250) );
  INVX4 INVX4_22 ( .A(u2_u1__abc_47660_n290_1), .Y(u2_u1__abc_47660_n292_1) );
  INVX4 INVX4_23 ( .A(u2_u2__abc_47660_n205), .Y(u2_u2__abc_47660_n207) );
  INVX4 INVX4_24 ( .A(u2_u2__abc_47660_n248), .Y(u2_u2__abc_47660_n250) );
  INVX4 INVX4_25 ( .A(u2_u2__abc_47660_n290_1), .Y(u2_u2__abc_47660_n292_1) );
  INVX4 INVX4_26 ( .A(u2_u3__abc_47660_n205), .Y(u2_u3__abc_47660_n207) );
  INVX4 INVX4_27 ( .A(u2_u3__abc_47660_n248), .Y(u2_u3__abc_47660_n250) );
  INVX4 INVX4_28 ( .A(u2_u3__abc_47660_n290_1), .Y(u2_u3__abc_47660_n292_1) );
  INVX4 INVX4_29 ( .A(u2_u4__abc_47660_n205), .Y(u2_u4__abc_47660_n207) );
  INVX4 INVX4_3 ( .A(cs_le_bF_buf2), .Y(u0__abc_49347_n4279) );
  INVX4 INVX4_30 ( .A(u2_u4__abc_47660_n248), .Y(u2_u4__abc_47660_n250) );
  INVX4 INVX4_31 ( .A(u2_u4__abc_47660_n290_1), .Y(u2_u4__abc_47660_n292_1) );
  INVX4 INVX4_32 ( .A(u2_u5__abc_47660_n205), .Y(u2_u5__abc_47660_n207) );
  INVX4 INVX4_33 ( .A(u2_u5__abc_47660_n248), .Y(u2_u5__abc_47660_n250) );
  INVX4 INVX4_34 ( .A(u2_u5__abc_47660_n290_1), .Y(u2_u5__abc_47660_n292_1) );
  INVX4 INVX4_35 ( .A(pack_le2), .Y(u3__abc_46775_n424) );
  INVX4 INVX4_36 ( .A(u3__abc_46775_n453), .Y(u3__abc_46775_n454) );
  INVX4 INVX4_37 ( .A(u3__abc_46775_n451), .Y(u3__abc_46775_n459) );
  INVX4 INVX4_38 ( .A(pack_le0), .Y(u3__abc_46775_n505) );
  INVX4 INVX4_39 ( .A(rst_i_bF_buf2), .Y(u3_u0__abc_48231_n514) );
  INVX4 INVX4_4 ( .A(u0__abc_49347_n4407), .Y(u0__abc_49347_n4409) );
  INVX4 INVX4_40 ( .A(u5__abc_54027_n369), .Y(u5__abc_54027_n370) );
  INVX4 INVX4_41 ( .A(u5_wb_wait), .Y(u5__abc_54027_n477) );
  INVX4 INVX4_42 ( .A(u5__abc_54027_n708), .Y(u5__abc_54027_n709_1) );
  INVX4 INVX4_43 ( .A(u5_cmd_asserted_bF_buf1), .Y(u5__abc_54027_n1312_1) );
  INVX4 INVX4_44 ( .A(u5_tmr_done), .Y(u5__abc_54027_n1383_1) );
  INVX4 INVX4_45 ( .A(rst_i_bF_buf2), .Y(u7__abc_47535_n99) );
  INVX4 INVX4_5 ( .A(rst_i_bF_buf2), .Y(u0_u0__abc_43300_n325) );
  INVX4 INVX4_6 ( .A(rst_i_bF_buf1), .Y(u0_u1__abc_43657_n324) );
  INVX4 INVX4_7 ( .A(rst_i_bF_buf0), .Y(u0_u2__abc_44109_n324) );
  INVX4 INVX4_8 ( .A(rst_i_bF_buf3), .Y(u0_u3__abc_44466_n328) );
  INVX4 INVX4_9 ( .A(rst_i_bF_buf2), .Y(u0_u4__abc_44844_n324) );
  INVX8 INVX8_1 ( .A(u0__abc_49347_n1175_bF_buf6), .Y(u0__abc_49347_n1176_1) );
  INVX8 INVX8_10 ( .A(u0_cs2_bF_buf5), .Y(u0__abc_49347_n2724) );
  INVX8 INVX8_11 ( .A(u0_cs3_bF_buf5), .Y(u0__abc_49347_n2725) );
  INVX8 INVX8_12 ( .A(u0_cs4_bF_buf5), .Y(u0__abc_49347_n2726) );
  INVX8 INVX8_13 ( .A(1'b0), .Y(u0__abc_49347_n2728) );
  INVX8 INVX8_14 ( .A(u0_cs5_bF_buf4), .Y(u0__abc_49347_n2730) );
  INVX8 INVX8_15 ( .A(u0_cs0_bF_buf4), .Y(u0__abc_49347_n2748) );
  INVX8 INVX8_16 ( .A(u0_rst_r3_bF_buf3), .Y(u0__abc_49347_n4304) );
  INVX8 INVX8_17 ( .A(u0__abc_49347_n4443_bF_buf3), .Y(u0__abc_49347_n4444) );
  INVX8 INVX8_18 ( .A(rst_i_bF_buf3), .Y(u0__abc_49347_n3188) );
  INVX8 INVX8_19 ( .A(u0_u0_rst_r2), .Y(u0_u0__abc_43300_n218) );
  INVX8 INVX8_2 ( .A(spec_req_cs_1_bF_buf3), .Y(u0__abc_49347_n1178_1) );
  INVX8 INVX8_20 ( .A(u0_u0_lmr_req_we_FF_INPUT_bF_buf3), .Y(u0_u0__abc_43300_n219_1) );
  INVX8 INVX8_21 ( .A(u0_u0_init_req_we_FF_INPUT_bF_buf3), .Y(u0_u0__abc_43300_n350) );
  INVX8 INVX8_22 ( .A(u0_u1_rst_r2), .Y(u0_u1__abc_43657_n219_1) );
  INVX8 INVX8_23 ( .A(u0_u2_rst_r2), .Y(u0_u2__abc_44109_n209) );
  INVX8 INVX8_24 ( .A(u0_u2_init_req_we_FF_INPUT_bF_buf3), .Y(u0_u2__abc_44109_n210_1) );
  INVX8 INVX8_25 ( .A(u0_u2_lmr_req_we_FF_INPUT_bF_buf3), .Y(u0_u2__abc_44109_n340) );
  INVX8 INVX8_26 ( .A(u0_u3_rst_r2_bF_buf5), .Y(u0_u3__abc_44466_n205_1) );
  INVX8 INVX8_27 ( .A(u0_u3_init_req_we_FF_INPUT_bF_buf4), .Y(u0_u3__abc_44466_n239_1) );
  INVX8 INVX8_28 ( .A(u0_u3_lmr_req_we_FF_INPUT_bF_buf4), .Y(u0_u3__abc_44466_n364) );
  INVX8 INVX8_29 ( .A(u0_u4_rst_r2), .Y(u0_u4__abc_44844_n209_1) );
  INVX8 INVX8_3 ( .A(spec_req_cs_2_bF_buf3), .Y(u0__abc_49347_n1179) );
  INVX8 INVX8_30 ( .A(u0_u5_rst_r2), .Y(u0_u5__abc_45296_n218) );
  INVX8 INVX8_31 ( .A(u1__abc_45852_n260_1), .Y(u1__abc_45852_n261) );
  INVX8 INVX8_32 ( .A(next_adr_bF_buf3), .Y(u1__abc_45852_n556) );
  INVX8 INVX8_33 ( .A(u1__abc_45852_n554_1_bF_buf3), .Y(u1__abc_45852_n562) );
  INVX8 INVX8_34 ( .A(wb_stb_i_bF_buf1), .Y(u1__abc_45852_n821) );
  INVX8 INVX8_35 ( .A(u1__abc_45852_n901_bF_buf3), .Y(u1__abc_45852_n903) );
  INVX8 INVX8_36 ( .A(u3__abc_46775_n277_1_bF_buf4), .Y(u3__abc_46775_n279) );
  INVX8 INVX8_37 ( .A(csc_5_bF_buf2), .Y(u3__abc_46775_n448) );
  INVX8 INVX8_38 ( .A(u3__abc_46775_n275_bF_buf3), .Y(u3__abc_46775_n625) );
  INVX8 INVX8_39 ( .A(rst_i_bF_buf1), .Y(u4__abc_49152_n191) );
  INVX8 INVX8_4 ( .A(spec_req_cs_3_bF_buf3), .Y(u0__abc_49347_n1180_1) );
  INVX8 INVX8_40 ( .A(rst_i_bF_buf0), .Y(u5__abc_54027_n1575) );
  INVX8 INVX8_41 ( .A(u6__abc_56056_n144_bF_buf3), .Y(u6__abc_56056_n154) );
  INVX8 INVX8_42 ( .A(rst_i_bF_buf3), .Y(u6__abc_56056_n167) );
  INVX8 INVX8_5 ( .A(spec_req_cs_4_bF_buf3), .Y(u0__abc_49347_n1181) );
  INVX8 INVX8_6 ( .A(spec_req_cs_6_bF_buf3), .Y(u0__abc_49347_n1183_1) );
  INVX8 INVX8_7 ( .A(spec_req_cs_5_bF_buf2), .Y(u0__abc_49347_n1185) );
  INVX8 INVX8_8 ( .A(spec_req_cs_0_bF_buf2), .Y(u0__abc_49347_n1203) );
  INVX8 INVX8_9 ( .A(u0_cs1_bF_buf5), .Y(u0__abc_49347_n2723) );
  OR2X2 OR2X2_1 ( .A(init_ack), .B(lmr_ack), .Y(lmr_sel) );
  OR2X2 OR2X2_10 ( .A(_abc_55805_n245_1), .B(cs_need_rfr_1_), .Y(_abc_55805_n252) );
  OR2X2 OR2X2_100 ( .A(lmr_sel_bF_buf1), .B(csc_5_bF_buf4), .Y(_abc_55805_n402) );
  OR2X2 OR2X2_1000 ( .A(u0__abc_49347_n4444_bF_buf0), .B(u0_csr_4_), .Y(u0__abc_49347_n4454) );
  OR2X2 OR2X2_1001 ( .A(u0__abc_49347_n4443_bF_buf3), .B(\wb_data_i[4] ), .Y(u0__abc_49347_n4455) );
  OR2X2 OR2X2_1002 ( .A(u0__abc_49347_n4444_bF_buf3), .B(u0_csr_5_), .Y(u0__abc_49347_n4457) );
  OR2X2 OR2X2_1003 ( .A(u0__abc_49347_n4443_bF_buf2), .B(\wb_data_i[5] ), .Y(u0__abc_49347_n4458) );
  OR2X2 OR2X2_1004 ( .A(u0__abc_49347_n4444_bF_buf2), .B(u0_csr_6_), .Y(u0__abc_49347_n4460) );
  OR2X2 OR2X2_1005 ( .A(u0__abc_49347_n4443_bF_buf1), .B(\wb_data_i[6] ), .Y(u0__abc_49347_n4461) );
  OR2X2 OR2X2_1006 ( .A(u0__abc_49347_n4444_bF_buf1), .B(u0_csr_7_), .Y(u0__abc_49347_n4463) );
  OR2X2 OR2X2_1007 ( .A(u0__abc_49347_n4443_bF_buf0), .B(\wb_data_i[7] ), .Y(u0__abc_49347_n4464) );
  OR2X2 OR2X2_1008 ( .A(u0__abc_49347_n4444_bF_buf0), .B(ref_int_0_), .Y(u0__abc_49347_n4466) );
  OR2X2 OR2X2_1009 ( .A(u0__abc_49347_n4443_bF_buf3), .B(\wb_data_i[8] ), .Y(u0__abc_49347_n4467) );
  OR2X2 OR2X2_101 ( .A(_abc_55805_n240_bF_buf0), .B(sp_csc_6_), .Y(_abc_55805_n404) );
  OR2X2 OR2X2_1010 ( .A(u0__abc_49347_n4444_bF_buf3), .B(ref_int_1_), .Y(u0__abc_49347_n4469) );
  OR2X2 OR2X2_1011 ( .A(u0__abc_49347_n4443_bF_buf2), .B(\wb_data_i[9] ), .Y(u0__abc_49347_n4470) );
  OR2X2 OR2X2_1012 ( .A(u0__abc_49347_n4444_bF_buf2), .B(ref_int_2_), .Y(u0__abc_49347_n4472) );
  OR2X2 OR2X2_1013 ( .A(u0__abc_49347_n4443_bF_buf1), .B(\wb_data_i[10] ), .Y(u0__abc_49347_n4473) );
  OR2X2 OR2X2_1014 ( .A(u0__abc_49347_n4444_bF_buf1), .B(rfr_ps_val_0_), .Y(u0__abc_49347_n4475) );
  OR2X2 OR2X2_1015 ( .A(u0__abc_49347_n4443_bF_buf0), .B(\wb_data_i[24] ), .Y(u0__abc_49347_n4476) );
  OR2X2 OR2X2_1016 ( .A(u0__abc_49347_n4444_bF_buf0), .B(rfr_ps_val_1_), .Y(u0__abc_49347_n4478) );
  OR2X2 OR2X2_1017 ( .A(u0__abc_49347_n4443_bF_buf3), .B(\wb_data_i[25] ), .Y(u0__abc_49347_n4479) );
  OR2X2 OR2X2_1018 ( .A(u0__abc_49347_n4444_bF_buf3), .B(rfr_ps_val_2_), .Y(u0__abc_49347_n4481) );
  OR2X2 OR2X2_1019 ( .A(u0__abc_49347_n4443_bF_buf2), .B(\wb_data_i[26] ), .Y(u0__abc_49347_n4482) );
  OR2X2 OR2X2_102 ( .A(lmr_sel_bF_buf0), .B(csc_6_), .Y(_abc_55805_n405) );
  OR2X2 OR2X2_1020 ( .A(u0__abc_49347_n4444_bF_buf2), .B(rfr_ps_val_3_), .Y(u0__abc_49347_n4484) );
  OR2X2 OR2X2_1021 ( .A(u0__abc_49347_n4443_bF_buf1), .B(\wb_data_i[27] ), .Y(u0__abc_49347_n4485) );
  OR2X2 OR2X2_1022 ( .A(u0__abc_49347_n4444_bF_buf1), .B(rfr_ps_val_4_), .Y(u0__abc_49347_n4487) );
  OR2X2 OR2X2_1023 ( .A(u0__abc_49347_n4443_bF_buf0), .B(\wb_data_i[28] ), .Y(u0__abc_49347_n4488) );
  OR2X2 OR2X2_1024 ( .A(u0__abc_49347_n4444_bF_buf0), .B(rfr_ps_val_5_), .Y(u0__abc_49347_n4490) );
  OR2X2 OR2X2_1025 ( .A(u0__abc_49347_n4443_bF_buf3), .B(\wb_data_i[29] ), .Y(u0__abc_49347_n4491) );
  OR2X2 OR2X2_1026 ( .A(u0__abc_49347_n4444_bF_buf3), .B(rfr_ps_val_6_), .Y(u0__abc_49347_n4493) );
  OR2X2 OR2X2_1027 ( .A(u0__abc_49347_n4443_bF_buf2), .B(\wb_data_i[30] ), .Y(u0__abc_49347_n4494) );
  OR2X2 OR2X2_1028 ( .A(u0__abc_49347_n4444_bF_buf2), .B(rfr_ps_val_7_), .Y(u0__abc_49347_n4496) );
  OR2X2 OR2X2_1029 ( .A(u0__abc_49347_n4443_bF_buf1), .B(\wb_data_i[31] ), .Y(u0__abc_49347_n4497) );
  OR2X2 OR2X2_103 ( .A(_abc_55805_n240_bF_buf5), .B(sp_csc_7_), .Y(_abc_55805_n407) );
  OR2X2 OR2X2_1030 ( .A(u0__abc_49347_n4520), .B(u0__abc_49347_n4517), .Y(u0__abc_49347_n4521) );
  OR2X2 OR2X2_1031 ( .A(u0__abc_49347_n4521), .B(u0__abc_49347_n4512), .Y(u0__abc_49347_n4522) );
  OR2X2 OR2X2_1032 ( .A(u0__abc_49347_n4522), .B(u0__abc_49347_n4508), .Y(u0__abc_49347_n4523) );
  OR2X2 OR2X2_1033 ( .A(u0__abc_49347_n4532), .B(u0__abc_49347_n4529), .Y(u0__abc_49347_n4533) );
  OR2X2 OR2X2_1034 ( .A(u0__abc_49347_n4533), .B(u0__abc_49347_n4527), .Y(u0__abc_49347_n4534) );
  OR2X2 OR2X2_1035 ( .A(u0__abc_49347_n4538), .B(u0__abc_49347_n4540), .Y(u0__abc_49347_n4541) );
  OR2X2 OR2X2_1036 ( .A(u0__abc_49347_n4541), .B(u0__abc_49347_n4536), .Y(u0__abc_49347_n4542) );
  OR2X2 OR2X2_1037 ( .A(u0__abc_49347_n4542), .B(u0__abc_49347_n4534), .Y(u0__abc_49347_n4543) );
  OR2X2 OR2X2_1038 ( .A(u0__abc_49347_n4543), .B(u0__abc_49347_n4523), .Y(u0__abc_49347_n4544) );
  OR2X2 OR2X2_1039 ( .A(u0__abc_49347_n4574), .B(u0__abc_49347_n4514), .Y(u0__abc_49347_n4575) );
  OR2X2 OR2X2_104 ( .A(lmr_sel_bF_buf6), .B(csc_7_), .Y(_abc_55805_n408) );
  OR2X2 OR2X2_1040 ( .A(u0__abc_49347_n4590), .B(u0__abc_49347_n4588), .Y(u0__abc_49347_n4591) );
  OR2X2 OR2X2_1041 ( .A(u0__abc_49347_n4591), .B(u0__abc_49347_n4587), .Y(u0__abc_49347_n4592) );
  OR2X2 OR2X2_1042 ( .A(u0__abc_49347_n4592), .B(u0__abc_49347_n4585), .Y(u0__abc_49347_n4593) );
  OR2X2 OR2X2_1043 ( .A(u0__abc_49347_n4595), .B(u0__abc_49347_n4594), .Y(u0__abc_49347_n4596) );
  OR2X2 OR2X2_1044 ( .A(u0__abc_49347_n4597), .B(u0__abc_49347_n4598), .Y(u0__abc_49347_n4599) );
  OR2X2 OR2X2_1045 ( .A(u0__abc_49347_n4596), .B(u0__abc_49347_n4599), .Y(u0__abc_49347_n4600) );
  OR2X2 OR2X2_1046 ( .A(u0__abc_49347_n4593), .B(u0__abc_49347_n4600), .Y(u0__abc_49347_n4601) );
  OR2X2 OR2X2_1047 ( .A(u0__abc_49347_n4583), .B(u0__abc_49347_n4601), .Y(u0__abc_49347_n4602) );
  OR2X2 OR2X2_1048 ( .A(u0__abc_49347_n4602), .B(u0__abc_49347_n4544), .Y(rf_dout_0_) );
  OR2X2 OR2X2_1049 ( .A(u0__abc_49347_n4605), .B(u0__abc_49347_n4606), .Y(u0__abc_49347_n4607) );
  OR2X2 OR2X2_105 ( .A(_abc_55805_n240_bF_buf4), .B(sp_csc_9_), .Y(_abc_55805_n413) );
  OR2X2 OR2X2_1050 ( .A(u0__abc_49347_n4607), .B(u0__abc_49347_n4604), .Y(u0__abc_49347_n4608) );
  OR2X2 OR2X2_1051 ( .A(u0__abc_49347_n4610), .B(u0__abc_49347_n4611), .Y(u0__abc_49347_n4612) );
  OR2X2 OR2X2_1052 ( .A(u0__abc_49347_n4612), .B(u0__abc_49347_n4609), .Y(u0__abc_49347_n4613) );
  OR2X2 OR2X2_1053 ( .A(u0__abc_49347_n4613), .B(u0__abc_49347_n4608), .Y(u0__abc_49347_n4614) );
  OR2X2 OR2X2_1054 ( .A(u0__abc_49347_n4616), .B(u0__abc_49347_n4617), .Y(u0__abc_49347_n4618) );
  OR2X2 OR2X2_1055 ( .A(u0__abc_49347_n4618), .B(u0__abc_49347_n4615), .Y(u0__abc_49347_n4619) );
  OR2X2 OR2X2_1056 ( .A(u0__abc_49347_n4614), .B(u0__abc_49347_n4619), .Y(u0__abc_49347_n4620) );
  OR2X2 OR2X2_1057 ( .A(u0__abc_49347_n4625), .B(u0__abc_49347_n4624), .Y(u0__abc_49347_n4626) );
  OR2X2 OR2X2_1058 ( .A(u0__abc_49347_n4626), .B(u0__abc_49347_n4623), .Y(u0__abc_49347_n4627) );
  OR2X2 OR2X2_1059 ( .A(u0__abc_49347_n4627), .B(u0__abc_49347_n4622), .Y(u0__abc_49347_n4628) );
  OR2X2 OR2X2_106 ( .A(lmr_sel_bF_buf5), .B(csc_9_), .Y(_abc_55805_n414) );
  OR2X2 OR2X2_1060 ( .A(u0__abc_49347_n4630), .B(u0__abc_49347_n4631), .Y(u0__abc_49347_n4632) );
  OR2X2 OR2X2_1061 ( .A(u0__abc_49347_n4632), .B(u0__abc_49347_n4629), .Y(u0__abc_49347_n4633) );
  OR2X2 OR2X2_1062 ( .A(u0__abc_49347_n4634), .B(u0__abc_49347_n4635), .Y(u0__abc_49347_n4636) );
  OR2X2 OR2X2_1063 ( .A(u0__abc_49347_n4633), .B(u0__abc_49347_n4636), .Y(u0__abc_49347_n4637) );
  OR2X2 OR2X2_1064 ( .A(u0__abc_49347_n4628), .B(u0__abc_49347_n4637), .Y(u0__abc_49347_n4638) );
  OR2X2 OR2X2_1065 ( .A(u0__abc_49347_n4621), .B(u0__abc_49347_n4638), .Y(u0__abc_49347_n4639) );
  OR2X2 OR2X2_1066 ( .A(u0__abc_49347_n4639), .B(u0__abc_49347_n4620), .Y(rf_dout_1_) );
  OR2X2 OR2X2_1067 ( .A(u0__abc_49347_n4644), .B(u0__abc_49347_n4643), .Y(u0__abc_49347_n4645) );
  OR2X2 OR2X2_1068 ( .A(u0__abc_49347_n4645), .B(u0__abc_49347_n4642), .Y(u0__abc_49347_n4646) );
  OR2X2 OR2X2_1069 ( .A(u0__abc_49347_n4646), .B(u0__abc_49347_n4641), .Y(u0__abc_49347_n4647) );
  OR2X2 OR2X2_107 ( .A(_abc_55805_n240_bF_buf3), .B(sp_csc_10_), .Y(_abc_55805_n416) );
  OR2X2 OR2X2_1070 ( .A(u0__abc_49347_n4650), .B(u0__abc_49347_n4649), .Y(u0__abc_49347_n4651) );
  OR2X2 OR2X2_1071 ( .A(u0__abc_49347_n4651), .B(u0__abc_49347_n4648), .Y(u0__abc_49347_n4652) );
  OR2X2 OR2X2_1072 ( .A(u0__abc_49347_n4654), .B(u0__abc_49347_n4655), .Y(u0__abc_49347_n4656) );
  OR2X2 OR2X2_1073 ( .A(u0__abc_49347_n4656), .B(u0__abc_49347_n4653), .Y(u0__abc_49347_n4657) );
  OR2X2 OR2X2_1074 ( .A(u0__abc_49347_n4657), .B(u0__abc_49347_n4652), .Y(u0__abc_49347_n4658) );
  OR2X2 OR2X2_1075 ( .A(u0__abc_49347_n4658), .B(u0__abc_49347_n4647), .Y(u0__abc_49347_n4659) );
  OR2X2 OR2X2_1076 ( .A(u0__abc_49347_n4664), .B(u0__abc_49347_n4663), .Y(u0__abc_49347_n4665) );
  OR2X2 OR2X2_1077 ( .A(u0__abc_49347_n4665), .B(u0__abc_49347_n4662), .Y(u0__abc_49347_n4666) );
  OR2X2 OR2X2_1078 ( .A(u0__abc_49347_n4666), .B(u0__abc_49347_n4661), .Y(u0__abc_49347_n4667) );
  OR2X2 OR2X2_1079 ( .A(u0__abc_49347_n4669), .B(u0__abc_49347_n4668), .Y(u0__abc_49347_n4670) );
  OR2X2 OR2X2_108 ( .A(lmr_sel_bF_buf4), .B(csc_10_), .Y(_abc_55805_n417) );
  OR2X2 OR2X2_1080 ( .A(u0__abc_49347_n4671), .B(u0__abc_49347_n4672), .Y(u0__abc_49347_n4673) );
  OR2X2 OR2X2_1081 ( .A(u0__abc_49347_n4670), .B(u0__abc_49347_n4673), .Y(u0__abc_49347_n4674) );
  OR2X2 OR2X2_1082 ( .A(u0__abc_49347_n4667), .B(u0__abc_49347_n4674), .Y(u0__abc_49347_n4675) );
  OR2X2 OR2X2_1083 ( .A(u0__abc_49347_n4660), .B(u0__abc_49347_n4675), .Y(u0__abc_49347_n4676) );
  OR2X2 OR2X2_1084 ( .A(u0__abc_49347_n4676), .B(u0__abc_49347_n4659), .Y(rf_dout_2_) );
  OR2X2 OR2X2_1085 ( .A(u0__abc_49347_n4681), .B(u0__abc_49347_n4680), .Y(u0__abc_49347_n4682) );
  OR2X2 OR2X2_1086 ( .A(u0__abc_49347_n4682), .B(u0__abc_49347_n4679), .Y(u0__abc_49347_n4683) );
  OR2X2 OR2X2_1087 ( .A(u0__abc_49347_n4683), .B(u0__abc_49347_n4678), .Y(u0__abc_49347_n4684) );
  OR2X2 OR2X2_1088 ( .A(u0__abc_49347_n4687), .B(u0__abc_49347_n4686), .Y(u0__abc_49347_n4688) );
  OR2X2 OR2X2_1089 ( .A(u0__abc_49347_n4688), .B(u0__abc_49347_n4685), .Y(u0__abc_49347_n4689) );
  OR2X2 OR2X2_109 ( .A(\wb_addr_i[31] ), .B(\wb_addr_i[30] ), .Y(_abc_55805_n482) );
  OR2X2 OR2X2_1090 ( .A(u0__abc_49347_n4691), .B(u0__abc_49347_n4692), .Y(u0__abc_49347_n4693) );
  OR2X2 OR2X2_1091 ( .A(u0__abc_49347_n4693), .B(u0__abc_49347_n4690), .Y(u0__abc_49347_n4694) );
  OR2X2 OR2X2_1092 ( .A(u0__abc_49347_n4694), .B(u0__abc_49347_n4689), .Y(u0__abc_49347_n4695) );
  OR2X2 OR2X2_1093 ( .A(u0__abc_49347_n4695), .B(u0__abc_49347_n4684), .Y(u0__abc_49347_n4696) );
  OR2X2 OR2X2_1094 ( .A(u0__abc_49347_n4701), .B(u0__abc_49347_n4700), .Y(u0__abc_49347_n4702) );
  OR2X2 OR2X2_1095 ( .A(u0__abc_49347_n4702), .B(u0__abc_49347_n4699), .Y(u0__abc_49347_n4703) );
  OR2X2 OR2X2_1096 ( .A(u0__abc_49347_n4703), .B(u0__abc_49347_n4698), .Y(u0__abc_49347_n4704) );
  OR2X2 OR2X2_1097 ( .A(u0__abc_49347_n4705), .B(u0__abc_49347_n4706), .Y(u0__abc_49347_n4707) );
  OR2X2 OR2X2_1098 ( .A(u0__abc_49347_n4708), .B(u0__abc_49347_n4709), .Y(u0__abc_49347_n4710) );
  OR2X2 OR2X2_1099 ( .A(u0__abc_49347_n4707), .B(u0__abc_49347_n4710), .Y(u0__abc_49347_n4711) );
  OR2X2 OR2X2_11 ( .A(_abc_55805_n240_bF_buf3), .B(spec_req_cs_2_bF_buf5), .Y(_abc_55805_n254) );
  OR2X2 OR2X2_110 ( .A(_abc_55805_n482), .B(\wb_addr_i[29] ), .Y(_abc_55805_n483) );
  OR2X2 OR2X2_1100 ( .A(u0__abc_49347_n4704), .B(u0__abc_49347_n4711), .Y(u0__abc_49347_n4712) );
  OR2X2 OR2X2_1101 ( .A(u0__abc_49347_n4697), .B(u0__abc_49347_n4712), .Y(u0__abc_49347_n4713) );
  OR2X2 OR2X2_1102 ( .A(u0__abc_49347_n4713), .B(u0__abc_49347_n4696), .Y(rf_dout_3_) );
  OR2X2 OR2X2_1103 ( .A(u0__abc_49347_n4716), .B(u0__abc_49347_n4717), .Y(u0__abc_49347_n4718) );
  OR2X2 OR2X2_1104 ( .A(u0__abc_49347_n4718), .B(u0__abc_49347_n4715), .Y(u0__abc_49347_n4719) );
  OR2X2 OR2X2_1105 ( .A(u0__abc_49347_n4721), .B(u0__abc_49347_n4722), .Y(u0__abc_49347_n4723) );
  OR2X2 OR2X2_1106 ( .A(u0__abc_49347_n4723), .B(u0__abc_49347_n4720), .Y(u0__abc_49347_n4724) );
  OR2X2 OR2X2_1107 ( .A(u0__abc_49347_n4724), .B(u0__abc_49347_n4719), .Y(u0__abc_49347_n4725) );
  OR2X2 OR2X2_1108 ( .A(u0__abc_49347_n4727), .B(u0__abc_49347_n4728), .Y(u0__abc_49347_n4729) );
  OR2X2 OR2X2_1109 ( .A(u0__abc_49347_n4729), .B(u0__abc_49347_n4726), .Y(u0__abc_49347_n4730) );
  OR2X2 OR2X2_111 ( .A(u0__abc_49347_n1101_1), .B(u0__abc_49347_n1102), .Y(u0__abc_49347_n1103_1) );
  OR2X2 OR2X2_1110 ( .A(u0__abc_49347_n4725), .B(u0__abc_49347_n4730), .Y(u0__abc_49347_n4731) );
  OR2X2 OR2X2_1111 ( .A(u0__abc_49347_n4736), .B(u0__abc_49347_n4735), .Y(u0__abc_49347_n4737) );
  OR2X2 OR2X2_1112 ( .A(u0__abc_49347_n4737), .B(u0__abc_49347_n4734), .Y(u0__abc_49347_n4738) );
  OR2X2 OR2X2_1113 ( .A(u0__abc_49347_n4738), .B(u0__abc_49347_n4733), .Y(u0__abc_49347_n4739) );
  OR2X2 OR2X2_1114 ( .A(u0__abc_49347_n4742), .B(u0__abc_49347_n4741), .Y(u0__abc_49347_n4743) );
  OR2X2 OR2X2_1115 ( .A(u0__abc_49347_n4743), .B(u0__abc_49347_n4740), .Y(u0__abc_49347_n4744) );
  OR2X2 OR2X2_1116 ( .A(u0__abc_49347_n4745), .B(u0__abc_49347_n4746), .Y(u0__abc_49347_n4747) );
  OR2X2 OR2X2_1117 ( .A(u0__abc_49347_n4744), .B(u0__abc_49347_n4747), .Y(u0__abc_49347_n4748) );
  OR2X2 OR2X2_1118 ( .A(u0__abc_49347_n4739), .B(u0__abc_49347_n4748), .Y(u0__abc_49347_n4749) );
  OR2X2 OR2X2_1119 ( .A(u0__abc_49347_n4732), .B(u0__abc_49347_n4749), .Y(u0__abc_49347_n4750) );
  OR2X2 OR2X2_112 ( .A(u0_sreq_cs_le), .B(spec_req_cs_0_bF_buf4), .Y(u0__abc_49347_n1107_1) );
  OR2X2 OR2X2_1120 ( .A(u0__abc_49347_n4750), .B(u0__abc_49347_n4731), .Y(rf_dout_4_) );
  OR2X2 OR2X2_1121 ( .A(u0__abc_49347_n4753), .B(u0__abc_49347_n4754), .Y(u0__abc_49347_n4755) );
  OR2X2 OR2X2_1122 ( .A(u0__abc_49347_n4755), .B(u0__abc_49347_n4752), .Y(u0__abc_49347_n4756) );
  OR2X2 OR2X2_1123 ( .A(u0__abc_49347_n4758), .B(u0__abc_49347_n4759), .Y(u0__abc_49347_n4760) );
  OR2X2 OR2X2_1124 ( .A(u0__abc_49347_n4760), .B(u0__abc_49347_n4757), .Y(u0__abc_49347_n4761) );
  OR2X2 OR2X2_1125 ( .A(u0__abc_49347_n4761), .B(u0__abc_49347_n4756), .Y(u0__abc_49347_n4762) );
  OR2X2 OR2X2_1126 ( .A(u0__abc_49347_n4764), .B(u0__abc_49347_n4765), .Y(u0__abc_49347_n4766) );
  OR2X2 OR2X2_1127 ( .A(u0__abc_49347_n4766), .B(u0__abc_49347_n4763), .Y(u0__abc_49347_n4767) );
  OR2X2 OR2X2_1128 ( .A(u0__abc_49347_n4762), .B(u0__abc_49347_n4767), .Y(u0__abc_49347_n4768) );
  OR2X2 OR2X2_1129 ( .A(u0__abc_49347_n4773), .B(u0__abc_49347_n4772), .Y(u0__abc_49347_n4774) );
  OR2X2 OR2X2_113 ( .A(u0__abc_49347_n1109_1), .B(u0__abc_49347_n1110), .Y(u0__abc_49347_n1111_1) );
  OR2X2 OR2X2_1130 ( .A(u0__abc_49347_n4774), .B(u0__abc_49347_n4771), .Y(u0__abc_49347_n4775) );
  OR2X2 OR2X2_1131 ( .A(u0__abc_49347_n4775), .B(u0__abc_49347_n4770), .Y(u0__abc_49347_n4776) );
  OR2X2 OR2X2_1132 ( .A(u0__abc_49347_n4778), .B(u0__abc_49347_n4779), .Y(u0__abc_49347_n4780) );
  OR2X2 OR2X2_1133 ( .A(u0__abc_49347_n4780), .B(u0__abc_49347_n4777), .Y(u0__abc_49347_n4781) );
  OR2X2 OR2X2_1134 ( .A(u0__abc_49347_n4782), .B(u0__abc_49347_n4783), .Y(u0__abc_49347_n4784) );
  OR2X2 OR2X2_1135 ( .A(u0__abc_49347_n4781), .B(u0__abc_49347_n4784), .Y(u0__abc_49347_n4785) );
  OR2X2 OR2X2_1136 ( .A(u0__abc_49347_n4776), .B(u0__abc_49347_n4785), .Y(u0__abc_49347_n4786) );
  OR2X2 OR2X2_1137 ( .A(u0__abc_49347_n4769), .B(u0__abc_49347_n4786), .Y(u0__abc_49347_n4787) );
  OR2X2 OR2X2_1138 ( .A(u0__abc_49347_n4787), .B(u0__abc_49347_n4768), .Y(rf_dout_5_) );
  OR2X2 OR2X2_1139 ( .A(u0__abc_49347_n4790), .B(u0__abc_49347_n4791), .Y(u0__abc_49347_n4792) );
  OR2X2 OR2X2_114 ( .A(u0__abc_49347_n1112), .B(u0__abc_49347_n1114), .Y(u0_spec_req_cs_1__FF_INPUT) );
  OR2X2 OR2X2_1140 ( .A(u0__abc_49347_n4792), .B(u0__abc_49347_n4789), .Y(u0__abc_49347_n4793) );
  OR2X2 OR2X2_1141 ( .A(u0__abc_49347_n4795), .B(u0__abc_49347_n4796), .Y(u0__abc_49347_n4797) );
  OR2X2 OR2X2_1142 ( .A(u0__abc_49347_n4797), .B(u0__abc_49347_n4794), .Y(u0__abc_49347_n4798) );
  OR2X2 OR2X2_1143 ( .A(u0__abc_49347_n4798), .B(u0__abc_49347_n4793), .Y(u0__abc_49347_n4799) );
  OR2X2 OR2X2_1144 ( .A(u0__abc_49347_n4801), .B(u0__abc_49347_n4802), .Y(u0__abc_49347_n4803) );
  OR2X2 OR2X2_1145 ( .A(u0__abc_49347_n4803), .B(u0__abc_49347_n4800), .Y(u0__abc_49347_n4804) );
  OR2X2 OR2X2_1146 ( .A(u0__abc_49347_n4799), .B(u0__abc_49347_n4804), .Y(u0__abc_49347_n4805) );
  OR2X2 OR2X2_1147 ( .A(u0__abc_49347_n4810), .B(u0__abc_49347_n4809), .Y(u0__abc_49347_n4811) );
  OR2X2 OR2X2_1148 ( .A(u0__abc_49347_n4811), .B(u0__abc_49347_n4808), .Y(u0__abc_49347_n4812) );
  OR2X2 OR2X2_1149 ( .A(u0__abc_49347_n4812), .B(u0__abc_49347_n4807), .Y(u0__abc_49347_n4813) );
  OR2X2 OR2X2_115 ( .A(u0__abc_49347_n1118_1), .B(u0__abc_49347_n1119), .Y(u0__abc_49347_n1120_1) );
  OR2X2 OR2X2_1150 ( .A(u0__abc_49347_n4816), .B(u0__abc_49347_n4815), .Y(u0__abc_49347_n4817) );
  OR2X2 OR2X2_1151 ( .A(u0__abc_49347_n4817), .B(u0__abc_49347_n4814), .Y(u0__abc_49347_n4818) );
  OR2X2 OR2X2_1152 ( .A(u0__abc_49347_n4820), .B(u0__abc_49347_n4819), .Y(u0__abc_49347_n4821) );
  OR2X2 OR2X2_1153 ( .A(u0__abc_49347_n4818), .B(u0__abc_49347_n4821), .Y(u0__abc_49347_n4822) );
  OR2X2 OR2X2_1154 ( .A(u0__abc_49347_n4813), .B(u0__abc_49347_n4822), .Y(u0__abc_49347_n4823) );
  OR2X2 OR2X2_1155 ( .A(u0__abc_49347_n4806), .B(u0__abc_49347_n4823), .Y(u0__abc_49347_n4824) );
  OR2X2 OR2X2_1156 ( .A(u0__abc_49347_n4824), .B(u0__abc_49347_n4805), .Y(rf_dout_6_) );
  OR2X2 OR2X2_1157 ( .A(u0__abc_49347_n4827), .B(u0__abc_49347_n4828), .Y(u0__abc_49347_n4829) );
  OR2X2 OR2X2_1158 ( .A(u0__abc_49347_n4829), .B(u0__abc_49347_n4826), .Y(u0__abc_49347_n4830) );
  OR2X2 OR2X2_1159 ( .A(u0__abc_49347_n4832), .B(u0__abc_49347_n4833), .Y(u0__abc_49347_n4834) );
  OR2X2 OR2X2_116 ( .A(u0__abc_49347_n1122_1), .B(u0__abc_49347_n1116_1), .Y(u0_spec_req_cs_2__FF_INPUT) );
  OR2X2 OR2X2_1160 ( .A(u0__abc_49347_n4834), .B(u0__abc_49347_n4831), .Y(u0__abc_49347_n4835) );
  OR2X2 OR2X2_1161 ( .A(u0__abc_49347_n4835), .B(u0__abc_49347_n4830), .Y(u0__abc_49347_n4836) );
  OR2X2 OR2X2_1162 ( .A(u0__abc_49347_n4838), .B(u0__abc_49347_n4839), .Y(u0__abc_49347_n4840) );
  OR2X2 OR2X2_1163 ( .A(u0__abc_49347_n4840), .B(u0__abc_49347_n4837), .Y(u0__abc_49347_n4841) );
  OR2X2 OR2X2_1164 ( .A(u0__abc_49347_n4836), .B(u0__abc_49347_n4841), .Y(u0__abc_49347_n4842) );
  OR2X2 OR2X2_1165 ( .A(u0__abc_49347_n4847), .B(u0__abc_49347_n4846), .Y(u0__abc_49347_n4848) );
  OR2X2 OR2X2_1166 ( .A(u0__abc_49347_n4848), .B(u0__abc_49347_n4845), .Y(u0__abc_49347_n4849) );
  OR2X2 OR2X2_1167 ( .A(u0__abc_49347_n4849), .B(u0__abc_49347_n4844), .Y(u0__abc_49347_n4850) );
  OR2X2 OR2X2_1168 ( .A(u0__abc_49347_n4852), .B(u0__abc_49347_n4853), .Y(u0__abc_49347_n4854) );
  OR2X2 OR2X2_1169 ( .A(u0__abc_49347_n4854), .B(u0__abc_49347_n4851), .Y(u0__abc_49347_n4855) );
  OR2X2 OR2X2_117 ( .A(u0__abc_49347_n1127), .B(u0__abc_49347_n1128_1), .Y(u0__abc_49347_n1129) );
  OR2X2 OR2X2_1170 ( .A(u0__abc_49347_n4857), .B(u0__abc_49347_n4856), .Y(u0__abc_49347_n4858) );
  OR2X2 OR2X2_1171 ( .A(u0__abc_49347_n4855), .B(u0__abc_49347_n4858), .Y(u0__abc_49347_n4859) );
  OR2X2 OR2X2_1172 ( .A(u0__abc_49347_n4850), .B(u0__abc_49347_n4859), .Y(u0__abc_49347_n4860) );
  OR2X2 OR2X2_1173 ( .A(u0__abc_49347_n4843), .B(u0__abc_49347_n4860), .Y(u0__abc_49347_n4861) );
  OR2X2 OR2X2_1174 ( .A(u0__abc_49347_n4861), .B(u0__abc_49347_n4842), .Y(rf_dout_7_) );
  OR2X2 OR2X2_1175 ( .A(u0__abc_49347_n4864), .B(u0__abc_49347_n4865), .Y(u0__abc_49347_n4866) );
  OR2X2 OR2X2_1176 ( .A(u0__abc_49347_n4866), .B(u0__abc_49347_n4863), .Y(u0__abc_49347_n4867) );
  OR2X2 OR2X2_1177 ( .A(u0__abc_49347_n4869), .B(u0__abc_49347_n4870), .Y(u0__abc_49347_n4871) );
  OR2X2 OR2X2_1178 ( .A(u0__abc_49347_n4871), .B(u0__abc_49347_n4868), .Y(u0__abc_49347_n4872) );
  OR2X2 OR2X2_1179 ( .A(u0__abc_49347_n4872), .B(u0__abc_49347_n4867), .Y(u0__abc_49347_n4873) );
  OR2X2 OR2X2_118 ( .A(u0__abc_49347_n1131), .B(u0__abc_49347_n1124_1), .Y(u0_spec_req_cs_3__FF_INPUT) );
  OR2X2 OR2X2_1180 ( .A(u0__abc_49347_n4875), .B(u0__abc_49347_n4876), .Y(u0__abc_49347_n4877) );
  OR2X2 OR2X2_1181 ( .A(u0__abc_49347_n4877), .B(u0__abc_49347_n4874), .Y(u0__abc_49347_n4878) );
  OR2X2 OR2X2_1182 ( .A(u0__abc_49347_n4873), .B(u0__abc_49347_n4878), .Y(u0__abc_49347_n4879) );
  OR2X2 OR2X2_1183 ( .A(u0__abc_49347_n4884), .B(u0__abc_49347_n4883), .Y(u0__abc_49347_n4885) );
  OR2X2 OR2X2_1184 ( .A(u0__abc_49347_n4885), .B(u0__abc_49347_n4882), .Y(u0__abc_49347_n4886) );
  OR2X2 OR2X2_1185 ( .A(u0__abc_49347_n4886), .B(u0__abc_49347_n4881), .Y(u0__abc_49347_n4887) );
  OR2X2 OR2X2_1186 ( .A(u0__abc_49347_n4889), .B(u0__abc_49347_n4890), .Y(u0__abc_49347_n4891) );
  OR2X2 OR2X2_1187 ( .A(u0__abc_49347_n4891), .B(u0__abc_49347_n4888), .Y(u0__abc_49347_n4892) );
  OR2X2 OR2X2_1188 ( .A(u0__abc_49347_n4893), .B(u0__abc_49347_n4894), .Y(u0__abc_49347_n4895) );
  OR2X2 OR2X2_1189 ( .A(u0__abc_49347_n4892), .B(u0__abc_49347_n4895), .Y(u0__abc_49347_n4896) );
  OR2X2 OR2X2_119 ( .A(u0__abc_49347_n1137_1), .B(u0__abc_49347_n1138), .Y(u0__abc_49347_n1139_1) );
  OR2X2 OR2X2_1190 ( .A(u0__abc_49347_n4887), .B(u0__abc_49347_n4896), .Y(u0__abc_49347_n4897) );
  OR2X2 OR2X2_1191 ( .A(u0__abc_49347_n4880), .B(u0__abc_49347_n4897), .Y(u0__abc_49347_n4898) );
  OR2X2 OR2X2_1192 ( .A(u0__abc_49347_n4898), .B(u0__abc_49347_n4879), .Y(rf_dout_8_) );
  OR2X2 OR2X2_1193 ( .A(u0__abc_49347_n4901), .B(u0__abc_49347_n4902), .Y(u0__abc_49347_n4903) );
  OR2X2 OR2X2_1194 ( .A(u0__abc_49347_n4903), .B(u0__abc_49347_n4900), .Y(u0__abc_49347_n4904) );
  OR2X2 OR2X2_1195 ( .A(u0__abc_49347_n4906), .B(u0__abc_49347_n4907), .Y(u0__abc_49347_n4908) );
  OR2X2 OR2X2_1196 ( .A(u0__abc_49347_n4908), .B(u0__abc_49347_n4905), .Y(u0__abc_49347_n4909) );
  OR2X2 OR2X2_1197 ( .A(u0__abc_49347_n4909), .B(u0__abc_49347_n4904), .Y(u0__abc_49347_n4910) );
  OR2X2 OR2X2_1198 ( .A(u0__abc_49347_n4913), .B(u0__abc_49347_n4912), .Y(u0__abc_49347_n4914) );
  OR2X2 OR2X2_1199 ( .A(u0__abc_49347_n4914), .B(u0__abc_49347_n4911), .Y(u0__abc_49347_n4915) );
  OR2X2 OR2X2_12 ( .A(lmr_sel_bF_buf4), .B(cs_2_), .Y(_abc_55805_n255) );
  OR2X2 OR2X2_120 ( .A(u0__abc_49347_n1141_1), .B(u0__abc_49347_n1133_1), .Y(u0_spec_req_cs_4__FF_INPUT) );
  OR2X2 OR2X2_1200 ( .A(u0__abc_49347_n4910), .B(u0__abc_49347_n4915), .Y(u0__abc_49347_n4916) );
  OR2X2 OR2X2_1201 ( .A(u0__abc_49347_n4921), .B(u0__abc_49347_n4920), .Y(u0__abc_49347_n4922) );
  OR2X2 OR2X2_1202 ( .A(u0__abc_49347_n4922), .B(u0__abc_49347_n4919), .Y(u0__abc_49347_n4923) );
  OR2X2 OR2X2_1203 ( .A(u0__abc_49347_n4923), .B(u0__abc_49347_n4918), .Y(u0__abc_49347_n4924) );
  OR2X2 OR2X2_1204 ( .A(u0__abc_49347_n4927), .B(u0__abc_49347_n4926), .Y(u0__abc_49347_n4928) );
  OR2X2 OR2X2_1205 ( .A(u0__abc_49347_n4928), .B(u0__abc_49347_n4925), .Y(u0__abc_49347_n4929) );
  OR2X2 OR2X2_1206 ( .A(u0__abc_49347_n4930), .B(u0__abc_49347_n4931), .Y(u0__abc_49347_n4932) );
  OR2X2 OR2X2_1207 ( .A(u0__abc_49347_n4929), .B(u0__abc_49347_n4932), .Y(u0__abc_49347_n4933) );
  OR2X2 OR2X2_1208 ( .A(u0__abc_49347_n4924), .B(u0__abc_49347_n4933), .Y(u0__abc_49347_n4934) );
  OR2X2 OR2X2_1209 ( .A(u0__abc_49347_n4917), .B(u0__abc_49347_n4934), .Y(u0__abc_49347_n4935) );
  OR2X2 OR2X2_121 ( .A(u0__abc_49347_n1144), .B(u0__abc_49347_n1145_1), .Y(u0__abc_49347_n1146) );
  OR2X2 OR2X2_1210 ( .A(u0__abc_49347_n4935), .B(u0__abc_49347_n4916), .Y(rf_dout_9_) );
  OR2X2 OR2X2_1211 ( .A(u0__abc_49347_n4940), .B(u0__abc_49347_n4939), .Y(u0__abc_49347_n4941) );
  OR2X2 OR2X2_1212 ( .A(u0__abc_49347_n4941), .B(u0__abc_49347_n4938), .Y(u0__abc_49347_n4942) );
  OR2X2 OR2X2_1213 ( .A(u0__abc_49347_n4942), .B(u0__abc_49347_n4937), .Y(u0__abc_49347_n4943) );
  OR2X2 OR2X2_1214 ( .A(u0__abc_49347_n4946), .B(u0__abc_49347_n4945), .Y(u0__abc_49347_n4947) );
  OR2X2 OR2X2_1215 ( .A(u0__abc_49347_n4947), .B(u0__abc_49347_n4944), .Y(u0__abc_49347_n4948) );
  OR2X2 OR2X2_1216 ( .A(u0__abc_49347_n4950), .B(u0__abc_49347_n4951), .Y(u0__abc_49347_n4952) );
  OR2X2 OR2X2_1217 ( .A(u0__abc_49347_n4952), .B(u0__abc_49347_n4949), .Y(u0__abc_49347_n4953) );
  OR2X2 OR2X2_1218 ( .A(u0__abc_49347_n4953), .B(u0__abc_49347_n4948), .Y(u0__abc_49347_n4954) );
  OR2X2 OR2X2_1219 ( .A(u0__abc_49347_n4954), .B(u0__abc_49347_n4943), .Y(u0__abc_49347_n4955) );
  OR2X2 OR2X2_122 ( .A(u0__abc_49347_n1151_1), .B(u0__abc_49347_n1143_1), .Y(u0_spec_req_cs_5__FF_INPUT) );
  OR2X2 OR2X2_1220 ( .A(u0__abc_49347_n4960), .B(u0__abc_49347_n4959), .Y(u0__abc_49347_n4961) );
  OR2X2 OR2X2_1221 ( .A(u0__abc_49347_n4961), .B(u0__abc_49347_n4958), .Y(u0__abc_49347_n4962) );
  OR2X2 OR2X2_1222 ( .A(u0__abc_49347_n4962), .B(u0__abc_49347_n4957), .Y(u0__abc_49347_n4963) );
  OR2X2 OR2X2_1223 ( .A(u0__abc_49347_n4965), .B(u0__abc_49347_n4964), .Y(u0__abc_49347_n4966) );
  OR2X2 OR2X2_1224 ( .A(u0__abc_49347_n4967), .B(u0__abc_49347_n4968), .Y(u0__abc_49347_n4969) );
  OR2X2 OR2X2_1225 ( .A(u0__abc_49347_n4966), .B(u0__abc_49347_n4969), .Y(u0__abc_49347_n4970) );
  OR2X2 OR2X2_1226 ( .A(u0__abc_49347_n4963), .B(u0__abc_49347_n4970), .Y(u0__abc_49347_n4971) );
  OR2X2 OR2X2_1227 ( .A(u0__abc_49347_n4956), .B(u0__abc_49347_n4971), .Y(u0__abc_49347_n4972) );
  OR2X2 OR2X2_1228 ( .A(u0__abc_49347_n4972), .B(u0__abc_49347_n4955), .Y(rf_dout_10_) );
  OR2X2 OR2X2_1229 ( .A(u0__abc_49347_n4975), .B(u0__abc_49347_n4976), .Y(u0__abc_49347_n4977) );
  OR2X2 OR2X2_123 ( .A(u0__abc_49347_n1155), .B(u0__abc_49347_n1156_1), .Y(u0__abc_49347_n1157) );
  OR2X2 OR2X2_1230 ( .A(u0__abc_49347_n4978), .B(u0__abc_49347_n4979), .Y(u0__abc_49347_n4980) );
  OR2X2 OR2X2_1231 ( .A(u0__abc_49347_n4977), .B(u0__abc_49347_n4980), .Y(u0__abc_49347_n4981) );
  OR2X2 OR2X2_1232 ( .A(u0__abc_49347_n4982), .B(u0__abc_49347_n4983), .Y(u0__abc_49347_n4984) );
  OR2X2 OR2X2_1233 ( .A(u0__abc_49347_n4986), .B(u0__abc_49347_n4985), .Y(u0__abc_49347_n4987) );
  OR2X2 OR2X2_1234 ( .A(u0__abc_49347_n4984), .B(u0__abc_49347_n4987), .Y(u0__abc_49347_n4988) );
  OR2X2 OR2X2_1235 ( .A(u0__abc_49347_n4988), .B(u0__abc_49347_n4981), .Y(u0__abc_49347_n4989) );
  OR2X2 OR2X2_1236 ( .A(u0__abc_49347_n4990), .B(u0__abc_49347_n4991), .Y(u0__abc_49347_n4992) );
  OR2X2 OR2X2_1237 ( .A(u0__abc_49347_n4994), .B(u0__abc_49347_n4993), .Y(u0__abc_49347_n4995) );
  OR2X2 OR2X2_1238 ( .A(u0__abc_49347_n4992), .B(u0__abc_49347_n4995), .Y(u0__abc_49347_n4996) );
  OR2X2 OR2X2_1239 ( .A(u0__abc_49347_n4998), .B(u0__abc_49347_n4997), .Y(u0__abc_49347_n4999) );
  OR2X2 OR2X2_124 ( .A(u0__abc_49347_n1160_1), .B(u0__abc_49347_n1161), .Y(u0_spec_req_cs_6__FF_INPUT) );
  OR2X2 OR2X2_1240 ( .A(u0__abc_49347_n5000), .B(u0__abc_49347_n5001), .Y(u0__abc_49347_n5002) );
  OR2X2 OR2X2_1241 ( .A(u0__abc_49347_n5002), .B(u0__abc_49347_n4999), .Y(u0__abc_49347_n5003) );
  OR2X2 OR2X2_1242 ( .A(u0__abc_49347_n4996), .B(u0__abc_49347_n5003), .Y(u0__abc_49347_n5004) );
  OR2X2 OR2X2_1243 ( .A(u0__abc_49347_n5004), .B(u0__abc_49347_n4989), .Y(u0__abc_49347_n5005) );
  OR2X2 OR2X2_1244 ( .A(u0__abc_49347_n5005), .B(u0__abc_49347_n4974), .Y(rf_dout_11_) );
  OR2X2 OR2X2_1245 ( .A(u0__abc_49347_n5009), .B(u0__abc_49347_n5008), .Y(u0__abc_49347_n5010) );
  OR2X2 OR2X2_1246 ( .A(u0__abc_49347_n5011), .B(u0__abc_49347_n5012), .Y(u0__abc_49347_n5013) );
  OR2X2 OR2X2_1247 ( .A(u0__abc_49347_n5010), .B(u0__abc_49347_n5013), .Y(u0__abc_49347_n5014) );
  OR2X2 OR2X2_1248 ( .A(u0__abc_49347_n5015), .B(u0__abc_49347_n5016), .Y(u0__abc_49347_n5017) );
  OR2X2 OR2X2_1249 ( .A(u0__abc_49347_n5018), .B(u0__abc_49347_n5019), .Y(u0__abc_49347_n5020) );
  OR2X2 OR2X2_125 ( .A(u0__abc_49347_n1100_1), .B(1'b0), .Y(u0__abc_49347_n1165) );
  OR2X2 OR2X2_1250 ( .A(u0__abc_49347_n5020), .B(u0__abc_49347_n5017), .Y(u0__abc_49347_n5021) );
  OR2X2 OR2X2_1251 ( .A(u0__abc_49347_n5014), .B(u0__abc_49347_n5021), .Y(u0__abc_49347_n5022) );
  OR2X2 OR2X2_1252 ( .A(u0__abc_49347_n5023), .B(u0__abc_49347_n5024), .Y(u0__abc_49347_n5025) );
  OR2X2 OR2X2_1253 ( .A(u0__abc_49347_n5026), .B(u0__abc_49347_n5027), .Y(u0__abc_49347_n5028) );
  OR2X2 OR2X2_1254 ( .A(u0__abc_49347_n5028), .B(u0__abc_49347_n5025), .Y(u0__abc_49347_n5029) );
  OR2X2 OR2X2_1255 ( .A(u0__abc_49347_n5030), .B(u0__abc_49347_n5031), .Y(u0__abc_49347_n5032) );
  OR2X2 OR2X2_1256 ( .A(u0__abc_49347_n5033), .B(u0__abc_49347_n5034), .Y(u0__abc_49347_n5035) );
  OR2X2 OR2X2_1257 ( .A(u0__abc_49347_n5035), .B(u0__abc_49347_n5032), .Y(u0__abc_49347_n5036) );
  OR2X2 OR2X2_1258 ( .A(u0__abc_49347_n5029), .B(u0__abc_49347_n5036), .Y(u0__abc_49347_n5037) );
  OR2X2 OR2X2_1259 ( .A(u0__abc_49347_n5022), .B(u0__abc_49347_n5037), .Y(u0__abc_49347_n5038) );
  OR2X2 OR2X2_126 ( .A(init_req), .B(1'b0), .Y(u0__abc_49347_n1166_1) );
  OR2X2 OR2X2_1260 ( .A(u0__abc_49347_n5038), .B(u0__abc_49347_n5007), .Y(rf_dout_12_) );
  OR2X2 OR2X2_1261 ( .A(u0__abc_49347_n5041), .B(u0__abc_49347_n5042), .Y(u0__abc_49347_n5043) );
  OR2X2 OR2X2_1262 ( .A(u0__abc_49347_n5045), .B(u0__abc_49347_n5044), .Y(u0__abc_49347_n5046) );
  OR2X2 OR2X2_1263 ( .A(u0__abc_49347_n5043), .B(u0__abc_49347_n5046), .Y(u0__abc_49347_n5047) );
  OR2X2 OR2X2_1264 ( .A(u0__abc_49347_n5048), .B(u0__abc_49347_n5049), .Y(u0__abc_49347_n5050) );
  OR2X2 OR2X2_1265 ( .A(u0__abc_49347_n5051), .B(u0__abc_49347_n5052), .Y(u0__abc_49347_n5053) );
  OR2X2 OR2X2_1266 ( .A(u0__abc_49347_n5050), .B(u0__abc_49347_n5053), .Y(u0__abc_49347_n5054) );
  OR2X2 OR2X2_1267 ( .A(u0__abc_49347_n5047), .B(u0__abc_49347_n5054), .Y(u0__abc_49347_n5055) );
  OR2X2 OR2X2_1268 ( .A(u0__abc_49347_n5056), .B(u0__abc_49347_n5057), .Y(u0__abc_49347_n5058) );
  OR2X2 OR2X2_1269 ( .A(u0__abc_49347_n5060), .B(u0__abc_49347_n5059), .Y(u0__abc_49347_n5061) );
  OR2X2 OR2X2_127 ( .A(u0__abc_49347_n1171), .B(u0__abc_49347_n1163), .Y(u0_spec_req_cs_7__FF_INPUT) );
  OR2X2 OR2X2_1270 ( .A(u0__abc_49347_n5058), .B(u0__abc_49347_n5061), .Y(u0__abc_49347_n5062) );
  OR2X2 OR2X2_1271 ( .A(u0__abc_49347_n5063), .B(u0__abc_49347_n5064), .Y(u0__abc_49347_n5065) );
  OR2X2 OR2X2_1272 ( .A(u0__abc_49347_n5066), .B(u0__abc_49347_n5067), .Y(u0__abc_49347_n5068) );
  OR2X2 OR2X2_1273 ( .A(u0__abc_49347_n5065), .B(u0__abc_49347_n5068), .Y(u0__abc_49347_n5069) );
  OR2X2 OR2X2_1274 ( .A(u0__abc_49347_n5069), .B(u0__abc_49347_n5062), .Y(u0__abc_49347_n5070) );
  OR2X2 OR2X2_1275 ( .A(u0__abc_49347_n5055), .B(u0__abc_49347_n5070), .Y(u0__abc_49347_n5071) );
  OR2X2 OR2X2_1276 ( .A(u0__abc_49347_n5071), .B(u0__abc_49347_n5040), .Y(rf_dout_13_) );
  OR2X2 OR2X2_1277 ( .A(u0__abc_49347_n5075), .B(u0__abc_49347_n5074), .Y(u0__abc_49347_n5076) );
  OR2X2 OR2X2_1278 ( .A(u0__abc_49347_n5077), .B(u0__abc_49347_n5078), .Y(u0__abc_49347_n5079) );
  OR2X2 OR2X2_1279 ( .A(u0__abc_49347_n5076), .B(u0__abc_49347_n5079), .Y(u0__abc_49347_n5080) );
  OR2X2 OR2X2_128 ( .A(cs_le_d), .B(u0_rf_we), .Y(u0__abc_49347_n1174_1) );
  OR2X2 OR2X2_1280 ( .A(u0__abc_49347_n5081), .B(u0__abc_49347_n5082), .Y(u0__abc_49347_n5083) );
  OR2X2 OR2X2_1281 ( .A(u0__abc_49347_n5084), .B(u0__abc_49347_n5085), .Y(u0__abc_49347_n5086) );
  OR2X2 OR2X2_1282 ( .A(u0__abc_49347_n5083), .B(u0__abc_49347_n5086), .Y(u0__abc_49347_n5087) );
  OR2X2 OR2X2_1283 ( .A(u0__abc_49347_n5087), .B(u0__abc_49347_n5080), .Y(u0__abc_49347_n5088) );
  OR2X2 OR2X2_1284 ( .A(u0__abc_49347_n5089), .B(u0__abc_49347_n5090), .Y(u0__abc_49347_n5091) );
  OR2X2 OR2X2_1285 ( .A(u0__abc_49347_n5092), .B(u0__abc_49347_n5093), .Y(u0__abc_49347_n5094) );
  OR2X2 OR2X2_1286 ( .A(u0__abc_49347_n5091), .B(u0__abc_49347_n5094), .Y(u0__abc_49347_n5095) );
  OR2X2 OR2X2_1287 ( .A(u0__abc_49347_n5096), .B(u0__abc_49347_n5097), .Y(u0__abc_49347_n5098) );
  OR2X2 OR2X2_1288 ( .A(u0__abc_49347_n5100), .B(u0__abc_49347_n5099), .Y(u0__abc_49347_n5101) );
  OR2X2 OR2X2_1289 ( .A(u0__abc_49347_n5098), .B(u0__abc_49347_n5101), .Y(u0__abc_49347_n5102) );
  OR2X2 OR2X2_129 ( .A(u0__abc_49347_n1183_1_bF_buf5), .B(1'b0), .Y(u0__abc_49347_n1184) );
  OR2X2 OR2X2_1290 ( .A(u0__abc_49347_n5102), .B(u0__abc_49347_n5095), .Y(u0__abc_49347_n5103) );
  OR2X2 OR2X2_1291 ( .A(u0__abc_49347_n5103), .B(u0__abc_49347_n5088), .Y(u0__abc_49347_n5104) );
  OR2X2 OR2X2_1292 ( .A(u0__abc_49347_n5104), .B(u0__abc_49347_n5073), .Y(rf_dout_14_) );
  OR2X2 OR2X2_1293 ( .A(u0__abc_49347_n5107), .B(u0__abc_49347_n5108), .Y(u0__abc_49347_n5109) );
  OR2X2 OR2X2_1294 ( .A(u0__abc_49347_n5111), .B(u0__abc_49347_n5110), .Y(u0__abc_49347_n5112) );
  OR2X2 OR2X2_1295 ( .A(u0__abc_49347_n5109), .B(u0__abc_49347_n5112), .Y(u0__abc_49347_n5113) );
  OR2X2 OR2X2_1296 ( .A(u0__abc_49347_n5114), .B(u0__abc_49347_n5115), .Y(u0__abc_49347_n5116) );
  OR2X2 OR2X2_1297 ( .A(u0__abc_49347_n5117), .B(u0__abc_49347_n5118), .Y(u0__abc_49347_n5119) );
  OR2X2 OR2X2_1298 ( .A(u0__abc_49347_n5116), .B(u0__abc_49347_n5119), .Y(u0__abc_49347_n5120) );
  OR2X2 OR2X2_1299 ( .A(u0__abc_49347_n5113), .B(u0__abc_49347_n5120), .Y(u0__abc_49347_n5121) );
  OR2X2 OR2X2_13 ( .A(_abc_55805_n256), .B(_abc_55805_n237_1), .Y(_abc_55805_n257) );
  OR2X2 OR2X2_130 ( .A(spec_req_cs_6_bF_buf2), .B(1'b0), .Y(u0__abc_49347_n1186) );
  OR2X2 OR2X2_1300 ( .A(u0__abc_49347_n5122), .B(u0__abc_49347_n5123), .Y(u0__abc_49347_n5124) );
  OR2X2 OR2X2_1301 ( .A(u0__abc_49347_n5126), .B(u0__abc_49347_n5125), .Y(u0__abc_49347_n5127) );
  OR2X2 OR2X2_1302 ( .A(u0__abc_49347_n5124), .B(u0__abc_49347_n5127), .Y(u0__abc_49347_n5128) );
  OR2X2 OR2X2_1303 ( .A(u0__abc_49347_n5129), .B(u0__abc_49347_n5130), .Y(u0__abc_49347_n5131) );
  OR2X2 OR2X2_1304 ( .A(u0__abc_49347_n5132), .B(u0__abc_49347_n5133), .Y(u0__abc_49347_n5134) );
  OR2X2 OR2X2_1305 ( .A(u0__abc_49347_n5131), .B(u0__abc_49347_n5134), .Y(u0__abc_49347_n5135) );
  OR2X2 OR2X2_1306 ( .A(u0__abc_49347_n5135), .B(u0__abc_49347_n5128), .Y(u0__abc_49347_n5136) );
  OR2X2 OR2X2_1307 ( .A(u0__abc_49347_n5121), .B(u0__abc_49347_n5136), .Y(u0__abc_49347_n5137) );
  OR2X2 OR2X2_1308 ( .A(u0__abc_49347_n5137), .B(u0__abc_49347_n5106), .Y(rf_dout_15_) );
  OR2X2 OR2X2_1309 ( .A(u0__abc_49347_n5141), .B(u0__abc_49347_n5140), .Y(u0__abc_49347_n5142) );
  OR2X2 OR2X2_131 ( .A(u0__abc_49347_n1188), .B(u0__abc_49347_n1182_1), .Y(u0__abc_49347_n1189) );
  OR2X2 OR2X2_1310 ( .A(u0__abc_49347_n5143), .B(u0__abc_49347_n5144), .Y(u0__abc_49347_n5145) );
  OR2X2 OR2X2_1311 ( .A(u0__abc_49347_n5142), .B(u0__abc_49347_n5145), .Y(u0__abc_49347_n5146) );
  OR2X2 OR2X2_1312 ( .A(u0__abc_49347_n5147), .B(u0__abc_49347_n5148), .Y(u0__abc_49347_n5149) );
  OR2X2 OR2X2_1313 ( .A(u0__abc_49347_n5150), .B(u0__abc_49347_n5151), .Y(u0__abc_49347_n5152) );
  OR2X2 OR2X2_1314 ( .A(u0__abc_49347_n5152), .B(u0__abc_49347_n5149), .Y(u0__abc_49347_n5153) );
  OR2X2 OR2X2_1315 ( .A(u0__abc_49347_n5146), .B(u0__abc_49347_n5153), .Y(u0__abc_49347_n5154) );
  OR2X2 OR2X2_1316 ( .A(u0__abc_49347_n5156), .B(u0__abc_49347_n5155), .Y(u0__abc_49347_n5157) );
  OR2X2 OR2X2_1317 ( .A(u0__abc_49347_n5158), .B(u0__abc_49347_n5159), .Y(u0__abc_49347_n5160) );
  OR2X2 OR2X2_1318 ( .A(u0__abc_49347_n5157), .B(u0__abc_49347_n5160), .Y(u0__abc_49347_n5161) );
  OR2X2 OR2X2_1319 ( .A(u0__abc_49347_n5162), .B(u0__abc_49347_n5163), .Y(u0__abc_49347_n5164) );
  OR2X2 OR2X2_132 ( .A(u0__abc_49347_n1190), .B(u0__abc_49347_n1191_1), .Y(u0__abc_49347_n1192_1) );
  OR2X2 OR2X2_1320 ( .A(u0__abc_49347_n5165), .B(u0__abc_49347_n5166), .Y(u0__abc_49347_n5167) );
  OR2X2 OR2X2_1321 ( .A(u0__abc_49347_n5164), .B(u0__abc_49347_n5167), .Y(u0__abc_49347_n5168) );
  OR2X2 OR2X2_1322 ( .A(u0__abc_49347_n5168), .B(u0__abc_49347_n5161), .Y(u0__abc_49347_n5169) );
  OR2X2 OR2X2_1323 ( .A(u0__abc_49347_n5154), .B(u0__abc_49347_n5169), .Y(u0__abc_49347_n5170) );
  OR2X2 OR2X2_1324 ( .A(u0__abc_49347_n5170), .B(u0__abc_49347_n5139), .Y(rf_dout_16_) );
  OR2X2 OR2X2_1325 ( .A(u0__abc_49347_n5174), .B(u0__abc_49347_n5173), .Y(u0__abc_49347_n5175) );
  OR2X2 OR2X2_1326 ( .A(u0__abc_49347_n5176), .B(u0__abc_49347_n5177), .Y(u0__abc_49347_n5178) );
  OR2X2 OR2X2_1327 ( .A(u0__abc_49347_n5178), .B(u0__abc_49347_n5175), .Y(u0__abc_49347_n5179) );
  OR2X2 OR2X2_1328 ( .A(u0__abc_49347_n5180), .B(u0__abc_49347_n5181), .Y(u0__abc_49347_n5182) );
  OR2X2 OR2X2_1329 ( .A(u0__abc_49347_n5183), .B(u0__abc_49347_n5184), .Y(u0__abc_49347_n5185) );
  OR2X2 OR2X2_133 ( .A(u0__abc_49347_n1193), .B(u0__abc_49347_n1194), .Y(u0__abc_49347_n1195) );
  OR2X2 OR2X2_1330 ( .A(u0__abc_49347_n5185), .B(u0__abc_49347_n5182), .Y(u0__abc_49347_n5186) );
  OR2X2 OR2X2_1331 ( .A(u0__abc_49347_n5179), .B(u0__abc_49347_n5186), .Y(u0__abc_49347_n5187) );
  OR2X2 OR2X2_1332 ( .A(u0__abc_49347_n5189), .B(u0__abc_49347_n5188), .Y(u0__abc_49347_n5190) );
  OR2X2 OR2X2_1333 ( .A(u0__abc_49347_n5191), .B(u0__abc_49347_n5192), .Y(u0__abc_49347_n5193) );
  OR2X2 OR2X2_1334 ( .A(u0__abc_49347_n5193), .B(u0__abc_49347_n5190), .Y(u0__abc_49347_n5194) );
  OR2X2 OR2X2_1335 ( .A(u0__abc_49347_n5195), .B(u0__abc_49347_n5196), .Y(u0__abc_49347_n5197) );
  OR2X2 OR2X2_1336 ( .A(u0__abc_49347_n5199), .B(u0__abc_49347_n5198), .Y(u0__abc_49347_n5200) );
  OR2X2 OR2X2_1337 ( .A(u0__abc_49347_n5197), .B(u0__abc_49347_n5200), .Y(u0__abc_49347_n5201) );
  OR2X2 OR2X2_1338 ( .A(u0__abc_49347_n5201), .B(u0__abc_49347_n5194), .Y(u0__abc_49347_n5202) );
  OR2X2 OR2X2_1339 ( .A(u0__abc_49347_n5187), .B(u0__abc_49347_n5202), .Y(u0__abc_49347_n5203) );
  OR2X2 OR2X2_134 ( .A(u0__abc_49347_n1196), .B(u0__abc_49347_n1197), .Y(u0__abc_49347_n1198) );
  OR2X2 OR2X2_1340 ( .A(u0__abc_49347_n5203), .B(u0__abc_49347_n5172), .Y(rf_dout_17_) );
  OR2X2 OR2X2_1341 ( .A(u0__abc_49347_n5206), .B(u0__abc_49347_n5207), .Y(u0__abc_49347_n5208) );
  OR2X2 OR2X2_1342 ( .A(u0__abc_49347_n5210), .B(u0__abc_49347_n5209), .Y(u0__abc_49347_n5211) );
  OR2X2 OR2X2_1343 ( .A(u0__abc_49347_n5208), .B(u0__abc_49347_n5211), .Y(u0__abc_49347_n5212) );
  OR2X2 OR2X2_1344 ( .A(u0__abc_49347_n5213), .B(u0__abc_49347_n5214), .Y(u0__abc_49347_n5215) );
  OR2X2 OR2X2_1345 ( .A(u0__abc_49347_n5216), .B(u0__abc_49347_n5217), .Y(u0__abc_49347_n5218) );
  OR2X2 OR2X2_1346 ( .A(u0__abc_49347_n5215), .B(u0__abc_49347_n5218), .Y(u0__abc_49347_n5219) );
  OR2X2 OR2X2_1347 ( .A(u0__abc_49347_n5219), .B(u0__abc_49347_n5212), .Y(u0__abc_49347_n5220) );
  OR2X2 OR2X2_1348 ( .A(u0__abc_49347_n5221), .B(u0__abc_49347_n5222), .Y(u0__abc_49347_n5223) );
  OR2X2 OR2X2_1349 ( .A(u0__abc_49347_n5224), .B(u0__abc_49347_n5225), .Y(u0__abc_49347_n5226) );
  OR2X2 OR2X2_135 ( .A(u0__abc_49347_n1200_1), .B(spec_req_cs_0_bF_buf3), .Y(u0__abc_49347_n1201_1) );
  OR2X2 OR2X2_1350 ( .A(u0__abc_49347_n5226), .B(u0__abc_49347_n5223), .Y(u0__abc_49347_n5227) );
  OR2X2 OR2X2_1351 ( .A(u0__abc_49347_n5228), .B(u0__abc_49347_n5229), .Y(u0__abc_49347_n5230) );
  OR2X2 OR2X2_1352 ( .A(u0__abc_49347_n5231), .B(u0__abc_49347_n5232), .Y(u0__abc_49347_n5233) );
  OR2X2 OR2X2_1353 ( .A(u0__abc_49347_n5233), .B(u0__abc_49347_n5230), .Y(u0__abc_49347_n5234) );
  OR2X2 OR2X2_1354 ( .A(u0__abc_49347_n5227), .B(u0__abc_49347_n5234), .Y(u0__abc_49347_n5235) );
  OR2X2 OR2X2_1355 ( .A(u0__abc_49347_n5235), .B(u0__abc_49347_n5220), .Y(u0__abc_49347_n5236) );
  OR2X2 OR2X2_1356 ( .A(u0__abc_49347_n5236), .B(u0__abc_49347_n5205), .Y(rf_dout_18_) );
  OR2X2 OR2X2_1357 ( .A(u0__abc_49347_n5239), .B(u0__abc_49347_n5240), .Y(u0__abc_49347_n5241) );
  OR2X2 OR2X2_1358 ( .A(u0__abc_49347_n5242), .B(u0__abc_49347_n5243), .Y(u0__abc_49347_n5244) );
  OR2X2 OR2X2_1359 ( .A(u0__abc_49347_n5244), .B(u0__abc_49347_n5241), .Y(u0__abc_49347_n5245) );
  OR2X2 OR2X2_136 ( .A(u0__abc_49347_n1199), .B(u0__abc_49347_n1201_1), .Y(u0__abc_49347_n1202) );
  OR2X2 OR2X2_1360 ( .A(u0__abc_49347_n5246), .B(u0__abc_49347_n5247), .Y(u0__abc_49347_n5248) );
  OR2X2 OR2X2_1361 ( .A(u0__abc_49347_n5250), .B(u0__abc_49347_n5249), .Y(u0__abc_49347_n5251) );
  OR2X2 OR2X2_1362 ( .A(u0__abc_49347_n5248), .B(u0__abc_49347_n5251), .Y(u0__abc_49347_n5252) );
  OR2X2 OR2X2_1363 ( .A(u0__abc_49347_n5252), .B(u0__abc_49347_n5245), .Y(u0__abc_49347_n5253) );
  OR2X2 OR2X2_1364 ( .A(u0__abc_49347_n5254), .B(u0__abc_49347_n5255), .Y(u0__abc_49347_n5256) );
  OR2X2 OR2X2_1365 ( .A(u0__abc_49347_n5258), .B(u0__abc_49347_n5257), .Y(u0__abc_49347_n5259) );
  OR2X2 OR2X2_1366 ( .A(u0__abc_49347_n5256), .B(u0__abc_49347_n5259), .Y(u0__abc_49347_n5260) );
  OR2X2 OR2X2_1367 ( .A(u0__abc_49347_n5261), .B(u0__abc_49347_n5262), .Y(u0__abc_49347_n5263) );
  OR2X2 OR2X2_1368 ( .A(u0__abc_49347_n5265), .B(u0__abc_49347_n5264), .Y(u0__abc_49347_n5266) );
  OR2X2 OR2X2_1369 ( .A(u0__abc_49347_n5263), .B(u0__abc_49347_n5266), .Y(u0__abc_49347_n5267) );
  OR2X2 OR2X2_137 ( .A(u0__abc_49347_n1203_bF_buf5), .B(u0_tms0_0_), .Y(u0__abc_49347_n1204) );
  OR2X2 OR2X2_1370 ( .A(u0__abc_49347_n5267), .B(u0__abc_49347_n5260), .Y(u0__abc_49347_n5268) );
  OR2X2 OR2X2_1371 ( .A(u0__abc_49347_n5253), .B(u0__abc_49347_n5268), .Y(u0__abc_49347_n5269) );
  OR2X2 OR2X2_1372 ( .A(u0__abc_49347_n5269), .B(u0__abc_49347_n5238), .Y(rf_dout_19_) );
  OR2X2 OR2X2_1373 ( .A(u0__abc_49347_n5273), .B(u0__abc_49347_n5272), .Y(u0__abc_49347_n5274) );
  OR2X2 OR2X2_1374 ( .A(u0__abc_49347_n5275), .B(u0__abc_49347_n5276), .Y(u0__abc_49347_n5277) );
  OR2X2 OR2X2_1375 ( .A(u0__abc_49347_n5274), .B(u0__abc_49347_n5277), .Y(u0__abc_49347_n5278) );
  OR2X2 OR2X2_1376 ( .A(u0__abc_49347_n5279), .B(u0__abc_49347_n5280), .Y(u0__abc_49347_n5281) );
  OR2X2 OR2X2_1377 ( .A(u0__abc_49347_n5282), .B(u0__abc_49347_n5283), .Y(u0__abc_49347_n5284) );
  OR2X2 OR2X2_1378 ( .A(u0__abc_49347_n5281), .B(u0__abc_49347_n5284), .Y(u0__abc_49347_n5285) );
  OR2X2 OR2X2_1379 ( .A(u0__abc_49347_n5278), .B(u0__abc_49347_n5285), .Y(u0__abc_49347_n5286) );
  OR2X2 OR2X2_138 ( .A(u0__abc_49347_n1206), .B(u0__abc_49347_n1177), .Y(u0_sp_tms_0__FF_INPUT) );
  OR2X2 OR2X2_1380 ( .A(u0__abc_49347_n5287), .B(u0__abc_49347_n5288), .Y(u0__abc_49347_n5289) );
  OR2X2 OR2X2_1381 ( .A(u0__abc_49347_n5290), .B(u0__abc_49347_n5291), .Y(u0__abc_49347_n5292) );
  OR2X2 OR2X2_1382 ( .A(u0__abc_49347_n5292), .B(u0__abc_49347_n5289), .Y(u0__abc_49347_n5293) );
  OR2X2 OR2X2_1383 ( .A(u0__abc_49347_n5295), .B(u0__abc_49347_n5294), .Y(u0__abc_49347_n5296) );
  OR2X2 OR2X2_1384 ( .A(u0__abc_49347_n5297), .B(u0__abc_49347_n5298), .Y(u0__abc_49347_n5299) );
  OR2X2 OR2X2_1385 ( .A(u0__abc_49347_n5299), .B(u0__abc_49347_n5296), .Y(u0__abc_49347_n5300) );
  OR2X2 OR2X2_1386 ( .A(u0__abc_49347_n5293), .B(u0__abc_49347_n5300), .Y(u0__abc_49347_n5301) );
  OR2X2 OR2X2_1387 ( .A(u0__abc_49347_n5286), .B(u0__abc_49347_n5301), .Y(u0__abc_49347_n5302) );
  OR2X2 OR2X2_1388 ( .A(u0__abc_49347_n5302), .B(u0__abc_49347_n5271), .Y(rf_dout_20_) );
  OR2X2 OR2X2_1389 ( .A(u0__abc_49347_n5305), .B(u0__abc_49347_n5306), .Y(u0__abc_49347_n5307) );
  OR2X2 OR2X2_139 ( .A(u0__abc_49347_n1183_1_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n1210_1) );
  OR2X2 OR2X2_1390 ( .A(u0__abc_49347_n5308), .B(u0__abc_49347_n5309), .Y(u0__abc_49347_n5310) );
  OR2X2 OR2X2_1391 ( .A(u0__abc_49347_n5307), .B(u0__abc_49347_n5310), .Y(u0__abc_49347_n5311) );
  OR2X2 OR2X2_1392 ( .A(u0__abc_49347_n5313), .B(u0__abc_49347_n5312), .Y(u0__abc_49347_n5314) );
  OR2X2 OR2X2_1393 ( .A(u0__abc_49347_n5315), .B(u0__abc_49347_n5316), .Y(u0__abc_49347_n5317) );
  OR2X2 OR2X2_1394 ( .A(u0__abc_49347_n5317), .B(u0__abc_49347_n5314), .Y(u0__abc_49347_n5318) );
  OR2X2 OR2X2_1395 ( .A(u0__abc_49347_n5311), .B(u0__abc_49347_n5318), .Y(u0__abc_49347_n5319) );
  OR2X2 OR2X2_1396 ( .A(u0__abc_49347_n5320), .B(u0__abc_49347_n5321), .Y(u0__abc_49347_n5322) );
  OR2X2 OR2X2_1397 ( .A(u0__abc_49347_n5323), .B(u0__abc_49347_n5324), .Y(u0__abc_49347_n5325) );
  OR2X2 OR2X2_1398 ( .A(u0__abc_49347_n5325), .B(u0__abc_49347_n5322), .Y(u0__abc_49347_n5326) );
  OR2X2 OR2X2_1399 ( .A(u0__abc_49347_n5328), .B(u0__abc_49347_n5327), .Y(u0__abc_49347_n5329) );
  OR2X2 OR2X2_14 ( .A(_abc_55805_n245_1), .B(cs_need_rfr_2_), .Y(_abc_55805_n258) );
  OR2X2 OR2X2_140 ( .A(spec_req_cs_6_bF_buf1), .B(1'b0), .Y(u0__abc_49347_n1211) );
  OR2X2 OR2X2_1400 ( .A(u0__abc_49347_n5330), .B(u0__abc_49347_n5331), .Y(u0__abc_49347_n5332) );
  OR2X2 OR2X2_1401 ( .A(u0__abc_49347_n5332), .B(u0__abc_49347_n5329), .Y(u0__abc_49347_n5333) );
  OR2X2 OR2X2_1402 ( .A(u0__abc_49347_n5326), .B(u0__abc_49347_n5333), .Y(u0__abc_49347_n5334) );
  OR2X2 OR2X2_1403 ( .A(u0__abc_49347_n5319), .B(u0__abc_49347_n5334), .Y(u0__abc_49347_n5335) );
  OR2X2 OR2X2_1404 ( .A(u0__abc_49347_n5335), .B(u0__abc_49347_n5304), .Y(rf_dout_21_) );
  OR2X2 OR2X2_1405 ( .A(u0__abc_49347_n5338), .B(u0__abc_49347_n5339), .Y(u0__abc_49347_n5340) );
  OR2X2 OR2X2_1406 ( .A(u0__abc_49347_n5342), .B(u0__abc_49347_n5341), .Y(u0__abc_49347_n5343) );
  OR2X2 OR2X2_1407 ( .A(u0__abc_49347_n5340), .B(u0__abc_49347_n5343), .Y(u0__abc_49347_n5344) );
  OR2X2 OR2X2_1408 ( .A(u0__abc_49347_n5346), .B(u0__abc_49347_n5345), .Y(u0__abc_49347_n5347) );
  OR2X2 OR2X2_1409 ( .A(u0__abc_49347_n5348), .B(u0__abc_49347_n5349), .Y(u0__abc_49347_n5350) );
  OR2X2 OR2X2_141 ( .A(u0__abc_49347_n1213), .B(u0__abc_49347_n1209_1), .Y(u0__abc_49347_n1214) );
  OR2X2 OR2X2_1410 ( .A(u0__abc_49347_n5347), .B(u0__abc_49347_n5350), .Y(u0__abc_49347_n5351) );
  OR2X2 OR2X2_1411 ( .A(u0__abc_49347_n5351), .B(u0__abc_49347_n5344), .Y(u0__abc_49347_n5352) );
  OR2X2 OR2X2_1412 ( .A(u0__abc_49347_n5353), .B(u0__abc_49347_n5354), .Y(u0__abc_49347_n5355) );
  OR2X2 OR2X2_1413 ( .A(u0__abc_49347_n5356), .B(u0__abc_49347_n5357), .Y(u0__abc_49347_n5358) );
  OR2X2 OR2X2_1414 ( .A(u0__abc_49347_n5358), .B(u0__abc_49347_n5355), .Y(u0__abc_49347_n5359) );
  OR2X2 OR2X2_1415 ( .A(u0__abc_49347_n5360), .B(u0__abc_49347_n5361), .Y(u0__abc_49347_n5362) );
  OR2X2 OR2X2_1416 ( .A(u0__abc_49347_n5363), .B(u0__abc_49347_n5364), .Y(u0__abc_49347_n5365) );
  OR2X2 OR2X2_1417 ( .A(u0__abc_49347_n5365), .B(u0__abc_49347_n5362), .Y(u0__abc_49347_n5366) );
  OR2X2 OR2X2_1418 ( .A(u0__abc_49347_n5359), .B(u0__abc_49347_n5366), .Y(u0__abc_49347_n5367) );
  OR2X2 OR2X2_1419 ( .A(u0__abc_49347_n5367), .B(u0__abc_49347_n5352), .Y(u0__abc_49347_n5368) );
  OR2X2 OR2X2_142 ( .A(u0__abc_49347_n1215), .B(u0__abc_49347_n1216), .Y(u0__abc_49347_n1217) );
  OR2X2 OR2X2_1420 ( .A(u0__abc_49347_n5368), .B(u0__abc_49347_n5337), .Y(rf_dout_22_) );
  OR2X2 OR2X2_1421 ( .A(u0__abc_49347_n5372), .B(u0__abc_49347_n5371), .Y(u0__abc_49347_n5373) );
  OR2X2 OR2X2_1422 ( .A(u0__abc_49347_n5375), .B(u0__abc_49347_n5374), .Y(u0__abc_49347_n5376) );
  OR2X2 OR2X2_1423 ( .A(u0__abc_49347_n5376), .B(u0__abc_49347_n5373), .Y(u0__abc_49347_n5377) );
  OR2X2 OR2X2_1424 ( .A(u0__abc_49347_n5379), .B(u0__abc_49347_n5378), .Y(u0__abc_49347_n5380) );
  OR2X2 OR2X2_1425 ( .A(u0__abc_49347_n5381), .B(u0__abc_49347_n5382), .Y(u0__abc_49347_n5383) );
  OR2X2 OR2X2_1426 ( .A(u0__abc_49347_n5380), .B(u0__abc_49347_n5383), .Y(u0__abc_49347_n5384) );
  OR2X2 OR2X2_1427 ( .A(u0__abc_49347_n5384), .B(u0__abc_49347_n5377), .Y(u0__abc_49347_n5385) );
  OR2X2 OR2X2_1428 ( .A(u0__abc_49347_n5386), .B(u0__abc_49347_n5387), .Y(u0__abc_49347_n5388) );
  OR2X2 OR2X2_1429 ( .A(u0__abc_49347_n5390), .B(u0__abc_49347_n5389), .Y(u0__abc_49347_n5391) );
  OR2X2 OR2X2_143 ( .A(u0__abc_49347_n1218_1), .B(u0__abc_49347_n1219_1), .Y(u0__abc_49347_n1220) );
  OR2X2 OR2X2_1430 ( .A(u0__abc_49347_n5388), .B(u0__abc_49347_n5391), .Y(u0__abc_49347_n5392) );
  OR2X2 OR2X2_1431 ( .A(u0__abc_49347_n5394), .B(u0__abc_49347_n5393), .Y(u0__abc_49347_n5395) );
  OR2X2 OR2X2_1432 ( .A(u0__abc_49347_n5396), .B(u0__abc_49347_n5397), .Y(u0__abc_49347_n5398) );
  OR2X2 OR2X2_1433 ( .A(u0__abc_49347_n5398), .B(u0__abc_49347_n5395), .Y(u0__abc_49347_n5399) );
  OR2X2 OR2X2_1434 ( .A(u0__abc_49347_n5392), .B(u0__abc_49347_n5399), .Y(u0__abc_49347_n5400) );
  OR2X2 OR2X2_1435 ( .A(u0__abc_49347_n5400), .B(u0__abc_49347_n5385), .Y(u0__abc_49347_n5401) );
  OR2X2 OR2X2_1436 ( .A(u0__abc_49347_n5401), .B(u0__abc_49347_n5370), .Y(rf_dout_23_) );
  OR2X2 OR2X2_1437 ( .A(u0__abc_49347_n5406), .B(u0__abc_49347_n5405), .Y(u0__abc_49347_n5407) );
  OR2X2 OR2X2_1438 ( .A(u0__abc_49347_n5407), .B(u0__abc_49347_n5404), .Y(u0__abc_49347_n5408) );
  OR2X2 OR2X2_1439 ( .A(u0__abc_49347_n5408), .B(u0__abc_49347_n5403), .Y(u0__abc_49347_n5409) );
  OR2X2 OR2X2_144 ( .A(u0__abc_49347_n1221), .B(u0__abc_49347_n1222), .Y(u0__abc_49347_n1223) );
  OR2X2 OR2X2_1440 ( .A(u0__abc_49347_n5412), .B(u0__abc_49347_n5411), .Y(u0__abc_49347_n5413) );
  OR2X2 OR2X2_1441 ( .A(u0__abc_49347_n5413), .B(u0__abc_49347_n5410), .Y(u0__abc_49347_n5414) );
  OR2X2 OR2X2_1442 ( .A(u0__abc_49347_n5416), .B(u0__abc_49347_n5417), .Y(u0__abc_49347_n5418) );
  OR2X2 OR2X2_1443 ( .A(u0__abc_49347_n5418), .B(u0__abc_49347_n5415), .Y(u0__abc_49347_n5419) );
  OR2X2 OR2X2_1444 ( .A(u0__abc_49347_n5419), .B(u0__abc_49347_n5414), .Y(u0__abc_49347_n5420) );
  OR2X2 OR2X2_1445 ( .A(u0__abc_49347_n5420), .B(u0__abc_49347_n5409), .Y(u0__abc_49347_n5421) );
  OR2X2 OR2X2_1446 ( .A(u0__abc_49347_n5423), .B(u0__abc_49347_n5424), .Y(u0__abc_49347_n5425) );
  OR2X2 OR2X2_1447 ( .A(u0__abc_49347_n5425), .B(u0__abc_49347_n5426), .Y(u0__abc_49347_n5427) );
  OR2X2 OR2X2_1448 ( .A(u0__abc_49347_n5428), .B(u0__abc_49347_n5429), .Y(u0__abc_49347_n5430) );
  OR2X2 OR2X2_1449 ( .A(u0__abc_49347_n5431), .B(u0__abc_49347_n5432), .Y(u0__abc_49347_n5433) );
  OR2X2 OR2X2_145 ( .A(u0__abc_49347_n1225), .B(spec_req_cs_0_bF_buf1), .Y(u0__abc_49347_n1226) );
  OR2X2 OR2X2_1450 ( .A(u0__abc_49347_n5430), .B(u0__abc_49347_n5433), .Y(u0__abc_49347_n5434) );
  OR2X2 OR2X2_1451 ( .A(u0__abc_49347_n5427), .B(u0__abc_49347_n5434), .Y(u0__abc_49347_n5435) );
  OR2X2 OR2X2_1452 ( .A(u0__abc_49347_n5422), .B(u0__abc_49347_n5435), .Y(u0__abc_49347_n5436) );
  OR2X2 OR2X2_1453 ( .A(u0__abc_49347_n5436), .B(u0__abc_49347_n5421), .Y(rf_dout_24_) );
  OR2X2 OR2X2_1454 ( .A(u0__abc_49347_n5440), .B(u0__abc_49347_n5441), .Y(u0__abc_49347_n5442) );
  OR2X2 OR2X2_1455 ( .A(u0__abc_49347_n5442), .B(u0__abc_49347_n5439), .Y(u0__abc_49347_n5443) );
  OR2X2 OR2X2_1456 ( .A(u0__abc_49347_n5445), .B(u0__abc_49347_n5446), .Y(u0__abc_49347_n5447) );
  OR2X2 OR2X2_1457 ( .A(u0__abc_49347_n5447), .B(u0__abc_49347_n5444), .Y(u0__abc_49347_n5448) );
  OR2X2 OR2X2_1458 ( .A(u0__abc_49347_n5448), .B(u0__abc_49347_n5443), .Y(u0__abc_49347_n5449) );
  OR2X2 OR2X2_1459 ( .A(u0__abc_49347_n5453), .B(u0__abc_49347_n5452), .Y(u0__abc_49347_n5454) );
  OR2X2 OR2X2_146 ( .A(u0__abc_49347_n1224), .B(u0__abc_49347_n1226), .Y(u0__abc_49347_n1227_1) );
  OR2X2 OR2X2_1460 ( .A(u0__abc_49347_n5454), .B(u0__abc_49347_n5451), .Y(u0__abc_49347_n5455) );
  OR2X2 OR2X2_1461 ( .A(u0__abc_49347_n5455), .B(u0__abc_49347_n5450), .Y(u0__abc_49347_n5456) );
  OR2X2 OR2X2_1462 ( .A(u0__abc_49347_n5458), .B(u0__abc_49347_n5459), .Y(u0__abc_49347_n5460) );
  OR2X2 OR2X2_1463 ( .A(u0__abc_49347_n5460), .B(u0__abc_49347_n5457), .Y(u0__abc_49347_n5461) );
  OR2X2 OR2X2_1464 ( .A(u0__abc_49347_n5462), .B(u0__abc_49347_n5463), .Y(u0__abc_49347_n5464) );
  OR2X2 OR2X2_1465 ( .A(u0__abc_49347_n5466), .B(u0__abc_49347_n5465), .Y(u0__abc_49347_n5467) );
  OR2X2 OR2X2_1466 ( .A(u0__abc_49347_n5467), .B(u0__abc_49347_n5464), .Y(u0__abc_49347_n5468) );
  OR2X2 OR2X2_1467 ( .A(u0__abc_49347_n5461), .B(u0__abc_49347_n5468), .Y(u0__abc_49347_n5469) );
  OR2X2 OR2X2_1468 ( .A(u0__abc_49347_n5469), .B(u0__abc_49347_n5456), .Y(u0__abc_49347_n5470) );
  OR2X2 OR2X2_1469 ( .A(u0__abc_49347_n5470), .B(u0__abc_49347_n5449), .Y(u0__abc_49347_n5471) );
  OR2X2 OR2X2_147 ( .A(u0__abc_49347_n1203_bF_buf4), .B(u0_tms0_1_), .Y(u0__abc_49347_n1228_1) );
  OR2X2 OR2X2_1470 ( .A(u0__abc_49347_n5471), .B(u0__abc_49347_n5438), .Y(rf_dout_25_) );
  OR2X2 OR2X2_1471 ( .A(u0__abc_49347_n5474), .B(u0__abc_49347_n5475), .Y(u0__abc_49347_n5476) );
  OR2X2 OR2X2_1472 ( .A(u0__abc_49347_n5477), .B(u0__abc_49347_n5478), .Y(u0__abc_49347_n5479) );
  OR2X2 OR2X2_1473 ( .A(u0__abc_49347_n5481), .B(u0__abc_49347_n5480), .Y(u0__abc_49347_n5482) );
  OR2X2 OR2X2_1474 ( .A(u0__abc_49347_n5479), .B(u0__abc_49347_n5482), .Y(u0__abc_49347_n5483) );
  OR2X2 OR2X2_1475 ( .A(u0__abc_49347_n5483), .B(u0__abc_49347_n5476), .Y(u0__abc_49347_n5484) );
  OR2X2 OR2X2_1476 ( .A(u0__abc_49347_n5486), .B(u0__abc_49347_n5487), .Y(u0__abc_49347_n5488) );
  OR2X2 OR2X2_1477 ( .A(u0__abc_49347_n5488), .B(u0__abc_49347_n5485), .Y(u0__abc_49347_n5489) );
  OR2X2 OR2X2_1478 ( .A(u0__abc_49347_n5490), .B(u0__abc_49347_n5491), .Y(u0__abc_49347_n5492) );
  OR2X2 OR2X2_1479 ( .A(u0__abc_49347_n5493), .B(u0__abc_49347_n5494), .Y(u0__abc_49347_n5495) );
  OR2X2 OR2X2_148 ( .A(u0__abc_49347_n1230), .B(u0__abc_49347_n1208), .Y(u0_sp_tms_1__FF_INPUT) );
  OR2X2 OR2X2_1480 ( .A(u0__abc_49347_n5492), .B(u0__abc_49347_n5495), .Y(u0__abc_49347_n5496) );
  OR2X2 OR2X2_1481 ( .A(u0__abc_49347_n5497), .B(u0__abc_49347_n5498), .Y(u0__abc_49347_n5499) );
  OR2X2 OR2X2_1482 ( .A(u0__abc_49347_n5500), .B(u0__abc_49347_n5501), .Y(u0__abc_49347_n5502) );
  OR2X2 OR2X2_1483 ( .A(u0__abc_49347_n5502), .B(u0__abc_49347_n5499), .Y(u0__abc_49347_n5503) );
  OR2X2 OR2X2_1484 ( .A(u0__abc_49347_n5496), .B(u0__abc_49347_n5503), .Y(u0__abc_49347_n5504) );
  OR2X2 OR2X2_1485 ( .A(u0__abc_49347_n5504), .B(u0__abc_49347_n5489), .Y(u0__abc_49347_n5505) );
  OR2X2 OR2X2_1486 ( .A(u0__abc_49347_n5505), .B(u0__abc_49347_n5484), .Y(u0__abc_49347_n5506) );
  OR2X2 OR2X2_1487 ( .A(u0__abc_49347_n5506), .B(u0__abc_49347_n5473), .Y(rf_dout_26_) );
  OR2X2 OR2X2_1488 ( .A(u0__abc_49347_n5510), .B(u0__abc_49347_n5511), .Y(u0__abc_49347_n5512) );
  OR2X2 OR2X2_1489 ( .A(u0__abc_49347_n5512), .B(u0__abc_49347_n5509), .Y(u0__abc_49347_n5513) );
  OR2X2 OR2X2_149 ( .A(u0__abc_49347_n1183_1_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n1234) );
  OR2X2 OR2X2_1490 ( .A(u0__abc_49347_n5516), .B(u0__abc_49347_n5515), .Y(u0__abc_49347_n5517) );
  OR2X2 OR2X2_1491 ( .A(u0__abc_49347_n5517), .B(u0__abc_49347_n5514), .Y(u0__abc_49347_n5518) );
  OR2X2 OR2X2_1492 ( .A(u0__abc_49347_n5513), .B(u0__abc_49347_n5518), .Y(u0__abc_49347_n5519) );
  OR2X2 OR2X2_1493 ( .A(u0__abc_49347_n5522), .B(u0__abc_49347_n5521), .Y(u0__abc_49347_n5523) );
  OR2X2 OR2X2_1494 ( .A(u0__abc_49347_n5523), .B(u0__abc_49347_n5520), .Y(u0__abc_49347_n5524) );
  OR2X2 OR2X2_1495 ( .A(u0__abc_49347_n5526), .B(u0__abc_49347_n5527), .Y(u0__abc_49347_n5528) );
  OR2X2 OR2X2_1496 ( .A(u0__abc_49347_n5528), .B(u0__abc_49347_n5525), .Y(u0__abc_49347_n5529) );
  OR2X2 OR2X2_1497 ( .A(u0__abc_49347_n5529), .B(u0__abc_49347_n5524), .Y(u0__abc_49347_n5530) );
  OR2X2 OR2X2_1498 ( .A(u0__abc_49347_n5533), .B(u0__abc_49347_n5532), .Y(u0__abc_49347_n5534) );
  OR2X2 OR2X2_1499 ( .A(u0__abc_49347_n5534), .B(u0__abc_49347_n5531), .Y(u0__abc_49347_n5535) );
  OR2X2 OR2X2_15 ( .A(_abc_55805_n240_bF_buf2), .B(spec_req_cs_3_bF_buf5), .Y(_abc_55805_n260) );
  OR2X2 OR2X2_150 ( .A(spec_req_cs_6_bF_buf0), .B(1'b0), .Y(u0__abc_49347_n1235) );
  OR2X2 OR2X2_1500 ( .A(u0__abc_49347_n5536), .B(u0__abc_49347_n5537), .Y(u0__abc_49347_n5538) );
  OR2X2 OR2X2_1501 ( .A(u0__abc_49347_n5535), .B(u0__abc_49347_n5538), .Y(u0__abc_49347_n5539) );
  OR2X2 OR2X2_1502 ( .A(u0__abc_49347_n5530), .B(u0__abc_49347_n5539), .Y(u0__abc_49347_n5540) );
  OR2X2 OR2X2_1503 ( .A(u0__abc_49347_n5540), .B(u0__abc_49347_n5519), .Y(u0__abc_49347_n5541) );
  OR2X2 OR2X2_1504 ( .A(u0__abc_49347_n5541), .B(u0__abc_49347_n5508), .Y(rf_dout_27_) );
  OR2X2 OR2X2_1505 ( .A(u0__abc_49347_n5545), .B(u0__abc_49347_n5546), .Y(u0__abc_49347_n5547) );
  OR2X2 OR2X2_1506 ( .A(u0__abc_49347_n5547), .B(u0__abc_49347_n5544), .Y(u0__abc_49347_n5548) );
  OR2X2 OR2X2_1507 ( .A(u0__abc_49347_n5550), .B(u0__abc_49347_n5551), .Y(u0__abc_49347_n5552) );
  OR2X2 OR2X2_1508 ( .A(u0__abc_49347_n5552), .B(u0__abc_49347_n5549), .Y(u0__abc_49347_n5553) );
  OR2X2 OR2X2_1509 ( .A(u0__abc_49347_n5553), .B(u0__abc_49347_n5548), .Y(u0__abc_49347_n5554) );
  OR2X2 OR2X2_151 ( .A(u0__abc_49347_n1237_1), .B(u0__abc_49347_n1233), .Y(u0__abc_49347_n1238) );
  OR2X2 OR2X2_1510 ( .A(u0__abc_49347_n5558), .B(u0__abc_49347_n5557), .Y(u0__abc_49347_n5559) );
  OR2X2 OR2X2_1511 ( .A(u0__abc_49347_n5559), .B(u0__abc_49347_n5556), .Y(u0__abc_49347_n5560) );
  OR2X2 OR2X2_1512 ( .A(u0__abc_49347_n5560), .B(u0__abc_49347_n5555), .Y(u0__abc_49347_n5561) );
  OR2X2 OR2X2_1513 ( .A(u0__abc_49347_n5563), .B(u0__abc_49347_n5564), .Y(u0__abc_49347_n5565) );
  OR2X2 OR2X2_1514 ( .A(u0__abc_49347_n5565), .B(u0__abc_49347_n5562), .Y(u0__abc_49347_n5566) );
  OR2X2 OR2X2_1515 ( .A(u0__abc_49347_n5567), .B(u0__abc_49347_n5568), .Y(u0__abc_49347_n5569) );
  OR2X2 OR2X2_1516 ( .A(u0__abc_49347_n5571), .B(u0__abc_49347_n5570), .Y(u0__abc_49347_n5572) );
  OR2X2 OR2X2_1517 ( .A(u0__abc_49347_n5572), .B(u0__abc_49347_n5569), .Y(u0__abc_49347_n5573) );
  OR2X2 OR2X2_1518 ( .A(u0__abc_49347_n5566), .B(u0__abc_49347_n5573), .Y(u0__abc_49347_n5574) );
  OR2X2 OR2X2_1519 ( .A(u0__abc_49347_n5574), .B(u0__abc_49347_n5561), .Y(u0__abc_49347_n5575) );
  OR2X2 OR2X2_152 ( .A(u0__abc_49347_n1239), .B(u0__abc_49347_n1240), .Y(u0__abc_49347_n1241) );
  OR2X2 OR2X2_1520 ( .A(u0__abc_49347_n5575), .B(u0__abc_49347_n5554), .Y(u0__abc_49347_n5576) );
  OR2X2 OR2X2_1521 ( .A(u0__abc_49347_n5576), .B(u0__abc_49347_n5543), .Y(rf_dout_28_) );
  OR2X2 OR2X2_1522 ( .A(u0__abc_49347_n5579), .B(u0__abc_49347_n5578), .Y(u0__abc_49347_n5580) );
  OR2X2 OR2X2_1523 ( .A(u0__abc_49347_n5582), .B(u0__abc_49347_n5581), .Y(u0__abc_49347_n5583) );
  OR2X2 OR2X2_1524 ( .A(u0__abc_49347_n5584), .B(u0__abc_49347_n5585), .Y(u0__abc_49347_n5586) );
  OR2X2 OR2X2_1525 ( .A(u0__abc_49347_n5586), .B(u0__abc_49347_n5583), .Y(u0__abc_49347_n5587) );
  OR2X2 OR2X2_1526 ( .A(u0__abc_49347_n5587), .B(u0__abc_49347_n5580), .Y(u0__abc_49347_n5588) );
  OR2X2 OR2X2_1527 ( .A(u0__abc_49347_n5590), .B(u0__abc_49347_n5591), .Y(u0__abc_49347_n5592) );
  OR2X2 OR2X2_1528 ( .A(u0__abc_49347_n5592), .B(u0__abc_49347_n5589), .Y(u0__abc_49347_n5593) );
  OR2X2 OR2X2_1529 ( .A(u0__abc_49347_n5595), .B(u0__abc_49347_n5596), .Y(u0__abc_49347_n5597) );
  OR2X2 OR2X2_153 ( .A(u0__abc_49347_n1242), .B(u0__abc_49347_n1243), .Y(u0__abc_49347_n1244) );
  OR2X2 OR2X2_1530 ( .A(u0__abc_49347_n5597), .B(u0__abc_49347_n5594), .Y(u0__abc_49347_n5598) );
  OR2X2 OR2X2_1531 ( .A(u0__abc_49347_n5593), .B(u0__abc_49347_n5598), .Y(u0__abc_49347_n5599) );
  OR2X2 OR2X2_1532 ( .A(u0__abc_49347_n5599), .B(u0__abc_49347_n5588), .Y(u0__abc_49347_n5600) );
  OR2X2 OR2X2_1533 ( .A(u0__abc_49347_n5604), .B(u0__abc_49347_n5603), .Y(u0__abc_49347_n5605) );
  OR2X2 OR2X2_1534 ( .A(u0__abc_49347_n5605), .B(u0__abc_49347_n5602), .Y(u0__abc_49347_n5606) );
  OR2X2 OR2X2_1535 ( .A(u0__abc_49347_n5607), .B(u0__abc_49347_n5608), .Y(u0__abc_49347_n5609) );
  OR2X2 OR2X2_1536 ( .A(u0__abc_49347_n5606), .B(u0__abc_49347_n5609), .Y(u0__abc_49347_n5610) );
  OR2X2 OR2X2_1537 ( .A(u0__abc_49347_n5601), .B(u0__abc_49347_n5610), .Y(u0__abc_49347_n5611) );
  OR2X2 OR2X2_1538 ( .A(u0__abc_49347_n5611), .B(u0__abc_49347_n5600), .Y(rf_dout_29_) );
  OR2X2 OR2X2_1539 ( .A(u0__abc_49347_n5614), .B(u0__abc_49347_n5615), .Y(u0__abc_49347_n5616) );
  OR2X2 OR2X2_154 ( .A(u0__abc_49347_n1245_1), .B(u0__abc_49347_n1246_1), .Y(u0__abc_49347_n1247) );
  OR2X2 OR2X2_1540 ( .A(u0__abc_49347_n5618), .B(u0__abc_49347_n5617), .Y(u0__abc_49347_n5619) );
  OR2X2 OR2X2_1541 ( .A(u0__abc_49347_n5620), .B(u0__abc_49347_n5621), .Y(u0__abc_49347_n5622) );
  OR2X2 OR2X2_1542 ( .A(u0__abc_49347_n5619), .B(u0__abc_49347_n5622), .Y(u0__abc_49347_n5623) );
  OR2X2 OR2X2_1543 ( .A(u0__abc_49347_n5623), .B(u0__abc_49347_n5616), .Y(u0__abc_49347_n5624) );
  OR2X2 OR2X2_1544 ( .A(u0__abc_49347_n5626), .B(u0__abc_49347_n5627), .Y(u0__abc_49347_n5628) );
  OR2X2 OR2X2_1545 ( .A(u0__abc_49347_n5628), .B(u0__abc_49347_n5625), .Y(u0__abc_49347_n5629) );
  OR2X2 OR2X2_1546 ( .A(u0__abc_49347_n5631), .B(u0__abc_49347_n5632), .Y(u0__abc_49347_n5633) );
  OR2X2 OR2X2_1547 ( .A(u0__abc_49347_n5633), .B(u0__abc_49347_n5630), .Y(u0__abc_49347_n5634) );
  OR2X2 OR2X2_1548 ( .A(u0__abc_49347_n5634), .B(u0__abc_49347_n5629), .Y(u0__abc_49347_n5635) );
  OR2X2 OR2X2_1549 ( .A(u0__abc_49347_n5638), .B(u0__abc_49347_n5637), .Y(u0__abc_49347_n5639) );
  OR2X2 OR2X2_155 ( .A(u0__abc_49347_n1249), .B(spec_req_cs_0_bF_buf0), .Y(u0__abc_49347_n1250) );
  OR2X2 OR2X2_1550 ( .A(u0__abc_49347_n5639), .B(u0__abc_49347_n5636), .Y(u0__abc_49347_n5640) );
  OR2X2 OR2X2_1551 ( .A(u0__abc_49347_n5641), .B(u0__abc_49347_n5642), .Y(u0__abc_49347_n5643) );
  OR2X2 OR2X2_1552 ( .A(u0__abc_49347_n5640), .B(u0__abc_49347_n5643), .Y(u0__abc_49347_n5644) );
  OR2X2 OR2X2_1553 ( .A(u0__abc_49347_n5635), .B(u0__abc_49347_n5644), .Y(u0__abc_49347_n5645) );
  OR2X2 OR2X2_1554 ( .A(u0__abc_49347_n5645), .B(u0__abc_49347_n5624), .Y(u0__abc_49347_n5646) );
  OR2X2 OR2X2_1555 ( .A(u0__abc_49347_n5646), .B(u0__abc_49347_n5613), .Y(rf_dout_30_) );
  OR2X2 OR2X2_1556 ( .A(u0__abc_49347_n5649), .B(u0__abc_49347_n5650), .Y(u0__abc_49347_n5651) );
  OR2X2 OR2X2_1557 ( .A(u0__abc_49347_n5653), .B(u0__abc_49347_n5652), .Y(u0__abc_49347_n5654) );
  OR2X2 OR2X2_1558 ( .A(u0__abc_49347_n5655), .B(u0__abc_49347_n5656), .Y(u0__abc_49347_n5657) );
  OR2X2 OR2X2_1559 ( .A(u0__abc_49347_n5657), .B(u0__abc_49347_n5654), .Y(u0__abc_49347_n5658) );
  OR2X2 OR2X2_156 ( .A(u0__abc_49347_n1248), .B(u0__abc_49347_n1250), .Y(u0__abc_49347_n1251) );
  OR2X2 OR2X2_1560 ( .A(u0__abc_49347_n5658), .B(u0__abc_49347_n5651), .Y(u0__abc_49347_n5659) );
  OR2X2 OR2X2_1561 ( .A(u0__abc_49347_n5663), .B(u0__abc_49347_n5662), .Y(u0__abc_49347_n5664) );
  OR2X2 OR2X2_1562 ( .A(u0__abc_49347_n5664), .B(u0__abc_49347_n5661), .Y(u0__abc_49347_n5665) );
  OR2X2 OR2X2_1563 ( .A(u0__abc_49347_n5665), .B(u0__abc_49347_n5660), .Y(u0__abc_49347_n5666) );
  OR2X2 OR2X2_1564 ( .A(u0__abc_49347_n5667), .B(u0__abc_49347_n5668), .Y(u0__abc_49347_n5669) );
  OR2X2 OR2X2_1565 ( .A(u0__abc_49347_n5669), .B(u0__abc_49347_n5670), .Y(u0__abc_49347_n5671) );
  OR2X2 OR2X2_1566 ( .A(u0__abc_49347_n5672), .B(u0__abc_49347_n5673), .Y(u0__abc_49347_n5674) );
  OR2X2 OR2X2_1567 ( .A(u0__abc_49347_n5675), .B(u0__abc_49347_n5676), .Y(u0__abc_49347_n5677) );
  OR2X2 OR2X2_1568 ( .A(u0__abc_49347_n5674), .B(u0__abc_49347_n5677), .Y(u0__abc_49347_n5678) );
  OR2X2 OR2X2_1569 ( .A(u0__abc_49347_n5671), .B(u0__abc_49347_n5678), .Y(u0__abc_49347_n5679) );
  OR2X2 OR2X2_157 ( .A(u0__abc_49347_n1203_bF_buf3), .B(u0_tms0_2_), .Y(u0__abc_49347_n1252) );
  OR2X2 OR2X2_1570 ( .A(u0__abc_49347_n5679), .B(u0__abc_49347_n5666), .Y(u0__abc_49347_n5680) );
  OR2X2 OR2X2_1571 ( .A(u0__abc_49347_n5680), .B(u0__abc_49347_n5659), .Y(u0__abc_49347_n5681) );
  OR2X2 OR2X2_1572 ( .A(u0__abc_49347_n5681), .B(u0__abc_49347_n5648), .Y(rf_dout_31_) );
  OR2X2 OR2X2_1573 ( .A(u0__abc_49347_n5743), .B(u0__abc_49347_n5745), .Y(u0__abc_49347_n5746) );
  OR2X2 OR2X2_1574 ( .A(u0__abc_49347_n5746), .B(u0__abc_49347_n5741), .Y(u0_sreq_cs_le_FF_INPUT) );
  OR2X2 OR2X2_1575 ( .A(u0_init_req4), .B(u0_init_req5), .Y(u0__abc_49347_n5748) );
  OR2X2 OR2X2_1576 ( .A(1'b0), .B(1'b0), .Y(u0__abc_49347_n5749) );
  OR2X2 OR2X2_1577 ( .A(u0__abc_49347_n5748), .B(u0__abc_49347_n5749), .Y(u0__abc_49347_n5750) );
  OR2X2 OR2X2_1578 ( .A(u0_init_req0), .B(u0_init_req1), .Y(u0__abc_49347_n5751) );
  OR2X2 OR2X2_1579 ( .A(u0_init_req2), .B(u0_init_req3), .Y(u0__abc_49347_n5752) );
  OR2X2 OR2X2_158 ( .A(u0__abc_49347_n1254_1), .B(u0__abc_49347_n1232), .Y(u0_sp_tms_2__FF_INPUT) );
  OR2X2 OR2X2_1580 ( .A(u0__abc_49347_n5751), .B(u0__abc_49347_n5752), .Y(u0__abc_49347_n5753) );
  OR2X2 OR2X2_1581 ( .A(u0__abc_49347_n5750), .B(u0__abc_49347_n5753), .Y(u0_init_req_FF_INPUT) );
  OR2X2 OR2X2_1582 ( .A(u0_lmr_req4), .B(u0_lmr_req5), .Y(u0__abc_49347_n5755) );
  OR2X2 OR2X2_1583 ( .A(1'b0), .B(1'b0), .Y(u0__abc_49347_n5756) );
  OR2X2 OR2X2_1584 ( .A(u0__abc_49347_n5755), .B(u0__abc_49347_n5756), .Y(u0__abc_49347_n5757) );
  OR2X2 OR2X2_1585 ( .A(u0_lmr_req0), .B(u0_lmr_req1), .Y(u0__abc_49347_n5758) );
  OR2X2 OR2X2_1586 ( .A(u0_lmr_req2), .B(u0_lmr_req3), .Y(u0__abc_49347_n5759) );
  OR2X2 OR2X2_1587 ( .A(u0__abc_49347_n5758), .B(u0__abc_49347_n5759), .Y(u0__abc_49347_n5760) );
  OR2X2 OR2X2_1588 ( .A(u0__abc_49347_n5757), .B(u0__abc_49347_n5760), .Y(u0_lmr_req_FF_INPUT) );
  OR2X2 OR2X2_1589 ( .A(u0_csc0_2_), .B(u0_csc0_1_), .Y(u0_u0__abc_43300_n201_1) );
  OR2X2 OR2X2_159 ( .A(u0__abc_49347_n1183_1_bF_buf2), .B(1'b0), .Y(u0__abc_49347_n1258) );
  OR2X2 OR2X2_1590 ( .A(u0_u0__abc_43300_n201_1), .B(u0_csc0_3_), .Y(u0_u0__abc_43300_n202_1) );
  OR2X2 OR2X2_1591 ( .A(u0_u0__abc_43300_n209), .B(u0_u0__abc_43300_n205_1), .Y(u0_u0_lmr_req_FF_INPUT) );
  OR2X2 OR2X2_1592 ( .A(u0_u0_addr_r_5_), .B(u0_u0_addr_r_3_), .Y(u0_u0__abc_43300_n212) );
  OR2X2 OR2X2_1593 ( .A(u0_u0__abc_43300_n212), .B(u0_u0_addr_r_6_), .Y(u0_u0__abc_43300_n213_1) );
  OR2X2 OR2X2_1594 ( .A(u0_u0_lmr_req_we_FF_INPUT_bF_buf4), .B(u0_tms0_0_), .Y(u0_u0__abc_43300_n217_1) );
  OR2X2 OR2X2_1595 ( .A(u0_u0__abc_43300_n219_1_bF_buf4), .B(\wb_data_i[0] ), .Y(u0_u0__abc_43300_n220_1) );
  OR2X2 OR2X2_1596 ( .A(u0_u0_lmr_req_we_FF_INPUT_bF_buf2), .B(u0_tms0_1_), .Y(u0_u0__abc_43300_n223_1) );
  OR2X2 OR2X2_1597 ( .A(u0_u0__abc_43300_n219_1_bF_buf3), .B(\wb_data_i[1] ), .Y(u0_u0__abc_43300_n224) );
  OR2X2 OR2X2_1598 ( .A(u0_u0_lmr_req_we_FF_INPUT_bF_buf1), .B(u0_tms0_2_), .Y(u0_u0__abc_43300_n227) );
  OR2X2 OR2X2_1599 ( .A(u0_u0__abc_43300_n219_1_bF_buf2), .B(\wb_data_i[2] ), .Y(u0_u0__abc_43300_n228_1) );
  OR2X2 OR2X2_16 ( .A(lmr_sel_bF_buf3), .B(cs_3_), .Y(_abc_55805_n261) );
  OR2X2 OR2X2_160 ( .A(spec_req_cs_6_bF_buf5), .B(1'b0), .Y(u0__abc_49347_n1259) );
  OR2X2 OR2X2_1600 ( .A(u0_u0_lmr_req_we_FF_INPUT_bF_buf0), .B(u0_tms0_3_), .Y(u0_u0__abc_43300_n231_1) );
  OR2X2 OR2X2_1601 ( .A(u0_u0__abc_43300_n219_1_bF_buf1), .B(\wb_data_i[3] ), .Y(u0_u0__abc_43300_n232_1) );
  OR2X2 OR2X2_1602 ( .A(u0_u0_lmr_req_we_FF_INPUT_bF_buf4), .B(u0_tms0_4_), .Y(u0_u0__abc_43300_n235_1) );
  OR2X2 OR2X2_1603 ( .A(u0_u0__abc_43300_n219_1_bF_buf0), .B(\wb_data_i[4] ), .Y(u0_u0__abc_43300_n236) );
  OR2X2 OR2X2_1604 ( .A(u0_u0_lmr_req_we_FF_INPUT_bF_buf3), .B(u0_tms0_5_), .Y(u0_u0__abc_43300_n239) );
  OR2X2 OR2X2_1605 ( .A(u0_u0__abc_43300_n219_1_bF_buf4), .B(\wb_data_i[5] ), .Y(u0_u0__abc_43300_n240_1) );
  OR2X2 OR2X2_1606 ( .A(u0_u0_lmr_req_we_FF_INPUT_bF_buf2), .B(u0_tms0_6_), .Y(u0_u0__abc_43300_n243_1) );
  OR2X2 OR2X2_1607 ( .A(u0_u0__abc_43300_n219_1_bF_buf3), .B(\wb_data_i[6] ), .Y(u0_u0__abc_43300_n244_1) );
  OR2X2 OR2X2_1608 ( .A(u0_u0_lmr_req_we_FF_INPUT_bF_buf1), .B(u0_tms0_7_), .Y(u0_u0__abc_43300_n247_1) );
  OR2X2 OR2X2_1609 ( .A(u0_u0__abc_43300_n219_1_bF_buf2), .B(\wb_data_i[7] ), .Y(u0_u0__abc_43300_n248) );
  OR2X2 OR2X2_161 ( .A(u0__abc_49347_n1261), .B(u0__abc_49347_n1257), .Y(u0__abc_49347_n1262) );
  OR2X2 OR2X2_1610 ( .A(u0_u0_lmr_req_we_FF_INPUT_bF_buf0), .B(u0_tms0_8_), .Y(u0_u0__abc_43300_n251) );
  OR2X2 OR2X2_1611 ( .A(u0_u0__abc_43300_n219_1_bF_buf1), .B(\wb_data_i[8] ), .Y(u0_u0__abc_43300_n252_1) );
  OR2X2 OR2X2_1612 ( .A(u0_u0_lmr_req_we_FF_INPUT_bF_buf4), .B(u0_tms0_9_), .Y(u0_u0__abc_43300_n255_1) );
  OR2X2 OR2X2_1613 ( .A(u0_u0__abc_43300_n219_1_bF_buf0), .B(\wb_data_i[9] ), .Y(u0_u0__abc_43300_n256) );
  OR2X2 OR2X2_1614 ( .A(u0_u0_lmr_req_we_FF_INPUT_bF_buf3), .B(u0_tms0_10_), .Y(u0_u0__abc_43300_n259) );
  OR2X2 OR2X2_1615 ( .A(u0_u0__abc_43300_n219_1_bF_buf4), .B(\wb_data_i[10] ), .Y(u0_u0__abc_43300_n260_1) );
  OR2X2 OR2X2_1616 ( .A(u0_u0_lmr_req_we_FF_INPUT_bF_buf2), .B(u0_tms0_11_), .Y(u0_u0__abc_43300_n263) );
  OR2X2 OR2X2_1617 ( .A(u0_u0__abc_43300_n219_1_bF_buf3), .B(\wb_data_i[11] ), .Y(u0_u0__abc_43300_n264) );
  OR2X2 OR2X2_1618 ( .A(u0_u0_lmr_req_we_FF_INPUT_bF_buf1), .B(u0_tms0_12_), .Y(u0_u0__abc_43300_n267) );
  OR2X2 OR2X2_1619 ( .A(u0_u0__abc_43300_n219_1_bF_buf2), .B(\wb_data_i[12] ), .Y(u0_u0__abc_43300_n268_1) );
  OR2X2 OR2X2_162 ( .A(u0__abc_49347_n1263_1), .B(u0__abc_49347_n1264_1), .Y(u0__abc_49347_n1265) );
  OR2X2 OR2X2_1620 ( .A(u0_u0_lmr_req_we_FF_INPUT_bF_buf0), .B(u0_tms0_13_), .Y(u0_u0__abc_43300_n271) );
  OR2X2 OR2X2_1621 ( .A(u0_u0__abc_43300_n219_1_bF_buf1), .B(\wb_data_i[13] ), .Y(u0_u0__abc_43300_n272) );
  OR2X2 OR2X2_1622 ( .A(u0_u0_lmr_req_we_FF_INPUT_bF_buf4), .B(u0_tms0_14_), .Y(u0_u0__abc_43300_n275_1) );
  OR2X2 OR2X2_1623 ( .A(u0_u0__abc_43300_n219_1_bF_buf0), .B(\wb_data_i[14] ), .Y(u0_u0__abc_43300_n276) );
  OR2X2 OR2X2_1624 ( .A(u0_u0_lmr_req_we_FF_INPUT_bF_buf3), .B(u0_tms0_15_), .Y(u0_u0__abc_43300_n279_1) );
  OR2X2 OR2X2_1625 ( .A(u0_u0__abc_43300_n219_1_bF_buf4), .B(\wb_data_i[15] ), .Y(u0_u0__abc_43300_n280) );
  OR2X2 OR2X2_1626 ( .A(u0_u0_lmr_req_we_FF_INPUT_bF_buf2), .B(u0_tms0_16_), .Y(u0_u0__abc_43300_n283_1) );
  OR2X2 OR2X2_1627 ( .A(u0_u0__abc_43300_n219_1_bF_buf3), .B(\wb_data_i[16] ), .Y(u0_u0__abc_43300_n284) );
  OR2X2 OR2X2_1628 ( .A(u0_u0_lmr_req_we_FF_INPUT_bF_buf1), .B(u0_tms0_17_), .Y(u0_u0__abc_43300_n287_1) );
  OR2X2 OR2X2_1629 ( .A(u0_u0__abc_43300_n219_1_bF_buf2), .B(\wb_data_i[17] ), .Y(u0_u0__abc_43300_n288) );
  OR2X2 OR2X2_163 ( .A(u0__abc_49347_n1266), .B(u0__abc_49347_n1267), .Y(u0__abc_49347_n1268) );
  OR2X2 OR2X2_1630 ( .A(u0_u0_lmr_req_we_FF_INPUT_bF_buf0), .B(u0_tms0_18_), .Y(u0_u0__abc_43300_n291) );
  OR2X2 OR2X2_1631 ( .A(u0_u0__abc_43300_n219_1_bF_buf1), .B(\wb_data_i[18] ), .Y(u0_u0__abc_43300_n292) );
  OR2X2 OR2X2_1632 ( .A(u0_u0_lmr_req_we_FF_INPUT_bF_buf4), .B(u0_tms0_19_), .Y(u0_u0__abc_43300_n295) );
  OR2X2 OR2X2_1633 ( .A(u0_u0__abc_43300_n219_1_bF_buf0), .B(\wb_data_i[19] ), .Y(u0_u0__abc_43300_n296_1) );
  OR2X2 OR2X2_1634 ( .A(u0_u0_lmr_req_we_FF_INPUT_bF_buf3), .B(u0_tms0_20_), .Y(u0_u0__abc_43300_n299) );
  OR2X2 OR2X2_1635 ( .A(u0_u0__abc_43300_n219_1_bF_buf4), .B(\wb_data_i[20] ), .Y(u0_u0__abc_43300_n300) );
  OR2X2 OR2X2_1636 ( .A(u0_u0_lmr_req_we_FF_INPUT_bF_buf2), .B(u0_tms0_21_), .Y(u0_u0__abc_43300_n303) );
  OR2X2 OR2X2_1637 ( .A(u0_u0__abc_43300_n219_1_bF_buf3), .B(\wb_data_i[21] ), .Y(u0_u0__abc_43300_n304) );
  OR2X2 OR2X2_1638 ( .A(u0_u0_lmr_req_we_FF_INPUT_bF_buf1), .B(u0_tms0_22_), .Y(u0_u0__abc_43300_n307) );
  OR2X2 OR2X2_1639 ( .A(u0_u0__abc_43300_n219_1_bF_buf2), .B(\wb_data_i[22] ), .Y(u0_u0__abc_43300_n308) );
  OR2X2 OR2X2_164 ( .A(u0__abc_49347_n1269), .B(u0__abc_49347_n1270), .Y(u0__abc_49347_n1271) );
  OR2X2 OR2X2_1640 ( .A(u0_u0_lmr_req_we_FF_INPUT_bF_buf0), .B(u0_tms0_23_), .Y(u0_u0__abc_43300_n311) );
  OR2X2 OR2X2_1641 ( .A(u0_u0__abc_43300_n219_1_bF_buf1), .B(\wb_data_i[23] ), .Y(u0_u0__abc_43300_n312_1) );
  OR2X2 OR2X2_1642 ( .A(u0_u0_lmr_req_we_FF_INPUT_bF_buf4), .B(u0_tms0_24_), .Y(u0_u0__abc_43300_n315_1) );
  OR2X2 OR2X2_1643 ( .A(u0_u0__abc_43300_n219_1_bF_buf0), .B(\wb_data_i[24] ), .Y(u0_u0__abc_43300_n316_1) );
  OR2X2 OR2X2_1644 ( .A(u0_u0_lmr_req_we_FF_INPUT_bF_buf3), .B(u0_tms0_25_), .Y(u0_u0__abc_43300_n319) );
  OR2X2 OR2X2_1645 ( .A(u0_u0__abc_43300_n219_1_bF_buf4), .B(\wb_data_i[25] ), .Y(u0_u0__abc_43300_n320) );
  OR2X2 OR2X2_1646 ( .A(u0_u0_lmr_req_we_FF_INPUT_bF_buf2), .B(u0_tms0_26_), .Y(u0_u0__abc_43300_n323_1) );
  OR2X2 OR2X2_1647 ( .A(u0_u0__abc_43300_n219_1_bF_buf3), .B(\wb_data_i[26] ), .Y(u0_u0__abc_43300_n324_1) );
  OR2X2 OR2X2_1648 ( .A(u0_u0_lmr_req_we_FF_INPUT_bF_buf1), .B(u0_tms0_27_), .Y(u0_u0__abc_43300_n327) );
  OR2X2 OR2X2_1649 ( .A(u0_u0__abc_43300_n219_1_bF_buf2), .B(\wb_data_i[27] ), .Y(u0_u0__abc_43300_n328) );
  OR2X2 OR2X2_165 ( .A(u0__abc_49347_n1273_1), .B(spec_req_cs_0_bF_buf5), .Y(u0__abc_49347_n1274) );
  OR2X2 OR2X2_1650 ( .A(u0_u0_lmr_req_we_FF_INPUT_bF_buf0), .B(u0_tms0_28_), .Y(u0_u0__abc_43300_n331) );
  OR2X2 OR2X2_1651 ( .A(u0_u0__abc_43300_n219_1_bF_buf1), .B(\wb_data_i[28] ), .Y(u0_u0__abc_43300_n332) );
  OR2X2 OR2X2_1652 ( .A(u0_u0_lmr_req_we_FF_INPUT_bF_buf4), .B(u0_tms0_29_), .Y(u0_u0__abc_43300_n335) );
  OR2X2 OR2X2_1653 ( .A(u0_u0__abc_43300_n219_1_bF_buf0), .B(\wb_data_i[29] ), .Y(u0_u0__abc_43300_n336) );
  OR2X2 OR2X2_1654 ( .A(u0_u0_lmr_req_we_FF_INPUT_bF_buf3), .B(u0_tms0_30_), .Y(u0_u0__abc_43300_n339) );
  OR2X2 OR2X2_1655 ( .A(u0_u0__abc_43300_n219_1_bF_buf4), .B(\wb_data_i[30] ), .Y(u0_u0__abc_43300_n340) );
  OR2X2 OR2X2_1656 ( .A(u0_u0_lmr_req_we_FF_INPUT_bF_buf2), .B(u0_tms0_31_), .Y(u0_u0__abc_43300_n343) );
  OR2X2 OR2X2_1657 ( .A(u0_u0__abc_43300_n219_1_bF_buf3), .B(\wb_data_i[31] ), .Y(u0_u0__abc_43300_n344) );
  OR2X2 OR2X2_1658 ( .A(u0_u0_init_req_we_FF_INPUT_bF_buf4), .B(u0_csc0_0_), .Y(u0_u0__abc_43300_n349) );
  OR2X2 OR2X2_1659 ( .A(u0_u0__abc_43300_n350_bF_buf4), .B(\wb_data_i[0] ), .Y(u0_u0__abc_43300_n351) );
  OR2X2 OR2X2_166 ( .A(u0__abc_49347_n1272_1), .B(u0__abc_49347_n1274), .Y(u0__abc_49347_n1275) );
  OR2X2 OR2X2_1660 ( .A(u0_u0_init_req_we_FF_INPUT_bF_buf2), .B(u0_csc0_1_), .Y(u0_u0__abc_43300_n354) );
  OR2X2 OR2X2_1661 ( .A(u0_u0__abc_43300_n350_bF_buf3), .B(\wb_data_i[1] ), .Y(u0_u0__abc_43300_n355) );
  OR2X2 OR2X2_1662 ( .A(u0_u0_init_req_we_FF_INPUT_bF_buf1), .B(u0_csc0_2_), .Y(u0_u0__abc_43300_n358) );
  OR2X2 OR2X2_1663 ( .A(u0_u0__abc_43300_n350_bF_buf2), .B(\wb_data_i[2] ), .Y(u0_u0__abc_43300_n359) );
  OR2X2 OR2X2_1664 ( .A(u0_u0_init_req_we_FF_INPUT_bF_buf0), .B(u0_csc0_3_), .Y(u0_u0__abc_43300_n362) );
  OR2X2 OR2X2_1665 ( .A(u0_u0__abc_43300_n350_bF_buf1), .B(\wb_data_i[3] ), .Y(u0_u0__abc_43300_n363) );
  OR2X2 OR2X2_1666 ( .A(u0_u0_init_req_we_FF_INPUT_bF_buf4), .B(u0_csc0_4_), .Y(u0_u0__abc_43300_n366) );
  OR2X2 OR2X2_1667 ( .A(u0_u0__abc_43300_n350_bF_buf0), .B(\wb_data_i[4] ), .Y(u0_u0__abc_43300_n367) );
  OR2X2 OR2X2_1668 ( .A(u0_u0_init_req_we_FF_INPUT_bF_buf3), .B(u0_csc0_5_), .Y(u0_u0__abc_43300_n370) );
  OR2X2 OR2X2_1669 ( .A(u0_u0__abc_43300_n350_bF_buf4), .B(\wb_data_i[5] ), .Y(u0_u0__abc_43300_n371) );
  OR2X2 OR2X2_167 ( .A(u0__abc_49347_n1203_bF_buf2), .B(u0_tms0_3_), .Y(u0__abc_49347_n1276) );
  OR2X2 OR2X2_1670 ( .A(u0_u0_init_req_we_FF_INPUT_bF_buf2), .B(u0_csc0_6_), .Y(u0_u0__abc_43300_n374) );
  OR2X2 OR2X2_1671 ( .A(u0_u0__abc_43300_n350_bF_buf3), .B(\wb_data_i[6] ), .Y(u0_u0__abc_43300_n375) );
  OR2X2 OR2X2_1672 ( .A(u0_u0_init_req_we_FF_INPUT_bF_buf1), .B(u0_csc0_7_), .Y(u0_u0__abc_43300_n378) );
  OR2X2 OR2X2_1673 ( .A(u0_u0__abc_43300_n350_bF_buf2), .B(\wb_data_i[7] ), .Y(u0_u0__abc_43300_n379) );
  OR2X2 OR2X2_1674 ( .A(u0_u0_init_req_we_FF_INPUT_bF_buf0), .B(u0_csc0_8_), .Y(u0_u0__abc_43300_n382) );
  OR2X2 OR2X2_1675 ( .A(u0_u0__abc_43300_n350_bF_buf1), .B(\wb_data_i[8] ), .Y(u0_u0__abc_43300_n383) );
  OR2X2 OR2X2_1676 ( .A(u0_u0_init_req_we_FF_INPUT_bF_buf4), .B(u0_csc0_9_), .Y(u0_u0__abc_43300_n386) );
  OR2X2 OR2X2_1677 ( .A(u0_u0__abc_43300_n350_bF_buf0), .B(\wb_data_i[9] ), .Y(u0_u0__abc_43300_n387) );
  OR2X2 OR2X2_1678 ( .A(u0_u0_init_req_we_FF_INPUT_bF_buf3), .B(u0_csc0_10_), .Y(u0_u0__abc_43300_n390) );
  OR2X2 OR2X2_1679 ( .A(u0_u0__abc_43300_n350_bF_buf4), .B(\wb_data_i[10] ), .Y(u0_u0__abc_43300_n391) );
  OR2X2 OR2X2_168 ( .A(u0__abc_49347_n1278), .B(u0__abc_49347_n1256), .Y(u0_sp_tms_3__FF_INPUT) );
  OR2X2 OR2X2_1680 ( .A(u0_u0_init_req_we_FF_INPUT_bF_buf2), .B(u0_csc0_11_), .Y(u0_u0__abc_43300_n394) );
  OR2X2 OR2X2_1681 ( .A(u0_u0__abc_43300_n350_bF_buf3), .B(\wb_data_i[11] ), .Y(u0_u0__abc_43300_n395) );
  OR2X2 OR2X2_1682 ( .A(u0_u0_init_req_we_FF_INPUT_bF_buf1), .B(u0_csc0_12_), .Y(u0_u0__abc_43300_n398) );
  OR2X2 OR2X2_1683 ( .A(u0_u0__abc_43300_n350_bF_buf2), .B(\wb_data_i[12] ), .Y(u0_u0__abc_43300_n399) );
  OR2X2 OR2X2_1684 ( .A(u0_u0_init_req_we_FF_INPUT_bF_buf0), .B(u0_csc0_13_), .Y(u0_u0__abc_43300_n402) );
  OR2X2 OR2X2_1685 ( .A(u0_u0__abc_43300_n350_bF_buf1), .B(\wb_data_i[13] ), .Y(u0_u0__abc_43300_n403) );
  OR2X2 OR2X2_1686 ( .A(u0_u0_init_req_we_FF_INPUT_bF_buf4), .B(u0_csc0_14_), .Y(u0_u0__abc_43300_n406) );
  OR2X2 OR2X2_1687 ( .A(u0_u0__abc_43300_n350_bF_buf0), .B(\wb_data_i[14] ), .Y(u0_u0__abc_43300_n407) );
  OR2X2 OR2X2_1688 ( .A(u0_u0_init_req_we_FF_INPUT_bF_buf3), .B(u0_csc0_15_), .Y(u0_u0__abc_43300_n410) );
  OR2X2 OR2X2_1689 ( .A(u0_u0__abc_43300_n350_bF_buf4), .B(\wb_data_i[15] ), .Y(u0_u0__abc_43300_n411) );
  OR2X2 OR2X2_169 ( .A(u0__abc_49347_n1183_1_bF_buf1), .B(1'b0), .Y(u0__abc_49347_n1282_1) );
  OR2X2 OR2X2_1690 ( .A(u0_u0_init_req_we_FF_INPUT_bF_buf2), .B(u0_csc0_16_), .Y(u0_u0__abc_43300_n414) );
  OR2X2 OR2X2_1691 ( .A(u0_u0__abc_43300_n350_bF_buf3), .B(\wb_data_i[16] ), .Y(u0_u0__abc_43300_n415) );
  OR2X2 OR2X2_1692 ( .A(u0_u0_init_req_we_FF_INPUT_bF_buf1), .B(u0_csc0_17_), .Y(u0_u0__abc_43300_n418) );
  OR2X2 OR2X2_1693 ( .A(u0_u0__abc_43300_n350_bF_buf2), .B(\wb_data_i[17] ), .Y(u0_u0__abc_43300_n419) );
  OR2X2 OR2X2_1694 ( .A(u0_u0_init_req_we_FF_INPUT_bF_buf0), .B(u0_csc0_18_), .Y(u0_u0__abc_43300_n422) );
  OR2X2 OR2X2_1695 ( .A(u0_u0__abc_43300_n350_bF_buf1), .B(\wb_data_i[18] ), .Y(u0_u0__abc_43300_n423) );
  OR2X2 OR2X2_1696 ( .A(u0_u0_init_req_we_FF_INPUT_bF_buf4), .B(u0_csc0_19_), .Y(u0_u0__abc_43300_n426) );
  OR2X2 OR2X2_1697 ( .A(u0_u0__abc_43300_n350_bF_buf0), .B(\wb_data_i[19] ), .Y(u0_u0__abc_43300_n427) );
  OR2X2 OR2X2_1698 ( .A(u0_u0_init_req_we_FF_INPUT_bF_buf3), .B(u0_csc0_20_), .Y(u0_u0__abc_43300_n430) );
  OR2X2 OR2X2_1699 ( .A(u0_u0__abc_43300_n350_bF_buf4), .B(\wb_data_i[20] ), .Y(u0_u0__abc_43300_n431) );
  OR2X2 OR2X2_17 ( .A(_abc_55805_n262), .B(_abc_55805_n237_1), .Y(_abc_55805_n263) );
  OR2X2 OR2X2_170 ( .A(spec_req_cs_6_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n1283) );
  OR2X2 OR2X2_1700 ( .A(u0_u0_init_req_we_FF_INPUT_bF_buf2), .B(u0_csc0_21_), .Y(u0_u0__abc_43300_n434) );
  OR2X2 OR2X2_1701 ( .A(u0_u0__abc_43300_n350_bF_buf3), .B(\wb_data_i[21] ), .Y(u0_u0__abc_43300_n435) );
  OR2X2 OR2X2_1702 ( .A(u0_u0_init_req_we_FF_INPUT_bF_buf1), .B(u0_csc0_22_), .Y(u0_u0__abc_43300_n438) );
  OR2X2 OR2X2_1703 ( .A(u0_u0__abc_43300_n350_bF_buf2), .B(\wb_data_i[22] ), .Y(u0_u0__abc_43300_n439) );
  OR2X2 OR2X2_1704 ( .A(u0_u0_init_req_we_FF_INPUT_bF_buf0), .B(u0_csc0_23_), .Y(u0_u0__abc_43300_n442) );
  OR2X2 OR2X2_1705 ( .A(u0_u0__abc_43300_n350_bF_buf1), .B(\wb_data_i[23] ), .Y(u0_u0__abc_43300_n443) );
  OR2X2 OR2X2_1706 ( .A(u0_u0_init_req_we_FF_INPUT_bF_buf4), .B(u0_csc0_24_), .Y(u0_u0__abc_43300_n446) );
  OR2X2 OR2X2_1707 ( .A(u0_u0__abc_43300_n350_bF_buf0), .B(\wb_data_i[24] ), .Y(u0_u0__abc_43300_n447) );
  OR2X2 OR2X2_1708 ( .A(u0_u0_init_req_we_FF_INPUT_bF_buf3), .B(u0_csc0_25_), .Y(u0_u0__abc_43300_n450) );
  OR2X2 OR2X2_1709 ( .A(u0_u0__abc_43300_n350_bF_buf4), .B(\wb_data_i[25] ), .Y(u0_u0__abc_43300_n451) );
  OR2X2 OR2X2_171 ( .A(u0__abc_49347_n1285), .B(u0__abc_49347_n1281_1), .Y(u0__abc_49347_n1286) );
  OR2X2 OR2X2_1710 ( .A(u0_u0_init_req_we_FF_INPUT_bF_buf2), .B(u0_csc0_26_), .Y(u0_u0__abc_43300_n454) );
  OR2X2 OR2X2_1711 ( .A(u0_u0__abc_43300_n350_bF_buf3), .B(\wb_data_i[26] ), .Y(u0_u0__abc_43300_n455) );
  OR2X2 OR2X2_1712 ( .A(u0_u0_init_req_we_FF_INPUT_bF_buf1), .B(u0_csc0_27_), .Y(u0_u0__abc_43300_n458) );
  OR2X2 OR2X2_1713 ( .A(u0_u0__abc_43300_n350_bF_buf2), .B(\wb_data_i[27] ), .Y(u0_u0__abc_43300_n459) );
  OR2X2 OR2X2_1714 ( .A(u0_u0_init_req_we_FF_INPUT_bF_buf0), .B(u0_csc0_28_), .Y(u0_u0__abc_43300_n462) );
  OR2X2 OR2X2_1715 ( .A(u0_u0__abc_43300_n350_bF_buf1), .B(\wb_data_i[28] ), .Y(u0_u0__abc_43300_n463) );
  OR2X2 OR2X2_1716 ( .A(u0_u0_init_req_we_FF_INPUT_bF_buf4), .B(u0_csc0_29_), .Y(u0_u0__abc_43300_n466) );
  OR2X2 OR2X2_1717 ( .A(u0_u0__abc_43300_n350_bF_buf0), .B(\wb_data_i[29] ), .Y(u0_u0__abc_43300_n467) );
  OR2X2 OR2X2_1718 ( .A(u0_u0_init_req_we_FF_INPUT_bF_buf3), .B(u0_csc0_30_), .Y(u0_u0__abc_43300_n470) );
  OR2X2 OR2X2_1719 ( .A(u0_u0__abc_43300_n350_bF_buf4), .B(\wb_data_i[30] ), .Y(u0_u0__abc_43300_n471) );
  OR2X2 OR2X2_172 ( .A(u0__abc_49347_n1287), .B(u0__abc_49347_n1288), .Y(u0__abc_49347_n1289) );
  OR2X2 OR2X2_1720 ( .A(u0_u0_init_req_we_FF_INPUT_bF_buf2), .B(u0_csc0_31_), .Y(u0_u0__abc_43300_n474) );
  OR2X2 OR2X2_1721 ( .A(u0_u0__abc_43300_n350_bF_buf3), .B(\wb_data_i[31] ), .Y(u0_u0__abc_43300_n475) );
  OR2X2 OR2X2_1722 ( .A(u0_u0__abc_43300_n481), .B(u0_u0__abc_43300_n479), .Y(u0_u0__abc_43300_n482) );
  OR2X2 OR2X2_1723 ( .A(u0_u0__abc_43300_n485), .B(u0_u0__abc_43300_n483), .Y(u0_u0__abc_43300_n486) );
  OR2X2 OR2X2_1724 ( .A(u0_u0__abc_43300_n492), .B(u0_u0__abc_43300_n484), .Y(u0_u0__abc_43300_n493) );
  OR2X2 OR2X2_1725 ( .A(u0_u0__abc_43300_n498), .B(u0_u0__abc_43300_n496), .Y(u0_u0__abc_43300_n499) );
  OR2X2 OR2X2_1726 ( .A(u0_u0__abc_43300_n502), .B(u0_u0__abc_43300_n500), .Y(u0_u0__abc_43300_n503) );
  OR2X2 OR2X2_1727 ( .A(u0_u0__abc_43300_n508), .B(u0_u0__abc_43300_n501), .Y(u0_u0__abc_43300_n509) );
  OR2X2 OR2X2_1728 ( .A(u0_u0__abc_43300_n516), .B(u0_u0__abc_43300_n517), .Y(u0_u0__abc_43300_n518) );
  OR2X2 OR2X2_1729 ( .A(u0_u0__abc_43300_n520), .B(u0_u0__abc_43300_n515), .Y(u0_u0__abc_43300_n521) );
  OR2X2 OR2X2_173 ( .A(u0__abc_49347_n1290_1), .B(u0__abc_49347_n1291_1), .Y(u0__abc_49347_n1292) );
  OR2X2 OR2X2_1730 ( .A(u0_u0__abc_43300_n525), .B(u0_u0__abc_43300_n489), .Y(u0_u0__abc_43300_n526) );
  OR2X2 OR2X2_1731 ( .A(u0_u0__abc_43300_n529), .B(u0_u0__abc_43300_n527), .Y(u0_u0__abc_43300_n530) );
  OR2X2 OR2X2_1732 ( .A(u0_u0__abc_43300_n534), .B(u0_u0__abc_43300_n532), .Y(u0_u0__abc_43300_n535) );
  OR2X2 OR2X2_1733 ( .A(u0_u0__abc_43300_n536), .B(u0_u0__abc_43300_n528), .Y(u0_u0__abc_43300_n537) );
  OR2X2 OR2X2_1734 ( .A(u0_u0__abc_43300_n540), .B(u0_u0__abc_43300_n533), .Y(u0_u0__abc_43300_n541) );
  OR2X2 OR2X2_1735 ( .A(u0_u0_inited), .B(u0_init_ack0), .Y(u0_u0_inited_FF_INPUT) );
  OR2X2 OR2X2_1736 ( .A(u0_u0__abc_43300_n554), .B(u0_u0__abc_43300_n550), .Y(u0_u0_init_req_FF_INPUT) );
  OR2X2 OR2X2_1737 ( .A(u0_csc1_2_), .B(u0_csc1_1_), .Y(u0_u1__abc_43657_n201_1) );
  OR2X2 OR2X2_1738 ( .A(u0_u1__abc_43657_n201_1), .B(u0_csc1_3_), .Y(u0_u1__abc_43657_n202) );
  OR2X2 OR2X2_1739 ( .A(u0_u1__abc_43657_n209_1), .B(u0_u1__abc_43657_n205), .Y(u0_u1_lmr_req_FF_INPUT) );
  OR2X2 OR2X2_174 ( .A(u0__abc_49347_n1293), .B(u0__abc_49347_n1294), .Y(u0__abc_49347_n1295) );
  OR2X2 OR2X2_1740 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf7), .B(u0_tms1_0_), .Y(u0_u1__abc_43657_n218_1) );
  OR2X2 OR2X2_1741 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf5), .B(u0_tms1_1_), .Y(u0_u1__abc_43657_n225_1) );
  OR2X2 OR2X2_1742 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf3), .B(u0_tms1_2_), .Y(u0_u1__abc_43657_n231_1) );
  OR2X2 OR2X2_1743 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf1), .B(u0_tms1_3_), .Y(u0_u1__abc_43657_n237_1) );
  OR2X2 OR2X2_1744 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf7), .B(u0_tms1_4_), .Y(u0_u1__abc_43657_n243_1) );
  OR2X2 OR2X2_1745 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf5), .B(u0_tms1_5_), .Y(u0_u1__abc_43657_n249_1) );
  OR2X2 OR2X2_1746 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf3), .B(u0_tms1_6_), .Y(u0_u1__abc_43657_n255) );
  OR2X2 OR2X2_1747 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf1), .B(u0_tms1_7_), .Y(u0_u1__abc_43657_n261_1) );
  OR2X2 OR2X2_1748 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf7), .B(u0_tms1_8_), .Y(u0_u1__abc_43657_n267_1) );
  OR2X2 OR2X2_1749 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf5), .B(u0_tms1_9_), .Y(u0_u1__abc_43657_n273) );
  OR2X2 OR2X2_175 ( .A(u0__abc_49347_n1297), .B(spec_req_cs_0_bF_buf4), .Y(u0__abc_49347_n1298) );
  OR2X2 OR2X2_1750 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf3), .B(u0_tms1_10_), .Y(u0_u1__abc_43657_n279) );
  OR2X2 OR2X2_1751 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf1), .B(u0_tms1_11_), .Y(u0_u1__abc_43657_n285) );
  OR2X2 OR2X2_1752 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf7), .B(u0_tms1_12_), .Y(u0_u1__abc_43657_n291) );
  OR2X2 OR2X2_1753 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf5), .B(u0_tms1_13_), .Y(u0_u1__abc_43657_n297_1) );
  OR2X2 OR2X2_1754 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf3), .B(u0_tms1_14_), .Y(u0_u1__abc_43657_n303) );
  OR2X2 OR2X2_1755 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf1), .B(u0_tms1_15_), .Y(u0_u1__abc_43657_n309_1) );
  OR2X2 OR2X2_1756 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf7), .B(u0_tms1_16_), .Y(u0_u1__abc_43657_n315_1) );
  OR2X2 OR2X2_1757 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf5), .B(u0_tms1_17_), .Y(u0_u1__abc_43657_n321) );
  OR2X2 OR2X2_1758 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf3), .B(u0_tms1_18_), .Y(u0_u1__abc_43657_n327) );
  OR2X2 OR2X2_1759 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf1), .B(u0_tms1_19_), .Y(u0_u1__abc_43657_n333) );
  OR2X2 OR2X2_176 ( .A(u0__abc_49347_n1296), .B(u0__abc_49347_n1298), .Y(u0__abc_49347_n1299_1) );
  OR2X2 OR2X2_1760 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf7), .B(u0_tms1_20_), .Y(u0_u1__abc_43657_n339) );
  OR2X2 OR2X2_1761 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf5), .B(u0_tms1_21_), .Y(u0_u1__abc_43657_n345) );
  OR2X2 OR2X2_1762 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf3), .B(u0_tms1_22_), .Y(u0_u1__abc_43657_n351) );
  OR2X2 OR2X2_1763 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf1), .B(u0_tms1_23_), .Y(u0_u1__abc_43657_n357) );
  OR2X2 OR2X2_1764 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf7), .B(u0_tms1_24_), .Y(u0_u1__abc_43657_n363) );
  OR2X2 OR2X2_1765 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf5), .B(u0_tms1_25_), .Y(u0_u1__abc_43657_n369) );
  OR2X2 OR2X2_1766 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf3), .B(u0_tms1_26_), .Y(u0_u1__abc_43657_n375) );
  OR2X2 OR2X2_1767 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf1), .B(u0_tms1_27_), .Y(u0_u1__abc_43657_n381) );
  OR2X2 OR2X2_1768 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf7), .B(u0_tms1_28_), .Y(u0_u1__abc_43657_n387) );
  OR2X2 OR2X2_1769 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf5), .B(u0_tms1_29_), .Y(u0_u1__abc_43657_n393) );
  OR2X2 OR2X2_177 ( .A(u0__abc_49347_n1203_bF_buf1), .B(u0_tms0_4_), .Y(u0__abc_49347_n1300_1) );
  OR2X2 OR2X2_1770 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf3), .B(u0_tms1_30_), .Y(u0_u1__abc_43657_n399) );
  OR2X2 OR2X2_1771 ( .A(u0_u1_lmr_req_we_FF_INPUT_bF_buf1), .B(u0_tms1_31_), .Y(u0_u1__abc_43657_n405) );
  OR2X2 OR2X2_1772 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf7), .B(u0_csc1_0_), .Y(u0_u1__abc_43657_n413) );
  OR2X2 OR2X2_1773 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf5), .B(u0_csc1_1_), .Y(u0_u1__abc_43657_n418) );
  OR2X2 OR2X2_1774 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf3), .B(u0_csc1_2_), .Y(u0_u1__abc_43657_n423) );
  OR2X2 OR2X2_1775 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf1), .B(u0_csc1_3_), .Y(u0_u1__abc_43657_n428) );
  OR2X2 OR2X2_1776 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf7), .B(u0_csc1_4_), .Y(u0_u1__abc_43657_n433) );
  OR2X2 OR2X2_1777 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf5), .B(u0_csc1_5_), .Y(u0_u1__abc_43657_n438) );
  OR2X2 OR2X2_1778 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf3), .B(u0_csc1_6_), .Y(u0_u1__abc_43657_n443) );
  OR2X2 OR2X2_1779 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf1), .B(u0_csc1_7_), .Y(u0_u1__abc_43657_n448) );
  OR2X2 OR2X2_178 ( .A(u0__abc_49347_n1302), .B(u0__abc_49347_n1280), .Y(u0_sp_tms_4__FF_INPUT) );
  OR2X2 OR2X2_1780 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf7), .B(u0_csc1_8_), .Y(u0_u1__abc_43657_n453) );
  OR2X2 OR2X2_1781 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf5), .B(u0_csc1_9_), .Y(u0_u1__abc_43657_n458) );
  OR2X2 OR2X2_1782 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf3), .B(u0_csc1_10_), .Y(u0_u1__abc_43657_n463) );
  OR2X2 OR2X2_1783 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf1), .B(u0_csc1_11_), .Y(u0_u1__abc_43657_n468) );
  OR2X2 OR2X2_1784 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf7), .B(u0_csc1_12_), .Y(u0_u1__abc_43657_n473) );
  OR2X2 OR2X2_1785 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf5), .B(u0_csc1_13_), .Y(u0_u1__abc_43657_n478) );
  OR2X2 OR2X2_1786 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf3), .B(u0_csc1_14_), .Y(u0_u1__abc_43657_n483) );
  OR2X2 OR2X2_1787 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf1), .B(u0_csc1_15_), .Y(u0_u1__abc_43657_n488) );
  OR2X2 OR2X2_1788 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf7), .B(u0_csc1_16_), .Y(u0_u1__abc_43657_n493) );
  OR2X2 OR2X2_1789 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf5), .B(u0_csc1_17_), .Y(u0_u1__abc_43657_n498) );
  OR2X2 OR2X2_179 ( .A(u0__abc_49347_n1183_1_bF_buf0), .B(1'b0), .Y(u0__abc_49347_n1306) );
  OR2X2 OR2X2_1790 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf3), .B(u0_csc1_18_), .Y(u0_u1__abc_43657_n503) );
  OR2X2 OR2X2_1791 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf1), .B(u0_csc1_19_), .Y(u0_u1__abc_43657_n508) );
  OR2X2 OR2X2_1792 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf7), .B(u0_csc1_20_), .Y(u0_u1__abc_43657_n513) );
  OR2X2 OR2X2_1793 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf5), .B(u0_csc1_21_), .Y(u0_u1__abc_43657_n518) );
  OR2X2 OR2X2_1794 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf3), .B(u0_csc1_22_), .Y(u0_u1__abc_43657_n523) );
  OR2X2 OR2X2_1795 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf1), .B(u0_csc1_23_), .Y(u0_u1__abc_43657_n528) );
  OR2X2 OR2X2_1796 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf7), .B(u0_csc1_24_), .Y(u0_u1__abc_43657_n533) );
  OR2X2 OR2X2_1797 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf5), .B(u0_csc1_25_), .Y(u0_u1__abc_43657_n538) );
  OR2X2 OR2X2_1798 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf3), .B(u0_csc1_26_), .Y(u0_u1__abc_43657_n543) );
  OR2X2 OR2X2_1799 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf1), .B(u0_csc1_27_), .Y(u0_u1__abc_43657_n548) );
  OR2X2 OR2X2_18 ( .A(_abc_55805_n245_1), .B(cs_need_rfr_3_), .Y(_abc_55805_n264) );
  OR2X2 OR2X2_180 ( .A(spec_req_cs_6_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n1307) );
  OR2X2 OR2X2_1800 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf7), .B(u0_csc1_28_), .Y(u0_u1__abc_43657_n553) );
  OR2X2 OR2X2_1801 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf5), .B(u0_csc1_29_), .Y(u0_u1__abc_43657_n558) );
  OR2X2 OR2X2_1802 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf3), .B(u0_csc1_30_), .Y(u0_u1__abc_43657_n563) );
  OR2X2 OR2X2_1803 ( .A(u0_u1_init_req_we_FF_INPUT_bF_buf1), .B(u0_csc1_31_), .Y(u0_u1__abc_43657_n568) );
  OR2X2 OR2X2_1804 ( .A(u0_u1__abc_43657_n576), .B(u0_u1__abc_43657_n574), .Y(u0_u1__abc_43657_n577) );
  OR2X2 OR2X2_1805 ( .A(u0_u1__abc_43657_n580), .B(u0_u1__abc_43657_n578), .Y(u0_u1__abc_43657_n581) );
  OR2X2 OR2X2_1806 ( .A(u0_u1__abc_43657_n587), .B(u0_u1__abc_43657_n579), .Y(u0_u1__abc_43657_n588) );
  OR2X2 OR2X2_1807 ( .A(u0_u1__abc_43657_n593), .B(u0_u1__abc_43657_n591), .Y(u0_u1__abc_43657_n594) );
  OR2X2 OR2X2_1808 ( .A(u0_u1__abc_43657_n597), .B(u0_u1__abc_43657_n595), .Y(u0_u1__abc_43657_n598) );
  OR2X2 OR2X2_1809 ( .A(u0_u1__abc_43657_n603), .B(u0_u1__abc_43657_n596), .Y(u0_u1__abc_43657_n604) );
  OR2X2 OR2X2_181 ( .A(u0__abc_49347_n1309_1), .B(u0__abc_49347_n1305), .Y(u0__abc_49347_n1310) );
  OR2X2 OR2X2_1810 ( .A(u0_u1__abc_43657_n611), .B(u0_u1__abc_43657_n612), .Y(u0_u1__abc_43657_n613) );
  OR2X2 OR2X2_1811 ( .A(u0_u1__abc_43657_n615), .B(u0_u1__abc_43657_n610), .Y(u0_u1__abc_43657_n616) );
  OR2X2 OR2X2_1812 ( .A(u0_u1__abc_43657_n620), .B(u0_u1__abc_43657_n584), .Y(u0_u1__abc_43657_n621) );
  OR2X2 OR2X2_1813 ( .A(u0_u1__abc_43657_n624), .B(u0_u1__abc_43657_n622), .Y(u0_u1__abc_43657_n625) );
  OR2X2 OR2X2_1814 ( .A(u0_u1__abc_43657_n629), .B(u0_u1__abc_43657_n627), .Y(u0_u1__abc_43657_n630) );
  OR2X2 OR2X2_1815 ( .A(u0_u1__abc_43657_n631), .B(u0_u1__abc_43657_n623), .Y(u0_u1__abc_43657_n632) );
  OR2X2 OR2X2_1816 ( .A(u0_u1__abc_43657_n635), .B(u0_u1__abc_43657_n628), .Y(u0_u1__abc_43657_n636) );
  OR2X2 OR2X2_1817 ( .A(u0_u1_inited), .B(u0_init_ack1), .Y(u0_u1_inited_FF_INPUT) );
  OR2X2 OR2X2_1818 ( .A(u0_u1__abc_43657_n649), .B(u0_u1__abc_43657_n645), .Y(u0_u1_init_req_FF_INPUT) );
  OR2X2 OR2X2_1819 ( .A(u0_u2_addr_r_4_), .B(u0_u2_addr_r_3_), .Y(u0_u2__abc_44109_n203) );
  OR2X2 OR2X2_182 ( .A(u0__abc_49347_n1311), .B(u0__abc_49347_n1312), .Y(u0__abc_49347_n1313) );
  OR2X2 OR2X2_1820 ( .A(u0_u2__abc_44109_n203), .B(u0_u2_addr_r_6_), .Y(u0_u2__abc_44109_n204_1) );
  OR2X2 OR2X2_1821 ( .A(u0_u2_init_req_we_FF_INPUT_bF_buf4), .B(u0_csc2_0_), .Y(u0_u2__abc_44109_n208_1) );
  OR2X2 OR2X2_1822 ( .A(u0_u2__abc_44109_n210_1_bF_buf4), .B(\wb_data_i[0] ), .Y(u0_u2__abc_44109_n211_1) );
  OR2X2 OR2X2_1823 ( .A(u0_u2_init_req_we_FF_INPUT_bF_buf2), .B(u0_csc2_1_), .Y(u0_u2__abc_44109_n214_1) );
  OR2X2 OR2X2_1824 ( .A(u0_u2__abc_44109_n210_1_bF_buf3), .B(\wb_data_i[1] ), .Y(u0_u2__abc_44109_n215) );
  OR2X2 OR2X2_1825 ( .A(u0_u2_init_req_we_FF_INPUT_bF_buf1), .B(u0_csc2_2_), .Y(u0_u2__abc_44109_n218) );
  OR2X2 OR2X2_1826 ( .A(u0_u2__abc_44109_n210_1_bF_buf2), .B(\wb_data_i[2] ), .Y(u0_u2__abc_44109_n219_1) );
  OR2X2 OR2X2_1827 ( .A(u0_u2_init_req_we_FF_INPUT_bF_buf0), .B(u0_csc2_3_), .Y(u0_u2__abc_44109_n222_1) );
  OR2X2 OR2X2_1828 ( .A(u0_u2__abc_44109_n210_1_bF_buf1), .B(\wb_data_i[3] ), .Y(u0_u2__abc_44109_n223_1) );
  OR2X2 OR2X2_1829 ( .A(u0_u2_init_req_we_FF_INPUT_bF_buf4), .B(u0_csc2_4_), .Y(u0_u2__abc_44109_n226_1) );
  OR2X2 OR2X2_183 ( .A(u0__abc_49347_n1314), .B(u0__abc_49347_n1315), .Y(u0__abc_49347_n1316) );
  OR2X2 OR2X2_1830 ( .A(u0_u2__abc_44109_n210_1_bF_buf0), .B(\wb_data_i[4] ), .Y(u0_u2__abc_44109_n227) );
  OR2X2 OR2X2_1831 ( .A(u0_u2_init_req_we_FF_INPUT_bF_buf3), .B(u0_csc2_5_), .Y(u0_u2__abc_44109_n230) );
  OR2X2 OR2X2_1832 ( .A(u0_u2__abc_44109_n210_1_bF_buf4), .B(\wb_data_i[5] ), .Y(u0_u2__abc_44109_n231_1) );
  OR2X2 OR2X2_1833 ( .A(u0_u2_init_req_we_FF_INPUT_bF_buf2), .B(u0_csc2_6_), .Y(u0_u2__abc_44109_n234_1) );
  OR2X2 OR2X2_1834 ( .A(u0_u2__abc_44109_n210_1_bF_buf3), .B(\wb_data_i[6] ), .Y(u0_u2__abc_44109_n235_1) );
  OR2X2 OR2X2_1835 ( .A(u0_u2_init_req_we_FF_INPUT_bF_buf1), .B(u0_csc2_7_), .Y(u0_u2__abc_44109_n238_1) );
  OR2X2 OR2X2_1836 ( .A(u0_u2__abc_44109_n210_1_bF_buf2), .B(\wb_data_i[7] ), .Y(u0_u2__abc_44109_n239) );
  OR2X2 OR2X2_1837 ( .A(u0_u2_init_req_we_FF_INPUT_bF_buf0), .B(u0_csc2_8_), .Y(u0_u2__abc_44109_n242) );
  OR2X2 OR2X2_1838 ( .A(u0_u2__abc_44109_n210_1_bF_buf1), .B(\wb_data_i[8] ), .Y(u0_u2__abc_44109_n243) );
  OR2X2 OR2X2_1839 ( .A(u0_u2_init_req_we_FF_INPUT_bF_buf4), .B(u0_csc2_9_), .Y(u0_u2__abc_44109_n246_1) );
  OR2X2 OR2X2_184 ( .A(u0__abc_49347_n1317_1), .B(u0__abc_49347_n1318_1), .Y(u0__abc_49347_n1319) );
  OR2X2 OR2X2_1840 ( .A(u0_u2__abc_44109_n210_1_bF_buf0), .B(\wb_data_i[9] ), .Y(u0_u2__abc_44109_n247) );
  OR2X2 OR2X2_1841 ( .A(u0_u2_init_req_we_FF_INPUT_bF_buf3), .B(u0_csc2_10_), .Y(u0_u2__abc_44109_n250_1) );
  OR2X2 OR2X2_1842 ( .A(u0_u2__abc_44109_n210_1_bF_buf4), .B(\wb_data_i[10] ), .Y(u0_u2__abc_44109_n251_1) );
  OR2X2 OR2X2_1843 ( .A(u0_u2_init_req_we_FF_INPUT_bF_buf2), .B(u0_csc2_11_), .Y(u0_u2__abc_44109_n254) );
  OR2X2 OR2X2_1844 ( .A(u0_u2__abc_44109_n210_1_bF_buf3), .B(\wb_data_i[11] ), .Y(u0_u2__abc_44109_n255) );
  OR2X2 OR2X2_1845 ( .A(u0_u2_init_req_we_FF_INPUT_bF_buf1), .B(u0_csc2_12_), .Y(u0_u2__abc_44109_n258_1) );
  OR2X2 OR2X2_1846 ( .A(u0_u2__abc_44109_n210_1_bF_buf2), .B(\wb_data_i[12] ), .Y(u0_u2__abc_44109_n259_1) );
  OR2X2 OR2X2_1847 ( .A(u0_u2_init_req_we_FF_INPUT_bF_buf0), .B(u0_csc2_13_), .Y(u0_u2__abc_44109_n262) );
  OR2X2 OR2X2_1848 ( .A(u0_u2__abc_44109_n210_1_bF_buf1), .B(\wb_data_i[13] ), .Y(u0_u2__abc_44109_n263_1) );
  OR2X2 OR2X2_1849 ( .A(u0_u2_init_req_we_FF_INPUT_bF_buf4), .B(u0_csc2_14_), .Y(u0_u2__abc_44109_n266) );
  OR2X2 OR2X2_185 ( .A(u0__abc_49347_n1321), .B(spec_req_cs_0_bF_buf3), .Y(u0__abc_49347_n1322) );
  OR2X2 OR2X2_1850 ( .A(u0_u2__abc_44109_n210_1_bF_buf0), .B(\wb_data_i[14] ), .Y(u0_u2__abc_44109_n267) );
  OR2X2 OR2X2_1851 ( .A(u0_u2_init_req_we_FF_INPUT_bF_buf3), .B(u0_csc2_15_), .Y(u0_u2__abc_44109_n270_1) );
  OR2X2 OR2X2_1852 ( .A(u0_u2__abc_44109_n210_1_bF_buf4), .B(\wb_data_i[15] ), .Y(u0_u2__abc_44109_n271) );
  OR2X2 OR2X2_1853 ( .A(u0_u2_init_req_we_FF_INPUT_bF_buf2), .B(u0_csc2_16_), .Y(u0_u2__abc_44109_n274_1) );
  OR2X2 OR2X2_1854 ( .A(u0_u2__abc_44109_n210_1_bF_buf3), .B(\wb_data_i[16] ), .Y(u0_u2__abc_44109_n275) );
  OR2X2 OR2X2_1855 ( .A(u0_u2_init_req_we_FF_INPUT_bF_buf1), .B(u0_csc2_17_), .Y(u0_u2__abc_44109_n278) );
  OR2X2 OR2X2_1856 ( .A(u0_u2__abc_44109_n210_1_bF_buf2), .B(\wb_data_i[17] ), .Y(u0_u2__abc_44109_n279) );
  OR2X2 OR2X2_1857 ( .A(u0_u2_init_req_we_FF_INPUT_bF_buf0), .B(u0_csc2_18_), .Y(u0_u2__abc_44109_n282) );
  OR2X2 OR2X2_1858 ( .A(u0_u2__abc_44109_n210_1_bF_buf1), .B(\wb_data_i[18] ), .Y(u0_u2__abc_44109_n283_1) );
  OR2X2 OR2X2_1859 ( .A(u0_u2_init_req_we_FF_INPUT_bF_buf4), .B(u0_csc2_19_), .Y(u0_u2__abc_44109_n286) );
  OR2X2 OR2X2_186 ( .A(u0__abc_49347_n1320), .B(u0__abc_49347_n1322), .Y(u0__abc_49347_n1323) );
  OR2X2 OR2X2_1860 ( .A(u0_u2__abc_44109_n210_1_bF_buf0), .B(\wb_data_i[19] ), .Y(u0_u2__abc_44109_n287_1) );
  OR2X2 OR2X2_1861 ( .A(u0_u2_init_req_we_FF_INPUT_bF_buf3), .B(u0_csc2_20_), .Y(u0_u2__abc_44109_n290) );
  OR2X2 OR2X2_1862 ( .A(u0_u2__abc_44109_n210_1_bF_buf4), .B(\wb_data_i[20] ), .Y(u0_u2__abc_44109_n291_1) );
  OR2X2 OR2X2_1863 ( .A(u0_u2_init_req_we_FF_INPUT_bF_buf2), .B(u0_csc2_21_), .Y(u0_u2__abc_44109_n294) );
  OR2X2 OR2X2_1864 ( .A(u0_u2__abc_44109_n210_1_bF_buf3), .B(\wb_data_i[21] ), .Y(u0_u2__abc_44109_n295_1) );
  OR2X2 OR2X2_1865 ( .A(u0_u2_init_req_we_FF_INPUT_bF_buf1), .B(u0_csc2_22_), .Y(u0_u2__abc_44109_n298) );
  OR2X2 OR2X2_1866 ( .A(u0_u2__abc_44109_n210_1_bF_buf2), .B(\wb_data_i[22] ), .Y(u0_u2__abc_44109_n299) );
  OR2X2 OR2X2_1867 ( .A(u0_u2_init_req_we_FF_INPUT_bF_buf0), .B(u0_csc2_23_), .Y(u0_u2__abc_44109_n302) );
  OR2X2 OR2X2_1868 ( .A(u0_u2__abc_44109_n210_1_bF_buf1), .B(\wb_data_i[23] ), .Y(u0_u2__abc_44109_n303) );
  OR2X2 OR2X2_1869 ( .A(u0_u2_init_req_we_FF_INPUT_bF_buf4), .B(u0_csc2_24_), .Y(u0_u2__abc_44109_n306_1) );
  OR2X2 OR2X2_187 ( .A(u0__abc_49347_n1203_bF_buf0), .B(u0_tms0_5_), .Y(u0__abc_49347_n1324) );
  OR2X2 OR2X2_1870 ( .A(u0_u2__abc_44109_n210_1_bF_buf0), .B(\wb_data_i[24] ), .Y(u0_u2__abc_44109_n307) );
  OR2X2 OR2X2_1871 ( .A(u0_u2_init_req_we_FF_INPUT_bF_buf3), .B(u0_csc2_25_), .Y(u0_u2__abc_44109_n310) );
  OR2X2 OR2X2_1872 ( .A(u0_u2__abc_44109_n210_1_bF_buf4), .B(\wb_data_i[25] ), .Y(u0_u2__abc_44109_n311) );
  OR2X2 OR2X2_1873 ( .A(u0_u2_init_req_we_FF_INPUT_bF_buf2), .B(u0_csc2_26_), .Y(u0_u2__abc_44109_n314) );
  OR2X2 OR2X2_1874 ( .A(u0_u2__abc_44109_n210_1_bF_buf3), .B(\wb_data_i[26] ), .Y(u0_u2__abc_44109_n315) );
  OR2X2 OR2X2_1875 ( .A(u0_u2_init_req_we_FF_INPUT_bF_buf1), .B(u0_csc2_27_), .Y(u0_u2__abc_44109_n318_1) );
  OR2X2 OR2X2_1876 ( .A(u0_u2__abc_44109_n210_1_bF_buf2), .B(\wb_data_i[27] ), .Y(u0_u2__abc_44109_n319) );
  OR2X2 OR2X2_1877 ( .A(u0_u2_init_req_we_FF_INPUT_bF_buf0), .B(u0_csc2_28_), .Y(u0_u2__abc_44109_n322_1) );
  OR2X2 OR2X2_1878 ( .A(u0_u2__abc_44109_n210_1_bF_buf1), .B(\wb_data_i[28] ), .Y(u0_u2__abc_44109_n323_1) );
  OR2X2 OR2X2_1879 ( .A(u0_u2_init_req_we_FF_INPUT_bF_buf4), .B(u0_csc2_29_), .Y(u0_u2__abc_44109_n326) );
  OR2X2 OR2X2_188 ( .A(u0__abc_49347_n1326_1), .B(u0__abc_49347_n1304), .Y(u0_sp_tms_5__FF_INPUT) );
  OR2X2 OR2X2_1880 ( .A(u0_u2__abc_44109_n210_1_bF_buf0), .B(\wb_data_i[29] ), .Y(u0_u2__abc_44109_n327) );
  OR2X2 OR2X2_1881 ( .A(u0_u2_init_req_we_FF_INPUT_bF_buf3), .B(u0_csc2_30_), .Y(u0_u2__abc_44109_n330) );
  OR2X2 OR2X2_1882 ( .A(u0_u2__abc_44109_n210_1_bF_buf4), .B(\wb_data_i[30] ), .Y(u0_u2__abc_44109_n331) );
  OR2X2 OR2X2_1883 ( .A(u0_u2_init_req_we_FF_INPUT_bF_buf2), .B(u0_csc2_31_), .Y(u0_u2__abc_44109_n334) );
  OR2X2 OR2X2_1884 ( .A(u0_u2__abc_44109_n210_1_bF_buf3), .B(\wb_data_i[31] ), .Y(u0_u2__abc_44109_n335) );
  OR2X2 OR2X2_1885 ( .A(u0_u2_lmr_req_we_FF_INPUT_bF_buf4), .B(u0_tms2_0_), .Y(u0_u2__abc_44109_n339) );
  OR2X2 OR2X2_1886 ( .A(u0_u2__abc_44109_n340_bF_buf4), .B(\wb_data_i[0] ), .Y(u0_u2__abc_44109_n341) );
  OR2X2 OR2X2_1887 ( .A(u0_u2_lmr_req_we_FF_INPUT_bF_buf2), .B(u0_tms2_1_), .Y(u0_u2__abc_44109_n344) );
  OR2X2 OR2X2_1888 ( .A(u0_u2__abc_44109_n340_bF_buf3), .B(\wb_data_i[1] ), .Y(u0_u2__abc_44109_n345) );
  OR2X2 OR2X2_1889 ( .A(u0_u2_lmr_req_we_FF_INPUT_bF_buf1), .B(u0_tms2_2_), .Y(u0_u2__abc_44109_n348) );
  OR2X2 OR2X2_189 ( .A(u0__abc_49347_n1183_1_bF_buf5), .B(1'b0), .Y(u0__abc_49347_n1330) );
  OR2X2 OR2X2_1890 ( .A(u0_u2__abc_44109_n340_bF_buf2), .B(\wb_data_i[2] ), .Y(u0_u2__abc_44109_n349) );
  OR2X2 OR2X2_1891 ( .A(u0_u2_lmr_req_we_FF_INPUT_bF_buf0), .B(u0_tms2_3_), .Y(u0_u2__abc_44109_n352) );
  OR2X2 OR2X2_1892 ( .A(u0_u2__abc_44109_n340_bF_buf1), .B(\wb_data_i[3] ), .Y(u0_u2__abc_44109_n353) );
  OR2X2 OR2X2_1893 ( .A(u0_u2_lmr_req_we_FF_INPUT_bF_buf4), .B(u0_tms2_4_), .Y(u0_u2__abc_44109_n356) );
  OR2X2 OR2X2_1894 ( .A(u0_u2__abc_44109_n340_bF_buf0), .B(\wb_data_i[4] ), .Y(u0_u2__abc_44109_n357) );
  OR2X2 OR2X2_1895 ( .A(u0_u2_lmr_req_we_FF_INPUT_bF_buf3), .B(u0_tms2_5_), .Y(u0_u2__abc_44109_n360) );
  OR2X2 OR2X2_1896 ( .A(u0_u2__abc_44109_n340_bF_buf4), .B(\wb_data_i[5] ), .Y(u0_u2__abc_44109_n361) );
  OR2X2 OR2X2_1897 ( .A(u0_u2_lmr_req_we_FF_INPUT_bF_buf2), .B(u0_tms2_6_), .Y(u0_u2__abc_44109_n364) );
  OR2X2 OR2X2_1898 ( .A(u0_u2__abc_44109_n340_bF_buf3), .B(\wb_data_i[6] ), .Y(u0_u2__abc_44109_n365) );
  OR2X2 OR2X2_1899 ( .A(u0_u2_lmr_req_we_FF_INPUT_bF_buf1), .B(u0_tms2_7_), .Y(u0_u2__abc_44109_n368) );
  OR2X2 OR2X2_19 ( .A(_abc_55805_n240_bF_buf1), .B(spec_req_cs_4_bF_buf5), .Y(_abc_55805_n266) );
  OR2X2 OR2X2_190 ( .A(spec_req_cs_6_bF_buf2), .B(1'b0), .Y(u0__abc_49347_n1331) );
  OR2X2 OR2X2_1900 ( .A(u0_u2__abc_44109_n340_bF_buf2), .B(\wb_data_i[7] ), .Y(u0_u2__abc_44109_n369) );
  OR2X2 OR2X2_1901 ( .A(u0_u2_lmr_req_we_FF_INPUT_bF_buf0), .B(u0_tms2_8_), .Y(u0_u2__abc_44109_n372) );
  OR2X2 OR2X2_1902 ( .A(u0_u2__abc_44109_n340_bF_buf1), .B(\wb_data_i[8] ), .Y(u0_u2__abc_44109_n373) );
  OR2X2 OR2X2_1903 ( .A(u0_u2_lmr_req_we_FF_INPUT_bF_buf4), .B(u0_tms2_9_), .Y(u0_u2__abc_44109_n376) );
  OR2X2 OR2X2_1904 ( .A(u0_u2__abc_44109_n340_bF_buf0), .B(\wb_data_i[9] ), .Y(u0_u2__abc_44109_n377) );
  OR2X2 OR2X2_1905 ( .A(u0_u2_lmr_req_we_FF_INPUT_bF_buf3), .B(u0_tms2_10_), .Y(u0_u2__abc_44109_n380) );
  OR2X2 OR2X2_1906 ( .A(u0_u2__abc_44109_n340_bF_buf4), .B(\wb_data_i[10] ), .Y(u0_u2__abc_44109_n381) );
  OR2X2 OR2X2_1907 ( .A(u0_u2_lmr_req_we_FF_INPUT_bF_buf2), .B(u0_tms2_11_), .Y(u0_u2__abc_44109_n384) );
  OR2X2 OR2X2_1908 ( .A(u0_u2__abc_44109_n340_bF_buf3), .B(\wb_data_i[11] ), .Y(u0_u2__abc_44109_n385) );
  OR2X2 OR2X2_1909 ( .A(u0_u2_lmr_req_we_FF_INPUT_bF_buf1), .B(u0_tms2_12_), .Y(u0_u2__abc_44109_n388) );
  OR2X2 OR2X2_191 ( .A(u0__abc_49347_n1333), .B(u0__abc_49347_n1329), .Y(u0__abc_49347_n1334) );
  OR2X2 OR2X2_1910 ( .A(u0_u2__abc_44109_n340_bF_buf2), .B(\wb_data_i[12] ), .Y(u0_u2__abc_44109_n389) );
  OR2X2 OR2X2_1911 ( .A(u0_u2_lmr_req_we_FF_INPUT_bF_buf0), .B(u0_tms2_13_), .Y(u0_u2__abc_44109_n392) );
  OR2X2 OR2X2_1912 ( .A(u0_u2__abc_44109_n340_bF_buf1), .B(\wb_data_i[13] ), .Y(u0_u2__abc_44109_n393) );
  OR2X2 OR2X2_1913 ( .A(u0_u2_lmr_req_we_FF_INPUT_bF_buf4), .B(u0_tms2_14_), .Y(u0_u2__abc_44109_n396) );
  OR2X2 OR2X2_1914 ( .A(u0_u2__abc_44109_n340_bF_buf0), .B(\wb_data_i[14] ), .Y(u0_u2__abc_44109_n397) );
  OR2X2 OR2X2_1915 ( .A(u0_u2_lmr_req_we_FF_INPUT_bF_buf3), .B(u0_tms2_15_), .Y(u0_u2__abc_44109_n400) );
  OR2X2 OR2X2_1916 ( .A(u0_u2__abc_44109_n340_bF_buf4), .B(\wb_data_i[15] ), .Y(u0_u2__abc_44109_n401) );
  OR2X2 OR2X2_1917 ( .A(u0_u2_lmr_req_we_FF_INPUT_bF_buf2), .B(u0_tms2_16_), .Y(u0_u2__abc_44109_n404) );
  OR2X2 OR2X2_1918 ( .A(u0_u2__abc_44109_n340_bF_buf3), .B(\wb_data_i[16] ), .Y(u0_u2__abc_44109_n405) );
  OR2X2 OR2X2_1919 ( .A(u0_u2_lmr_req_we_FF_INPUT_bF_buf1), .B(u0_tms2_17_), .Y(u0_u2__abc_44109_n408) );
  OR2X2 OR2X2_192 ( .A(u0__abc_49347_n1335_1), .B(u0__abc_49347_n1336_1), .Y(u0__abc_49347_n1337) );
  OR2X2 OR2X2_1920 ( .A(u0_u2__abc_44109_n340_bF_buf2), .B(\wb_data_i[17] ), .Y(u0_u2__abc_44109_n409) );
  OR2X2 OR2X2_1921 ( .A(u0_u2_lmr_req_we_FF_INPUT_bF_buf0), .B(u0_tms2_18_), .Y(u0_u2__abc_44109_n412) );
  OR2X2 OR2X2_1922 ( .A(u0_u2__abc_44109_n340_bF_buf1), .B(\wb_data_i[18] ), .Y(u0_u2__abc_44109_n413) );
  OR2X2 OR2X2_1923 ( .A(u0_u2_lmr_req_we_FF_INPUT_bF_buf4), .B(u0_tms2_19_), .Y(u0_u2__abc_44109_n416) );
  OR2X2 OR2X2_1924 ( .A(u0_u2__abc_44109_n340_bF_buf0), .B(\wb_data_i[19] ), .Y(u0_u2__abc_44109_n417) );
  OR2X2 OR2X2_1925 ( .A(u0_u2_lmr_req_we_FF_INPUT_bF_buf3), .B(u0_tms2_20_), .Y(u0_u2__abc_44109_n420) );
  OR2X2 OR2X2_1926 ( .A(u0_u2__abc_44109_n340_bF_buf4), .B(\wb_data_i[20] ), .Y(u0_u2__abc_44109_n421) );
  OR2X2 OR2X2_1927 ( .A(u0_u2_lmr_req_we_FF_INPUT_bF_buf2), .B(u0_tms2_21_), .Y(u0_u2__abc_44109_n424) );
  OR2X2 OR2X2_1928 ( .A(u0_u2__abc_44109_n340_bF_buf3), .B(\wb_data_i[21] ), .Y(u0_u2__abc_44109_n425) );
  OR2X2 OR2X2_1929 ( .A(u0_u2_lmr_req_we_FF_INPUT_bF_buf1), .B(u0_tms2_22_), .Y(u0_u2__abc_44109_n428) );
  OR2X2 OR2X2_193 ( .A(u0__abc_49347_n1338), .B(u0__abc_49347_n1339), .Y(u0__abc_49347_n1340) );
  OR2X2 OR2X2_1930 ( .A(u0_u2__abc_44109_n340_bF_buf2), .B(\wb_data_i[22] ), .Y(u0_u2__abc_44109_n429) );
  OR2X2 OR2X2_1931 ( .A(u0_u2_lmr_req_we_FF_INPUT_bF_buf0), .B(u0_tms2_23_), .Y(u0_u2__abc_44109_n432) );
  OR2X2 OR2X2_1932 ( .A(u0_u2__abc_44109_n340_bF_buf1), .B(\wb_data_i[23] ), .Y(u0_u2__abc_44109_n433) );
  OR2X2 OR2X2_1933 ( .A(u0_u2_lmr_req_we_FF_INPUT_bF_buf4), .B(u0_tms2_24_), .Y(u0_u2__abc_44109_n436) );
  OR2X2 OR2X2_1934 ( .A(u0_u2__abc_44109_n340_bF_buf0), .B(\wb_data_i[24] ), .Y(u0_u2__abc_44109_n437) );
  OR2X2 OR2X2_1935 ( .A(u0_u2_lmr_req_we_FF_INPUT_bF_buf3), .B(u0_tms2_25_), .Y(u0_u2__abc_44109_n440) );
  OR2X2 OR2X2_1936 ( .A(u0_u2__abc_44109_n340_bF_buf4), .B(\wb_data_i[25] ), .Y(u0_u2__abc_44109_n441) );
  OR2X2 OR2X2_1937 ( .A(u0_u2_lmr_req_we_FF_INPUT_bF_buf2), .B(u0_tms2_26_), .Y(u0_u2__abc_44109_n444) );
  OR2X2 OR2X2_1938 ( .A(u0_u2__abc_44109_n340_bF_buf3), .B(\wb_data_i[26] ), .Y(u0_u2__abc_44109_n445) );
  OR2X2 OR2X2_1939 ( .A(u0_u2_lmr_req_we_FF_INPUT_bF_buf1), .B(u0_tms2_27_), .Y(u0_u2__abc_44109_n448) );
  OR2X2 OR2X2_194 ( .A(u0__abc_49347_n1341), .B(u0__abc_49347_n1342), .Y(u0__abc_49347_n1343) );
  OR2X2 OR2X2_1940 ( .A(u0_u2__abc_44109_n340_bF_buf2), .B(\wb_data_i[27] ), .Y(u0_u2__abc_44109_n449) );
  OR2X2 OR2X2_1941 ( .A(u0_u2_lmr_req_we_FF_INPUT_bF_buf0), .B(u0_tms2_28_), .Y(u0_u2__abc_44109_n452) );
  OR2X2 OR2X2_1942 ( .A(u0_u2__abc_44109_n340_bF_buf1), .B(\wb_data_i[28] ), .Y(u0_u2__abc_44109_n453) );
  OR2X2 OR2X2_1943 ( .A(u0_u2_lmr_req_we_FF_INPUT_bF_buf4), .B(u0_tms2_29_), .Y(u0_u2__abc_44109_n456) );
  OR2X2 OR2X2_1944 ( .A(u0_u2__abc_44109_n340_bF_buf0), .B(\wb_data_i[29] ), .Y(u0_u2__abc_44109_n457) );
  OR2X2 OR2X2_1945 ( .A(u0_u2_lmr_req_we_FF_INPUT_bF_buf3), .B(u0_tms2_30_), .Y(u0_u2__abc_44109_n460) );
  OR2X2 OR2X2_1946 ( .A(u0_u2__abc_44109_n340_bF_buf4), .B(\wb_data_i[30] ), .Y(u0_u2__abc_44109_n461) );
  OR2X2 OR2X2_1947 ( .A(u0_u2_lmr_req_we_FF_INPUT_bF_buf2), .B(u0_tms2_31_), .Y(u0_u2__abc_44109_n464) );
  OR2X2 OR2X2_1948 ( .A(u0_u2__abc_44109_n340_bF_buf3), .B(\wb_data_i[31] ), .Y(u0_u2__abc_44109_n465) );
  OR2X2 OR2X2_1949 ( .A(u0_csc2_1_), .B(u0_csc2_2_), .Y(u0_u2__abc_44109_n468) );
  OR2X2 OR2X2_195 ( .A(u0__abc_49347_n1345_1), .B(spec_req_cs_0_bF_buf2), .Y(u0__abc_49347_n1346) );
  OR2X2 OR2X2_1950 ( .A(u0_u2__abc_44109_n468), .B(u0_csc2_3_), .Y(u0_u2__abc_44109_n469) );
  OR2X2 OR2X2_1951 ( .A(u0_u2__abc_44109_n476), .B(u0_u2__abc_44109_n472), .Y(u0_u2_lmr_req_FF_INPUT) );
  OR2X2 OR2X2_1952 ( .A(u0_u2__abc_44109_n483), .B(u0_u2__abc_44109_n479), .Y(u0_u2_init_req_FF_INPUT) );
  OR2X2 OR2X2_1953 ( .A(u0_u2_inited), .B(u0_init_ack2), .Y(u0_u2_inited_FF_INPUT) );
  OR2X2 OR2X2_1954 ( .A(u0_u2__abc_44109_n489), .B(u0_u2__abc_44109_n487), .Y(u0_u2__abc_44109_n490) );
  OR2X2 OR2X2_1955 ( .A(u0_u2__abc_44109_n493), .B(u0_u2__abc_44109_n491), .Y(u0_u2__abc_44109_n494) );
  OR2X2 OR2X2_1956 ( .A(u0_u2__abc_44109_n500), .B(u0_u2__abc_44109_n492), .Y(u0_u2__abc_44109_n501) );
  OR2X2 OR2X2_1957 ( .A(u0_u2__abc_44109_n506), .B(u0_u2__abc_44109_n504), .Y(u0_u2__abc_44109_n507) );
  OR2X2 OR2X2_1958 ( .A(u0_u2__abc_44109_n510), .B(u0_u2__abc_44109_n508), .Y(u0_u2__abc_44109_n511) );
  OR2X2 OR2X2_1959 ( .A(u0_u2__abc_44109_n516), .B(u0_u2__abc_44109_n509), .Y(u0_u2__abc_44109_n517) );
  OR2X2 OR2X2_196 ( .A(u0__abc_49347_n1344_1), .B(u0__abc_49347_n1346), .Y(u0__abc_49347_n1347) );
  OR2X2 OR2X2_1960 ( .A(u0_u2__abc_44109_n524), .B(u0_u2__abc_44109_n525), .Y(u0_u2__abc_44109_n526) );
  OR2X2 OR2X2_1961 ( .A(u0_u2__abc_44109_n528), .B(u0_u2__abc_44109_n523), .Y(u0_u2__abc_44109_n529) );
  OR2X2 OR2X2_1962 ( .A(u0_u2__abc_44109_n533), .B(u0_u2__abc_44109_n497), .Y(u0_u2__abc_44109_n534) );
  OR2X2 OR2X2_1963 ( .A(u0_u2__abc_44109_n537), .B(u0_u2__abc_44109_n535), .Y(u0_u2__abc_44109_n538) );
  OR2X2 OR2X2_1964 ( .A(u0_u2__abc_44109_n542), .B(u0_u2__abc_44109_n540), .Y(u0_u2__abc_44109_n543) );
  OR2X2 OR2X2_1965 ( .A(u0_u2__abc_44109_n544), .B(u0_u2__abc_44109_n536), .Y(u0_u2__abc_44109_n545) );
  OR2X2 OR2X2_1966 ( .A(u0_u2__abc_44109_n548), .B(u0_u2__abc_44109_n541), .Y(u0_u2__abc_44109_n549) );
  OR2X2 OR2X2_1967 ( .A(u0_u3_init_req_we_FF_INPUT_bF_buf5), .B(u0_csc3_0_), .Y(u0_u3__abc_44466_n214_1) );
  OR2X2 OR2X2_1968 ( .A(u0_u3__abc_44466_n220_1), .B(u0_u3__abc_44466_n221_1), .Y(u0_u3__abc_44466_n222) );
  OR2X2 OR2X2_1969 ( .A(u0_u3__abc_44466_n219), .B(u0_u3__abc_44466_n222), .Y(u0_u3_csc_0__FF_INPUT) );
  OR2X2 OR2X2_197 ( .A(u0__abc_49347_n1203_bF_buf5), .B(u0_tms0_6_), .Y(u0__abc_49347_n1348) );
  OR2X2 OR2X2_1970 ( .A(u0_u3_init_req_we_FF_INPUT_bF_buf3), .B(u0_csc3_1_), .Y(u0_u3__abc_44466_n224_1) );
  OR2X2 OR2X2_1971 ( .A(u0_u3__abc_44466_n229_1), .B(u0_u3__abc_44466_n220_1), .Y(u0_u3_csc_1__FF_INPUT) );
  OR2X2 OR2X2_1972 ( .A(u0_u3_init_req_we_FF_INPUT_bF_buf1), .B(u0_csc3_2_), .Y(u0_u3__abc_44466_n231) );
  OR2X2 OR2X2_1973 ( .A(u0_u3__abc_44466_n236_1), .B(u0_u3__abc_44466_n221_1), .Y(u0_u3_csc_2__FF_INPUT) );
  OR2X2 OR2X2_1974 ( .A(u0_u3__abc_44466_n240), .B(u0_u3__abc_44466_n238_1), .Y(u0_u3__abc_44466_n241_1) );
  OR2X2 OR2X2_1975 ( .A(u0_u3_init_req_we_FF_INPUT_bF_buf3), .B(u0_csc3_4_), .Y(u0_u3__abc_44466_n243) );
  OR2X2 OR2X2_1976 ( .A(u0_u3__abc_44466_n247), .B(u0_u3_rst_r2_bF_buf2), .Y(u0_u3__abc_44466_n248) );
  OR2X2 OR2X2_1977 ( .A(u0_u3__abc_44466_n205_1_bF_buf0), .B(_auto_iopadmap_cc_313_execute_56321_0_), .Y(u0_u3__abc_44466_n249) );
  OR2X2 OR2X2_1978 ( .A(u0_u3_init_req_we_FF_INPUT_bF_buf1), .B(u0_csc3_5_), .Y(u0_u3__abc_44466_n251) );
  OR2X2 OR2X2_1979 ( .A(u0_u3__abc_44466_n255_1), .B(u0_u3_rst_r2_bF_buf1), .Y(u0_u3__abc_44466_n256_1) );
  OR2X2 OR2X2_198 ( .A(u0__abc_49347_n1350), .B(u0__abc_49347_n1328), .Y(u0_sp_tms_6__FF_INPUT) );
  OR2X2 OR2X2_1980 ( .A(u0_u3__abc_44466_n205_1_bF_buf4), .B(_auto_iopadmap_cc_313_execute_56321_1_), .Y(u0_u3__abc_44466_n257) );
  OR2X2 OR2X2_1981 ( .A(u0_u3__abc_44466_n260_1), .B(u0_u3__abc_44466_n259), .Y(u0_u3__abc_44466_n261) );
  OR2X2 OR2X2_1982 ( .A(u0_u3__abc_44466_n264_1), .B(u0_u3__abc_44466_n263_1), .Y(u0_u3__abc_44466_n265_1) );
  OR2X2 OR2X2_1983 ( .A(u0_u3__abc_44466_n268), .B(u0_u3__abc_44466_n267_1), .Y(u0_u3__abc_44466_n269) );
  OR2X2 OR2X2_1984 ( .A(u0_u3__abc_44466_n272_1), .B(u0_u3__abc_44466_n271), .Y(u0_u3__abc_44466_n273) );
  OR2X2 OR2X2_1985 ( .A(u0_u3__abc_44466_n276), .B(u0_u3__abc_44466_n275), .Y(u0_u3__abc_44466_n277) );
  OR2X2 OR2X2_1986 ( .A(u0_u3__abc_44466_n280_1), .B(u0_u3__abc_44466_n279), .Y(u0_u3__abc_44466_n281) );
  OR2X2 OR2X2_1987 ( .A(u0_u3__abc_44466_n284), .B(u0_u3__abc_44466_n283), .Y(u0_u3__abc_44466_n285_1) );
  OR2X2 OR2X2_1988 ( .A(u0_u3__abc_44466_n288), .B(u0_u3__abc_44466_n287_1), .Y(u0_u3__abc_44466_n289_1) );
  OR2X2 OR2X2_1989 ( .A(u0_u3__abc_44466_n292), .B(u0_u3__abc_44466_n291_1), .Y(u0_u3__abc_44466_n293) );
  OR2X2 OR2X2_199 ( .A(u0__abc_49347_n1183_1_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n1354_1) );
  OR2X2 OR2X2_1990 ( .A(u0_u3__abc_44466_n296), .B(u0_u3__abc_44466_n295_1), .Y(u0_u3__abc_44466_n297_1) );
  OR2X2 OR2X2_1991 ( .A(u0_u3__abc_44466_n300), .B(u0_u3__abc_44466_n299_1), .Y(u0_u3__abc_44466_n301_1) );
  OR2X2 OR2X2_1992 ( .A(u0_u3__abc_44466_n304), .B(u0_u3__abc_44466_n303), .Y(u0_u3__abc_44466_n305) );
  OR2X2 OR2X2_1993 ( .A(u0_u3__abc_44466_n308_1), .B(u0_u3__abc_44466_n307), .Y(u0_u3__abc_44466_n309) );
  OR2X2 OR2X2_1994 ( .A(u0_u3__abc_44466_n312), .B(u0_u3__abc_44466_n311), .Y(u0_u3__abc_44466_n313) );
  OR2X2 OR2X2_1995 ( .A(u0_u3__abc_44466_n316), .B(u0_u3__abc_44466_n315), .Y(u0_u3__abc_44466_n317) );
  OR2X2 OR2X2_1996 ( .A(u0_u3__abc_44466_n320), .B(u0_u3__abc_44466_n319), .Y(u0_u3__abc_44466_n321) );
  OR2X2 OR2X2_1997 ( .A(u0_u3__abc_44466_n324_1), .B(u0_u3__abc_44466_n323), .Y(u0_u3__abc_44466_n325) );
  OR2X2 OR2X2_1998 ( .A(u0_u3__abc_44466_n328_1), .B(u0_u3__abc_44466_n327_1), .Y(u0_u3__abc_44466_n329) );
  OR2X2 OR2X2_1999 ( .A(u0_u3__abc_44466_n332), .B(u0_u3__abc_44466_n331), .Y(u0_u3__abc_44466_n333) );
  OR2X2 OR2X2_2 ( .A(susp_sel), .B(rfr_ack), .Y(_abc_55805_n237_1) );
  OR2X2 OR2X2_20 ( .A(lmr_sel_bF_buf2), .B(cs_4_), .Y(_abc_55805_n267) );
  OR2X2 OR2X2_200 ( .A(spec_req_cs_6_bF_buf1), .B(1'b0), .Y(u0__abc_49347_n1355) );
  OR2X2 OR2X2_2000 ( .A(u0_u3__abc_44466_n336), .B(u0_u3__abc_44466_n335), .Y(u0_u3__abc_44466_n337) );
  OR2X2 OR2X2_2001 ( .A(u0_u3__abc_44466_n340), .B(u0_u3__abc_44466_n339), .Y(u0_u3__abc_44466_n341) );
  OR2X2 OR2X2_2002 ( .A(u0_u3__abc_44466_n344), .B(u0_u3__abc_44466_n343), .Y(u0_u3__abc_44466_n345) );
  OR2X2 OR2X2_2003 ( .A(u0_u3__abc_44466_n348), .B(u0_u3__abc_44466_n347), .Y(u0_u3__abc_44466_n349) );
  OR2X2 OR2X2_2004 ( .A(u0_u3__abc_44466_n352), .B(u0_u3__abc_44466_n351), .Y(u0_u3__abc_44466_n353) );
  OR2X2 OR2X2_2005 ( .A(u0_u3__abc_44466_n356), .B(u0_u3__abc_44466_n355), .Y(u0_u3__abc_44466_n357) );
  OR2X2 OR2X2_2006 ( .A(u0_u3__abc_44466_n360), .B(u0_u3__abc_44466_n359), .Y(u0_u3__abc_44466_n361) );
  OR2X2 OR2X2_2007 ( .A(u0_u3__abc_44466_n366), .B(u0_u3_rst_r2_bF_buf0), .Y(u0_u3__abc_44466_n367) );
  OR2X2 OR2X2_2008 ( .A(u0_u3__abc_44466_n367), .B(u0_u3__abc_44466_n365), .Y(u0_u3_tms_0__FF_INPUT) );
  OR2X2 OR2X2_2009 ( .A(u0_u3__abc_44466_n370), .B(u0_u3_rst_r2_bF_buf5), .Y(u0_u3__abc_44466_n371) );
  OR2X2 OR2X2_201 ( .A(u0__abc_49347_n1357), .B(u0__abc_49347_n1353_1), .Y(u0__abc_49347_n1358) );
  OR2X2 OR2X2_2010 ( .A(u0_u3__abc_44466_n371), .B(u0_u3__abc_44466_n369), .Y(u0_u3_tms_1__FF_INPUT) );
  OR2X2 OR2X2_2011 ( .A(u0_u3__abc_44466_n374), .B(u0_u3_rst_r2_bF_buf4), .Y(u0_u3__abc_44466_n375) );
  OR2X2 OR2X2_2012 ( .A(u0_u3__abc_44466_n375), .B(u0_u3__abc_44466_n373), .Y(u0_u3_tms_2__FF_INPUT) );
  OR2X2 OR2X2_2013 ( .A(u0_u3__abc_44466_n378), .B(u0_u3_rst_r2_bF_buf3), .Y(u0_u3__abc_44466_n379) );
  OR2X2 OR2X2_2014 ( .A(u0_u3__abc_44466_n379), .B(u0_u3__abc_44466_n377), .Y(u0_u3_tms_3__FF_INPUT) );
  OR2X2 OR2X2_2015 ( .A(u0_u3__abc_44466_n382), .B(u0_u3_rst_r2_bF_buf2), .Y(u0_u3__abc_44466_n383) );
  OR2X2 OR2X2_2016 ( .A(u0_u3__abc_44466_n383), .B(u0_u3__abc_44466_n381), .Y(u0_u3_tms_4__FF_INPUT) );
  OR2X2 OR2X2_2017 ( .A(u0_u3__abc_44466_n386), .B(u0_u3_rst_r2_bF_buf1), .Y(u0_u3__abc_44466_n387) );
  OR2X2 OR2X2_2018 ( .A(u0_u3__abc_44466_n387), .B(u0_u3__abc_44466_n385), .Y(u0_u3_tms_5__FF_INPUT) );
  OR2X2 OR2X2_2019 ( .A(u0_u3__abc_44466_n390), .B(u0_u3_rst_r2_bF_buf0), .Y(u0_u3__abc_44466_n391) );
  OR2X2 OR2X2_202 ( .A(u0__abc_49347_n1359), .B(u0__abc_49347_n1360), .Y(u0__abc_49347_n1361) );
  OR2X2 OR2X2_2020 ( .A(u0_u3__abc_44466_n391), .B(u0_u3__abc_44466_n389), .Y(u0_u3_tms_6__FF_INPUT) );
  OR2X2 OR2X2_2021 ( .A(u0_u3__abc_44466_n394), .B(u0_u3_rst_r2_bF_buf5), .Y(u0_u3__abc_44466_n395) );
  OR2X2 OR2X2_2022 ( .A(u0_u3__abc_44466_n395), .B(u0_u3__abc_44466_n393), .Y(u0_u3_tms_7__FF_INPUT) );
  OR2X2 OR2X2_2023 ( .A(u0_u3__abc_44466_n398), .B(u0_u3_rst_r2_bF_buf4), .Y(u0_u3__abc_44466_n399) );
  OR2X2 OR2X2_2024 ( .A(u0_u3__abc_44466_n399), .B(u0_u3__abc_44466_n397), .Y(u0_u3_tms_8__FF_INPUT) );
  OR2X2 OR2X2_2025 ( .A(u0_u3__abc_44466_n402), .B(u0_u3_rst_r2_bF_buf3), .Y(u0_u3__abc_44466_n403) );
  OR2X2 OR2X2_2026 ( .A(u0_u3__abc_44466_n403), .B(u0_u3__abc_44466_n401), .Y(u0_u3_tms_9__FF_INPUT) );
  OR2X2 OR2X2_2027 ( .A(u0_u3__abc_44466_n406), .B(u0_u3_rst_r2_bF_buf2), .Y(u0_u3__abc_44466_n407) );
  OR2X2 OR2X2_2028 ( .A(u0_u3__abc_44466_n407), .B(u0_u3__abc_44466_n405), .Y(u0_u3_tms_10__FF_INPUT) );
  OR2X2 OR2X2_2029 ( .A(u0_u3__abc_44466_n410), .B(u0_u3_rst_r2_bF_buf1), .Y(u0_u3__abc_44466_n411) );
  OR2X2 OR2X2_203 ( .A(u0__abc_49347_n1362_1), .B(u0__abc_49347_n1363_1), .Y(u0__abc_49347_n1364) );
  OR2X2 OR2X2_2030 ( .A(u0_u3__abc_44466_n411), .B(u0_u3__abc_44466_n409), .Y(u0_u3_tms_11__FF_INPUT) );
  OR2X2 OR2X2_2031 ( .A(u0_u3__abc_44466_n414), .B(u0_u3_rst_r2_bF_buf0), .Y(u0_u3__abc_44466_n415) );
  OR2X2 OR2X2_2032 ( .A(u0_u3__abc_44466_n415), .B(u0_u3__abc_44466_n413), .Y(u0_u3_tms_12__FF_INPUT) );
  OR2X2 OR2X2_2033 ( .A(u0_u3__abc_44466_n418), .B(u0_u3_rst_r2_bF_buf5), .Y(u0_u3__abc_44466_n419) );
  OR2X2 OR2X2_2034 ( .A(u0_u3__abc_44466_n419), .B(u0_u3__abc_44466_n417), .Y(u0_u3_tms_13__FF_INPUT) );
  OR2X2 OR2X2_2035 ( .A(u0_u3__abc_44466_n422), .B(u0_u3_rst_r2_bF_buf4), .Y(u0_u3__abc_44466_n423) );
  OR2X2 OR2X2_2036 ( .A(u0_u3__abc_44466_n423), .B(u0_u3__abc_44466_n421), .Y(u0_u3_tms_14__FF_INPUT) );
  OR2X2 OR2X2_2037 ( .A(u0_u3__abc_44466_n426), .B(u0_u3_rst_r2_bF_buf3), .Y(u0_u3__abc_44466_n427) );
  OR2X2 OR2X2_2038 ( .A(u0_u3__abc_44466_n427), .B(u0_u3__abc_44466_n425), .Y(u0_u3_tms_15__FF_INPUT) );
  OR2X2 OR2X2_2039 ( .A(u0_u3__abc_44466_n430), .B(u0_u3_rst_r2_bF_buf2), .Y(u0_u3__abc_44466_n431) );
  OR2X2 OR2X2_204 ( .A(u0__abc_49347_n1365), .B(u0__abc_49347_n1366), .Y(u0__abc_49347_n1367) );
  OR2X2 OR2X2_2040 ( .A(u0_u3__abc_44466_n431), .B(u0_u3__abc_44466_n429), .Y(u0_u3_tms_16__FF_INPUT) );
  OR2X2 OR2X2_2041 ( .A(u0_u3__abc_44466_n434), .B(u0_u3_rst_r2_bF_buf1), .Y(u0_u3__abc_44466_n435) );
  OR2X2 OR2X2_2042 ( .A(u0_u3__abc_44466_n435), .B(u0_u3__abc_44466_n433), .Y(u0_u3_tms_17__FF_INPUT) );
  OR2X2 OR2X2_2043 ( .A(u0_u3__abc_44466_n438), .B(u0_u3_rst_r2_bF_buf0), .Y(u0_u3__abc_44466_n439) );
  OR2X2 OR2X2_2044 ( .A(u0_u3__abc_44466_n439), .B(u0_u3__abc_44466_n437), .Y(u0_u3_tms_18__FF_INPUT) );
  OR2X2 OR2X2_2045 ( .A(u0_u3__abc_44466_n442), .B(u0_u3_rst_r2_bF_buf5), .Y(u0_u3__abc_44466_n443) );
  OR2X2 OR2X2_2046 ( .A(u0_u3__abc_44466_n443), .B(u0_u3__abc_44466_n441), .Y(u0_u3_tms_19__FF_INPUT) );
  OR2X2 OR2X2_2047 ( .A(u0_u3__abc_44466_n446), .B(u0_u3_rst_r2_bF_buf4), .Y(u0_u3__abc_44466_n447) );
  OR2X2 OR2X2_2048 ( .A(u0_u3__abc_44466_n447), .B(u0_u3__abc_44466_n445), .Y(u0_u3_tms_20__FF_INPUT) );
  OR2X2 OR2X2_2049 ( .A(u0_u3__abc_44466_n450), .B(u0_u3_rst_r2_bF_buf3), .Y(u0_u3__abc_44466_n451) );
  OR2X2 OR2X2_205 ( .A(u0__abc_49347_n1369), .B(spec_req_cs_0_bF_buf1), .Y(u0__abc_49347_n1370) );
  OR2X2 OR2X2_2050 ( .A(u0_u3__abc_44466_n451), .B(u0_u3__abc_44466_n449), .Y(u0_u3_tms_21__FF_INPUT) );
  OR2X2 OR2X2_2051 ( .A(u0_u3__abc_44466_n454), .B(u0_u3_rst_r2_bF_buf2), .Y(u0_u3__abc_44466_n455) );
  OR2X2 OR2X2_2052 ( .A(u0_u3__abc_44466_n455), .B(u0_u3__abc_44466_n453), .Y(u0_u3_tms_22__FF_INPUT) );
  OR2X2 OR2X2_2053 ( .A(u0_u3__abc_44466_n458), .B(u0_u3_rst_r2_bF_buf1), .Y(u0_u3__abc_44466_n459) );
  OR2X2 OR2X2_2054 ( .A(u0_u3__abc_44466_n459), .B(u0_u3__abc_44466_n457), .Y(u0_u3_tms_23__FF_INPUT) );
  OR2X2 OR2X2_2055 ( .A(u0_u3__abc_44466_n462), .B(u0_u3_rst_r2_bF_buf0), .Y(u0_u3__abc_44466_n463) );
  OR2X2 OR2X2_2056 ( .A(u0_u3__abc_44466_n463), .B(u0_u3__abc_44466_n461), .Y(u0_u3_tms_24__FF_INPUT) );
  OR2X2 OR2X2_2057 ( .A(u0_u3__abc_44466_n466), .B(u0_u3_rst_r2_bF_buf5), .Y(u0_u3__abc_44466_n467) );
  OR2X2 OR2X2_2058 ( .A(u0_u3__abc_44466_n467), .B(u0_u3__abc_44466_n465), .Y(u0_u3_tms_25__FF_INPUT) );
  OR2X2 OR2X2_2059 ( .A(u0_u3__abc_44466_n470), .B(u0_u3_rst_r2_bF_buf4), .Y(u0_u3__abc_44466_n471) );
  OR2X2 OR2X2_206 ( .A(u0__abc_49347_n1368), .B(u0__abc_49347_n1370), .Y(u0__abc_49347_n1371_1) );
  OR2X2 OR2X2_2060 ( .A(u0_u3__abc_44466_n471), .B(u0_u3__abc_44466_n469), .Y(u0_u3_tms_26__FF_INPUT) );
  OR2X2 OR2X2_2061 ( .A(u0_u3__abc_44466_n474), .B(u0_u3_rst_r2_bF_buf3), .Y(u0_u3__abc_44466_n475) );
  OR2X2 OR2X2_2062 ( .A(u0_u3__abc_44466_n475), .B(u0_u3__abc_44466_n473), .Y(u0_u3_tms_27__FF_INPUT) );
  OR2X2 OR2X2_2063 ( .A(u0_u3__abc_44466_n478), .B(u0_u3_rst_r2_bF_buf2), .Y(u0_u3__abc_44466_n479) );
  OR2X2 OR2X2_2064 ( .A(u0_u3__abc_44466_n479), .B(u0_u3__abc_44466_n477), .Y(u0_u3_tms_28__FF_INPUT) );
  OR2X2 OR2X2_2065 ( .A(u0_u3__abc_44466_n482), .B(u0_u3_rst_r2_bF_buf1), .Y(u0_u3__abc_44466_n483) );
  OR2X2 OR2X2_2066 ( .A(u0_u3__abc_44466_n483), .B(u0_u3__abc_44466_n481), .Y(u0_u3_tms_29__FF_INPUT) );
  OR2X2 OR2X2_2067 ( .A(u0_u3__abc_44466_n486), .B(u0_u3_rst_r2_bF_buf0), .Y(u0_u3__abc_44466_n487) );
  OR2X2 OR2X2_2068 ( .A(u0_u3__abc_44466_n487), .B(u0_u3__abc_44466_n485), .Y(u0_u3_tms_30__FF_INPUT) );
  OR2X2 OR2X2_2069 ( .A(u0_u3__abc_44466_n490), .B(u0_u3_rst_r2_bF_buf5), .Y(u0_u3__abc_44466_n491) );
  OR2X2 OR2X2_207 ( .A(u0__abc_49347_n1203_bF_buf4), .B(u0_tms0_7_), .Y(u0__abc_49347_n1372_1) );
  OR2X2 OR2X2_2070 ( .A(u0_u3__abc_44466_n491), .B(u0_u3__abc_44466_n489), .Y(u0_u3_tms_31__FF_INPUT) );
  OR2X2 OR2X2_2071 ( .A(u0_csc3_1_), .B(u0_csc3_2_), .Y(u0_u3__abc_44466_n493) );
  OR2X2 OR2X2_2072 ( .A(u0_u3__abc_44466_n493), .B(u0_csc3_3_), .Y(u0_u3__abc_44466_n494) );
  OR2X2 OR2X2_2073 ( .A(u0_u3__abc_44466_n501), .B(u0_u3__abc_44466_n497), .Y(u0_u3_lmr_req_FF_INPUT) );
  OR2X2 OR2X2_2074 ( .A(u0_u3__abc_44466_n508), .B(u0_u3__abc_44466_n504), .Y(u0_u3_init_req_FF_INPUT) );
  OR2X2 OR2X2_2075 ( .A(u0_u3_inited), .B(u0_init_ack3), .Y(u0_u3_inited_FF_INPUT) );
  OR2X2 OR2X2_2076 ( .A(u0_u3__abc_44466_n514), .B(u0_u3__abc_44466_n512), .Y(u0_u3__abc_44466_n515) );
  OR2X2 OR2X2_2077 ( .A(u0_u3__abc_44466_n518), .B(u0_u3__abc_44466_n516), .Y(u0_u3__abc_44466_n519) );
  OR2X2 OR2X2_2078 ( .A(u0_u3__abc_44466_n525), .B(u0_u3__abc_44466_n517), .Y(u0_u3__abc_44466_n526) );
  OR2X2 OR2X2_2079 ( .A(u0_u3__abc_44466_n531), .B(u0_u3__abc_44466_n529), .Y(u0_u3__abc_44466_n532) );
  OR2X2 OR2X2_208 ( .A(u0__abc_49347_n1374), .B(u0__abc_49347_n1352), .Y(u0_sp_tms_7__FF_INPUT) );
  OR2X2 OR2X2_2080 ( .A(u0_u3__abc_44466_n535), .B(u0_u3__abc_44466_n533), .Y(u0_u3__abc_44466_n536) );
  OR2X2 OR2X2_2081 ( .A(u0_u3__abc_44466_n541), .B(u0_u3__abc_44466_n534), .Y(u0_u3__abc_44466_n542) );
  OR2X2 OR2X2_2082 ( .A(u0_u3__abc_44466_n549), .B(u0_u3__abc_44466_n550), .Y(u0_u3__abc_44466_n551) );
  OR2X2 OR2X2_2083 ( .A(u0_u3__abc_44466_n553), .B(u0_u3__abc_44466_n548), .Y(u0_u3__abc_44466_n554) );
  OR2X2 OR2X2_2084 ( .A(u0_u3__abc_44466_n558), .B(u0_u3__abc_44466_n522), .Y(u0_u3__abc_44466_n559) );
  OR2X2 OR2X2_2085 ( .A(u0_u3__abc_44466_n562), .B(u0_u3__abc_44466_n560), .Y(u0_u3__abc_44466_n563) );
  OR2X2 OR2X2_2086 ( .A(u0_u3__abc_44466_n567), .B(u0_u3__abc_44466_n565), .Y(u0_u3__abc_44466_n568) );
  OR2X2 OR2X2_2087 ( .A(u0_u3__abc_44466_n569), .B(u0_u3__abc_44466_n561), .Y(u0_u3__abc_44466_n570) );
  OR2X2 OR2X2_2088 ( .A(u0_u3__abc_44466_n573), .B(u0_u3__abc_44466_n566), .Y(u0_u3__abc_44466_n574) );
  OR2X2 OR2X2_2089 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf7), .B(u0_tms4_0_), .Y(u0_u4__abc_44844_n208) );
  OR2X2 OR2X2_209 ( .A(u0__abc_49347_n1183_1_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n1378) );
  OR2X2 OR2X2_2090 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf5), .B(u0_tms4_1_), .Y(u0_u4__abc_44844_n215_1) );
  OR2X2 OR2X2_2091 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf3), .B(u0_tms4_2_), .Y(u0_u4__abc_44844_n221_1) );
  OR2X2 OR2X2_2092 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf1), .B(u0_tms4_3_), .Y(u0_u4__abc_44844_n227_1) );
  OR2X2 OR2X2_2093 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf7), .B(u0_tms4_4_), .Y(u0_u4__abc_44844_n233_1) );
  OR2X2 OR2X2_2094 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf5), .B(u0_tms4_5_), .Y(u0_u4__abc_44844_n239_1) );
  OR2X2 OR2X2_2095 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf3), .B(u0_tms4_6_), .Y(u0_u4__abc_44844_n245_1) );
  OR2X2 OR2X2_2096 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf1), .B(u0_tms4_7_), .Y(u0_u4__abc_44844_n251_1) );
  OR2X2 OR2X2_2097 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf7), .B(u0_tms4_8_), .Y(u0_u4__abc_44844_n257) );
  OR2X2 OR2X2_2098 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf5), .B(u0_tms4_9_), .Y(u0_u4__abc_44844_n263_1) );
  OR2X2 OR2X2_2099 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf3), .B(u0_tms4_10_), .Y(u0_u4__abc_44844_n269) );
  OR2X2 OR2X2_21 ( .A(_abc_55805_n268), .B(_abc_55805_n237_1), .Y(_abc_55805_n269) );
  OR2X2 OR2X2_210 ( .A(spec_req_cs_6_bF_buf0), .B(1'b0), .Y(u0__abc_49347_n1379) );
  OR2X2 OR2X2_2100 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf1), .B(u0_tms4_11_), .Y(u0_u4__abc_44844_n275) );
  OR2X2 OR2X2_2101 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf7), .B(u0_tms4_12_), .Y(u0_u4__abc_44844_n281_1) );
  OR2X2 OR2X2_2102 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf5), .B(u0_tms4_13_), .Y(u0_u4__abc_44844_n287_1) );
  OR2X2 OR2X2_2103 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf3), .B(u0_tms4_14_), .Y(u0_u4__abc_44844_n293_1) );
  OR2X2 OR2X2_2104 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf1), .B(u0_tms4_15_), .Y(u0_u4__abc_44844_n299) );
  OR2X2 OR2X2_2105 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf7), .B(u0_tms4_16_), .Y(u0_u4__abc_44844_n305) );
  OR2X2 OR2X2_2106 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf5), .B(u0_tms4_17_), .Y(u0_u4__abc_44844_n311) );
  OR2X2 OR2X2_2107 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf3), .B(u0_tms4_18_), .Y(u0_u4__abc_44844_n317) );
  OR2X2 OR2X2_2108 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf1), .B(u0_tms4_19_), .Y(u0_u4__abc_44844_n323_1) );
  OR2X2 OR2X2_2109 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf7), .B(u0_tms4_20_), .Y(u0_u4__abc_44844_n329) );
  OR2X2 OR2X2_211 ( .A(u0__abc_49347_n1381_1), .B(u0__abc_49347_n1377), .Y(u0__abc_49347_n1382) );
  OR2X2 OR2X2_2110 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf5), .B(u0_tms4_21_), .Y(u0_u4__abc_44844_n335) );
  OR2X2 OR2X2_2111 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf3), .B(u0_tms4_22_), .Y(u0_u4__abc_44844_n341) );
  OR2X2 OR2X2_2112 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf1), .B(u0_tms4_23_), .Y(u0_u4__abc_44844_n347) );
  OR2X2 OR2X2_2113 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf7), .B(u0_tms4_24_), .Y(u0_u4__abc_44844_n353) );
  OR2X2 OR2X2_2114 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf5), .B(u0_tms4_25_), .Y(u0_u4__abc_44844_n359) );
  OR2X2 OR2X2_2115 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf3), .B(u0_tms4_26_), .Y(u0_u4__abc_44844_n365) );
  OR2X2 OR2X2_2116 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf1), .B(u0_tms4_27_), .Y(u0_u4__abc_44844_n371) );
  OR2X2 OR2X2_2117 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf7), .B(u0_tms4_28_), .Y(u0_u4__abc_44844_n377) );
  OR2X2 OR2X2_2118 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf5), .B(u0_tms4_29_), .Y(u0_u4__abc_44844_n383) );
  OR2X2 OR2X2_2119 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf3), .B(u0_tms4_30_), .Y(u0_u4__abc_44844_n389) );
  OR2X2 OR2X2_212 ( .A(u0__abc_49347_n1383), .B(u0__abc_49347_n1384), .Y(u0__abc_49347_n1385) );
  OR2X2 OR2X2_2120 ( .A(u0_u4_lmr_req_we_FF_INPUT_bF_buf1), .B(u0_tms4_31_), .Y(u0_u4__abc_44844_n395) );
  OR2X2 OR2X2_2121 ( .A(u0_csc4_2_), .B(u0_csc4_1_), .Y(u0_u4__abc_44844_n401) );
  OR2X2 OR2X2_2122 ( .A(u0_u4__abc_44844_n401), .B(u0_csc4_3_), .Y(u0_u4__abc_44844_n402) );
  OR2X2 OR2X2_2123 ( .A(u0_u4__abc_44844_n409), .B(u0_u4__abc_44844_n405), .Y(u0_u4_lmr_req_FF_INPUT) );
  OR2X2 OR2X2_2124 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf7), .B(u0_csc4_0_), .Y(u0_u4__abc_44844_n413) );
  OR2X2 OR2X2_2125 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf5), .B(u0_csc4_1_), .Y(u0_u4__abc_44844_n418) );
  OR2X2 OR2X2_2126 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf3), .B(u0_csc4_2_), .Y(u0_u4__abc_44844_n423) );
  OR2X2 OR2X2_2127 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf1), .B(u0_csc4_3_), .Y(u0_u4__abc_44844_n428) );
  OR2X2 OR2X2_2128 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf7), .B(u0_csc4_4_), .Y(u0_u4__abc_44844_n433) );
  OR2X2 OR2X2_2129 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf5), .B(u0_csc4_5_), .Y(u0_u4__abc_44844_n438) );
  OR2X2 OR2X2_213 ( .A(u0__abc_49347_n1386), .B(u0__abc_49347_n1387), .Y(u0__abc_49347_n1388) );
  OR2X2 OR2X2_2130 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf3), .B(u0_csc4_6_), .Y(u0_u4__abc_44844_n443) );
  OR2X2 OR2X2_2131 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf1), .B(u0_csc4_7_), .Y(u0_u4__abc_44844_n448) );
  OR2X2 OR2X2_2132 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf7), .B(u0_csc4_8_), .Y(u0_u4__abc_44844_n453) );
  OR2X2 OR2X2_2133 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf5), .B(u0_csc4_9_), .Y(u0_u4__abc_44844_n458) );
  OR2X2 OR2X2_2134 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf3), .B(u0_csc4_10_), .Y(u0_u4__abc_44844_n463) );
  OR2X2 OR2X2_2135 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf1), .B(u0_csc4_11_), .Y(u0_u4__abc_44844_n468) );
  OR2X2 OR2X2_2136 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf7), .B(u0_csc4_12_), .Y(u0_u4__abc_44844_n473) );
  OR2X2 OR2X2_2137 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf5), .B(u0_csc4_13_), .Y(u0_u4__abc_44844_n478) );
  OR2X2 OR2X2_2138 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf3), .B(u0_csc4_14_), .Y(u0_u4__abc_44844_n483) );
  OR2X2 OR2X2_2139 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf1), .B(u0_csc4_15_), .Y(u0_u4__abc_44844_n488) );
  OR2X2 OR2X2_214 ( .A(u0__abc_49347_n1389_1), .B(u0__abc_49347_n1390_1), .Y(u0__abc_49347_n1391) );
  OR2X2 OR2X2_2140 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf7), .B(u0_csc4_16_), .Y(u0_u4__abc_44844_n493) );
  OR2X2 OR2X2_2141 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf5), .B(u0_csc4_17_), .Y(u0_u4__abc_44844_n498) );
  OR2X2 OR2X2_2142 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf3), .B(u0_csc4_18_), .Y(u0_u4__abc_44844_n503) );
  OR2X2 OR2X2_2143 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf1), .B(u0_csc4_19_), .Y(u0_u4__abc_44844_n508) );
  OR2X2 OR2X2_2144 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf7), .B(u0_csc4_20_), .Y(u0_u4__abc_44844_n513) );
  OR2X2 OR2X2_2145 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf5), .B(u0_csc4_21_), .Y(u0_u4__abc_44844_n518) );
  OR2X2 OR2X2_2146 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf3), .B(u0_csc4_22_), .Y(u0_u4__abc_44844_n523) );
  OR2X2 OR2X2_2147 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf1), .B(u0_csc4_23_), .Y(u0_u4__abc_44844_n528) );
  OR2X2 OR2X2_2148 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf7), .B(u0_csc4_24_), .Y(u0_u4__abc_44844_n533) );
  OR2X2 OR2X2_2149 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf5), .B(u0_csc4_25_), .Y(u0_u4__abc_44844_n538) );
  OR2X2 OR2X2_215 ( .A(u0__abc_49347_n1393), .B(spec_req_cs_0_bF_buf0), .Y(u0__abc_49347_n1394) );
  OR2X2 OR2X2_2150 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf3), .B(u0_csc4_26_), .Y(u0_u4__abc_44844_n543) );
  OR2X2 OR2X2_2151 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf1), .B(u0_csc4_27_), .Y(u0_u4__abc_44844_n548) );
  OR2X2 OR2X2_2152 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf7), .B(u0_csc4_28_), .Y(u0_u4__abc_44844_n553) );
  OR2X2 OR2X2_2153 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf5), .B(u0_csc4_29_), .Y(u0_u4__abc_44844_n558) );
  OR2X2 OR2X2_2154 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf3), .B(u0_csc4_30_), .Y(u0_u4__abc_44844_n563) );
  OR2X2 OR2X2_2155 ( .A(u0_u4_init_req_we_FF_INPUT_bF_buf1), .B(u0_csc4_31_), .Y(u0_u4__abc_44844_n568) );
  OR2X2 OR2X2_2156 ( .A(u0_u4__abc_44844_n578), .B(u0_u4__abc_44844_n574), .Y(u0_u4_init_req_FF_INPUT) );
  OR2X2 OR2X2_2157 ( .A(u0_u4_inited), .B(u0_init_ack4), .Y(u0_u4_inited_FF_INPUT) );
  OR2X2 OR2X2_2158 ( .A(u0_u4__abc_44844_n584), .B(u0_u4__abc_44844_n582), .Y(u0_u4__abc_44844_n585) );
  OR2X2 OR2X2_2159 ( .A(u0_u4__abc_44844_n588), .B(u0_u4__abc_44844_n586), .Y(u0_u4__abc_44844_n589) );
  OR2X2 OR2X2_216 ( .A(u0__abc_49347_n1392), .B(u0__abc_49347_n1394), .Y(u0__abc_49347_n1395) );
  OR2X2 OR2X2_2160 ( .A(u0_u4__abc_44844_n595), .B(u0_u4__abc_44844_n587), .Y(u0_u4__abc_44844_n596) );
  OR2X2 OR2X2_2161 ( .A(u0_u4__abc_44844_n601), .B(u0_u4__abc_44844_n599), .Y(u0_u4__abc_44844_n602) );
  OR2X2 OR2X2_2162 ( .A(u0_u4__abc_44844_n605), .B(u0_u4__abc_44844_n603), .Y(u0_u4__abc_44844_n606) );
  OR2X2 OR2X2_2163 ( .A(u0_u4__abc_44844_n611), .B(u0_u4__abc_44844_n604), .Y(u0_u4__abc_44844_n612) );
  OR2X2 OR2X2_2164 ( .A(u0_u4__abc_44844_n619), .B(u0_u4__abc_44844_n620), .Y(u0_u4__abc_44844_n621) );
  OR2X2 OR2X2_2165 ( .A(u0_u4__abc_44844_n623), .B(u0_u4__abc_44844_n618), .Y(u0_u4__abc_44844_n624) );
  OR2X2 OR2X2_2166 ( .A(u0_u4__abc_44844_n628), .B(u0_u4__abc_44844_n592), .Y(u0_u4__abc_44844_n629) );
  OR2X2 OR2X2_2167 ( .A(u0_u4__abc_44844_n632), .B(u0_u4__abc_44844_n630), .Y(u0_u4__abc_44844_n633) );
  OR2X2 OR2X2_2168 ( .A(u0_u4__abc_44844_n637), .B(u0_u4__abc_44844_n635), .Y(u0_u4__abc_44844_n638) );
  OR2X2 OR2X2_2169 ( .A(u0_u4__abc_44844_n639), .B(u0_u4__abc_44844_n631), .Y(u0_u4__abc_44844_n640) );
  OR2X2 OR2X2_217 ( .A(u0__abc_49347_n1203_bF_buf3), .B(u0_tms0_8_), .Y(u0__abc_49347_n1396) );
  OR2X2 OR2X2_2170 ( .A(u0_u4__abc_44844_n643), .B(u0_u4__abc_44844_n636), .Y(u0_u4__abc_44844_n644) );
  OR2X2 OR2X2_2171 ( .A(u0_csc5_2_), .B(u0_csc5_1_), .Y(u0_u5__abc_45296_n201_1) );
  OR2X2 OR2X2_2172 ( .A(u0_u5__abc_45296_n201_1), .B(u0_csc5_3_), .Y(u0_u5__abc_45296_n202_1) );
  OR2X2 OR2X2_2173 ( .A(u0_u5__abc_45296_n209), .B(u0_u5__abc_45296_n205_1), .Y(u0_u5_lmr_req_FF_INPUT) );
  OR2X2 OR2X2_2174 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf7), .B(u0_tms5_0_), .Y(u0_u5__abc_45296_n217_1) );
  OR2X2 OR2X2_2175 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf5), .B(u0_tms5_1_), .Y(u0_u5__abc_45296_n224) );
  OR2X2 OR2X2_2176 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf3), .B(u0_tms5_2_), .Y(u0_u5__abc_45296_n230) );
  OR2X2 OR2X2_2177 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf1), .B(u0_tms5_3_), .Y(u0_u5__abc_45296_n236) );
  OR2X2 OR2X2_2178 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf7), .B(u0_tms5_4_), .Y(u0_u5__abc_45296_n242) );
  OR2X2 OR2X2_2179 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf5), .B(u0_tms5_5_), .Y(u0_u5__abc_45296_n248) );
  OR2X2 OR2X2_218 ( .A(u0__abc_49347_n1398_1), .B(u0__abc_49347_n1376), .Y(u0_sp_tms_8__FF_INPUT) );
  OR2X2 OR2X2_2180 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf3), .B(u0_tms5_6_), .Y(u0_u5__abc_45296_n254) );
  OR2X2 OR2X2_2181 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf1), .B(u0_tms5_7_), .Y(u0_u5__abc_45296_n260_1) );
  OR2X2 OR2X2_2182 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf7), .B(u0_tms5_8_), .Y(u0_u5__abc_45296_n266_1) );
  OR2X2 OR2X2_2183 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf5), .B(u0_tms5_9_), .Y(u0_u5__abc_45296_n272) );
  OR2X2 OR2X2_2184 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf3), .B(u0_tms5_10_), .Y(u0_u5__abc_45296_n278) );
  OR2X2 OR2X2_2185 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf1), .B(u0_tms5_11_), .Y(u0_u5__abc_45296_n284) );
  OR2X2 OR2X2_2186 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf7), .B(u0_tms5_12_), .Y(u0_u5__abc_45296_n290) );
  OR2X2 OR2X2_2187 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf5), .B(u0_tms5_13_), .Y(u0_u5__abc_45296_n296_1) );
  OR2X2 OR2X2_2188 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf3), .B(u0_tms5_14_), .Y(u0_u5__abc_45296_n302) );
  OR2X2 OR2X2_2189 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf1), .B(u0_tms5_15_), .Y(u0_u5__abc_45296_n308) );
  OR2X2 OR2X2_219 ( .A(u0__abc_49347_n1183_1_bF_buf2), .B(1'b0), .Y(u0__abc_49347_n1402) );
  OR2X2 OR2X2_2190 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf7), .B(u0_tms5_16_), .Y(u0_u5__abc_45296_n314_1) );
  OR2X2 OR2X2_2191 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf5), .B(u0_tms5_17_), .Y(u0_u5__abc_45296_n320) );
  OR2X2 OR2X2_2192 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf3), .B(u0_tms5_18_), .Y(u0_u5__abc_45296_n326) );
  OR2X2 OR2X2_2193 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf1), .B(u0_tms5_19_), .Y(u0_u5__abc_45296_n332) );
  OR2X2 OR2X2_2194 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf7), .B(u0_tms5_20_), .Y(u0_u5__abc_45296_n338) );
  OR2X2 OR2X2_2195 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf5), .B(u0_tms5_21_), .Y(u0_u5__abc_45296_n344) );
  OR2X2 OR2X2_2196 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf3), .B(u0_tms5_22_), .Y(u0_u5__abc_45296_n350) );
  OR2X2 OR2X2_2197 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf1), .B(u0_tms5_23_), .Y(u0_u5__abc_45296_n356) );
  OR2X2 OR2X2_2198 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf7), .B(u0_tms5_24_), .Y(u0_u5__abc_45296_n362) );
  OR2X2 OR2X2_2199 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf5), .B(u0_tms5_25_), .Y(u0_u5__abc_45296_n368) );
  OR2X2 OR2X2_22 ( .A(_abc_55805_n245_1), .B(cs_need_rfr_4_), .Y(_abc_55805_n270) );
  OR2X2 OR2X2_220 ( .A(spec_req_cs_6_bF_buf5), .B(1'b0), .Y(u0__abc_49347_n1403) );
  OR2X2 OR2X2_2200 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf3), .B(u0_tms5_26_), .Y(u0_u5__abc_45296_n374) );
  OR2X2 OR2X2_2201 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf1), .B(u0_tms5_27_), .Y(u0_u5__abc_45296_n380) );
  OR2X2 OR2X2_2202 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf7), .B(u0_tms5_28_), .Y(u0_u5__abc_45296_n386) );
  OR2X2 OR2X2_2203 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf5), .B(u0_tms5_29_), .Y(u0_u5__abc_45296_n392) );
  OR2X2 OR2X2_2204 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf3), .B(u0_tms5_30_), .Y(u0_u5__abc_45296_n398) );
  OR2X2 OR2X2_2205 ( .A(u0_u5_lmr_req_we_FF_INPUT_bF_buf1), .B(u0_tms5_31_), .Y(u0_u5__abc_45296_n404) );
  OR2X2 OR2X2_2206 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf7), .B(u0_csc5_0_), .Y(u0_u5__abc_45296_n412) );
  OR2X2 OR2X2_2207 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf5), .B(u0_csc5_1_), .Y(u0_u5__abc_45296_n417) );
  OR2X2 OR2X2_2208 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf3), .B(u0_csc5_2_), .Y(u0_u5__abc_45296_n422) );
  OR2X2 OR2X2_2209 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf1), .B(u0_csc5_3_), .Y(u0_u5__abc_45296_n427) );
  OR2X2 OR2X2_221 ( .A(u0__abc_49347_n1405), .B(u0__abc_49347_n1401), .Y(u0__abc_49347_n1406) );
  OR2X2 OR2X2_2210 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf7), .B(u0_csc5_4_), .Y(u0_u5__abc_45296_n432) );
  OR2X2 OR2X2_2211 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf5), .B(u0_csc5_5_), .Y(u0_u5__abc_45296_n437) );
  OR2X2 OR2X2_2212 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf3), .B(u0_csc5_6_), .Y(u0_u5__abc_45296_n442) );
  OR2X2 OR2X2_2213 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf1), .B(u0_csc5_7_), .Y(u0_u5__abc_45296_n447) );
  OR2X2 OR2X2_2214 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf7), .B(u0_csc5_8_), .Y(u0_u5__abc_45296_n452) );
  OR2X2 OR2X2_2215 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf5), .B(u0_csc5_9_), .Y(u0_u5__abc_45296_n457) );
  OR2X2 OR2X2_2216 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf3), .B(u0_csc5_10_), .Y(u0_u5__abc_45296_n462) );
  OR2X2 OR2X2_2217 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf1), .B(u0_csc5_11_), .Y(u0_u5__abc_45296_n467) );
  OR2X2 OR2X2_2218 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf7), .B(u0_csc5_12_), .Y(u0_u5__abc_45296_n472) );
  OR2X2 OR2X2_2219 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf5), .B(u0_csc5_13_), .Y(u0_u5__abc_45296_n477) );
  OR2X2 OR2X2_222 ( .A(u0__abc_49347_n1407_1), .B(u0__abc_49347_n1408_1), .Y(u0__abc_49347_n1409) );
  OR2X2 OR2X2_2220 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf3), .B(u0_csc5_14_), .Y(u0_u5__abc_45296_n482) );
  OR2X2 OR2X2_2221 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf1), .B(u0_csc5_15_), .Y(u0_u5__abc_45296_n487) );
  OR2X2 OR2X2_2222 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf7), .B(u0_csc5_16_), .Y(u0_u5__abc_45296_n492) );
  OR2X2 OR2X2_2223 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf5), .B(u0_csc5_17_), .Y(u0_u5__abc_45296_n497) );
  OR2X2 OR2X2_2224 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf3), .B(u0_csc5_18_), .Y(u0_u5__abc_45296_n502) );
  OR2X2 OR2X2_2225 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf1), .B(u0_csc5_19_), .Y(u0_u5__abc_45296_n507) );
  OR2X2 OR2X2_2226 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf7), .B(u0_csc5_20_), .Y(u0_u5__abc_45296_n512) );
  OR2X2 OR2X2_2227 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf5), .B(u0_csc5_21_), .Y(u0_u5__abc_45296_n517) );
  OR2X2 OR2X2_2228 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf3), .B(u0_csc5_22_), .Y(u0_u5__abc_45296_n522) );
  OR2X2 OR2X2_2229 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf1), .B(u0_csc5_23_), .Y(u0_u5__abc_45296_n527) );
  OR2X2 OR2X2_223 ( .A(u0__abc_49347_n1410), .B(u0__abc_49347_n1411), .Y(u0__abc_49347_n1412) );
  OR2X2 OR2X2_2230 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf7), .B(u0_csc5_24_), .Y(u0_u5__abc_45296_n532) );
  OR2X2 OR2X2_2231 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf5), .B(u0_csc5_25_), .Y(u0_u5__abc_45296_n537) );
  OR2X2 OR2X2_2232 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf3), .B(u0_csc5_26_), .Y(u0_u5__abc_45296_n542) );
  OR2X2 OR2X2_2233 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf1), .B(u0_csc5_27_), .Y(u0_u5__abc_45296_n547) );
  OR2X2 OR2X2_2234 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf7), .B(u0_csc5_28_), .Y(u0_u5__abc_45296_n552) );
  OR2X2 OR2X2_2235 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf5), .B(u0_csc5_29_), .Y(u0_u5__abc_45296_n557) );
  OR2X2 OR2X2_2236 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf3), .B(u0_csc5_30_), .Y(u0_u5__abc_45296_n562) );
  OR2X2 OR2X2_2237 ( .A(u0_u5_init_req_we_FF_INPUT_bF_buf1), .B(u0_csc5_31_), .Y(u0_u5__abc_45296_n567) );
  OR2X2 OR2X2_2238 ( .A(u0_u5__abc_45296_n575), .B(u0_u5__abc_45296_n573), .Y(u0_u5__abc_45296_n576) );
  OR2X2 OR2X2_2239 ( .A(u0_u5__abc_45296_n579), .B(u0_u5__abc_45296_n577), .Y(u0_u5__abc_45296_n580) );
  OR2X2 OR2X2_224 ( .A(u0__abc_49347_n1413), .B(u0__abc_49347_n1414), .Y(u0__abc_49347_n1415) );
  OR2X2 OR2X2_2240 ( .A(u0_u5__abc_45296_n586), .B(u0_u5__abc_45296_n578), .Y(u0_u5__abc_45296_n587) );
  OR2X2 OR2X2_2241 ( .A(u0_u5__abc_45296_n592), .B(u0_u5__abc_45296_n590), .Y(u0_u5__abc_45296_n593) );
  OR2X2 OR2X2_2242 ( .A(u0_u5__abc_45296_n596), .B(u0_u5__abc_45296_n594), .Y(u0_u5__abc_45296_n597) );
  OR2X2 OR2X2_2243 ( .A(u0_u5__abc_45296_n602), .B(u0_u5__abc_45296_n595), .Y(u0_u5__abc_45296_n603) );
  OR2X2 OR2X2_2244 ( .A(u0_u5__abc_45296_n610), .B(u0_u5__abc_45296_n611), .Y(u0_u5__abc_45296_n612) );
  OR2X2 OR2X2_2245 ( .A(u0_u5__abc_45296_n614), .B(u0_u5__abc_45296_n609), .Y(u0_u5__abc_45296_n615) );
  OR2X2 OR2X2_2246 ( .A(u0_u5__abc_45296_n619), .B(u0_u5__abc_45296_n583), .Y(u0_u5__abc_45296_n620) );
  OR2X2 OR2X2_2247 ( .A(u0_u5__abc_45296_n623), .B(u0_u5__abc_45296_n621), .Y(u0_u5__abc_45296_n624) );
  OR2X2 OR2X2_2248 ( .A(u0_u5__abc_45296_n628), .B(u0_u5__abc_45296_n626), .Y(u0_u5__abc_45296_n629) );
  OR2X2 OR2X2_2249 ( .A(u0_u5__abc_45296_n630), .B(u0_u5__abc_45296_n622), .Y(u0_u5__abc_45296_n631) );
  OR2X2 OR2X2_225 ( .A(u0__abc_49347_n1417_1), .B(spec_req_cs_0_bF_buf5), .Y(u0__abc_49347_n1418) );
  OR2X2 OR2X2_2250 ( .A(u0_u5__abc_45296_n634), .B(u0_u5__abc_45296_n627), .Y(u0_u5__abc_45296_n635) );
  OR2X2 OR2X2_2251 ( .A(u0_u5_inited), .B(u0_init_ack5), .Y(u0_u5_inited_FF_INPUT) );
  OR2X2 OR2X2_2252 ( .A(u0_u5__abc_45296_n648), .B(u0_u5__abc_45296_n644), .Y(u0_u5_init_req_FF_INPUT) );
  OR2X2 OR2X2_2253 ( .A(csc_s_4_), .B(csc_s_5_bF_buf4), .Y(u1__abc_45852_n260_1) );
  OR2X2 OR2X2_2254 ( .A(u1__abc_45852_n262_1), .B(u1__abc_45852_n265_1), .Y(page_size_10_) );
  OR2X2 OR2X2_2255 ( .A(u1__abc_45852_n263), .B(csc_s_7_), .Y(u1__abc_45852_n268) );
  OR2X2 OR2X2_2256 ( .A(u1__abc_45852_n269), .B(csc_s_5_bF_buf3), .Y(u1__abc_45852_n270) );
  OR2X2 OR2X2_2257 ( .A(u1__abc_45852_n268), .B(u1__abc_45852_n270), .Y(u1__abc_45852_n271_1) );
  OR2X2 OR2X2_2258 ( .A(csc_s_7_), .B(csc_s_6_), .Y(u1__abc_45852_n272_1) );
  OR2X2 OR2X2_2259 ( .A(u1__abc_45852_n260_1), .B(u1__abc_45852_n272_1), .Y(u1__abc_45852_n273_1) );
  OR2X2 OR2X2_226 ( .A(u0__abc_49347_n1416_1), .B(u0__abc_49347_n1418), .Y(u0__abc_49347_n1419) );
  OR2X2 OR2X2_2260 ( .A(u1__abc_45852_n285_1), .B(u1__abc_45852_n286_1), .Y(u1__abc_45852_n287_1) );
  OR2X2 OR2X2_2261 ( .A(u1__abc_45852_n287_1), .B(u1__abc_45852_n283), .Y(u1__abc_45852_n288) );
  OR2X2 OR2X2_2262 ( .A(u1__abc_45852_n288), .B(u1_bas), .Y(u1__abc_45852_n289) );
  OR2X2 OR2X2_2263 ( .A(u1__abc_45852_n295), .B(u1__abc_45852_n294_1), .Y(u1__abc_45852_n296) );
  OR2X2 OR2X2_2264 ( .A(u1__abc_45852_n296), .B(u1__abc_45852_n293_1), .Y(u1__abc_45852_n297) );
  OR2X2 OR2X2_2265 ( .A(u1__abc_45852_n262_1), .B(u1__abc_45852_n277), .Y(u1__abc_45852_n303) );
  OR2X2 OR2X2_2266 ( .A(u1__abc_45852_n305), .B(u1__abc_45852_n306_1), .Y(u1__abc_45852_n307_1) );
  OR2X2 OR2X2_2267 ( .A(u1__abc_45852_n307_1), .B(u1__abc_45852_n304), .Y(u1__abc_45852_n308_1) );
  OR2X2 OR2X2_2268 ( .A(u1__abc_45852_n308_1), .B(u1__abc_45852_n302), .Y(u1__abc_45852_n309) );
  OR2X2 OR2X2_2269 ( .A(u1__abc_45852_n301_1), .B(u1__abc_45852_n309), .Y(u1__abc_45852_n310) );
  OR2X2 OR2X2_227 ( .A(u0__abc_49347_n1203_bF_buf2), .B(u0_tms0_9_), .Y(u0__abc_49347_n1420) );
  OR2X2 OR2X2_2270 ( .A(u1__abc_45852_n310), .B(u1__abc_45852_n290), .Y(u1__abc_45852_n311) );
  OR2X2 OR2X2_2271 ( .A(u1__abc_45852_n313_1), .B(u1__abc_45852_n282), .Y(u1_bank_adr_0__FF_INPUT) );
  OR2X2 OR2X2_2272 ( .A(u1__abc_45852_n317), .B(u1__abc_45852_n318), .Y(u1__abc_45852_n319) );
  OR2X2 OR2X2_2273 ( .A(u1__abc_45852_n319), .B(u1__abc_45852_n316), .Y(u1__abc_45852_n320_1) );
  OR2X2 OR2X2_2274 ( .A(u1__abc_45852_n320_1), .B(u1_bas), .Y(u1__abc_45852_n321_1) );
  OR2X2 OR2X2_2275 ( .A(u1__abc_45852_n325), .B(u1__abc_45852_n326), .Y(u1__abc_45852_n327_1) );
  OR2X2 OR2X2_2276 ( .A(u1__abc_45852_n327_1), .B(u1__abc_45852_n324), .Y(u1__abc_45852_n328_1) );
  OR2X2 OR2X2_2277 ( .A(u1__abc_45852_n328_1), .B(u1__abc_45852_n323), .Y(u1__abc_45852_n329_1) );
  OR2X2 OR2X2_2278 ( .A(u1__abc_45852_n322_1), .B(u1__abc_45852_n329_1), .Y(u1__abc_45852_n330) );
  OR2X2 OR2X2_2279 ( .A(u1__abc_45852_n330), .B(u1__abc_45852_n290), .Y(u1__abc_45852_n331) );
  OR2X2 OR2X2_228 ( .A(u0__abc_49347_n1422), .B(u0__abc_49347_n1400), .Y(u0_sp_tms_9__FF_INPUT) );
  OR2X2 OR2X2_2280 ( .A(u1__abc_45852_n333_1), .B(u1__abc_45852_n315_1), .Y(u1_bank_adr_1__FF_INPUT) );
  OR2X2 OR2X2_2281 ( .A(u1__abc_45852_n338), .B(u1__abc_45852_n337), .Y(u1__abc_45852_n339_1) );
  OR2X2 OR2X2_2282 ( .A(u1__abc_45852_n339_1), .B(u1__abc_45852_n336), .Y(u1__abc_45852_n340_1) );
  OR2X2 OR2X2_2283 ( .A(u1__abc_45852_n340_1), .B(u1_bas), .Y(u1__abc_45852_n341_1) );
  OR2X2 OR2X2_2284 ( .A(u1__abc_45852_n288), .B(u1__abc_45852_n290), .Y(u1__abc_45852_n342) );
  OR2X2 OR2X2_2285 ( .A(u1__abc_45852_n344), .B(u1__abc_45852_n335_1), .Y(u1_row_adr_0__FF_INPUT) );
  OR2X2 OR2X2_2286 ( .A(u1__abc_45852_n349), .B(u1__abc_45852_n348), .Y(u1__abc_45852_n350) );
  OR2X2 OR2X2_2287 ( .A(u1__abc_45852_n350), .B(u1__abc_45852_n347_1), .Y(u1__abc_45852_n351_1) );
  OR2X2 OR2X2_2288 ( .A(u1__abc_45852_n351_1), .B(u1_bas), .Y(u1__abc_45852_n352_1) );
  OR2X2 OR2X2_2289 ( .A(u1__abc_45852_n320_1), .B(u1__abc_45852_n290), .Y(u1__abc_45852_n353_1) );
  OR2X2 OR2X2_229 ( .A(u0__abc_49347_n1183_1_bF_buf1), .B(1'b0), .Y(u0__abc_49347_n1426_1) );
  OR2X2 OR2X2_2290 ( .A(u1__abc_45852_n355), .B(u1__abc_45852_n346_1), .Y(u1_row_adr_1__FF_INPUT) );
  OR2X2 OR2X2_2291 ( .A(u1__abc_45852_n362), .B(u1__abc_45852_n361), .Y(u1__abc_45852_n363_1) );
  OR2X2 OR2X2_2292 ( .A(u1__abc_45852_n364_1), .B(u1__abc_45852_n360), .Y(u1__abc_45852_n365_1) );
  OR2X2 OR2X2_2293 ( .A(u1__abc_45852_n367), .B(u1__abc_45852_n368), .Y(u1__abc_45852_n369_1) );
  OR2X2 OR2X2_2294 ( .A(u1__abc_45852_n366), .B(u1__abc_45852_n369_1), .Y(u1__abc_45852_n370_1) );
  OR2X2 OR2X2_2295 ( .A(u1__abc_45852_n365_1), .B(u1__abc_45852_n370_1), .Y(u1__abc_45852_n371_1) );
  OR2X2 OR2X2_2296 ( .A(u1__abc_45852_n359_1), .B(u1__abc_45852_n371_1), .Y(u1__abc_45852_n372) );
  OR2X2 OR2X2_2297 ( .A(u1__abc_45852_n372), .B(u1_bas), .Y(u1__abc_45852_n373) );
  OR2X2 OR2X2_2298 ( .A(u1__abc_45852_n340_1), .B(u1__abc_45852_n290), .Y(u1__abc_45852_n374) );
  OR2X2 OR2X2_2299 ( .A(u1__abc_45852_n376_1), .B(u1__abc_45852_n357_1), .Y(u1_row_adr_2__FF_INPUT) );
  OR2X2 OR2X2_23 ( .A(_abc_55805_n240_bF_buf0), .B(spec_req_cs_5_bF_buf5), .Y(_abc_55805_n272) );
  OR2X2 OR2X2_230 ( .A(spec_req_cs_6_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n1427) );
  OR2X2 OR2X2_2300 ( .A(u1__abc_45852_n382_1), .B(u1__abc_45852_n381_1), .Y(u1__abc_45852_n383_1) );
  OR2X2 OR2X2_2301 ( .A(u1__abc_45852_n383_1), .B(u1__abc_45852_n380), .Y(u1__abc_45852_n384) );
  OR2X2 OR2X2_2302 ( .A(u1__abc_45852_n384), .B(u1__abc_45852_n379), .Y(u1__abc_45852_n385) );
  OR2X2 OR2X2_2303 ( .A(u1__abc_45852_n385), .B(u1_bas), .Y(u1__abc_45852_n386) );
  OR2X2 OR2X2_2304 ( .A(u1__abc_45852_n351_1), .B(u1__abc_45852_n290), .Y(u1__abc_45852_n387_1) );
  OR2X2 OR2X2_2305 ( .A(u1__abc_45852_n389_1), .B(u1__abc_45852_n378), .Y(u1_row_adr_3__FF_INPUT) );
  OR2X2 OR2X2_2306 ( .A(u1__abc_45852_n394_1), .B(u1__abc_45852_n393_1), .Y(u1__abc_45852_n395_1) );
  OR2X2 OR2X2_2307 ( .A(u1__abc_45852_n397), .B(u1__abc_45852_n398), .Y(u1__abc_45852_n399_1) );
  OR2X2 OR2X2_2308 ( .A(u1__abc_45852_n396), .B(u1__abc_45852_n399_1), .Y(u1__abc_45852_n400_1) );
  OR2X2 OR2X2_2309 ( .A(u1__abc_45852_n395_1), .B(u1__abc_45852_n400_1), .Y(u1__abc_45852_n401_1) );
  OR2X2 OR2X2_231 ( .A(u0__abc_49347_n1429), .B(u0__abc_49347_n1425_1), .Y(u0__abc_49347_n1430) );
  OR2X2 OR2X2_2310 ( .A(u1__abc_45852_n392), .B(u1__abc_45852_n401_1), .Y(u1__abc_45852_n402) );
  OR2X2 OR2X2_2311 ( .A(u1__abc_45852_n402), .B(u1_bas), .Y(u1__abc_45852_n403) );
  OR2X2 OR2X2_2312 ( .A(u1__abc_45852_n372), .B(u1__abc_45852_n290), .Y(u1__abc_45852_n404) );
  OR2X2 OR2X2_2313 ( .A(u1__abc_45852_n406_1), .B(u1__abc_45852_n391), .Y(u1_row_adr_4__FF_INPUT) );
  OR2X2 OR2X2_2314 ( .A(u1__abc_45852_n385), .B(u1__abc_45852_n290), .Y(u1__abc_45852_n409) );
  OR2X2 OR2X2_2315 ( .A(u1__abc_45852_n412_1), .B(u1__abc_45852_n411_1), .Y(u1__abc_45852_n413_1) );
  OR2X2 OR2X2_2316 ( .A(u1__abc_45852_n415), .B(u1__abc_45852_n416), .Y(u1__abc_45852_n417_1) );
  OR2X2 OR2X2_2317 ( .A(u1__abc_45852_n414), .B(u1__abc_45852_n417_1), .Y(u1__abc_45852_n418_1) );
  OR2X2 OR2X2_2318 ( .A(u1__abc_45852_n413_1), .B(u1__abc_45852_n418_1), .Y(u1__abc_45852_n419_1) );
  OR2X2 OR2X2_2319 ( .A(u1__abc_45852_n410), .B(u1__abc_45852_n419_1), .Y(u1__abc_45852_n420_1) );
  OR2X2 OR2X2_232 ( .A(u0__abc_49347_n1431), .B(u0__abc_49347_n1432), .Y(u0__abc_49347_n1433) );
  OR2X2 OR2X2_2320 ( .A(u1__abc_45852_n420_1), .B(u1_bas), .Y(u1__abc_45852_n421_1) );
  OR2X2 OR2X2_2321 ( .A(u1__abc_45852_n423_1), .B(u1__abc_45852_n408), .Y(u1_row_adr_5__FF_INPUT) );
  OR2X2 OR2X2_2322 ( .A(u1__abc_45852_n428_1), .B(u1__abc_45852_n427_1), .Y(u1__abc_45852_n429_1) );
  OR2X2 OR2X2_2323 ( .A(u1__abc_45852_n429_1), .B(u1__abc_45852_n426_1), .Y(u1__abc_45852_n430_1) );
  OR2X2 OR2X2_2324 ( .A(u1__abc_45852_n430_1), .B(u1_bas), .Y(u1__abc_45852_n431_1) );
  OR2X2 OR2X2_2325 ( .A(u1__abc_45852_n402), .B(u1__abc_45852_n290), .Y(u1__abc_45852_n432_1) );
  OR2X2 OR2X2_2326 ( .A(u1__abc_45852_n434_1), .B(u1__abc_45852_n425_1), .Y(u1_row_adr_6__FF_INPUT) );
  OR2X2 OR2X2_2327 ( .A(u1__abc_45852_n420_1), .B(u1__abc_45852_n290), .Y(u1__abc_45852_n437_1) );
  OR2X2 OR2X2_2328 ( .A(u1__abc_45852_n440_1), .B(u1__abc_45852_n439_1), .Y(u1__abc_45852_n441_1) );
  OR2X2 OR2X2_2329 ( .A(u1__abc_45852_n441_1), .B(u1__abc_45852_n438_1), .Y(u1__abc_45852_n442_1) );
  OR2X2 OR2X2_233 ( .A(u0__abc_49347_n1434_1), .B(u0__abc_49347_n1435_1), .Y(u0__abc_49347_n1436) );
  OR2X2 OR2X2_2330 ( .A(u1__abc_45852_n442_1), .B(u1_bas), .Y(u1__abc_45852_n443_1) );
  OR2X2 OR2X2_2331 ( .A(u1__abc_45852_n445_1), .B(u1__abc_45852_n436_1), .Y(u1_row_adr_7__FF_INPUT) );
  OR2X2 OR2X2_2332 ( .A(u1__abc_45852_n451_1), .B(u1__abc_45852_n450_1), .Y(u1__abc_45852_n452_1) );
  OR2X2 OR2X2_2333 ( .A(u1__abc_45852_n452_1), .B(u1__abc_45852_n449_1), .Y(u1__abc_45852_n453_1) );
  OR2X2 OR2X2_2334 ( .A(u1__abc_45852_n453_1), .B(u1__abc_45852_n448_1), .Y(u1__abc_45852_n454_1) );
  OR2X2 OR2X2_2335 ( .A(u1__abc_45852_n454_1), .B(u1_bas), .Y(u1__abc_45852_n455_1) );
  OR2X2 OR2X2_2336 ( .A(u1__abc_45852_n430_1), .B(u1__abc_45852_n290), .Y(u1__abc_45852_n456_1) );
  OR2X2 OR2X2_2337 ( .A(u1__abc_45852_n458_1), .B(u1__abc_45852_n447_1), .Y(u1_row_adr_8__FF_INPUT) );
  OR2X2 OR2X2_2338 ( .A(u1__abc_45852_n442_1), .B(u1__abc_45852_n290), .Y(u1__abc_45852_n461_1) );
  OR2X2 OR2X2_2339 ( .A(u1__abc_45852_n464_1), .B(u1__abc_45852_n465_1), .Y(u1__abc_45852_n466_1) );
  OR2X2 OR2X2_234 ( .A(u0__abc_49347_n1437), .B(u0__abc_49347_n1438), .Y(u0__abc_49347_n1439) );
  OR2X2 OR2X2_2340 ( .A(u1__abc_45852_n463_1), .B(u1__abc_45852_n466_1), .Y(u1__abc_45852_n467) );
  OR2X2 OR2X2_2341 ( .A(u1__abc_45852_n306_1), .B(u1_bas), .Y(u1__abc_45852_n468_1) );
  OR2X2 OR2X2_2342 ( .A(u1__abc_45852_n467), .B(u1__abc_45852_n468_1), .Y(u1__abc_45852_n469) );
  OR2X2 OR2X2_2343 ( .A(u1__abc_45852_n469), .B(u1__abc_45852_n462_1), .Y(u1__abc_45852_n470_1) );
  OR2X2 OR2X2_2344 ( .A(u1__abc_45852_n472_1), .B(u1__abc_45852_n460_1), .Y(u1_row_adr_9__FF_INPUT) );
  OR2X2 OR2X2_2345 ( .A(u1__abc_45852_n454_1), .B(u1__abc_45852_n290), .Y(u1__abc_45852_n475) );
  OR2X2 OR2X2_2346 ( .A(u1__abc_45852_n326), .B(u1_bas), .Y(u1__abc_45852_n479) );
  OR2X2 OR2X2_2347 ( .A(u1__abc_45852_n479), .B(u1__abc_45852_n478), .Y(u1__abc_45852_n480) );
  OR2X2 OR2X2_2348 ( .A(u1__abc_45852_n481), .B(u1__abc_45852_n302), .Y(u1__abc_45852_n482) );
  OR2X2 OR2X2_2349 ( .A(u1__abc_45852_n482), .B(u1__abc_45852_n483_1), .Y(u1__abc_45852_n484) );
  OR2X2 OR2X2_235 ( .A(u0__abc_49347_n1441), .B(spec_req_cs_0_bF_buf4), .Y(u0__abc_49347_n1442) );
  OR2X2 OR2X2_2350 ( .A(u1__abc_45852_n484), .B(u1__abc_45852_n480), .Y(u1__abc_45852_n485) );
  OR2X2 OR2X2_2351 ( .A(u1__abc_45852_n485), .B(u1__abc_45852_n476_1), .Y(u1__abc_45852_n486) );
  OR2X2 OR2X2_2352 ( .A(u1__abc_45852_n488_1), .B(u1__abc_45852_n474_1), .Y(u1_row_adr_10__FF_INPUT) );
  OR2X2 OR2X2_2353 ( .A(u1__abc_45852_n467), .B(u1__abc_45852_n290), .Y(u1__abc_45852_n491) );
  OR2X2 OR2X2_2354 ( .A(u1__abc_45852_n491), .B(u1__abc_45852_n462_1), .Y(u1__abc_45852_n492) );
  OR2X2 OR2X2_2355 ( .A(u1__abc_45852_n324), .B(u1_bas), .Y(u1__abc_45852_n496_1) );
  OR2X2 OR2X2_2356 ( .A(u1__abc_45852_n496_1), .B(u1__abc_45852_n495), .Y(u1__abc_45852_n497) );
  OR2X2 OR2X2_2357 ( .A(u1__abc_45852_n497), .B(u1__abc_45852_n494_1), .Y(u1__abc_45852_n498) );
  OR2X2 OR2X2_2358 ( .A(u1__abc_45852_n498), .B(u1__abc_45852_n493), .Y(u1__abc_45852_n499) );
  OR2X2 OR2X2_2359 ( .A(u1__abc_45852_n501), .B(u1__abc_45852_n490_1), .Y(u1_row_adr_11__FF_INPUT) );
  OR2X2 OR2X2_236 ( .A(u0__abc_49347_n1440), .B(u0__abc_49347_n1442), .Y(u0__abc_49347_n1443_1) );
  OR2X2 OR2X2_2360 ( .A(u1__abc_45852_n478), .B(u1__abc_45852_n290), .Y(u1__abc_45852_n505) );
  OR2X2 OR2X2_2361 ( .A(u1__abc_45852_n505), .B(u1__abc_45852_n504), .Y(u1__abc_45852_n506_1) );
  OR2X2 OR2X2_2362 ( .A(u1__abc_45852_n476_1), .B(u1__abc_45852_n506_1), .Y(u1__abc_45852_n507) );
  OR2X2 OR2X2_2363 ( .A(u1__abc_45852_n325), .B(u1_bas), .Y(u1__abc_45852_n510) );
  OR2X2 OR2X2_2364 ( .A(u1__abc_45852_n510), .B(u1__abc_45852_n509), .Y(u1__abc_45852_n511) );
  OR2X2 OR2X2_2365 ( .A(u1__abc_45852_n508_1), .B(u1__abc_45852_n511), .Y(u1__abc_45852_n512_1) );
  OR2X2 OR2X2_2366 ( .A(u1__abc_45852_n514_1), .B(u1__abc_45852_n503), .Y(u1_row_adr_12__FF_INPUT) );
  OR2X2 OR2X2_2367 ( .A(u1__abc_45852_n517), .B(u1__abc_45852_n518_1), .Y(u1__abc_45852_n519) );
  OR2X2 OR2X2_2368 ( .A(u1__abc_45852_n520_1), .B(\wb_addr_i[2] ), .Y(u1__abc_45852_n521) );
  OR2X2 OR2X2_2369 ( .A(u1__abc_45852_n519), .B(u1_col_adr_0_), .Y(u1__abc_45852_n522) );
  OR2X2 OR2X2_237 ( .A(u0__abc_49347_n1203_bF_buf1), .B(u0_tms0_10_), .Y(u0__abc_49347_n1444_1) );
  OR2X2 OR2X2_2370 ( .A(u1__abc_45852_n520_1), .B(\wb_addr_i[3] ), .Y(u1__abc_45852_n524_1) );
  OR2X2 OR2X2_2371 ( .A(u1__abc_45852_n519), .B(u1_col_adr_1_), .Y(u1__abc_45852_n525) );
  OR2X2 OR2X2_2372 ( .A(u1__abc_45852_n520_1), .B(\wb_addr_i[4] ), .Y(u1__abc_45852_n527) );
  OR2X2 OR2X2_2373 ( .A(u1__abc_45852_n519), .B(u1_col_adr_2_), .Y(u1__abc_45852_n528) );
  OR2X2 OR2X2_2374 ( .A(u1__abc_45852_n520_1), .B(\wb_addr_i[5] ), .Y(u1__abc_45852_n530_1) );
  OR2X2 OR2X2_2375 ( .A(u1__abc_45852_n519), .B(u1_col_adr_3_), .Y(u1__abc_45852_n531) );
  OR2X2 OR2X2_2376 ( .A(u1__abc_45852_n520_1), .B(\wb_addr_i[6] ), .Y(u1__abc_45852_n533) );
  OR2X2 OR2X2_2377 ( .A(u1__abc_45852_n519), .B(u1_col_adr_4_), .Y(u1__abc_45852_n534) );
  OR2X2 OR2X2_2378 ( .A(u1__abc_45852_n520_1), .B(\wb_addr_i[7] ), .Y(u1__abc_45852_n536_1) );
  OR2X2 OR2X2_2379 ( .A(u1__abc_45852_n519), .B(u1_col_adr_5_), .Y(u1__abc_45852_n537) );
  OR2X2 OR2X2_238 ( .A(u0__abc_49347_n1446), .B(u0__abc_49347_n1424), .Y(u0_sp_tms_10__FF_INPUT) );
  OR2X2 OR2X2_2380 ( .A(u1__abc_45852_n520_1), .B(\wb_addr_i[8] ), .Y(u1__abc_45852_n539) );
  OR2X2 OR2X2_2381 ( .A(u1__abc_45852_n519), .B(u1_col_adr_6_), .Y(u1__abc_45852_n540) );
  OR2X2 OR2X2_2382 ( .A(u1__abc_45852_n520_1), .B(\wb_addr_i[9] ), .Y(u1__abc_45852_n542_1) );
  OR2X2 OR2X2_2383 ( .A(u1__abc_45852_n519), .B(u1_col_adr_7_), .Y(u1__abc_45852_n543) );
  OR2X2 OR2X2_2384 ( .A(u1__abc_45852_n548_1), .B(u1__abc_45852_n545), .Y(u1_col_adr_8__FF_INPUT) );
  OR2X2 OR2X2_2385 ( .A(u1__abc_45852_n552), .B(u1__abc_45852_n550_1), .Y(u1_col_adr_9__FF_INPUT) );
  OR2X2 OR2X2_2386 ( .A(cs_le_bF_buf3), .B(wb_we_i), .Y(u1__abc_45852_n554_1) );
  OR2X2 OR2X2_2387 ( .A(u1_acs_addr_0_), .B(next_adr_bF_buf4), .Y(u1__abc_45852_n555) );
  OR2X2 OR2X2_2388 ( .A(u1__abc_45852_n556_bF_buf3), .B(u1_acs_addr_pl1_0_), .Y(u1__abc_45852_n557_1) );
  OR2X2 OR2X2_2389 ( .A(u1__abc_45852_n558), .B(u1__abc_45852_n554_1_bF_buf4), .Y(u1__abc_45852_n559) );
  OR2X2 OR2X2_239 ( .A(u0__abc_49347_n1183_1_bF_buf0), .B(1'b0), .Y(u0__abc_49347_n1450) );
  OR2X2 OR2X2_2390 ( .A(u1__abc_45852_n562_bF_buf3), .B(u1__abc_45852_n563), .Y(u1__abc_45852_n564_1) );
  OR2X2 OR2X2_2391 ( .A(u1__abc_45852_n564_1), .B(u1__abc_45852_n561), .Y(u1__abc_45852_n565) );
  OR2X2 OR2X2_2392 ( .A(u1__abc_45852_n565), .B(u1__abc_45852_n560_1), .Y(u1__abc_45852_n566) );
  OR2X2 OR2X2_2393 ( .A(next_adr_bF_buf2), .B(u1_acs_addr_1_), .Y(u1__abc_45852_n568) );
  OR2X2 OR2X2_2394 ( .A(u1__abc_45852_n556_bF_buf2), .B(u1_acs_addr_pl1_1_), .Y(u1__abc_45852_n569) );
  OR2X2 OR2X2_2395 ( .A(u1__abc_45852_n570_1), .B(u1__abc_45852_n554_1_bF_buf2), .Y(u1__abc_45852_n571) );
  OR2X2 OR2X2_2396 ( .A(u1__abc_45852_n562_bF_buf2), .B(u1__abc_45852_n574), .Y(u1__abc_45852_n575) );
  OR2X2 OR2X2_2397 ( .A(u1__abc_45852_n575), .B(u1__abc_45852_n573_1), .Y(u1__abc_45852_n576_1) );
  OR2X2 OR2X2_2398 ( .A(u1__abc_45852_n576_1), .B(u1__abc_45852_n572), .Y(u1__abc_45852_n577) );
  OR2X2 OR2X2_2399 ( .A(next_adr_bF_buf1), .B(u1_acs_addr_2_), .Y(u1__abc_45852_n579_1) );
  OR2X2 OR2X2_24 ( .A(lmr_sel_bF_buf1), .B(cs_5_), .Y(_abc_55805_n273) );
  OR2X2 OR2X2_240 ( .A(spec_req_cs_6_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n1451) );
  OR2X2 OR2X2_2400 ( .A(u1__abc_45852_n556_bF_buf1), .B(u1_acs_addr_pl1_2_), .Y(u1__abc_45852_n580) );
  OR2X2 OR2X2_2401 ( .A(u1__abc_45852_n581), .B(u1__abc_45852_n554_1_bF_buf1), .Y(u1__abc_45852_n582_1) );
  OR2X2 OR2X2_2402 ( .A(u1__abc_45852_n562_bF_buf1), .B(u1__abc_45852_n585_1), .Y(u1__abc_45852_n586) );
  OR2X2 OR2X2_2403 ( .A(u1__abc_45852_n586), .B(u1__abc_45852_n584), .Y(u1__abc_45852_n587) );
  OR2X2 OR2X2_2404 ( .A(u1__abc_45852_n587), .B(u1__abc_45852_n583), .Y(u1__abc_45852_n588_1) );
  OR2X2 OR2X2_2405 ( .A(next_adr_bF_buf0), .B(u1_acs_addr_3_), .Y(u1__abc_45852_n590_1) );
  OR2X2 OR2X2_2406 ( .A(u1__abc_45852_n556_bF_buf0), .B(u1_acs_addr_pl1_3_), .Y(u1__abc_45852_n591) );
  OR2X2 OR2X2_2407 ( .A(u1__abc_45852_n592), .B(u1__abc_45852_n554_1_bF_buf0), .Y(u1__abc_45852_n593) );
  OR2X2 OR2X2_2408 ( .A(u1__abc_45852_n562_bF_buf0), .B(u1__abc_45852_n596), .Y(u1__abc_45852_n597_1) );
  OR2X2 OR2X2_2409 ( .A(u1__abc_45852_n597_1), .B(u1__abc_45852_n595_1), .Y(u1__abc_45852_n598) );
  OR2X2 OR2X2_241 ( .A(u0__abc_49347_n1453_1), .B(u0__abc_49347_n1449), .Y(u0__abc_49347_n1454) );
  OR2X2 OR2X2_2410 ( .A(u1__abc_45852_n598), .B(u1__abc_45852_n594), .Y(u1__abc_45852_n599_1) );
  OR2X2 OR2X2_2411 ( .A(next_adr_bF_buf4), .B(u1_acs_addr_4_), .Y(u1__abc_45852_n601_1) );
  OR2X2 OR2X2_2412 ( .A(u1__abc_45852_n556_bF_buf3), .B(u1_acs_addr_pl1_4_), .Y(u1__abc_45852_n602) );
  OR2X2 OR2X2_2413 ( .A(u1__abc_45852_n603), .B(u1__abc_45852_n554_1_bF_buf4), .Y(u1__abc_45852_n604) );
  OR2X2 OR2X2_2414 ( .A(u1__abc_45852_n562_bF_buf3), .B(u1__abc_45852_n607), .Y(u1__abc_45852_n608) );
  OR2X2 OR2X2_2415 ( .A(u1__abc_45852_n608), .B(u1__abc_45852_n606), .Y(u1__abc_45852_n609) );
  OR2X2 OR2X2_2416 ( .A(u1__abc_45852_n609), .B(u1__abc_45852_n605), .Y(u1__abc_45852_n610) );
  OR2X2 OR2X2_2417 ( .A(next_adr_bF_buf3), .B(u1_acs_addr_5_), .Y(u1__abc_45852_n612) );
  OR2X2 OR2X2_2418 ( .A(u1__abc_45852_n556_bF_buf2), .B(u1_acs_addr_pl1_5_), .Y(u1__abc_45852_n613) );
  OR2X2 OR2X2_2419 ( .A(u1__abc_45852_n614), .B(u1__abc_45852_n554_1_bF_buf3), .Y(u1__abc_45852_n615) );
  OR2X2 OR2X2_242 ( .A(u0__abc_49347_n1455), .B(u0__abc_49347_n1456), .Y(u0__abc_49347_n1457) );
  OR2X2 OR2X2_2420 ( .A(u1__abc_45852_n562_bF_buf2), .B(u1__abc_45852_n618), .Y(u1__abc_45852_n619) );
  OR2X2 OR2X2_2421 ( .A(u1__abc_45852_n619), .B(u1__abc_45852_n617), .Y(u1__abc_45852_n620) );
  OR2X2 OR2X2_2422 ( .A(u1__abc_45852_n620), .B(u1__abc_45852_n616), .Y(u1__abc_45852_n621) );
  OR2X2 OR2X2_2423 ( .A(next_adr_bF_buf2), .B(u1_acs_addr_6_), .Y(u1__abc_45852_n623) );
  OR2X2 OR2X2_2424 ( .A(u1__abc_45852_n556_bF_buf1), .B(u1_acs_addr_pl1_6_), .Y(u1__abc_45852_n624) );
  OR2X2 OR2X2_2425 ( .A(u1__abc_45852_n625), .B(u1__abc_45852_n554_1_bF_buf2), .Y(u1__abc_45852_n626) );
  OR2X2 OR2X2_2426 ( .A(u1__abc_45852_n562_bF_buf1), .B(u1__abc_45852_n629), .Y(u1__abc_45852_n630) );
  OR2X2 OR2X2_2427 ( .A(u1__abc_45852_n630), .B(u1__abc_45852_n628), .Y(u1__abc_45852_n631) );
  OR2X2 OR2X2_2428 ( .A(u1__abc_45852_n631), .B(u1__abc_45852_n627), .Y(u1__abc_45852_n632) );
  OR2X2 OR2X2_2429 ( .A(next_adr_bF_buf1), .B(u1_acs_addr_7_), .Y(u1__abc_45852_n634) );
  OR2X2 OR2X2_243 ( .A(u0__abc_49347_n1458), .B(u0__abc_49347_n1459), .Y(u0__abc_49347_n1460) );
  OR2X2 OR2X2_2430 ( .A(u1__abc_45852_n556_bF_buf0), .B(u1_acs_addr_pl1_7_), .Y(u1__abc_45852_n635) );
  OR2X2 OR2X2_2431 ( .A(u1__abc_45852_n636), .B(u1__abc_45852_n554_1_bF_buf1), .Y(u1__abc_45852_n637) );
  OR2X2 OR2X2_2432 ( .A(u1__abc_45852_n562_bF_buf0), .B(u1__abc_45852_n640), .Y(u1__abc_45852_n641) );
  OR2X2 OR2X2_2433 ( .A(u1__abc_45852_n641), .B(u1__abc_45852_n639), .Y(u1__abc_45852_n642) );
  OR2X2 OR2X2_2434 ( .A(u1__abc_45852_n642), .B(u1__abc_45852_n638), .Y(u1__abc_45852_n643) );
  OR2X2 OR2X2_2435 ( .A(next_adr_bF_buf0), .B(u1_acs_addr_8_), .Y(u1__abc_45852_n645) );
  OR2X2 OR2X2_2436 ( .A(u1__abc_45852_n556_bF_buf3), .B(u1_acs_addr_pl1_8_), .Y(u1__abc_45852_n646) );
  OR2X2 OR2X2_2437 ( .A(u1__abc_45852_n647), .B(u1__abc_45852_n554_1_bF_buf0), .Y(u1__abc_45852_n648) );
  OR2X2 OR2X2_2438 ( .A(u1__abc_45852_n562_bF_buf3), .B(u1__abc_45852_n651), .Y(u1__abc_45852_n652) );
  OR2X2 OR2X2_2439 ( .A(u1__abc_45852_n652), .B(u1__abc_45852_n650), .Y(u1__abc_45852_n653) );
  OR2X2 OR2X2_244 ( .A(u0__abc_49347_n1461_1), .B(u0__abc_49347_n1462_1), .Y(u0__abc_49347_n1463) );
  OR2X2 OR2X2_2440 ( .A(u1__abc_45852_n653), .B(u1__abc_45852_n649), .Y(u1__abc_45852_n654) );
  OR2X2 OR2X2_2441 ( .A(next_adr_bF_buf4), .B(u1_acs_addr_9_), .Y(u1__abc_45852_n656) );
  OR2X2 OR2X2_2442 ( .A(u1__abc_45852_n556_bF_buf2), .B(u1_acs_addr_pl1_9_), .Y(u1__abc_45852_n657) );
  OR2X2 OR2X2_2443 ( .A(u1__abc_45852_n658), .B(u1__abc_45852_n554_1_bF_buf4), .Y(u1__abc_45852_n659) );
  OR2X2 OR2X2_2444 ( .A(u1__abc_45852_n562_bF_buf2), .B(u1__abc_45852_n662), .Y(u1__abc_45852_n663) );
  OR2X2 OR2X2_2445 ( .A(u1__abc_45852_n663), .B(u1__abc_45852_n661), .Y(u1__abc_45852_n664) );
  OR2X2 OR2X2_2446 ( .A(u1__abc_45852_n664), .B(u1__abc_45852_n660), .Y(u1__abc_45852_n665) );
  OR2X2 OR2X2_2447 ( .A(next_adr_bF_buf3), .B(u1_acs_addr_10_), .Y(u1__abc_45852_n667) );
  OR2X2 OR2X2_2448 ( .A(u1__abc_45852_n556_bF_buf1), .B(u1_acs_addr_pl1_10_), .Y(u1__abc_45852_n668) );
  OR2X2 OR2X2_2449 ( .A(u1__abc_45852_n669), .B(u1__abc_45852_n554_1_bF_buf3), .Y(u1__abc_45852_n670) );
  OR2X2 OR2X2_245 ( .A(u0__abc_49347_n1465), .B(spec_req_cs_0_bF_buf3), .Y(u0__abc_49347_n1466) );
  OR2X2 OR2X2_2450 ( .A(u1__abc_45852_n562_bF_buf1), .B(u1__abc_45852_n673), .Y(u1__abc_45852_n674) );
  OR2X2 OR2X2_2451 ( .A(u1__abc_45852_n674), .B(u1__abc_45852_n672), .Y(u1__abc_45852_n675) );
  OR2X2 OR2X2_2452 ( .A(u1__abc_45852_n675), .B(u1__abc_45852_n671), .Y(u1__abc_45852_n676) );
  OR2X2 OR2X2_2453 ( .A(next_adr_bF_buf2), .B(u1_acs_addr_11_), .Y(u1__abc_45852_n678) );
  OR2X2 OR2X2_2454 ( .A(u1__abc_45852_n556_bF_buf0), .B(u1_acs_addr_pl1_11_), .Y(u1__abc_45852_n679) );
  OR2X2 OR2X2_2455 ( .A(u1__abc_45852_n680), .B(u1__abc_45852_n554_1_bF_buf2), .Y(u1__abc_45852_n681) );
  OR2X2 OR2X2_2456 ( .A(u1__abc_45852_n562_bF_buf0), .B(u1__abc_45852_n684), .Y(u1__abc_45852_n685) );
  OR2X2 OR2X2_2457 ( .A(u1__abc_45852_n685), .B(u1__abc_45852_n683), .Y(u1__abc_45852_n686) );
  OR2X2 OR2X2_2458 ( .A(u1__abc_45852_n686), .B(u1__abc_45852_n682), .Y(u1__abc_45852_n687) );
  OR2X2 OR2X2_2459 ( .A(next_adr_bF_buf1), .B(u1_acs_addr_12_), .Y(u1__abc_45852_n689) );
  OR2X2 OR2X2_246 ( .A(u0__abc_49347_n1464), .B(u0__abc_49347_n1466), .Y(u0__abc_49347_n1467) );
  OR2X2 OR2X2_2460 ( .A(u1__abc_45852_n556_bF_buf3), .B(u1_acs_addr_pl1_12_), .Y(u1__abc_45852_n690) );
  OR2X2 OR2X2_2461 ( .A(u1__abc_45852_n691), .B(u1__abc_45852_n554_1_bF_buf1), .Y(u1__abc_45852_n692) );
  OR2X2 OR2X2_2462 ( .A(u1__abc_45852_n562_bF_buf3), .B(u1__abc_45852_n695), .Y(u1__abc_45852_n696) );
  OR2X2 OR2X2_2463 ( .A(u1__abc_45852_n696), .B(u1__abc_45852_n694), .Y(u1__abc_45852_n697) );
  OR2X2 OR2X2_2464 ( .A(u1__abc_45852_n697), .B(u1__abc_45852_n693), .Y(u1__abc_45852_n698) );
  OR2X2 OR2X2_2465 ( .A(next_adr_bF_buf0), .B(u1_acs_addr_13_), .Y(u1__abc_45852_n700) );
  OR2X2 OR2X2_2466 ( .A(u1__abc_45852_n556_bF_buf2), .B(u1_acs_addr_pl1_13_), .Y(u1__abc_45852_n701) );
  OR2X2 OR2X2_2467 ( .A(u1__abc_45852_n702), .B(u1__abc_45852_n554_1_bF_buf0), .Y(u1__abc_45852_n703) );
  OR2X2 OR2X2_2468 ( .A(u1__abc_45852_n562_bF_buf2), .B(u1__abc_45852_n706), .Y(u1__abc_45852_n707) );
  OR2X2 OR2X2_2469 ( .A(u1__abc_45852_n707), .B(u1__abc_45852_n705), .Y(u1__abc_45852_n708) );
  OR2X2 OR2X2_247 ( .A(u0__abc_49347_n1203_bF_buf0), .B(u0_tms0_11_), .Y(u0__abc_49347_n1468) );
  OR2X2 OR2X2_2470 ( .A(u1__abc_45852_n708), .B(u1__abc_45852_n704), .Y(u1__abc_45852_n709) );
  OR2X2 OR2X2_2471 ( .A(next_adr_bF_buf4), .B(u1_acs_addr_14_), .Y(u1__abc_45852_n711) );
  OR2X2 OR2X2_2472 ( .A(u1__abc_45852_n556_bF_buf1), .B(u1_acs_addr_pl1_14_), .Y(u1__abc_45852_n712) );
  OR2X2 OR2X2_2473 ( .A(u1__abc_45852_n713), .B(u1__abc_45852_n554_1_bF_buf4), .Y(u1__abc_45852_n714) );
  OR2X2 OR2X2_2474 ( .A(u1__abc_45852_n562_bF_buf1), .B(u1__abc_45852_n717), .Y(u1__abc_45852_n718) );
  OR2X2 OR2X2_2475 ( .A(u1__abc_45852_n718), .B(u1__abc_45852_n716), .Y(u1__abc_45852_n719) );
  OR2X2 OR2X2_2476 ( .A(u1__abc_45852_n719), .B(u1__abc_45852_n715), .Y(u1__abc_45852_n720) );
  OR2X2 OR2X2_2477 ( .A(next_adr_bF_buf3), .B(u1_acs_addr_15_), .Y(u1__abc_45852_n722) );
  OR2X2 OR2X2_2478 ( .A(u1__abc_45852_n556_bF_buf0), .B(u1_acs_addr_pl1_15_), .Y(u1__abc_45852_n723) );
  OR2X2 OR2X2_2479 ( .A(u1__abc_45852_n724), .B(u1__abc_45852_n554_1_bF_buf3), .Y(u1__abc_45852_n725) );
  OR2X2 OR2X2_248 ( .A(u0__abc_49347_n1470_1), .B(u0__abc_49347_n1448), .Y(u0_sp_tms_11__FF_INPUT) );
  OR2X2 OR2X2_2480 ( .A(u1__abc_45852_n562_bF_buf0), .B(u1__abc_45852_n728), .Y(u1__abc_45852_n729) );
  OR2X2 OR2X2_2481 ( .A(u1__abc_45852_n729), .B(u1__abc_45852_n727), .Y(u1__abc_45852_n730) );
  OR2X2 OR2X2_2482 ( .A(u1__abc_45852_n730), .B(u1__abc_45852_n726), .Y(u1__abc_45852_n731) );
  OR2X2 OR2X2_2483 ( .A(next_adr_bF_buf2), .B(u1_acs_addr_16_), .Y(u1__abc_45852_n733) );
  OR2X2 OR2X2_2484 ( .A(u1__abc_45852_n556_bF_buf3), .B(u1_acs_addr_pl1_16_), .Y(u1__abc_45852_n734) );
  OR2X2 OR2X2_2485 ( .A(u1__abc_45852_n735), .B(u1__abc_45852_n554_1_bF_buf2), .Y(u1__abc_45852_n736) );
  OR2X2 OR2X2_2486 ( .A(u1__abc_45852_n562_bF_buf3), .B(u1__abc_45852_n739), .Y(u1__abc_45852_n740) );
  OR2X2 OR2X2_2487 ( .A(u1__abc_45852_n740), .B(u1__abc_45852_n738), .Y(u1__abc_45852_n741) );
  OR2X2 OR2X2_2488 ( .A(u1__abc_45852_n741), .B(u1__abc_45852_n737), .Y(u1__abc_45852_n742) );
  OR2X2 OR2X2_2489 ( .A(next_adr_bF_buf1), .B(u1_acs_addr_17_), .Y(u1__abc_45852_n744) );
  OR2X2 OR2X2_249 ( .A(u0__abc_49347_n1183_1_bF_buf5), .B(1'b0), .Y(u0__abc_49347_n1474) );
  OR2X2 OR2X2_2490 ( .A(u1__abc_45852_n556_bF_buf2), .B(u1_acs_addr_pl1_17_), .Y(u1__abc_45852_n745) );
  OR2X2 OR2X2_2491 ( .A(u1__abc_45852_n746), .B(u1__abc_45852_n554_1_bF_buf1), .Y(u1__abc_45852_n747) );
  OR2X2 OR2X2_2492 ( .A(u1__abc_45852_n562_bF_buf2), .B(u1__abc_45852_n750), .Y(u1__abc_45852_n751) );
  OR2X2 OR2X2_2493 ( .A(u1__abc_45852_n751), .B(u1__abc_45852_n749), .Y(u1__abc_45852_n752) );
  OR2X2 OR2X2_2494 ( .A(u1__abc_45852_n752), .B(u1__abc_45852_n748), .Y(u1__abc_45852_n753) );
  OR2X2 OR2X2_2495 ( .A(next_adr_bF_buf0), .B(u1_acs_addr_18_), .Y(u1__abc_45852_n755) );
  OR2X2 OR2X2_2496 ( .A(u1__abc_45852_n556_bF_buf1), .B(u1_acs_addr_pl1_18_), .Y(u1__abc_45852_n756) );
  OR2X2 OR2X2_2497 ( .A(u1__abc_45852_n757), .B(u1__abc_45852_n554_1_bF_buf0), .Y(u1__abc_45852_n758) );
  OR2X2 OR2X2_2498 ( .A(u1__abc_45852_n562_bF_buf1), .B(u1__abc_45852_n761), .Y(u1__abc_45852_n762) );
  OR2X2 OR2X2_2499 ( .A(u1__abc_45852_n762), .B(u1__abc_45852_n760), .Y(u1__abc_45852_n763) );
  OR2X2 OR2X2_25 ( .A(_abc_55805_n274), .B(_abc_55805_n237_1), .Y(_abc_55805_n275) );
  OR2X2 OR2X2_250 ( .A(spec_req_cs_6_bF_buf2), .B(1'b0), .Y(u0__abc_49347_n1475) );
  OR2X2 OR2X2_2500 ( .A(u1__abc_45852_n763), .B(u1__abc_45852_n759), .Y(u1__abc_45852_n764) );
  OR2X2 OR2X2_2501 ( .A(next_adr_bF_buf4), .B(u1_acs_addr_19_), .Y(u1__abc_45852_n766) );
  OR2X2 OR2X2_2502 ( .A(u1__abc_45852_n556_bF_buf0), .B(u1_acs_addr_pl1_19_), .Y(u1__abc_45852_n767) );
  OR2X2 OR2X2_2503 ( .A(u1__abc_45852_n768), .B(u1__abc_45852_n554_1_bF_buf4), .Y(u1__abc_45852_n769) );
  OR2X2 OR2X2_2504 ( .A(u1__abc_45852_n562_bF_buf0), .B(u1__abc_45852_n772), .Y(u1__abc_45852_n773) );
  OR2X2 OR2X2_2505 ( .A(u1__abc_45852_n773), .B(u1__abc_45852_n771), .Y(u1__abc_45852_n774) );
  OR2X2 OR2X2_2506 ( .A(u1__abc_45852_n774), .B(u1__abc_45852_n770), .Y(u1__abc_45852_n775) );
  OR2X2 OR2X2_2507 ( .A(next_adr_bF_buf3), .B(u1_acs_addr_20_), .Y(u1__abc_45852_n777) );
  OR2X2 OR2X2_2508 ( .A(u1__abc_45852_n556_bF_buf3), .B(u1_acs_addr_pl1_20_), .Y(u1__abc_45852_n778) );
  OR2X2 OR2X2_2509 ( .A(u1__abc_45852_n779), .B(u1__abc_45852_n554_1_bF_buf3), .Y(u1__abc_45852_n780) );
  OR2X2 OR2X2_251 ( .A(u0__abc_49347_n1477), .B(u0__abc_49347_n1473), .Y(u0__abc_49347_n1478) );
  OR2X2 OR2X2_2510 ( .A(u1__abc_45852_n562_bF_buf3), .B(u1__abc_45852_n783), .Y(u1__abc_45852_n784) );
  OR2X2 OR2X2_2511 ( .A(u1__abc_45852_n784), .B(u1__abc_45852_n782), .Y(u1__abc_45852_n785) );
  OR2X2 OR2X2_2512 ( .A(u1__abc_45852_n785), .B(u1__abc_45852_n781), .Y(u1__abc_45852_n786) );
  OR2X2 OR2X2_2513 ( .A(next_adr_bF_buf2), .B(u1_acs_addr_21_), .Y(u1__abc_45852_n788) );
  OR2X2 OR2X2_2514 ( .A(u1__abc_45852_n556_bF_buf2), .B(u1_acs_addr_pl1_21_), .Y(u1__abc_45852_n789) );
  OR2X2 OR2X2_2515 ( .A(u1__abc_45852_n790), .B(u1__abc_45852_n554_1_bF_buf2), .Y(u1__abc_45852_n791) );
  OR2X2 OR2X2_2516 ( .A(u1__abc_45852_n562_bF_buf2), .B(u1__abc_45852_n794), .Y(u1__abc_45852_n795) );
  OR2X2 OR2X2_2517 ( .A(u1__abc_45852_n795), .B(u1__abc_45852_n793), .Y(u1__abc_45852_n796) );
  OR2X2 OR2X2_2518 ( .A(u1__abc_45852_n796), .B(u1__abc_45852_n792), .Y(u1__abc_45852_n797) );
  OR2X2 OR2X2_2519 ( .A(next_adr_bF_buf1), .B(u1_acs_addr_22_), .Y(u1__abc_45852_n799) );
  OR2X2 OR2X2_252 ( .A(u0__abc_49347_n1479_1), .B(u0__abc_49347_n1480_1), .Y(u0__abc_49347_n1481) );
  OR2X2 OR2X2_2520 ( .A(u1__abc_45852_n556_bF_buf1), .B(u1_acs_addr_pl1_22_), .Y(u1__abc_45852_n800) );
  OR2X2 OR2X2_2521 ( .A(u1__abc_45852_n801), .B(u1__abc_45852_n554_1_bF_buf1), .Y(u1__abc_45852_n802) );
  OR2X2 OR2X2_2522 ( .A(u1__abc_45852_n562_bF_buf1), .B(u1__abc_45852_n804), .Y(u1__abc_45852_n805) );
  OR2X2 OR2X2_2523 ( .A(u1__abc_45852_n805), .B(u1__abc_45852_n477_1), .Y(u1__abc_45852_n806) );
  OR2X2 OR2X2_2524 ( .A(u1__abc_45852_n806), .B(u1__abc_45852_n803), .Y(u1__abc_45852_n807) );
  OR2X2 OR2X2_2525 ( .A(next_adr_bF_buf0), .B(u1_acs_addr_23_), .Y(u1__abc_45852_n809) );
  OR2X2 OR2X2_2526 ( .A(u1__abc_45852_n556_bF_buf0), .B(u1_acs_addr_pl1_23_), .Y(u1__abc_45852_n810) );
  OR2X2 OR2X2_2527 ( .A(u1__abc_45852_n811), .B(u1__abc_45852_n554_1_bF_buf0), .Y(u1__abc_45852_n812) );
  OR2X2 OR2X2_2528 ( .A(u1__abc_45852_n562_bF_buf0), .B(u1__abc_45852_n815), .Y(u1__abc_45852_n816) );
  OR2X2 OR2X2_2529 ( .A(u1__abc_45852_n816), .B(u1__abc_45852_n814), .Y(u1__abc_45852_n817) );
  OR2X2 OR2X2_253 ( .A(u0__abc_49347_n1482), .B(u0__abc_49347_n1483), .Y(u0__abc_49347_n1484) );
  OR2X2 OR2X2_2530 ( .A(u1__abc_45852_n817), .B(u1__abc_45852_n813), .Y(u1__abc_45852_n818) );
  OR2X2 OR2X2_2531 ( .A(wb_stb_i_bF_buf2), .B(u1_sram_addr_0_), .Y(u1__abc_45852_n820) );
  OR2X2 OR2X2_2532 ( .A(u1__abc_45852_n821_bF_buf3), .B(\wb_addr_i[2] ), .Y(u1__abc_45852_n822) );
  OR2X2 OR2X2_2533 ( .A(wb_stb_i_bF_buf0), .B(u1_sram_addr_1_), .Y(u1__abc_45852_n824) );
  OR2X2 OR2X2_2534 ( .A(u1__abc_45852_n821_bF_buf2), .B(\wb_addr_i[3] ), .Y(u1__abc_45852_n825) );
  OR2X2 OR2X2_2535 ( .A(wb_stb_i_bF_buf5), .B(u1_sram_addr_2_), .Y(u1__abc_45852_n827) );
  OR2X2 OR2X2_2536 ( .A(u1__abc_45852_n821_bF_buf1), .B(\wb_addr_i[4] ), .Y(u1__abc_45852_n828) );
  OR2X2 OR2X2_2537 ( .A(wb_stb_i_bF_buf4), .B(u1_sram_addr_3_), .Y(u1__abc_45852_n830) );
  OR2X2 OR2X2_2538 ( .A(u1__abc_45852_n821_bF_buf0), .B(\wb_addr_i[5] ), .Y(u1__abc_45852_n831) );
  OR2X2 OR2X2_2539 ( .A(wb_stb_i_bF_buf3), .B(u1_sram_addr_4_), .Y(u1__abc_45852_n833) );
  OR2X2 OR2X2_254 ( .A(u0__abc_49347_n1485), .B(u0__abc_49347_n1486), .Y(u0__abc_49347_n1487) );
  OR2X2 OR2X2_2540 ( .A(u1__abc_45852_n821_bF_buf3), .B(\wb_addr_i[6] ), .Y(u1__abc_45852_n834) );
  OR2X2 OR2X2_2541 ( .A(wb_stb_i_bF_buf2), .B(u1_sram_addr_5_), .Y(u1__abc_45852_n836) );
  OR2X2 OR2X2_2542 ( .A(u1__abc_45852_n821_bF_buf2), .B(\wb_addr_i[7] ), .Y(u1__abc_45852_n837) );
  OR2X2 OR2X2_2543 ( .A(wb_stb_i_bF_buf1), .B(u1_sram_addr_6_), .Y(u1__abc_45852_n839) );
  OR2X2 OR2X2_2544 ( .A(u1__abc_45852_n821_bF_buf1), .B(\wb_addr_i[8] ), .Y(u1__abc_45852_n840) );
  OR2X2 OR2X2_2545 ( .A(wb_stb_i_bF_buf0), .B(u1_sram_addr_7_), .Y(u1__abc_45852_n842) );
  OR2X2 OR2X2_2546 ( .A(u1__abc_45852_n821_bF_buf0), .B(\wb_addr_i[9] ), .Y(u1__abc_45852_n843) );
  OR2X2 OR2X2_2547 ( .A(wb_stb_i_bF_buf5), .B(u1_sram_addr_8_), .Y(u1__abc_45852_n845) );
  OR2X2 OR2X2_2548 ( .A(u1__abc_45852_n821_bF_buf3), .B(\wb_addr_i[10] ), .Y(u1__abc_45852_n846) );
  OR2X2 OR2X2_2549 ( .A(wb_stb_i_bF_buf4), .B(u1_sram_addr_9_), .Y(u1__abc_45852_n848) );
  OR2X2 OR2X2_255 ( .A(u0__abc_49347_n1489_1), .B(spec_req_cs_0_bF_buf2), .Y(u0__abc_49347_n1490) );
  OR2X2 OR2X2_2550 ( .A(u1__abc_45852_n821_bF_buf2), .B(\wb_addr_i[11] ), .Y(u1__abc_45852_n849) );
  OR2X2 OR2X2_2551 ( .A(wb_stb_i_bF_buf3), .B(u1_sram_addr_10_), .Y(u1__abc_45852_n851) );
  OR2X2 OR2X2_2552 ( .A(u1__abc_45852_n821_bF_buf1), .B(\wb_addr_i[12] ), .Y(u1__abc_45852_n852) );
  OR2X2 OR2X2_2553 ( .A(wb_stb_i_bF_buf2), .B(u1_sram_addr_11_), .Y(u1__abc_45852_n854) );
  OR2X2 OR2X2_2554 ( .A(u1__abc_45852_n821_bF_buf0), .B(\wb_addr_i[13] ), .Y(u1__abc_45852_n855) );
  OR2X2 OR2X2_2555 ( .A(wb_stb_i_bF_buf1), .B(u1_sram_addr_12_), .Y(u1__abc_45852_n857) );
  OR2X2 OR2X2_2556 ( .A(u1__abc_45852_n821_bF_buf3), .B(\wb_addr_i[14] ), .Y(u1__abc_45852_n858) );
  OR2X2 OR2X2_2557 ( .A(wb_stb_i_bF_buf0), .B(u1_sram_addr_13_), .Y(u1__abc_45852_n860) );
  OR2X2 OR2X2_2558 ( .A(u1__abc_45852_n821_bF_buf2), .B(\wb_addr_i[15] ), .Y(u1__abc_45852_n861) );
  OR2X2 OR2X2_2559 ( .A(wb_stb_i_bF_buf5), .B(u1_sram_addr_14_), .Y(u1__abc_45852_n863) );
  OR2X2 OR2X2_256 ( .A(u0__abc_49347_n1488_1), .B(u0__abc_49347_n1490), .Y(u0__abc_49347_n1491) );
  OR2X2 OR2X2_2560 ( .A(u1__abc_45852_n821_bF_buf1), .B(\wb_addr_i[16] ), .Y(u1__abc_45852_n864) );
  OR2X2 OR2X2_2561 ( .A(wb_stb_i_bF_buf4), .B(u1_sram_addr_15_), .Y(u1__abc_45852_n866) );
  OR2X2 OR2X2_2562 ( .A(u1__abc_45852_n821_bF_buf0), .B(\wb_addr_i[17] ), .Y(u1__abc_45852_n867) );
  OR2X2 OR2X2_2563 ( .A(wb_stb_i_bF_buf3), .B(u1_sram_addr_16_), .Y(u1__abc_45852_n869) );
  OR2X2 OR2X2_2564 ( .A(u1__abc_45852_n821_bF_buf3), .B(\wb_addr_i[18] ), .Y(u1__abc_45852_n870) );
  OR2X2 OR2X2_2565 ( .A(wb_stb_i_bF_buf2), .B(u1_sram_addr_17_), .Y(u1__abc_45852_n872) );
  OR2X2 OR2X2_2566 ( .A(u1__abc_45852_n821_bF_buf2), .B(\wb_addr_i[19] ), .Y(u1__abc_45852_n873) );
  OR2X2 OR2X2_2567 ( .A(wb_stb_i_bF_buf1), .B(u1_sram_addr_18_), .Y(u1__abc_45852_n875) );
  OR2X2 OR2X2_2568 ( .A(u1__abc_45852_n821_bF_buf1), .B(\wb_addr_i[20] ), .Y(u1__abc_45852_n876) );
  OR2X2 OR2X2_2569 ( .A(wb_stb_i_bF_buf0), .B(u1_sram_addr_19_), .Y(u1__abc_45852_n878) );
  OR2X2 OR2X2_257 ( .A(u0__abc_49347_n1203_bF_buf5), .B(u0_tms0_12_), .Y(u0__abc_49347_n1492) );
  OR2X2 OR2X2_2570 ( .A(u1__abc_45852_n821_bF_buf0), .B(\wb_addr_i[21] ), .Y(u1__abc_45852_n879) );
  OR2X2 OR2X2_2571 ( .A(wb_stb_i_bF_buf5), .B(u1_sram_addr_20_), .Y(u1__abc_45852_n881) );
  OR2X2 OR2X2_2572 ( .A(u1__abc_45852_n821_bF_buf3), .B(\wb_addr_i[22] ), .Y(u1__abc_45852_n882) );
  OR2X2 OR2X2_2573 ( .A(wb_stb_i_bF_buf4), .B(u1_sram_addr_21_), .Y(u1__abc_45852_n884) );
  OR2X2 OR2X2_2574 ( .A(u1__abc_45852_n821_bF_buf2), .B(wb_addr_i_23_bF_buf3), .Y(u1__abc_45852_n885) );
  OR2X2 OR2X2_2575 ( .A(wb_stb_i_bF_buf3), .B(u1_sram_addr_22_), .Y(u1__abc_45852_n887) );
  OR2X2 OR2X2_2576 ( .A(u1__abc_45852_n821_bF_buf1), .B(\wb_addr_i[24] ), .Y(u1__abc_45852_n888) );
  OR2X2 OR2X2_2577 ( .A(wb_stb_i_bF_buf2), .B(u1_sram_addr_23_), .Y(u1__abc_45852_n890) );
  OR2X2 OR2X2_2578 ( .A(u1__abc_45852_n821_bF_buf0), .B(wb_addr_i_25_bF_buf2), .Y(u1__abc_45852_n891) );
  OR2X2 OR2X2_2579 ( .A(csc_s_3_), .B(csc_s_1_), .Y(u1__abc_45852_n893) );
  OR2X2 OR2X2_258 ( .A(u0__abc_49347_n1494), .B(u0__abc_49347_n1472), .Y(u0_sp_tms_12__FF_INPUT) );
  OR2X2 OR2X2_2580 ( .A(u1__abc_45852_n893_bF_buf4), .B(u1__abc_45852_n894), .Y(u1__abc_45852_n895) );
  OR2X2 OR2X2_2581 ( .A(csc_s_2_bF_buf2), .B(csc_s_3_), .Y(u1__abc_45852_n898) );
  OR2X2 OR2X2_2582 ( .A(u1__abc_45852_n904), .B(u1__abc_45852_n902), .Y(u1__abc_45852_n905) );
  OR2X2 OR2X2_2583 ( .A(u1__abc_45852_n905), .B(u1__abc_45852_n897_bF_buf3), .Y(u1__abc_45852_n906) );
  OR2X2 OR2X2_2584 ( .A(u1__abc_45852_n910), .B(row_adr_0_bF_buf5), .Y(u1__abc_45852_n911) );
  OR2X2 OR2X2_2585 ( .A(u1_col_adr_0_), .B(row_sel), .Y(u1__abc_45852_n912) );
  OR2X2 OR2X2_2586 ( .A(u1__abc_45852_n913), .B(u1__abc_45852_n909), .Y(u1__abc_45852_n914) );
  OR2X2 OR2X2_2587 ( .A(u1__abc_45852_n917), .B(tms_s_0_), .Y(u1__abc_45852_n918) );
  OR2X2 OR2X2_2588 ( .A(u1__abc_45852_n907), .B(u1__abc_45852_n920), .Y(mc_addr_d_0_) );
  OR2X2 OR2X2_2589 ( .A(u1__abc_45852_n893_bF_buf2), .B(u1__abc_45852_n922), .Y(u1__abc_45852_n923) );
  OR2X2 OR2X2_259 ( .A(u0__abc_49347_n1183_1_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n1498_1) );
  OR2X2 OR2X2_2590 ( .A(u1__abc_45852_n925), .B(u1__abc_45852_n924), .Y(u1__abc_45852_n926) );
  OR2X2 OR2X2_2591 ( .A(u1__abc_45852_n926), .B(u1__abc_45852_n897_bF_buf2), .Y(u1__abc_45852_n927) );
  OR2X2 OR2X2_2592 ( .A(u1__abc_45852_n910), .B(row_adr_1_bF_buf5), .Y(u1__abc_45852_n929) );
  OR2X2 OR2X2_2593 ( .A(u1_col_adr_1_), .B(row_sel), .Y(u1__abc_45852_n930) );
  OR2X2 OR2X2_2594 ( .A(u1__abc_45852_n931), .B(u1__abc_45852_n909), .Y(u1__abc_45852_n932) );
  OR2X2 OR2X2_2595 ( .A(u1__abc_45852_n917), .B(tms_s_1_), .Y(u1__abc_45852_n933) );
  OR2X2 OR2X2_2596 ( .A(u1__abc_45852_n928), .B(u1__abc_45852_n935), .Y(mc_addr_d_1_) );
  OR2X2 OR2X2_2597 ( .A(u1__abc_45852_n893_bF_buf1), .B(u1__abc_45852_n937), .Y(u1__abc_45852_n938) );
  OR2X2 OR2X2_2598 ( .A(u1__abc_45852_n940), .B(u1__abc_45852_n939), .Y(u1__abc_45852_n941) );
  OR2X2 OR2X2_2599 ( .A(u1__abc_45852_n941), .B(u1__abc_45852_n897_bF_buf1), .Y(u1__abc_45852_n942) );
  OR2X2 OR2X2_26 ( .A(_abc_55805_n245_1), .B(cs_need_rfr_5_), .Y(_abc_55805_n276) );
  OR2X2 OR2X2_260 ( .A(spec_req_cs_6_bF_buf1), .B(1'b0), .Y(u0__abc_49347_n1499) );
  OR2X2 OR2X2_2600 ( .A(u1__abc_45852_n910), .B(row_adr_2_bF_buf5), .Y(u1__abc_45852_n944) );
  OR2X2 OR2X2_2601 ( .A(u1_col_adr_2_), .B(row_sel), .Y(u1__abc_45852_n945) );
  OR2X2 OR2X2_2602 ( .A(u1__abc_45852_n946), .B(u1__abc_45852_n909), .Y(u1__abc_45852_n947) );
  OR2X2 OR2X2_2603 ( .A(u1__abc_45852_n917), .B(tms_s_2_), .Y(u1__abc_45852_n948) );
  OR2X2 OR2X2_2604 ( .A(u1__abc_45852_n943), .B(u1__abc_45852_n950), .Y(mc_addr_d_2_) );
  OR2X2 OR2X2_2605 ( .A(u1__abc_45852_n893_bF_buf0), .B(u1__abc_45852_n952), .Y(u1__abc_45852_n953) );
  OR2X2 OR2X2_2606 ( .A(u1__abc_45852_n955), .B(u1__abc_45852_n954), .Y(u1__abc_45852_n956) );
  OR2X2 OR2X2_2607 ( .A(u1__abc_45852_n956), .B(u1__abc_45852_n897_bF_buf0), .Y(u1__abc_45852_n957) );
  OR2X2 OR2X2_2608 ( .A(u1__abc_45852_n910), .B(row_adr_3_bF_buf5), .Y(u1__abc_45852_n959) );
  OR2X2 OR2X2_2609 ( .A(u1_col_adr_3_), .B(row_sel), .Y(u1__abc_45852_n960) );
  OR2X2 OR2X2_261 ( .A(u0__abc_49347_n1501), .B(u0__abc_49347_n1497_1), .Y(u0__abc_49347_n1502) );
  OR2X2 OR2X2_2610 ( .A(u1__abc_45852_n961), .B(u1__abc_45852_n909), .Y(u1__abc_45852_n962) );
  OR2X2 OR2X2_2611 ( .A(u1__abc_45852_n917), .B(tms_s_3_), .Y(u1__abc_45852_n963) );
  OR2X2 OR2X2_2612 ( .A(u1__abc_45852_n958), .B(u1__abc_45852_n965), .Y(mc_addr_d_3_) );
  OR2X2 OR2X2_2613 ( .A(u1__abc_45852_n893_bF_buf4), .B(u1__abc_45852_n967), .Y(u1__abc_45852_n968) );
  OR2X2 OR2X2_2614 ( .A(u1__abc_45852_n970), .B(u1__abc_45852_n969), .Y(u1__abc_45852_n971) );
  OR2X2 OR2X2_2615 ( .A(u1__abc_45852_n971), .B(u1__abc_45852_n897_bF_buf3), .Y(u1__abc_45852_n972) );
  OR2X2 OR2X2_2616 ( .A(u1__abc_45852_n910), .B(row_adr_4_bF_buf5), .Y(u1__abc_45852_n974) );
  OR2X2 OR2X2_2617 ( .A(u1_col_adr_4_), .B(row_sel), .Y(u1__abc_45852_n975) );
  OR2X2 OR2X2_2618 ( .A(u1__abc_45852_n976), .B(u1__abc_45852_n909), .Y(u1__abc_45852_n977) );
  OR2X2 OR2X2_2619 ( .A(u1__abc_45852_n917), .B(tms_s_4_), .Y(u1__abc_45852_n978) );
  OR2X2 OR2X2_262 ( .A(u0__abc_49347_n1503), .B(u0__abc_49347_n1504), .Y(u0__abc_49347_n1505) );
  OR2X2 OR2X2_2620 ( .A(u1__abc_45852_n973), .B(u1__abc_45852_n980), .Y(mc_addr_d_4_) );
  OR2X2 OR2X2_2621 ( .A(u1__abc_45852_n893_bF_buf3), .B(u1__abc_45852_n982), .Y(u1__abc_45852_n983) );
  OR2X2 OR2X2_2622 ( .A(u1__abc_45852_n985), .B(u1__abc_45852_n984), .Y(u1__abc_45852_n986) );
  OR2X2 OR2X2_2623 ( .A(u1__abc_45852_n986), .B(u1__abc_45852_n897_bF_buf2), .Y(u1__abc_45852_n987) );
  OR2X2 OR2X2_2624 ( .A(u1__abc_45852_n910), .B(row_adr_5_bF_buf5), .Y(u1__abc_45852_n989) );
  OR2X2 OR2X2_2625 ( .A(u1_col_adr_5_), .B(row_sel), .Y(u1__abc_45852_n990) );
  OR2X2 OR2X2_2626 ( .A(u1__abc_45852_n991), .B(u1__abc_45852_n909), .Y(u1__abc_45852_n992) );
  OR2X2 OR2X2_2627 ( .A(u1__abc_45852_n917), .B(tms_s_5_), .Y(u1__abc_45852_n993) );
  OR2X2 OR2X2_2628 ( .A(u1__abc_45852_n988), .B(u1__abc_45852_n995), .Y(mc_addr_d_5_) );
  OR2X2 OR2X2_2629 ( .A(u1__abc_45852_n893_bF_buf2), .B(u1__abc_45852_n997), .Y(u1__abc_45852_n998) );
  OR2X2 OR2X2_263 ( .A(u0__abc_49347_n1506_1), .B(u0__abc_49347_n1507_1), .Y(u0__abc_49347_n1508) );
  OR2X2 OR2X2_2630 ( .A(u1__abc_45852_n1000), .B(u1__abc_45852_n999), .Y(u1__abc_45852_n1001) );
  OR2X2 OR2X2_2631 ( .A(u1__abc_45852_n1001), .B(u1__abc_45852_n897_bF_buf1), .Y(u1__abc_45852_n1002) );
  OR2X2 OR2X2_2632 ( .A(u1__abc_45852_n910), .B(row_adr_6_bF_buf5), .Y(u1__abc_45852_n1004) );
  OR2X2 OR2X2_2633 ( .A(u1_col_adr_6_), .B(row_sel), .Y(u1__abc_45852_n1005) );
  OR2X2 OR2X2_2634 ( .A(u1__abc_45852_n1006), .B(u1__abc_45852_n909), .Y(u1__abc_45852_n1007) );
  OR2X2 OR2X2_2635 ( .A(u1__abc_45852_n917), .B(tms_s_6_), .Y(u1__abc_45852_n1008) );
  OR2X2 OR2X2_2636 ( .A(u1__abc_45852_n1003), .B(u1__abc_45852_n1010), .Y(mc_addr_d_6_) );
  OR2X2 OR2X2_2637 ( .A(u1__abc_45852_n893_bF_buf1), .B(u1__abc_45852_n1012), .Y(u1__abc_45852_n1013) );
  OR2X2 OR2X2_2638 ( .A(u1__abc_45852_n1015), .B(u1__abc_45852_n1014), .Y(u1__abc_45852_n1016) );
  OR2X2 OR2X2_2639 ( .A(u1__abc_45852_n1016), .B(u1__abc_45852_n897_bF_buf0), .Y(u1__abc_45852_n1017) );
  OR2X2 OR2X2_264 ( .A(u0__abc_49347_n1509), .B(u0__abc_49347_n1510), .Y(u0__abc_49347_n1511) );
  OR2X2 OR2X2_2640 ( .A(u1__abc_45852_n910), .B(row_adr_7_bF_buf5), .Y(u1__abc_45852_n1019) );
  OR2X2 OR2X2_2641 ( .A(u1_col_adr_7_), .B(row_sel), .Y(u1__abc_45852_n1020) );
  OR2X2 OR2X2_2642 ( .A(u1__abc_45852_n1021), .B(u1__abc_45852_n909), .Y(u1__abc_45852_n1022) );
  OR2X2 OR2X2_2643 ( .A(u1__abc_45852_n917), .B(tms_s_7_), .Y(u1__abc_45852_n1023) );
  OR2X2 OR2X2_2644 ( .A(u1__abc_45852_n1018), .B(u1__abc_45852_n1025), .Y(mc_addr_d_7_) );
  OR2X2 OR2X2_2645 ( .A(u1__abc_45852_n893_bF_buf0), .B(u1__abc_45852_n1027), .Y(u1__abc_45852_n1028) );
  OR2X2 OR2X2_2646 ( .A(u1__abc_45852_n1030), .B(u1__abc_45852_n1029), .Y(u1__abc_45852_n1031) );
  OR2X2 OR2X2_2647 ( .A(u1__abc_45852_n1031), .B(u1__abc_45852_n897_bF_buf3), .Y(u1__abc_45852_n1032) );
  OR2X2 OR2X2_2648 ( .A(u1__abc_45852_n910), .B(row_adr_8_bF_buf5), .Y(u1__abc_45852_n1034) );
  OR2X2 OR2X2_2649 ( .A(u1_col_adr_8_), .B(row_sel), .Y(u1__abc_45852_n1035) );
  OR2X2 OR2X2_265 ( .A(u0__abc_49347_n1513), .B(spec_req_cs_0_bF_buf1), .Y(u0__abc_49347_n1514) );
  OR2X2 OR2X2_2650 ( .A(u1__abc_45852_n1036), .B(u1__abc_45852_n909), .Y(u1__abc_45852_n1037) );
  OR2X2 OR2X2_2651 ( .A(u1__abc_45852_n917), .B(tms_s_8_), .Y(u1__abc_45852_n1038) );
  OR2X2 OR2X2_2652 ( .A(u1__abc_45852_n1033), .B(u1__abc_45852_n1040), .Y(mc_addr_d_8_) );
  OR2X2 OR2X2_2653 ( .A(u1__abc_45852_n893_bF_buf4), .B(u1__abc_45852_n1042), .Y(u1__abc_45852_n1043) );
  OR2X2 OR2X2_2654 ( .A(u1__abc_45852_n1045), .B(u1__abc_45852_n1044), .Y(u1__abc_45852_n1046) );
  OR2X2 OR2X2_2655 ( .A(u1__abc_45852_n1046), .B(u1__abc_45852_n897_bF_buf2), .Y(u1__abc_45852_n1047) );
  OR2X2 OR2X2_2656 ( .A(u1__abc_45852_n910), .B(row_adr_9_bF_buf5), .Y(u1__abc_45852_n1049) );
  OR2X2 OR2X2_2657 ( .A(u1_col_adr_9_), .B(row_sel), .Y(u1__abc_45852_n1050) );
  OR2X2 OR2X2_2658 ( .A(u1__abc_45852_n1051), .B(u1__abc_45852_n909), .Y(u1__abc_45852_n1052) );
  OR2X2 OR2X2_2659 ( .A(u1__abc_45852_n917), .B(tms_s_9_), .Y(u1__abc_45852_n1053) );
  OR2X2 OR2X2_266 ( .A(u0__abc_49347_n1512), .B(u0__abc_49347_n1514), .Y(u0__abc_49347_n1515_1) );
  OR2X2 OR2X2_2660 ( .A(u1__abc_45852_n1048), .B(u1__abc_45852_n1055), .Y(mc_addr_d_9_) );
  OR2X2 OR2X2_2661 ( .A(u1__abc_45852_n917), .B(tms_s_11_), .Y(u1__abc_45852_n1057) );
  OR2X2 OR2X2_2662 ( .A(u1__abc_45852_n909), .B(u1__abc_45852_n1058), .Y(u1__abc_45852_n1059) );
  OR2X2 OR2X2_2663 ( .A(u1__abc_45852_n893_bF_buf3), .B(u1__abc_45852_n1062), .Y(u1__abc_45852_n1063) );
  OR2X2 OR2X2_2664 ( .A(u1__abc_45852_n903_bF_buf1), .B(u1_sram_addr_11_), .Y(u1__abc_45852_n1064) );
  OR2X2 OR2X2_2665 ( .A(u1__abc_45852_n901_bF_buf3), .B(\wb_addr_i[13] ), .Y(u1__abc_45852_n1065) );
  OR2X2 OR2X2_2666 ( .A(u1__abc_45852_n1066), .B(u1__abc_45852_n897_bF_buf1), .Y(u1__abc_45852_n1067) );
  OR2X2 OR2X2_2667 ( .A(u1__abc_45852_n1068), .B(u1__abc_45852_n1061), .Y(mc_addr_d_11_) );
  OR2X2 OR2X2_2668 ( .A(u1__abc_45852_n917), .B(tms_s_12_), .Y(u1__abc_45852_n1070) );
  OR2X2 OR2X2_2669 ( .A(u1__abc_45852_n909), .B(u1__abc_45852_n1071), .Y(u1__abc_45852_n1072) );
  OR2X2 OR2X2_267 ( .A(u0__abc_49347_n1203_bF_buf4), .B(u0_tms0_13_), .Y(u0__abc_49347_n1516_1) );
  OR2X2 OR2X2_2670 ( .A(u1__abc_45852_n893_bF_buf2), .B(u1__abc_45852_n1075), .Y(u1__abc_45852_n1076) );
  OR2X2 OR2X2_2671 ( .A(u1__abc_45852_n903_bF_buf0), .B(u1_sram_addr_12_), .Y(u1__abc_45852_n1077) );
  OR2X2 OR2X2_2672 ( .A(u1__abc_45852_n901_bF_buf2), .B(\wb_addr_i[14] ), .Y(u1__abc_45852_n1078) );
  OR2X2 OR2X2_2673 ( .A(u1__abc_45852_n1079), .B(u1__abc_45852_n897_bF_buf0), .Y(u1__abc_45852_n1080) );
  OR2X2 OR2X2_2674 ( .A(u1__abc_45852_n1081), .B(u1__abc_45852_n1074), .Y(mc_addr_d_12_) );
  OR2X2 OR2X2_2675 ( .A(u1__abc_45852_n893_bF_buf1), .B(u1__abc_45852_n1084), .Y(u1__abc_45852_n1085) );
  OR2X2 OR2X2_2676 ( .A(u1__abc_45852_n903_bF_buf3), .B(u1_sram_addr_13_), .Y(u1__abc_45852_n1086) );
  OR2X2 OR2X2_2677 ( .A(u1__abc_45852_n901_bF_buf1), .B(\wb_addr_i[15] ), .Y(u1__abc_45852_n1087) );
  OR2X2 OR2X2_2678 ( .A(u1__abc_45852_n1088), .B(u1__abc_45852_n897_bF_buf3), .Y(u1__abc_45852_n1089) );
  OR2X2 OR2X2_2679 ( .A(u1__abc_45852_n1090), .B(u1__abc_45852_n1083), .Y(mc_addr_d_13_) );
  OR2X2 OR2X2_268 ( .A(u0__abc_49347_n1518), .B(u0__abc_49347_n1496), .Y(u0_sp_tms_13__FF_INPUT) );
  OR2X2 OR2X2_2680 ( .A(u1__abc_45852_n893_bF_buf0), .B(u1__abc_45852_n1093), .Y(u1__abc_45852_n1094) );
  OR2X2 OR2X2_2681 ( .A(u1__abc_45852_n903_bF_buf2), .B(u1_sram_addr_14_), .Y(u1__abc_45852_n1095) );
  OR2X2 OR2X2_2682 ( .A(u1__abc_45852_n901_bF_buf0), .B(\wb_addr_i[16] ), .Y(u1__abc_45852_n1096) );
  OR2X2 OR2X2_2683 ( .A(u1__abc_45852_n1097), .B(u1__abc_45852_n897_bF_buf2), .Y(u1__abc_45852_n1098) );
  OR2X2 OR2X2_2684 ( .A(u1__abc_45852_n1099), .B(u1__abc_45852_n1092), .Y(mc_addr_d_14_) );
  OR2X2 OR2X2_2685 ( .A(u1__abc_45852_n893_bF_buf4), .B(u1__abc_45852_n1101), .Y(u1__abc_45852_n1102) );
  OR2X2 OR2X2_2686 ( .A(u1__abc_45852_n1104), .B(u1__abc_45852_n897_bF_buf1), .Y(u1__abc_45852_n1105) );
  OR2X2 OR2X2_2687 ( .A(u1__abc_45852_n1105), .B(u1__abc_45852_n1103), .Y(u1__abc_45852_n1106) );
  OR2X2 OR2X2_2688 ( .A(u1__abc_45852_n893_bF_buf3), .B(u1__abc_45852_n1108), .Y(u1__abc_45852_n1109) );
  OR2X2 OR2X2_2689 ( .A(u1__abc_45852_n1111), .B(u1__abc_45852_n1110), .Y(u1__abc_45852_n1112) );
  OR2X2 OR2X2_269 ( .A(u0__abc_49347_n1183_1_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n1522) );
  OR2X2 OR2X2_2690 ( .A(u1__abc_45852_n1112), .B(u1__abc_45852_n897_bF_buf0), .Y(u1__abc_45852_n1113) );
  OR2X2 OR2X2_2691 ( .A(u1__abc_45852_n893_bF_buf2), .B(u1__abc_45852_n1115), .Y(u1__abc_45852_n1116) );
  OR2X2 OR2X2_2692 ( .A(u1__abc_45852_n1118), .B(u1__abc_45852_n1117), .Y(u1__abc_45852_n1119) );
  OR2X2 OR2X2_2693 ( .A(u1__abc_45852_n1119), .B(u1__abc_45852_n897_bF_buf3), .Y(u1__abc_45852_n1120) );
  OR2X2 OR2X2_2694 ( .A(u1__abc_45852_n893_bF_buf1), .B(u1__abc_45852_n1122), .Y(u1__abc_45852_n1123) );
  OR2X2 OR2X2_2695 ( .A(u1__abc_45852_n1125), .B(u1__abc_45852_n1124), .Y(u1__abc_45852_n1126) );
  OR2X2 OR2X2_2696 ( .A(u1__abc_45852_n1126), .B(u1__abc_45852_n897_bF_buf2), .Y(u1__abc_45852_n1127) );
  OR2X2 OR2X2_2697 ( .A(u1__abc_45852_n893_bF_buf0), .B(u1__abc_45852_n1129), .Y(u1__abc_45852_n1130) );
  OR2X2 OR2X2_2698 ( .A(u1__abc_45852_n1132), .B(u1__abc_45852_n1131), .Y(u1__abc_45852_n1133) );
  OR2X2 OR2X2_2699 ( .A(u1__abc_45852_n1133), .B(u1__abc_45852_n897_bF_buf1), .Y(u1__abc_45852_n1134) );
  OR2X2 OR2X2_27 ( .A(_abc_55805_n240_bF_buf5), .B(spec_req_cs_6_bF_buf5), .Y(_abc_55805_n278) );
  OR2X2 OR2X2_270 ( .A(spec_req_cs_6_bF_buf0), .B(1'b0), .Y(u0__abc_49347_n1523) );
  OR2X2 OR2X2_2700 ( .A(u1__abc_45852_n893_bF_buf4), .B(u1__abc_45852_n1136), .Y(u1__abc_45852_n1137) );
  OR2X2 OR2X2_2701 ( .A(u1__abc_45852_n1139), .B(u1__abc_45852_n1138), .Y(u1__abc_45852_n1140) );
  OR2X2 OR2X2_2702 ( .A(u1__abc_45852_n1140), .B(u1__abc_45852_n897_bF_buf0), .Y(u1__abc_45852_n1141) );
  OR2X2 OR2X2_2703 ( .A(u1__abc_45852_n893_bF_buf3), .B(u1__abc_45852_n1143), .Y(u1__abc_45852_n1144) );
  OR2X2 OR2X2_2704 ( .A(u1__abc_45852_n1146), .B(u1__abc_45852_n1145), .Y(u1__abc_45852_n1147) );
  OR2X2 OR2X2_2705 ( .A(u1__abc_45852_n1147), .B(u1__abc_45852_n897_bF_buf3), .Y(u1__abc_45852_n1148) );
  OR2X2 OR2X2_2706 ( .A(u1__abc_45852_n893_bF_buf2), .B(u1__abc_45852_n1150), .Y(u1__abc_45852_n1151) );
  OR2X2 OR2X2_2707 ( .A(u1__abc_45852_n1153), .B(u1__abc_45852_n1152), .Y(u1__abc_45852_n1154) );
  OR2X2 OR2X2_2708 ( .A(u1__abc_45852_n1154), .B(u1__abc_45852_n897_bF_buf2), .Y(u1__abc_45852_n1155) );
  OR2X2 OR2X2_2709 ( .A(u1__abc_45852_n893_bF_buf1), .B(u1__abc_45852_n1157), .Y(u1__abc_45852_n1158) );
  OR2X2 OR2X2_271 ( .A(u0__abc_49347_n1525_1), .B(u0__abc_49347_n1521), .Y(u0__abc_49347_n1526) );
  OR2X2 OR2X2_2710 ( .A(u1__abc_45852_n1160), .B(u1__abc_45852_n1159), .Y(u1__abc_45852_n1161) );
  OR2X2 OR2X2_2711 ( .A(u1__abc_45852_n1161), .B(u1__abc_45852_n897_bF_buf1), .Y(u1__abc_45852_n1162) );
  OR2X2 OR2X2_2712 ( .A(u1__abc_45852_n901_bF_buf0), .B(\wb_addr_i[12] ), .Y(u1__abc_45852_n1164) );
  OR2X2 OR2X2_2713 ( .A(u1__abc_45852_n903_bF_buf0), .B(u1_sram_addr_10_), .Y(u1__abc_45852_n1165) );
  OR2X2 OR2X2_2714 ( .A(u1__abc_45852_n1166), .B(u1__abc_45852_n897_bF_buf0), .Y(u1__abc_45852_n1167) );
  OR2X2 OR2X2_2715 ( .A(u1__abc_45852_n893_bF_buf0), .B(u1__abc_45852_n1168), .Y(u1__abc_45852_n1169) );
  OR2X2 OR2X2_2716 ( .A(row_sel), .B(cmd_a10), .Y(u1__abc_45852_n1171) );
  OR2X2 OR2X2_2717 ( .A(u1__abc_45852_n910), .B(row_adr_10_bF_buf5), .Y(u1__abc_45852_n1172) );
  OR2X2 OR2X2_2718 ( .A(u1__abc_45852_n1173), .B(u1__abc_45852_n909), .Y(u1__abc_45852_n1174) );
  OR2X2 OR2X2_2719 ( .A(u1__abc_45852_n917), .B(tms_s_10_), .Y(u1__abc_45852_n1175) );
  OR2X2 OR2X2_272 ( .A(u0__abc_49347_n1527), .B(u0__abc_49347_n1528), .Y(u0__abc_49347_n1529) );
  OR2X2 OR2X2_2720 ( .A(u1__abc_45852_n1177), .B(rfr_ack), .Y(u1__abc_45852_n1178) );
  OR2X2 OR2X2_2721 ( .A(u1__abc_45852_n1170), .B(u1__abc_45852_n1178), .Y(mc_addr_d_10_) );
  OR2X2 OR2X2_2722 ( .A(u1_u0__abc_45749_n51), .B(u1_acs_addr_13_), .Y(u1_u0__abc_45749_n54) );
  OR2X2 OR2X2_2723 ( .A(u1_u0__abc_45749_n52_1), .B(u1_acs_addr_14_), .Y(u1_u0__abc_45749_n58) );
  OR2X2 OR2X2_2724 ( .A(u1_u0__abc_45749_n56_1), .B(u1_acs_addr_15_), .Y(u1_u0__abc_45749_n60_1) );
  OR2X2 OR2X2_2725 ( .A(u1_u0__abc_45749_n62_1), .B(u1_acs_addr_16_), .Y(u1_u0__abc_45749_n67_1) );
  OR2X2 OR2X2_2726 ( .A(u1_u0__abc_45749_n65), .B(u1_acs_addr_17_), .Y(u1_u0__abc_45749_n69) );
  OR2X2 OR2X2_2727 ( .A(u1_u0__abc_45749_n71_1), .B(u1_acs_addr_18_), .Y(u1_u0__abc_45749_n76) );
  OR2X2 OR2X2_2728 ( .A(u1_u0__abc_45749_n74_1), .B(u1_acs_addr_19_), .Y(u1_u0__abc_45749_n78_1) );
  OR2X2 OR2X2_2729 ( .A(u1_u0__abc_45749_n81), .B(u1_acs_addr_20_), .Y(u1_u0__abc_45749_n86) );
  OR2X2 OR2X2_273 ( .A(u0__abc_49347_n1530), .B(u0__abc_49347_n1531), .Y(u0__abc_49347_n1532) );
  OR2X2 OR2X2_2730 ( .A(u1_u0__abc_45749_n84), .B(u1_acs_addr_21_), .Y(u1_u0__abc_45749_n88) );
  OR2X2 OR2X2_2731 ( .A(u1_u0__abc_45749_n90), .B(u1_acs_addr_22_), .Y(u1_u0__abc_45749_n95) );
  OR2X2 OR2X2_2732 ( .A(u1_u0__abc_45749_n93), .B(u1_acs_addr_23_), .Y(u1_u0__abc_45749_n97) );
  OR2X2 OR2X2_2733 ( .A(u1_u0_inc_next), .B(u1_acs_addr_12_), .Y(u1_u0__abc_45749_n102) );
  OR2X2 OR2X2_2734 ( .A(u1_acs_addr_0_), .B(u1_acs_addr_1_), .Y(u1_u0__abc_45749_n106) );
  OR2X2 OR2X2_2735 ( .A(u1_u0__abc_45749_n104), .B(u1_acs_addr_2_), .Y(u1_u0__abc_45749_n110) );
  OR2X2 OR2X2_2736 ( .A(u1_u0__abc_45749_n108), .B(u1_acs_addr_3_), .Y(u1_u0__abc_45749_n114) );
  OR2X2 OR2X2_2737 ( .A(u1_u0__abc_45749_n112), .B(u1_acs_addr_4_), .Y(u1_u0__abc_45749_n118) );
  OR2X2 OR2X2_2738 ( .A(u1_u0__abc_45749_n116), .B(u1_acs_addr_5_), .Y(u1_u0__abc_45749_n120) );
  OR2X2 OR2X2_2739 ( .A(u1_u0__abc_45749_n122), .B(u1_acs_addr_6_), .Y(u1_u0__abc_45749_n127) );
  OR2X2 OR2X2_274 ( .A(u0__abc_49347_n1533_1), .B(u0__abc_49347_n1534_1), .Y(u0__abc_49347_n1535) );
  OR2X2 OR2X2_2740 ( .A(u1_u0__abc_45749_n125), .B(u1_acs_addr_7_), .Y(u1_u0__abc_45749_n129) );
  OR2X2 OR2X2_2741 ( .A(u1_u0__abc_45749_n132), .B(u1_acs_addr_8_), .Y(u1_u0__abc_45749_n137) );
  OR2X2 OR2X2_2742 ( .A(u1_u0__abc_45749_n135), .B(u1_acs_addr_9_), .Y(u1_u0__abc_45749_n139) );
  OR2X2 OR2X2_2743 ( .A(u1_u0__abc_45749_n141), .B(u1_acs_addr_10_), .Y(u1_u0__abc_45749_n146) );
  OR2X2 OR2X2_2744 ( .A(u1_u0__abc_45749_n144), .B(u1_acs_addr_11_), .Y(u1_u0__abc_45749_n150) );
  OR2X2 OR2X2_2745 ( .A(u2__abc_48153_n80), .B(rfr_ack), .Y(u2_bank_clr_all_0) );
  OR2X2 OR2X2_2746 ( .A(u2__abc_48153_n82_1), .B(rfr_ack), .Y(u2_bank_clr_all_1) );
  OR2X2 OR2X2_2747 ( .A(u2__abc_48153_n84_1), .B(rfr_ack), .Y(u2_bank_clr_all_2) );
  OR2X2 OR2X2_2748 ( .A(u2__abc_48153_n86), .B(rfr_ack), .Y(u2_bank_clr_all_3) );
  OR2X2 OR2X2_2749 ( .A(u2__abc_48153_n88_1), .B(rfr_ack), .Y(u2_bank_clr_all_4) );
  OR2X2 OR2X2_275 ( .A(u0__abc_49347_n1537), .B(spec_req_cs_0_bF_buf0), .Y(u0__abc_49347_n1538) );
  OR2X2 OR2X2_2750 ( .A(u2__abc_48153_n90), .B(rfr_ack), .Y(u2_bank_clr_all_5) );
  OR2X2 OR2X2_2751 ( .A(u2__abc_48153_n96), .B(u2__abc_48153_n97), .Y(u2__abc_48153_n98) );
  OR2X2 OR2X2_2752 ( .A(u2__abc_48153_n99), .B(u2__abc_48153_n100), .Y(u2__abc_48153_n101) );
  OR2X2 OR2X2_2753 ( .A(u2__abc_48153_n98), .B(u2__abc_48153_n101), .Y(u2__abc_48153_n102) );
  OR2X2 OR2X2_2754 ( .A(u2__abc_48153_n103), .B(u2__abc_48153_n104), .Y(u2__abc_48153_n105) );
  OR2X2 OR2X2_2755 ( .A(u2__abc_48153_n106), .B(u2__abc_48153_n107), .Y(u2__abc_48153_n108) );
  OR2X2 OR2X2_2756 ( .A(u2__abc_48153_n105), .B(u2__abc_48153_n108), .Y(u2__abc_48153_n109) );
  OR2X2 OR2X2_2757 ( .A(u2__abc_48153_n102), .B(u2__abc_48153_n109), .Y(u2_bank_open_FF_INPUT) );
  OR2X2 OR2X2_2758 ( .A(u2__abc_48153_n111), .B(u2__abc_48153_n112), .Y(u2__abc_48153_n113) );
  OR2X2 OR2X2_2759 ( .A(u2__abc_48153_n114), .B(u2__abc_48153_n115), .Y(u2__abc_48153_n116) );
  OR2X2 OR2X2_276 ( .A(u0__abc_49347_n1536), .B(u0__abc_49347_n1538), .Y(u0__abc_49347_n1539) );
  OR2X2 OR2X2_2760 ( .A(u2__abc_48153_n113), .B(u2__abc_48153_n116), .Y(u2__abc_48153_n117) );
  OR2X2 OR2X2_2761 ( .A(u2__abc_48153_n118), .B(u2__abc_48153_n119), .Y(u2__abc_48153_n120) );
  OR2X2 OR2X2_2762 ( .A(u2__abc_48153_n121), .B(u2__abc_48153_n122), .Y(u2__abc_48153_n123) );
  OR2X2 OR2X2_2763 ( .A(u2__abc_48153_n120), .B(u2__abc_48153_n123), .Y(u2__abc_48153_n124) );
  OR2X2 OR2X2_2764 ( .A(u2__abc_48153_n117), .B(u2__abc_48153_n124), .Y(u2_row_same_FF_INPUT) );
  OR2X2 OR2X2_2765 ( .A(u2_u0__abc_47660_n137_bF_buf4), .B(u2_u0_b3_last_row_0_), .Y(u2_u0__abc_47660_n138) );
  OR2X2 OR2X2_2766 ( .A(u2_u0__abc_47660_n137_bF_buf2), .B(u2_u0_b3_last_row_1_), .Y(u2_u0__abc_47660_n143) );
  OR2X2 OR2X2_2767 ( .A(u2_u0__abc_47660_n137_bF_buf0), .B(u2_u0_b3_last_row_2_), .Y(u2_u0__abc_47660_n148) );
  OR2X2 OR2X2_2768 ( .A(u2_u0__abc_47660_n137_bF_buf3), .B(u2_u0_b3_last_row_3_), .Y(u2_u0__abc_47660_n153) );
  OR2X2 OR2X2_2769 ( .A(u2_u0__abc_47660_n137_bF_buf1), .B(u2_u0_b3_last_row_4_), .Y(u2_u0__abc_47660_n158) );
  OR2X2 OR2X2_277 ( .A(u0__abc_49347_n1203_bF_buf3), .B(u0_tms0_14_), .Y(u0__abc_49347_n1540) );
  OR2X2 OR2X2_2770 ( .A(u2_u0__abc_47660_n137_bF_buf4), .B(u2_u0_b3_last_row_5_), .Y(u2_u0__abc_47660_n163) );
  OR2X2 OR2X2_2771 ( .A(u2_u0__abc_47660_n137_bF_buf2), .B(u2_u0_b3_last_row_6_), .Y(u2_u0__abc_47660_n168) );
  OR2X2 OR2X2_2772 ( .A(u2_u0__abc_47660_n137_bF_buf0), .B(u2_u0_b3_last_row_7_), .Y(u2_u0__abc_47660_n173) );
  OR2X2 OR2X2_2773 ( .A(u2_u0__abc_47660_n137_bF_buf3), .B(u2_u0_b3_last_row_8_), .Y(u2_u0__abc_47660_n178) );
  OR2X2 OR2X2_2774 ( .A(u2_u0__abc_47660_n137_bF_buf1), .B(u2_u0_b3_last_row_9_), .Y(u2_u0__abc_47660_n183) );
  OR2X2 OR2X2_2775 ( .A(u2_u0__abc_47660_n137_bF_buf4), .B(u2_u0_b3_last_row_10_), .Y(u2_u0__abc_47660_n188) );
  OR2X2 OR2X2_2776 ( .A(u2_u0__abc_47660_n137_bF_buf2), .B(u2_u0_b3_last_row_11_), .Y(u2_u0__abc_47660_n193) );
  OR2X2 OR2X2_2777 ( .A(u2_u0__abc_47660_n137_bF_buf0), .B(u2_u0_b3_last_row_12_), .Y(u2_u0__abc_47660_n198) );
  OR2X2 OR2X2_2778 ( .A(u2_u0__abc_47660_n205), .B(u2_u0_b2_last_row_0_), .Y(u2_u0__abc_47660_n206) );
  OR2X2 OR2X2_2779 ( .A(u2_u0__abc_47660_n207), .B(row_adr_0_bF_buf3), .Y(u2_u0__abc_47660_n208) );
  OR2X2 OR2X2_278 ( .A(u0__abc_49347_n1542_1), .B(u0__abc_49347_n1520), .Y(u0_sp_tms_14__FF_INPUT) );
  OR2X2 OR2X2_2780 ( .A(u2_u0__abc_47660_n205), .B(u2_u0_b2_last_row_1_), .Y(u2_u0__abc_47660_n210) );
  OR2X2 OR2X2_2781 ( .A(u2_u0__abc_47660_n207), .B(row_adr_1_bF_buf3), .Y(u2_u0__abc_47660_n211) );
  OR2X2 OR2X2_2782 ( .A(u2_u0__abc_47660_n205), .B(u2_u0_b2_last_row_2_), .Y(u2_u0__abc_47660_n213) );
  OR2X2 OR2X2_2783 ( .A(u2_u0__abc_47660_n207), .B(row_adr_2_bF_buf3), .Y(u2_u0__abc_47660_n214) );
  OR2X2 OR2X2_2784 ( .A(u2_u0__abc_47660_n205), .B(u2_u0_b2_last_row_3_), .Y(u2_u0__abc_47660_n216) );
  OR2X2 OR2X2_2785 ( .A(u2_u0__abc_47660_n207), .B(row_adr_3_bF_buf3), .Y(u2_u0__abc_47660_n217) );
  OR2X2 OR2X2_2786 ( .A(u2_u0__abc_47660_n205), .B(u2_u0_b2_last_row_4_), .Y(u2_u0__abc_47660_n219) );
  OR2X2 OR2X2_2787 ( .A(u2_u0__abc_47660_n207), .B(row_adr_4_bF_buf3), .Y(u2_u0__abc_47660_n220) );
  OR2X2 OR2X2_2788 ( .A(u2_u0__abc_47660_n205), .B(u2_u0_b2_last_row_5_), .Y(u2_u0__abc_47660_n222) );
  OR2X2 OR2X2_2789 ( .A(u2_u0__abc_47660_n207), .B(row_adr_5_bF_buf3), .Y(u2_u0__abc_47660_n223) );
  OR2X2 OR2X2_279 ( .A(u0__abc_49347_n1183_1_bF_buf2), .B(1'b0), .Y(u0__abc_49347_n1546) );
  OR2X2 OR2X2_2790 ( .A(u2_u0__abc_47660_n205), .B(u2_u0_b2_last_row_6_), .Y(u2_u0__abc_47660_n225) );
  OR2X2 OR2X2_2791 ( .A(u2_u0__abc_47660_n207), .B(row_adr_6_bF_buf3), .Y(u2_u0__abc_47660_n226) );
  OR2X2 OR2X2_2792 ( .A(u2_u0__abc_47660_n205), .B(u2_u0_b2_last_row_7_), .Y(u2_u0__abc_47660_n228) );
  OR2X2 OR2X2_2793 ( .A(u2_u0__abc_47660_n207), .B(row_adr_7_bF_buf3), .Y(u2_u0__abc_47660_n229) );
  OR2X2 OR2X2_2794 ( .A(u2_u0__abc_47660_n205), .B(u2_u0_b2_last_row_8_), .Y(u2_u0__abc_47660_n231) );
  OR2X2 OR2X2_2795 ( .A(u2_u0__abc_47660_n207), .B(row_adr_8_bF_buf3), .Y(u2_u0__abc_47660_n232) );
  OR2X2 OR2X2_2796 ( .A(u2_u0__abc_47660_n205), .B(u2_u0_b2_last_row_9_), .Y(u2_u0__abc_47660_n234) );
  OR2X2 OR2X2_2797 ( .A(u2_u0__abc_47660_n207), .B(row_adr_9_bF_buf3), .Y(u2_u0__abc_47660_n235) );
  OR2X2 OR2X2_2798 ( .A(u2_u0__abc_47660_n205), .B(u2_u0_b2_last_row_10_), .Y(u2_u0__abc_47660_n237) );
  OR2X2 OR2X2_2799 ( .A(u2_u0__abc_47660_n207), .B(row_adr_10_bF_buf3), .Y(u2_u0__abc_47660_n238) );
  OR2X2 OR2X2_28 ( .A(lmr_sel_bF_buf0), .B(cs_6_), .Y(_abc_55805_n279) );
  OR2X2 OR2X2_280 ( .A(spec_req_cs_6_bF_buf5), .B(1'b0), .Y(u0__abc_49347_n1547) );
  OR2X2 OR2X2_2800 ( .A(u2_u0__abc_47660_n205), .B(u2_u0_b2_last_row_11_), .Y(u2_u0__abc_47660_n240) );
  OR2X2 OR2X2_2801 ( .A(u2_u0__abc_47660_n207), .B(row_adr_11_bF_buf3), .Y(u2_u0__abc_47660_n241) );
  OR2X2 OR2X2_2802 ( .A(u2_u0__abc_47660_n205), .B(u2_u0_b2_last_row_12_), .Y(u2_u0__abc_47660_n243) );
  OR2X2 OR2X2_2803 ( .A(u2_u0__abc_47660_n207), .B(row_adr_12_bF_buf3), .Y(u2_u0__abc_47660_n244) );
  OR2X2 OR2X2_2804 ( .A(u2_u0__abc_47660_n248), .B(u2_u0_b1_last_row_0_), .Y(u2_u0__abc_47660_n249) );
  OR2X2 OR2X2_2805 ( .A(u2_u0__abc_47660_n250), .B(row_adr_0_bF_buf2), .Y(u2_u0__abc_47660_n251) );
  OR2X2 OR2X2_2806 ( .A(u2_u0__abc_47660_n248), .B(u2_u0_b1_last_row_1_), .Y(u2_u0__abc_47660_n253) );
  OR2X2 OR2X2_2807 ( .A(u2_u0__abc_47660_n250), .B(row_adr_1_bF_buf2), .Y(u2_u0__abc_47660_n254) );
  OR2X2 OR2X2_2808 ( .A(u2_u0__abc_47660_n248), .B(u2_u0_b1_last_row_2_), .Y(u2_u0__abc_47660_n256) );
  OR2X2 OR2X2_2809 ( .A(u2_u0__abc_47660_n250), .B(row_adr_2_bF_buf2), .Y(u2_u0__abc_47660_n257) );
  OR2X2 OR2X2_281 ( .A(u0__abc_49347_n1549), .B(u0__abc_49347_n1545), .Y(u0__abc_49347_n1550) );
  OR2X2 OR2X2_2810 ( .A(u2_u0__abc_47660_n248), .B(u2_u0_b1_last_row_3_), .Y(u2_u0__abc_47660_n259) );
  OR2X2 OR2X2_2811 ( .A(u2_u0__abc_47660_n250), .B(row_adr_3_bF_buf2), .Y(u2_u0__abc_47660_n260) );
  OR2X2 OR2X2_2812 ( .A(u2_u0__abc_47660_n248), .B(u2_u0_b1_last_row_4_), .Y(u2_u0__abc_47660_n262) );
  OR2X2 OR2X2_2813 ( .A(u2_u0__abc_47660_n250), .B(row_adr_4_bF_buf2), .Y(u2_u0__abc_47660_n263) );
  OR2X2 OR2X2_2814 ( .A(u2_u0__abc_47660_n248), .B(u2_u0_b1_last_row_5_), .Y(u2_u0__abc_47660_n265) );
  OR2X2 OR2X2_2815 ( .A(u2_u0__abc_47660_n250), .B(row_adr_5_bF_buf2), .Y(u2_u0__abc_47660_n266) );
  OR2X2 OR2X2_2816 ( .A(u2_u0__abc_47660_n248), .B(u2_u0_b1_last_row_6_), .Y(u2_u0__abc_47660_n268) );
  OR2X2 OR2X2_2817 ( .A(u2_u0__abc_47660_n250), .B(row_adr_6_bF_buf2), .Y(u2_u0__abc_47660_n269) );
  OR2X2 OR2X2_2818 ( .A(u2_u0__abc_47660_n248), .B(u2_u0_b1_last_row_7_), .Y(u2_u0__abc_47660_n271) );
  OR2X2 OR2X2_2819 ( .A(u2_u0__abc_47660_n250), .B(row_adr_7_bF_buf2), .Y(u2_u0__abc_47660_n272) );
  OR2X2 OR2X2_282 ( .A(u0__abc_49347_n1551_1), .B(u0__abc_49347_n1552_1), .Y(u0__abc_49347_n1553) );
  OR2X2 OR2X2_2820 ( .A(u2_u0__abc_47660_n248), .B(u2_u0_b1_last_row_8_), .Y(u2_u0__abc_47660_n274) );
  OR2X2 OR2X2_2821 ( .A(u2_u0__abc_47660_n250), .B(row_adr_8_bF_buf2), .Y(u2_u0__abc_47660_n275_1) );
  OR2X2 OR2X2_2822 ( .A(u2_u0__abc_47660_n248), .B(u2_u0_b1_last_row_9_), .Y(u2_u0__abc_47660_n277) );
  OR2X2 OR2X2_2823 ( .A(u2_u0__abc_47660_n250), .B(row_adr_9_bF_buf2), .Y(u2_u0__abc_47660_n278_1) );
  OR2X2 OR2X2_2824 ( .A(u2_u0__abc_47660_n248), .B(u2_u0_b1_last_row_10_), .Y(u2_u0__abc_47660_n280) );
  OR2X2 OR2X2_2825 ( .A(u2_u0__abc_47660_n250), .B(row_adr_10_bF_buf2), .Y(u2_u0__abc_47660_n281) );
  OR2X2 OR2X2_2826 ( .A(u2_u0__abc_47660_n248), .B(u2_u0_b1_last_row_11_), .Y(u2_u0__abc_47660_n283_1) );
  OR2X2 OR2X2_2827 ( .A(u2_u0__abc_47660_n250), .B(row_adr_11_bF_buf2), .Y(u2_u0__abc_47660_n284) );
  OR2X2 OR2X2_2828 ( .A(u2_u0__abc_47660_n248), .B(u2_u0_b1_last_row_12_), .Y(u2_u0__abc_47660_n286_1) );
  OR2X2 OR2X2_2829 ( .A(u2_u0__abc_47660_n250), .B(row_adr_12_bF_buf2), .Y(u2_u0__abc_47660_n287_1) );
  OR2X2 OR2X2_283 ( .A(u0__abc_49347_n1554), .B(u0__abc_49347_n1555), .Y(u0__abc_49347_n1556) );
  OR2X2 OR2X2_2830 ( .A(u2_u0__abc_47660_n290_1), .B(u2_u0_b0_last_row_0_), .Y(u2_u0__abc_47660_n291) );
  OR2X2 OR2X2_2831 ( .A(u2_u0__abc_47660_n292_1), .B(row_adr_0_bF_buf1), .Y(u2_u0__abc_47660_n293) );
  OR2X2 OR2X2_2832 ( .A(u2_u0__abc_47660_n290_1), .B(u2_u0_b0_last_row_1_), .Y(u2_u0__abc_47660_n295) );
  OR2X2 OR2X2_2833 ( .A(u2_u0__abc_47660_n292_1), .B(row_adr_1_bF_buf1), .Y(u2_u0__abc_47660_n296_1) );
  OR2X2 OR2X2_2834 ( .A(u2_u0__abc_47660_n290_1), .B(u2_u0_b0_last_row_2_), .Y(u2_u0__abc_47660_n298) );
  OR2X2 OR2X2_2835 ( .A(u2_u0__abc_47660_n292_1), .B(row_adr_2_bF_buf1), .Y(u2_u0__abc_47660_n299) );
  OR2X2 OR2X2_2836 ( .A(u2_u0__abc_47660_n290_1), .B(u2_u0_b0_last_row_3_), .Y(u2_u0__abc_47660_n301) );
  OR2X2 OR2X2_2837 ( .A(u2_u0__abc_47660_n292_1), .B(row_adr_3_bF_buf1), .Y(u2_u0__abc_47660_n302) );
  OR2X2 OR2X2_2838 ( .A(u2_u0__abc_47660_n290_1), .B(u2_u0_b0_last_row_4_), .Y(u2_u0__abc_47660_n304_1) );
  OR2X2 OR2X2_2839 ( .A(u2_u0__abc_47660_n292_1), .B(row_adr_4_bF_buf1), .Y(u2_u0__abc_47660_n305_1) );
  OR2X2 OR2X2_284 ( .A(u0__abc_49347_n1557), .B(u0__abc_49347_n1558), .Y(u0__abc_49347_n1559) );
  OR2X2 OR2X2_2840 ( .A(u2_u0__abc_47660_n290_1), .B(u2_u0_b0_last_row_5_), .Y(u2_u0__abc_47660_n307) );
  OR2X2 OR2X2_2841 ( .A(u2_u0__abc_47660_n292_1), .B(row_adr_5_bF_buf1), .Y(u2_u0__abc_47660_n308) );
  OR2X2 OR2X2_2842 ( .A(u2_u0__abc_47660_n290_1), .B(u2_u0_b0_last_row_6_), .Y(u2_u0__abc_47660_n310) );
  OR2X2 OR2X2_2843 ( .A(u2_u0__abc_47660_n292_1), .B(row_adr_6_bF_buf1), .Y(u2_u0__abc_47660_n311) );
  OR2X2 OR2X2_2844 ( .A(u2_u0__abc_47660_n290_1), .B(u2_u0_b0_last_row_7_), .Y(u2_u0__abc_47660_n313) );
  OR2X2 OR2X2_2845 ( .A(u2_u0__abc_47660_n292_1), .B(row_adr_7_bF_buf1), .Y(u2_u0__abc_47660_n314) );
  OR2X2 OR2X2_2846 ( .A(u2_u0__abc_47660_n290_1), .B(u2_u0_b0_last_row_8_), .Y(u2_u0__abc_47660_n316) );
  OR2X2 OR2X2_2847 ( .A(u2_u0__abc_47660_n292_1), .B(row_adr_8_bF_buf1), .Y(u2_u0__abc_47660_n317) );
  OR2X2 OR2X2_2848 ( .A(u2_u0__abc_47660_n290_1), .B(u2_u0_b0_last_row_9_), .Y(u2_u0__abc_47660_n319) );
  OR2X2 OR2X2_2849 ( .A(u2_u0__abc_47660_n292_1), .B(row_adr_9_bF_buf1), .Y(u2_u0__abc_47660_n320) );
  OR2X2 OR2X2_285 ( .A(u0__abc_49347_n1561_1), .B(spec_req_cs_0_bF_buf5), .Y(u0__abc_49347_n1562) );
  OR2X2 OR2X2_2850 ( .A(u2_u0__abc_47660_n290_1), .B(u2_u0_b0_last_row_10_), .Y(u2_u0__abc_47660_n322) );
  OR2X2 OR2X2_2851 ( .A(u2_u0__abc_47660_n292_1), .B(row_adr_10_bF_buf1), .Y(u2_u0__abc_47660_n323) );
  OR2X2 OR2X2_2852 ( .A(u2_u0__abc_47660_n290_1), .B(u2_u0_b0_last_row_11_), .Y(u2_u0__abc_47660_n325) );
  OR2X2 OR2X2_2853 ( .A(u2_u0__abc_47660_n292_1), .B(row_adr_11_bF_buf1), .Y(u2_u0__abc_47660_n326) );
  OR2X2 OR2X2_2854 ( .A(u2_u0__abc_47660_n290_1), .B(u2_u0_b0_last_row_12_), .Y(u2_u0__abc_47660_n328) );
  OR2X2 OR2X2_2855 ( .A(u2_u0__abc_47660_n292_1), .B(row_adr_12_bF_buf1), .Y(u2_u0__abc_47660_n329) );
  OR2X2 OR2X2_2856 ( .A(u2_u0__abc_47660_n331), .B(row_adr_12_bF_buf0), .Y(u2_u0__abc_47660_n332) );
  OR2X2 OR2X2_2857 ( .A(u2_u0__abc_47660_n333), .B(row_adr_11_bF_buf0), .Y(u2_u0__abc_47660_n334) );
  OR2X2 OR2X2_2858 ( .A(u2_u0__abc_47660_n199), .B(u2_u0_b0_last_row_12_), .Y(u2_u0__abc_47660_n335) );
  OR2X2 OR2X2_2859 ( .A(u2_u0__abc_47660_n194), .B(u2_u0_b0_last_row_11_), .Y(u2_u0__abc_47660_n338) );
  OR2X2 OR2X2_286 ( .A(u0__abc_49347_n1560_1), .B(u0__abc_49347_n1562), .Y(u0__abc_49347_n1563) );
  OR2X2 OR2X2_2860 ( .A(u2_u0__abc_47660_n339), .B(row_adr_9_bF_buf0), .Y(u2_u0__abc_47660_n340) );
  OR2X2 OR2X2_2861 ( .A(u2_u0__abc_47660_n184), .B(u2_u0_b0_last_row_9_), .Y(u2_u0__abc_47660_n342) );
  OR2X2 OR2X2_2862 ( .A(u2_u0__abc_47660_n343), .B(row_adr_7_bF_buf0), .Y(u2_u0__abc_47660_n344) );
  OR2X2 OR2X2_2863 ( .A(u2_u0__abc_47660_n164), .B(u2_u0_b0_last_row_5_), .Y(u2_u0__abc_47660_n348) );
  OR2X2 OR2X2_2864 ( .A(u2_u0__abc_47660_n159), .B(u2_u0_b0_last_row_4_), .Y(u2_u0__abc_47660_n350) );
  OR2X2 OR2X2_2865 ( .A(u2_u0__abc_47660_n351), .B(row_adr_4_bF_buf0), .Y(u2_u0__abc_47660_n352) );
  OR2X2 OR2X2_2866 ( .A(u2_u0__abc_47660_n355), .B(row_adr_0_bF_buf0), .Y(u2_u0__abc_47660_n356) );
  OR2X2 OR2X2_2867 ( .A(u2_u0__abc_47660_n139), .B(u2_u0_b0_last_row_0_), .Y(u2_u0__abc_47660_n357) );
  OR2X2 OR2X2_2868 ( .A(u2_u0__abc_47660_n144), .B(u2_u0_b0_last_row_1_), .Y(u2_u0__abc_47660_n359) );
  OR2X2 OR2X2_2869 ( .A(u2_u0__abc_47660_n360), .B(row_adr_5_bF_buf0), .Y(u2_u0__abc_47660_n361) );
  OR2X2 OR2X2_287 ( .A(u0__abc_49347_n1203_bF_buf2), .B(u0_tms0_15_), .Y(u0__abc_49347_n1564) );
  OR2X2 OR2X2_2870 ( .A(u2_u0__abc_47660_n366), .B(row_adr_10_bF_buf0), .Y(u2_u0__abc_47660_n367) );
  OR2X2 OR2X2_2871 ( .A(u2_u0__abc_47660_n189), .B(u2_u0_b0_last_row_10_), .Y(u2_u0__abc_47660_n368) );
  OR2X2 OR2X2_2872 ( .A(u2_u0__abc_47660_n372), .B(u2_u0__abc_47660_n370), .Y(u2_u0__abc_47660_n373) );
  OR2X2 OR2X2_2873 ( .A(u2_u0__abc_47660_n154), .B(u2_u0_b0_last_row_3_), .Y(u2_u0__abc_47660_n375) );
  OR2X2 OR2X2_2874 ( .A(u2_u0__abc_47660_n376), .B(row_adr_2_bF_buf0), .Y(u2_u0__abc_47660_n377) );
  OR2X2 OR2X2_2875 ( .A(u2_u0__abc_47660_n379), .B(row_adr_1_bF_buf0), .Y(u2_u0__abc_47660_n380) );
  OR2X2 OR2X2_2876 ( .A(u2_u0__abc_47660_n149), .B(u2_u0_b0_last_row_2_), .Y(u2_u0__abc_47660_n381) );
  OR2X2 OR2X2_2877 ( .A(u2_u0__abc_47660_n384), .B(row_adr_3_bF_buf0), .Y(u2_u0__abc_47660_n385) );
  OR2X2 OR2X2_2878 ( .A(u2_u0__abc_47660_n174), .B(u2_u0_b0_last_row_7_), .Y(u2_u0__abc_47660_n386) );
  OR2X2 OR2X2_2879 ( .A(u2_u0__abc_47660_n390), .B(u2_u0__abc_47660_n388), .Y(u2_u0__abc_47660_n391) );
  OR2X2 OR2X2_288 ( .A(u0__abc_49347_n1566), .B(u0__abc_49347_n1544), .Y(u0_sp_tms_15__FF_INPUT) );
  OR2X2 OR2X2_2880 ( .A(u2_u0__abc_47660_n396), .B(row_adr_12_bF_buf6), .Y(u2_u0__abc_47660_n397) );
  OR2X2 OR2X2_2881 ( .A(u2_u0__abc_47660_n398), .B(row_adr_11_bF_buf6), .Y(u2_u0__abc_47660_n399) );
  OR2X2 OR2X2_2882 ( .A(u2_u0__abc_47660_n199), .B(u2_u0_b2_last_row_12_), .Y(u2_u0__abc_47660_n400) );
  OR2X2 OR2X2_2883 ( .A(u2_u0__abc_47660_n194), .B(u2_u0_b2_last_row_11_), .Y(u2_u0__abc_47660_n403) );
  OR2X2 OR2X2_2884 ( .A(u2_u0__abc_47660_n404), .B(row_adr_9_bF_buf6), .Y(u2_u0__abc_47660_n405) );
  OR2X2 OR2X2_2885 ( .A(u2_u0__abc_47660_n184), .B(u2_u0_b2_last_row_9_), .Y(u2_u0__abc_47660_n407) );
  OR2X2 OR2X2_2886 ( .A(u2_u0__abc_47660_n408), .B(row_adr_7_bF_buf6), .Y(u2_u0__abc_47660_n409) );
  OR2X2 OR2X2_2887 ( .A(u2_u0__abc_47660_n164), .B(u2_u0_b2_last_row_5_), .Y(u2_u0__abc_47660_n413) );
  OR2X2 OR2X2_2888 ( .A(u2_u0__abc_47660_n159), .B(u2_u0_b2_last_row_4_), .Y(u2_u0__abc_47660_n415) );
  OR2X2 OR2X2_2889 ( .A(u2_u0__abc_47660_n416), .B(row_adr_4_bF_buf6), .Y(u2_u0__abc_47660_n417) );
  OR2X2 OR2X2_289 ( .A(u0__abc_49347_n1183_1_bF_buf1), .B(1'b0), .Y(u0__abc_49347_n1570_1) );
  OR2X2 OR2X2_2890 ( .A(u2_u0__abc_47660_n420), .B(row_adr_0_bF_buf6), .Y(u2_u0__abc_47660_n421) );
  OR2X2 OR2X2_2891 ( .A(u2_u0__abc_47660_n139), .B(u2_u0_b2_last_row_0_), .Y(u2_u0__abc_47660_n422) );
  OR2X2 OR2X2_2892 ( .A(u2_u0__abc_47660_n144), .B(u2_u0_b2_last_row_1_), .Y(u2_u0__abc_47660_n424) );
  OR2X2 OR2X2_2893 ( .A(u2_u0__abc_47660_n425), .B(row_adr_5_bF_buf6), .Y(u2_u0__abc_47660_n426) );
  OR2X2 OR2X2_2894 ( .A(u2_u0__abc_47660_n431), .B(row_adr_10_bF_buf6), .Y(u2_u0__abc_47660_n432) );
  OR2X2 OR2X2_2895 ( .A(u2_u0__abc_47660_n189), .B(u2_u0_b2_last_row_10_), .Y(u2_u0__abc_47660_n433) );
  OR2X2 OR2X2_2896 ( .A(u2_u0__abc_47660_n437), .B(u2_u0__abc_47660_n435), .Y(u2_u0__abc_47660_n438) );
  OR2X2 OR2X2_2897 ( .A(u2_u0__abc_47660_n154), .B(u2_u0_b2_last_row_3_), .Y(u2_u0__abc_47660_n440) );
  OR2X2 OR2X2_2898 ( .A(u2_u0__abc_47660_n441), .B(row_adr_2_bF_buf6), .Y(u2_u0__abc_47660_n442) );
  OR2X2 OR2X2_2899 ( .A(u2_u0__abc_47660_n444), .B(row_adr_1_bF_buf6), .Y(u2_u0__abc_47660_n445) );
  OR2X2 OR2X2_29 ( .A(_abc_55805_n280), .B(_abc_55805_n237_1), .Y(_abc_55805_n281) );
  OR2X2 OR2X2_290 ( .A(spec_req_cs_6_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n1571) );
  OR2X2 OR2X2_2900 ( .A(u2_u0__abc_47660_n149), .B(u2_u0_b2_last_row_2_), .Y(u2_u0__abc_47660_n446) );
  OR2X2 OR2X2_2901 ( .A(u2_u0__abc_47660_n449), .B(row_adr_3_bF_buf6), .Y(u2_u0__abc_47660_n450) );
  OR2X2 OR2X2_2902 ( .A(u2_u0__abc_47660_n174), .B(u2_u0_b2_last_row_7_), .Y(u2_u0__abc_47660_n451) );
  OR2X2 OR2X2_2903 ( .A(u2_u0__abc_47660_n455), .B(u2_u0__abc_47660_n453), .Y(u2_u0__abc_47660_n456) );
  OR2X2 OR2X2_2904 ( .A(u2_u0__abc_47660_n395), .B(u2_u0__abc_47660_n460), .Y(u2_u0__abc_47660_n461) );
  OR2X2 OR2X2_2905 ( .A(u2_u0__abc_47660_n462), .B(row_adr_12_bF_buf5), .Y(u2_u0__abc_47660_n463) );
  OR2X2 OR2X2_2906 ( .A(u2_u0__abc_47660_n464), .B(row_adr_11_bF_buf5), .Y(u2_u0__abc_47660_n465) );
  OR2X2 OR2X2_2907 ( .A(u2_u0__abc_47660_n199), .B(u2_u0_b1_last_row_12_), .Y(u2_u0__abc_47660_n466) );
  OR2X2 OR2X2_2908 ( .A(u2_u0__abc_47660_n194), .B(u2_u0_b1_last_row_11_), .Y(u2_u0__abc_47660_n469) );
  OR2X2 OR2X2_2909 ( .A(u2_u0__abc_47660_n470), .B(row_adr_9_bF_buf5), .Y(u2_u0__abc_47660_n471) );
  OR2X2 OR2X2_291 ( .A(u0__abc_49347_n1573), .B(u0__abc_49347_n1569_1), .Y(u0__abc_49347_n1574) );
  OR2X2 OR2X2_2910 ( .A(u2_u0__abc_47660_n184), .B(u2_u0_b1_last_row_9_), .Y(u2_u0__abc_47660_n473) );
  OR2X2 OR2X2_2911 ( .A(u2_u0__abc_47660_n474), .B(row_adr_7_bF_buf5), .Y(u2_u0__abc_47660_n475) );
  OR2X2 OR2X2_2912 ( .A(u2_u0__abc_47660_n164), .B(u2_u0_b1_last_row_5_), .Y(u2_u0__abc_47660_n479) );
  OR2X2 OR2X2_2913 ( .A(u2_u0__abc_47660_n159), .B(u2_u0_b1_last_row_4_), .Y(u2_u0__abc_47660_n481) );
  OR2X2 OR2X2_2914 ( .A(u2_u0__abc_47660_n482), .B(row_adr_4_bF_buf5), .Y(u2_u0__abc_47660_n483) );
  OR2X2 OR2X2_2915 ( .A(u2_u0__abc_47660_n486), .B(row_adr_0_bF_buf5), .Y(u2_u0__abc_47660_n487) );
  OR2X2 OR2X2_2916 ( .A(u2_u0__abc_47660_n139), .B(u2_u0_b1_last_row_0_), .Y(u2_u0__abc_47660_n488) );
  OR2X2 OR2X2_2917 ( .A(u2_u0__abc_47660_n144), .B(u2_u0_b1_last_row_1_), .Y(u2_u0__abc_47660_n490) );
  OR2X2 OR2X2_2918 ( .A(u2_u0__abc_47660_n491), .B(row_adr_5_bF_buf5), .Y(u2_u0__abc_47660_n492) );
  OR2X2 OR2X2_2919 ( .A(u2_u0__abc_47660_n497), .B(row_adr_10_bF_buf5), .Y(u2_u0__abc_47660_n498) );
  OR2X2 OR2X2_292 ( .A(u0__abc_49347_n1575), .B(u0__abc_49347_n1576), .Y(u0__abc_49347_n1577) );
  OR2X2 OR2X2_2920 ( .A(u2_u0__abc_47660_n189), .B(u2_u0_b1_last_row_10_), .Y(u2_u0__abc_47660_n499) );
  OR2X2 OR2X2_2921 ( .A(u2_u0__abc_47660_n503), .B(u2_u0__abc_47660_n501), .Y(u2_u0__abc_47660_n504) );
  OR2X2 OR2X2_2922 ( .A(u2_u0__abc_47660_n154), .B(u2_u0_b1_last_row_3_), .Y(u2_u0__abc_47660_n506) );
  OR2X2 OR2X2_2923 ( .A(u2_u0__abc_47660_n507), .B(row_adr_2_bF_buf5), .Y(u2_u0__abc_47660_n508) );
  OR2X2 OR2X2_2924 ( .A(u2_u0__abc_47660_n510), .B(row_adr_1_bF_buf5), .Y(u2_u0__abc_47660_n511) );
  OR2X2 OR2X2_2925 ( .A(u2_u0__abc_47660_n149), .B(u2_u0_b1_last_row_2_), .Y(u2_u0__abc_47660_n512) );
  OR2X2 OR2X2_2926 ( .A(u2_u0__abc_47660_n515), .B(row_adr_3_bF_buf5), .Y(u2_u0__abc_47660_n516) );
  OR2X2 OR2X2_2927 ( .A(u2_u0__abc_47660_n174), .B(u2_u0_b1_last_row_7_), .Y(u2_u0__abc_47660_n517) );
  OR2X2 OR2X2_2928 ( .A(u2_u0__abc_47660_n521), .B(u2_u0__abc_47660_n519), .Y(u2_u0__abc_47660_n522) );
  OR2X2 OR2X2_2929 ( .A(u2_u0__abc_47660_n527), .B(row_adr_9_bF_buf4), .Y(u2_u0__abc_47660_n528) );
  OR2X2 OR2X2_293 ( .A(u0__abc_49347_n1578_1), .B(u0__abc_49347_n1579_1), .Y(u0__abc_49347_n1580) );
  OR2X2 OR2X2_2930 ( .A(u2_u0__abc_47660_n189), .B(u2_u0_b3_last_row_10_), .Y(u2_u0__abc_47660_n529) );
  OR2X2 OR2X2_2931 ( .A(u2_u0__abc_47660_n184), .B(u2_u0_b3_last_row_9_), .Y(u2_u0__abc_47660_n530) );
  OR2X2 OR2X2_2932 ( .A(u2_u0__abc_47660_n194), .B(u2_u0_b3_last_row_11_), .Y(u2_u0__abc_47660_n533) );
  OR2X2 OR2X2_2933 ( .A(u2_u0__abc_47660_n534), .B(row_adr_11_bF_buf4), .Y(u2_u0__abc_47660_n535) );
  OR2X2 OR2X2_2934 ( .A(u2_u0__abc_47660_n199), .B(u2_u0_b3_last_row_12_), .Y(u2_u0__abc_47660_n537) );
  OR2X2 OR2X2_2935 ( .A(u2_u0__abc_47660_n538), .B(row_adr_8_bF_buf4), .Y(u2_u0__abc_47660_n539) );
  OR2X2 OR2X2_2936 ( .A(u2_u0__abc_47660_n159), .B(u2_u0_b3_last_row_4_), .Y(u2_u0__abc_47660_n543) );
  OR2X2 OR2X2_2937 ( .A(u2_u0__abc_47660_n544), .B(row_adr_4_bF_buf4), .Y(u2_u0__abc_47660_n545) );
  OR2X2 OR2X2_2938 ( .A(u2_u0__abc_47660_n547), .B(row_adr_3_bF_buf4), .Y(u2_u0__abc_47660_n548) );
  OR2X2 OR2X2_2939 ( .A(u2_u0__abc_47660_n551), .B(row_adr_0_bF_buf4), .Y(u2_u0__abc_47660_n552) );
  OR2X2 OR2X2_294 ( .A(u0__abc_49347_n1581), .B(u0__abc_49347_n1582), .Y(u0__abc_49347_n1583) );
  OR2X2 OR2X2_2940 ( .A(u2_u0__abc_47660_n139), .B(u2_u0_b3_last_row_0_), .Y(u2_u0__abc_47660_n553) );
  OR2X2 OR2X2_2941 ( .A(u2_u0__abc_47660_n555), .B(row_adr_2_bF_buf4), .Y(u2_u0__abc_47660_n556) );
  OR2X2 OR2X2_2942 ( .A(u2_u0__abc_47660_n149), .B(u2_u0_b3_last_row_2_), .Y(u2_u0__abc_47660_n557) );
  OR2X2 OR2X2_2943 ( .A(u2_u0__abc_47660_n174), .B(u2_u0_b3_last_row_7_), .Y(u2_u0__abc_47660_n562) );
  OR2X2 OR2X2_2944 ( .A(u2_u0__abc_47660_n563), .B(row_adr_7_bF_buf4), .Y(u2_u0__abc_47660_n564) );
  OR2X2 OR2X2_2945 ( .A(u2_u0__abc_47660_n566), .B(row_adr_10_bF_buf4), .Y(u2_u0__abc_47660_n567) );
  OR2X2 OR2X2_2946 ( .A(u2_u0__abc_47660_n179), .B(u2_u0_b3_last_row_8_), .Y(u2_u0__abc_47660_n568) );
  OR2X2 OR2X2_2947 ( .A(u2_u0__abc_47660_n169), .B(u2_u0_b3_last_row_6_), .Y(u2_u0__abc_47660_n571) );
  OR2X2 OR2X2_2948 ( .A(u2_u0__abc_47660_n572), .B(row_adr_6_bF_buf4), .Y(u2_u0__abc_47660_n573) );
  OR2X2 OR2X2_2949 ( .A(u2_u0__abc_47660_n575), .B(row_adr_5_bF_buf4), .Y(u2_u0__abc_47660_n576) );
  OR2X2 OR2X2_295 ( .A(u0__abc_49347_n1585), .B(spec_req_cs_0_bF_buf4), .Y(u0__abc_49347_n1586) );
  OR2X2 OR2X2_2950 ( .A(u2_u0__abc_47660_n154), .B(u2_u0_b3_last_row_3_), .Y(u2_u0__abc_47660_n577) );
  OR2X2 OR2X2_2951 ( .A(u2_u0__abc_47660_n164), .B(u2_u0_b3_last_row_5_), .Y(u2_u0__abc_47660_n580) );
  OR2X2 OR2X2_2952 ( .A(u2_u0__abc_47660_n581), .B(row_adr_1_bF_buf4), .Y(u2_u0__abc_47660_n582) );
  OR2X2 OR2X2_2953 ( .A(u2_u0__abc_47660_n144), .B(u2_u0_b3_last_row_1_), .Y(u2_u0__abc_47660_n584) );
  OR2X2 OR2X2_2954 ( .A(u2_u0__abc_47660_n585), .B(row_adr_12_bF_buf4), .Y(u2_u0__abc_47660_n586) );
  OR2X2 OR2X2_2955 ( .A(u2_u0__abc_47660_n526), .B(u2_u0__abc_47660_n591), .Y(u2_u0__abc_47660_n592) );
  OR2X2 OR2X2_2956 ( .A(u2_u0__abc_47660_n461), .B(u2_u0__abc_47660_n592), .Y(u2_row_same_0) );
  OR2X2 OR2X2_2957 ( .A(u2_u0__abc_47660_n594), .B(u2_u0__abc_47660_n595), .Y(u2_u0__abc_47660_n596) );
  OR2X2 OR2X2_2958 ( .A(u2_u0__abc_47660_n598), .B(u2_u0__abc_47660_n597), .Y(u2_u0__abc_47660_n599) );
  OR2X2 OR2X2_2959 ( .A(u2_u0__abc_47660_n596), .B(u2_u0__abc_47660_n599), .Y(u2_bank_open_0) );
  OR2X2 OR2X2_296 ( .A(u0__abc_49347_n1584), .B(u0__abc_49347_n1586), .Y(u0__abc_49347_n1587_1) );
  OR2X2 OR2X2_2960 ( .A(u2_u0__abc_47660_n608), .B(u2_u0__abc_47660_n137_bF_buf3), .Y(u2_u0_bank3_open_FF_INPUT) );
  OR2X2 OR2X2_2961 ( .A(u2_u0__abc_47660_n611), .B(u2_u0__abc_47660_n610), .Y(u2_u0__abc_47660_n612) );
  OR2X2 OR2X2_2962 ( .A(u2_u0__abc_47660_n614), .B(u2_u0__abc_47660_n205), .Y(u2_u0_bank2_open_FF_INPUT) );
  OR2X2 OR2X2_2963 ( .A(u2_u0__abc_47660_n616), .B(u2_u0__abc_47660_n610), .Y(u2_u0__abc_47660_n617) );
  OR2X2 OR2X2_2964 ( .A(u2_u0__abc_47660_n619), .B(u2_u0__abc_47660_n248), .Y(u2_u0_bank1_open_FF_INPUT) );
  OR2X2 OR2X2_2965 ( .A(u2_u0__abc_47660_n621), .B(u2_u0__abc_47660_n610), .Y(u2_u0__abc_47660_n622) );
  OR2X2 OR2X2_2966 ( .A(u2_u0__abc_47660_n624), .B(u2_u0__abc_47660_n290_1), .Y(u2_u0_bank0_open_FF_INPUT) );
  OR2X2 OR2X2_2967 ( .A(u2_u1__abc_47660_n137_bF_buf4), .B(u2_u1_b3_last_row_0_), .Y(u2_u1__abc_47660_n138) );
  OR2X2 OR2X2_2968 ( .A(u2_u1__abc_47660_n137_bF_buf2), .B(u2_u1_b3_last_row_1_), .Y(u2_u1__abc_47660_n143) );
  OR2X2 OR2X2_2969 ( .A(u2_u1__abc_47660_n137_bF_buf0), .B(u2_u1_b3_last_row_2_), .Y(u2_u1__abc_47660_n148) );
  OR2X2 OR2X2_297 ( .A(u0__abc_49347_n1203_bF_buf1), .B(u0_tms0_16_), .Y(u0__abc_49347_n1588_1) );
  OR2X2 OR2X2_2970 ( .A(u2_u1__abc_47660_n137_bF_buf3), .B(u2_u1_b3_last_row_3_), .Y(u2_u1__abc_47660_n153) );
  OR2X2 OR2X2_2971 ( .A(u2_u1__abc_47660_n137_bF_buf1), .B(u2_u1_b3_last_row_4_), .Y(u2_u1__abc_47660_n158) );
  OR2X2 OR2X2_2972 ( .A(u2_u1__abc_47660_n137_bF_buf4), .B(u2_u1_b3_last_row_5_), .Y(u2_u1__abc_47660_n163) );
  OR2X2 OR2X2_2973 ( .A(u2_u1__abc_47660_n137_bF_buf2), .B(u2_u1_b3_last_row_6_), .Y(u2_u1__abc_47660_n168) );
  OR2X2 OR2X2_2974 ( .A(u2_u1__abc_47660_n137_bF_buf0), .B(u2_u1_b3_last_row_7_), .Y(u2_u1__abc_47660_n173) );
  OR2X2 OR2X2_2975 ( .A(u2_u1__abc_47660_n137_bF_buf3), .B(u2_u1_b3_last_row_8_), .Y(u2_u1__abc_47660_n178) );
  OR2X2 OR2X2_2976 ( .A(u2_u1__abc_47660_n137_bF_buf1), .B(u2_u1_b3_last_row_9_), .Y(u2_u1__abc_47660_n183) );
  OR2X2 OR2X2_2977 ( .A(u2_u1__abc_47660_n137_bF_buf4), .B(u2_u1_b3_last_row_10_), .Y(u2_u1__abc_47660_n188) );
  OR2X2 OR2X2_2978 ( .A(u2_u1__abc_47660_n137_bF_buf2), .B(u2_u1_b3_last_row_11_), .Y(u2_u1__abc_47660_n193) );
  OR2X2 OR2X2_2979 ( .A(u2_u1__abc_47660_n137_bF_buf0), .B(u2_u1_b3_last_row_12_), .Y(u2_u1__abc_47660_n198) );
  OR2X2 OR2X2_298 ( .A(u0__abc_49347_n1590), .B(u0__abc_49347_n1568), .Y(u0_sp_tms_16__FF_INPUT) );
  OR2X2 OR2X2_2980 ( .A(u2_u1__abc_47660_n205), .B(u2_u1_b2_last_row_0_), .Y(u2_u1__abc_47660_n206) );
  OR2X2 OR2X2_2981 ( .A(u2_u1__abc_47660_n207), .B(row_adr_0_bF_buf2), .Y(u2_u1__abc_47660_n208) );
  OR2X2 OR2X2_2982 ( .A(u2_u1__abc_47660_n205), .B(u2_u1_b2_last_row_1_), .Y(u2_u1__abc_47660_n210) );
  OR2X2 OR2X2_2983 ( .A(u2_u1__abc_47660_n207), .B(row_adr_1_bF_buf2), .Y(u2_u1__abc_47660_n211) );
  OR2X2 OR2X2_2984 ( .A(u2_u1__abc_47660_n205), .B(u2_u1_b2_last_row_2_), .Y(u2_u1__abc_47660_n213) );
  OR2X2 OR2X2_2985 ( .A(u2_u1__abc_47660_n207), .B(row_adr_2_bF_buf2), .Y(u2_u1__abc_47660_n214) );
  OR2X2 OR2X2_2986 ( .A(u2_u1__abc_47660_n205), .B(u2_u1_b2_last_row_3_), .Y(u2_u1__abc_47660_n216) );
  OR2X2 OR2X2_2987 ( .A(u2_u1__abc_47660_n207), .B(row_adr_3_bF_buf2), .Y(u2_u1__abc_47660_n217) );
  OR2X2 OR2X2_2988 ( .A(u2_u1__abc_47660_n205), .B(u2_u1_b2_last_row_4_), .Y(u2_u1__abc_47660_n219) );
  OR2X2 OR2X2_2989 ( .A(u2_u1__abc_47660_n207), .B(row_adr_4_bF_buf2), .Y(u2_u1__abc_47660_n220) );
  OR2X2 OR2X2_299 ( .A(u0__abc_49347_n1183_1_bF_buf0), .B(1'b0), .Y(u0__abc_49347_n1594) );
  OR2X2 OR2X2_2990 ( .A(u2_u1__abc_47660_n205), .B(u2_u1_b2_last_row_5_), .Y(u2_u1__abc_47660_n222) );
  OR2X2 OR2X2_2991 ( .A(u2_u1__abc_47660_n207), .B(row_adr_5_bF_buf2), .Y(u2_u1__abc_47660_n223) );
  OR2X2 OR2X2_2992 ( .A(u2_u1__abc_47660_n205), .B(u2_u1_b2_last_row_6_), .Y(u2_u1__abc_47660_n225) );
  OR2X2 OR2X2_2993 ( .A(u2_u1__abc_47660_n207), .B(row_adr_6_bF_buf2), .Y(u2_u1__abc_47660_n226) );
  OR2X2 OR2X2_2994 ( .A(u2_u1__abc_47660_n205), .B(u2_u1_b2_last_row_7_), .Y(u2_u1__abc_47660_n228) );
  OR2X2 OR2X2_2995 ( .A(u2_u1__abc_47660_n207), .B(row_adr_7_bF_buf2), .Y(u2_u1__abc_47660_n229) );
  OR2X2 OR2X2_2996 ( .A(u2_u1__abc_47660_n205), .B(u2_u1_b2_last_row_8_), .Y(u2_u1__abc_47660_n231) );
  OR2X2 OR2X2_2997 ( .A(u2_u1__abc_47660_n207), .B(row_adr_8_bF_buf2), .Y(u2_u1__abc_47660_n232) );
  OR2X2 OR2X2_2998 ( .A(u2_u1__abc_47660_n205), .B(u2_u1_b2_last_row_9_), .Y(u2_u1__abc_47660_n234) );
  OR2X2 OR2X2_2999 ( .A(u2_u1__abc_47660_n207), .B(row_adr_9_bF_buf2), .Y(u2_u1__abc_47660_n235) );
  OR2X2 OR2X2_3 ( .A(_abc_55805_n240_bF_buf5), .B(spec_req_cs_0_bF_buf5), .Y(_abc_55805_n241_1) );
  OR2X2 OR2X2_30 ( .A(_abc_55805_n245_1), .B(cs_need_rfr_6_), .Y(_abc_55805_n282) );
  OR2X2 OR2X2_300 ( .A(spec_req_cs_6_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n1595) );
  OR2X2 OR2X2_3000 ( .A(u2_u1__abc_47660_n205), .B(u2_u1_b2_last_row_10_), .Y(u2_u1__abc_47660_n237) );
  OR2X2 OR2X2_3001 ( .A(u2_u1__abc_47660_n207), .B(row_adr_10_bF_buf2), .Y(u2_u1__abc_47660_n238) );
  OR2X2 OR2X2_3002 ( .A(u2_u1__abc_47660_n205), .B(u2_u1_b2_last_row_11_), .Y(u2_u1__abc_47660_n240) );
  OR2X2 OR2X2_3003 ( .A(u2_u1__abc_47660_n207), .B(row_adr_11_bF_buf2), .Y(u2_u1__abc_47660_n241) );
  OR2X2 OR2X2_3004 ( .A(u2_u1__abc_47660_n205), .B(u2_u1_b2_last_row_12_), .Y(u2_u1__abc_47660_n243) );
  OR2X2 OR2X2_3005 ( .A(u2_u1__abc_47660_n207), .B(row_adr_12_bF_buf2), .Y(u2_u1__abc_47660_n244) );
  OR2X2 OR2X2_3006 ( .A(u2_u1__abc_47660_n248), .B(u2_u1_b1_last_row_0_), .Y(u2_u1__abc_47660_n249) );
  OR2X2 OR2X2_3007 ( .A(u2_u1__abc_47660_n250), .B(row_adr_0_bF_buf1), .Y(u2_u1__abc_47660_n251) );
  OR2X2 OR2X2_3008 ( .A(u2_u1__abc_47660_n248), .B(u2_u1_b1_last_row_1_), .Y(u2_u1__abc_47660_n253) );
  OR2X2 OR2X2_3009 ( .A(u2_u1__abc_47660_n250), .B(row_adr_1_bF_buf1), .Y(u2_u1__abc_47660_n254) );
  OR2X2 OR2X2_301 ( .A(u0__abc_49347_n1597_1), .B(u0__abc_49347_n1593), .Y(u0__abc_49347_n1598) );
  OR2X2 OR2X2_3010 ( .A(u2_u1__abc_47660_n248), .B(u2_u1_b1_last_row_2_), .Y(u2_u1__abc_47660_n256) );
  OR2X2 OR2X2_3011 ( .A(u2_u1__abc_47660_n250), .B(row_adr_2_bF_buf1), .Y(u2_u1__abc_47660_n257) );
  OR2X2 OR2X2_3012 ( .A(u2_u1__abc_47660_n248), .B(u2_u1_b1_last_row_3_), .Y(u2_u1__abc_47660_n259) );
  OR2X2 OR2X2_3013 ( .A(u2_u1__abc_47660_n250), .B(row_adr_3_bF_buf1), .Y(u2_u1__abc_47660_n260) );
  OR2X2 OR2X2_3014 ( .A(u2_u1__abc_47660_n248), .B(u2_u1_b1_last_row_4_), .Y(u2_u1__abc_47660_n262) );
  OR2X2 OR2X2_3015 ( .A(u2_u1__abc_47660_n250), .B(row_adr_4_bF_buf1), .Y(u2_u1__abc_47660_n263) );
  OR2X2 OR2X2_3016 ( .A(u2_u1__abc_47660_n248), .B(u2_u1_b1_last_row_5_), .Y(u2_u1__abc_47660_n265) );
  OR2X2 OR2X2_3017 ( .A(u2_u1__abc_47660_n250), .B(row_adr_5_bF_buf1), .Y(u2_u1__abc_47660_n266) );
  OR2X2 OR2X2_3018 ( .A(u2_u1__abc_47660_n248), .B(u2_u1_b1_last_row_6_), .Y(u2_u1__abc_47660_n268) );
  OR2X2 OR2X2_3019 ( .A(u2_u1__abc_47660_n250), .B(row_adr_6_bF_buf1), .Y(u2_u1__abc_47660_n269) );
  OR2X2 OR2X2_302 ( .A(u0__abc_49347_n1599), .B(u0__abc_49347_n1600), .Y(u0__abc_49347_n1601) );
  OR2X2 OR2X2_3020 ( .A(u2_u1__abc_47660_n248), .B(u2_u1_b1_last_row_7_), .Y(u2_u1__abc_47660_n271) );
  OR2X2 OR2X2_3021 ( .A(u2_u1__abc_47660_n250), .B(row_adr_7_bF_buf1), .Y(u2_u1__abc_47660_n272) );
  OR2X2 OR2X2_3022 ( .A(u2_u1__abc_47660_n248), .B(u2_u1_b1_last_row_8_), .Y(u2_u1__abc_47660_n274) );
  OR2X2 OR2X2_3023 ( .A(u2_u1__abc_47660_n250), .B(row_adr_8_bF_buf1), .Y(u2_u1__abc_47660_n275_1) );
  OR2X2 OR2X2_3024 ( .A(u2_u1__abc_47660_n248), .B(u2_u1_b1_last_row_9_), .Y(u2_u1__abc_47660_n277) );
  OR2X2 OR2X2_3025 ( .A(u2_u1__abc_47660_n250), .B(row_adr_9_bF_buf1), .Y(u2_u1__abc_47660_n278_1) );
  OR2X2 OR2X2_3026 ( .A(u2_u1__abc_47660_n248), .B(u2_u1_b1_last_row_10_), .Y(u2_u1__abc_47660_n280) );
  OR2X2 OR2X2_3027 ( .A(u2_u1__abc_47660_n250), .B(row_adr_10_bF_buf1), .Y(u2_u1__abc_47660_n281) );
  OR2X2 OR2X2_3028 ( .A(u2_u1__abc_47660_n248), .B(u2_u1_b1_last_row_11_), .Y(u2_u1__abc_47660_n283_1) );
  OR2X2 OR2X2_3029 ( .A(u2_u1__abc_47660_n250), .B(row_adr_11_bF_buf1), .Y(u2_u1__abc_47660_n284) );
  OR2X2 OR2X2_303 ( .A(u0__abc_49347_n1602), .B(u0__abc_49347_n1603), .Y(u0__abc_49347_n1604) );
  OR2X2 OR2X2_3030 ( .A(u2_u1__abc_47660_n248), .B(u2_u1_b1_last_row_12_), .Y(u2_u1__abc_47660_n286_1) );
  OR2X2 OR2X2_3031 ( .A(u2_u1__abc_47660_n250), .B(row_adr_12_bF_buf1), .Y(u2_u1__abc_47660_n287_1) );
  OR2X2 OR2X2_3032 ( .A(u2_u1__abc_47660_n290_1), .B(u2_u1_b0_last_row_0_), .Y(u2_u1__abc_47660_n291) );
  OR2X2 OR2X2_3033 ( .A(u2_u1__abc_47660_n292_1), .B(row_adr_0_bF_buf0), .Y(u2_u1__abc_47660_n293) );
  OR2X2 OR2X2_3034 ( .A(u2_u1__abc_47660_n290_1), .B(u2_u1_b0_last_row_1_), .Y(u2_u1__abc_47660_n295) );
  OR2X2 OR2X2_3035 ( .A(u2_u1__abc_47660_n292_1), .B(row_adr_1_bF_buf0), .Y(u2_u1__abc_47660_n296_1) );
  OR2X2 OR2X2_3036 ( .A(u2_u1__abc_47660_n290_1), .B(u2_u1_b0_last_row_2_), .Y(u2_u1__abc_47660_n298) );
  OR2X2 OR2X2_3037 ( .A(u2_u1__abc_47660_n292_1), .B(row_adr_2_bF_buf0), .Y(u2_u1__abc_47660_n299) );
  OR2X2 OR2X2_3038 ( .A(u2_u1__abc_47660_n290_1), .B(u2_u1_b0_last_row_3_), .Y(u2_u1__abc_47660_n301) );
  OR2X2 OR2X2_3039 ( .A(u2_u1__abc_47660_n292_1), .B(row_adr_3_bF_buf0), .Y(u2_u1__abc_47660_n302) );
  OR2X2 OR2X2_304 ( .A(u0__abc_49347_n1605_1), .B(u0__abc_49347_n1606_1), .Y(u0__abc_49347_n1607) );
  OR2X2 OR2X2_3040 ( .A(u2_u1__abc_47660_n290_1), .B(u2_u1_b0_last_row_4_), .Y(u2_u1__abc_47660_n304_1) );
  OR2X2 OR2X2_3041 ( .A(u2_u1__abc_47660_n292_1), .B(row_adr_4_bF_buf0), .Y(u2_u1__abc_47660_n305_1) );
  OR2X2 OR2X2_3042 ( .A(u2_u1__abc_47660_n290_1), .B(u2_u1_b0_last_row_5_), .Y(u2_u1__abc_47660_n307) );
  OR2X2 OR2X2_3043 ( .A(u2_u1__abc_47660_n292_1), .B(row_adr_5_bF_buf0), .Y(u2_u1__abc_47660_n308) );
  OR2X2 OR2X2_3044 ( .A(u2_u1__abc_47660_n290_1), .B(u2_u1_b0_last_row_6_), .Y(u2_u1__abc_47660_n310) );
  OR2X2 OR2X2_3045 ( .A(u2_u1__abc_47660_n292_1), .B(row_adr_6_bF_buf0), .Y(u2_u1__abc_47660_n311) );
  OR2X2 OR2X2_3046 ( .A(u2_u1__abc_47660_n290_1), .B(u2_u1_b0_last_row_7_), .Y(u2_u1__abc_47660_n313) );
  OR2X2 OR2X2_3047 ( .A(u2_u1__abc_47660_n292_1), .B(row_adr_7_bF_buf0), .Y(u2_u1__abc_47660_n314) );
  OR2X2 OR2X2_3048 ( .A(u2_u1__abc_47660_n290_1), .B(u2_u1_b0_last_row_8_), .Y(u2_u1__abc_47660_n316) );
  OR2X2 OR2X2_3049 ( .A(u2_u1__abc_47660_n292_1), .B(row_adr_8_bF_buf0), .Y(u2_u1__abc_47660_n317) );
  OR2X2 OR2X2_305 ( .A(u0__abc_49347_n1609), .B(spec_req_cs_0_bF_buf3), .Y(u0__abc_49347_n1610) );
  OR2X2 OR2X2_3050 ( .A(u2_u1__abc_47660_n290_1), .B(u2_u1_b0_last_row_9_), .Y(u2_u1__abc_47660_n319) );
  OR2X2 OR2X2_3051 ( .A(u2_u1__abc_47660_n292_1), .B(row_adr_9_bF_buf0), .Y(u2_u1__abc_47660_n320) );
  OR2X2 OR2X2_3052 ( .A(u2_u1__abc_47660_n290_1), .B(u2_u1_b0_last_row_10_), .Y(u2_u1__abc_47660_n322) );
  OR2X2 OR2X2_3053 ( .A(u2_u1__abc_47660_n292_1), .B(row_adr_10_bF_buf0), .Y(u2_u1__abc_47660_n323) );
  OR2X2 OR2X2_3054 ( .A(u2_u1__abc_47660_n290_1), .B(u2_u1_b0_last_row_11_), .Y(u2_u1__abc_47660_n325) );
  OR2X2 OR2X2_3055 ( .A(u2_u1__abc_47660_n292_1), .B(row_adr_11_bF_buf0), .Y(u2_u1__abc_47660_n326) );
  OR2X2 OR2X2_3056 ( .A(u2_u1__abc_47660_n290_1), .B(u2_u1_b0_last_row_12_), .Y(u2_u1__abc_47660_n328) );
  OR2X2 OR2X2_3057 ( .A(u2_u1__abc_47660_n292_1), .B(row_adr_12_bF_buf0), .Y(u2_u1__abc_47660_n329) );
  OR2X2 OR2X2_3058 ( .A(u2_u1__abc_47660_n331), .B(row_adr_12_bF_buf6), .Y(u2_u1__abc_47660_n332) );
  OR2X2 OR2X2_3059 ( .A(u2_u1__abc_47660_n333), .B(row_adr_11_bF_buf6), .Y(u2_u1__abc_47660_n334) );
  OR2X2 OR2X2_306 ( .A(u0__abc_49347_n1608), .B(u0__abc_49347_n1610), .Y(u0__abc_49347_n1611) );
  OR2X2 OR2X2_3060 ( .A(u2_u1__abc_47660_n199), .B(u2_u1_b0_last_row_12_), .Y(u2_u1__abc_47660_n335) );
  OR2X2 OR2X2_3061 ( .A(u2_u1__abc_47660_n194), .B(u2_u1_b0_last_row_11_), .Y(u2_u1__abc_47660_n338) );
  OR2X2 OR2X2_3062 ( .A(u2_u1__abc_47660_n339), .B(row_adr_9_bF_buf6), .Y(u2_u1__abc_47660_n340) );
  OR2X2 OR2X2_3063 ( .A(u2_u1__abc_47660_n184), .B(u2_u1_b0_last_row_9_), .Y(u2_u1__abc_47660_n342) );
  OR2X2 OR2X2_3064 ( .A(u2_u1__abc_47660_n343), .B(row_adr_7_bF_buf6), .Y(u2_u1__abc_47660_n344) );
  OR2X2 OR2X2_3065 ( .A(u2_u1__abc_47660_n164), .B(u2_u1_b0_last_row_5_), .Y(u2_u1__abc_47660_n348) );
  OR2X2 OR2X2_3066 ( .A(u2_u1__abc_47660_n159), .B(u2_u1_b0_last_row_4_), .Y(u2_u1__abc_47660_n350) );
  OR2X2 OR2X2_3067 ( .A(u2_u1__abc_47660_n351), .B(row_adr_4_bF_buf6), .Y(u2_u1__abc_47660_n352) );
  OR2X2 OR2X2_3068 ( .A(u2_u1__abc_47660_n355), .B(row_adr_0_bF_buf6), .Y(u2_u1__abc_47660_n356) );
  OR2X2 OR2X2_3069 ( .A(u2_u1__abc_47660_n139), .B(u2_u1_b0_last_row_0_), .Y(u2_u1__abc_47660_n357) );
  OR2X2 OR2X2_307 ( .A(u0__abc_49347_n1203_bF_buf0), .B(u0_tms0_17_), .Y(u0__abc_49347_n1612) );
  OR2X2 OR2X2_3070 ( .A(u2_u1__abc_47660_n144), .B(u2_u1_b0_last_row_1_), .Y(u2_u1__abc_47660_n359) );
  OR2X2 OR2X2_3071 ( .A(u2_u1__abc_47660_n360), .B(row_adr_5_bF_buf6), .Y(u2_u1__abc_47660_n361) );
  OR2X2 OR2X2_3072 ( .A(u2_u1__abc_47660_n366), .B(row_adr_10_bF_buf6), .Y(u2_u1__abc_47660_n367) );
  OR2X2 OR2X2_3073 ( .A(u2_u1__abc_47660_n189), .B(u2_u1_b0_last_row_10_), .Y(u2_u1__abc_47660_n368) );
  OR2X2 OR2X2_3074 ( .A(u2_u1__abc_47660_n372), .B(u2_u1__abc_47660_n370), .Y(u2_u1__abc_47660_n373) );
  OR2X2 OR2X2_3075 ( .A(u2_u1__abc_47660_n154), .B(u2_u1_b0_last_row_3_), .Y(u2_u1__abc_47660_n375) );
  OR2X2 OR2X2_3076 ( .A(u2_u1__abc_47660_n376), .B(row_adr_2_bF_buf6), .Y(u2_u1__abc_47660_n377) );
  OR2X2 OR2X2_3077 ( .A(u2_u1__abc_47660_n379), .B(row_adr_1_bF_buf6), .Y(u2_u1__abc_47660_n380) );
  OR2X2 OR2X2_3078 ( .A(u2_u1__abc_47660_n149), .B(u2_u1_b0_last_row_2_), .Y(u2_u1__abc_47660_n381) );
  OR2X2 OR2X2_3079 ( .A(u2_u1__abc_47660_n384), .B(row_adr_3_bF_buf6), .Y(u2_u1__abc_47660_n385) );
  OR2X2 OR2X2_308 ( .A(u0__abc_49347_n1614_1), .B(u0__abc_49347_n1592), .Y(u0_sp_tms_17__FF_INPUT) );
  OR2X2 OR2X2_3080 ( .A(u2_u1__abc_47660_n174), .B(u2_u1_b0_last_row_7_), .Y(u2_u1__abc_47660_n386) );
  OR2X2 OR2X2_3081 ( .A(u2_u1__abc_47660_n390), .B(u2_u1__abc_47660_n388), .Y(u2_u1__abc_47660_n391) );
  OR2X2 OR2X2_3082 ( .A(u2_u1__abc_47660_n396), .B(row_adr_12_bF_buf5), .Y(u2_u1__abc_47660_n397) );
  OR2X2 OR2X2_3083 ( .A(u2_u1__abc_47660_n398), .B(row_adr_11_bF_buf5), .Y(u2_u1__abc_47660_n399) );
  OR2X2 OR2X2_3084 ( .A(u2_u1__abc_47660_n199), .B(u2_u1_b2_last_row_12_), .Y(u2_u1__abc_47660_n400) );
  OR2X2 OR2X2_3085 ( .A(u2_u1__abc_47660_n194), .B(u2_u1_b2_last_row_11_), .Y(u2_u1__abc_47660_n403) );
  OR2X2 OR2X2_3086 ( .A(u2_u1__abc_47660_n404), .B(row_adr_9_bF_buf5), .Y(u2_u1__abc_47660_n405) );
  OR2X2 OR2X2_3087 ( .A(u2_u1__abc_47660_n184), .B(u2_u1_b2_last_row_9_), .Y(u2_u1__abc_47660_n407) );
  OR2X2 OR2X2_3088 ( .A(u2_u1__abc_47660_n408), .B(row_adr_7_bF_buf5), .Y(u2_u1__abc_47660_n409) );
  OR2X2 OR2X2_3089 ( .A(u2_u1__abc_47660_n164), .B(u2_u1_b2_last_row_5_), .Y(u2_u1__abc_47660_n413) );
  OR2X2 OR2X2_309 ( .A(u0__abc_49347_n1183_1_bF_buf5), .B(1'b0), .Y(u0__abc_49347_n1618) );
  OR2X2 OR2X2_3090 ( .A(u2_u1__abc_47660_n159), .B(u2_u1_b2_last_row_4_), .Y(u2_u1__abc_47660_n415) );
  OR2X2 OR2X2_3091 ( .A(u2_u1__abc_47660_n416), .B(row_adr_4_bF_buf5), .Y(u2_u1__abc_47660_n417) );
  OR2X2 OR2X2_3092 ( .A(u2_u1__abc_47660_n420), .B(row_adr_0_bF_buf5), .Y(u2_u1__abc_47660_n421) );
  OR2X2 OR2X2_3093 ( .A(u2_u1__abc_47660_n139), .B(u2_u1_b2_last_row_0_), .Y(u2_u1__abc_47660_n422) );
  OR2X2 OR2X2_3094 ( .A(u2_u1__abc_47660_n144), .B(u2_u1_b2_last_row_1_), .Y(u2_u1__abc_47660_n424) );
  OR2X2 OR2X2_3095 ( .A(u2_u1__abc_47660_n425), .B(row_adr_5_bF_buf5), .Y(u2_u1__abc_47660_n426) );
  OR2X2 OR2X2_3096 ( .A(u2_u1__abc_47660_n431), .B(row_adr_10_bF_buf5), .Y(u2_u1__abc_47660_n432) );
  OR2X2 OR2X2_3097 ( .A(u2_u1__abc_47660_n189), .B(u2_u1_b2_last_row_10_), .Y(u2_u1__abc_47660_n433) );
  OR2X2 OR2X2_3098 ( .A(u2_u1__abc_47660_n437), .B(u2_u1__abc_47660_n435), .Y(u2_u1__abc_47660_n438) );
  OR2X2 OR2X2_3099 ( .A(u2_u1__abc_47660_n154), .B(u2_u1_b2_last_row_3_), .Y(u2_u1__abc_47660_n440) );
  OR2X2 OR2X2_31 ( .A(_abc_55805_n240_bF_buf4), .B(spec_req_cs_7_), .Y(_abc_55805_n284) );
  OR2X2 OR2X2_310 ( .A(spec_req_cs_6_bF_buf2), .B(1'b0), .Y(u0__abc_49347_n1619) );
  OR2X2 OR2X2_3100 ( .A(u2_u1__abc_47660_n441), .B(row_adr_2_bF_buf5), .Y(u2_u1__abc_47660_n442) );
  OR2X2 OR2X2_3101 ( .A(u2_u1__abc_47660_n444), .B(row_adr_1_bF_buf5), .Y(u2_u1__abc_47660_n445) );
  OR2X2 OR2X2_3102 ( .A(u2_u1__abc_47660_n149), .B(u2_u1_b2_last_row_2_), .Y(u2_u1__abc_47660_n446) );
  OR2X2 OR2X2_3103 ( .A(u2_u1__abc_47660_n449), .B(row_adr_3_bF_buf5), .Y(u2_u1__abc_47660_n450) );
  OR2X2 OR2X2_3104 ( .A(u2_u1__abc_47660_n174), .B(u2_u1_b2_last_row_7_), .Y(u2_u1__abc_47660_n451) );
  OR2X2 OR2X2_3105 ( .A(u2_u1__abc_47660_n455), .B(u2_u1__abc_47660_n453), .Y(u2_u1__abc_47660_n456) );
  OR2X2 OR2X2_3106 ( .A(u2_u1__abc_47660_n395), .B(u2_u1__abc_47660_n460), .Y(u2_u1__abc_47660_n461) );
  OR2X2 OR2X2_3107 ( .A(u2_u1__abc_47660_n462), .B(row_adr_12_bF_buf4), .Y(u2_u1__abc_47660_n463) );
  OR2X2 OR2X2_3108 ( .A(u2_u1__abc_47660_n464), .B(row_adr_11_bF_buf4), .Y(u2_u1__abc_47660_n465) );
  OR2X2 OR2X2_3109 ( .A(u2_u1__abc_47660_n199), .B(u2_u1_b1_last_row_12_), .Y(u2_u1__abc_47660_n466) );
  OR2X2 OR2X2_311 ( .A(u0__abc_49347_n1621), .B(u0__abc_49347_n1617), .Y(u0__abc_49347_n1622) );
  OR2X2 OR2X2_3110 ( .A(u2_u1__abc_47660_n194), .B(u2_u1_b1_last_row_11_), .Y(u2_u1__abc_47660_n469) );
  OR2X2 OR2X2_3111 ( .A(u2_u1__abc_47660_n470), .B(row_adr_9_bF_buf4), .Y(u2_u1__abc_47660_n471) );
  OR2X2 OR2X2_3112 ( .A(u2_u1__abc_47660_n184), .B(u2_u1_b1_last_row_9_), .Y(u2_u1__abc_47660_n473) );
  OR2X2 OR2X2_3113 ( .A(u2_u1__abc_47660_n474), .B(row_adr_7_bF_buf4), .Y(u2_u1__abc_47660_n475) );
  OR2X2 OR2X2_3114 ( .A(u2_u1__abc_47660_n164), .B(u2_u1_b1_last_row_5_), .Y(u2_u1__abc_47660_n479) );
  OR2X2 OR2X2_3115 ( .A(u2_u1__abc_47660_n159), .B(u2_u1_b1_last_row_4_), .Y(u2_u1__abc_47660_n481) );
  OR2X2 OR2X2_3116 ( .A(u2_u1__abc_47660_n482), .B(row_adr_4_bF_buf4), .Y(u2_u1__abc_47660_n483) );
  OR2X2 OR2X2_3117 ( .A(u2_u1__abc_47660_n486), .B(row_adr_0_bF_buf4), .Y(u2_u1__abc_47660_n487) );
  OR2X2 OR2X2_3118 ( .A(u2_u1__abc_47660_n139), .B(u2_u1_b1_last_row_0_), .Y(u2_u1__abc_47660_n488) );
  OR2X2 OR2X2_3119 ( .A(u2_u1__abc_47660_n144), .B(u2_u1_b1_last_row_1_), .Y(u2_u1__abc_47660_n490) );
  OR2X2 OR2X2_312 ( .A(u0__abc_49347_n1623_1), .B(u0__abc_49347_n1624_1), .Y(u0__abc_49347_n1625) );
  OR2X2 OR2X2_3120 ( .A(u2_u1__abc_47660_n491), .B(row_adr_5_bF_buf4), .Y(u2_u1__abc_47660_n492) );
  OR2X2 OR2X2_3121 ( .A(u2_u1__abc_47660_n497), .B(row_adr_10_bF_buf4), .Y(u2_u1__abc_47660_n498) );
  OR2X2 OR2X2_3122 ( .A(u2_u1__abc_47660_n189), .B(u2_u1_b1_last_row_10_), .Y(u2_u1__abc_47660_n499) );
  OR2X2 OR2X2_3123 ( .A(u2_u1__abc_47660_n503), .B(u2_u1__abc_47660_n501), .Y(u2_u1__abc_47660_n504) );
  OR2X2 OR2X2_3124 ( .A(u2_u1__abc_47660_n154), .B(u2_u1_b1_last_row_3_), .Y(u2_u1__abc_47660_n506) );
  OR2X2 OR2X2_3125 ( .A(u2_u1__abc_47660_n507), .B(row_adr_2_bF_buf4), .Y(u2_u1__abc_47660_n508) );
  OR2X2 OR2X2_3126 ( .A(u2_u1__abc_47660_n510), .B(row_adr_1_bF_buf4), .Y(u2_u1__abc_47660_n511) );
  OR2X2 OR2X2_3127 ( .A(u2_u1__abc_47660_n149), .B(u2_u1_b1_last_row_2_), .Y(u2_u1__abc_47660_n512) );
  OR2X2 OR2X2_3128 ( .A(u2_u1__abc_47660_n515), .B(row_adr_3_bF_buf4), .Y(u2_u1__abc_47660_n516) );
  OR2X2 OR2X2_3129 ( .A(u2_u1__abc_47660_n174), .B(u2_u1_b1_last_row_7_), .Y(u2_u1__abc_47660_n517) );
  OR2X2 OR2X2_313 ( .A(u0__abc_49347_n1626), .B(u0__abc_49347_n1627), .Y(u0__abc_49347_n1628) );
  OR2X2 OR2X2_3130 ( .A(u2_u1__abc_47660_n521), .B(u2_u1__abc_47660_n519), .Y(u2_u1__abc_47660_n522) );
  OR2X2 OR2X2_3131 ( .A(u2_u1__abc_47660_n527), .B(row_adr_9_bF_buf3), .Y(u2_u1__abc_47660_n528) );
  OR2X2 OR2X2_3132 ( .A(u2_u1__abc_47660_n189), .B(u2_u1_b3_last_row_10_), .Y(u2_u1__abc_47660_n529) );
  OR2X2 OR2X2_3133 ( .A(u2_u1__abc_47660_n184), .B(u2_u1_b3_last_row_9_), .Y(u2_u1__abc_47660_n530) );
  OR2X2 OR2X2_3134 ( .A(u2_u1__abc_47660_n194), .B(u2_u1_b3_last_row_11_), .Y(u2_u1__abc_47660_n533) );
  OR2X2 OR2X2_3135 ( .A(u2_u1__abc_47660_n534), .B(row_adr_11_bF_buf3), .Y(u2_u1__abc_47660_n535) );
  OR2X2 OR2X2_3136 ( .A(u2_u1__abc_47660_n199), .B(u2_u1_b3_last_row_12_), .Y(u2_u1__abc_47660_n537) );
  OR2X2 OR2X2_3137 ( .A(u2_u1__abc_47660_n538), .B(row_adr_8_bF_buf3), .Y(u2_u1__abc_47660_n539) );
  OR2X2 OR2X2_3138 ( .A(u2_u1__abc_47660_n159), .B(u2_u1_b3_last_row_4_), .Y(u2_u1__abc_47660_n543) );
  OR2X2 OR2X2_3139 ( .A(u2_u1__abc_47660_n544), .B(row_adr_4_bF_buf3), .Y(u2_u1__abc_47660_n545) );
  OR2X2 OR2X2_314 ( .A(u0__abc_49347_n1629), .B(u0__abc_49347_n1630), .Y(u0__abc_49347_n1631) );
  OR2X2 OR2X2_3140 ( .A(u2_u1__abc_47660_n547), .B(row_adr_3_bF_buf3), .Y(u2_u1__abc_47660_n548) );
  OR2X2 OR2X2_3141 ( .A(u2_u1__abc_47660_n551), .B(row_adr_0_bF_buf3), .Y(u2_u1__abc_47660_n552) );
  OR2X2 OR2X2_3142 ( .A(u2_u1__abc_47660_n139), .B(u2_u1_b3_last_row_0_), .Y(u2_u1__abc_47660_n553) );
  OR2X2 OR2X2_3143 ( .A(u2_u1__abc_47660_n555), .B(row_adr_2_bF_buf3), .Y(u2_u1__abc_47660_n556) );
  OR2X2 OR2X2_3144 ( .A(u2_u1__abc_47660_n149), .B(u2_u1_b3_last_row_2_), .Y(u2_u1__abc_47660_n557) );
  OR2X2 OR2X2_3145 ( .A(u2_u1__abc_47660_n174), .B(u2_u1_b3_last_row_7_), .Y(u2_u1__abc_47660_n562) );
  OR2X2 OR2X2_3146 ( .A(u2_u1__abc_47660_n563), .B(row_adr_7_bF_buf3), .Y(u2_u1__abc_47660_n564) );
  OR2X2 OR2X2_3147 ( .A(u2_u1__abc_47660_n566), .B(row_adr_10_bF_buf3), .Y(u2_u1__abc_47660_n567) );
  OR2X2 OR2X2_3148 ( .A(u2_u1__abc_47660_n179), .B(u2_u1_b3_last_row_8_), .Y(u2_u1__abc_47660_n568) );
  OR2X2 OR2X2_3149 ( .A(u2_u1__abc_47660_n169), .B(u2_u1_b3_last_row_6_), .Y(u2_u1__abc_47660_n571) );
  OR2X2 OR2X2_315 ( .A(u0__abc_49347_n1633_1), .B(spec_req_cs_0_bF_buf2), .Y(u0__abc_49347_n1634) );
  OR2X2 OR2X2_3150 ( .A(u2_u1__abc_47660_n572), .B(row_adr_6_bF_buf3), .Y(u2_u1__abc_47660_n573) );
  OR2X2 OR2X2_3151 ( .A(u2_u1__abc_47660_n575), .B(row_adr_5_bF_buf3), .Y(u2_u1__abc_47660_n576) );
  OR2X2 OR2X2_3152 ( .A(u2_u1__abc_47660_n154), .B(u2_u1_b3_last_row_3_), .Y(u2_u1__abc_47660_n577) );
  OR2X2 OR2X2_3153 ( .A(u2_u1__abc_47660_n164), .B(u2_u1_b3_last_row_5_), .Y(u2_u1__abc_47660_n580) );
  OR2X2 OR2X2_3154 ( .A(u2_u1__abc_47660_n581), .B(row_adr_1_bF_buf3), .Y(u2_u1__abc_47660_n582) );
  OR2X2 OR2X2_3155 ( .A(u2_u1__abc_47660_n144), .B(u2_u1_b3_last_row_1_), .Y(u2_u1__abc_47660_n584) );
  OR2X2 OR2X2_3156 ( .A(u2_u1__abc_47660_n585), .B(row_adr_12_bF_buf3), .Y(u2_u1__abc_47660_n586) );
  OR2X2 OR2X2_3157 ( .A(u2_u1__abc_47660_n526), .B(u2_u1__abc_47660_n591), .Y(u2_u1__abc_47660_n592) );
  OR2X2 OR2X2_3158 ( .A(u2_u1__abc_47660_n461), .B(u2_u1__abc_47660_n592), .Y(u2_row_same_1) );
  OR2X2 OR2X2_3159 ( .A(u2_u1__abc_47660_n594), .B(u2_u1__abc_47660_n595), .Y(u2_u1__abc_47660_n596) );
  OR2X2 OR2X2_316 ( .A(u0__abc_49347_n1632_1), .B(u0__abc_49347_n1634), .Y(u0__abc_49347_n1635) );
  OR2X2 OR2X2_3160 ( .A(u2_u1__abc_47660_n598), .B(u2_u1__abc_47660_n597), .Y(u2_u1__abc_47660_n599) );
  OR2X2 OR2X2_3161 ( .A(u2_u1__abc_47660_n596), .B(u2_u1__abc_47660_n599), .Y(u2_bank_open_1) );
  OR2X2 OR2X2_3162 ( .A(u2_u1__abc_47660_n608), .B(u2_u1__abc_47660_n137_bF_buf3), .Y(u2_u1_bank3_open_FF_INPUT) );
  OR2X2 OR2X2_3163 ( .A(u2_u1__abc_47660_n611), .B(u2_u1__abc_47660_n610), .Y(u2_u1__abc_47660_n612) );
  OR2X2 OR2X2_3164 ( .A(u2_u1__abc_47660_n614), .B(u2_u1__abc_47660_n205), .Y(u2_u1_bank2_open_FF_INPUT) );
  OR2X2 OR2X2_3165 ( .A(u2_u1__abc_47660_n616), .B(u2_u1__abc_47660_n610), .Y(u2_u1__abc_47660_n617) );
  OR2X2 OR2X2_3166 ( .A(u2_u1__abc_47660_n619), .B(u2_u1__abc_47660_n248), .Y(u2_u1_bank1_open_FF_INPUT) );
  OR2X2 OR2X2_3167 ( .A(u2_u1__abc_47660_n621), .B(u2_u1__abc_47660_n610), .Y(u2_u1__abc_47660_n622) );
  OR2X2 OR2X2_3168 ( .A(u2_u1__abc_47660_n624), .B(u2_u1__abc_47660_n290_1), .Y(u2_u1_bank0_open_FF_INPUT) );
  OR2X2 OR2X2_3169 ( .A(u2_u2__abc_47660_n137_bF_buf4), .B(u2_u2_b3_last_row_0_), .Y(u2_u2__abc_47660_n138) );
  OR2X2 OR2X2_317 ( .A(u0__abc_49347_n1203_bF_buf5), .B(u0_tms0_18_), .Y(u0__abc_49347_n1636) );
  OR2X2 OR2X2_3170 ( .A(u2_u2__abc_47660_n137_bF_buf2), .B(u2_u2_b3_last_row_1_), .Y(u2_u2__abc_47660_n143) );
  OR2X2 OR2X2_3171 ( .A(u2_u2__abc_47660_n137_bF_buf0), .B(u2_u2_b3_last_row_2_), .Y(u2_u2__abc_47660_n148) );
  OR2X2 OR2X2_3172 ( .A(u2_u2__abc_47660_n137_bF_buf3), .B(u2_u2_b3_last_row_3_), .Y(u2_u2__abc_47660_n153) );
  OR2X2 OR2X2_3173 ( .A(u2_u2__abc_47660_n137_bF_buf1), .B(u2_u2_b3_last_row_4_), .Y(u2_u2__abc_47660_n158) );
  OR2X2 OR2X2_3174 ( .A(u2_u2__abc_47660_n137_bF_buf4), .B(u2_u2_b3_last_row_5_), .Y(u2_u2__abc_47660_n163) );
  OR2X2 OR2X2_3175 ( .A(u2_u2__abc_47660_n137_bF_buf2), .B(u2_u2_b3_last_row_6_), .Y(u2_u2__abc_47660_n168) );
  OR2X2 OR2X2_3176 ( .A(u2_u2__abc_47660_n137_bF_buf0), .B(u2_u2_b3_last_row_7_), .Y(u2_u2__abc_47660_n173) );
  OR2X2 OR2X2_3177 ( .A(u2_u2__abc_47660_n137_bF_buf3), .B(u2_u2_b3_last_row_8_), .Y(u2_u2__abc_47660_n178) );
  OR2X2 OR2X2_3178 ( .A(u2_u2__abc_47660_n137_bF_buf1), .B(u2_u2_b3_last_row_9_), .Y(u2_u2__abc_47660_n183) );
  OR2X2 OR2X2_3179 ( .A(u2_u2__abc_47660_n137_bF_buf4), .B(u2_u2_b3_last_row_10_), .Y(u2_u2__abc_47660_n188) );
  OR2X2 OR2X2_318 ( .A(u0__abc_49347_n1638), .B(u0__abc_49347_n1616), .Y(u0_sp_tms_18__FF_INPUT) );
  OR2X2 OR2X2_3180 ( .A(u2_u2__abc_47660_n137_bF_buf2), .B(u2_u2_b3_last_row_11_), .Y(u2_u2__abc_47660_n193) );
  OR2X2 OR2X2_3181 ( .A(u2_u2__abc_47660_n137_bF_buf0), .B(u2_u2_b3_last_row_12_), .Y(u2_u2__abc_47660_n198) );
  OR2X2 OR2X2_3182 ( .A(u2_u2__abc_47660_n205), .B(u2_u2_b2_last_row_0_), .Y(u2_u2__abc_47660_n206) );
  OR2X2 OR2X2_3183 ( .A(u2_u2__abc_47660_n207), .B(row_adr_0_bF_buf1), .Y(u2_u2__abc_47660_n208) );
  OR2X2 OR2X2_3184 ( .A(u2_u2__abc_47660_n205), .B(u2_u2_b2_last_row_1_), .Y(u2_u2__abc_47660_n210) );
  OR2X2 OR2X2_3185 ( .A(u2_u2__abc_47660_n207), .B(row_adr_1_bF_buf1), .Y(u2_u2__abc_47660_n211) );
  OR2X2 OR2X2_3186 ( .A(u2_u2__abc_47660_n205), .B(u2_u2_b2_last_row_2_), .Y(u2_u2__abc_47660_n213) );
  OR2X2 OR2X2_3187 ( .A(u2_u2__abc_47660_n207), .B(row_adr_2_bF_buf1), .Y(u2_u2__abc_47660_n214) );
  OR2X2 OR2X2_3188 ( .A(u2_u2__abc_47660_n205), .B(u2_u2_b2_last_row_3_), .Y(u2_u2__abc_47660_n216) );
  OR2X2 OR2X2_3189 ( .A(u2_u2__abc_47660_n207), .B(row_adr_3_bF_buf1), .Y(u2_u2__abc_47660_n217) );
  OR2X2 OR2X2_319 ( .A(u0__abc_49347_n1183_1_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n1642_1) );
  OR2X2 OR2X2_3190 ( .A(u2_u2__abc_47660_n205), .B(u2_u2_b2_last_row_4_), .Y(u2_u2__abc_47660_n219) );
  OR2X2 OR2X2_3191 ( .A(u2_u2__abc_47660_n207), .B(row_adr_4_bF_buf1), .Y(u2_u2__abc_47660_n220) );
  OR2X2 OR2X2_3192 ( .A(u2_u2__abc_47660_n205), .B(u2_u2_b2_last_row_5_), .Y(u2_u2__abc_47660_n222) );
  OR2X2 OR2X2_3193 ( .A(u2_u2__abc_47660_n207), .B(row_adr_5_bF_buf1), .Y(u2_u2__abc_47660_n223) );
  OR2X2 OR2X2_3194 ( .A(u2_u2__abc_47660_n205), .B(u2_u2_b2_last_row_6_), .Y(u2_u2__abc_47660_n225) );
  OR2X2 OR2X2_3195 ( .A(u2_u2__abc_47660_n207), .B(row_adr_6_bF_buf1), .Y(u2_u2__abc_47660_n226) );
  OR2X2 OR2X2_3196 ( .A(u2_u2__abc_47660_n205), .B(u2_u2_b2_last_row_7_), .Y(u2_u2__abc_47660_n228) );
  OR2X2 OR2X2_3197 ( .A(u2_u2__abc_47660_n207), .B(row_adr_7_bF_buf1), .Y(u2_u2__abc_47660_n229) );
  OR2X2 OR2X2_3198 ( .A(u2_u2__abc_47660_n205), .B(u2_u2_b2_last_row_8_), .Y(u2_u2__abc_47660_n231) );
  OR2X2 OR2X2_3199 ( .A(u2_u2__abc_47660_n207), .B(row_adr_8_bF_buf1), .Y(u2_u2__abc_47660_n232) );
  OR2X2 OR2X2_32 ( .A(lmr_sel_bF_buf6), .B(cs_7_), .Y(_abc_55805_n285) );
  OR2X2 OR2X2_320 ( .A(spec_req_cs_6_bF_buf1), .B(1'b0), .Y(u0__abc_49347_n1643) );
  OR2X2 OR2X2_3200 ( .A(u2_u2__abc_47660_n205), .B(u2_u2_b2_last_row_9_), .Y(u2_u2__abc_47660_n234) );
  OR2X2 OR2X2_3201 ( .A(u2_u2__abc_47660_n207), .B(row_adr_9_bF_buf1), .Y(u2_u2__abc_47660_n235) );
  OR2X2 OR2X2_3202 ( .A(u2_u2__abc_47660_n205), .B(u2_u2_b2_last_row_10_), .Y(u2_u2__abc_47660_n237) );
  OR2X2 OR2X2_3203 ( .A(u2_u2__abc_47660_n207), .B(row_adr_10_bF_buf1), .Y(u2_u2__abc_47660_n238) );
  OR2X2 OR2X2_3204 ( .A(u2_u2__abc_47660_n205), .B(u2_u2_b2_last_row_11_), .Y(u2_u2__abc_47660_n240) );
  OR2X2 OR2X2_3205 ( .A(u2_u2__abc_47660_n207), .B(row_adr_11_bF_buf1), .Y(u2_u2__abc_47660_n241) );
  OR2X2 OR2X2_3206 ( .A(u2_u2__abc_47660_n205), .B(u2_u2_b2_last_row_12_), .Y(u2_u2__abc_47660_n243) );
  OR2X2 OR2X2_3207 ( .A(u2_u2__abc_47660_n207), .B(row_adr_12_bF_buf1), .Y(u2_u2__abc_47660_n244) );
  OR2X2 OR2X2_3208 ( .A(u2_u2__abc_47660_n248), .B(u2_u2_b1_last_row_0_), .Y(u2_u2__abc_47660_n249) );
  OR2X2 OR2X2_3209 ( .A(u2_u2__abc_47660_n250), .B(row_adr_0_bF_buf0), .Y(u2_u2__abc_47660_n251) );
  OR2X2 OR2X2_321 ( .A(u0__abc_49347_n1645), .B(u0__abc_49347_n1641_1), .Y(u0__abc_49347_n1646) );
  OR2X2 OR2X2_3210 ( .A(u2_u2__abc_47660_n248), .B(u2_u2_b1_last_row_1_), .Y(u2_u2__abc_47660_n253) );
  OR2X2 OR2X2_3211 ( .A(u2_u2__abc_47660_n250), .B(row_adr_1_bF_buf0), .Y(u2_u2__abc_47660_n254) );
  OR2X2 OR2X2_3212 ( .A(u2_u2__abc_47660_n248), .B(u2_u2_b1_last_row_2_), .Y(u2_u2__abc_47660_n256) );
  OR2X2 OR2X2_3213 ( .A(u2_u2__abc_47660_n250), .B(row_adr_2_bF_buf0), .Y(u2_u2__abc_47660_n257) );
  OR2X2 OR2X2_3214 ( .A(u2_u2__abc_47660_n248), .B(u2_u2_b1_last_row_3_), .Y(u2_u2__abc_47660_n259) );
  OR2X2 OR2X2_3215 ( .A(u2_u2__abc_47660_n250), .B(row_adr_3_bF_buf0), .Y(u2_u2__abc_47660_n260) );
  OR2X2 OR2X2_3216 ( .A(u2_u2__abc_47660_n248), .B(u2_u2_b1_last_row_4_), .Y(u2_u2__abc_47660_n262) );
  OR2X2 OR2X2_3217 ( .A(u2_u2__abc_47660_n250), .B(row_adr_4_bF_buf0), .Y(u2_u2__abc_47660_n263) );
  OR2X2 OR2X2_3218 ( .A(u2_u2__abc_47660_n248), .B(u2_u2_b1_last_row_5_), .Y(u2_u2__abc_47660_n265) );
  OR2X2 OR2X2_3219 ( .A(u2_u2__abc_47660_n250), .B(row_adr_5_bF_buf0), .Y(u2_u2__abc_47660_n266) );
  OR2X2 OR2X2_322 ( .A(u0__abc_49347_n1647), .B(u0__abc_49347_n1648), .Y(u0__abc_49347_n1649) );
  OR2X2 OR2X2_3220 ( .A(u2_u2__abc_47660_n248), .B(u2_u2_b1_last_row_6_), .Y(u2_u2__abc_47660_n268) );
  OR2X2 OR2X2_3221 ( .A(u2_u2__abc_47660_n250), .B(row_adr_6_bF_buf0), .Y(u2_u2__abc_47660_n269) );
  OR2X2 OR2X2_3222 ( .A(u2_u2__abc_47660_n248), .B(u2_u2_b1_last_row_7_), .Y(u2_u2__abc_47660_n271) );
  OR2X2 OR2X2_3223 ( .A(u2_u2__abc_47660_n250), .B(row_adr_7_bF_buf0), .Y(u2_u2__abc_47660_n272) );
  OR2X2 OR2X2_3224 ( .A(u2_u2__abc_47660_n248), .B(u2_u2_b1_last_row_8_), .Y(u2_u2__abc_47660_n274) );
  OR2X2 OR2X2_3225 ( .A(u2_u2__abc_47660_n250), .B(row_adr_8_bF_buf0), .Y(u2_u2__abc_47660_n275_1) );
  OR2X2 OR2X2_3226 ( .A(u2_u2__abc_47660_n248), .B(u2_u2_b1_last_row_9_), .Y(u2_u2__abc_47660_n277) );
  OR2X2 OR2X2_3227 ( .A(u2_u2__abc_47660_n250), .B(row_adr_9_bF_buf0), .Y(u2_u2__abc_47660_n278_1) );
  OR2X2 OR2X2_3228 ( .A(u2_u2__abc_47660_n248), .B(u2_u2_b1_last_row_10_), .Y(u2_u2__abc_47660_n280) );
  OR2X2 OR2X2_3229 ( .A(u2_u2__abc_47660_n250), .B(row_adr_10_bF_buf0), .Y(u2_u2__abc_47660_n281) );
  OR2X2 OR2X2_323 ( .A(u0__abc_49347_n1650_1), .B(u0__abc_49347_n1651_1), .Y(u0__abc_49347_n1652) );
  OR2X2 OR2X2_3230 ( .A(u2_u2__abc_47660_n248), .B(u2_u2_b1_last_row_11_), .Y(u2_u2__abc_47660_n283_1) );
  OR2X2 OR2X2_3231 ( .A(u2_u2__abc_47660_n250), .B(row_adr_11_bF_buf0), .Y(u2_u2__abc_47660_n284) );
  OR2X2 OR2X2_3232 ( .A(u2_u2__abc_47660_n248), .B(u2_u2_b1_last_row_12_), .Y(u2_u2__abc_47660_n286_1) );
  OR2X2 OR2X2_3233 ( .A(u2_u2__abc_47660_n250), .B(row_adr_12_bF_buf0), .Y(u2_u2__abc_47660_n287_1) );
  OR2X2 OR2X2_3234 ( .A(u2_u2__abc_47660_n290_1), .B(u2_u2_b0_last_row_0_), .Y(u2_u2__abc_47660_n291) );
  OR2X2 OR2X2_3235 ( .A(u2_u2__abc_47660_n292_1), .B(row_adr_0_bF_buf6), .Y(u2_u2__abc_47660_n293) );
  OR2X2 OR2X2_3236 ( .A(u2_u2__abc_47660_n290_1), .B(u2_u2_b0_last_row_1_), .Y(u2_u2__abc_47660_n295) );
  OR2X2 OR2X2_3237 ( .A(u2_u2__abc_47660_n292_1), .B(row_adr_1_bF_buf6), .Y(u2_u2__abc_47660_n296_1) );
  OR2X2 OR2X2_3238 ( .A(u2_u2__abc_47660_n290_1), .B(u2_u2_b0_last_row_2_), .Y(u2_u2__abc_47660_n298) );
  OR2X2 OR2X2_3239 ( .A(u2_u2__abc_47660_n292_1), .B(row_adr_2_bF_buf6), .Y(u2_u2__abc_47660_n299) );
  OR2X2 OR2X2_324 ( .A(u0__abc_49347_n1653), .B(u0__abc_49347_n1654), .Y(u0__abc_49347_n1655) );
  OR2X2 OR2X2_3240 ( .A(u2_u2__abc_47660_n290_1), .B(u2_u2_b0_last_row_3_), .Y(u2_u2__abc_47660_n301) );
  OR2X2 OR2X2_3241 ( .A(u2_u2__abc_47660_n292_1), .B(row_adr_3_bF_buf6), .Y(u2_u2__abc_47660_n302) );
  OR2X2 OR2X2_3242 ( .A(u2_u2__abc_47660_n290_1), .B(u2_u2_b0_last_row_4_), .Y(u2_u2__abc_47660_n304_1) );
  OR2X2 OR2X2_3243 ( .A(u2_u2__abc_47660_n292_1), .B(row_adr_4_bF_buf6), .Y(u2_u2__abc_47660_n305_1) );
  OR2X2 OR2X2_3244 ( .A(u2_u2__abc_47660_n290_1), .B(u2_u2_b0_last_row_5_), .Y(u2_u2__abc_47660_n307) );
  OR2X2 OR2X2_3245 ( .A(u2_u2__abc_47660_n292_1), .B(row_adr_5_bF_buf6), .Y(u2_u2__abc_47660_n308) );
  OR2X2 OR2X2_3246 ( .A(u2_u2__abc_47660_n290_1), .B(u2_u2_b0_last_row_6_), .Y(u2_u2__abc_47660_n310) );
  OR2X2 OR2X2_3247 ( .A(u2_u2__abc_47660_n292_1), .B(row_adr_6_bF_buf6), .Y(u2_u2__abc_47660_n311) );
  OR2X2 OR2X2_3248 ( .A(u2_u2__abc_47660_n290_1), .B(u2_u2_b0_last_row_7_), .Y(u2_u2__abc_47660_n313) );
  OR2X2 OR2X2_3249 ( .A(u2_u2__abc_47660_n292_1), .B(row_adr_7_bF_buf6), .Y(u2_u2__abc_47660_n314) );
  OR2X2 OR2X2_325 ( .A(u0__abc_49347_n1657), .B(spec_req_cs_0_bF_buf1), .Y(u0__abc_49347_n1658) );
  OR2X2 OR2X2_3250 ( .A(u2_u2__abc_47660_n290_1), .B(u2_u2_b0_last_row_8_), .Y(u2_u2__abc_47660_n316) );
  OR2X2 OR2X2_3251 ( .A(u2_u2__abc_47660_n292_1), .B(row_adr_8_bF_buf6), .Y(u2_u2__abc_47660_n317) );
  OR2X2 OR2X2_3252 ( .A(u2_u2__abc_47660_n290_1), .B(u2_u2_b0_last_row_9_), .Y(u2_u2__abc_47660_n319) );
  OR2X2 OR2X2_3253 ( .A(u2_u2__abc_47660_n292_1), .B(row_adr_9_bF_buf6), .Y(u2_u2__abc_47660_n320) );
  OR2X2 OR2X2_3254 ( .A(u2_u2__abc_47660_n290_1), .B(u2_u2_b0_last_row_10_), .Y(u2_u2__abc_47660_n322) );
  OR2X2 OR2X2_3255 ( .A(u2_u2__abc_47660_n292_1), .B(row_adr_10_bF_buf6), .Y(u2_u2__abc_47660_n323) );
  OR2X2 OR2X2_3256 ( .A(u2_u2__abc_47660_n290_1), .B(u2_u2_b0_last_row_11_), .Y(u2_u2__abc_47660_n325) );
  OR2X2 OR2X2_3257 ( .A(u2_u2__abc_47660_n292_1), .B(row_adr_11_bF_buf6), .Y(u2_u2__abc_47660_n326) );
  OR2X2 OR2X2_3258 ( .A(u2_u2__abc_47660_n290_1), .B(u2_u2_b0_last_row_12_), .Y(u2_u2__abc_47660_n328) );
  OR2X2 OR2X2_3259 ( .A(u2_u2__abc_47660_n292_1), .B(row_adr_12_bF_buf6), .Y(u2_u2__abc_47660_n329) );
  OR2X2 OR2X2_326 ( .A(u0__abc_49347_n1656), .B(u0__abc_49347_n1658), .Y(u0__abc_49347_n1659_1) );
  OR2X2 OR2X2_3260 ( .A(u2_u2__abc_47660_n331), .B(row_adr_12_bF_buf5), .Y(u2_u2__abc_47660_n332) );
  OR2X2 OR2X2_3261 ( .A(u2_u2__abc_47660_n333), .B(row_adr_11_bF_buf5), .Y(u2_u2__abc_47660_n334) );
  OR2X2 OR2X2_3262 ( .A(u2_u2__abc_47660_n199), .B(u2_u2_b0_last_row_12_), .Y(u2_u2__abc_47660_n335) );
  OR2X2 OR2X2_3263 ( .A(u2_u2__abc_47660_n194), .B(u2_u2_b0_last_row_11_), .Y(u2_u2__abc_47660_n338) );
  OR2X2 OR2X2_3264 ( .A(u2_u2__abc_47660_n339), .B(row_adr_9_bF_buf5), .Y(u2_u2__abc_47660_n340) );
  OR2X2 OR2X2_3265 ( .A(u2_u2__abc_47660_n184), .B(u2_u2_b0_last_row_9_), .Y(u2_u2__abc_47660_n342) );
  OR2X2 OR2X2_3266 ( .A(u2_u2__abc_47660_n343), .B(row_adr_7_bF_buf5), .Y(u2_u2__abc_47660_n344) );
  OR2X2 OR2X2_3267 ( .A(u2_u2__abc_47660_n164), .B(u2_u2_b0_last_row_5_), .Y(u2_u2__abc_47660_n348) );
  OR2X2 OR2X2_3268 ( .A(u2_u2__abc_47660_n159), .B(u2_u2_b0_last_row_4_), .Y(u2_u2__abc_47660_n350) );
  OR2X2 OR2X2_3269 ( .A(u2_u2__abc_47660_n351), .B(row_adr_4_bF_buf5), .Y(u2_u2__abc_47660_n352) );
  OR2X2 OR2X2_327 ( .A(u0__abc_49347_n1203_bF_buf4), .B(u0_tms0_19_), .Y(u0__abc_49347_n1660_1) );
  OR2X2 OR2X2_3270 ( .A(u2_u2__abc_47660_n355), .B(row_adr_0_bF_buf5), .Y(u2_u2__abc_47660_n356) );
  OR2X2 OR2X2_3271 ( .A(u2_u2__abc_47660_n139), .B(u2_u2_b0_last_row_0_), .Y(u2_u2__abc_47660_n357) );
  OR2X2 OR2X2_3272 ( .A(u2_u2__abc_47660_n144), .B(u2_u2_b0_last_row_1_), .Y(u2_u2__abc_47660_n359) );
  OR2X2 OR2X2_3273 ( .A(u2_u2__abc_47660_n360), .B(row_adr_5_bF_buf5), .Y(u2_u2__abc_47660_n361) );
  OR2X2 OR2X2_3274 ( .A(u2_u2__abc_47660_n366), .B(row_adr_10_bF_buf5), .Y(u2_u2__abc_47660_n367) );
  OR2X2 OR2X2_3275 ( .A(u2_u2__abc_47660_n189), .B(u2_u2_b0_last_row_10_), .Y(u2_u2__abc_47660_n368) );
  OR2X2 OR2X2_3276 ( .A(u2_u2__abc_47660_n372), .B(u2_u2__abc_47660_n370), .Y(u2_u2__abc_47660_n373) );
  OR2X2 OR2X2_3277 ( .A(u2_u2__abc_47660_n154), .B(u2_u2_b0_last_row_3_), .Y(u2_u2__abc_47660_n375) );
  OR2X2 OR2X2_3278 ( .A(u2_u2__abc_47660_n376), .B(row_adr_2_bF_buf5), .Y(u2_u2__abc_47660_n377) );
  OR2X2 OR2X2_3279 ( .A(u2_u2__abc_47660_n379), .B(row_adr_1_bF_buf5), .Y(u2_u2__abc_47660_n380) );
  OR2X2 OR2X2_328 ( .A(u0__abc_49347_n1662), .B(u0__abc_49347_n1640), .Y(u0_sp_tms_19__FF_INPUT) );
  OR2X2 OR2X2_3280 ( .A(u2_u2__abc_47660_n149), .B(u2_u2_b0_last_row_2_), .Y(u2_u2__abc_47660_n381) );
  OR2X2 OR2X2_3281 ( .A(u2_u2__abc_47660_n384), .B(row_adr_3_bF_buf5), .Y(u2_u2__abc_47660_n385) );
  OR2X2 OR2X2_3282 ( .A(u2_u2__abc_47660_n174), .B(u2_u2_b0_last_row_7_), .Y(u2_u2__abc_47660_n386) );
  OR2X2 OR2X2_3283 ( .A(u2_u2__abc_47660_n390), .B(u2_u2__abc_47660_n388), .Y(u2_u2__abc_47660_n391) );
  OR2X2 OR2X2_3284 ( .A(u2_u2__abc_47660_n396), .B(row_adr_12_bF_buf4), .Y(u2_u2__abc_47660_n397) );
  OR2X2 OR2X2_3285 ( .A(u2_u2__abc_47660_n398), .B(row_adr_11_bF_buf4), .Y(u2_u2__abc_47660_n399) );
  OR2X2 OR2X2_3286 ( .A(u2_u2__abc_47660_n199), .B(u2_u2_b2_last_row_12_), .Y(u2_u2__abc_47660_n400) );
  OR2X2 OR2X2_3287 ( .A(u2_u2__abc_47660_n194), .B(u2_u2_b2_last_row_11_), .Y(u2_u2__abc_47660_n403) );
  OR2X2 OR2X2_3288 ( .A(u2_u2__abc_47660_n404), .B(row_adr_9_bF_buf4), .Y(u2_u2__abc_47660_n405) );
  OR2X2 OR2X2_3289 ( .A(u2_u2__abc_47660_n184), .B(u2_u2_b2_last_row_9_), .Y(u2_u2__abc_47660_n407) );
  OR2X2 OR2X2_329 ( .A(u0__abc_49347_n1183_1_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n1666) );
  OR2X2 OR2X2_3290 ( .A(u2_u2__abc_47660_n408), .B(row_adr_7_bF_buf4), .Y(u2_u2__abc_47660_n409) );
  OR2X2 OR2X2_3291 ( .A(u2_u2__abc_47660_n164), .B(u2_u2_b2_last_row_5_), .Y(u2_u2__abc_47660_n413) );
  OR2X2 OR2X2_3292 ( .A(u2_u2__abc_47660_n159), .B(u2_u2_b2_last_row_4_), .Y(u2_u2__abc_47660_n415) );
  OR2X2 OR2X2_3293 ( .A(u2_u2__abc_47660_n416), .B(row_adr_4_bF_buf4), .Y(u2_u2__abc_47660_n417) );
  OR2X2 OR2X2_3294 ( .A(u2_u2__abc_47660_n420), .B(row_adr_0_bF_buf4), .Y(u2_u2__abc_47660_n421) );
  OR2X2 OR2X2_3295 ( .A(u2_u2__abc_47660_n139), .B(u2_u2_b2_last_row_0_), .Y(u2_u2__abc_47660_n422) );
  OR2X2 OR2X2_3296 ( .A(u2_u2__abc_47660_n144), .B(u2_u2_b2_last_row_1_), .Y(u2_u2__abc_47660_n424) );
  OR2X2 OR2X2_3297 ( .A(u2_u2__abc_47660_n425), .B(row_adr_5_bF_buf4), .Y(u2_u2__abc_47660_n426) );
  OR2X2 OR2X2_3298 ( .A(u2_u2__abc_47660_n431), .B(row_adr_10_bF_buf4), .Y(u2_u2__abc_47660_n432) );
  OR2X2 OR2X2_3299 ( .A(u2_u2__abc_47660_n189), .B(u2_u2_b2_last_row_10_), .Y(u2_u2__abc_47660_n433) );
  OR2X2 OR2X2_33 ( .A(_abc_55805_n286), .B(_abc_55805_n237_1), .Y(_abc_55805_n287) );
  OR2X2 OR2X2_330 ( .A(spec_req_cs_6_bF_buf0), .B(1'b0), .Y(u0__abc_49347_n1667) );
  OR2X2 OR2X2_3300 ( .A(u2_u2__abc_47660_n437), .B(u2_u2__abc_47660_n435), .Y(u2_u2__abc_47660_n438) );
  OR2X2 OR2X2_3301 ( .A(u2_u2__abc_47660_n154), .B(u2_u2_b2_last_row_3_), .Y(u2_u2__abc_47660_n440) );
  OR2X2 OR2X2_3302 ( .A(u2_u2__abc_47660_n441), .B(row_adr_2_bF_buf4), .Y(u2_u2__abc_47660_n442) );
  OR2X2 OR2X2_3303 ( .A(u2_u2__abc_47660_n444), .B(row_adr_1_bF_buf4), .Y(u2_u2__abc_47660_n445) );
  OR2X2 OR2X2_3304 ( .A(u2_u2__abc_47660_n149), .B(u2_u2_b2_last_row_2_), .Y(u2_u2__abc_47660_n446) );
  OR2X2 OR2X2_3305 ( .A(u2_u2__abc_47660_n449), .B(row_adr_3_bF_buf4), .Y(u2_u2__abc_47660_n450) );
  OR2X2 OR2X2_3306 ( .A(u2_u2__abc_47660_n174), .B(u2_u2_b2_last_row_7_), .Y(u2_u2__abc_47660_n451) );
  OR2X2 OR2X2_3307 ( .A(u2_u2__abc_47660_n455), .B(u2_u2__abc_47660_n453), .Y(u2_u2__abc_47660_n456) );
  OR2X2 OR2X2_3308 ( .A(u2_u2__abc_47660_n395), .B(u2_u2__abc_47660_n460), .Y(u2_u2__abc_47660_n461) );
  OR2X2 OR2X2_3309 ( .A(u2_u2__abc_47660_n462), .B(row_adr_12_bF_buf3), .Y(u2_u2__abc_47660_n463) );
  OR2X2 OR2X2_331 ( .A(u0__abc_49347_n1669_1), .B(u0__abc_49347_n1665), .Y(u0__abc_49347_n1670) );
  OR2X2 OR2X2_3310 ( .A(u2_u2__abc_47660_n464), .B(row_adr_11_bF_buf3), .Y(u2_u2__abc_47660_n465) );
  OR2X2 OR2X2_3311 ( .A(u2_u2__abc_47660_n199), .B(u2_u2_b1_last_row_12_), .Y(u2_u2__abc_47660_n466) );
  OR2X2 OR2X2_3312 ( .A(u2_u2__abc_47660_n194), .B(u2_u2_b1_last_row_11_), .Y(u2_u2__abc_47660_n469) );
  OR2X2 OR2X2_3313 ( .A(u2_u2__abc_47660_n470), .B(row_adr_9_bF_buf3), .Y(u2_u2__abc_47660_n471) );
  OR2X2 OR2X2_3314 ( .A(u2_u2__abc_47660_n184), .B(u2_u2_b1_last_row_9_), .Y(u2_u2__abc_47660_n473) );
  OR2X2 OR2X2_3315 ( .A(u2_u2__abc_47660_n474), .B(row_adr_7_bF_buf3), .Y(u2_u2__abc_47660_n475) );
  OR2X2 OR2X2_3316 ( .A(u2_u2__abc_47660_n164), .B(u2_u2_b1_last_row_5_), .Y(u2_u2__abc_47660_n479) );
  OR2X2 OR2X2_3317 ( .A(u2_u2__abc_47660_n159), .B(u2_u2_b1_last_row_4_), .Y(u2_u2__abc_47660_n481) );
  OR2X2 OR2X2_3318 ( .A(u2_u2__abc_47660_n482), .B(row_adr_4_bF_buf3), .Y(u2_u2__abc_47660_n483) );
  OR2X2 OR2X2_3319 ( .A(u2_u2__abc_47660_n486), .B(row_adr_0_bF_buf3), .Y(u2_u2__abc_47660_n487) );
  OR2X2 OR2X2_332 ( .A(u0__abc_49347_n1671), .B(u0__abc_49347_n1672), .Y(u0__abc_49347_n1673) );
  OR2X2 OR2X2_3320 ( .A(u2_u2__abc_47660_n139), .B(u2_u2_b1_last_row_0_), .Y(u2_u2__abc_47660_n488) );
  OR2X2 OR2X2_3321 ( .A(u2_u2__abc_47660_n144), .B(u2_u2_b1_last_row_1_), .Y(u2_u2__abc_47660_n490) );
  OR2X2 OR2X2_3322 ( .A(u2_u2__abc_47660_n491), .B(row_adr_5_bF_buf3), .Y(u2_u2__abc_47660_n492) );
  OR2X2 OR2X2_3323 ( .A(u2_u2__abc_47660_n497), .B(row_adr_10_bF_buf3), .Y(u2_u2__abc_47660_n498) );
  OR2X2 OR2X2_3324 ( .A(u2_u2__abc_47660_n189), .B(u2_u2_b1_last_row_10_), .Y(u2_u2__abc_47660_n499) );
  OR2X2 OR2X2_3325 ( .A(u2_u2__abc_47660_n503), .B(u2_u2__abc_47660_n501), .Y(u2_u2__abc_47660_n504) );
  OR2X2 OR2X2_3326 ( .A(u2_u2__abc_47660_n154), .B(u2_u2_b1_last_row_3_), .Y(u2_u2__abc_47660_n506) );
  OR2X2 OR2X2_3327 ( .A(u2_u2__abc_47660_n507), .B(row_adr_2_bF_buf3), .Y(u2_u2__abc_47660_n508) );
  OR2X2 OR2X2_3328 ( .A(u2_u2__abc_47660_n510), .B(row_adr_1_bF_buf3), .Y(u2_u2__abc_47660_n511) );
  OR2X2 OR2X2_3329 ( .A(u2_u2__abc_47660_n149), .B(u2_u2_b1_last_row_2_), .Y(u2_u2__abc_47660_n512) );
  OR2X2 OR2X2_333 ( .A(u0__abc_49347_n1674), .B(u0__abc_49347_n1675), .Y(u0__abc_49347_n1676) );
  OR2X2 OR2X2_3330 ( .A(u2_u2__abc_47660_n515), .B(row_adr_3_bF_buf3), .Y(u2_u2__abc_47660_n516) );
  OR2X2 OR2X2_3331 ( .A(u2_u2__abc_47660_n174), .B(u2_u2_b1_last_row_7_), .Y(u2_u2__abc_47660_n517) );
  OR2X2 OR2X2_3332 ( .A(u2_u2__abc_47660_n521), .B(u2_u2__abc_47660_n519), .Y(u2_u2__abc_47660_n522) );
  OR2X2 OR2X2_3333 ( .A(u2_u2__abc_47660_n527), .B(row_adr_9_bF_buf2), .Y(u2_u2__abc_47660_n528) );
  OR2X2 OR2X2_3334 ( .A(u2_u2__abc_47660_n189), .B(u2_u2_b3_last_row_10_), .Y(u2_u2__abc_47660_n529) );
  OR2X2 OR2X2_3335 ( .A(u2_u2__abc_47660_n184), .B(u2_u2_b3_last_row_9_), .Y(u2_u2__abc_47660_n530) );
  OR2X2 OR2X2_3336 ( .A(u2_u2__abc_47660_n194), .B(u2_u2_b3_last_row_11_), .Y(u2_u2__abc_47660_n533) );
  OR2X2 OR2X2_3337 ( .A(u2_u2__abc_47660_n534), .B(row_adr_11_bF_buf2), .Y(u2_u2__abc_47660_n535) );
  OR2X2 OR2X2_3338 ( .A(u2_u2__abc_47660_n199), .B(u2_u2_b3_last_row_12_), .Y(u2_u2__abc_47660_n537) );
  OR2X2 OR2X2_3339 ( .A(u2_u2__abc_47660_n538), .B(row_adr_8_bF_buf2), .Y(u2_u2__abc_47660_n539) );
  OR2X2 OR2X2_334 ( .A(u0__abc_49347_n1677_1), .B(u0__abc_49347_n1678_1), .Y(u0__abc_49347_n1679) );
  OR2X2 OR2X2_3340 ( .A(u2_u2__abc_47660_n159), .B(u2_u2_b3_last_row_4_), .Y(u2_u2__abc_47660_n543) );
  OR2X2 OR2X2_3341 ( .A(u2_u2__abc_47660_n544), .B(row_adr_4_bF_buf2), .Y(u2_u2__abc_47660_n545) );
  OR2X2 OR2X2_3342 ( .A(u2_u2__abc_47660_n547), .B(row_adr_3_bF_buf2), .Y(u2_u2__abc_47660_n548) );
  OR2X2 OR2X2_3343 ( .A(u2_u2__abc_47660_n551), .B(row_adr_0_bF_buf2), .Y(u2_u2__abc_47660_n552) );
  OR2X2 OR2X2_3344 ( .A(u2_u2__abc_47660_n139), .B(u2_u2_b3_last_row_0_), .Y(u2_u2__abc_47660_n553) );
  OR2X2 OR2X2_3345 ( .A(u2_u2__abc_47660_n555), .B(row_adr_2_bF_buf2), .Y(u2_u2__abc_47660_n556) );
  OR2X2 OR2X2_3346 ( .A(u2_u2__abc_47660_n149), .B(u2_u2_b3_last_row_2_), .Y(u2_u2__abc_47660_n557) );
  OR2X2 OR2X2_3347 ( .A(u2_u2__abc_47660_n174), .B(u2_u2_b3_last_row_7_), .Y(u2_u2__abc_47660_n562) );
  OR2X2 OR2X2_3348 ( .A(u2_u2__abc_47660_n563), .B(row_adr_7_bF_buf2), .Y(u2_u2__abc_47660_n564) );
  OR2X2 OR2X2_3349 ( .A(u2_u2__abc_47660_n566), .B(row_adr_10_bF_buf2), .Y(u2_u2__abc_47660_n567) );
  OR2X2 OR2X2_335 ( .A(u0__abc_49347_n1681), .B(spec_req_cs_0_bF_buf0), .Y(u0__abc_49347_n1682) );
  OR2X2 OR2X2_3350 ( .A(u2_u2__abc_47660_n179), .B(u2_u2_b3_last_row_8_), .Y(u2_u2__abc_47660_n568) );
  OR2X2 OR2X2_3351 ( .A(u2_u2__abc_47660_n169), .B(u2_u2_b3_last_row_6_), .Y(u2_u2__abc_47660_n571) );
  OR2X2 OR2X2_3352 ( .A(u2_u2__abc_47660_n572), .B(row_adr_6_bF_buf2), .Y(u2_u2__abc_47660_n573) );
  OR2X2 OR2X2_3353 ( .A(u2_u2__abc_47660_n575), .B(row_adr_5_bF_buf2), .Y(u2_u2__abc_47660_n576) );
  OR2X2 OR2X2_3354 ( .A(u2_u2__abc_47660_n154), .B(u2_u2_b3_last_row_3_), .Y(u2_u2__abc_47660_n577) );
  OR2X2 OR2X2_3355 ( .A(u2_u2__abc_47660_n164), .B(u2_u2_b3_last_row_5_), .Y(u2_u2__abc_47660_n580) );
  OR2X2 OR2X2_3356 ( .A(u2_u2__abc_47660_n581), .B(row_adr_1_bF_buf2), .Y(u2_u2__abc_47660_n582) );
  OR2X2 OR2X2_3357 ( .A(u2_u2__abc_47660_n144), .B(u2_u2_b3_last_row_1_), .Y(u2_u2__abc_47660_n584) );
  OR2X2 OR2X2_3358 ( .A(u2_u2__abc_47660_n585), .B(row_adr_12_bF_buf2), .Y(u2_u2__abc_47660_n586) );
  OR2X2 OR2X2_3359 ( .A(u2_u2__abc_47660_n526), .B(u2_u2__abc_47660_n591), .Y(u2_u2__abc_47660_n592) );
  OR2X2 OR2X2_336 ( .A(u0__abc_49347_n1680), .B(u0__abc_49347_n1682), .Y(u0__abc_49347_n1683) );
  OR2X2 OR2X2_3360 ( .A(u2_u2__abc_47660_n461), .B(u2_u2__abc_47660_n592), .Y(u2_row_same_2) );
  OR2X2 OR2X2_3361 ( .A(u2_u2__abc_47660_n594), .B(u2_u2__abc_47660_n595), .Y(u2_u2__abc_47660_n596) );
  OR2X2 OR2X2_3362 ( .A(u2_u2__abc_47660_n598), .B(u2_u2__abc_47660_n597), .Y(u2_u2__abc_47660_n599) );
  OR2X2 OR2X2_3363 ( .A(u2_u2__abc_47660_n596), .B(u2_u2__abc_47660_n599), .Y(u2_bank_open_2) );
  OR2X2 OR2X2_3364 ( .A(u2_u2__abc_47660_n608), .B(u2_u2__abc_47660_n137_bF_buf3), .Y(u2_u2_bank3_open_FF_INPUT) );
  OR2X2 OR2X2_3365 ( .A(u2_u2__abc_47660_n611), .B(u2_u2__abc_47660_n610), .Y(u2_u2__abc_47660_n612) );
  OR2X2 OR2X2_3366 ( .A(u2_u2__abc_47660_n614), .B(u2_u2__abc_47660_n205), .Y(u2_u2_bank2_open_FF_INPUT) );
  OR2X2 OR2X2_3367 ( .A(u2_u2__abc_47660_n616), .B(u2_u2__abc_47660_n610), .Y(u2_u2__abc_47660_n617) );
  OR2X2 OR2X2_3368 ( .A(u2_u2__abc_47660_n619), .B(u2_u2__abc_47660_n248), .Y(u2_u2_bank1_open_FF_INPUT) );
  OR2X2 OR2X2_3369 ( .A(u2_u2__abc_47660_n621), .B(u2_u2__abc_47660_n610), .Y(u2_u2__abc_47660_n622) );
  OR2X2 OR2X2_337 ( .A(u0__abc_49347_n1203_bF_buf3), .B(u0_tms0_20_), .Y(u0__abc_49347_n1684) );
  OR2X2 OR2X2_3370 ( .A(u2_u2__abc_47660_n624), .B(u2_u2__abc_47660_n290_1), .Y(u2_u2_bank0_open_FF_INPUT) );
  OR2X2 OR2X2_3371 ( .A(u2_u3__abc_47660_n137_bF_buf4), .B(u2_u3_b3_last_row_0_), .Y(u2_u3__abc_47660_n138) );
  OR2X2 OR2X2_3372 ( .A(u2_u3__abc_47660_n137_bF_buf2), .B(u2_u3_b3_last_row_1_), .Y(u2_u3__abc_47660_n143) );
  OR2X2 OR2X2_3373 ( .A(u2_u3__abc_47660_n137_bF_buf0), .B(u2_u3_b3_last_row_2_), .Y(u2_u3__abc_47660_n148) );
  OR2X2 OR2X2_3374 ( .A(u2_u3__abc_47660_n137_bF_buf3), .B(u2_u3_b3_last_row_3_), .Y(u2_u3__abc_47660_n153) );
  OR2X2 OR2X2_3375 ( .A(u2_u3__abc_47660_n137_bF_buf1), .B(u2_u3_b3_last_row_4_), .Y(u2_u3__abc_47660_n158) );
  OR2X2 OR2X2_3376 ( .A(u2_u3__abc_47660_n137_bF_buf4), .B(u2_u3_b3_last_row_5_), .Y(u2_u3__abc_47660_n163) );
  OR2X2 OR2X2_3377 ( .A(u2_u3__abc_47660_n137_bF_buf2), .B(u2_u3_b3_last_row_6_), .Y(u2_u3__abc_47660_n168) );
  OR2X2 OR2X2_3378 ( .A(u2_u3__abc_47660_n137_bF_buf0), .B(u2_u3_b3_last_row_7_), .Y(u2_u3__abc_47660_n173) );
  OR2X2 OR2X2_3379 ( .A(u2_u3__abc_47660_n137_bF_buf3), .B(u2_u3_b3_last_row_8_), .Y(u2_u3__abc_47660_n178) );
  OR2X2 OR2X2_338 ( .A(u0__abc_49347_n1686_1), .B(u0__abc_49347_n1664), .Y(u0_sp_tms_20__FF_INPUT) );
  OR2X2 OR2X2_3380 ( .A(u2_u3__abc_47660_n137_bF_buf1), .B(u2_u3_b3_last_row_9_), .Y(u2_u3__abc_47660_n183) );
  OR2X2 OR2X2_3381 ( .A(u2_u3__abc_47660_n137_bF_buf4), .B(u2_u3_b3_last_row_10_), .Y(u2_u3__abc_47660_n188) );
  OR2X2 OR2X2_3382 ( .A(u2_u3__abc_47660_n137_bF_buf2), .B(u2_u3_b3_last_row_11_), .Y(u2_u3__abc_47660_n193) );
  OR2X2 OR2X2_3383 ( .A(u2_u3__abc_47660_n137_bF_buf0), .B(u2_u3_b3_last_row_12_), .Y(u2_u3__abc_47660_n198) );
  OR2X2 OR2X2_3384 ( .A(u2_u3__abc_47660_n205), .B(u2_u3_b2_last_row_0_), .Y(u2_u3__abc_47660_n206) );
  OR2X2 OR2X2_3385 ( .A(u2_u3__abc_47660_n207), .B(row_adr_0_bF_buf0), .Y(u2_u3__abc_47660_n208) );
  OR2X2 OR2X2_3386 ( .A(u2_u3__abc_47660_n205), .B(u2_u3_b2_last_row_1_), .Y(u2_u3__abc_47660_n210) );
  OR2X2 OR2X2_3387 ( .A(u2_u3__abc_47660_n207), .B(row_adr_1_bF_buf0), .Y(u2_u3__abc_47660_n211) );
  OR2X2 OR2X2_3388 ( .A(u2_u3__abc_47660_n205), .B(u2_u3_b2_last_row_2_), .Y(u2_u3__abc_47660_n213) );
  OR2X2 OR2X2_3389 ( .A(u2_u3__abc_47660_n207), .B(row_adr_2_bF_buf0), .Y(u2_u3__abc_47660_n214) );
  OR2X2 OR2X2_339 ( .A(u0__abc_49347_n1183_1_bF_buf2), .B(1'b0), .Y(u0__abc_49347_n1690) );
  OR2X2 OR2X2_3390 ( .A(u2_u3__abc_47660_n205), .B(u2_u3_b2_last_row_3_), .Y(u2_u3__abc_47660_n216) );
  OR2X2 OR2X2_3391 ( .A(u2_u3__abc_47660_n207), .B(row_adr_3_bF_buf0), .Y(u2_u3__abc_47660_n217) );
  OR2X2 OR2X2_3392 ( .A(u2_u3__abc_47660_n205), .B(u2_u3_b2_last_row_4_), .Y(u2_u3__abc_47660_n219) );
  OR2X2 OR2X2_3393 ( .A(u2_u3__abc_47660_n207), .B(row_adr_4_bF_buf0), .Y(u2_u3__abc_47660_n220) );
  OR2X2 OR2X2_3394 ( .A(u2_u3__abc_47660_n205), .B(u2_u3_b2_last_row_5_), .Y(u2_u3__abc_47660_n222) );
  OR2X2 OR2X2_3395 ( .A(u2_u3__abc_47660_n207), .B(row_adr_5_bF_buf0), .Y(u2_u3__abc_47660_n223) );
  OR2X2 OR2X2_3396 ( .A(u2_u3__abc_47660_n205), .B(u2_u3_b2_last_row_6_), .Y(u2_u3__abc_47660_n225) );
  OR2X2 OR2X2_3397 ( .A(u2_u3__abc_47660_n207), .B(row_adr_6_bF_buf0), .Y(u2_u3__abc_47660_n226) );
  OR2X2 OR2X2_3398 ( .A(u2_u3__abc_47660_n205), .B(u2_u3_b2_last_row_7_), .Y(u2_u3__abc_47660_n228) );
  OR2X2 OR2X2_3399 ( .A(u2_u3__abc_47660_n207), .B(row_adr_7_bF_buf0), .Y(u2_u3__abc_47660_n229) );
  OR2X2 OR2X2_34 ( .A(_abc_55805_n245_1), .B(cs_need_rfr_7_), .Y(_abc_55805_n288) );
  OR2X2 OR2X2_340 ( .A(spec_req_cs_6_bF_buf5), .B(1'b0), .Y(u0__abc_49347_n1691) );
  OR2X2 OR2X2_3400 ( .A(u2_u3__abc_47660_n205), .B(u2_u3_b2_last_row_8_), .Y(u2_u3__abc_47660_n231) );
  OR2X2 OR2X2_3401 ( .A(u2_u3__abc_47660_n207), .B(row_adr_8_bF_buf0), .Y(u2_u3__abc_47660_n232) );
  OR2X2 OR2X2_3402 ( .A(u2_u3__abc_47660_n205), .B(u2_u3_b2_last_row_9_), .Y(u2_u3__abc_47660_n234) );
  OR2X2 OR2X2_3403 ( .A(u2_u3__abc_47660_n207), .B(row_adr_9_bF_buf0), .Y(u2_u3__abc_47660_n235) );
  OR2X2 OR2X2_3404 ( .A(u2_u3__abc_47660_n205), .B(u2_u3_b2_last_row_10_), .Y(u2_u3__abc_47660_n237) );
  OR2X2 OR2X2_3405 ( .A(u2_u3__abc_47660_n207), .B(row_adr_10_bF_buf0), .Y(u2_u3__abc_47660_n238) );
  OR2X2 OR2X2_3406 ( .A(u2_u3__abc_47660_n205), .B(u2_u3_b2_last_row_11_), .Y(u2_u3__abc_47660_n240) );
  OR2X2 OR2X2_3407 ( .A(u2_u3__abc_47660_n207), .B(row_adr_11_bF_buf0), .Y(u2_u3__abc_47660_n241) );
  OR2X2 OR2X2_3408 ( .A(u2_u3__abc_47660_n205), .B(u2_u3_b2_last_row_12_), .Y(u2_u3__abc_47660_n243) );
  OR2X2 OR2X2_3409 ( .A(u2_u3__abc_47660_n207), .B(row_adr_12_bF_buf0), .Y(u2_u3__abc_47660_n244) );
  OR2X2 OR2X2_341 ( .A(u0__abc_49347_n1693), .B(u0__abc_49347_n1689), .Y(u0__abc_49347_n1694) );
  OR2X2 OR2X2_3410 ( .A(u2_u3__abc_47660_n248), .B(u2_u3_b1_last_row_0_), .Y(u2_u3__abc_47660_n249) );
  OR2X2 OR2X2_3411 ( .A(u2_u3__abc_47660_n250), .B(row_adr_0_bF_buf6), .Y(u2_u3__abc_47660_n251) );
  OR2X2 OR2X2_3412 ( .A(u2_u3__abc_47660_n248), .B(u2_u3_b1_last_row_1_), .Y(u2_u3__abc_47660_n253) );
  OR2X2 OR2X2_3413 ( .A(u2_u3__abc_47660_n250), .B(row_adr_1_bF_buf6), .Y(u2_u3__abc_47660_n254) );
  OR2X2 OR2X2_3414 ( .A(u2_u3__abc_47660_n248), .B(u2_u3_b1_last_row_2_), .Y(u2_u3__abc_47660_n256) );
  OR2X2 OR2X2_3415 ( .A(u2_u3__abc_47660_n250), .B(row_adr_2_bF_buf6), .Y(u2_u3__abc_47660_n257) );
  OR2X2 OR2X2_3416 ( .A(u2_u3__abc_47660_n248), .B(u2_u3_b1_last_row_3_), .Y(u2_u3__abc_47660_n259) );
  OR2X2 OR2X2_3417 ( .A(u2_u3__abc_47660_n250), .B(row_adr_3_bF_buf6), .Y(u2_u3__abc_47660_n260) );
  OR2X2 OR2X2_3418 ( .A(u2_u3__abc_47660_n248), .B(u2_u3_b1_last_row_4_), .Y(u2_u3__abc_47660_n262) );
  OR2X2 OR2X2_3419 ( .A(u2_u3__abc_47660_n250), .B(row_adr_4_bF_buf6), .Y(u2_u3__abc_47660_n263) );
  OR2X2 OR2X2_342 ( .A(u0__abc_49347_n1695_1), .B(u0__abc_49347_n1696_1), .Y(u0__abc_49347_n1697) );
  OR2X2 OR2X2_3420 ( .A(u2_u3__abc_47660_n248), .B(u2_u3_b1_last_row_5_), .Y(u2_u3__abc_47660_n265) );
  OR2X2 OR2X2_3421 ( .A(u2_u3__abc_47660_n250), .B(row_adr_5_bF_buf6), .Y(u2_u3__abc_47660_n266) );
  OR2X2 OR2X2_3422 ( .A(u2_u3__abc_47660_n248), .B(u2_u3_b1_last_row_6_), .Y(u2_u3__abc_47660_n268) );
  OR2X2 OR2X2_3423 ( .A(u2_u3__abc_47660_n250), .B(row_adr_6_bF_buf6), .Y(u2_u3__abc_47660_n269) );
  OR2X2 OR2X2_3424 ( .A(u2_u3__abc_47660_n248), .B(u2_u3_b1_last_row_7_), .Y(u2_u3__abc_47660_n271) );
  OR2X2 OR2X2_3425 ( .A(u2_u3__abc_47660_n250), .B(row_adr_7_bF_buf6), .Y(u2_u3__abc_47660_n272) );
  OR2X2 OR2X2_3426 ( .A(u2_u3__abc_47660_n248), .B(u2_u3_b1_last_row_8_), .Y(u2_u3__abc_47660_n274) );
  OR2X2 OR2X2_3427 ( .A(u2_u3__abc_47660_n250), .B(row_adr_8_bF_buf6), .Y(u2_u3__abc_47660_n275_1) );
  OR2X2 OR2X2_3428 ( .A(u2_u3__abc_47660_n248), .B(u2_u3_b1_last_row_9_), .Y(u2_u3__abc_47660_n277) );
  OR2X2 OR2X2_3429 ( .A(u2_u3__abc_47660_n250), .B(row_adr_9_bF_buf6), .Y(u2_u3__abc_47660_n278_1) );
  OR2X2 OR2X2_343 ( .A(u0__abc_49347_n1698), .B(u0__abc_49347_n1699), .Y(u0__abc_49347_n1700) );
  OR2X2 OR2X2_3430 ( .A(u2_u3__abc_47660_n248), .B(u2_u3_b1_last_row_10_), .Y(u2_u3__abc_47660_n280) );
  OR2X2 OR2X2_3431 ( .A(u2_u3__abc_47660_n250), .B(row_adr_10_bF_buf6), .Y(u2_u3__abc_47660_n281) );
  OR2X2 OR2X2_3432 ( .A(u2_u3__abc_47660_n248), .B(u2_u3_b1_last_row_11_), .Y(u2_u3__abc_47660_n283_1) );
  OR2X2 OR2X2_3433 ( .A(u2_u3__abc_47660_n250), .B(row_adr_11_bF_buf6), .Y(u2_u3__abc_47660_n284) );
  OR2X2 OR2X2_3434 ( .A(u2_u3__abc_47660_n248), .B(u2_u3_b1_last_row_12_), .Y(u2_u3__abc_47660_n286_1) );
  OR2X2 OR2X2_3435 ( .A(u2_u3__abc_47660_n250), .B(row_adr_12_bF_buf6), .Y(u2_u3__abc_47660_n287_1) );
  OR2X2 OR2X2_3436 ( .A(u2_u3__abc_47660_n290_1), .B(u2_u3_b0_last_row_0_), .Y(u2_u3__abc_47660_n291) );
  OR2X2 OR2X2_3437 ( .A(u2_u3__abc_47660_n292_1), .B(row_adr_0_bF_buf5), .Y(u2_u3__abc_47660_n293) );
  OR2X2 OR2X2_3438 ( .A(u2_u3__abc_47660_n290_1), .B(u2_u3_b0_last_row_1_), .Y(u2_u3__abc_47660_n295) );
  OR2X2 OR2X2_3439 ( .A(u2_u3__abc_47660_n292_1), .B(row_adr_1_bF_buf5), .Y(u2_u3__abc_47660_n296_1) );
  OR2X2 OR2X2_344 ( .A(u0__abc_49347_n1701), .B(u0__abc_49347_n1702), .Y(u0__abc_49347_n1703) );
  OR2X2 OR2X2_3440 ( .A(u2_u3__abc_47660_n290_1), .B(u2_u3_b0_last_row_2_), .Y(u2_u3__abc_47660_n298) );
  OR2X2 OR2X2_3441 ( .A(u2_u3__abc_47660_n292_1), .B(row_adr_2_bF_buf5), .Y(u2_u3__abc_47660_n299) );
  OR2X2 OR2X2_3442 ( .A(u2_u3__abc_47660_n290_1), .B(u2_u3_b0_last_row_3_), .Y(u2_u3__abc_47660_n301) );
  OR2X2 OR2X2_3443 ( .A(u2_u3__abc_47660_n292_1), .B(row_adr_3_bF_buf5), .Y(u2_u3__abc_47660_n302) );
  OR2X2 OR2X2_3444 ( .A(u2_u3__abc_47660_n290_1), .B(u2_u3_b0_last_row_4_), .Y(u2_u3__abc_47660_n304_1) );
  OR2X2 OR2X2_3445 ( .A(u2_u3__abc_47660_n292_1), .B(row_adr_4_bF_buf5), .Y(u2_u3__abc_47660_n305_1) );
  OR2X2 OR2X2_3446 ( .A(u2_u3__abc_47660_n290_1), .B(u2_u3_b0_last_row_5_), .Y(u2_u3__abc_47660_n307) );
  OR2X2 OR2X2_3447 ( .A(u2_u3__abc_47660_n292_1), .B(row_adr_5_bF_buf5), .Y(u2_u3__abc_47660_n308) );
  OR2X2 OR2X2_3448 ( .A(u2_u3__abc_47660_n290_1), .B(u2_u3_b0_last_row_6_), .Y(u2_u3__abc_47660_n310) );
  OR2X2 OR2X2_3449 ( .A(u2_u3__abc_47660_n292_1), .B(row_adr_6_bF_buf5), .Y(u2_u3__abc_47660_n311) );
  OR2X2 OR2X2_345 ( .A(u0__abc_49347_n1705_1), .B(spec_req_cs_0_bF_buf5), .Y(u0__abc_49347_n1706) );
  OR2X2 OR2X2_3450 ( .A(u2_u3__abc_47660_n290_1), .B(u2_u3_b0_last_row_7_), .Y(u2_u3__abc_47660_n313) );
  OR2X2 OR2X2_3451 ( .A(u2_u3__abc_47660_n292_1), .B(row_adr_7_bF_buf5), .Y(u2_u3__abc_47660_n314) );
  OR2X2 OR2X2_3452 ( .A(u2_u3__abc_47660_n290_1), .B(u2_u3_b0_last_row_8_), .Y(u2_u3__abc_47660_n316) );
  OR2X2 OR2X2_3453 ( .A(u2_u3__abc_47660_n292_1), .B(row_adr_8_bF_buf5), .Y(u2_u3__abc_47660_n317) );
  OR2X2 OR2X2_3454 ( .A(u2_u3__abc_47660_n290_1), .B(u2_u3_b0_last_row_9_), .Y(u2_u3__abc_47660_n319) );
  OR2X2 OR2X2_3455 ( .A(u2_u3__abc_47660_n292_1), .B(row_adr_9_bF_buf5), .Y(u2_u3__abc_47660_n320) );
  OR2X2 OR2X2_3456 ( .A(u2_u3__abc_47660_n290_1), .B(u2_u3_b0_last_row_10_), .Y(u2_u3__abc_47660_n322) );
  OR2X2 OR2X2_3457 ( .A(u2_u3__abc_47660_n292_1), .B(row_adr_10_bF_buf5), .Y(u2_u3__abc_47660_n323) );
  OR2X2 OR2X2_3458 ( .A(u2_u3__abc_47660_n290_1), .B(u2_u3_b0_last_row_11_), .Y(u2_u3__abc_47660_n325) );
  OR2X2 OR2X2_3459 ( .A(u2_u3__abc_47660_n292_1), .B(row_adr_11_bF_buf5), .Y(u2_u3__abc_47660_n326) );
  OR2X2 OR2X2_346 ( .A(u0__abc_49347_n1704_1), .B(u0__abc_49347_n1706), .Y(u0__abc_49347_n1707) );
  OR2X2 OR2X2_3460 ( .A(u2_u3__abc_47660_n290_1), .B(u2_u3_b0_last_row_12_), .Y(u2_u3__abc_47660_n328) );
  OR2X2 OR2X2_3461 ( .A(u2_u3__abc_47660_n292_1), .B(row_adr_12_bF_buf5), .Y(u2_u3__abc_47660_n329) );
  OR2X2 OR2X2_3462 ( .A(u2_u3__abc_47660_n331), .B(row_adr_12_bF_buf4), .Y(u2_u3__abc_47660_n332) );
  OR2X2 OR2X2_3463 ( .A(u2_u3__abc_47660_n333), .B(row_adr_11_bF_buf4), .Y(u2_u3__abc_47660_n334) );
  OR2X2 OR2X2_3464 ( .A(u2_u3__abc_47660_n199), .B(u2_u3_b0_last_row_12_), .Y(u2_u3__abc_47660_n335) );
  OR2X2 OR2X2_3465 ( .A(u2_u3__abc_47660_n194), .B(u2_u3_b0_last_row_11_), .Y(u2_u3__abc_47660_n338) );
  OR2X2 OR2X2_3466 ( .A(u2_u3__abc_47660_n339), .B(row_adr_9_bF_buf4), .Y(u2_u3__abc_47660_n340) );
  OR2X2 OR2X2_3467 ( .A(u2_u3__abc_47660_n184), .B(u2_u3_b0_last_row_9_), .Y(u2_u3__abc_47660_n342) );
  OR2X2 OR2X2_3468 ( .A(u2_u3__abc_47660_n343), .B(row_adr_7_bF_buf4), .Y(u2_u3__abc_47660_n344) );
  OR2X2 OR2X2_3469 ( .A(u2_u3__abc_47660_n164), .B(u2_u3_b0_last_row_5_), .Y(u2_u3__abc_47660_n348) );
  OR2X2 OR2X2_347 ( .A(u0__abc_49347_n1203_bF_buf2), .B(u0_tms0_21_), .Y(u0__abc_49347_n1708) );
  OR2X2 OR2X2_3470 ( .A(u2_u3__abc_47660_n159), .B(u2_u3_b0_last_row_4_), .Y(u2_u3__abc_47660_n350) );
  OR2X2 OR2X2_3471 ( .A(u2_u3__abc_47660_n351), .B(row_adr_4_bF_buf4), .Y(u2_u3__abc_47660_n352) );
  OR2X2 OR2X2_3472 ( .A(u2_u3__abc_47660_n355), .B(row_adr_0_bF_buf4), .Y(u2_u3__abc_47660_n356) );
  OR2X2 OR2X2_3473 ( .A(u2_u3__abc_47660_n139), .B(u2_u3_b0_last_row_0_), .Y(u2_u3__abc_47660_n357) );
  OR2X2 OR2X2_3474 ( .A(u2_u3__abc_47660_n144), .B(u2_u3_b0_last_row_1_), .Y(u2_u3__abc_47660_n359) );
  OR2X2 OR2X2_3475 ( .A(u2_u3__abc_47660_n360), .B(row_adr_5_bF_buf4), .Y(u2_u3__abc_47660_n361) );
  OR2X2 OR2X2_3476 ( .A(u2_u3__abc_47660_n366), .B(row_adr_10_bF_buf4), .Y(u2_u3__abc_47660_n367) );
  OR2X2 OR2X2_3477 ( .A(u2_u3__abc_47660_n189), .B(u2_u3_b0_last_row_10_), .Y(u2_u3__abc_47660_n368) );
  OR2X2 OR2X2_3478 ( .A(u2_u3__abc_47660_n372), .B(u2_u3__abc_47660_n370), .Y(u2_u3__abc_47660_n373) );
  OR2X2 OR2X2_3479 ( .A(u2_u3__abc_47660_n154), .B(u2_u3_b0_last_row_3_), .Y(u2_u3__abc_47660_n375) );
  OR2X2 OR2X2_348 ( .A(u0__abc_49347_n1710), .B(u0__abc_49347_n1688), .Y(u0_sp_tms_21__FF_INPUT) );
  OR2X2 OR2X2_3480 ( .A(u2_u3__abc_47660_n376), .B(row_adr_2_bF_buf4), .Y(u2_u3__abc_47660_n377) );
  OR2X2 OR2X2_3481 ( .A(u2_u3__abc_47660_n379), .B(row_adr_1_bF_buf4), .Y(u2_u3__abc_47660_n380) );
  OR2X2 OR2X2_3482 ( .A(u2_u3__abc_47660_n149), .B(u2_u3_b0_last_row_2_), .Y(u2_u3__abc_47660_n381) );
  OR2X2 OR2X2_3483 ( .A(u2_u3__abc_47660_n384), .B(row_adr_3_bF_buf4), .Y(u2_u3__abc_47660_n385) );
  OR2X2 OR2X2_3484 ( .A(u2_u3__abc_47660_n174), .B(u2_u3_b0_last_row_7_), .Y(u2_u3__abc_47660_n386) );
  OR2X2 OR2X2_3485 ( .A(u2_u3__abc_47660_n390), .B(u2_u3__abc_47660_n388), .Y(u2_u3__abc_47660_n391) );
  OR2X2 OR2X2_3486 ( .A(u2_u3__abc_47660_n396), .B(row_adr_12_bF_buf3), .Y(u2_u3__abc_47660_n397) );
  OR2X2 OR2X2_3487 ( .A(u2_u3__abc_47660_n398), .B(row_adr_11_bF_buf3), .Y(u2_u3__abc_47660_n399) );
  OR2X2 OR2X2_3488 ( .A(u2_u3__abc_47660_n199), .B(u2_u3_b2_last_row_12_), .Y(u2_u3__abc_47660_n400) );
  OR2X2 OR2X2_3489 ( .A(u2_u3__abc_47660_n194), .B(u2_u3_b2_last_row_11_), .Y(u2_u3__abc_47660_n403) );
  OR2X2 OR2X2_349 ( .A(u0__abc_49347_n1183_1_bF_buf1), .B(1'b0), .Y(u0__abc_49347_n1714_1) );
  OR2X2 OR2X2_3490 ( .A(u2_u3__abc_47660_n404), .B(row_adr_9_bF_buf3), .Y(u2_u3__abc_47660_n405) );
  OR2X2 OR2X2_3491 ( .A(u2_u3__abc_47660_n184), .B(u2_u3_b2_last_row_9_), .Y(u2_u3__abc_47660_n407) );
  OR2X2 OR2X2_3492 ( .A(u2_u3__abc_47660_n408), .B(row_adr_7_bF_buf3), .Y(u2_u3__abc_47660_n409) );
  OR2X2 OR2X2_3493 ( .A(u2_u3__abc_47660_n164), .B(u2_u3_b2_last_row_5_), .Y(u2_u3__abc_47660_n413) );
  OR2X2 OR2X2_3494 ( .A(u2_u3__abc_47660_n159), .B(u2_u3_b2_last_row_4_), .Y(u2_u3__abc_47660_n415) );
  OR2X2 OR2X2_3495 ( .A(u2_u3__abc_47660_n416), .B(row_adr_4_bF_buf3), .Y(u2_u3__abc_47660_n417) );
  OR2X2 OR2X2_3496 ( .A(u2_u3__abc_47660_n420), .B(row_adr_0_bF_buf3), .Y(u2_u3__abc_47660_n421) );
  OR2X2 OR2X2_3497 ( .A(u2_u3__abc_47660_n139), .B(u2_u3_b2_last_row_0_), .Y(u2_u3__abc_47660_n422) );
  OR2X2 OR2X2_3498 ( .A(u2_u3__abc_47660_n144), .B(u2_u3_b2_last_row_1_), .Y(u2_u3__abc_47660_n424) );
  OR2X2 OR2X2_3499 ( .A(u2_u3__abc_47660_n425), .B(row_adr_5_bF_buf3), .Y(u2_u3__abc_47660_n426) );
  OR2X2 OR2X2_35 ( .A(_abc_55805_n240_bF_buf3), .B(sp_tms_0_), .Y(_abc_55805_n290) );
  OR2X2 OR2X2_350 ( .A(spec_req_cs_6_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n1715) );
  OR2X2 OR2X2_3500 ( .A(u2_u3__abc_47660_n431), .B(row_adr_10_bF_buf3), .Y(u2_u3__abc_47660_n432) );
  OR2X2 OR2X2_3501 ( .A(u2_u3__abc_47660_n189), .B(u2_u3_b2_last_row_10_), .Y(u2_u3__abc_47660_n433) );
  OR2X2 OR2X2_3502 ( .A(u2_u3__abc_47660_n437), .B(u2_u3__abc_47660_n435), .Y(u2_u3__abc_47660_n438) );
  OR2X2 OR2X2_3503 ( .A(u2_u3__abc_47660_n154), .B(u2_u3_b2_last_row_3_), .Y(u2_u3__abc_47660_n440) );
  OR2X2 OR2X2_3504 ( .A(u2_u3__abc_47660_n441), .B(row_adr_2_bF_buf3), .Y(u2_u3__abc_47660_n442) );
  OR2X2 OR2X2_3505 ( .A(u2_u3__abc_47660_n444), .B(row_adr_1_bF_buf3), .Y(u2_u3__abc_47660_n445) );
  OR2X2 OR2X2_3506 ( .A(u2_u3__abc_47660_n149), .B(u2_u3_b2_last_row_2_), .Y(u2_u3__abc_47660_n446) );
  OR2X2 OR2X2_3507 ( .A(u2_u3__abc_47660_n449), .B(row_adr_3_bF_buf3), .Y(u2_u3__abc_47660_n450) );
  OR2X2 OR2X2_3508 ( .A(u2_u3__abc_47660_n174), .B(u2_u3_b2_last_row_7_), .Y(u2_u3__abc_47660_n451) );
  OR2X2 OR2X2_3509 ( .A(u2_u3__abc_47660_n455), .B(u2_u3__abc_47660_n453), .Y(u2_u3__abc_47660_n456) );
  OR2X2 OR2X2_351 ( .A(u0__abc_49347_n1717), .B(u0__abc_49347_n1713_1), .Y(u0__abc_49347_n1718) );
  OR2X2 OR2X2_3510 ( .A(u2_u3__abc_47660_n395), .B(u2_u3__abc_47660_n460), .Y(u2_u3__abc_47660_n461) );
  OR2X2 OR2X2_3511 ( .A(u2_u3__abc_47660_n462), .B(row_adr_12_bF_buf2), .Y(u2_u3__abc_47660_n463) );
  OR2X2 OR2X2_3512 ( .A(u2_u3__abc_47660_n464), .B(row_adr_11_bF_buf2), .Y(u2_u3__abc_47660_n465) );
  OR2X2 OR2X2_3513 ( .A(u2_u3__abc_47660_n199), .B(u2_u3_b1_last_row_12_), .Y(u2_u3__abc_47660_n466) );
  OR2X2 OR2X2_3514 ( .A(u2_u3__abc_47660_n194), .B(u2_u3_b1_last_row_11_), .Y(u2_u3__abc_47660_n469) );
  OR2X2 OR2X2_3515 ( .A(u2_u3__abc_47660_n470), .B(row_adr_9_bF_buf2), .Y(u2_u3__abc_47660_n471) );
  OR2X2 OR2X2_3516 ( .A(u2_u3__abc_47660_n184), .B(u2_u3_b1_last_row_9_), .Y(u2_u3__abc_47660_n473) );
  OR2X2 OR2X2_3517 ( .A(u2_u3__abc_47660_n474), .B(row_adr_7_bF_buf2), .Y(u2_u3__abc_47660_n475) );
  OR2X2 OR2X2_3518 ( .A(u2_u3__abc_47660_n164), .B(u2_u3_b1_last_row_5_), .Y(u2_u3__abc_47660_n479) );
  OR2X2 OR2X2_3519 ( .A(u2_u3__abc_47660_n159), .B(u2_u3_b1_last_row_4_), .Y(u2_u3__abc_47660_n481) );
  OR2X2 OR2X2_352 ( .A(u0__abc_49347_n1719), .B(u0__abc_49347_n1720), .Y(u0__abc_49347_n1721) );
  OR2X2 OR2X2_3520 ( .A(u2_u3__abc_47660_n482), .B(row_adr_4_bF_buf2), .Y(u2_u3__abc_47660_n483) );
  OR2X2 OR2X2_3521 ( .A(u2_u3__abc_47660_n486), .B(row_adr_0_bF_buf2), .Y(u2_u3__abc_47660_n487) );
  OR2X2 OR2X2_3522 ( .A(u2_u3__abc_47660_n139), .B(u2_u3_b1_last_row_0_), .Y(u2_u3__abc_47660_n488) );
  OR2X2 OR2X2_3523 ( .A(u2_u3__abc_47660_n144), .B(u2_u3_b1_last_row_1_), .Y(u2_u3__abc_47660_n490) );
  OR2X2 OR2X2_3524 ( .A(u2_u3__abc_47660_n491), .B(row_adr_5_bF_buf2), .Y(u2_u3__abc_47660_n492) );
  OR2X2 OR2X2_3525 ( .A(u2_u3__abc_47660_n497), .B(row_adr_10_bF_buf2), .Y(u2_u3__abc_47660_n498) );
  OR2X2 OR2X2_3526 ( .A(u2_u3__abc_47660_n189), .B(u2_u3_b1_last_row_10_), .Y(u2_u3__abc_47660_n499) );
  OR2X2 OR2X2_3527 ( .A(u2_u3__abc_47660_n503), .B(u2_u3__abc_47660_n501), .Y(u2_u3__abc_47660_n504) );
  OR2X2 OR2X2_3528 ( .A(u2_u3__abc_47660_n154), .B(u2_u3_b1_last_row_3_), .Y(u2_u3__abc_47660_n506) );
  OR2X2 OR2X2_3529 ( .A(u2_u3__abc_47660_n507), .B(row_adr_2_bF_buf2), .Y(u2_u3__abc_47660_n508) );
  OR2X2 OR2X2_353 ( .A(u0__abc_49347_n1722_1), .B(u0__abc_49347_n1723_1), .Y(u0__abc_49347_n1724) );
  OR2X2 OR2X2_3530 ( .A(u2_u3__abc_47660_n510), .B(row_adr_1_bF_buf2), .Y(u2_u3__abc_47660_n511) );
  OR2X2 OR2X2_3531 ( .A(u2_u3__abc_47660_n149), .B(u2_u3_b1_last_row_2_), .Y(u2_u3__abc_47660_n512) );
  OR2X2 OR2X2_3532 ( .A(u2_u3__abc_47660_n515), .B(row_adr_3_bF_buf2), .Y(u2_u3__abc_47660_n516) );
  OR2X2 OR2X2_3533 ( .A(u2_u3__abc_47660_n174), .B(u2_u3_b1_last_row_7_), .Y(u2_u3__abc_47660_n517) );
  OR2X2 OR2X2_3534 ( .A(u2_u3__abc_47660_n521), .B(u2_u3__abc_47660_n519), .Y(u2_u3__abc_47660_n522) );
  OR2X2 OR2X2_3535 ( .A(u2_u3__abc_47660_n527), .B(row_adr_9_bF_buf1), .Y(u2_u3__abc_47660_n528) );
  OR2X2 OR2X2_3536 ( .A(u2_u3__abc_47660_n189), .B(u2_u3_b3_last_row_10_), .Y(u2_u3__abc_47660_n529) );
  OR2X2 OR2X2_3537 ( .A(u2_u3__abc_47660_n184), .B(u2_u3_b3_last_row_9_), .Y(u2_u3__abc_47660_n530) );
  OR2X2 OR2X2_3538 ( .A(u2_u3__abc_47660_n194), .B(u2_u3_b3_last_row_11_), .Y(u2_u3__abc_47660_n533) );
  OR2X2 OR2X2_3539 ( .A(u2_u3__abc_47660_n534), .B(row_adr_11_bF_buf1), .Y(u2_u3__abc_47660_n535) );
  OR2X2 OR2X2_354 ( .A(u0__abc_49347_n1725), .B(u0__abc_49347_n1726), .Y(u0__abc_49347_n1727) );
  OR2X2 OR2X2_3540 ( .A(u2_u3__abc_47660_n199), .B(u2_u3_b3_last_row_12_), .Y(u2_u3__abc_47660_n537) );
  OR2X2 OR2X2_3541 ( .A(u2_u3__abc_47660_n538), .B(row_adr_8_bF_buf1), .Y(u2_u3__abc_47660_n539) );
  OR2X2 OR2X2_3542 ( .A(u2_u3__abc_47660_n159), .B(u2_u3_b3_last_row_4_), .Y(u2_u3__abc_47660_n543) );
  OR2X2 OR2X2_3543 ( .A(u2_u3__abc_47660_n544), .B(row_adr_4_bF_buf1), .Y(u2_u3__abc_47660_n545) );
  OR2X2 OR2X2_3544 ( .A(u2_u3__abc_47660_n547), .B(row_adr_3_bF_buf1), .Y(u2_u3__abc_47660_n548) );
  OR2X2 OR2X2_3545 ( .A(u2_u3__abc_47660_n551), .B(row_adr_0_bF_buf1), .Y(u2_u3__abc_47660_n552) );
  OR2X2 OR2X2_3546 ( .A(u2_u3__abc_47660_n139), .B(u2_u3_b3_last_row_0_), .Y(u2_u3__abc_47660_n553) );
  OR2X2 OR2X2_3547 ( .A(u2_u3__abc_47660_n555), .B(row_adr_2_bF_buf1), .Y(u2_u3__abc_47660_n556) );
  OR2X2 OR2X2_3548 ( .A(u2_u3__abc_47660_n149), .B(u2_u3_b3_last_row_2_), .Y(u2_u3__abc_47660_n557) );
  OR2X2 OR2X2_3549 ( .A(u2_u3__abc_47660_n174), .B(u2_u3_b3_last_row_7_), .Y(u2_u3__abc_47660_n562) );
  OR2X2 OR2X2_355 ( .A(u0__abc_49347_n1729), .B(spec_req_cs_0_bF_buf4), .Y(u0__abc_49347_n1730) );
  OR2X2 OR2X2_3550 ( .A(u2_u3__abc_47660_n563), .B(row_adr_7_bF_buf1), .Y(u2_u3__abc_47660_n564) );
  OR2X2 OR2X2_3551 ( .A(u2_u3__abc_47660_n566), .B(row_adr_10_bF_buf1), .Y(u2_u3__abc_47660_n567) );
  OR2X2 OR2X2_3552 ( .A(u2_u3__abc_47660_n179), .B(u2_u3_b3_last_row_8_), .Y(u2_u3__abc_47660_n568) );
  OR2X2 OR2X2_3553 ( .A(u2_u3__abc_47660_n169), .B(u2_u3_b3_last_row_6_), .Y(u2_u3__abc_47660_n571) );
  OR2X2 OR2X2_3554 ( .A(u2_u3__abc_47660_n572), .B(row_adr_6_bF_buf1), .Y(u2_u3__abc_47660_n573) );
  OR2X2 OR2X2_3555 ( .A(u2_u3__abc_47660_n575), .B(row_adr_5_bF_buf1), .Y(u2_u3__abc_47660_n576) );
  OR2X2 OR2X2_3556 ( .A(u2_u3__abc_47660_n154), .B(u2_u3_b3_last_row_3_), .Y(u2_u3__abc_47660_n577) );
  OR2X2 OR2X2_3557 ( .A(u2_u3__abc_47660_n164), .B(u2_u3_b3_last_row_5_), .Y(u2_u3__abc_47660_n580) );
  OR2X2 OR2X2_3558 ( .A(u2_u3__abc_47660_n581), .B(row_adr_1_bF_buf1), .Y(u2_u3__abc_47660_n582) );
  OR2X2 OR2X2_3559 ( .A(u2_u3__abc_47660_n144), .B(u2_u3_b3_last_row_1_), .Y(u2_u3__abc_47660_n584) );
  OR2X2 OR2X2_356 ( .A(u0__abc_49347_n1728), .B(u0__abc_49347_n1730), .Y(u0__abc_49347_n1731_1) );
  OR2X2 OR2X2_3560 ( .A(u2_u3__abc_47660_n585), .B(row_adr_12_bF_buf1), .Y(u2_u3__abc_47660_n586) );
  OR2X2 OR2X2_3561 ( .A(u2_u3__abc_47660_n526), .B(u2_u3__abc_47660_n591), .Y(u2_u3__abc_47660_n592) );
  OR2X2 OR2X2_3562 ( .A(u2_u3__abc_47660_n461), .B(u2_u3__abc_47660_n592), .Y(u2_row_same_3) );
  OR2X2 OR2X2_3563 ( .A(u2_u3__abc_47660_n594), .B(u2_u3__abc_47660_n595), .Y(u2_u3__abc_47660_n596) );
  OR2X2 OR2X2_3564 ( .A(u2_u3__abc_47660_n598), .B(u2_u3__abc_47660_n597), .Y(u2_u3__abc_47660_n599) );
  OR2X2 OR2X2_3565 ( .A(u2_u3__abc_47660_n596), .B(u2_u3__abc_47660_n599), .Y(u2_bank_open_3) );
  OR2X2 OR2X2_3566 ( .A(u2_u3__abc_47660_n608), .B(u2_u3__abc_47660_n137_bF_buf3), .Y(u2_u3_bank3_open_FF_INPUT) );
  OR2X2 OR2X2_3567 ( .A(u2_u3__abc_47660_n611), .B(u2_u3__abc_47660_n610), .Y(u2_u3__abc_47660_n612) );
  OR2X2 OR2X2_3568 ( .A(u2_u3__abc_47660_n614), .B(u2_u3__abc_47660_n205), .Y(u2_u3_bank2_open_FF_INPUT) );
  OR2X2 OR2X2_3569 ( .A(u2_u3__abc_47660_n616), .B(u2_u3__abc_47660_n610), .Y(u2_u3__abc_47660_n617) );
  OR2X2 OR2X2_357 ( .A(u0__abc_49347_n1203_bF_buf1), .B(u0_tms0_22_), .Y(u0__abc_49347_n1732_1) );
  OR2X2 OR2X2_3570 ( .A(u2_u3__abc_47660_n619), .B(u2_u3__abc_47660_n248), .Y(u2_u3_bank1_open_FF_INPUT) );
  OR2X2 OR2X2_3571 ( .A(u2_u3__abc_47660_n621), .B(u2_u3__abc_47660_n610), .Y(u2_u3__abc_47660_n622) );
  OR2X2 OR2X2_3572 ( .A(u2_u3__abc_47660_n624), .B(u2_u3__abc_47660_n290_1), .Y(u2_u3_bank0_open_FF_INPUT) );
  OR2X2 OR2X2_3573 ( .A(u2_u4__abc_47660_n137_bF_buf4), .B(u2_u4_b3_last_row_0_), .Y(u2_u4__abc_47660_n138) );
  OR2X2 OR2X2_3574 ( .A(u2_u4__abc_47660_n137_bF_buf2), .B(u2_u4_b3_last_row_1_), .Y(u2_u4__abc_47660_n143) );
  OR2X2 OR2X2_3575 ( .A(u2_u4__abc_47660_n137_bF_buf0), .B(u2_u4_b3_last_row_2_), .Y(u2_u4__abc_47660_n148) );
  OR2X2 OR2X2_3576 ( .A(u2_u4__abc_47660_n137_bF_buf3), .B(u2_u4_b3_last_row_3_), .Y(u2_u4__abc_47660_n153) );
  OR2X2 OR2X2_3577 ( .A(u2_u4__abc_47660_n137_bF_buf1), .B(u2_u4_b3_last_row_4_), .Y(u2_u4__abc_47660_n158) );
  OR2X2 OR2X2_3578 ( .A(u2_u4__abc_47660_n137_bF_buf4), .B(u2_u4_b3_last_row_5_), .Y(u2_u4__abc_47660_n163) );
  OR2X2 OR2X2_3579 ( .A(u2_u4__abc_47660_n137_bF_buf2), .B(u2_u4_b3_last_row_6_), .Y(u2_u4__abc_47660_n168) );
  OR2X2 OR2X2_358 ( .A(u0__abc_49347_n1734), .B(u0__abc_49347_n1712), .Y(u0_sp_tms_22__FF_INPUT) );
  OR2X2 OR2X2_3580 ( .A(u2_u4__abc_47660_n137_bF_buf0), .B(u2_u4_b3_last_row_7_), .Y(u2_u4__abc_47660_n173) );
  OR2X2 OR2X2_3581 ( .A(u2_u4__abc_47660_n137_bF_buf3), .B(u2_u4_b3_last_row_8_), .Y(u2_u4__abc_47660_n178) );
  OR2X2 OR2X2_3582 ( .A(u2_u4__abc_47660_n137_bF_buf1), .B(u2_u4_b3_last_row_9_), .Y(u2_u4__abc_47660_n183) );
  OR2X2 OR2X2_3583 ( .A(u2_u4__abc_47660_n137_bF_buf4), .B(u2_u4_b3_last_row_10_), .Y(u2_u4__abc_47660_n188) );
  OR2X2 OR2X2_3584 ( .A(u2_u4__abc_47660_n137_bF_buf2), .B(u2_u4_b3_last_row_11_), .Y(u2_u4__abc_47660_n193) );
  OR2X2 OR2X2_3585 ( .A(u2_u4__abc_47660_n137_bF_buf0), .B(u2_u4_b3_last_row_12_), .Y(u2_u4__abc_47660_n198) );
  OR2X2 OR2X2_3586 ( .A(u2_u4__abc_47660_n205), .B(u2_u4_b2_last_row_0_), .Y(u2_u4__abc_47660_n206) );
  OR2X2 OR2X2_3587 ( .A(u2_u4__abc_47660_n207), .B(row_adr_0_bF_buf6), .Y(u2_u4__abc_47660_n208) );
  OR2X2 OR2X2_3588 ( .A(u2_u4__abc_47660_n205), .B(u2_u4_b2_last_row_1_), .Y(u2_u4__abc_47660_n210) );
  OR2X2 OR2X2_3589 ( .A(u2_u4__abc_47660_n207), .B(row_adr_1_bF_buf6), .Y(u2_u4__abc_47660_n211) );
  OR2X2 OR2X2_359 ( .A(u0__abc_49347_n1183_1_bF_buf0), .B(1'b0), .Y(u0__abc_49347_n1738) );
  OR2X2 OR2X2_3590 ( .A(u2_u4__abc_47660_n205), .B(u2_u4_b2_last_row_2_), .Y(u2_u4__abc_47660_n213) );
  OR2X2 OR2X2_3591 ( .A(u2_u4__abc_47660_n207), .B(row_adr_2_bF_buf6), .Y(u2_u4__abc_47660_n214) );
  OR2X2 OR2X2_3592 ( .A(u2_u4__abc_47660_n205), .B(u2_u4_b2_last_row_3_), .Y(u2_u4__abc_47660_n216) );
  OR2X2 OR2X2_3593 ( .A(u2_u4__abc_47660_n207), .B(row_adr_3_bF_buf6), .Y(u2_u4__abc_47660_n217) );
  OR2X2 OR2X2_3594 ( .A(u2_u4__abc_47660_n205), .B(u2_u4_b2_last_row_4_), .Y(u2_u4__abc_47660_n219) );
  OR2X2 OR2X2_3595 ( .A(u2_u4__abc_47660_n207), .B(row_adr_4_bF_buf6), .Y(u2_u4__abc_47660_n220) );
  OR2X2 OR2X2_3596 ( .A(u2_u4__abc_47660_n205), .B(u2_u4_b2_last_row_5_), .Y(u2_u4__abc_47660_n222) );
  OR2X2 OR2X2_3597 ( .A(u2_u4__abc_47660_n207), .B(row_adr_5_bF_buf6), .Y(u2_u4__abc_47660_n223) );
  OR2X2 OR2X2_3598 ( .A(u2_u4__abc_47660_n205), .B(u2_u4_b2_last_row_6_), .Y(u2_u4__abc_47660_n225) );
  OR2X2 OR2X2_3599 ( .A(u2_u4__abc_47660_n207), .B(row_adr_6_bF_buf6), .Y(u2_u4__abc_47660_n226) );
  OR2X2 OR2X2_36 ( .A(lmr_sel_bF_buf5), .B(tms_0_), .Y(_abc_55805_n291) );
  OR2X2 OR2X2_360 ( .A(spec_req_cs_6_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n1739) );
  OR2X2 OR2X2_3600 ( .A(u2_u4__abc_47660_n205), .B(u2_u4_b2_last_row_7_), .Y(u2_u4__abc_47660_n228) );
  OR2X2 OR2X2_3601 ( .A(u2_u4__abc_47660_n207), .B(row_adr_7_bF_buf6), .Y(u2_u4__abc_47660_n229) );
  OR2X2 OR2X2_3602 ( .A(u2_u4__abc_47660_n205), .B(u2_u4_b2_last_row_8_), .Y(u2_u4__abc_47660_n231) );
  OR2X2 OR2X2_3603 ( .A(u2_u4__abc_47660_n207), .B(row_adr_8_bF_buf6), .Y(u2_u4__abc_47660_n232) );
  OR2X2 OR2X2_3604 ( .A(u2_u4__abc_47660_n205), .B(u2_u4_b2_last_row_9_), .Y(u2_u4__abc_47660_n234) );
  OR2X2 OR2X2_3605 ( .A(u2_u4__abc_47660_n207), .B(row_adr_9_bF_buf6), .Y(u2_u4__abc_47660_n235) );
  OR2X2 OR2X2_3606 ( .A(u2_u4__abc_47660_n205), .B(u2_u4_b2_last_row_10_), .Y(u2_u4__abc_47660_n237) );
  OR2X2 OR2X2_3607 ( .A(u2_u4__abc_47660_n207), .B(row_adr_10_bF_buf6), .Y(u2_u4__abc_47660_n238) );
  OR2X2 OR2X2_3608 ( .A(u2_u4__abc_47660_n205), .B(u2_u4_b2_last_row_11_), .Y(u2_u4__abc_47660_n240) );
  OR2X2 OR2X2_3609 ( .A(u2_u4__abc_47660_n207), .B(row_adr_11_bF_buf6), .Y(u2_u4__abc_47660_n241) );
  OR2X2 OR2X2_361 ( .A(u0__abc_49347_n1741_1), .B(u0__abc_49347_n1737), .Y(u0__abc_49347_n1742) );
  OR2X2 OR2X2_3610 ( .A(u2_u4__abc_47660_n205), .B(u2_u4_b2_last_row_12_), .Y(u2_u4__abc_47660_n243) );
  OR2X2 OR2X2_3611 ( .A(u2_u4__abc_47660_n207), .B(row_adr_12_bF_buf6), .Y(u2_u4__abc_47660_n244) );
  OR2X2 OR2X2_3612 ( .A(u2_u4__abc_47660_n248), .B(u2_u4_b1_last_row_0_), .Y(u2_u4__abc_47660_n249) );
  OR2X2 OR2X2_3613 ( .A(u2_u4__abc_47660_n250), .B(row_adr_0_bF_buf5), .Y(u2_u4__abc_47660_n251) );
  OR2X2 OR2X2_3614 ( .A(u2_u4__abc_47660_n248), .B(u2_u4_b1_last_row_1_), .Y(u2_u4__abc_47660_n253) );
  OR2X2 OR2X2_3615 ( .A(u2_u4__abc_47660_n250), .B(row_adr_1_bF_buf5), .Y(u2_u4__abc_47660_n254) );
  OR2X2 OR2X2_3616 ( .A(u2_u4__abc_47660_n248), .B(u2_u4_b1_last_row_2_), .Y(u2_u4__abc_47660_n256) );
  OR2X2 OR2X2_3617 ( .A(u2_u4__abc_47660_n250), .B(row_adr_2_bF_buf5), .Y(u2_u4__abc_47660_n257) );
  OR2X2 OR2X2_3618 ( .A(u2_u4__abc_47660_n248), .B(u2_u4_b1_last_row_3_), .Y(u2_u4__abc_47660_n259) );
  OR2X2 OR2X2_3619 ( .A(u2_u4__abc_47660_n250), .B(row_adr_3_bF_buf5), .Y(u2_u4__abc_47660_n260) );
  OR2X2 OR2X2_362 ( .A(u0__abc_49347_n1743), .B(u0__abc_49347_n1744), .Y(u0__abc_49347_n1745) );
  OR2X2 OR2X2_3620 ( .A(u2_u4__abc_47660_n248), .B(u2_u4_b1_last_row_4_), .Y(u2_u4__abc_47660_n262) );
  OR2X2 OR2X2_3621 ( .A(u2_u4__abc_47660_n250), .B(row_adr_4_bF_buf5), .Y(u2_u4__abc_47660_n263) );
  OR2X2 OR2X2_3622 ( .A(u2_u4__abc_47660_n248), .B(u2_u4_b1_last_row_5_), .Y(u2_u4__abc_47660_n265) );
  OR2X2 OR2X2_3623 ( .A(u2_u4__abc_47660_n250), .B(row_adr_5_bF_buf5), .Y(u2_u4__abc_47660_n266) );
  OR2X2 OR2X2_3624 ( .A(u2_u4__abc_47660_n248), .B(u2_u4_b1_last_row_6_), .Y(u2_u4__abc_47660_n268) );
  OR2X2 OR2X2_3625 ( .A(u2_u4__abc_47660_n250), .B(row_adr_6_bF_buf5), .Y(u2_u4__abc_47660_n269) );
  OR2X2 OR2X2_3626 ( .A(u2_u4__abc_47660_n248), .B(u2_u4_b1_last_row_7_), .Y(u2_u4__abc_47660_n271) );
  OR2X2 OR2X2_3627 ( .A(u2_u4__abc_47660_n250), .B(row_adr_7_bF_buf5), .Y(u2_u4__abc_47660_n272) );
  OR2X2 OR2X2_3628 ( .A(u2_u4__abc_47660_n248), .B(u2_u4_b1_last_row_8_), .Y(u2_u4__abc_47660_n274) );
  OR2X2 OR2X2_3629 ( .A(u2_u4__abc_47660_n250), .B(row_adr_8_bF_buf5), .Y(u2_u4__abc_47660_n275_1) );
  OR2X2 OR2X2_363 ( .A(u0__abc_49347_n1746), .B(u0__abc_49347_n1747), .Y(u0__abc_49347_n1748) );
  OR2X2 OR2X2_3630 ( .A(u2_u4__abc_47660_n248), .B(u2_u4_b1_last_row_9_), .Y(u2_u4__abc_47660_n277) );
  OR2X2 OR2X2_3631 ( .A(u2_u4__abc_47660_n250), .B(row_adr_9_bF_buf5), .Y(u2_u4__abc_47660_n278_1) );
  OR2X2 OR2X2_3632 ( .A(u2_u4__abc_47660_n248), .B(u2_u4_b1_last_row_10_), .Y(u2_u4__abc_47660_n280) );
  OR2X2 OR2X2_3633 ( .A(u2_u4__abc_47660_n250), .B(row_adr_10_bF_buf5), .Y(u2_u4__abc_47660_n281) );
  OR2X2 OR2X2_3634 ( .A(u2_u4__abc_47660_n248), .B(u2_u4_b1_last_row_11_), .Y(u2_u4__abc_47660_n283_1) );
  OR2X2 OR2X2_3635 ( .A(u2_u4__abc_47660_n250), .B(row_adr_11_bF_buf5), .Y(u2_u4__abc_47660_n284) );
  OR2X2 OR2X2_3636 ( .A(u2_u4__abc_47660_n248), .B(u2_u4_b1_last_row_12_), .Y(u2_u4__abc_47660_n286_1) );
  OR2X2 OR2X2_3637 ( .A(u2_u4__abc_47660_n250), .B(row_adr_12_bF_buf5), .Y(u2_u4__abc_47660_n287_1) );
  OR2X2 OR2X2_3638 ( .A(u2_u4__abc_47660_n290_1), .B(u2_u4_b0_last_row_0_), .Y(u2_u4__abc_47660_n291) );
  OR2X2 OR2X2_3639 ( .A(u2_u4__abc_47660_n292_1), .B(row_adr_0_bF_buf4), .Y(u2_u4__abc_47660_n293) );
  OR2X2 OR2X2_364 ( .A(u0__abc_49347_n1749_1), .B(u0__abc_49347_n1750_1), .Y(u0__abc_49347_n1751_1) );
  OR2X2 OR2X2_3640 ( .A(u2_u4__abc_47660_n290_1), .B(u2_u4_b0_last_row_1_), .Y(u2_u4__abc_47660_n295) );
  OR2X2 OR2X2_3641 ( .A(u2_u4__abc_47660_n292_1), .B(row_adr_1_bF_buf4), .Y(u2_u4__abc_47660_n296_1) );
  OR2X2 OR2X2_3642 ( .A(u2_u4__abc_47660_n290_1), .B(u2_u4_b0_last_row_2_), .Y(u2_u4__abc_47660_n298) );
  OR2X2 OR2X2_3643 ( .A(u2_u4__abc_47660_n292_1), .B(row_adr_2_bF_buf4), .Y(u2_u4__abc_47660_n299) );
  OR2X2 OR2X2_3644 ( .A(u2_u4__abc_47660_n290_1), .B(u2_u4_b0_last_row_3_), .Y(u2_u4__abc_47660_n301) );
  OR2X2 OR2X2_3645 ( .A(u2_u4__abc_47660_n292_1), .B(row_adr_3_bF_buf4), .Y(u2_u4__abc_47660_n302) );
  OR2X2 OR2X2_3646 ( .A(u2_u4__abc_47660_n290_1), .B(u2_u4_b0_last_row_4_), .Y(u2_u4__abc_47660_n304_1) );
  OR2X2 OR2X2_3647 ( .A(u2_u4__abc_47660_n292_1), .B(row_adr_4_bF_buf4), .Y(u2_u4__abc_47660_n305_1) );
  OR2X2 OR2X2_3648 ( .A(u2_u4__abc_47660_n290_1), .B(u2_u4_b0_last_row_5_), .Y(u2_u4__abc_47660_n307) );
  OR2X2 OR2X2_3649 ( .A(u2_u4__abc_47660_n292_1), .B(row_adr_5_bF_buf4), .Y(u2_u4__abc_47660_n308) );
  OR2X2 OR2X2_365 ( .A(u0__abc_49347_n1753), .B(spec_req_cs_0_bF_buf3), .Y(u0__abc_49347_n1754_1) );
  OR2X2 OR2X2_3650 ( .A(u2_u4__abc_47660_n290_1), .B(u2_u4_b0_last_row_6_), .Y(u2_u4__abc_47660_n310) );
  OR2X2 OR2X2_3651 ( .A(u2_u4__abc_47660_n292_1), .B(row_adr_6_bF_buf4), .Y(u2_u4__abc_47660_n311) );
  OR2X2 OR2X2_3652 ( .A(u2_u4__abc_47660_n290_1), .B(u2_u4_b0_last_row_7_), .Y(u2_u4__abc_47660_n313) );
  OR2X2 OR2X2_3653 ( .A(u2_u4__abc_47660_n292_1), .B(row_adr_7_bF_buf4), .Y(u2_u4__abc_47660_n314) );
  OR2X2 OR2X2_3654 ( .A(u2_u4__abc_47660_n290_1), .B(u2_u4_b0_last_row_8_), .Y(u2_u4__abc_47660_n316) );
  OR2X2 OR2X2_3655 ( .A(u2_u4__abc_47660_n292_1), .B(row_adr_8_bF_buf4), .Y(u2_u4__abc_47660_n317) );
  OR2X2 OR2X2_3656 ( .A(u2_u4__abc_47660_n290_1), .B(u2_u4_b0_last_row_9_), .Y(u2_u4__abc_47660_n319) );
  OR2X2 OR2X2_3657 ( .A(u2_u4__abc_47660_n292_1), .B(row_adr_9_bF_buf4), .Y(u2_u4__abc_47660_n320) );
  OR2X2 OR2X2_3658 ( .A(u2_u4__abc_47660_n290_1), .B(u2_u4_b0_last_row_10_), .Y(u2_u4__abc_47660_n322) );
  OR2X2 OR2X2_3659 ( .A(u2_u4__abc_47660_n292_1), .B(row_adr_10_bF_buf4), .Y(u2_u4__abc_47660_n323) );
  OR2X2 OR2X2_366 ( .A(u0__abc_49347_n1752), .B(u0__abc_49347_n1754_1), .Y(u0__abc_49347_n1755) );
  OR2X2 OR2X2_3660 ( .A(u2_u4__abc_47660_n290_1), .B(u2_u4_b0_last_row_11_), .Y(u2_u4__abc_47660_n325) );
  OR2X2 OR2X2_3661 ( .A(u2_u4__abc_47660_n292_1), .B(row_adr_11_bF_buf4), .Y(u2_u4__abc_47660_n326) );
  OR2X2 OR2X2_3662 ( .A(u2_u4__abc_47660_n290_1), .B(u2_u4_b0_last_row_12_), .Y(u2_u4__abc_47660_n328) );
  OR2X2 OR2X2_3663 ( .A(u2_u4__abc_47660_n292_1), .B(row_adr_12_bF_buf4), .Y(u2_u4__abc_47660_n329) );
  OR2X2 OR2X2_3664 ( .A(u2_u4__abc_47660_n331), .B(row_adr_12_bF_buf3), .Y(u2_u4__abc_47660_n332) );
  OR2X2 OR2X2_3665 ( .A(u2_u4__abc_47660_n333), .B(row_adr_11_bF_buf3), .Y(u2_u4__abc_47660_n334) );
  OR2X2 OR2X2_3666 ( .A(u2_u4__abc_47660_n199), .B(u2_u4_b0_last_row_12_), .Y(u2_u4__abc_47660_n335) );
  OR2X2 OR2X2_3667 ( .A(u2_u4__abc_47660_n194), .B(u2_u4_b0_last_row_11_), .Y(u2_u4__abc_47660_n338) );
  OR2X2 OR2X2_3668 ( .A(u2_u4__abc_47660_n339), .B(row_adr_9_bF_buf3), .Y(u2_u4__abc_47660_n340) );
  OR2X2 OR2X2_3669 ( .A(u2_u4__abc_47660_n184), .B(u2_u4_b0_last_row_9_), .Y(u2_u4__abc_47660_n342) );
  OR2X2 OR2X2_367 ( .A(u0__abc_49347_n1203_bF_buf0), .B(u0_tms0_23_), .Y(u0__abc_49347_n1756_1) );
  OR2X2 OR2X2_3670 ( .A(u2_u4__abc_47660_n343), .B(row_adr_7_bF_buf3), .Y(u2_u4__abc_47660_n344) );
  OR2X2 OR2X2_3671 ( .A(u2_u4__abc_47660_n164), .B(u2_u4_b0_last_row_5_), .Y(u2_u4__abc_47660_n348) );
  OR2X2 OR2X2_3672 ( .A(u2_u4__abc_47660_n159), .B(u2_u4_b0_last_row_4_), .Y(u2_u4__abc_47660_n350) );
  OR2X2 OR2X2_3673 ( .A(u2_u4__abc_47660_n351), .B(row_adr_4_bF_buf3), .Y(u2_u4__abc_47660_n352) );
  OR2X2 OR2X2_3674 ( .A(u2_u4__abc_47660_n355), .B(row_adr_0_bF_buf3), .Y(u2_u4__abc_47660_n356) );
  OR2X2 OR2X2_3675 ( .A(u2_u4__abc_47660_n139), .B(u2_u4_b0_last_row_0_), .Y(u2_u4__abc_47660_n357) );
  OR2X2 OR2X2_3676 ( .A(u2_u4__abc_47660_n144), .B(u2_u4_b0_last_row_1_), .Y(u2_u4__abc_47660_n359) );
  OR2X2 OR2X2_3677 ( .A(u2_u4__abc_47660_n360), .B(row_adr_5_bF_buf3), .Y(u2_u4__abc_47660_n361) );
  OR2X2 OR2X2_3678 ( .A(u2_u4__abc_47660_n366), .B(row_adr_10_bF_buf3), .Y(u2_u4__abc_47660_n367) );
  OR2X2 OR2X2_3679 ( .A(u2_u4__abc_47660_n189), .B(u2_u4_b0_last_row_10_), .Y(u2_u4__abc_47660_n368) );
  OR2X2 OR2X2_368 ( .A(u0__abc_49347_n1758), .B(u0__abc_49347_n1736), .Y(u0_sp_tms_23__FF_INPUT) );
  OR2X2 OR2X2_3680 ( .A(u2_u4__abc_47660_n372), .B(u2_u4__abc_47660_n370), .Y(u2_u4__abc_47660_n373) );
  OR2X2 OR2X2_3681 ( .A(u2_u4__abc_47660_n154), .B(u2_u4_b0_last_row_3_), .Y(u2_u4__abc_47660_n375) );
  OR2X2 OR2X2_3682 ( .A(u2_u4__abc_47660_n376), .B(row_adr_2_bF_buf3), .Y(u2_u4__abc_47660_n377) );
  OR2X2 OR2X2_3683 ( .A(u2_u4__abc_47660_n379), .B(row_adr_1_bF_buf3), .Y(u2_u4__abc_47660_n380) );
  OR2X2 OR2X2_3684 ( .A(u2_u4__abc_47660_n149), .B(u2_u4_b0_last_row_2_), .Y(u2_u4__abc_47660_n381) );
  OR2X2 OR2X2_3685 ( .A(u2_u4__abc_47660_n384), .B(row_adr_3_bF_buf3), .Y(u2_u4__abc_47660_n385) );
  OR2X2 OR2X2_3686 ( .A(u2_u4__abc_47660_n174), .B(u2_u4_b0_last_row_7_), .Y(u2_u4__abc_47660_n386) );
  OR2X2 OR2X2_3687 ( .A(u2_u4__abc_47660_n390), .B(u2_u4__abc_47660_n388), .Y(u2_u4__abc_47660_n391) );
  OR2X2 OR2X2_3688 ( .A(u2_u4__abc_47660_n396), .B(row_adr_12_bF_buf2), .Y(u2_u4__abc_47660_n397) );
  OR2X2 OR2X2_3689 ( .A(u2_u4__abc_47660_n398), .B(row_adr_11_bF_buf2), .Y(u2_u4__abc_47660_n399) );
  OR2X2 OR2X2_369 ( .A(u0__abc_49347_n1183_1_bF_buf5), .B(1'b0), .Y(u0__abc_49347_n1762) );
  OR2X2 OR2X2_3690 ( .A(u2_u4__abc_47660_n199), .B(u2_u4_b2_last_row_12_), .Y(u2_u4__abc_47660_n400) );
  OR2X2 OR2X2_3691 ( .A(u2_u4__abc_47660_n194), .B(u2_u4_b2_last_row_11_), .Y(u2_u4__abc_47660_n403) );
  OR2X2 OR2X2_3692 ( .A(u2_u4__abc_47660_n404), .B(row_adr_9_bF_buf2), .Y(u2_u4__abc_47660_n405) );
  OR2X2 OR2X2_3693 ( .A(u2_u4__abc_47660_n184), .B(u2_u4_b2_last_row_9_), .Y(u2_u4__abc_47660_n407) );
  OR2X2 OR2X2_3694 ( .A(u2_u4__abc_47660_n408), .B(row_adr_7_bF_buf2), .Y(u2_u4__abc_47660_n409) );
  OR2X2 OR2X2_3695 ( .A(u2_u4__abc_47660_n164), .B(u2_u4_b2_last_row_5_), .Y(u2_u4__abc_47660_n413) );
  OR2X2 OR2X2_3696 ( .A(u2_u4__abc_47660_n159), .B(u2_u4_b2_last_row_4_), .Y(u2_u4__abc_47660_n415) );
  OR2X2 OR2X2_3697 ( .A(u2_u4__abc_47660_n416), .B(row_adr_4_bF_buf2), .Y(u2_u4__abc_47660_n417) );
  OR2X2 OR2X2_3698 ( .A(u2_u4__abc_47660_n420), .B(row_adr_0_bF_buf2), .Y(u2_u4__abc_47660_n421) );
  OR2X2 OR2X2_3699 ( .A(u2_u4__abc_47660_n139), .B(u2_u4_b2_last_row_0_), .Y(u2_u4__abc_47660_n422) );
  OR2X2 OR2X2_37 ( .A(_abc_55805_n240_bF_buf2), .B(sp_tms_1_), .Y(_abc_55805_n293) );
  OR2X2 OR2X2_370 ( .A(spec_req_cs_6_bF_buf2), .B(1'b0), .Y(u0__abc_49347_n1763_1) );
  OR2X2 OR2X2_3700 ( .A(u2_u4__abc_47660_n144), .B(u2_u4_b2_last_row_1_), .Y(u2_u4__abc_47660_n424) );
  OR2X2 OR2X2_3701 ( .A(u2_u4__abc_47660_n425), .B(row_adr_5_bF_buf2), .Y(u2_u4__abc_47660_n426) );
  OR2X2 OR2X2_3702 ( .A(u2_u4__abc_47660_n431), .B(row_adr_10_bF_buf2), .Y(u2_u4__abc_47660_n432) );
  OR2X2 OR2X2_3703 ( .A(u2_u4__abc_47660_n189), .B(u2_u4_b2_last_row_10_), .Y(u2_u4__abc_47660_n433) );
  OR2X2 OR2X2_3704 ( .A(u2_u4__abc_47660_n437), .B(u2_u4__abc_47660_n435), .Y(u2_u4__abc_47660_n438) );
  OR2X2 OR2X2_3705 ( .A(u2_u4__abc_47660_n154), .B(u2_u4_b2_last_row_3_), .Y(u2_u4__abc_47660_n440) );
  OR2X2 OR2X2_3706 ( .A(u2_u4__abc_47660_n441), .B(row_adr_2_bF_buf2), .Y(u2_u4__abc_47660_n442) );
  OR2X2 OR2X2_3707 ( .A(u2_u4__abc_47660_n444), .B(row_adr_1_bF_buf2), .Y(u2_u4__abc_47660_n445) );
  OR2X2 OR2X2_3708 ( .A(u2_u4__abc_47660_n149), .B(u2_u4_b2_last_row_2_), .Y(u2_u4__abc_47660_n446) );
  OR2X2 OR2X2_3709 ( .A(u2_u4__abc_47660_n449), .B(row_adr_3_bF_buf2), .Y(u2_u4__abc_47660_n450) );
  OR2X2 OR2X2_371 ( .A(u0__abc_49347_n1765), .B(u0__abc_49347_n1761), .Y(u0__abc_49347_n1766_1) );
  OR2X2 OR2X2_3710 ( .A(u2_u4__abc_47660_n174), .B(u2_u4_b2_last_row_7_), .Y(u2_u4__abc_47660_n451) );
  OR2X2 OR2X2_3711 ( .A(u2_u4__abc_47660_n455), .B(u2_u4__abc_47660_n453), .Y(u2_u4__abc_47660_n456) );
  OR2X2 OR2X2_3712 ( .A(u2_u4__abc_47660_n395), .B(u2_u4__abc_47660_n460), .Y(u2_u4__abc_47660_n461) );
  OR2X2 OR2X2_3713 ( .A(u2_u4__abc_47660_n462), .B(row_adr_12_bF_buf1), .Y(u2_u4__abc_47660_n463) );
  OR2X2 OR2X2_3714 ( .A(u2_u4__abc_47660_n464), .B(row_adr_11_bF_buf1), .Y(u2_u4__abc_47660_n465) );
  OR2X2 OR2X2_3715 ( .A(u2_u4__abc_47660_n199), .B(u2_u4_b1_last_row_12_), .Y(u2_u4__abc_47660_n466) );
  OR2X2 OR2X2_3716 ( .A(u2_u4__abc_47660_n194), .B(u2_u4_b1_last_row_11_), .Y(u2_u4__abc_47660_n469) );
  OR2X2 OR2X2_3717 ( .A(u2_u4__abc_47660_n470), .B(row_adr_9_bF_buf1), .Y(u2_u4__abc_47660_n471) );
  OR2X2 OR2X2_3718 ( .A(u2_u4__abc_47660_n184), .B(u2_u4_b1_last_row_9_), .Y(u2_u4__abc_47660_n473) );
  OR2X2 OR2X2_3719 ( .A(u2_u4__abc_47660_n474), .B(row_adr_7_bF_buf1), .Y(u2_u4__abc_47660_n475) );
  OR2X2 OR2X2_372 ( .A(u0__abc_49347_n1767_1), .B(u0__abc_49347_n1768), .Y(u0__abc_49347_n1769) );
  OR2X2 OR2X2_3720 ( .A(u2_u4__abc_47660_n164), .B(u2_u4_b1_last_row_5_), .Y(u2_u4__abc_47660_n479) );
  OR2X2 OR2X2_3721 ( .A(u2_u4__abc_47660_n159), .B(u2_u4_b1_last_row_4_), .Y(u2_u4__abc_47660_n481) );
  OR2X2 OR2X2_3722 ( .A(u2_u4__abc_47660_n482), .B(row_adr_4_bF_buf1), .Y(u2_u4__abc_47660_n483) );
  OR2X2 OR2X2_3723 ( .A(u2_u4__abc_47660_n486), .B(row_adr_0_bF_buf1), .Y(u2_u4__abc_47660_n487) );
  OR2X2 OR2X2_3724 ( .A(u2_u4__abc_47660_n139), .B(u2_u4_b1_last_row_0_), .Y(u2_u4__abc_47660_n488) );
  OR2X2 OR2X2_3725 ( .A(u2_u4__abc_47660_n144), .B(u2_u4_b1_last_row_1_), .Y(u2_u4__abc_47660_n490) );
  OR2X2 OR2X2_3726 ( .A(u2_u4__abc_47660_n491), .B(row_adr_5_bF_buf1), .Y(u2_u4__abc_47660_n492) );
  OR2X2 OR2X2_3727 ( .A(u2_u4__abc_47660_n497), .B(row_adr_10_bF_buf1), .Y(u2_u4__abc_47660_n498) );
  OR2X2 OR2X2_3728 ( .A(u2_u4__abc_47660_n189), .B(u2_u4_b1_last_row_10_), .Y(u2_u4__abc_47660_n499) );
  OR2X2 OR2X2_3729 ( .A(u2_u4__abc_47660_n503), .B(u2_u4__abc_47660_n501), .Y(u2_u4__abc_47660_n504) );
  OR2X2 OR2X2_373 ( .A(u0__abc_49347_n1770), .B(u0__abc_49347_n1771_1), .Y(u0__abc_49347_n1772_1) );
  OR2X2 OR2X2_3730 ( .A(u2_u4__abc_47660_n154), .B(u2_u4_b1_last_row_3_), .Y(u2_u4__abc_47660_n506) );
  OR2X2 OR2X2_3731 ( .A(u2_u4__abc_47660_n507), .B(row_adr_2_bF_buf1), .Y(u2_u4__abc_47660_n508) );
  OR2X2 OR2X2_3732 ( .A(u2_u4__abc_47660_n510), .B(row_adr_1_bF_buf1), .Y(u2_u4__abc_47660_n511) );
  OR2X2 OR2X2_3733 ( .A(u2_u4__abc_47660_n149), .B(u2_u4_b1_last_row_2_), .Y(u2_u4__abc_47660_n512) );
  OR2X2 OR2X2_3734 ( .A(u2_u4__abc_47660_n515), .B(row_adr_3_bF_buf1), .Y(u2_u4__abc_47660_n516) );
  OR2X2 OR2X2_3735 ( .A(u2_u4__abc_47660_n174), .B(u2_u4_b1_last_row_7_), .Y(u2_u4__abc_47660_n517) );
  OR2X2 OR2X2_3736 ( .A(u2_u4__abc_47660_n521), .B(u2_u4__abc_47660_n519), .Y(u2_u4__abc_47660_n522) );
  OR2X2 OR2X2_3737 ( .A(u2_u4__abc_47660_n527), .B(row_adr_9_bF_buf0), .Y(u2_u4__abc_47660_n528) );
  OR2X2 OR2X2_3738 ( .A(u2_u4__abc_47660_n189), .B(u2_u4_b3_last_row_10_), .Y(u2_u4__abc_47660_n529) );
  OR2X2 OR2X2_3739 ( .A(u2_u4__abc_47660_n184), .B(u2_u4_b3_last_row_9_), .Y(u2_u4__abc_47660_n530) );
  OR2X2 OR2X2_374 ( .A(u0__abc_49347_n1773_1), .B(u0__abc_49347_n1774_1), .Y(u0__abc_49347_n1775_1) );
  OR2X2 OR2X2_3740 ( .A(u2_u4__abc_47660_n194), .B(u2_u4_b3_last_row_11_), .Y(u2_u4__abc_47660_n533) );
  OR2X2 OR2X2_3741 ( .A(u2_u4__abc_47660_n534), .B(row_adr_11_bF_buf0), .Y(u2_u4__abc_47660_n535) );
  OR2X2 OR2X2_3742 ( .A(u2_u4__abc_47660_n199), .B(u2_u4_b3_last_row_12_), .Y(u2_u4__abc_47660_n537) );
  OR2X2 OR2X2_3743 ( .A(u2_u4__abc_47660_n538), .B(row_adr_8_bF_buf0), .Y(u2_u4__abc_47660_n539) );
  OR2X2 OR2X2_3744 ( .A(u2_u4__abc_47660_n159), .B(u2_u4_b3_last_row_4_), .Y(u2_u4__abc_47660_n543) );
  OR2X2 OR2X2_3745 ( .A(u2_u4__abc_47660_n544), .B(row_adr_4_bF_buf0), .Y(u2_u4__abc_47660_n545) );
  OR2X2 OR2X2_3746 ( .A(u2_u4__abc_47660_n547), .B(row_adr_3_bF_buf0), .Y(u2_u4__abc_47660_n548) );
  OR2X2 OR2X2_3747 ( .A(u2_u4__abc_47660_n551), .B(row_adr_0_bF_buf0), .Y(u2_u4__abc_47660_n552) );
  OR2X2 OR2X2_3748 ( .A(u2_u4__abc_47660_n139), .B(u2_u4_b3_last_row_0_), .Y(u2_u4__abc_47660_n553) );
  OR2X2 OR2X2_3749 ( .A(u2_u4__abc_47660_n555), .B(row_adr_2_bF_buf0), .Y(u2_u4__abc_47660_n556) );
  OR2X2 OR2X2_375 ( .A(u0__abc_49347_n1777_1), .B(spec_req_cs_0_bF_buf2), .Y(u0__abc_49347_n1778_1) );
  OR2X2 OR2X2_3750 ( .A(u2_u4__abc_47660_n149), .B(u2_u4_b3_last_row_2_), .Y(u2_u4__abc_47660_n557) );
  OR2X2 OR2X2_3751 ( .A(u2_u4__abc_47660_n174), .B(u2_u4_b3_last_row_7_), .Y(u2_u4__abc_47660_n562) );
  OR2X2 OR2X2_3752 ( .A(u2_u4__abc_47660_n563), .B(row_adr_7_bF_buf0), .Y(u2_u4__abc_47660_n564) );
  OR2X2 OR2X2_3753 ( .A(u2_u4__abc_47660_n566), .B(row_adr_10_bF_buf0), .Y(u2_u4__abc_47660_n567) );
  OR2X2 OR2X2_3754 ( .A(u2_u4__abc_47660_n179), .B(u2_u4_b3_last_row_8_), .Y(u2_u4__abc_47660_n568) );
  OR2X2 OR2X2_3755 ( .A(u2_u4__abc_47660_n169), .B(u2_u4_b3_last_row_6_), .Y(u2_u4__abc_47660_n571) );
  OR2X2 OR2X2_3756 ( .A(u2_u4__abc_47660_n572), .B(row_adr_6_bF_buf0), .Y(u2_u4__abc_47660_n573) );
  OR2X2 OR2X2_3757 ( .A(u2_u4__abc_47660_n575), .B(row_adr_5_bF_buf0), .Y(u2_u4__abc_47660_n576) );
  OR2X2 OR2X2_3758 ( .A(u2_u4__abc_47660_n154), .B(u2_u4_b3_last_row_3_), .Y(u2_u4__abc_47660_n577) );
  OR2X2 OR2X2_3759 ( .A(u2_u4__abc_47660_n164), .B(u2_u4_b3_last_row_5_), .Y(u2_u4__abc_47660_n580) );
  OR2X2 OR2X2_376 ( .A(u0__abc_49347_n1776_1), .B(u0__abc_49347_n1778_1), .Y(u0__abc_49347_n1779_1) );
  OR2X2 OR2X2_3760 ( .A(u2_u4__abc_47660_n581), .B(row_adr_1_bF_buf0), .Y(u2_u4__abc_47660_n582) );
  OR2X2 OR2X2_3761 ( .A(u2_u4__abc_47660_n144), .B(u2_u4_b3_last_row_1_), .Y(u2_u4__abc_47660_n584) );
  OR2X2 OR2X2_3762 ( .A(u2_u4__abc_47660_n585), .B(row_adr_12_bF_buf0), .Y(u2_u4__abc_47660_n586) );
  OR2X2 OR2X2_3763 ( .A(u2_u4__abc_47660_n526), .B(u2_u4__abc_47660_n591), .Y(u2_u4__abc_47660_n592) );
  OR2X2 OR2X2_3764 ( .A(u2_u4__abc_47660_n461), .B(u2_u4__abc_47660_n592), .Y(u2_row_same_4) );
  OR2X2 OR2X2_3765 ( .A(u2_u4__abc_47660_n594), .B(u2_u4__abc_47660_n595), .Y(u2_u4__abc_47660_n596) );
  OR2X2 OR2X2_3766 ( .A(u2_u4__abc_47660_n598), .B(u2_u4__abc_47660_n597), .Y(u2_u4__abc_47660_n599) );
  OR2X2 OR2X2_3767 ( .A(u2_u4__abc_47660_n596), .B(u2_u4__abc_47660_n599), .Y(u2_bank_open_4) );
  OR2X2 OR2X2_3768 ( .A(u2_u4__abc_47660_n608), .B(u2_u4__abc_47660_n137_bF_buf3), .Y(u2_u4_bank3_open_FF_INPUT) );
  OR2X2 OR2X2_3769 ( .A(u2_u4__abc_47660_n611), .B(u2_u4__abc_47660_n610), .Y(u2_u4__abc_47660_n612) );
  OR2X2 OR2X2_377 ( .A(u0__abc_49347_n1203_bF_buf5), .B(u0_tms0_24_), .Y(u0__abc_49347_n1780_1) );
  OR2X2 OR2X2_3770 ( .A(u2_u4__abc_47660_n614), .B(u2_u4__abc_47660_n205), .Y(u2_u4_bank2_open_FF_INPUT) );
  OR2X2 OR2X2_3771 ( .A(u2_u4__abc_47660_n616), .B(u2_u4__abc_47660_n610), .Y(u2_u4__abc_47660_n617) );
  OR2X2 OR2X2_3772 ( .A(u2_u4__abc_47660_n619), .B(u2_u4__abc_47660_n248), .Y(u2_u4_bank1_open_FF_INPUT) );
  OR2X2 OR2X2_3773 ( .A(u2_u4__abc_47660_n621), .B(u2_u4__abc_47660_n610), .Y(u2_u4__abc_47660_n622) );
  OR2X2 OR2X2_3774 ( .A(u2_u4__abc_47660_n624), .B(u2_u4__abc_47660_n290_1), .Y(u2_u4_bank0_open_FF_INPUT) );
  OR2X2 OR2X2_3775 ( .A(u2_u5__abc_47660_n137_bF_buf4), .B(u2_u5_b3_last_row_0_), .Y(u2_u5__abc_47660_n138) );
  OR2X2 OR2X2_3776 ( .A(u2_u5__abc_47660_n137_bF_buf2), .B(u2_u5_b3_last_row_1_), .Y(u2_u5__abc_47660_n143) );
  OR2X2 OR2X2_3777 ( .A(u2_u5__abc_47660_n137_bF_buf0), .B(u2_u5_b3_last_row_2_), .Y(u2_u5__abc_47660_n148) );
  OR2X2 OR2X2_3778 ( .A(u2_u5__abc_47660_n137_bF_buf3), .B(u2_u5_b3_last_row_3_), .Y(u2_u5__abc_47660_n153) );
  OR2X2 OR2X2_3779 ( .A(u2_u5__abc_47660_n137_bF_buf1), .B(u2_u5_b3_last_row_4_), .Y(u2_u5__abc_47660_n158) );
  OR2X2 OR2X2_378 ( .A(u0__abc_49347_n1782_1), .B(u0__abc_49347_n1760_1), .Y(u0_sp_tms_24__FF_INPUT) );
  OR2X2 OR2X2_3780 ( .A(u2_u5__abc_47660_n137_bF_buf4), .B(u2_u5_b3_last_row_5_), .Y(u2_u5__abc_47660_n163) );
  OR2X2 OR2X2_3781 ( .A(u2_u5__abc_47660_n137_bF_buf2), .B(u2_u5_b3_last_row_6_), .Y(u2_u5__abc_47660_n168) );
  OR2X2 OR2X2_3782 ( .A(u2_u5__abc_47660_n137_bF_buf0), .B(u2_u5_b3_last_row_7_), .Y(u2_u5__abc_47660_n173) );
  OR2X2 OR2X2_3783 ( .A(u2_u5__abc_47660_n137_bF_buf3), .B(u2_u5_b3_last_row_8_), .Y(u2_u5__abc_47660_n178) );
  OR2X2 OR2X2_3784 ( .A(u2_u5__abc_47660_n137_bF_buf1), .B(u2_u5_b3_last_row_9_), .Y(u2_u5__abc_47660_n183) );
  OR2X2 OR2X2_3785 ( .A(u2_u5__abc_47660_n137_bF_buf4), .B(u2_u5_b3_last_row_10_), .Y(u2_u5__abc_47660_n188) );
  OR2X2 OR2X2_3786 ( .A(u2_u5__abc_47660_n137_bF_buf2), .B(u2_u5_b3_last_row_11_), .Y(u2_u5__abc_47660_n193) );
  OR2X2 OR2X2_3787 ( .A(u2_u5__abc_47660_n137_bF_buf0), .B(u2_u5_b3_last_row_12_), .Y(u2_u5__abc_47660_n198) );
  OR2X2 OR2X2_3788 ( .A(u2_u5__abc_47660_n205), .B(u2_u5_b2_last_row_0_), .Y(u2_u5__abc_47660_n206) );
  OR2X2 OR2X2_3789 ( .A(u2_u5__abc_47660_n207), .B(row_adr_0_bF_buf5), .Y(u2_u5__abc_47660_n208) );
  OR2X2 OR2X2_379 ( .A(u0__abc_49347_n1183_1_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n1786_1) );
  OR2X2 OR2X2_3790 ( .A(u2_u5__abc_47660_n205), .B(u2_u5_b2_last_row_1_), .Y(u2_u5__abc_47660_n210) );
  OR2X2 OR2X2_3791 ( .A(u2_u5__abc_47660_n207), .B(row_adr_1_bF_buf5), .Y(u2_u5__abc_47660_n211) );
  OR2X2 OR2X2_3792 ( .A(u2_u5__abc_47660_n205), .B(u2_u5_b2_last_row_2_), .Y(u2_u5__abc_47660_n213) );
  OR2X2 OR2X2_3793 ( .A(u2_u5__abc_47660_n207), .B(row_adr_2_bF_buf5), .Y(u2_u5__abc_47660_n214) );
  OR2X2 OR2X2_3794 ( .A(u2_u5__abc_47660_n205), .B(u2_u5_b2_last_row_3_), .Y(u2_u5__abc_47660_n216) );
  OR2X2 OR2X2_3795 ( .A(u2_u5__abc_47660_n207), .B(row_adr_3_bF_buf5), .Y(u2_u5__abc_47660_n217) );
  OR2X2 OR2X2_3796 ( .A(u2_u5__abc_47660_n205), .B(u2_u5_b2_last_row_4_), .Y(u2_u5__abc_47660_n219) );
  OR2X2 OR2X2_3797 ( .A(u2_u5__abc_47660_n207), .B(row_adr_4_bF_buf5), .Y(u2_u5__abc_47660_n220) );
  OR2X2 OR2X2_3798 ( .A(u2_u5__abc_47660_n205), .B(u2_u5_b2_last_row_5_), .Y(u2_u5__abc_47660_n222) );
  OR2X2 OR2X2_3799 ( .A(u2_u5__abc_47660_n207), .B(row_adr_5_bF_buf5), .Y(u2_u5__abc_47660_n223) );
  OR2X2 OR2X2_38 ( .A(lmr_sel_bF_buf4), .B(tms_1_), .Y(_abc_55805_n294) );
  OR2X2 OR2X2_380 ( .A(spec_req_cs_6_bF_buf1), .B(1'b0), .Y(u0__abc_49347_n1787_1) );
  OR2X2 OR2X2_3800 ( .A(u2_u5__abc_47660_n205), .B(u2_u5_b2_last_row_6_), .Y(u2_u5__abc_47660_n225) );
  OR2X2 OR2X2_3801 ( .A(u2_u5__abc_47660_n207), .B(row_adr_6_bF_buf5), .Y(u2_u5__abc_47660_n226) );
  OR2X2 OR2X2_3802 ( .A(u2_u5__abc_47660_n205), .B(u2_u5_b2_last_row_7_), .Y(u2_u5__abc_47660_n228) );
  OR2X2 OR2X2_3803 ( .A(u2_u5__abc_47660_n207), .B(row_adr_7_bF_buf5), .Y(u2_u5__abc_47660_n229) );
  OR2X2 OR2X2_3804 ( .A(u2_u5__abc_47660_n205), .B(u2_u5_b2_last_row_8_), .Y(u2_u5__abc_47660_n231) );
  OR2X2 OR2X2_3805 ( .A(u2_u5__abc_47660_n207), .B(row_adr_8_bF_buf5), .Y(u2_u5__abc_47660_n232) );
  OR2X2 OR2X2_3806 ( .A(u2_u5__abc_47660_n205), .B(u2_u5_b2_last_row_9_), .Y(u2_u5__abc_47660_n234) );
  OR2X2 OR2X2_3807 ( .A(u2_u5__abc_47660_n207), .B(row_adr_9_bF_buf5), .Y(u2_u5__abc_47660_n235) );
  OR2X2 OR2X2_3808 ( .A(u2_u5__abc_47660_n205), .B(u2_u5_b2_last_row_10_), .Y(u2_u5__abc_47660_n237) );
  OR2X2 OR2X2_3809 ( .A(u2_u5__abc_47660_n207), .B(row_adr_10_bF_buf5), .Y(u2_u5__abc_47660_n238) );
  OR2X2 OR2X2_381 ( .A(u0__abc_49347_n1789_1), .B(u0__abc_49347_n1785_1), .Y(u0__abc_49347_n1790_1) );
  OR2X2 OR2X2_3810 ( .A(u2_u5__abc_47660_n205), .B(u2_u5_b2_last_row_11_), .Y(u2_u5__abc_47660_n240) );
  OR2X2 OR2X2_3811 ( .A(u2_u5__abc_47660_n207), .B(row_adr_11_bF_buf5), .Y(u2_u5__abc_47660_n241) );
  OR2X2 OR2X2_3812 ( .A(u2_u5__abc_47660_n205), .B(u2_u5_b2_last_row_12_), .Y(u2_u5__abc_47660_n243) );
  OR2X2 OR2X2_3813 ( .A(u2_u5__abc_47660_n207), .B(row_adr_12_bF_buf5), .Y(u2_u5__abc_47660_n244) );
  OR2X2 OR2X2_3814 ( .A(u2_u5__abc_47660_n248), .B(u2_u5_b1_last_row_0_), .Y(u2_u5__abc_47660_n249) );
  OR2X2 OR2X2_3815 ( .A(u2_u5__abc_47660_n250), .B(row_adr_0_bF_buf4), .Y(u2_u5__abc_47660_n251) );
  OR2X2 OR2X2_3816 ( .A(u2_u5__abc_47660_n248), .B(u2_u5_b1_last_row_1_), .Y(u2_u5__abc_47660_n253) );
  OR2X2 OR2X2_3817 ( .A(u2_u5__abc_47660_n250), .B(row_adr_1_bF_buf4), .Y(u2_u5__abc_47660_n254) );
  OR2X2 OR2X2_3818 ( .A(u2_u5__abc_47660_n248), .B(u2_u5_b1_last_row_2_), .Y(u2_u5__abc_47660_n256) );
  OR2X2 OR2X2_3819 ( .A(u2_u5__abc_47660_n250), .B(row_adr_2_bF_buf4), .Y(u2_u5__abc_47660_n257) );
  OR2X2 OR2X2_382 ( .A(u0__abc_49347_n1791_1), .B(u0__abc_49347_n1792_1), .Y(u0__abc_49347_n1793_1) );
  OR2X2 OR2X2_3820 ( .A(u2_u5__abc_47660_n248), .B(u2_u5_b1_last_row_3_), .Y(u2_u5__abc_47660_n259) );
  OR2X2 OR2X2_3821 ( .A(u2_u5__abc_47660_n250), .B(row_adr_3_bF_buf4), .Y(u2_u5__abc_47660_n260) );
  OR2X2 OR2X2_3822 ( .A(u2_u5__abc_47660_n248), .B(u2_u5_b1_last_row_4_), .Y(u2_u5__abc_47660_n262) );
  OR2X2 OR2X2_3823 ( .A(u2_u5__abc_47660_n250), .B(row_adr_4_bF_buf4), .Y(u2_u5__abc_47660_n263) );
  OR2X2 OR2X2_3824 ( .A(u2_u5__abc_47660_n248), .B(u2_u5_b1_last_row_5_), .Y(u2_u5__abc_47660_n265) );
  OR2X2 OR2X2_3825 ( .A(u2_u5__abc_47660_n250), .B(row_adr_5_bF_buf4), .Y(u2_u5__abc_47660_n266) );
  OR2X2 OR2X2_3826 ( .A(u2_u5__abc_47660_n248), .B(u2_u5_b1_last_row_6_), .Y(u2_u5__abc_47660_n268) );
  OR2X2 OR2X2_3827 ( .A(u2_u5__abc_47660_n250), .B(row_adr_6_bF_buf4), .Y(u2_u5__abc_47660_n269) );
  OR2X2 OR2X2_3828 ( .A(u2_u5__abc_47660_n248), .B(u2_u5_b1_last_row_7_), .Y(u2_u5__abc_47660_n271) );
  OR2X2 OR2X2_3829 ( .A(u2_u5__abc_47660_n250), .B(row_adr_7_bF_buf4), .Y(u2_u5__abc_47660_n272) );
  OR2X2 OR2X2_383 ( .A(u0__abc_49347_n1794_1), .B(u0__abc_49347_n1795_1), .Y(u0__abc_49347_n1796_1) );
  OR2X2 OR2X2_3830 ( .A(u2_u5__abc_47660_n248), .B(u2_u5_b1_last_row_8_), .Y(u2_u5__abc_47660_n274) );
  OR2X2 OR2X2_3831 ( .A(u2_u5__abc_47660_n250), .B(row_adr_8_bF_buf4), .Y(u2_u5__abc_47660_n275_1) );
  OR2X2 OR2X2_3832 ( .A(u2_u5__abc_47660_n248), .B(u2_u5_b1_last_row_9_), .Y(u2_u5__abc_47660_n277) );
  OR2X2 OR2X2_3833 ( .A(u2_u5__abc_47660_n250), .B(row_adr_9_bF_buf4), .Y(u2_u5__abc_47660_n278_1) );
  OR2X2 OR2X2_3834 ( .A(u2_u5__abc_47660_n248), .B(u2_u5_b1_last_row_10_), .Y(u2_u5__abc_47660_n280) );
  OR2X2 OR2X2_3835 ( .A(u2_u5__abc_47660_n250), .B(row_adr_10_bF_buf4), .Y(u2_u5__abc_47660_n281) );
  OR2X2 OR2X2_3836 ( .A(u2_u5__abc_47660_n248), .B(u2_u5_b1_last_row_11_), .Y(u2_u5__abc_47660_n283_1) );
  OR2X2 OR2X2_3837 ( .A(u2_u5__abc_47660_n250), .B(row_adr_11_bF_buf4), .Y(u2_u5__abc_47660_n284) );
  OR2X2 OR2X2_3838 ( .A(u2_u5__abc_47660_n248), .B(u2_u5_b1_last_row_12_), .Y(u2_u5__abc_47660_n286_1) );
  OR2X2 OR2X2_3839 ( .A(u2_u5__abc_47660_n250), .B(row_adr_12_bF_buf4), .Y(u2_u5__abc_47660_n287_1) );
  OR2X2 OR2X2_384 ( .A(u0__abc_49347_n1797_1), .B(u0__abc_49347_n1798_1), .Y(u0__abc_49347_n1799_1) );
  OR2X2 OR2X2_3840 ( .A(u2_u5__abc_47660_n290_1), .B(u2_u5_b0_last_row_0_), .Y(u2_u5__abc_47660_n291) );
  OR2X2 OR2X2_3841 ( .A(u2_u5__abc_47660_n292_1), .B(row_adr_0_bF_buf3), .Y(u2_u5__abc_47660_n293) );
  OR2X2 OR2X2_3842 ( .A(u2_u5__abc_47660_n290_1), .B(u2_u5_b0_last_row_1_), .Y(u2_u5__abc_47660_n295) );
  OR2X2 OR2X2_3843 ( .A(u2_u5__abc_47660_n292_1), .B(row_adr_1_bF_buf3), .Y(u2_u5__abc_47660_n296_1) );
  OR2X2 OR2X2_3844 ( .A(u2_u5__abc_47660_n290_1), .B(u2_u5_b0_last_row_2_), .Y(u2_u5__abc_47660_n298) );
  OR2X2 OR2X2_3845 ( .A(u2_u5__abc_47660_n292_1), .B(row_adr_2_bF_buf3), .Y(u2_u5__abc_47660_n299) );
  OR2X2 OR2X2_3846 ( .A(u2_u5__abc_47660_n290_1), .B(u2_u5_b0_last_row_3_), .Y(u2_u5__abc_47660_n301) );
  OR2X2 OR2X2_3847 ( .A(u2_u5__abc_47660_n292_1), .B(row_adr_3_bF_buf3), .Y(u2_u5__abc_47660_n302) );
  OR2X2 OR2X2_3848 ( .A(u2_u5__abc_47660_n290_1), .B(u2_u5_b0_last_row_4_), .Y(u2_u5__abc_47660_n304_1) );
  OR2X2 OR2X2_3849 ( .A(u2_u5__abc_47660_n292_1), .B(row_adr_4_bF_buf3), .Y(u2_u5__abc_47660_n305_1) );
  OR2X2 OR2X2_385 ( .A(u0__abc_49347_n1801_1), .B(spec_req_cs_0_bF_buf1), .Y(u0__abc_49347_n1802_1) );
  OR2X2 OR2X2_3850 ( .A(u2_u5__abc_47660_n290_1), .B(u2_u5_b0_last_row_5_), .Y(u2_u5__abc_47660_n307) );
  OR2X2 OR2X2_3851 ( .A(u2_u5__abc_47660_n292_1), .B(row_adr_5_bF_buf3), .Y(u2_u5__abc_47660_n308) );
  OR2X2 OR2X2_3852 ( .A(u2_u5__abc_47660_n290_1), .B(u2_u5_b0_last_row_6_), .Y(u2_u5__abc_47660_n310) );
  OR2X2 OR2X2_3853 ( .A(u2_u5__abc_47660_n292_1), .B(row_adr_6_bF_buf3), .Y(u2_u5__abc_47660_n311) );
  OR2X2 OR2X2_3854 ( .A(u2_u5__abc_47660_n290_1), .B(u2_u5_b0_last_row_7_), .Y(u2_u5__abc_47660_n313) );
  OR2X2 OR2X2_3855 ( .A(u2_u5__abc_47660_n292_1), .B(row_adr_7_bF_buf3), .Y(u2_u5__abc_47660_n314) );
  OR2X2 OR2X2_3856 ( .A(u2_u5__abc_47660_n290_1), .B(u2_u5_b0_last_row_8_), .Y(u2_u5__abc_47660_n316) );
  OR2X2 OR2X2_3857 ( .A(u2_u5__abc_47660_n292_1), .B(row_adr_8_bF_buf3), .Y(u2_u5__abc_47660_n317) );
  OR2X2 OR2X2_3858 ( .A(u2_u5__abc_47660_n290_1), .B(u2_u5_b0_last_row_9_), .Y(u2_u5__abc_47660_n319) );
  OR2X2 OR2X2_3859 ( .A(u2_u5__abc_47660_n292_1), .B(row_adr_9_bF_buf3), .Y(u2_u5__abc_47660_n320) );
  OR2X2 OR2X2_386 ( .A(u0__abc_49347_n1800_1), .B(u0__abc_49347_n1802_1), .Y(u0__abc_49347_n1803_1) );
  OR2X2 OR2X2_3860 ( .A(u2_u5__abc_47660_n290_1), .B(u2_u5_b0_last_row_10_), .Y(u2_u5__abc_47660_n322) );
  OR2X2 OR2X2_3861 ( .A(u2_u5__abc_47660_n292_1), .B(row_adr_10_bF_buf3), .Y(u2_u5__abc_47660_n323) );
  OR2X2 OR2X2_3862 ( .A(u2_u5__abc_47660_n290_1), .B(u2_u5_b0_last_row_11_), .Y(u2_u5__abc_47660_n325) );
  OR2X2 OR2X2_3863 ( .A(u2_u5__abc_47660_n292_1), .B(row_adr_11_bF_buf3), .Y(u2_u5__abc_47660_n326) );
  OR2X2 OR2X2_3864 ( .A(u2_u5__abc_47660_n290_1), .B(u2_u5_b0_last_row_12_), .Y(u2_u5__abc_47660_n328) );
  OR2X2 OR2X2_3865 ( .A(u2_u5__abc_47660_n292_1), .B(row_adr_12_bF_buf3), .Y(u2_u5__abc_47660_n329) );
  OR2X2 OR2X2_3866 ( .A(u2_u5__abc_47660_n331), .B(row_adr_12_bF_buf2), .Y(u2_u5__abc_47660_n332) );
  OR2X2 OR2X2_3867 ( .A(u2_u5__abc_47660_n333), .B(row_adr_11_bF_buf2), .Y(u2_u5__abc_47660_n334) );
  OR2X2 OR2X2_3868 ( .A(u2_u5__abc_47660_n199), .B(u2_u5_b0_last_row_12_), .Y(u2_u5__abc_47660_n335) );
  OR2X2 OR2X2_3869 ( .A(u2_u5__abc_47660_n194), .B(u2_u5_b0_last_row_11_), .Y(u2_u5__abc_47660_n338) );
  OR2X2 OR2X2_387 ( .A(u0__abc_49347_n1203_bF_buf4), .B(u0_tms0_25_), .Y(u0__abc_49347_n1804_1) );
  OR2X2 OR2X2_3870 ( .A(u2_u5__abc_47660_n339), .B(row_adr_9_bF_buf2), .Y(u2_u5__abc_47660_n340) );
  OR2X2 OR2X2_3871 ( .A(u2_u5__abc_47660_n184), .B(u2_u5_b0_last_row_9_), .Y(u2_u5__abc_47660_n342) );
  OR2X2 OR2X2_3872 ( .A(u2_u5__abc_47660_n343), .B(row_adr_7_bF_buf2), .Y(u2_u5__abc_47660_n344) );
  OR2X2 OR2X2_3873 ( .A(u2_u5__abc_47660_n164), .B(u2_u5_b0_last_row_5_), .Y(u2_u5__abc_47660_n348) );
  OR2X2 OR2X2_3874 ( .A(u2_u5__abc_47660_n159), .B(u2_u5_b0_last_row_4_), .Y(u2_u5__abc_47660_n350) );
  OR2X2 OR2X2_3875 ( .A(u2_u5__abc_47660_n351), .B(row_adr_4_bF_buf2), .Y(u2_u5__abc_47660_n352) );
  OR2X2 OR2X2_3876 ( .A(u2_u5__abc_47660_n355), .B(row_adr_0_bF_buf2), .Y(u2_u5__abc_47660_n356) );
  OR2X2 OR2X2_3877 ( .A(u2_u5__abc_47660_n139), .B(u2_u5_b0_last_row_0_), .Y(u2_u5__abc_47660_n357) );
  OR2X2 OR2X2_3878 ( .A(u2_u5__abc_47660_n144), .B(u2_u5_b0_last_row_1_), .Y(u2_u5__abc_47660_n359) );
  OR2X2 OR2X2_3879 ( .A(u2_u5__abc_47660_n360), .B(row_adr_5_bF_buf2), .Y(u2_u5__abc_47660_n361) );
  OR2X2 OR2X2_388 ( .A(u0__abc_49347_n1806_1), .B(u0__abc_49347_n1784_1), .Y(u0_sp_tms_25__FF_INPUT) );
  OR2X2 OR2X2_3880 ( .A(u2_u5__abc_47660_n366), .B(row_adr_10_bF_buf2), .Y(u2_u5__abc_47660_n367) );
  OR2X2 OR2X2_3881 ( .A(u2_u5__abc_47660_n189), .B(u2_u5_b0_last_row_10_), .Y(u2_u5__abc_47660_n368) );
  OR2X2 OR2X2_3882 ( .A(u2_u5__abc_47660_n372), .B(u2_u5__abc_47660_n370), .Y(u2_u5__abc_47660_n373) );
  OR2X2 OR2X2_3883 ( .A(u2_u5__abc_47660_n154), .B(u2_u5_b0_last_row_3_), .Y(u2_u5__abc_47660_n375) );
  OR2X2 OR2X2_3884 ( .A(u2_u5__abc_47660_n376), .B(row_adr_2_bF_buf2), .Y(u2_u5__abc_47660_n377) );
  OR2X2 OR2X2_3885 ( .A(u2_u5__abc_47660_n379), .B(row_adr_1_bF_buf2), .Y(u2_u5__abc_47660_n380) );
  OR2X2 OR2X2_3886 ( .A(u2_u5__abc_47660_n149), .B(u2_u5_b0_last_row_2_), .Y(u2_u5__abc_47660_n381) );
  OR2X2 OR2X2_3887 ( .A(u2_u5__abc_47660_n384), .B(row_adr_3_bF_buf2), .Y(u2_u5__abc_47660_n385) );
  OR2X2 OR2X2_3888 ( .A(u2_u5__abc_47660_n174), .B(u2_u5_b0_last_row_7_), .Y(u2_u5__abc_47660_n386) );
  OR2X2 OR2X2_3889 ( .A(u2_u5__abc_47660_n390), .B(u2_u5__abc_47660_n388), .Y(u2_u5__abc_47660_n391) );
  OR2X2 OR2X2_389 ( .A(u0__abc_49347_n1183_1_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n1810_1) );
  OR2X2 OR2X2_3890 ( .A(u2_u5__abc_47660_n396), .B(row_adr_12_bF_buf1), .Y(u2_u5__abc_47660_n397) );
  OR2X2 OR2X2_3891 ( .A(u2_u5__abc_47660_n398), .B(row_adr_11_bF_buf1), .Y(u2_u5__abc_47660_n399) );
  OR2X2 OR2X2_3892 ( .A(u2_u5__abc_47660_n199), .B(u2_u5_b2_last_row_12_), .Y(u2_u5__abc_47660_n400) );
  OR2X2 OR2X2_3893 ( .A(u2_u5__abc_47660_n194), .B(u2_u5_b2_last_row_11_), .Y(u2_u5__abc_47660_n403) );
  OR2X2 OR2X2_3894 ( .A(u2_u5__abc_47660_n404), .B(row_adr_9_bF_buf1), .Y(u2_u5__abc_47660_n405) );
  OR2X2 OR2X2_3895 ( .A(u2_u5__abc_47660_n184), .B(u2_u5_b2_last_row_9_), .Y(u2_u5__abc_47660_n407) );
  OR2X2 OR2X2_3896 ( .A(u2_u5__abc_47660_n408), .B(row_adr_7_bF_buf1), .Y(u2_u5__abc_47660_n409) );
  OR2X2 OR2X2_3897 ( .A(u2_u5__abc_47660_n164), .B(u2_u5_b2_last_row_5_), .Y(u2_u5__abc_47660_n413) );
  OR2X2 OR2X2_3898 ( .A(u2_u5__abc_47660_n159), .B(u2_u5_b2_last_row_4_), .Y(u2_u5__abc_47660_n415) );
  OR2X2 OR2X2_3899 ( .A(u2_u5__abc_47660_n416), .B(row_adr_4_bF_buf1), .Y(u2_u5__abc_47660_n417) );
  OR2X2 OR2X2_39 ( .A(_abc_55805_n240_bF_buf1), .B(sp_tms_2_), .Y(_abc_55805_n296) );
  OR2X2 OR2X2_390 ( .A(spec_req_cs_6_bF_buf0), .B(1'b0), .Y(u0__abc_49347_n1811_1) );
  OR2X2 OR2X2_3900 ( .A(u2_u5__abc_47660_n420), .B(row_adr_0_bF_buf1), .Y(u2_u5__abc_47660_n421) );
  OR2X2 OR2X2_3901 ( .A(u2_u5__abc_47660_n139), .B(u2_u5_b2_last_row_0_), .Y(u2_u5__abc_47660_n422) );
  OR2X2 OR2X2_3902 ( .A(u2_u5__abc_47660_n144), .B(u2_u5_b2_last_row_1_), .Y(u2_u5__abc_47660_n424) );
  OR2X2 OR2X2_3903 ( .A(u2_u5__abc_47660_n425), .B(row_adr_5_bF_buf1), .Y(u2_u5__abc_47660_n426) );
  OR2X2 OR2X2_3904 ( .A(u2_u5__abc_47660_n431), .B(row_adr_10_bF_buf1), .Y(u2_u5__abc_47660_n432) );
  OR2X2 OR2X2_3905 ( .A(u2_u5__abc_47660_n189), .B(u2_u5_b2_last_row_10_), .Y(u2_u5__abc_47660_n433) );
  OR2X2 OR2X2_3906 ( .A(u2_u5__abc_47660_n437), .B(u2_u5__abc_47660_n435), .Y(u2_u5__abc_47660_n438) );
  OR2X2 OR2X2_3907 ( .A(u2_u5__abc_47660_n154), .B(u2_u5_b2_last_row_3_), .Y(u2_u5__abc_47660_n440) );
  OR2X2 OR2X2_3908 ( .A(u2_u5__abc_47660_n441), .B(row_adr_2_bF_buf1), .Y(u2_u5__abc_47660_n442) );
  OR2X2 OR2X2_3909 ( .A(u2_u5__abc_47660_n444), .B(row_adr_1_bF_buf1), .Y(u2_u5__abc_47660_n445) );
  OR2X2 OR2X2_391 ( .A(u0__abc_49347_n1813_1), .B(u0__abc_49347_n1809_1), .Y(u0__abc_49347_n1814_1) );
  OR2X2 OR2X2_3910 ( .A(u2_u5__abc_47660_n149), .B(u2_u5_b2_last_row_2_), .Y(u2_u5__abc_47660_n446) );
  OR2X2 OR2X2_3911 ( .A(u2_u5__abc_47660_n449), .B(row_adr_3_bF_buf1), .Y(u2_u5__abc_47660_n450) );
  OR2X2 OR2X2_3912 ( .A(u2_u5__abc_47660_n174), .B(u2_u5_b2_last_row_7_), .Y(u2_u5__abc_47660_n451) );
  OR2X2 OR2X2_3913 ( .A(u2_u5__abc_47660_n455), .B(u2_u5__abc_47660_n453), .Y(u2_u5__abc_47660_n456) );
  OR2X2 OR2X2_3914 ( .A(u2_u5__abc_47660_n395), .B(u2_u5__abc_47660_n460), .Y(u2_u5__abc_47660_n461) );
  OR2X2 OR2X2_3915 ( .A(u2_u5__abc_47660_n462), .B(row_adr_12_bF_buf0), .Y(u2_u5__abc_47660_n463) );
  OR2X2 OR2X2_3916 ( .A(u2_u5__abc_47660_n464), .B(row_adr_11_bF_buf0), .Y(u2_u5__abc_47660_n465) );
  OR2X2 OR2X2_3917 ( .A(u2_u5__abc_47660_n199), .B(u2_u5_b1_last_row_12_), .Y(u2_u5__abc_47660_n466) );
  OR2X2 OR2X2_3918 ( .A(u2_u5__abc_47660_n194), .B(u2_u5_b1_last_row_11_), .Y(u2_u5__abc_47660_n469) );
  OR2X2 OR2X2_3919 ( .A(u2_u5__abc_47660_n470), .B(row_adr_9_bF_buf0), .Y(u2_u5__abc_47660_n471) );
  OR2X2 OR2X2_392 ( .A(u0__abc_49347_n1815_1), .B(u0__abc_49347_n1816_1), .Y(u0__abc_49347_n1817_1) );
  OR2X2 OR2X2_3920 ( .A(u2_u5__abc_47660_n184), .B(u2_u5_b1_last_row_9_), .Y(u2_u5__abc_47660_n473) );
  OR2X2 OR2X2_3921 ( .A(u2_u5__abc_47660_n474), .B(row_adr_7_bF_buf0), .Y(u2_u5__abc_47660_n475) );
  OR2X2 OR2X2_3922 ( .A(u2_u5__abc_47660_n164), .B(u2_u5_b1_last_row_5_), .Y(u2_u5__abc_47660_n479) );
  OR2X2 OR2X2_3923 ( .A(u2_u5__abc_47660_n159), .B(u2_u5_b1_last_row_4_), .Y(u2_u5__abc_47660_n481) );
  OR2X2 OR2X2_3924 ( .A(u2_u5__abc_47660_n482), .B(row_adr_4_bF_buf0), .Y(u2_u5__abc_47660_n483) );
  OR2X2 OR2X2_3925 ( .A(u2_u5__abc_47660_n486), .B(row_adr_0_bF_buf0), .Y(u2_u5__abc_47660_n487) );
  OR2X2 OR2X2_3926 ( .A(u2_u5__abc_47660_n139), .B(u2_u5_b1_last_row_0_), .Y(u2_u5__abc_47660_n488) );
  OR2X2 OR2X2_3927 ( .A(u2_u5__abc_47660_n144), .B(u2_u5_b1_last_row_1_), .Y(u2_u5__abc_47660_n490) );
  OR2X2 OR2X2_3928 ( .A(u2_u5__abc_47660_n491), .B(row_adr_5_bF_buf0), .Y(u2_u5__abc_47660_n492) );
  OR2X2 OR2X2_3929 ( .A(u2_u5__abc_47660_n497), .B(row_adr_10_bF_buf0), .Y(u2_u5__abc_47660_n498) );
  OR2X2 OR2X2_393 ( .A(u0__abc_49347_n1818_1), .B(u0__abc_49347_n1819_1), .Y(u0__abc_49347_n1820_1) );
  OR2X2 OR2X2_3930 ( .A(u2_u5__abc_47660_n189), .B(u2_u5_b1_last_row_10_), .Y(u2_u5__abc_47660_n499) );
  OR2X2 OR2X2_3931 ( .A(u2_u5__abc_47660_n503), .B(u2_u5__abc_47660_n501), .Y(u2_u5__abc_47660_n504) );
  OR2X2 OR2X2_3932 ( .A(u2_u5__abc_47660_n154), .B(u2_u5_b1_last_row_3_), .Y(u2_u5__abc_47660_n506) );
  OR2X2 OR2X2_3933 ( .A(u2_u5__abc_47660_n507), .B(row_adr_2_bF_buf0), .Y(u2_u5__abc_47660_n508) );
  OR2X2 OR2X2_3934 ( .A(u2_u5__abc_47660_n510), .B(row_adr_1_bF_buf0), .Y(u2_u5__abc_47660_n511) );
  OR2X2 OR2X2_3935 ( .A(u2_u5__abc_47660_n149), .B(u2_u5_b1_last_row_2_), .Y(u2_u5__abc_47660_n512) );
  OR2X2 OR2X2_3936 ( .A(u2_u5__abc_47660_n515), .B(row_adr_3_bF_buf0), .Y(u2_u5__abc_47660_n516) );
  OR2X2 OR2X2_3937 ( .A(u2_u5__abc_47660_n174), .B(u2_u5_b1_last_row_7_), .Y(u2_u5__abc_47660_n517) );
  OR2X2 OR2X2_3938 ( .A(u2_u5__abc_47660_n521), .B(u2_u5__abc_47660_n519), .Y(u2_u5__abc_47660_n522) );
  OR2X2 OR2X2_3939 ( .A(u2_u5__abc_47660_n527), .B(row_adr_9_bF_buf6), .Y(u2_u5__abc_47660_n528) );
  OR2X2 OR2X2_394 ( .A(u0__abc_49347_n1821_1), .B(u0__abc_49347_n1822_1), .Y(u0__abc_49347_n1823_1) );
  OR2X2 OR2X2_3940 ( .A(u2_u5__abc_47660_n189), .B(u2_u5_b3_last_row_10_), .Y(u2_u5__abc_47660_n529) );
  OR2X2 OR2X2_3941 ( .A(u2_u5__abc_47660_n184), .B(u2_u5_b3_last_row_9_), .Y(u2_u5__abc_47660_n530) );
  OR2X2 OR2X2_3942 ( .A(u2_u5__abc_47660_n194), .B(u2_u5_b3_last_row_11_), .Y(u2_u5__abc_47660_n533) );
  OR2X2 OR2X2_3943 ( .A(u2_u5__abc_47660_n534), .B(row_adr_11_bF_buf6), .Y(u2_u5__abc_47660_n535) );
  OR2X2 OR2X2_3944 ( .A(u2_u5__abc_47660_n199), .B(u2_u5_b3_last_row_12_), .Y(u2_u5__abc_47660_n537) );
  OR2X2 OR2X2_3945 ( .A(u2_u5__abc_47660_n538), .B(row_adr_8_bF_buf6), .Y(u2_u5__abc_47660_n539) );
  OR2X2 OR2X2_3946 ( .A(u2_u5__abc_47660_n159), .B(u2_u5_b3_last_row_4_), .Y(u2_u5__abc_47660_n543) );
  OR2X2 OR2X2_3947 ( .A(u2_u5__abc_47660_n544), .B(row_adr_4_bF_buf6), .Y(u2_u5__abc_47660_n545) );
  OR2X2 OR2X2_3948 ( .A(u2_u5__abc_47660_n547), .B(row_adr_3_bF_buf6), .Y(u2_u5__abc_47660_n548) );
  OR2X2 OR2X2_3949 ( .A(u2_u5__abc_47660_n551), .B(row_adr_0_bF_buf6), .Y(u2_u5__abc_47660_n552) );
  OR2X2 OR2X2_395 ( .A(u0__abc_49347_n1825_1), .B(spec_req_cs_0_bF_buf0), .Y(u0__abc_49347_n1826_1) );
  OR2X2 OR2X2_3950 ( .A(u2_u5__abc_47660_n139), .B(u2_u5_b3_last_row_0_), .Y(u2_u5__abc_47660_n553) );
  OR2X2 OR2X2_3951 ( .A(u2_u5__abc_47660_n555), .B(row_adr_2_bF_buf6), .Y(u2_u5__abc_47660_n556) );
  OR2X2 OR2X2_3952 ( .A(u2_u5__abc_47660_n149), .B(u2_u5_b3_last_row_2_), .Y(u2_u5__abc_47660_n557) );
  OR2X2 OR2X2_3953 ( .A(u2_u5__abc_47660_n174), .B(u2_u5_b3_last_row_7_), .Y(u2_u5__abc_47660_n562) );
  OR2X2 OR2X2_3954 ( .A(u2_u5__abc_47660_n563), .B(row_adr_7_bF_buf6), .Y(u2_u5__abc_47660_n564) );
  OR2X2 OR2X2_3955 ( .A(u2_u5__abc_47660_n566), .B(row_adr_10_bF_buf6), .Y(u2_u5__abc_47660_n567) );
  OR2X2 OR2X2_3956 ( .A(u2_u5__abc_47660_n179), .B(u2_u5_b3_last_row_8_), .Y(u2_u5__abc_47660_n568) );
  OR2X2 OR2X2_3957 ( .A(u2_u5__abc_47660_n169), .B(u2_u5_b3_last_row_6_), .Y(u2_u5__abc_47660_n571) );
  OR2X2 OR2X2_3958 ( .A(u2_u5__abc_47660_n572), .B(row_adr_6_bF_buf6), .Y(u2_u5__abc_47660_n573) );
  OR2X2 OR2X2_3959 ( .A(u2_u5__abc_47660_n575), .B(row_adr_5_bF_buf6), .Y(u2_u5__abc_47660_n576) );
  OR2X2 OR2X2_396 ( .A(u0__abc_49347_n1824_1), .B(u0__abc_49347_n1826_1), .Y(u0__abc_49347_n1827_1) );
  OR2X2 OR2X2_3960 ( .A(u2_u5__abc_47660_n154), .B(u2_u5_b3_last_row_3_), .Y(u2_u5__abc_47660_n577) );
  OR2X2 OR2X2_3961 ( .A(u2_u5__abc_47660_n164), .B(u2_u5_b3_last_row_5_), .Y(u2_u5__abc_47660_n580) );
  OR2X2 OR2X2_3962 ( .A(u2_u5__abc_47660_n581), .B(row_adr_1_bF_buf6), .Y(u2_u5__abc_47660_n582) );
  OR2X2 OR2X2_3963 ( .A(u2_u5__abc_47660_n144), .B(u2_u5_b3_last_row_1_), .Y(u2_u5__abc_47660_n584) );
  OR2X2 OR2X2_3964 ( .A(u2_u5__abc_47660_n585), .B(row_adr_12_bF_buf6), .Y(u2_u5__abc_47660_n586) );
  OR2X2 OR2X2_3965 ( .A(u2_u5__abc_47660_n526), .B(u2_u5__abc_47660_n591), .Y(u2_u5__abc_47660_n592) );
  OR2X2 OR2X2_3966 ( .A(u2_u5__abc_47660_n461), .B(u2_u5__abc_47660_n592), .Y(u2_row_same_5) );
  OR2X2 OR2X2_3967 ( .A(u2_u5__abc_47660_n594), .B(u2_u5__abc_47660_n595), .Y(u2_u5__abc_47660_n596) );
  OR2X2 OR2X2_3968 ( .A(u2_u5__abc_47660_n598), .B(u2_u5__abc_47660_n597), .Y(u2_u5__abc_47660_n599) );
  OR2X2 OR2X2_3969 ( .A(u2_u5__abc_47660_n596), .B(u2_u5__abc_47660_n599), .Y(u2_bank_open_5) );
  OR2X2 OR2X2_397 ( .A(u0__abc_49347_n1203_bF_buf3), .B(u0_tms0_26_), .Y(u0__abc_49347_n1828_1) );
  OR2X2 OR2X2_3970 ( .A(u2_u5__abc_47660_n608), .B(u2_u5__abc_47660_n137_bF_buf3), .Y(u2_u5_bank3_open_FF_INPUT) );
  OR2X2 OR2X2_3971 ( .A(u2_u5__abc_47660_n611), .B(u2_u5__abc_47660_n610), .Y(u2_u5__abc_47660_n612) );
  OR2X2 OR2X2_3972 ( .A(u2_u5__abc_47660_n614), .B(u2_u5__abc_47660_n205), .Y(u2_u5_bank2_open_FF_INPUT) );
  OR2X2 OR2X2_3973 ( .A(u2_u5__abc_47660_n616), .B(u2_u5__abc_47660_n610), .Y(u2_u5__abc_47660_n617) );
  OR2X2 OR2X2_3974 ( .A(u2_u5__abc_47660_n619), .B(u2_u5__abc_47660_n248), .Y(u2_u5_bank1_open_FF_INPUT) );
  OR2X2 OR2X2_3975 ( .A(u2_u5__abc_47660_n621), .B(u2_u5__abc_47660_n610), .Y(u2_u5__abc_47660_n622) );
  OR2X2 OR2X2_3976 ( .A(u2_u5__abc_47660_n624), .B(u2_u5__abc_47660_n290_1), .Y(u2_u5_bank0_open_FF_INPUT) );
  OR2X2 OR2X2_3977 ( .A(csc_3_), .B(csc_2_), .Y(u3__abc_46775_n275) );
  OR2X2 OR2X2_3978 ( .A(mem_ack_r), .B(csc_1_), .Y(u3__abc_46775_n276) );
  OR2X2 OR2X2_3979 ( .A(u3__abc_46775_n275_bF_buf4), .B(u3__abc_46775_n276), .Y(u3__abc_46775_n277_1) );
  OR2X2 OR2X2_398 ( .A(u0__abc_49347_n1830_1), .B(u0__abc_49347_n1808_1), .Y(u0_sp_tms_26__FF_INPUT) );
  OR2X2 OR2X2_3980 ( .A(u3__abc_46775_n277_1_bF_buf5), .B(mc_dp_od_0_), .Y(u3__abc_46775_n278_1) );
  OR2X2 OR2X2_3981 ( .A(\wb_data_i[3] ), .B(\wb_data_i[2] ), .Y(u3__abc_46775_n280) );
  OR2X2 OR2X2_3982 ( .A(u3__abc_46775_n285_1), .B(\wb_data_i[0] ), .Y(u3__abc_46775_n286_1) );
  OR2X2 OR2X2_3983 ( .A(u3__abc_46775_n287_1), .B(\wb_data_i[1] ), .Y(u3__abc_46775_n288) );
  OR2X2 OR2X2_3984 ( .A(u3__abc_46775_n284), .B(u3__abc_46775_n289), .Y(u3__abc_46775_n292_1) );
  OR2X2 OR2X2_3985 ( .A(\wb_data_i[7] ), .B(\wb_data_i[6] ), .Y(u3__abc_46775_n295_1) );
  OR2X2 OR2X2_3986 ( .A(u3__abc_46775_n300_1), .B(\wb_data_i[4] ), .Y(u3__abc_46775_n301_1) );
  OR2X2 OR2X2_3987 ( .A(u3__abc_46775_n302_1), .B(\wb_data_i[5] ), .Y(u3__abc_46775_n303) );
  OR2X2 OR2X2_3988 ( .A(u3__abc_46775_n306_1), .B(u3__abc_46775_n307_1), .Y(u3__abc_46775_n308) );
  OR2X2 OR2X2_3989 ( .A(u3__abc_46775_n294), .B(u3__abc_46775_n309), .Y(u3__abc_46775_n310_1) );
  OR2X2 OR2X2_399 ( .A(u0__abc_49347_n1183_1_bF_buf2), .B(1'b0), .Y(u0__abc_49347_n1834_1) );
  OR2X2 OR2X2_3990 ( .A(u3__abc_46775_n293), .B(u3__abc_46775_n308), .Y(u3__abc_46775_n311_1) );
  OR2X2 OR2X2_3991 ( .A(u3__abc_46775_n312_1), .B(u3__abc_46775_n279_bF_buf5), .Y(u3__abc_46775_n313) );
  OR2X2 OR2X2_3992 ( .A(u3__abc_46775_n277_1_bF_buf3), .B(mc_dp_od_1_), .Y(u3__abc_46775_n315_1) );
  OR2X2 OR2X2_3993 ( .A(\wb_data_i[11] ), .B(\wb_data_i[10] ), .Y(u3__abc_46775_n316_1) );
  OR2X2 OR2X2_3994 ( .A(u3__abc_46775_n320_1), .B(\wb_data_i[8] ), .Y(u3__abc_46775_n321_1) );
  OR2X2 OR2X2_3995 ( .A(u3__abc_46775_n322_1), .B(\wb_data_i[9] ), .Y(u3__abc_46775_n323) );
  OR2X2 OR2X2_3996 ( .A(u3__abc_46775_n325_1), .B(u3__abc_46775_n319), .Y(u3__abc_46775_n328) );
  OR2X2 OR2X2_3997 ( .A(\wb_data_i[15] ), .B(\wb_data_i[14] ), .Y(u3__abc_46775_n331_1) );
  OR2X2 OR2X2_3998 ( .A(u3__abc_46775_n336_1), .B(\wb_data_i[12] ), .Y(u3__abc_46775_n337_1) );
  OR2X2 OR2X2_3999 ( .A(u3__abc_46775_n338), .B(\wb_data_i[13] ), .Y(u3__abc_46775_n339) );
  OR2X2 OR2X2_4 ( .A(lmr_sel_bF_buf6), .B(cs_0_), .Y(_abc_55805_n242_1) );
  OR2X2 OR2X2_40 ( .A(lmr_sel_bF_buf3), .B(tms_2_), .Y(_abc_55805_n297) );
  OR2X2 OR2X2_400 ( .A(spec_req_cs_6_bF_buf5), .B(1'b0), .Y(u0__abc_49347_n1835_1) );
  OR2X2 OR2X2_4000 ( .A(u3__abc_46775_n342_1), .B(u3__abc_46775_n343), .Y(u3__abc_46775_n344) );
  OR2X2 OR2X2_4001 ( .A(u3__abc_46775_n330_1), .B(u3__abc_46775_n345_1), .Y(u3__abc_46775_n346_1) );
  OR2X2 OR2X2_4002 ( .A(u3__abc_46775_n329), .B(u3__abc_46775_n344), .Y(u3__abc_46775_n347_1) );
  OR2X2 OR2X2_4003 ( .A(u3__abc_46775_n348), .B(u3__abc_46775_n279_bF_buf4), .Y(u3__abc_46775_n349) );
  OR2X2 OR2X2_4004 ( .A(\wb_data_i[19] ), .B(\wb_data_i[18] ), .Y(u3__abc_46775_n351_1) );
  OR2X2 OR2X2_4005 ( .A(u3__abc_46775_n355_1), .B(\wb_data_i[16] ), .Y(u3__abc_46775_n356_1) );
  OR2X2 OR2X2_4006 ( .A(u3__abc_46775_n357_1), .B(\wb_data_i[17] ), .Y(u3__abc_46775_n358) );
  OR2X2 OR2X2_4007 ( .A(u3__abc_46775_n360_1), .B(u3__abc_46775_n354), .Y(u3__abc_46775_n363) );
  OR2X2 OR2X2_4008 ( .A(\wb_data_i[23] ), .B(\wb_data_i[22] ), .Y(u3__abc_46775_n365_1) );
  OR2X2 OR2X2_4009 ( .A(u3__abc_46775_n370_1), .B(\wb_data_i[20] ), .Y(u3__abc_46775_n371_1) );
  OR2X2 OR2X2_401 ( .A(u0__abc_49347_n1837_1), .B(u0__abc_49347_n1833_1), .Y(u0__abc_49347_n1838_1) );
  OR2X2 OR2X2_4010 ( .A(u3__abc_46775_n372_1), .B(\wb_data_i[21] ), .Y(u3__abc_46775_n373_1) );
  OR2X2 OR2X2_4011 ( .A(u3__abc_46775_n376), .B(u3__abc_46775_n377), .Y(u3__abc_46775_n378) );
  OR2X2 OR2X2_4012 ( .A(u3__abc_46775_n382), .B(u3__abc_46775_n380), .Y(u3__abc_46775_n383) );
  OR2X2 OR2X2_4013 ( .A(u3__abc_46775_n384), .B(u3__abc_46775_n385), .Y(u3_mc_dp_o_2__FF_INPUT) );
  OR2X2 OR2X2_4014 ( .A(\wb_data_i[27] ), .B(\wb_data_i[26] ), .Y(u3__abc_46775_n387) );
  OR2X2 OR2X2_4015 ( .A(u3__abc_46775_n391), .B(\wb_data_i[24] ), .Y(u3__abc_46775_n392_1) );
  OR2X2 OR2X2_4016 ( .A(u3__abc_46775_n393_1), .B(\wb_data_i[25] ), .Y(u3__abc_46775_n394) );
  OR2X2 OR2X2_4017 ( .A(u3__abc_46775_n396), .B(u3__abc_46775_n390_1), .Y(u3__abc_46775_n399) );
  OR2X2 OR2X2_4018 ( .A(\wb_data_i[31] ), .B(\wb_data_i[30] ), .Y(u3__abc_46775_n401) );
  OR2X2 OR2X2_4019 ( .A(u3__abc_46775_n406), .B(\wb_data_i[28] ), .Y(u3__abc_46775_n407) );
  OR2X2 OR2X2_402 ( .A(u0__abc_49347_n1839_1), .B(u0__abc_49347_n1840_1), .Y(u0__abc_49347_n1841_1) );
  OR2X2 OR2X2_4020 ( .A(u3__abc_46775_n408), .B(\wb_data_i[29] ), .Y(u3__abc_46775_n409) );
  OR2X2 OR2X2_4021 ( .A(u3__abc_46775_n412), .B(u3__abc_46775_n413_1), .Y(u3__abc_46775_n414_1) );
  OR2X2 OR2X2_4022 ( .A(u3__abc_46775_n418), .B(u3__abc_46775_n416_1), .Y(u3__abc_46775_n419_1) );
  OR2X2 OR2X2_4023 ( .A(u3__abc_46775_n420), .B(u3__abc_46775_n421_1), .Y(u3_mc_dp_o_3__FF_INPUT) );
  OR2X2 OR2X2_4024 ( .A(u3_byte2_0_), .B(pack_le2), .Y(u3__abc_46775_n423) );
  OR2X2 OR2X2_4025 ( .A(u3__abc_46775_n424), .B(mc_data_ir_0_), .Y(u3__abc_46775_n425) );
  OR2X2 OR2X2_4026 ( .A(pack_le2), .B(u3_byte2_1_), .Y(u3__abc_46775_n427) );
  OR2X2 OR2X2_4027 ( .A(u3__abc_46775_n424), .B(mc_data_ir_1_), .Y(u3__abc_46775_n428) );
  OR2X2 OR2X2_4028 ( .A(pack_le2), .B(u3_byte2_2_), .Y(u3__abc_46775_n430) );
  OR2X2 OR2X2_4029 ( .A(u3__abc_46775_n424), .B(mc_data_ir_2_), .Y(u3__abc_46775_n431) );
  OR2X2 OR2X2_403 ( .A(u0__abc_49347_n1842_1), .B(u0__abc_49347_n1843_1), .Y(u0__abc_49347_n1844_1) );
  OR2X2 OR2X2_4030 ( .A(pack_le2), .B(u3_byte2_3_), .Y(u3__abc_46775_n433) );
  OR2X2 OR2X2_4031 ( .A(u3__abc_46775_n424), .B(mc_data_ir_3_), .Y(u3__abc_46775_n434) );
  OR2X2 OR2X2_4032 ( .A(pack_le2), .B(u3_byte2_4_), .Y(u3__abc_46775_n436) );
  OR2X2 OR2X2_4033 ( .A(u3__abc_46775_n424), .B(mc_data_ir_4_), .Y(u3__abc_46775_n437) );
  OR2X2 OR2X2_4034 ( .A(pack_le2), .B(u3_byte2_5_), .Y(u3__abc_46775_n439) );
  OR2X2 OR2X2_4035 ( .A(u3__abc_46775_n424), .B(mc_data_ir_5_), .Y(u3__abc_46775_n440) );
  OR2X2 OR2X2_4036 ( .A(pack_le2), .B(u3_byte2_6_), .Y(u3__abc_46775_n442) );
  OR2X2 OR2X2_4037 ( .A(u3__abc_46775_n424), .B(mc_data_ir_6_), .Y(u3__abc_46775_n443) );
  OR2X2 OR2X2_4038 ( .A(pack_le2), .B(u3_byte2_7_), .Y(u3__abc_46775_n445) );
  OR2X2 OR2X2_4039 ( .A(u3__abc_46775_n424), .B(mc_data_ir_7_), .Y(u3__abc_46775_n446) );
  OR2X2 OR2X2_404 ( .A(u0__abc_49347_n1845_1), .B(u0__abc_49347_n1846_1), .Y(u0__abc_49347_n1847_1) );
  OR2X2 OR2X2_4040 ( .A(u3__abc_46775_n454), .B(mc_data_ir_8_), .Y(u3__abc_46775_n455) );
  OR2X2 OR2X2_4041 ( .A(u3__abc_46775_n453), .B(u3_byte1_0_), .Y(u3__abc_46775_n456) );
  OR2X2 OR2X2_4042 ( .A(u3__abc_46775_n457), .B(u3__abc_46775_n451), .Y(u3__abc_46775_n458) );
  OR2X2 OR2X2_4043 ( .A(u3__abc_46775_n459), .B(mc_data_ir_0_), .Y(u3__abc_46775_n460) );
  OR2X2 OR2X2_4044 ( .A(u3__abc_46775_n454), .B(mc_data_ir_9_), .Y(u3__abc_46775_n462) );
  OR2X2 OR2X2_4045 ( .A(u3__abc_46775_n453), .B(u3_byte1_1_), .Y(u3__abc_46775_n463) );
  OR2X2 OR2X2_4046 ( .A(u3__abc_46775_n464), .B(u3__abc_46775_n451), .Y(u3__abc_46775_n465) );
  OR2X2 OR2X2_4047 ( .A(u3__abc_46775_n459), .B(mc_data_ir_1_), .Y(u3__abc_46775_n466) );
  OR2X2 OR2X2_4048 ( .A(u3__abc_46775_n454), .B(mc_data_ir_10_), .Y(u3__abc_46775_n468) );
  OR2X2 OR2X2_4049 ( .A(u3__abc_46775_n453), .B(u3_byte1_2_), .Y(u3__abc_46775_n469) );
  OR2X2 OR2X2_405 ( .A(u0__abc_49347_n1849_1), .B(spec_req_cs_0_bF_buf5), .Y(u0__abc_49347_n1850_1) );
  OR2X2 OR2X2_4050 ( .A(u3__abc_46775_n470), .B(u3__abc_46775_n451), .Y(u3__abc_46775_n471) );
  OR2X2 OR2X2_4051 ( .A(u3__abc_46775_n459), .B(mc_data_ir_2_), .Y(u3__abc_46775_n472) );
  OR2X2 OR2X2_4052 ( .A(u3__abc_46775_n454), .B(mc_data_ir_11_), .Y(u3__abc_46775_n474) );
  OR2X2 OR2X2_4053 ( .A(u3__abc_46775_n453), .B(u3_byte1_3_), .Y(u3__abc_46775_n475) );
  OR2X2 OR2X2_4054 ( .A(u3__abc_46775_n476), .B(u3__abc_46775_n451), .Y(u3__abc_46775_n477) );
  OR2X2 OR2X2_4055 ( .A(u3__abc_46775_n459), .B(mc_data_ir_3_), .Y(u3__abc_46775_n478) );
  OR2X2 OR2X2_4056 ( .A(u3__abc_46775_n454), .B(mc_data_ir_12_), .Y(u3__abc_46775_n480) );
  OR2X2 OR2X2_4057 ( .A(u3__abc_46775_n453), .B(u3_byte1_4_), .Y(u3__abc_46775_n481) );
  OR2X2 OR2X2_4058 ( .A(u3__abc_46775_n482), .B(u3__abc_46775_n451), .Y(u3__abc_46775_n483) );
  OR2X2 OR2X2_4059 ( .A(u3__abc_46775_n459), .B(mc_data_ir_4_), .Y(u3__abc_46775_n484) );
  OR2X2 OR2X2_406 ( .A(u0__abc_49347_n1848_1), .B(u0__abc_49347_n1850_1), .Y(u0__abc_49347_n1851_1) );
  OR2X2 OR2X2_4060 ( .A(u3__abc_46775_n454), .B(mc_data_ir_13_), .Y(u3__abc_46775_n486) );
  OR2X2 OR2X2_4061 ( .A(u3__abc_46775_n453), .B(u3_byte1_5_), .Y(u3__abc_46775_n487) );
  OR2X2 OR2X2_4062 ( .A(u3__abc_46775_n488), .B(u3__abc_46775_n451), .Y(u3__abc_46775_n489) );
  OR2X2 OR2X2_4063 ( .A(u3__abc_46775_n459), .B(mc_data_ir_5_), .Y(u3__abc_46775_n490) );
  OR2X2 OR2X2_4064 ( .A(u3__abc_46775_n454), .B(mc_data_ir_14_), .Y(u3__abc_46775_n492) );
  OR2X2 OR2X2_4065 ( .A(u3__abc_46775_n453), .B(u3_byte1_6_), .Y(u3__abc_46775_n493) );
  OR2X2 OR2X2_4066 ( .A(u3__abc_46775_n494), .B(u3__abc_46775_n451), .Y(u3__abc_46775_n495) );
  OR2X2 OR2X2_4067 ( .A(u3__abc_46775_n459), .B(mc_data_ir_6_), .Y(u3__abc_46775_n496) );
  OR2X2 OR2X2_4068 ( .A(u3__abc_46775_n454), .B(mc_data_ir_15_), .Y(u3__abc_46775_n498) );
  OR2X2 OR2X2_4069 ( .A(u3__abc_46775_n453), .B(u3_byte1_7_), .Y(u3__abc_46775_n499) );
  OR2X2 OR2X2_407 ( .A(u0__abc_49347_n1203_bF_buf2), .B(u0_tms0_27_), .Y(u0__abc_49347_n1852_1) );
  OR2X2 OR2X2_4070 ( .A(u3__abc_46775_n500), .B(u3__abc_46775_n451), .Y(u3__abc_46775_n501) );
  OR2X2 OR2X2_4071 ( .A(u3__abc_46775_n459), .B(mc_data_ir_7_), .Y(u3__abc_46775_n502) );
  OR2X2 OR2X2_4072 ( .A(pack_le0), .B(u3_byte0_0_), .Y(u3__abc_46775_n504) );
  OR2X2 OR2X2_4073 ( .A(u3__abc_46775_n505), .B(mc_data_ir_0_), .Y(u3__abc_46775_n506) );
  OR2X2 OR2X2_4074 ( .A(pack_le0), .B(u3_byte0_1_), .Y(u3__abc_46775_n508) );
  OR2X2 OR2X2_4075 ( .A(u3__abc_46775_n505), .B(mc_data_ir_1_), .Y(u3__abc_46775_n509) );
  OR2X2 OR2X2_4076 ( .A(pack_le0), .B(u3_byte0_2_), .Y(u3__abc_46775_n511) );
  OR2X2 OR2X2_4077 ( .A(u3__abc_46775_n505), .B(mc_data_ir_2_), .Y(u3__abc_46775_n512) );
  OR2X2 OR2X2_4078 ( .A(pack_le0), .B(u3_byte0_3_), .Y(u3__abc_46775_n514) );
  OR2X2 OR2X2_4079 ( .A(u3__abc_46775_n505), .B(mc_data_ir_3_), .Y(u3__abc_46775_n515) );
  OR2X2 OR2X2_408 ( .A(u0__abc_49347_n1854_1), .B(u0__abc_49347_n1832_1), .Y(u0_sp_tms_27__FF_INPUT) );
  OR2X2 OR2X2_4080 ( .A(pack_le0), .B(u3_byte0_4_), .Y(u3__abc_46775_n517) );
  OR2X2 OR2X2_4081 ( .A(u3__abc_46775_n505), .B(mc_data_ir_4_), .Y(u3__abc_46775_n518) );
  OR2X2 OR2X2_4082 ( .A(pack_le0), .B(u3_byte0_5_), .Y(u3__abc_46775_n520) );
  OR2X2 OR2X2_4083 ( .A(u3__abc_46775_n505), .B(mc_data_ir_5_), .Y(u3__abc_46775_n521) );
  OR2X2 OR2X2_4084 ( .A(pack_le0), .B(u3_byte0_6_), .Y(u3__abc_46775_n523) );
  OR2X2 OR2X2_4085 ( .A(u3__abc_46775_n505), .B(mc_data_ir_6_), .Y(u3__abc_46775_n524) );
  OR2X2 OR2X2_4086 ( .A(pack_le0), .B(u3_byte0_7_), .Y(u3__abc_46775_n526) );
  OR2X2 OR2X2_4087 ( .A(u3__abc_46775_n505), .B(mc_data_ir_7_), .Y(u3__abc_46775_n527) );
  OR2X2 OR2X2_4088 ( .A(u3__abc_46775_n279_bF_buf1), .B(\wb_data_i[0] ), .Y(u3__abc_46775_n529) );
  OR2X2 OR2X2_4089 ( .A(u3__abc_46775_n277_1_bF_buf0), .B(mc_data_od_0_), .Y(u3__abc_46775_n530) );
  OR2X2 OR2X2_409 ( .A(u0__abc_49347_n1183_1_bF_buf1), .B(1'b0), .Y(u0__abc_49347_n1980) );
  OR2X2 OR2X2_4090 ( .A(u3__abc_46775_n279_bF_buf0), .B(\wb_data_i[1] ), .Y(u3__abc_46775_n532) );
  OR2X2 OR2X2_4091 ( .A(u3__abc_46775_n277_1_bF_buf5), .B(mc_data_od_1_), .Y(u3__abc_46775_n533) );
  OR2X2 OR2X2_4092 ( .A(u3__abc_46775_n279_bF_buf5), .B(\wb_data_i[2] ), .Y(u3__abc_46775_n535) );
  OR2X2 OR2X2_4093 ( .A(u3__abc_46775_n277_1_bF_buf4), .B(mc_data_od_2_), .Y(u3__abc_46775_n536) );
  OR2X2 OR2X2_4094 ( .A(u3__abc_46775_n279_bF_buf4), .B(\wb_data_i[3] ), .Y(u3__abc_46775_n538) );
  OR2X2 OR2X2_4095 ( .A(u3__abc_46775_n277_1_bF_buf3), .B(mc_data_od_3_), .Y(u3__abc_46775_n539) );
  OR2X2 OR2X2_4096 ( .A(u3__abc_46775_n279_bF_buf3), .B(\wb_data_i[4] ), .Y(u3__abc_46775_n541) );
  OR2X2 OR2X2_4097 ( .A(u3__abc_46775_n277_1_bF_buf2), .B(mc_data_od_4_), .Y(u3__abc_46775_n542) );
  OR2X2 OR2X2_4098 ( .A(u3__abc_46775_n279_bF_buf2), .B(\wb_data_i[5] ), .Y(u3__abc_46775_n544) );
  OR2X2 OR2X2_4099 ( .A(u3__abc_46775_n277_1_bF_buf1), .B(mc_data_od_5_), .Y(u3__abc_46775_n545) );
  OR2X2 OR2X2_41 ( .A(_abc_55805_n240_bF_buf0), .B(sp_tms_3_), .Y(_abc_55805_n299) );
  OR2X2 OR2X2_410 ( .A(spec_req_cs_6_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n1981_1) );
  OR2X2 OR2X2_4100 ( .A(u3__abc_46775_n279_bF_buf1), .B(\wb_data_i[6] ), .Y(u3__abc_46775_n547) );
  OR2X2 OR2X2_4101 ( .A(u3__abc_46775_n277_1_bF_buf0), .B(mc_data_od_6_), .Y(u3__abc_46775_n548) );
  OR2X2 OR2X2_4102 ( .A(u3__abc_46775_n279_bF_buf0), .B(\wb_data_i[7] ), .Y(u3__abc_46775_n550) );
  OR2X2 OR2X2_4103 ( .A(u3__abc_46775_n277_1_bF_buf5), .B(mc_data_od_7_), .Y(u3__abc_46775_n551) );
  OR2X2 OR2X2_4104 ( .A(u3__abc_46775_n279_bF_buf5), .B(\wb_data_i[8] ), .Y(u3__abc_46775_n553) );
  OR2X2 OR2X2_4105 ( .A(u3__abc_46775_n277_1_bF_buf4), .B(mc_data_od_8_), .Y(u3__abc_46775_n554) );
  OR2X2 OR2X2_4106 ( .A(u3__abc_46775_n279_bF_buf4), .B(\wb_data_i[9] ), .Y(u3__abc_46775_n556) );
  OR2X2 OR2X2_4107 ( .A(u3__abc_46775_n277_1_bF_buf3), .B(mc_data_od_9_), .Y(u3__abc_46775_n557) );
  OR2X2 OR2X2_4108 ( .A(u3__abc_46775_n279_bF_buf3), .B(\wb_data_i[10] ), .Y(u3__abc_46775_n559) );
  OR2X2 OR2X2_4109 ( .A(u3__abc_46775_n277_1_bF_buf2), .B(mc_data_od_10_), .Y(u3__abc_46775_n560) );
  OR2X2 OR2X2_411 ( .A(u0__abc_49347_n1983_1), .B(u0__abc_49347_n1979_1), .Y(u0__abc_49347_n1984_1) );
  OR2X2 OR2X2_4110 ( .A(u3__abc_46775_n279_bF_buf2), .B(\wb_data_i[11] ), .Y(u3__abc_46775_n562) );
  OR2X2 OR2X2_4111 ( .A(u3__abc_46775_n277_1_bF_buf1), .B(mc_data_od_11_), .Y(u3__abc_46775_n563) );
  OR2X2 OR2X2_4112 ( .A(u3__abc_46775_n279_bF_buf1), .B(\wb_data_i[12] ), .Y(u3__abc_46775_n565) );
  OR2X2 OR2X2_4113 ( .A(u3__abc_46775_n277_1_bF_buf0), .B(mc_data_od_12_), .Y(u3__abc_46775_n566) );
  OR2X2 OR2X2_4114 ( .A(u3__abc_46775_n279_bF_buf0), .B(\wb_data_i[13] ), .Y(u3__abc_46775_n568) );
  OR2X2 OR2X2_4115 ( .A(u3__abc_46775_n277_1_bF_buf5), .B(mc_data_od_13_), .Y(u3__abc_46775_n569) );
  OR2X2 OR2X2_4116 ( .A(u3__abc_46775_n279_bF_buf5), .B(\wb_data_i[14] ), .Y(u3__abc_46775_n571) );
  OR2X2 OR2X2_4117 ( .A(u3__abc_46775_n277_1_bF_buf4), .B(mc_data_od_14_), .Y(u3__abc_46775_n572) );
  OR2X2 OR2X2_4118 ( .A(u3__abc_46775_n279_bF_buf4), .B(\wb_data_i[15] ), .Y(u3__abc_46775_n574) );
  OR2X2 OR2X2_4119 ( .A(u3__abc_46775_n277_1_bF_buf3), .B(mc_data_od_15_), .Y(u3__abc_46775_n575) );
  OR2X2 OR2X2_412 ( .A(u0__abc_49347_n1985), .B(u0__abc_49347_n1986), .Y(u0__abc_49347_n1987) );
  OR2X2 OR2X2_4120 ( .A(u3__abc_46775_n279_bF_buf3), .B(\wb_data_i[16] ), .Y(u3__abc_46775_n577) );
  OR2X2 OR2X2_4121 ( .A(u3__abc_46775_n277_1_bF_buf2), .B(mc_data_od_16_), .Y(u3__abc_46775_n578) );
  OR2X2 OR2X2_4122 ( .A(u3__abc_46775_n279_bF_buf2), .B(\wb_data_i[17] ), .Y(u3__abc_46775_n580) );
  OR2X2 OR2X2_4123 ( .A(u3__abc_46775_n277_1_bF_buf1), .B(mc_data_od_17_), .Y(u3__abc_46775_n581) );
  OR2X2 OR2X2_4124 ( .A(u3__abc_46775_n279_bF_buf1), .B(\wb_data_i[18] ), .Y(u3__abc_46775_n583) );
  OR2X2 OR2X2_4125 ( .A(u3__abc_46775_n277_1_bF_buf0), .B(mc_data_od_18_), .Y(u3__abc_46775_n584) );
  OR2X2 OR2X2_4126 ( .A(u3__abc_46775_n279_bF_buf0), .B(\wb_data_i[19] ), .Y(u3__abc_46775_n586) );
  OR2X2 OR2X2_4127 ( .A(u3__abc_46775_n277_1_bF_buf5), .B(mc_data_od_19_), .Y(u3__abc_46775_n587) );
  OR2X2 OR2X2_4128 ( .A(u3__abc_46775_n279_bF_buf5), .B(\wb_data_i[20] ), .Y(u3__abc_46775_n589) );
  OR2X2 OR2X2_4129 ( .A(u3__abc_46775_n277_1_bF_buf4), .B(mc_data_od_20_), .Y(u3__abc_46775_n590) );
  OR2X2 OR2X2_413 ( .A(u0__abc_49347_n1988), .B(u0__abc_49347_n1989), .Y(u0__abc_49347_n1990) );
  OR2X2 OR2X2_4130 ( .A(u3__abc_46775_n279_bF_buf4), .B(\wb_data_i[21] ), .Y(u3__abc_46775_n592) );
  OR2X2 OR2X2_4131 ( .A(u3__abc_46775_n277_1_bF_buf3), .B(mc_data_od_21_), .Y(u3__abc_46775_n593) );
  OR2X2 OR2X2_4132 ( .A(u3__abc_46775_n279_bF_buf3), .B(\wb_data_i[22] ), .Y(u3__abc_46775_n595) );
  OR2X2 OR2X2_4133 ( .A(u3__abc_46775_n277_1_bF_buf2), .B(mc_data_od_22_), .Y(u3__abc_46775_n596) );
  OR2X2 OR2X2_4134 ( .A(u3__abc_46775_n279_bF_buf2), .B(\wb_data_i[23] ), .Y(u3__abc_46775_n598) );
  OR2X2 OR2X2_4135 ( .A(u3__abc_46775_n277_1_bF_buf1), .B(mc_data_od_23_), .Y(u3__abc_46775_n599) );
  OR2X2 OR2X2_4136 ( .A(u3__abc_46775_n279_bF_buf1), .B(\wb_data_i[24] ), .Y(u3__abc_46775_n601) );
  OR2X2 OR2X2_4137 ( .A(u3__abc_46775_n277_1_bF_buf0), .B(mc_data_od_24_), .Y(u3__abc_46775_n602) );
  OR2X2 OR2X2_4138 ( .A(u3__abc_46775_n279_bF_buf0), .B(\wb_data_i[25] ), .Y(u3__abc_46775_n604) );
  OR2X2 OR2X2_4139 ( .A(u3__abc_46775_n277_1_bF_buf5), .B(mc_data_od_25_), .Y(u3__abc_46775_n605) );
  OR2X2 OR2X2_414 ( .A(u0__abc_49347_n1991), .B(u0__abc_49347_n1992), .Y(u0__abc_49347_n1993) );
  OR2X2 OR2X2_4140 ( .A(u3__abc_46775_n279_bF_buf5), .B(\wb_data_i[26] ), .Y(u3__abc_46775_n607) );
  OR2X2 OR2X2_4141 ( .A(u3__abc_46775_n277_1_bF_buf4), .B(mc_data_od_26_), .Y(u3__abc_46775_n608) );
  OR2X2 OR2X2_4142 ( .A(u3__abc_46775_n279_bF_buf4), .B(\wb_data_i[27] ), .Y(u3__abc_46775_n610) );
  OR2X2 OR2X2_4143 ( .A(u3__abc_46775_n277_1_bF_buf3), .B(mc_data_od_27_), .Y(u3__abc_46775_n611) );
  OR2X2 OR2X2_4144 ( .A(u3__abc_46775_n279_bF_buf3), .B(\wb_data_i[28] ), .Y(u3__abc_46775_n613) );
  OR2X2 OR2X2_4145 ( .A(u3__abc_46775_n277_1_bF_buf2), .B(mc_data_od_28_), .Y(u3__abc_46775_n614) );
  OR2X2 OR2X2_4146 ( .A(u3__abc_46775_n279_bF_buf2), .B(\wb_data_i[29] ), .Y(u3__abc_46775_n616) );
  OR2X2 OR2X2_4147 ( .A(u3__abc_46775_n277_1_bF_buf1), .B(mc_data_od_29_), .Y(u3__abc_46775_n617) );
  OR2X2 OR2X2_4148 ( .A(u3__abc_46775_n279_bF_buf1), .B(\wb_data_i[30] ), .Y(u3__abc_46775_n619) );
  OR2X2 OR2X2_4149 ( .A(u3__abc_46775_n277_1_bF_buf0), .B(mc_data_od_30_), .Y(u3__abc_46775_n620) );
  OR2X2 OR2X2_415 ( .A(u0__abc_49347_n1995), .B(spec_req_cs_0_bF_buf4), .Y(u0__abc_49347_n1996) );
  OR2X2 OR2X2_4150 ( .A(u3__abc_46775_n279_bF_buf0), .B(\wb_data_i[31] ), .Y(u3__abc_46775_n622) );
  OR2X2 OR2X2_4151 ( .A(u3__abc_46775_n277_1_bF_buf5), .B(mc_data_od_31_), .Y(u3__abc_46775_n623) );
  OR2X2 OR2X2_4152 ( .A(csc_5_bF_buf1), .B(u3_byte0_0_), .Y(u3__abc_46775_n626) );
  OR2X2 OR2X2_4153 ( .A(u3__abc_46775_n448_bF_buf1), .B(mc_data_ir_0_), .Y(u3__abc_46775_n627) );
  OR2X2 OR2X2_4154 ( .A(u3__abc_46775_n628), .B(u3__abc_46775_n625_bF_buf4), .Y(u3__abc_46775_n629) );
  OR2X2 OR2X2_4155 ( .A(u3__abc_46775_n275_bF_buf2), .B(u3_rd_fifo_out_0_), .Y(u3__abc_46775_n630) );
  OR2X2 OR2X2_4156 ( .A(csc_5_bF_buf0), .B(u3_byte0_1_), .Y(u3__abc_46775_n632) );
  OR2X2 OR2X2_4157 ( .A(u3__abc_46775_n448_bF_buf0), .B(mc_data_ir_1_), .Y(u3__abc_46775_n633) );
  OR2X2 OR2X2_4158 ( .A(u3__abc_46775_n634), .B(u3__abc_46775_n625_bF_buf3), .Y(u3__abc_46775_n635) );
  OR2X2 OR2X2_4159 ( .A(u3__abc_46775_n275_bF_buf1), .B(u3_rd_fifo_out_1_), .Y(u3__abc_46775_n636) );
  OR2X2 OR2X2_416 ( .A(u0__abc_49347_n1994), .B(u0__abc_49347_n1996), .Y(u0__abc_49347_n1997) );
  OR2X2 OR2X2_4160 ( .A(csc_5_bF_buf4), .B(u3_byte0_2_), .Y(u3__abc_46775_n638) );
  OR2X2 OR2X2_4161 ( .A(u3__abc_46775_n448_bF_buf3), .B(mc_data_ir_2_), .Y(u3__abc_46775_n639) );
  OR2X2 OR2X2_4162 ( .A(u3__abc_46775_n640), .B(u3__abc_46775_n625_bF_buf2), .Y(u3__abc_46775_n641) );
  OR2X2 OR2X2_4163 ( .A(u3__abc_46775_n275_bF_buf0), .B(u3_rd_fifo_out_2_), .Y(u3__abc_46775_n642) );
  OR2X2 OR2X2_4164 ( .A(csc_5_bF_buf3), .B(u3_byte0_3_), .Y(u3__abc_46775_n644) );
  OR2X2 OR2X2_4165 ( .A(u3__abc_46775_n448_bF_buf2), .B(mc_data_ir_3_), .Y(u3__abc_46775_n645) );
  OR2X2 OR2X2_4166 ( .A(u3__abc_46775_n646), .B(u3__abc_46775_n625_bF_buf1), .Y(u3__abc_46775_n647) );
  OR2X2 OR2X2_4167 ( .A(u3__abc_46775_n275_bF_buf4), .B(u3_rd_fifo_out_3_), .Y(u3__abc_46775_n648) );
  OR2X2 OR2X2_4168 ( .A(csc_5_bF_buf2), .B(u3_byte0_4_), .Y(u3__abc_46775_n650) );
  OR2X2 OR2X2_4169 ( .A(u3__abc_46775_n448_bF_buf1), .B(mc_data_ir_4_), .Y(u3__abc_46775_n651) );
  OR2X2 OR2X2_417 ( .A(u0__abc_49347_n1203_bF_buf1), .B(u0_csc0_1_), .Y(u0__abc_49347_n1998) );
  OR2X2 OR2X2_4170 ( .A(u3__abc_46775_n652), .B(u3__abc_46775_n625_bF_buf0), .Y(u3__abc_46775_n653) );
  OR2X2 OR2X2_4171 ( .A(u3__abc_46775_n275_bF_buf3), .B(u3_rd_fifo_out_4_), .Y(u3__abc_46775_n654) );
  OR2X2 OR2X2_4172 ( .A(csc_5_bF_buf1), .B(u3_byte0_5_), .Y(u3__abc_46775_n656) );
  OR2X2 OR2X2_4173 ( .A(u3__abc_46775_n448_bF_buf0), .B(mc_data_ir_5_), .Y(u3__abc_46775_n657) );
  OR2X2 OR2X2_4174 ( .A(u3__abc_46775_n658), .B(u3__abc_46775_n625_bF_buf4), .Y(u3__abc_46775_n659) );
  OR2X2 OR2X2_4175 ( .A(u3__abc_46775_n275_bF_buf2), .B(u3_rd_fifo_out_5_), .Y(u3__abc_46775_n660) );
  OR2X2 OR2X2_4176 ( .A(csc_5_bF_buf0), .B(u3_byte0_6_), .Y(u3__abc_46775_n662) );
  OR2X2 OR2X2_4177 ( .A(u3__abc_46775_n448_bF_buf3), .B(mc_data_ir_6_), .Y(u3__abc_46775_n663) );
  OR2X2 OR2X2_4178 ( .A(u3__abc_46775_n664), .B(u3__abc_46775_n625_bF_buf3), .Y(u3__abc_46775_n665) );
  OR2X2 OR2X2_4179 ( .A(u3__abc_46775_n275_bF_buf1), .B(u3_rd_fifo_out_6_), .Y(u3__abc_46775_n666) );
  OR2X2 OR2X2_418 ( .A(u0__abc_49347_n2000), .B(u0__abc_49347_n1978), .Y(u0_sp_csc_1__FF_INPUT) );
  OR2X2 OR2X2_4180 ( .A(csc_5_bF_buf4), .B(u3_byte0_7_), .Y(u3__abc_46775_n668) );
  OR2X2 OR2X2_4181 ( .A(u3__abc_46775_n448_bF_buf2), .B(mc_data_ir_7_), .Y(u3__abc_46775_n669) );
  OR2X2 OR2X2_4182 ( .A(u3__abc_46775_n670), .B(u3__abc_46775_n625_bF_buf2), .Y(u3__abc_46775_n671) );
  OR2X2 OR2X2_4183 ( .A(u3__abc_46775_n275_bF_buf0), .B(u3_rd_fifo_out_7_), .Y(u3__abc_46775_n672) );
  OR2X2 OR2X2_4184 ( .A(csc_5_bF_buf3), .B(u3_byte1_0_), .Y(u3__abc_46775_n674) );
  OR2X2 OR2X2_4185 ( .A(u3__abc_46775_n448_bF_buf1), .B(mc_data_ir_8_), .Y(u3__abc_46775_n675) );
  OR2X2 OR2X2_4186 ( .A(u3__abc_46775_n676), .B(u3__abc_46775_n625_bF_buf1), .Y(u3__abc_46775_n677) );
  OR2X2 OR2X2_4187 ( .A(u3__abc_46775_n275_bF_buf4), .B(u3_rd_fifo_out_8_), .Y(u3__abc_46775_n678) );
  OR2X2 OR2X2_4188 ( .A(csc_5_bF_buf2), .B(u3_byte1_1_), .Y(u3__abc_46775_n680) );
  OR2X2 OR2X2_4189 ( .A(u3__abc_46775_n448_bF_buf0), .B(mc_data_ir_9_), .Y(u3__abc_46775_n681) );
  OR2X2 OR2X2_419 ( .A(u0__abc_49347_n1183_1_bF_buf0), .B(1'b0), .Y(u0__abc_49347_n2004) );
  OR2X2 OR2X2_4190 ( .A(u3__abc_46775_n682), .B(u3__abc_46775_n625_bF_buf0), .Y(u3__abc_46775_n683) );
  OR2X2 OR2X2_4191 ( .A(u3__abc_46775_n275_bF_buf3), .B(u3_rd_fifo_out_9_), .Y(u3__abc_46775_n684) );
  OR2X2 OR2X2_4192 ( .A(csc_5_bF_buf1), .B(u3_byte1_2_), .Y(u3__abc_46775_n686) );
  OR2X2 OR2X2_4193 ( .A(u3__abc_46775_n448_bF_buf3), .B(mc_data_ir_10_), .Y(u3__abc_46775_n687) );
  OR2X2 OR2X2_4194 ( .A(u3__abc_46775_n688), .B(u3__abc_46775_n625_bF_buf4), .Y(u3__abc_46775_n689) );
  OR2X2 OR2X2_4195 ( .A(u3__abc_46775_n275_bF_buf2), .B(u3_rd_fifo_out_10_), .Y(u3__abc_46775_n690) );
  OR2X2 OR2X2_4196 ( .A(csc_5_bF_buf0), .B(u3_byte1_3_), .Y(u3__abc_46775_n692) );
  OR2X2 OR2X2_4197 ( .A(u3__abc_46775_n448_bF_buf2), .B(mc_data_ir_11_), .Y(u3__abc_46775_n693) );
  OR2X2 OR2X2_4198 ( .A(u3__abc_46775_n694), .B(u3__abc_46775_n625_bF_buf3), .Y(u3__abc_46775_n695) );
  OR2X2 OR2X2_4199 ( .A(u3__abc_46775_n275_bF_buf1), .B(u3_rd_fifo_out_11_), .Y(u3__abc_46775_n696) );
  OR2X2 OR2X2_42 ( .A(lmr_sel_bF_buf2), .B(tms_3_), .Y(_abc_55805_n300) );
  OR2X2 OR2X2_420 ( .A(spec_req_cs_6_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n2005) );
  OR2X2 OR2X2_4200 ( .A(csc_5_bF_buf4), .B(u3_byte1_4_), .Y(u3__abc_46775_n698) );
  OR2X2 OR2X2_4201 ( .A(u3__abc_46775_n448_bF_buf1), .B(mc_data_ir_12_), .Y(u3__abc_46775_n699) );
  OR2X2 OR2X2_4202 ( .A(u3__abc_46775_n700), .B(u3__abc_46775_n625_bF_buf2), .Y(u3__abc_46775_n701) );
  OR2X2 OR2X2_4203 ( .A(u3__abc_46775_n275_bF_buf0), .B(u3_rd_fifo_out_12_), .Y(u3__abc_46775_n702) );
  OR2X2 OR2X2_4204 ( .A(csc_5_bF_buf3), .B(u3_byte1_5_), .Y(u3__abc_46775_n704) );
  OR2X2 OR2X2_4205 ( .A(u3__abc_46775_n448_bF_buf0), .B(mc_data_ir_13_), .Y(u3__abc_46775_n705) );
  OR2X2 OR2X2_4206 ( .A(u3__abc_46775_n706), .B(u3__abc_46775_n625_bF_buf1), .Y(u3__abc_46775_n707) );
  OR2X2 OR2X2_4207 ( .A(u3__abc_46775_n275_bF_buf4), .B(u3_rd_fifo_out_13_), .Y(u3__abc_46775_n708) );
  OR2X2 OR2X2_4208 ( .A(csc_5_bF_buf2), .B(u3_byte1_6_), .Y(u3__abc_46775_n710) );
  OR2X2 OR2X2_4209 ( .A(u3__abc_46775_n448_bF_buf3), .B(mc_data_ir_14_), .Y(u3__abc_46775_n711) );
  OR2X2 OR2X2_421 ( .A(u0__abc_49347_n2007), .B(u0__abc_49347_n2003), .Y(u0__abc_49347_n2008) );
  OR2X2 OR2X2_4210 ( .A(u3__abc_46775_n712), .B(u3__abc_46775_n625_bF_buf0), .Y(u3__abc_46775_n713) );
  OR2X2 OR2X2_4211 ( .A(u3__abc_46775_n275_bF_buf3), .B(u3_rd_fifo_out_14_), .Y(u3__abc_46775_n714) );
  OR2X2 OR2X2_4212 ( .A(csc_5_bF_buf1), .B(u3_byte1_7_), .Y(u3__abc_46775_n716) );
  OR2X2 OR2X2_4213 ( .A(u3__abc_46775_n448_bF_buf2), .B(mc_data_ir_15_), .Y(u3__abc_46775_n717) );
  OR2X2 OR2X2_4214 ( .A(u3__abc_46775_n718), .B(u3__abc_46775_n625_bF_buf4), .Y(u3__abc_46775_n719) );
  OR2X2 OR2X2_4215 ( .A(u3__abc_46775_n275_bF_buf2), .B(u3_rd_fifo_out_15_), .Y(u3__abc_46775_n720) );
  OR2X2 OR2X2_4216 ( .A(u3__abc_46775_n722), .B(u3__abc_46775_n723), .Y(u3__abc_46775_n724) );
  OR2X2 OR2X2_4217 ( .A(u3__abc_46775_n725), .B(u3__abc_46775_n625_bF_buf3), .Y(u3__abc_46775_n726) );
  OR2X2 OR2X2_4218 ( .A(u3__abc_46775_n726), .B(u3__abc_46775_n724), .Y(u3__abc_46775_n727) );
  OR2X2 OR2X2_4219 ( .A(u3__abc_46775_n275_bF_buf1), .B(u3_rd_fifo_out_16_), .Y(u3__abc_46775_n728) );
  OR2X2 OR2X2_422 ( .A(u0__abc_49347_n2009), .B(u0__abc_49347_n2010), .Y(u0__abc_49347_n2011) );
  OR2X2 OR2X2_4220 ( .A(u3__abc_46775_n730), .B(u3__abc_46775_n731), .Y(u3__abc_46775_n732) );
  OR2X2 OR2X2_4221 ( .A(u3__abc_46775_n733), .B(u3__abc_46775_n625_bF_buf2), .Y(u3__abc_46775_n734) );
  OR2X2 OR2X2_4222 ( .A(u3__abc_46775_n734), .B(u3__abc_46775_n732), .Y(u3__abc_46775_n735) );
  OR2X2 OR2X2_4223 ( .A(u3__abc_46775_n275_bF_buf0), .B(u3_rd_fifo_out_17_), .Y(u3__abc_46775_n736) );
  OR2X2 OR2X2_4224 ( .A(u3__abc_46775_n738), .B(u3__abc_46775_n739), .Y(u3__abc_46775_n740) );
  OR2X2 OR2X2_4225 ( .A(u3__abc_46775_n741), .B(u3__abc_46775_n625_bF_buf1), .Y(u3__abc_46775_n742) );
  OR2X2 OR2X2_4226 ( .A(u3__abc_46775_n742), .B(u3__abc_46775_n740), .Y(u3__abc_46775_n743) );
  OR2X2 OR2X2_4227 ( .A(u3__abc_46775_n275_bF_buf4), .B(u3_rd_fifo_out_18_), .Y(u3__abc_46775_n744) );
  OR2X2 OR2X2_4228 ( .A(u3__abc_46775_n746), .B(u3__abc_46775_n747), .Y(u3__abc_46775_n748) );
  OR2X2 OR2X2_4229 ( .A(u3__abc_46775_n749), .B(u3__abc_46775_n625_bF_buf0), .Y(u3__abc_46775_n750) );
  OR2X2 OR2X2_423 ( .A(u0__abc_49347_n2012), .B(u0__abc_49347_n2013), .Y(u0__abc_49347_n2014) );
  OR2X2 OR2X2_4230 ( .A(u3__abc_46775_n750), .B(u3__abc_46775_n748), .Y(u3__abc_46775_n751) );
  OR2X2 OR2X2_4231 ( .A(u3__abc_46775_n275_bF_buf3), .B(u3_rd_fifo_out_19_), .Y(u3__abc_46775_n752) );
  OR2X2 OR2X2_4232 ( .A(u3__abc_46775_n754), .B(u3__abc_46775_n755), .Y(u3__abc_46775_n756) );
  OR2X2 OR2X2_4233 ( .A(u3__abc_46775_n757), .B(u3__abc_46775_n625_bF_buf4), .Y(u3__abc_46775_n758) );
  OR2X2 OR2X2_4234 ( .A(u3__abc_46775_n758), .B(u3__abc_46775_n756), .Y(u3__abc_46775_n759) );
  OR2X2 OR2X2_4235 ( .A(u3__abc_46775_n275_bF_buf2), .B(u3_rd_fifo_out_20_), .Y(u3__abc_46775_n760) );
  OR2X2 OR2X2_4236 ( .A(u3__abc_46775_n762), .B(u3__abc_46775_n763), .Y(u3__abc_46775_n764) );
  OR2X2 OR2X2_4237 ( .A(u3__abc_46775_n765), .B(u3__abc_46775_n625_bF_buf3), .Y(u3__abc_46775_n766) );
  OR2X2 OR2X2_4238 ( .A(u3__abc_46775_n766), .B(u3__abc_46775_n764), .Y(u3__abc_46775_n767) );
  OR2X2 OR2X2_4239 ( .A(u3__abc_46775_n275_bF_buf1), .B(u3_rd_fifo_out_21_), .Y(u3__abc_46775_n768) );
  OR2X2 OR2X2_424 ( .A(u0__abc_49347_n2015), .B(u0__abc_49347_n2016), .Y(u0__abc_49347_n2017) );
  OR2X2 OR2X2_4240 ( .A(u3__abc_46775_n770), .B(u3__abc_46775_n771), .Y(u3__abc_46775_n772) );
  OR2X2 OR2X2_4241 ( .A(u3__abc_46775_n773), .B(u3__abc_46775_n625_bF_buf2), .Y(u3__abc_46775_n774) );
  OR2X2 OR2X2_4242 ( .A(u3__abc_46775_n774), .B(u3__abc_46775_n772), .Y(u3__abc_46775_n775) );
  OR2X2 OR2X2_4243 ( .A(u3__abc_46775_n275_bF_buf0), .B(u3_rd_fifo_out_22_), .Y(u3__abc_46775_n776) );
  OR2X2 OR2X2_4244 ( .A(u3__abc_46775_n778), .B(u3__abc_46775_n779), .Y(u3__abc_46775_n780) );
  OR2X2 OR2X2_4245 ( .A(u3__abc_46775_n781), .B(u3__abc_46775_n625_bF_buf1), .Y(u3__abc_46775_n782) );
  OR2X2 OR2X2_4246 ( .A(u3__abc_46775_n782), .B(u3__abc_46775_n780), .Y(u3__abc_46775_n783) );
  OR2X2 OR2X2_4247 ( .A(u3__abc_46775_n275_bF_buf4), .B(u3_rd_fifo_out_23_), .Y(u3__abc_46775_n784) );
  OR2X2 OR2X2_4248 ( .A(u3__abc_46775_n786), .B(u3__abc_46775_n787), .Y(u3__abc_46775_n788) );
  OR2X2 OR2X2_4249 ( .A(u3__abc_46775_n789), .B(u3__abc_46775_n625_bF_buf0), .Y(u3__abc_46775_n790) );
  OR2X2 OR2X2_425 ( .A(u0__abc_49347_n2019), .B(spec_req_cs_0_bF_buf3), .Y(u0__abc_49347_n2020) );
  OR2X2 OR2X2_4250 ( .A(u3__abc_46775_n790), .B(u3__abc_46775_n788), .Y(u3__abc_46775_n791) );
  OR2X2 OR2X2_4251 ( .A(u3__abc_46775_n275_bF_buf3), .B(u3_rd_fifo_out_24_), .Y(u3__abc_46775_n792) );
  OR2X2 OR2X2_4252 ( .A(u3__abc_46775_n794), .B(u3__abc_46775_n795), .Y(u3__abc_46775_n796) );
  OR2X2 OR2X2_4253 ( .A(u3__abc_46775_n797), .B(u3__abc_46775_n625_bF_buf4), .Y(u3__abc_46775_n798) );
  OR2X2 OR2X2_4254 ( .A(u3__abc_46775_n798), .B(u3__abc_46775_n796), .Y(u3__abc_46775_n799) );
  OR2X2 OR2X2_4255 ( .A(u3__abc_46775_n275_bF_buf2), .B(u3_rd_fifo_out_25_), .Y(u3__abc_46775_n800) );
  OR2X2 OR2X2_4256 ( .A(u3__abc_46775_n802), .B(u3__abc_46775_n803), .Y(u3__abc_46775_n804) );
  OR2X2 OR2X2_4257 ( .A(u3__abc_46775_n805), .B(u3__abc_46775_n625_bF_buf3), .Y(u3__abc_46775_n806) );
  OR2X2 OR2X2_4258 ( .A(u3__abc_46775_n806), .B(u3__abc_46775_n804), .Y(u3__abc_46775_n807) );
  OR2X2 OR2X2_4259 ( .A(u3__abc_46775_n275_bF_buf1), .B(u3_rd_fifo_out_26_), .Y(u3__abc_46775_n808) );
  OR2X2 OR2X2_426 ( .A(u0__abc_49347_n2018), .B(u0__abc_49347_n2020), .Y(u0__abc_49347_n2021) );
  OR2X2 OR2X2_4260 ( .A(u3__abc_46775_n810), .B(u3__abc_46775_n811), .Y(u3__abc_46775_n812) );
  OR2X2 OR2X2_4261 ( .A(u3__abc_46775_n813), .B(u3__abc_46775_n625_bF_buf2), .Y(u3__abc_46775_n814) );
  OR2X2 OR2X2_4262 ( .A(u3__abc_46775_n814), .B(u3__abc_46775_n812), .Y(u3__abc_46775_n815) );
  OR2X2 OR2X2_4263 ( .A(u3__abc_46775_n275_bF_buf0), .B(u3_rd_fifo_out_27_), .Y(u3__abc_46775_n816) );
  OR2X2 OR2X2_4264 ( .A(u3__abc_46775_n818), .B(u3__abc_46775_n819), .Y(u3__abc_46775_n820) );
  OR2X2 OR2X2_4265 ( .A(u3__abc_46775_n821), .B(u3__abc_46775_n625_bF_buf1), .Y(u3__abc_46775_n822) );
  OR2X2 OR2X2_4266 ( .A(u3__abc_46775_n822), .B(u3__abc_46775_n820), .Y(u3__abc_46775_n823) );
  OR2X2 OR2X2_4267 ( .A(u3__abc_46775_n275_bF_buf4), .B(u3_rd_fifo_out_28_), .Y(u3__abc_46775_n824) );
  OR2X2 OR2X2_4268 ( .A(u3__abc_46775_n826), .B(u3__abc_46775_n827), .Y(u3__abc_46775_n828) );
  OR2X2 OR2X2_4269 ( .A(u3__abc_46775_n829), .B(u3__abc_46775_n625_bF_buf0), .Y(u3__abc_46775_n830) );
  OR2X2 OR2X2_427 ( .A(u0__abc_49347_n1203_bF_buf0), .B(u0_csc0_2_), .Y(u0__abc_49347_n2022) );
  OR2X2 OR2X2_4270 ( .A(u3__abc_46775_n830), .B(u3__abc_46775_n828), .Y(u3__abc_46775_n831) );
  OR2X2 OR2X2_4271 ( .A(u3__abc_46775_n275_bF_buf3), .B(u3_rd_fifo_out_29_), .Y(u3__abc_46775_n832) );
  OR2X2 OR2X2_4272 ( .A(u3__abc_46775_n834), .B(u3__abc_46775_n835), .Y(u3__abc_46775_n836) );
  OR2X2 OR2X2_4273 ( .A(u3__abc_46775_n837), .B(u3__abc_46775_n625_bF_buf4), .Y(u3__abc_46775_n838) );
  OR2X2 OR2X2_4274 ( .A(u3__abc_46775_n838), .B(u3__abc_46775_n836), .Y(u3__abc_46775_n839) );
  OR2X2 OR2X2_4275 ( .A(u3__abc_46775_n275_bF_buf2), .B(u3_rd_fifo_out_30_), .Y(u3__abc_46775_n840) );
  OR2X2 OR2X2_4276 ( .A(u3__abc_46775_n842), .B(u3__abc_46775_n843), .Y(u3__abc_46775_n844) );
  OR2X2 OR2X2_4277 ( .A(u3__abc_46775_n845), .B(u3__abc_46775_n625_bF_buf3), .Y(u3__abc_46775_n846) );
  OR2X2 OR2X2_4278 ( .A(u3__abc_46775_n846), .B(u3__abc_46775_n844), .Y(u3__abc_46775_n847) );
  OR2X2 OR2X2_4279 ( .A(u3__abc_46775_n275_bF_buf1), .B(u3_rd_fifo_out_31_), .Y(u3__abc_46775_n848) );
  OR2X2 OR2X2_428 ( .A(u0__abc_49347_n2024), .B(u0__abc_49347_n2002), .Y(u0_sp_csc_2__FF_INPUT) );
  OR2X2 OR2X2_4280 ( .A(u3__abc_46775_n851), .B(u3__abc_46775_n850), .Y(u3_rd_fifo_clr) );
  OR2X2 OR2X2_4281 ( .A(u3_rd_fifo_out_14_), .B(u3_rd_fifo_out_15_), .Y(u3__abc_46775_n854) );
  OR2X2 OR2X2_4282 ( .A(u3__abc_46775_n861), .B(u3__abc_46775_n863), .Y(u3__abc_46775_n864) );
  OR2X2 OR2X2_4283 ( .A(u3__abc_46775_n864), .B(u3__abc_46775_n859), .Y(u3__abc_46775_n865) );
  OR2X2 OR2X2_4284 ( .A(u3__abc_46775_n862), .B(u3_rd_fifo_out_9_), .Y(u3__abc_46775_n866) );
  OR2X2 OR2X2_4285 ( .A(u3__abc_46775_n860), .B(u3_rd_fifo_out_8_), .Y(u3__abc_46775_n867) );
  OR2X2 OR2X2_4286 ( .A(u3__abc_46775_n868), .B(u3_rd_fifo_out_33_), .Y(u3__abc_46775_n869) );
  OR2X2 OR2X2_4287 ( .A(u3__abc_46775_n870), .B(u3__abc_46775_n858), .Y(u3__abc_46775_n871) );
  OR2X2 OR2X2_4288 ( .A(u3__abc_46775_n868), .B(u3__abc_46775_n859), .Y(u3__abc_46775_n872) );
  OR2X2 OR2X2_4289 ( .A(u3__abc_46775_n864), .B(u3_rd_fifo_out_33_), .Y(u3__abc_46775_n873) );
  OR2X2 OR2X2_429 ( .A(u0__abc_49347_n1183_1_bF_buf5), .B(1'b0), .Y(u0__abc_49347_n2028) );
  OR2X2 OR2X2_4290 ( .A(u3__abc_46775_n874), .B(u3__abc_46775_n857), .Y(u3__abc_46775_n875) );
  OR2X2 OR2X2_4291 ( .A(u3_rd_fifo_out_12_), .B(u3_rd_fifo_out_13_), .Y(u3__abc_46775_n878) );
  OR2X2 OR2X2_4292 ( .A(u3__abc_46775_n883), .B(u3_rd_fifo_out_10_), .Y(u3__abc_46775_n886) );
  OR2X2 OR2X2_4293 ( .A(u3__abc_46775_n889), .B(u3__abc_46775_n890), .Y(u3__abc_46775_n891) );
  OR2X2 OR2X2_4294 ( .A(u3__abc_46775_n877), .B(u3__abc_46775_n892), .Y(u3__abc_46775_n893) );
  OR2X2 OR2X2_4295 ( .A(u3__abc_46775_n876), .B(u3__abc_46775_n891), .Y(u3__abc_46775_n894) );
  OR2X2 OR2X2_4296 ( .A(u3_rd_fifo_out_22_), .B(u3_rd_fifo_out_23_), .Y(u3__abc_46775_n897) );
  OR2X2 OR2X2_4297 ( .A(u3_rd_fifo_out_16_), .B(u3_rd_fifo_out_17_), .Y(u3__abc_46775_n903) );
  OR2X2 OR2X2_4298 ( .A(u3__abc_46775_n906), .B(u3__abc_46775_n902), .Y(u3__abc_46775_n907) );
  OR2X2 OR2X2_4299 ( .A(u3__abc_46775_n910), .B(u3__abc_46775_n904), .Y(u3__abc_46775_n911) );
  OR2X2 OR2X2_43 ( .A(_abc_55805_n240_bF_buf5), .B(sp_tms_4_), .Y(_abc_55805_n302) );
  OR2X2 OR2X2_430 ( .A(spec_req_cs_6_bF_buf2), .B(1'b0), .Y(u0__abc_49347_n2029) );
  OR2X2 OR2X2_4300 ( .A(u3__abc_46775_n911), .B(u3_rd_fifo_out_34_), .Y(u3__abc_46775_n912) );
  OR2X2 OR2X2_4301 ( .A(u3__abc_46775_n913), .B(u3__abc_46775_n901), .Y(u3__abc_46775_n914) );
  OR2X2 OR2X2_4302 ( .A(u3__abc_46775_n915), .B(u3__abc_46775_n916), .Y(u3__abc_46775_n917) );
  OR2X2 OR2X2_4303 ( .A(u3__abc_46775_n917), .B(u3__abc_46775_n900), .Y(u3__abc_46775_n918) );
  OR2X2 OR2X2_4304 ( .A(u3_rd_fifo_out_20_), .B(u3_rd_fifo_out_21_), .Y(u3__abc_46775_n921) );
  OR2X2 OR2X2_4305 ( .A(u3__abc_46775_n926), .B(u3_rd_fifo_out_18_), .Y(u3__abc_46775_n929) );
  OR2X2 OR2X2_4306 ( .A(u3__abc_46775_n932), .B(u3__abc_46775_n933), .Y(u3__abc_46775_n934) );
  OR2X2 OR2X2_4307 ( .A(u3__abc_46775_n920), .B(u3__abc_46775_n935), .Y(u3__abc_46775_n936) );
  OR2X2 OR2X2_4308 ( .A(u3__abc_46775_n919), .B(u3__abc_46775_n934), .Y(u3__abc_46775_n937) );
  OR2X2 OR2X2_4309 ( .A(u3__abc_46775_n896), .B(u3__abc_46775_n939), .Y(u3__abc_46775_n940) );
  OR2X2 OR2X2_431 ( .A(u0__abc_49347_n2031), .B(u0__abc_49347_n2027), .Y(u0__abc_49347_n2032) );
  OR2X2 OR2X2_4310 ( .A(u3_rd_fifo_out_6_), .B(u3_rd_fifo_out_7_), .Y(u3__abc_46775_n941) );
  OR2X2 OR2X2_4311 ( .A(u3_rd_fifo_out_0_), .B(u3_rd_fifo_out_1_), .Y(u3__abc_46775_n947) );
  OR2X2 OR2X2_4312 ( .A(u3__abc_46775_n950), .B(u3__abc_46775_n946), .Y(u3__abc_46775_n951) );
  OR2X2 OR2X2_4313 ( .A(u3__abc_46775_n954), .B(u3__abc_46775_n948), .Y(u3__abc_46775_n955) );
  OR2X2 OR2X2_4314 ( .A(u3__abc_46775_n955), .B(u3_rd_fifo_out_32_), .Y(u3__abc_46775_n956) );
  OR2X2 OR2X2_4315 ( .A(u3__abc_46775_n957), .B(u3__abc_46775_n945), .Y(u3__abc_46775_n958) );
  OR2X2 OR2X2_4316 ( .A(u3__abc_46775_n959), .B(u3__abc_46775_n960), .Y(u3__abc_46775_n961) );
  OR2X2 OR2X2_4317 ( .A(u3__abc_46775_n961), .B(u3__abc_46775_n944), .Y(u3__abc_46775_n962) );
  OR2X2 OR2X2_4318 ( .A(u3_rd_fifo_out_4_), .B(u3_rd_fifo_out_5_), .Y(u3__abc_46775_n965) );
  OR2X2 OR2X2_4319 ( .A(u3__abc_46775_n970), .B(u3_rd_fifo_out_2_), .Y(u3__abc_46775_n973) );
  OR2X2 OR2X2_432 ( .A(u0__abc_49347_n2033), .B(u0__abc_49347_n2034), .Y(u0__abc_49347_n2035) );
  OR2X2 OR2X2_4320 ( .A(u3__abc_46775_n976), .B(u3__abc_46775_n977), .Y(u3__abc_46775_n978) );
  OR2X2 OR2X2_4321 ( .A(u3__abc_46775_n964), .B(u3__abc_46775_n979), .Y(u3__abc_46775_n980) );
  OR2X2 OR2X2_4322 ( .A(u3__abc_46775_n963), .B(u3__abc_46775_n978), .Y(u3__abc_46775_n981) );
  OR2X2 OR2X2_4323 ( .A(u3_rd_fifo_out_30_), .B(u3_rd_fifo_out_31_), .Y(u3__abc_46775_n984) );
  OR2X2 OR2X2_4324 ( .A(u3_rd_fifo_out_24_), .B(u3_rd_fifo_out_25_), .Y(u3__abc_46775_n990) );
  OR2X2 OR2X2_4325 ( .A(u3__abc_46775_n993), .B(u3__abc_46775_n989), .Y(u3__abc_46775_n994) );
  OR2X2 OR2X2_4326 ( .A(u3__abc_46775_n995), .B(u3_rd_fifo_out_25_), .Y(u3__abc_46775_n996) );
  OR2X2 OR2X2_4327 ( .A(u3__abc_46775_n997), .B(u3_rd_fifo_out_24_), .Y(u3__abc_46775_n998) );
  OR2X2 OR2X2_4328 ( .A(u3__abc_46775_n999), .B(u3_rd_fifo_out_35_), .Y(u3__abc_46775_n1000) );
  OR2X2 OR2X2_4329 ( .A(u3__abc_46775_n1001), .B(u3__abc_46775_n988), .Y(u3__abc_46775_n1002) );
  OR2X2 OR2X2_433 ( .A(u0__abc_49347_n2036), .B(u0__abc_49347_n2037), .Y(u0__abc_49347_n2038) );
  OR2X2 OR2X2_4330 ( .A(u3__abc_46775_n1003), .B(u3__abc_46775_n1004), .Y(u3__abc_46775_n1005) );
  OR2X2 OR2X2_4331 ( .A(u3__abc_46775_n1005), .B(u3__abc_46775_n987), .Y(u3__abc_46775_n1006) );
  OR2X2 OR2X2_4332 ( .A(u3_rd_fifo_out_28_), .B(u3_rd_fifo_out_29_), .Y(u3__abc_46775_n1009) );
  OR2X2 OR2X2_4333 ( .A(u3__abc_46775_n1014), .B(u3_rd_fifo_out_26_), .Y(u3__abc_46775_n1017) );
  OR2X2 OR2X2_4334 ( .A(u3__abc_46775_n1020), .B(u3__abc_46775_n1021), .Y(u3__abc_46775_n1022) );
  OR2X2 OR2X2_4335 ( .A(u3__abc_46775_n1008), .B(u3__abc_46775_n1023), .Y(u3__abc_46775_n1024) );
  OR2X2 OR2X2_4336 ( .A(u3__abc_46775_n1007), .B(u3__abc_46775_n1022), .Y(u3__abc_46775_n1025) );
  OR2X2 OR2X2_4337 ( .A(u3__abc_46775_n983), .B(u3__abc_46775_n1027), .Y(u3__abc_46775_n1028) );
  OR2X2 OR2X2_4338 ( .A(u3__abc_46775_n940), .B(u3__abc_46775_n1028), .Y(u3__abc_46775_n1029) );
  OR2X2 OR2X2_4339 ( .A(u3_u0__abc_48231_n382_bF_buf7), .B(u3_u0_r3_0_), .Y(u3_u0__abc_48231_n383) );
  OR2X2 OR2X2_434 ( .A(u0__abc_49347_n2039), .B(u0__abc_49347_n2040), .Y(u0__abc_49347_n2041) );
  OR2X2 OR2X2_4340 ( .A(u3_u0__abc_48231_n382_bF_buf5), .B(u3_u0_r3_1_), .Y(u3_u0__abc_48231_n388_1) );
  OR2X2 OR2X2_4341 ( .A(u3_u0__abc_48231_n382_bF_buf3), .B(u3_u0_r3_2_), .Y(u3_u0__abc_48231_n393) );
  OR2X2 OR2X2_4342 ( .A(u3_u0__abc_48231_n382_bF_buf1), .B(u3_u0_r3_3_), .Y(u3_u0__abc_48231_n398) );
  OR2X2 OR2X2_4343 ( .A(u3_u0__abc_48231_n382_bF_buf7), .B(u3_u0_r3_4_), .Y(u3_u0__abc_48231_n403) );
  OR2X2 OR2X2_4344 ( .A(u3_u0__abc_48231_n382_bF_buf5), .B(u3_u0_r3_5_), .Y(u3_u0__abc_48231_n408_1) );
  OR2X2 OR2X2_4345 ( .A(u3_u0__abc_48231_n382_bF_buf3), .B(u3_u0_r3_6_), .Y(u3_u0__abc_48231_n413) );
  OR2X2 OR2X2_4346 ( .A(u3_u0__abc_48231_n382_bF_buf1), .B(u3_u0_r3_7_), .Y(u3_u0__abc_48231_n418) );
  OR2X2 OR2X2_4347 ( .A(u3_u0__abc_48231_n382_bF_buf7), .B(u3_u0_r3_8_), .Y(u3_u0__abc_48231_n423) );
  OR2X2 OR2X2_4348 ( .A(u3_u0__abc_48231_n382_bF_buf5), .B(u3_u0_r3_9_), .Y(u3_u0__abc_48231_n428_1) );
  OR2X2 OR2X2_4349 ( .A(u3_u0__abc_48231_n382_bF_buf3), .B(u3_u0_r3_10_), .Y(u3_u0__abc_48231_n433) );
  OR2X2 OR2X2_435 ( .A(u0__abc_49347_n2043), .B(spec_req_cs_0_bF_buf2), .Y(u0__abc_49347_n2044) );
  OR2X2 OR2X2_4350 ( .A(u3_u0__abc_48231_n382_bF_buf1), .B(u3_u0_r3_11_), .Y(u3_u0__abc_48231_n438) );
  OR2X2 OR2X2_4351 ( .A(u3_u0__abc_48231_n382_bF_buf7), .B(u3_u0_r3_12_), .Y(u3_u0__abc_48231_n443) );
  OR2X2 OR2X2_4352 ( .A(u3_u0__abc_48231_n382_bF_buf5), .B(u3_u0_r3_13_), .Y(u3_u0__abc_48231_n448_1) );
  OR2X2 OR2X2_4353 ( .A(u3_u0__abc_48231_n382_bF_buf3), .B(u3_u0_r3_14_), .Y(u3_u0__abc_48231_n453) );
  OR2X2 OR2X2_4354 ( .A(u3_u0__abc_48231_n382_bF_buf1), .B(u3_u0_r3_15_), .Y(u3_u0__abc_48231_n458) );
  OR2X2 OR2X2_4355 ( .A(u3_u0__abc_48231_n382_bF_buf7), .B(u3_u0_r3_16_), .Y(u3_u0__abc_48231_n463) );
  OR2X2 OR2X2_4356 ( .A(u3_u0__abc_48231_n382_bF_buf5), .B(u3_u0_r3_17_), .Y(u3_u0__abc_48231_n468_1) );
  OR2X2 OR2X2_4357 ( .A(u3_u0__abc_48231_n382_bF_buf3), .B(u3_u0_r3_18_), .Y(u3_u0__abc_48231_n473) );
  OR2X2 OR2X2_4358 ( .A(u3_u0__abc_48231_n382_bF_buf1), .B(u3_u0_r3_19_), .Y(u3_u0__abc_48231_n478) );
  OR2X2 OR2X2_4359 ( .A(u3_u0__abc_48231_n382_bF_buf7), .B(u3_u0_r3_20_), .Y(u3_u0__abc_48231_n483) );
  OR2X2 OR2X2_436 ( .A(u0__abc_49347_n2042), .B(u0__abc_49347_n2044), .Y(u0__abc_49347_n2045) );
  OR2X2 OR2X2_4360 ( .A(u3_u0__abc_48231_n382_bF_buf5), .B(u3_u0_r3_21_), .Y(u3_u0__abc_48231_n488_1) );
  OR2X2 OR2X2_4361 ( .A(u3_u0__abc_48231_n382_bF_buf3), .B(u3_u0_r3_22_), .Y(u3_u0__abc_48231_n493) );
  OR2X2 OR2X2_4362 ( .A(u3_u0__abc_48231_n382_bF_buf1), .B(u3_u0_r3_23_), .Y(u3_u0__abc_48231_n498) );
  OR2X2 OR2X2_4363 ( .A(u3_u0__abc_48231_n382_bF_buf7), .B(u3_u0_r3_24_), .Y(u3_u0__abc_48231_n503) );
  OR2X2 OR2X2_4364 ( .A(u3_u0__abc_48231_n382_bF_buf5), .B(u3_u0_r3_25_), .Y(u3_u0__abc_48231_n508_1) );
  OR2X2 OR2X2_4365 ( .A(u3_u0__abc_48231_n382_bF_buf3), .B(u3_u0_r3_26_), .Y(u3_u0__abc_48231_n513_1) );
  OR2X2 OR2X2_4366 ( .A(u3_u0__abc_48231_n382_bF_buf1), .B(u3_u0_r3_27_), .Y(u3_u0__abc_48231_n518) );
  OR2X2 OR2X2_4367 ( .A(u3_u0__abc_48231_n382_bF_buf7), .B(u3_u0_r3_28_), .Y(u3_u0__abc_48231_n523) );
  OR2X2 OR2X2_4368 ( .A(u3_u0__abc_48231_n382_bF_buf5), .B(u3_u0_r3_29_), .Y(u3_u0__abc_48231_n528) );
  OR2X2 OR2X2_4369 ( .A(u3_u0__abc_48231_n382_bF_buf3), .B(u3_u0_r3_30_), .Y(u3_u0__abc_48231_n533) );
  OR2X2 OR2X2_437 ( .A(u0__abc_49347_n1203_bF_buf5), .B(u0_csc0_3_), .Y(u0__abc_49347_n2046) );
  OR2X2 OR2X2_4370 ( .A(u3_u0__abc_48231_n382_bF_buf1), .B(u3_u0_r3_31_), .Y(u3_u0__abc_48231_n538) );
  OR2X2 OR2X2_4371 ( .A(u3_u0__abc_48231_n382_bF_buf7), .B(u3_u0_r3_32_), .Y(u3_u0__abc_48231_n543) );
  OR2X2 OR2X2_4372 ( .A(u3_u0__abc_48231_n382_bF_buf5), .B(u3_u0_r3_33_), .Y(u3_u0__abc_48231_n548) );
  OR2X2 OR2X2_4373 ( .A(u3_u0__abc_48231_n382_bF_buf3), .B(u3_u0_r3_34_), .Y(u3_u0__abc_48231_n553) );
  OR2X2 OR2X2_4374 ( .A(u3_u0__abc_48231_n382_bF_buf1), .B(u3_u0_r3_35_), .Y(u3_u0__abc_48231_n558) );
  OR2X2 OR2X2_4375 ( .A(u3_u0__abc_48231_n563_bF_buf7), .B(u3_u0_r2_0_), .Y(u3_u0__abc_48231_n564) );
  OR2X2 OR2X2_4376 ( .A(u3_u0__abc_48231_n563_bF_buf5), .B(u3_u0_r2_1_), .Y(u3_u0__abc_48231_n568) );
  OR2X2 OR2X2_4377 ( .A(u3_u0__abc_48231_n563_bF_buf3), .B(u3_u0_r2_2_), .Y(u3_u0__abc_48231_n572) );
  OR2X2 OR2X2_4378 ( .A(u3_u0__abc_48231_n563_bF_buf1), .B(u3_u0_r2_3_), .Y(u3_u0__abc_48231_n576) );
  OR2X2 OR2X2_4379 ( .A(u3_u0__abc_48231_n563_bF_buf7), .B(u3_u0_r2_4_), .Y(u3_u0__abc_48231_n580) );
  OR2X2 OR2X2_438 ( .A(u0__abc_49347_n2048), .B(u0__abc_49347_n2026), .Y(u0_sp_csc_3__FF_INPUT) );
  OR2X2 OR2X2_4380 ( .A(u3_u0__abc_48231_n563_bF_buf5), .B(u3_u0_r2_5_), .Y(u3_u0__abc_48231_n584) );
  OR2X2 OR2X2_4381 ( .A(u3_u0__abc_48231_n563_bF_buf3), .B(u3_u0_r2_6_), .Y(u3_u0__abc_48231_n588) );
  OR2X2 OR2X2_4382 ( .A(u3_u0__abc_48231_n563_bF_buf1), .B(u3_u0_r2_7_), .Y(u3_u0__abc_48231_n592) );
  OR2X2 OR2X2_4383 ( .A(u3_u0__abc_48231_n563_bF_buf7), .B(u3_u0_r2_8_), .Y(u3_u0__abc_48231_n596) );
  OR2X2 OR2X2_4384 ( .A(u3_u0__abc_48231_n563_bF_buf5), .B(u3_u0_r2_9_), .Y(u3_u0__abc_48231_n600) );
  OR2X2 OR2X2_4385 ( .A(u3_u0__abc_48231_n563_bF_buf3), .B(u3_u0_r2_10_), .Y(u3_u0__abc_48231_n604) );
  OR2X2 OR2X2_4386 ( .A(u3_u0__abc_48231_n563_bF_buf1), .B(u3_u0_r2_11_), .Y(u3_u0__abc_48231_n608) );
  OR2X2 OR2X2_4387 ( .A(u3_u0__abc_48231_n563_bF_buf7), .B(u3_u0_r2_12_), .Y(u3_u0__abc_48231_n612) );
  OR2X2 OR2X2_4388 ( .A(u3_u0__abc_48231_n563_bF_buf5), .B(u3_u0_r2_13_), .Y(u3_u0__abc_48231_n616) );
  OR2X2 OR2X2_4389 ( .A(u3_u0__abc_48231_n563_bF_buf3), .B(u3_u0_r2_14_), .Y(u3_u0__abc_48231_n620) );
  OR2X2 OR2X2_439 ( .A(u0__abc_49347_n1183_1_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n2052) );
  OR2X2 OR2X2_4390 ( .A(u3_u0__abc_48231_n563_bF_buf1), .B(u3_u0_r2_15_), .Y(u3_u0__abc_48231_n624) );
  OR2X2 OR2X2_4391 ( .A(u3_u0__abc_48231_n563_bF_buf7), .B(u3_u0_r2_16_), .Y(u3_u0__abc_48231_n628) );
  OR2X2 OR2X2_4392 ( .A(u3_u0__abc_48231_n563_bF_buf5), .B(u3_u0_r2_17_), .Y(u3_u0__abc_48231_n632) );
  OR2X2 OR2X2_4393 ( .A(u3_u0__abc_48231_n563_bF_buf3), .B(u3_u0_r2_18_), .Y(u3_u0__abc_48231_n636) );
  OR2X2 OR2X2_4394 ( .A(u3_u0__abc_48231_n563_bF_buf1), .B(u3_u0_r2_19_), .Y(u3_u0__abc_48231_n640) );
  OR2X2 OR2X2_4395 ( .A(u3_u0__abc_48231_n563_bF_buf7), .B(u3_u0_r2_20_), .Y(u3_u0__abc_48231_n644) );
  OR2X2 OR2X2_4396 ( .A(u3_u0__abc_48231_n563_bF_buf5), .B(u3_u0_r2_21_), .Y(u3_u0__abc_48231_n648) );
  OR2X2 OR2X2_4397 ( .A(u3_u0__abc_48231_n563_bF_buf3), .B(u3_u0_r2_22_), .Y(u3_u0__abc_48231_n652) );
  OR2X2 OR2X2_4398 ( .A(u3_u0__abc_48231_n563_bF_buf1), .B(u3_u0_r2_23_), .Y(u3_u0__abc_48231_n656) );
  OR2X2 OR2X2_4399 ( .A(u3_u0__abc_48231_n563_bF_buf7), .B(u3_u0_r2_24_), .Y(u3_u0__abc_48231_n660) );
  OR2X2 OR2X2_44 ( .A(lmr_sel_bF_buf1), .B(tms_4_), .Y(_abc_55805_n303) );
  OR2X2 OR2X2_440 ( .A(spec_req_cs_6_bF_buf1), .B(1'b0), .Y(u0__abc_49347_n2053) );
  OR2X2 OR2X2_4400 ( .A(u3_u0__abc_48231_n563_bF_buf5), .B(u3_u0_r2_25_), .Y(u3_u0__abc_48231_n664) );
  OR2X2 OR2X2_4401 ( .A(u3_u0__abc_48231_n563_bF_buf3), .B(u3_u0_r2_26_), .Y(u3_u0__abc_48231_n668) );
  OR2X2 OR2X2_4402 ( .A(u3_u0__abc_48231_n563_bF_buf1), .B(u3_u0_r2_27_), .Y(u3_u0__abc_48231_n672) );
  OR2X2 OR2X2_4403 ( .A(u3_u0__abc_48231_n563_bF_buf7), .B(u3_u0_r2_28_), .Y(u3_u0__abc_48231_n676) );
  OR2X2 OR2X2_4404 ( .A(u3_u0__abc_48231_n563_bF_buf5), .B(u3_u0_r2_29_), .Y(u3_u0__abc_48231_n680) );
  OR2X2 OR2X2_4405 ( .A(u3_u0__abc_48231_n563_bF_buf3), .B(u3_u0_r2_30_), .Y(u3_u0__abc_48231_n684) );
  OR2X2 OR2X2_4406 ( .A(u3_u0__abc_48231_n563_bF_buf1), .B(u3_u0_r2_31_), .Y(u3_u0__abc_48231_n688) );
  OR2X2 OR2X2_4407 ( .A(u3_u0__abc_48231_n563_bF_buf7), .B(u3_u0_r2_32_), .Y(u3_u0__abc_48231_n692) );
  OR2X2 OR2X2_4408 ( .A(u3_u0__abc_48231_n563_bF_buf5), .B(u3_u0_r2_33_), .Y(u3_u0__abc_48231_n696) );
  OR2X2 OR2X2_4409 ( .A(u3_u0__abc_48231_n563_bF_buf3), .B(u3_u0_r2_34_), .Y(u3_u0__abc_48231_n700) );
  OR2X2 OR2X2_441 ( .A(u0__abc_49347_n2055), .B(u0__abc_49347_n2051_1), .Y(u0__abc_49347_n2056) );
  OR2X2 OR2X2_4410 ( .A(u3_u0__abc_48231_n563_bF_buf1), .B(u3_u0_r2_35_), .Y(u3_u0__abc_48231_n704) );
  OR2X2 OR2X2_4411 ( .A(u3_u0__abc_48231_n708_bF_buf7), .B(u3_u0_r1_0_), .Y(u3_u0__abc_48231_n709) );
  OR2X2 OR2X2_4412 ( .A(u3_u0__abc_48231_n708_bF_buf5), .B(u3_u0_r1_1_), .Y(u3_u0__abc_48231_n713) );
  OR2X2 OR2X2_4413 ( .A(u3_u0__abc_48231_n708_bF_buf3), .B(u3_u0_r1_2_), .Y(u3_u0__abc_48231_n717) );
  OR2X2 OR2X2_4414 ( .A(u3_u0__abc_48231_n708_bF_buf1), .B(u3_u0_r1_3_), .Y(u3_u0__abc_48231_n721) );
  OR2X2 OR2X2_4415 ( .A(u3_u0__abc_48231_n708_bF_buf7), .B(u3_u0_r1_4_), .Y(u3_u0__abc_48231_n725) );
  OR2X2 OR2X2_4416 ( .A(u3_u0__abc_48231_n708_bF_buf5), .B(u3_u0_r1_5_), .Y(u3_u0__abc_48231_n729) );
  OR2X2 OR2X2_4417 ( .A(u3_u0__abc_48231_n708_bF_buf3), .B(u3_u0_r1_6_), .Y(u3_u0__abc_48231_n733) );
  OR2X2 OR2X2_4418 ( .A(u3_u0__abc_48231_n708_bF_buf1), .B(u3_u0_r1_7_), .Y(u3_u0__abc_48231_n737) );
  OR2X2 OR2X2_4419 ( .A(u3_u0__abc_48231_n708_bF_buf7), .B(u3_u0_r1_8_), .Y(u3_u0__abc_48231_n741) );
  OR2X2 OR2X2_442 ( .A(u0__abc_49347_n2057), .B(u0__abc_49347_n2058), .Y(u0__abc_49347_n2059) );
  OR2X2 OR2X2_4420 ( .A(u3_u0__abc_48231_n708_bF_buf5), .B(u3_u0_r1_9_), .Y(u3_u0__abc_48231_n745) );
  OR2X2 OR2X2_4421 ( .A(u3_u0__abc_48231_n708_bF_buf3), .B(u3_u0_r1_10_), .Y(u3_u0__abc_48231_n749) );
  OR2X2 OR2X2_4422 ( .A(u3_u0__abc_48231_n708_bF_buf1), .B(u3_u0_r1_11_), .Y(u3_u0__abc_48231_n753) );
  OR2X2 OR2X2_4423 ( .A(u3_u0__abc_48231_n708_bF_buf7), .B(u3_u0_r1_12_), .Y(u3_u0__abc_48231_n757) );
  OR2X2 OR2X2_4424 ( .A(u3_u0__abc_48231_n708_bF_buf5), .B(u3_u0_r1_13_), .Y(u3_u0__abc_48231_n761) );
  OR2X2 OR2X2_4425 ( .A(u3_u0__abc_48231_n708_bF_buf3), .B(u3_u0_r1_14_), .Y(u3_u0__abc_48231_n765) );
  OR2X2 OR2X2_4426 ( .A(u3_u0__abc_48231_n708_bF_buf1), .B(u3_u0_r1_15_), .Y(u3_u0__abc_48231_n769) );
  OR2X2 OR2X2_4427 ( .A(u3_u0__abc_48231_n708_bF_buf7), .B(u3_u0_r1_16_), .Y(u3_u0__abc_48231_n773) );
  OR2X2 OR2X2_4428 ( .A(u3_u0__abc_48231_n708_bF_buf5), .B(u3_u0_r1_17_), .Y(u3_u0__abc_48231_n777) );
  OR2X2 OR2X2_4429 ( .A(u3_u0__abc_48231_n708_bF_buf3), .B(u3_u0_r1_18_), .Y(u3_u0__abc_48231_n781) );
  OR2X2 OR2X2_443 ( .A(u0__abc_49347_n2060), .B(u0__abc_49347_n2061), .Y(u0__abc_49347_n2062) );
  OR2X2 OR2X2_4430 ( .A(u3_u0__abc_48231_n708_bF_buf1), .B(u3_u0_r1_19_), .Y(u3_u0__abc_48231_n785) );
  OR2X2 OR2X2_4431 ( .A(u3_u0__abc_48231_n708_bF_buf7), .B(u3_u0_r1_20_), .Y(u3_u0__abc_48231_n789) );
  OR2X2 OR2X2_4432 ( .A(u3_u0__abc_48231_n708_bF_buf5), .B(u3_u0_r1_21_), .Y(u3_u0__abc_48231_n793) );
  OR2X2 OR2X2_4433 ( .A(u3_u0__abc_48231_n708_bF_buf3), .B(u3_u0_r1_22_), .Y(u3_u0__abc_48231_n797) );
  OR2X2 OR2X2_4434 ( .A(u3_u0__abc_48231_n708_bF_buf1), .B(u3_u0_r1_23_), .Y(u3_u0__abc_48231_n801) );
  OR2X2 OR2X2_4435 ( .A(u3_u0__abc_48231_n708_bF_buf7), .B(u3_u0_r1_24_), .Y(u3_u0__abc_48231_n805) );
  OR2X2 OR2X2_4436 ( .A(u3_u0__abc_48231_n708_bF_buf5), .B(u3_u0_r1_25_), .Y(u3_u0__abc_48231_n809) );
  OR2X2 OR2X2_4437 ( .A(u3_u0__abc_48231_n708_bF_buf3), .B(u3_u0_r1_26_), .Y(u3_u0__abc_48231_n813) );
  OR2X2 OR2X2_4438 ( .A(u3_u0__abc_48231_n708_bF_buf1), .B(u3_u0_r1_27_), .Y(u3_u0__abc_48231_n817) );
  OR2X2 OR2X2_4439 ( .A(u3_u0__abc_48231_n708_bF_buf7), .B(u3_u0_r1_28_), .Y(u3_u0__abc_48231_n821) );
  OR2X2 OR2X2_444 ( .A(u0__abc_49347_n2063), .B(u0__abc_49347_n2064), .Y(u0__abc_49347_n2065) );
  OR2X2 OR2X2_4440 ( .A(u3_u0__abc_48231_n708_bF_buf5), .B(u3_u0_r1_29_), .Y(u3_u0__abc_48231_n825) );
  OR2X2 OR2X2_4441 ( .A(u3_u0__abc_48231_n708_bF_buf3), .B(u3_u0_r1_30_), .Y(u3_u0__abc_48231_n829) );
  OR2X2 OR2X2_4442 ( .A(u3_u0__abc_48231_n708_bF_buf1), .B(u3_u0_r1_31_), .Y(u3_u0__abc_48231_n833) );
  OR2X2 OR2X2_4443 ( .A(u3_u0__abc_48231_n708_bF_buf7), .B(u3_u0_r1_32_), .Y(u3_u0__abc_48231_n837) );
  OR2X2 OR2X2_4444 ( .A(u3_u0__abc_48231_n708_bF_buf5), .B(u3_u0_r1_33_), .Y(u3_u0__abc_48231_n841) );
  OR2X2 OR2X2_4445 ( .A(u3_u0__abc_48231_n708_bF_buf3), .B(u3_u0_r1_34_), .Y(u3_u0__abc_48231_n845) );
  OR2X2 OR2X2_4446 ( .A(u3_u0__abc_48231_n708_bF_buf1), .B(u3_u0_r1_35_), .Y(u3_u0__abc_48231_n849) );
  OR2X2 OR2X2_4447 ( .A(u3_u0__abc_48231_n853_bF_buf7), .B(u3_u0_r0_0_), .Y(u3_u0__abc_48231_n854) );
  OR2X2 OR2X2_4448 ( .A(u3_u0__abc_48231_n853_bF_buf5), .B(u3_u0_r0_1_), .Y(u3_u0__abc_48231_n858) );
  OR2X2 OR2X2_4449 ( .A(u3_u0__abc_48231_n853_bF_buf3), .B(u3_u0_r0_2_), .Y(u3_u0__abc_48231_n862) );
  OR2X2 OR2X2_445 ( .A(u0__abc_49347_n2067), .B(spec_req_cs_0_bF_buf1), .Y(u0__abc_49347_n2068) );
  OR2X2 OR2X2_4450 ( .A(u3_u0__abc_48231_n853_bF_buf1), .B(u3_u0_r0_3_), .Y(u3_u0__abc_48231_n866) );
  OR2X2 OR2X2_4451 ( .A(u3_u0__abc_48231_n853_bF_buf7), .B(u3_u0_r0_4_), .Y(u3_u0__abc_48231_n870) );
  OR2X2 OR2X2_4452 ( .A(u3_u0__abc_48231_n853_bF_buf5), .B(u3_u0_r0_5_), .Y(u3_u0__abc_48231_n874) );
  OR2X2 OR2X2_4453 ( .A(u3_u0__abc_48231_n853_bF_buf3), .B(u3_u0_r0_6_), .Y(u3_u0__abc_48231_n878) );
  OR2X2 OR2X2_4454 ( .A(u3_u0__abc_48231_n853_bF_buf1), .B(u3_u0_r0_7_), .Y(u3_u0__abc_48231_n882) );
  OR2X2 OR2X2_4455 ( .A(u3_u0__abc_48231_n853_bF_buf7), .B(u3_u0_r0_8_), .Y(u3_u0__abc_48231_n886) );
  OR2X2 OR2X2_4456 ( .A(u3_u0__abc_48231_n853_bF_buf5), .B(u3_u0_r0_9_), .Y(u3_u0__abc_48231_n890) );
  OR2X2 OR2X2_4457 ( .A(u3_u0__abc_48231_n853_bF_buf3), .B(u3_u0_r0_10_), .Y(u3_u0__abc_48231_n894) );
  OR2X2 OR2X2_4458 ( .A(u3_u0__abc_48231_n853_bF_buf1), .B(u3_u0_r0_11_), .Y(u3_u0__abc_48231_n898) );
  OR2X2 OR2X2_4459 ( .A(u3_u0__abc_48231_n853_bF_buf7), .B(u3_u0_r0_12_), .Y(u3_u0__abc_48231_n902) );
  OR2X2 OR2X2_446 ( .A(u0__abc_49347_n2066), .B(u0__abc_49347_n2068), .Y(u0__abc_49347_n2069) );
  OR2X2 OR2X2_4460 ( .A(u3_u0__abc_48231_n853_bF_buf5), .B(u3_u0_r0_13_), .Y(u3_u0__abc_48231_n906) );
  OR2X2 OR2X2_4461 ( .A(u3_u0__abc_48231_n853_bF_buf3), .B(u3_u0_r0_14_), .Y(u3_u0__abc_48231_n910) );
  OR2X2 OR2X2_4462 ( .A(u3_u0__abc_48231_n853_bF_buf1), .B(u3_u0_r0_15_), .Y(u3_u0__abc_48231_n914) );
  OR2X2 OR2X2_4463 ( .A(u3_u0__abc_48231_n853_bF_buf7), .B(u3_u0_r0_16_), .Y(u3_u0__abc_48231_n918) );
  OR2X2 OR2X2_4464 ( .A(u3_u0__abc_48231_n853_bF_buf5), .B(u3_u0_r0_17_), .Y(u3_u0__abc_48231_n922) );
  OR2X2 OR2X2_4465 ( .A(u3_u0__abc_48231_n853_bF_buf3), .B(u3_u0_r0_18_), .Y(u3_u0__abc_48231_n926) );
  OR2X2 OR2X2_4466 ( .A(u3_u0__abc_48231_n853_bF_buf1), .B(u3_u0_r0_19_), .Y(u3_u0__abc_48231_n930) );
  OR2X2 OR2X2_4467 ( .A(u3_u0__abc_48231_n853_bF_buf7), .B(u3_u0_r0_20_), .Y(u3_u0__abc_48231_n934) );
  OR2X2 OR2X2_4468 ( .A(u3_u0__abc_48231_n853_bF_buf5), .B(u3_u0_r0_21_), .Y(u3_u0__abc_48231_n938) );
  OR2X2 OR2X2_4469 ( .A(u3_u0__abc_48231_n853_bF_buf3), .B(u3_u0_r0_22_), .Y(u3_u0__abc_48231_n942) );
  OR2X2 OR2X2_447 ( .A(u0__abc_49347_n1203_bF_buf4), .B(u0_csc0_4_), .Y(u0__abc_49347_n2070) );
  OR2X2 OR2X2_4470 ( .A(u3_u0__abc_48231_n853_bF_buf1), .B(u3_u0_r0_23_), .Y(u3_u0__abc_48231_n946) );
  OR2X2 OR2X2_4471 ( .A(u3_u0__abc_48231_n853_bF_buf7), .B(u3_u0_r0_24_), .Y(u3_u0__abc_48231_n950) );
  OR2X2 OR2X2_4472 ( .A(u3_u0__abc_48231_n853_bF_buf5), .B(u3_u0_r0_25_), .Y(u3_u0__abc_48231_n954) );
  OR2X2 OR2X2_4473 ( .A(u3_u0__abc_48231_n853_bF_buf3), .B(u3_u0_r0_26_), .Y(u3_u0__abc_48231_n958) );
  OR2X2 OR2X2_4474 ( .A(u3_u0__abc_48231_n853_bF_buf1), .B(u3_u0_r0_27_), .Y(u3_u0__abc_48231_n962) );
  OR2X2 OR2X2_4475 ( .A(u3_u0__abc_48231_n853_bF_buf7), .B(u3_u0_r0_28_), .Y(u3_u0__abc_48231_n966) );
  OR2X2 OR2X2_4476 ( .A(u3_u0__abc_48231_n853_bF_buf5), .B(u3_u0_r0_29_), .Y(u3_u0__abc_48231_n970) );
  OR2X2 OR2X2_4477 ( .A(u3_u0__abc_48231_n853_bF_buf3), .B(u3_u0_r0_30_), .Y(u3_u0__abc_48231_n974) );
  OR2X2 OR2X2_4478 ( .A(u3_u0__abc_48231_n853_bF_buf1), .B(u3_u0_r0_31_), .Y(u3_u0__abc_48231_n978) );
  OR2X2 OR2X2_4479 ( .A(u3_u0__abc_48231_n853_bF_buf7), .B(u3_u0_r0_32_), .Y(u3_u0__abc_48231_n982) );
  OR2X2 OR2X2_448 ( .A(u0__abc_49347_n2072_1), .B(u0__abc_49347_n2050), .Y(u0_sp_csc_4__FF_INPUT) );
  OR2X2 OR2X2_4480 ( .A(u3_u0__abc_48231_n853_bF_buf5), .B(u3_u0_r0_33_), .Y(u3_u0__abc_48231_n986) );
  OR2X2 OR2X2_4481 ( .A(u3_u0__abc_48231_n853_bF_buf3), .B(u3_u0_r0_34_), .Y(u3_u0__abc_48231_n990) );
  OR2X2 OR2X2_4482 ( .A(u3_u0__abc_48231_n853_bF_buf1), .B(u3_u0_r0_35_), .Y(u3_u0__abc_48231_n994) );
  OR2X2 OR2X2_4483 ( .A(u3_u0__abc_48231_n382_bF_buf7), .B(u3_rd_fifo_clr), .Y(u3_u0__abc_48231_n1000) );
  OR2X2 OR2X2_4484 ( .A(u3_u0__abc_48231_n1000), .B(u3_u0__abc_48231_n999), .Y(u3_u0_wr_adr_0__FF_INPUT) );
  OR2X2 OR2X2_4485 ( .A(u3_u0__abc_48231_n1003), .B(u3_u0__abc_48231_n853_bF_buf7), .Y(u3_u0__abc_48231_n1004) );
  OR2X2 OR2X2_4486 ( .A(u3_u0__abc_48231_n1006), .B(u3_u0__abc_48231_n708_bF_buf7), .Y(u3_u0__abc_48231_n1007) );
  OR2X2 OR2X2_4487 ( .A(u3_u0__abc_48231_n1009), .B(u3_u0__abc_48231_n563_bF_buf7), .Y(u3_u0__abc_48231_n1010) );
  OR2X2 OR2X2_4488 ( .A(u3_u0__abc_48231_n1014), .B(u3_rd_fifo_clr), .Y(u3_u0__abc_48231_n1015) );
  OR2X2 OR2X2_4489 ( .A(u3_u0__abc_48231_n1015), .B(u3_u0__abc_48231_n1013), .Y(u3_u0_rd_adr_0__FF_INPUT) );
  OR2X2 OR2X2_449 ( .A(u0__abc_49347_n1183_1_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n2076) );
  OR2X2 OR2X2_4490 ( .A(u3_u0__abc_48231_n1018), .B(u3_u0__abc_48231_n1017), .Y(u3_u0__abc_48231_n1019) );
  OR2X2 OR2X2_4491 ( .A(u3_u0__abc_48231_n1022), .B(u3_u0__abc_48231_n1021), .Y(u3_u0__abc_48231_n1023) );
  OR2X2 OR2X2_4492 ( .A(u3_u0__abc_48231_n1026), .B(u3_u0__abc_48231_n1025), .Y(u3_u0__abc_48231_n1027) );
  OR2X2 OR2X2_4493 ( .A(u3_u0_rd_adr_3_), .B(u3_u0_rd_adr_1_), .Y(u3_u0__abc_48231_n1036) );
  OR2X2 OR2X2_4494 ( .A(u3_u0__abc_48231_n1032), .B(u3_u0_rd_adr_2_), .Y(u3_u0__abc_48231_n1037) );
  OR2X2 OR2X2_4495 ( .A(u3_u0__abc_48231_n1037), .B(u3_u0__abc_48231_n1036), .Y(u3_u0__abc_48231_n1038) );
  OR2X2 OR2X2_4496 ( .A(u3_u0__abc_48231_n1030), .B(u3_u0_rd_adr_0_), .Y(u3_u0__abc_48231_n1039) );
  OR2X2 OR2X2_4497 ( .A(u3_u0__abc_48231_n1039), .B(u3_u0__abc_48231_n1036), .Y(u3_u0__abc_48231_n1040) );
  OR2X2 OR2X2_4498 ( .A(u3_u0__abc_48231_n1051), .B(u3_u0__abc_48231_n1052), .Y(u3_u0__abc_48231_n1053) );
  OR2X2 OR2X2_4499 ( .A(u3_u0__abc_48231_n1053), .B(u3_u0__abc_48231_n1048), .Y(u3_u0__abc_48231_n1054) );
  OR2X2 OR2X2_45 ( .A(_abc_55805_n240_bF_buf4), .B(sp_tms_5_), .Y(_abc_55805_n305) );
  OR2X2 OR2X2_450 ( .A(spec_req_cs_6_bF_buf0), .B(1'b0), .Y(u0__abc_49347_n2077) );
  OR2X2 OR2X2_4500 ( .A(u3_u0__abc_48231_n1054), .B(u3_u0__abc_48231_n1043), .Y(u3_rd_fifo_out_0_) );
  OR2X2 OR2X2_4501 ( .A(u3_u0__abc_48231_n1058), .B(u3_u0__abc_48231_n1059), .Y(u3_u0__abc_48231_n1060) );
  OR2X2 OR2X2_4502 ( .A(u3_u0__abc_48231_n1060), .B(u3_u0__abc_48231_n1057), .Y(u3_u0__abc_48231_n1061) );
  OR2X2 OR2X2_4503 ( .A(u3_u0__abc_48231_n1061), .B(u3_u0__abc_48231_n1056), .Y(u3_rd_fifo_out_1_) );
  OR2X2 OR2X2_4504 ( .A(u3_u0__abc_48231_n1065), .B(u3_u0__abc_48231_n1066), .Y(u3_u0__abc_48231_n1067) );
  OR2X2 OR2X2_4505 ( .A(u3_u0__abc_48231_n1067), .B(u3_u0__abc_48231_n1064), .Y(u3_u0__abc_48231_n1068) );
  OR2X2 OR2X2_4506 ( .A(u3_u0__abc_48231_n1068), .B(u3_u0__abc_48231_n1063), .Y(u3_rd_fifo_out_2_) );
  OR2X2 OR2X2_4507 ( .A(u3_u0__abc_48231_n1072), .B(u3_u0__abc_48231_n1073), .Y(u3_u0__abc_48231_n1074) );
  OR2X2 OR2X2_4508 ( .A(u3_u0__abc_48231_n1074), .B(u3_u0__abc_48231_n1071), .Y(u3_u0__abc_48231_n1075) );
  OR2X2 OR2X2_4509 ( .A(u3_u0__abc_48231_n1075), .B(u3_u0__abc_48231_n1070), .Y(u3_rd_fifo_out_3_) );
  OR2X2 OR2X2_451 ( .A(u0__abc_49347_n2079), .B(u0__abc_49347_n2075), .Y(u0__abc_49347_n2080) );
  OR2X2 OR2X2_4510 ( .A(u3_u0__abc_48231_n1079), .B(u3_u0__abc_48231_n1080), .Y(u3_u0__abc_48231_n1081) );
  OR2X2 OR2X2_4511 ( .A(u3_u0__abc_48231_n1081), .B(u3_u0__abc_48231_n1078), .Y(u3_u0__abc_48231_n1082) );
  OR2X2 OR2X2_4512 ( .A(u3_u0__abc_48231_n1082), .B(u3_u0__abc_48231_n1077), .Y(u3_rd_fifo_out_4_) );
  OR2X2 OR2X2_4513 ( .A(u3_u0__abc_48231_n1086), .B(u3_u0__abc_48231_n1087), .Y(u3_u0__abc_48231_n1088) );
  OR2X2 OR2X2_4514 ( .A(u3_u0__abc_48231_n1088), .B(u3_u0__abc_48231_n1085), .Y(u3_u0__abc_48231_n1089) );
  OR2X2 OR2X2_4515 ( .A(u3_u0__abc_48231_n1089), .B(u3_u0__abc_48231_n1084), .Y(u3_rd_fifo_out_5_) );
  OR2X2 OR2X2_4516 ( .A(u3_u0__abc_48231_n1093), .B(u3_u0__abc_48231_n1094), .Y(u3_u0__abc_48231_n1095) );
  OR2X2 OR2X2_4517 ( .A(u3_u0__abc_48231_n1095), .B(u3_u0__abc_48231_n1092), .Y(u3_u0__abc_48231_n1096) );
  OR2X2 OR2X2_4518 ( .A(u3_u0__abc_48231_n1096), .B(u3_u0__abc_48231_n1091), .Y(u3_rd_fifo_out_6_) );
  OR2X2 OR2X2_4519 ( .A(u3_u0__abc_48231_n1100), .B(u3_u0__abc_48231_n1101), .Y(u3_u0__abc_48231_n1102) );
  OR2X2 OR2X2_452 ( .A(u0__abc_49347_n2081), .B(u0__abc_49347_n2082), .Y(u0__abc_49347_n2083) );
  OR2X2 OR2X2_4520 ( .A(u3_u0__abc_48231_n1102), .B(u3_u0__abc_48231_n1099), .Y(u3_u0__abc_48231_n1103) );
  OR2X2 OR2X2_4521 ( .A(u3_u0__abc_48231_n1103), .B(u3_u0__abc_48231_n1098), .Y(u3_rd_fifo_out_7_) );
  OR2X2 OR2X2_4522 ( .A(u3_u0__abc_48231_n1107), .B(u3_u0__abc_48231_n1108), .Y(u3_u0__abc_48231_n1109) );
  OR2X2 OR2X2_4523 ( .A(u3_u0__abc_48231_n1109), .B(u3_u0__abc_48231_n1106), .Y(u3_u0__abc_48231_n1110) );
  OR2X2 OR2X2_4524 ( .A(u3_u0__abc_48231_n1110), .B(u3_u0__abc_48231_n1105), .Y(u3_rd_fifo_out_8_) );
  OR2X2 OR2X2_4525 ( .A(u3_u0__abc_48231_n1114), .B(u3_u0__abc_48231_n1115), .Y(u3_u0__abc_48231_n1116) );
  OR2X2 OR2X2_4526 ( .A(u3_u0__abc_48231_n1116), .B(u3_u0__abc_48231_n1113), .Y(u3_u0__abc_48231_n1117) );
  OR2X2 OR2X2_4527 ( .A(u3_u0__abc_48231_n1117), .B(u3_u0__abc_48231_n1112), .Y(u3_rd_fifo_out_9_) );
  OR2X2 OR2X2_4528 ( .A(u3_u0__abc_48231_n1121), .B(u3_u0__abc_48231_n1122), .Y(u3_u0__abc_48231_n1123) );
  OR2X2 OR2X2_4529 ( .A(u3_u0__abc_48231_n1123), .B(u3_u0__abc_48231_n1120), .Y(u3_u0__abc_48231_n1124) );
  OR2X2 OR2X2_453 ( .A(u0__abc_49347_n2084), .B(u0__abc_49347_n2085), .Y(u0__abc_49347_n2086) );
  OR2X2 OR2X2_4530 ( .A(u3_u0__abc_48231_n1124), .B(u3_u0__abc_48231_n1119), .Y(u3_rd_fifo_out_10_) );
  OR2X2 OR2X2_4531 ( .A(u3_u0__abc_48231_n1128), .B(u3_u0__abc_48231_n1129), .Y(u3_u0__abc_48231_n1130) );
  OR2X2 OR2X2_4532 ( .A(u3_u0__abc_48231_n1130), .B(u3_u0__abc_48231_n1127), .Y(u3_u0__abc_48231_n1131) );
  OR2X2 OR2X2_4533 ( .A(u3_u0__abc_48231_n1131), .B(u3_u0__abc_48231_n1126), .Y(u3_rd_fifo_out_11_) );
  OR2X2 OR2X2_4534 ( .A(u3_u0__abc_48231_n1135), .B(u3_u0__abc_48231_n1136), .Y(u3_u0__abc_48231_n1137) );
  OR2X2 OR2X2_4535 ( .A(u3_u0__abc_48231_n1137), .B(u3_u0__abc_48231_n1134), .Y(u3_u0__abc_48231_n1138) );
  OR2X2 OR2X2_4536 ( .A(u3_u0__abc_48231_n1138), .B(u3_u0__abc_48231_n1133), .Y(u3_rd_fifo_out_12_) );
  OR2X2 OR2X2_4537 ( .A(u3_u0__abc_48231_n1142), .B(u3_u0__abc_48231_n1143), .Y(u3_u0__abc_48231_n1144) );
  OR2X2 OR2X2_4538 ( .A(u3_u0__abc_48231_n1144), .B(u3_u0__abc_48231_n1141), .Y(u3_u0__abc_48231_n1145) );
  OR2X2 OR2X2_4539 ( .A(u3_u0__abc_48231_n1145), .B(u3_u0__abc_48231_n1140), .Y(u3_rd_fifo_out_13_) );
  OR2X2 OR2X2_454 ( .A(u0__abc_49347_n2087), .B(u0__abc_49347_n2088), .Y(u0__abc_49347_n2089) );
  OR2X2 OR2X2_4540 ( .A(u3_u0__abc_48231_n1149), .B(u3_u0__abc_48231_n1150), .Y(u3_u0__abc_48231_n1151) );
  OR2X2 OR2X2_4541 ( .A(u3_u0__abc_48231_n1151), .B(u3_u0__abc_48231_n1148), .Y(u3_u0__abc_48231_n1152) );
  OR2X2 OR2X2_4542 ( .A(u3_u0__abc_48231_n1152), .B(u3_u0__abc_48231_n1147), .Y(u3_rd_fifo_out_14_) );
  OR2X2 OR2X2_4543 ( .A(u3_u0__abc_48231_n1156), .B(u3_u0__abc_48231_n1157), .Y(u3_u0__abc_48231_n1158) );
  OR2X2 OR2X2_4544 ( .A(u3_u0__abc_48231_n1158), .B(u3_u0__abc_48231_n1155), .Y(u3_u0__abc_48231_n1159) );
  OR2X2 OR2X2_4545 ( .A(u3_u0__abc_48231_n1159), .B(u3_u0__abc_48231_n1154), .Y(u3_rd_fifo_out_15_) );
  OR2X2 OR2X2_4546 ( .A(u3_u0__abc_48231_n1163), .B(u3_u0__abc_48231_n1164), .Y(u3_u0__abc_48231_n1165) );
  OR2X2 OR2X2_4547 ( .A(u3_u0__abc_48231_n1165), .B(u3_u0__abc_48231_n1162), .Y(u3_u0__abc_48231_n1166) );
  OR2X2 OR2X2_4548 ( .A(u3_u0__abc_48231_n1166), .B(u3_u0__abc_48231_n1161), .Y(u3_rd_fifo_out_16_) );
  OR2X2 OR2X2_4549 ( .A(u3_u0__abc_48231_n1170), .B(u3_u0__abc_48231_n1171), .Y(u3_u0__abc_48231_n1172) );
  OR2X2 OR2X2_455 ( .A(u0__abc_49347_n2091), .B(spec_req_cs_0_bF_buf0), .Y(u0__abc_49347_n2092) );
  OR2X2 OR2X2_4550 ( .A(u3_u0__abc_48231_n1172), .B(u3_u0__abc_48231_n1169), .Y(u3_u0__abc_48231_n1173) );
  OR2X2 OR2X2_4551 ( .A(u3_u0__abc_48231_n1173), .B(u3_u0__abc_48231_n1168), .Y(u3_rd_fifo_out_17_) );
  OR2X2 OR2X2_4552 ( .A(u3_u0__abc_48231_n1177), .B(u3_u0__abc_48231_n1178), .Y(u3_u0__abc_48231_n1179) );
  OR2X2 OR2X2_4553 ( .A(u3_u0__abc_48231_n1179), .B(u3_u0__abc_48231_n1176), .Y(u3_u0__abc_48231_n1180) );
  OR2X2 OR2X2_4554 ( .A(u3_u0__abc_48231_n1180), .B(u3_u0__abc_48231_n1175), .Y(u3_rd_fifo_out_18_) );
  OR2X2 OR2X2_4555 ( .A(u3_u0__abc_48231_n1184), .B(u3_u0__abc_48231_n1185), .Y(u3_u0__abc_48231_n1186) );
  OR2X2 OR2X2_4556 ( .A(u3_u0__abc_48231_n1186), .B(u3_u0__abc_48231_n1183), .Y(u3_u0__abc_48231_n1187) );
  OR2X2 OR2X2_4557 ( .A(u3_u0__abc_48231_n1187), .B(u3_u0__abc_48231_n1182), .Y(u3_rd_fifo_out_19_) );
  OR2X2 OR2X2_4558 ( .A(u3_u0__abc_48231_n1191), .B(u3_u0__abc_48231_n1192), .Y(u3_u0__abc_48231_n1193) );
  OR2X2 OR2X2_4559 ( .A(u3_u0__abc_48231_n1193), .B(u3_u0__abc_48231_n1190), .Y(u3_u0__abc_48231_n1194) );
  OR2X2 OR2X2_456 ( .A(u0__abc_49347_n2090), .B(u0__abc_49347_n2092), .Y(u0__abc_49347_n2093) );
  OR2X2 OR2X2_4560 ( .A(u3_u0__abc_48231_n1194), .B(u3_u0__abc_48231_n1189), .Y(u3_rd_fifo_out_20_) );
  OR2X2 OR2X2_4561 ( .A(u3_u0__abc_48231_n1198), .B(u3_u0__abc_48231_n1199), .Y(u3_u0__abc_48231_n1200) );
  OR2X2 OR2X2_4562 ( .A(u3_u0__abc_48231_n1200), .B(u3_u0__abc_48231_n1197), .Y(u3_u0__abc_48231_n1201) );
  OR2X2 OR2X2_4563 ( .A(u3_u0__abc_48231_n1201), .B(u3_u0__abc_48231_n1196), .Y(u3_rd_fifo_out_21_) );
  OR2X2 OR2X2_4564 ( .A(u3_u0__abc_48231_n1205), .B(u3_u0__abc_48231_n1206), .Y(u3_u0__abc_48231_n1207) );
  OR2X2 OR2X2_4565 ( .A(u3_u0__abc_48231_n1207), .B(u3_u0__abc_48231_n1204), .Y(u3_u0__abc_48231_n1208) );
  OR2X2 OR2X2_4566 ( .A(u3_u0__abc_48231_n1208), .B(u3_u0__abc_48231_n1203), .Y(u3_rd_fifo_out_22_) );
  OR2X2 OR2X2_4567 ( .A(u3_u0__abc_48231_n1212), .B(u3_u0__abc_48231_n1213), .Y(u3_u0__abc_48231_n1214) );
  OR2X2 OR2X2_4568 ( .A(u3_u0__abc_48231_n1214), .B(u3_u0__abc_48231_n1211), .Y(u3_u0__abc_48231_n1215) );
  OR2X2 OR2X2_4569 ( .A(u3_u0__abc_48231_n1215), .B(u3_u0__abc_48231_n1210), .Y(u3_rd_fifo_out_23_) );
  OR2X2 OR2X2_457 ( .A(u0__abc_49347_n1203_bF_buf3), .B(u0_csc0_5_), .Y(u0__abc_49347_n2094) );
  OR2X2 OR2X2_4570 ( .A(u3_u0__abc_48231_n1219), .B(u3_u0__abc_48231_n1220), .Y(u3_u0__abc_48231_n1221) );
  OR2X2 OR2X2_4571 ( .A(u3_u0__abc_48231_n1221), .B(u3_u0__abc_48231_n1218), .Y(u3_u0__abc_48231_n1222) );
  OR2X2 OR2X2_4572 ( .A(u3_u0__abc_48231_n1222), .B(u3_u0__abc_48231_n1217), .Y(u3_rd_fifo_out_24_) );
  OR2X2 OR2X2_4573 ( .A(u3_u0__abc_48231_n1226), .B(u3_u0__abc_48231_n1227), .Y(u3_u0__abc_48231_n1228) );
  OR2X2 OR2X2_4574 ( .A(u3_u0__abc_48231_n1228), .B(u3_u0__abc_48231_n1225), .Y(u3_u0__abc_48231_n1229) );
  OR2X2 OR2X2_4575 ( .A(u3_u0__abc_48231_n1229), .B(u3_u0__abc_48231_n1224), .Y(u3_rd_fifo_out_25_) );
  OR2X2 OR2X2_4576 ( .A(u3_u0__abc_48231_n1233), .B(u3_u0__abc_48231_n1234), .Y(u3_u0__abc_48231_n1235) );
  OR2X2 OR2X2_4577 ( .A(u3_u0__abc_48231_n1235), .B(u3_u0__abc_48231_n1232), .Y(u3_u0__abc_48231_n1236) );
  OR2X2 OR2X2_4578 ( .A(u3_u0__abc_48231_n1236), .B(u3_u0__abc_48231_n1231), .Y(u3_rd_fifo_out_26_) );
  OR2X2 OR2X2_4579 ( .A(u3_u0__abc_48231_n1240), .B(u3_u0__abc_48231_n1241), .Y(u3_u0__abc_48231_n1242) );
  OR2X2 OR2X2_458 ( .A(u0__abc_49347_n2096), .B(u0__abc_49347_n2074), .Y(u0_sp_csc_5__FF_INPUT) );
  OR2X2 OR2X2_4580 ( .A(u3_u0__abc_48231_n1242), .B(u3_u0__abc_48231_n1239), .Y(u3_u0__abc_48231_n1243) );
  OR2X2 OR2X2_4581 ( .A(u3_u0__abc_48231_n1243), .B(u3_u0__abc_48231_n1238), .Y(u3_rd_fifo_out_27_) );
  OR2X2 OR2X2_4582 ( .A(u3_u0__abc_48231_n1247), .B(u3_u0__abc_48231_n1248), .Y(u3_u0__abc_48231_n1249) );
  OR2X2 OR2X2_4583 ( .A(u3_u0__abc_48231_n1249), .B(u3_u0__abc_48231_n1246), .Y(u3_u0__abc_48231_n1250) );
  OR2X2 OR2X2_4584 ( .A(u3_u0__abc_48231_n1250), .B(u3_u0__abc_48231_n1245), .Y(u3_rd_fifo_out_28_) );
  OR2X2 OR2X2_4585 ( .A(u3_u0__abc_48231_n1254), .B(u3_u0__abc_48231_n1255), .Y(u3_u0__abc_48231_n1256) );
  OR2X2 OR2X2_4586 ( .A(u3_u0__abc_48231_n1256), .B(u3_u0__abc_48231_n1253), .Y(u3_u0__abc_48231_n1257) );
  OR2X2 OR2X2_4587 ( .A(u3_u0__abc_48231_n1257), .B(u3_u0__abc_48231_n1252), .Y(u3_rd_fifo_out_29_) );
  OR2X2 OR2X2_4588 ( .A(u3_u0__abc_48231_n1261), .B(u3_u0__abc_48231_n1262), .Y(u3_u0__abc_48231_n1263) );
  OR2X2 OR2X2_4589 ( .A(u3_u0__abc_48231_n1263), .B(u3_u0__abc_48231_n1260), .Y(u3_u0__abc_48231_n1264) );
  OR2X2 OR2X2_459 ( .A(u0__abc_49347_n1183_1_bF_buf2), .B(1'b0), .Y(u0__abc_49347_n2100) );
  OR2X2 OR2X2_4590 ( .A(u3_u0__abc_48231_n1264), .B(u3_u0__abc_48231_n1259), .Y(u3_rd_fifo_out_30_) );
  OR2X2 OR2X2_4591 ( .A(u3_u0__abc_48231_n1268), .B(u3_u0__abc_48231_n1269), .Y(u3_u0__abc_48231_n1270) );
  OR2X2 OR2X2_4592 ( .A(u3_u0__abc_48231_n1270), .B(u3_u0__abc_48231_n1267), .Y(u3_u0__abc_48231_n1271) );
  OR2X2 OR2X2_4593 ( .A(u3_u0__abc_48231_n1271), .B(u3_u0__abc_48231_n1266), .Y(u3_rd_fifo_out_31_) );
  OR2X2 OR2X2_4594 ( .A(u3_u0__abc_48231_n1275), .B(u3_u0__abc_48231_n1276), .Y(u3_u0__abc_48231_n1277) );
  OR2X2 OR2X2_4595 ( .A(u3_u0__abc_48231_n1277), .B(u3_u0__abc_48231_n1274), .Y(u3_u0__abc_48231_n1278) );
  OR2X2 OR2X2_4596 ( .A(u3_u0__abc_48231_n1278), .B(u3_u0__abc_48231_n1273), .Y(u3_rd_fifo_out_32_) );
  OR2X2 OR2X2_4597 ( .A(u3_u0__abc_48231_n1282), .B(u3_u0__abc_48231_n1283), .Y(u3_u0__abc_48231_n1284) );
  OR2X2 OR2X2_4598 ( .A(u3_u0__abc_48231_n1284), .B(u3_u0__abc_48231_n1281), .Y(u3_u0__abc_48231_n1285) );
  OR2X2 OR2X2_4599 ( .A(u3_u0__abc_48231_n1285), .B(u3_u0__abc_48231_n1280), .Y(u3_rd_fifo_out_33_) );
  OR2X2 OR2X2_46 ( .A(lmr_sel_bF_buf0), .B(tms_5_), .Y(_abc_55805_n306) );
  OR2X2 OR2X2_460 ( .A(spec_req_cs_6_bF_buf5), .B(1'b0), .Y(u0__abc_49347_n2101) );
  OR2X2 OR2X2_4600 ( .A(u3_u0__abc_48231_n1289), .B(u3_u0__abc_48231_n1290), .Y(u3_u0__abc_48231_n1291) );
  OR2X2 OR2X2_4601 ( .A(u3_u0__abc_48231_n1291), .B(u3_u0__abc_48231_n1288), .Y(u3_u0__abc_48231_n1292) );
  OR2X2 OR2X2_4602 ( .A(u3_u0__abc_48231_n1292), .B(u3_u0__abc_48231_n1287), .Y(u3_rd_fifo_out_34_) );
  OR2X2 OR2X2_4603 ( .A(u3_u0__abc_48231_n1296), .B(u3_u0__abc_48231_n1297), .Y(u3_u0__abc_48231_n1298) );
  OR2X2 OR2X2_4604 ( .A(u3_u0__abc_48231_n1298), .B(u3_u0__abc_48231_n1295), .Y(u3_u0__abc_48231_n1299) );
  OR2X2 OR2X2_4605 ( .A(u3_u0__abc_48231_n1299), .B(u3_u0__abc_48231_n1294), .Y(u3_rd_fifo_out_35_) );
  OR2X2 OR2X2_4606 ( .A(cs_need_rfr_6_), .B(cs_need_rfr_7_), .Y(u4__abc_49152_n65) );
  OR2X2 OR2X2_4607 ( .A(cs_need_rfr_4_), .B(cs_need_rfr_5_), .Y(u4__abc_49152_n66_1) );
  OR2X2 OR2X2_4608 ( .A(u4__abc_49152_n65), .B(u4__abc_49152_n66_1), .Y(u4__abc_49152_n67) );
  OR2X2 OR2X2_4609 ( .A(cs_need_rfr_2_), .B(cs_need_rfr_3_), .Y(u4__abc_49152_n68) );
  OR2X2 OR2X2_461 ( .A(u0__abc_49347_n2103), .B(u0__abc_49347_n2099), .Y(u0__abc_49347_n2104) );
  OR2X2 OR2X2_4610 ( .A(cs_need_rfr_0_), .B(cs_need_rfr_1_), .Y(u4__abc_49152_n69_1) );
  OR2X2 OR2X2_4611 ( .A(u4__abc_49152_n68), .B(u4__abc_49152_n69_1), .Y(u4__abc_49152_n70) );
  OR2X2 OR2X2_4612 ( .A(u4__abc_49152_n67), .B(u4__abc_49152_n70), .Y(u4_rfr_en_FF_INPUT) );
  OR2X2 OR2X2_4613 ( .A(u4__abc_49152_n73_1), .B(u4__abc_49152_n75), .Y(u4__abc_49152_n76_1) );
  OR2X2 OR2X2_4614 ( .A(u4__abc_49152_n78), .B(u4__abc_49152_n80), .Y(u4__abc_49152_n81) );
  OR2X2 OR2X2_4615 ( .A(u4__abc_49152_n76_1), .B(u4__abc_49152_n81), .Y(u4__abc_49152_n82_1) );
  OR2X2 OR2X2_4616 ( .A(u4__abc_49152_n84), .B(u4__abc_49152_n86), .Y(u4__abc_49152_n87) );
  OR2X2 OR2X2_4617 ( .A(u4__abc_49152_n89), .B(u4__abc_49152_n91), .Y(u4__abc_49152_n92) );
  OR2X2 OR2X2_4618 ( .A(u4__abc_49152_n87), .B(u4__abc_49152_n92), .Y(u4__abc_49152_n93_1) );
  OR2X2 OR2X2_4619 ( .A(u4__abc_49152_n82_1), .B(u4__abc_49152_n93_1), .Y(u4__abc_49152_n94) );
  OR2X2 OR2X2_462 ( .A(u0__abc_49347_n2105), .B(u0__abc_49347_n2106), .Y(u0__abc_49347_n2107) );
  OR2X2 OR2X2_4620 ( .A(u4__abc_49152_n96), .B(u4__abc_49152_n98), .Y(u4__abc_49152_n99) );
  OR2X2 OR2X2_4621 ( .A(u4__abc_49152_n101_1), .B(u4__abc_49152_n103), .Y(u4__abc_49152_n104_1) );
  OR2X2 OR2X2_4622 ( .A(u4__abc_49152_n99), .B(u4__abc_49152_n104_1), .Y(u4__abc_49152_n105) );
  OR2X2 OR2X2_4623 ( .A(u4__abc_49152_n107), .B(u4__abc_49152_n109), .Y(u4__abc_49152_n110) );
  OR2X2 OR2X2_4624 ( .A(u4_ps_cnt_3_), .B(rfr_ps_val_3_), .Y(u4__abc_49152_n111) );
  OR2X2 OR2X2_4625 ( .A(u4__abc_49152_n110), .B(u4__abc_49152_n114), .Y(u4__abc_49152_n115) );
  OR2X2 OR2X2_4626 ( .A(u4__abc_49152_n105), .B(u4__abc_49152_n115), .Y(u4__abc_49152_n116) );
  OR2X2 OR2X2_4627 ( .A(u4__abc_49152_n94), .B(u4__abc_49152_n116), .Y(u4__abc_49152_n117) );
  OR2X2 OR2X2_4628 ( .A(u4_rfr_clr), .B(rfr_req), .Y(u4__abc_49152_n120) );
  OR2X2 OR2X2_4629 ( .A(u4_rfr_ce), .B(u4_rfr_cnt_0_), .Y(u4__abc_49152_n124_1) );
  OR2X2 OR2X2_463 ( .A(u0__abc_49347_n2108_1), .B(u0__abc_49347_n2109), .Y(u0__abc_49347_n2110) );
  OR2X2 OR2X2_4630 ( .A(u4__abc_49152_n122), .B(u4_rfr_cnt_1_), .Y(u4__abc_49152_n130) );
  OR2X2 OR2X2_4631 ( .A(u4__abc_49152_n128), .B(u4_rfr_cnt_2_), .Y(u4__abc_49152_n133) );
  OR2X2 OR2X2_4632 ( .A(u4__abc_49152_n135), .B(u4_rfr_cnt_3_), .Y(u4__abc_49152_n142) );
  OR2X2 OR2X2_4633 ( .A(u4__abc_49152_n140), .B(u4_rfr_cnt_4_), .Y(u4__abc_49152_n147) );
  OR2X2 OR2X2_4634 ( .A(u4__abc_49152_n145), .B(u4_rfr_cnt_5_), .Y(u4__abc_49152_n150) );
  OR2X2 OR2X2_4635 ( .A(u4__abc_49152_n152), .B(u4_rfr_cnt_6_), .Y(u4__abc_49152_n158) );
  OR2X2 OR2X2_4636 ( .A(u4__abc_49152_n156), .B(u4_rfr_cnt_7_), .Y(u4__abc_49152_n161) );
  OR2X2 OR2X2_4637 ( .A(u4__abc_49152_n117), .B(u4__abc_49152_n174), .Y(u4__abc_49152_n175) );
  OR2X2 OR2X2_4638 ( .A(u4_ps_cnt_0_), .B(u4_rfr_en), .Y(u4__abc_49152_n177) );
  OR2X2 OR2X2_4639 ( .A(u4__abc_49152_n178), .B(u4_ps_cnt_1_), .Y(u4__abc_49152_n182) );
  OR2X2 OR2X2_464 ( .A(u0__abc_49347_n2111), .B(u0__abc_49347_n2112), .Y(u0__abc_49347_n2113) );
  OR2X2 OR2X2_4640 ( .A(u4__abc_49152_n187), .B(u4__abc_49152_n188), .Y(u4__abc_49152_n189_1) );
  OR2X2 OR2X2_4641 ( .A(u4__abc_49152_n192), .B(u4_ps_cnt_3_), .Y(u4__abc_49152_n193) );
  OR2X2 OR2X2_4642 ( .A(u4__abc_49152_n194), .B(u4_ps_cnt_4_), .Y(u4__abc_49152_n198) );
  OR2X2 OR2X2_4643 ( .A(u4__abc_49152_n200), .B(u4_ps_cnt_5_), .Y(u4__abc_49152_n204) );
  OR2X2 OR2X2_4644 ( .A(u4__abc_49152_n205), .B(u4_ps_cnt_6_), .Y(u4__abc_49152_n209) );
  OR2X2 OR2X2_4645 ( .A(u4__abc_49152_n215), .B(u4_ps_cnt_7_), .Y(u4__abc_49152_n221) );
  OR2X2 OR2X2_4646 ( .A(u4__abc_49152_n227), .B(u4__abc_49152_n232), .Y(u4__abc_49152_n233) );
  OR2X2 OR2X2_4647 ( .A(u4__abc_49152_n236), .B(u4__abc_49152_n238), .Y(u4__abc_49152_n239) );
  OR2X2 OR2X2_4648 ( .A(u4__abc_49152_n239), .B(ref_int_2_), .Y(u4__abc_49152_n240) );
  OR2X2 OR2X2_4649 ( .A(u4__abc_49152_n240), .B(u4__abc_49152_n233), .Y(u4__abc_49152_n241) );
  OR2X2 OR2X2_465 ( .A(u0__abc_49347_n2115), .B(spec_req_cs_0_bF_buf5), .Y(u0__abc_49347_n2116) );
  OR2X2 OR2X2_4650 ( .A(u4__abc_49152_n162), .B(u4__abc_49152_n234), .Y(u4__abc_49152_n242) );
  OR2X2 OR2X2_4651 ( .A(u4__abc_49152_n249), .B(u4__abc_49152_n246), .Y(u4__abc_49152_n250) );
  OR2X2 OR2X2_4652 ( .A(u4__abc_49152_n250), .B(u4__abc_49152_n245), .Y(u4__abc_49152_n251) );
  OR2X2 OR2X2_4653 ( .A(u4__abc_49152_n252), .B(u4__abc_49152_n256), .Y(u4_rfr_clr_FF_INPUT) );
  OR2X2 OR2X2_4654 ( .A(u5_burst_cnt_1_), .B(u5_burst_cnt_2_), .Y(u5__abc_54027_n250) );
  OR2X2 OR2X2_4655 ( .A(u5__abc_54027_n250), .B(u5_burst_cnt_0_), .Y(u5__abc_54027_n251) );
  OR2X2 OR2X2_4656 ( .A(u5__abc_54027_n251), .B(u5_burst_cnt_3_), .Y(u5__abc_54027_n252_1) );
  OR2X2 OR2X2_4657 ( .A(u5__abc_54027_n309), .B(u5__abc_54027_n291), .Y(init_ack) );
  OR2X2 OR2X2_4658 ( .A(u5__abc_54027_n322_1), .B(u5__abc_54027_n318), .Y(dv) );
  OR2X2 OR2X2_4659 ( .A(u5_timer_3_), .B(u5_timer_2_), .Y(u5__abc_54027_n325) );
  OR2X2 OR2X2_466 ( .A(u0__abc_49347_n2114), .B(u0__abc_49347_n2116), .Y(u0__abc_49347_n2117) );
  OR2X2 OR2X2_4660 ( .A(u5_timer_1_), .B(u5_timer_0_), .Y(u5__abc_54027_n331) );
  OR2X2 OR2X2_4661 ( .A(u5_timer_7_), .B(u5_timer_6_), .Y(u5__abc_54027_n332) );
  OR2X2 OR2X2_4662 ( .A(u5__abc_54027_n331), .B(u5__abc_54027_n332), .Y(u5__abc_54027_n333_1) );
  OR2X2 OR2X2_4663 ( .A(u5__abc_54027_n345), .B(u5__abc_54027_n348), .Y(u5__abc_54027_n349) );
  OR2X2 OR2X2_4664 ( .A(u5__abc_54027_n354), .B(u5__abc_54027_n355), .Y(u5__abc_54027_n356) );
  OR2X2 OR2X2_4665 ( .A(u5__abc_54027_n356), .B(u5__abc_54027_n352), .Y(u5__abc_54027_n357) );
  OR2X2 OR2X2_4666 ( .A(u5__abc_54027_n357), .B(u5__abc_54027_n349), .Y(u5_rfr_ack_d) );
  OR2X2 OR2X2_4667 ( .A(u5__abc_54027_n395), .B(u5__abc_54027_n394_1), .Y(u5__abc_54027_n396) );
  OR2X2 OR2X2_4668 ( .A(u5__abc_54027_n399), .B(u5__abc_54027_n394_1), .Y(u5__abc_54027_n400) );
  OR2X2 OR2X2_4669 ( .A(u5_state_2_), .B(u5_state_3_), .Y(u5__abc_54027_n409) );
  OR2X2 OR2X2_467 ( .A(u0__abc_49347_n1203_bF_buf2), .B(u0_csc0_6_), .Y(u0__abc_49347_n2118) );
  OR2X2 OR2X2_4670 ( .A(u5__abc_54027_n286), .B(u5_state_1_), .Y(u5__abc_54027_n410) );
  OR2X2 OR2X2_4671 ( .A(u5__abc_54027_n410), .B(u5__abc_54027_n409), .Y(u5__abc_54027_n411) );
  OR2X2 OR2X2_4672 ( .A(u5_state_5_), .B(u5_state_4_), .Y(u5__abc_54027_n412) );
  OR2X2 OR2X2_4673 ( .A(u5__abc_54027_n412), .B(u5__abc_54027_n267), .Y(u5__abc_54027_n413) );
  OR2X2 OR2X2_4674 ( .A(u5__abc_54027_n411), .B(u5__abc_54027_n413), .Y(u5__abc_54027_n414) );
  OR2X2 OR2X2_4675 ( .A(u5__abc_54027_n304), .B(u5__abc_54027_n460), .Y(u5__abc_54027_n461_1) );
  OR2X2 OR2X2_4676 ( .A(u5__abc_54027_n472), .B(tms_s_9_), .Y(u5__abc_54027_n473) );
  OR2X2 OR2X2_4677 ( .A(u5__abc_54027_n478_1), .B(u5__abc_54027_n479), .Y(u5__abc_54027_n480) );
  OR2X2 OR2X2_4678 ( .A(u5__abc_54027_n473), .B(u5__abc_54027_n480), .Y(u5__abc_54027_n481) );
  OR2X2 OR2X2_4679 ( .A(u5__abc_54027_n474), .B(u5_cke_r), .Y(u5__abc_54027_n482) );
  OR2X2 OR2X2_468 ( .A(u0__abc_49347_n2120), .B(u0__abc_49347_n2098), .Y(u0_sp_csc_6__FF_INPUT) );
  OR2X2 OR2X2_4680 ( .A(u5__abc_54027_n485), .B(u5__abc_54027_n421), .Y(u5__abc_54027_n486_1) );
  OR2X2 OR2X2_4681 ( .A(u5__abc_54027_n484_1), .B(u5__abc_54027_n486_1), .Y(u5__abc_54027_n487) );
  OR2X2 OR2X2_4682 ( .A(obct_cs_6_), .B(obct_cs_7_), .Y(u5__abc_54027_n493_1) );
  OR2X2 OR2X2_4683 ( .A(obct_cs_4_), .B(obct_cs_5_), .Y(u5__abc_54027_n494) );
  OR2X2 OR2X2_4684 ( .A(u5__abc_54027_n493_1), .B(u5__abc_54027_n494), .Y(u5__abc_54027_n495_1) );
  OR2X2 OR2X2_4685 ( .A(obct_cs_2_), .B(obct_cs_3_), .Y(u5__abc_54027_n496) );
  OR2X2 OR2X2_4686 ( .A(obct_cs_0_), .B(obct_cs_1_), .Y(u5__abc_54027_n497) );
  OR2X2 OR2X2_4687 ( .A(u5__abc_54027_n496), .B(u5__abc_54027_n497), .Y(u5__abc_54027_n498) );
  OR2X2 OR2X2_4688 ( .A(u5__abc_54027_n495_1), .B(u5__abc_54027_n498), .Y(u5__abc_54027_n499) );
  OR2X2 OR2X2_4689 ( .A(u5__abc_54027_n517), .B(u5__abc_54027_n414), .Y(u5__abc_54027_n518) );
  OR2X2 OR2X2_469 ( .A(u0__abc_49347_n1183_1_bF_buf1), .B(1'b0), .Y(u0__abc_49347_n2124) );
  OR2X2 OR2X2_4690 ( .A(u5__abc_54027_n453), .B(u5__abc_54027_n520), .Y(u5__abc_54027_n521) );
  OR2X2 OR2X2_4691 ( .A(u5__abc_54027_n530), .B(u5__abc_54027_n466), .Y(u5_cmd_0_) );
  OR2X2 OR2X2_4692 ( .A(u5__abc_54027_n534), .B(u5__abc_54027_n532_1), .Y(u5_we_) );
  OR2X2 OR2X2_4693 ( .A(u5__abc_54027_n539), .B(u5__abc_54027_n466), .Y(u5_cmd_1_) );
  OR2X2 OR2X2_4694 ( .A(u5__abc_54027_n542), .B(u5__abc_54027_n541), .Y(cas_) );
  OR2X2 OR2X2_4695 ( .A(u5__abc_54027_n363), .B(u5__abc_54027_n545_1), .Y(u5__abc_54027_n546) );
  OR2X2 OR2X2_4696 ( .A(u5__abc_54027_n466), .B(u5__abc_54027_n551), .Y(u5_cmd_2_) );
  OR2X2 OR2X2_4697 ( .A(u5__abc_54027_n554), .B(u5__abc_54027_n553_1), .Y(ras_) );
  OR2X2 OR2X2_4698 ( .A(u5__abc_54027_n558), .B(u5__abc_54027_n421), .Y(u5__abc_54027_n559) );
  OR2X2 OR2X2_4699 ( .A(u5_rfr_ack_d), .B(u5__abc_54027_n564), .Y(u5__abc_54027_n565) );
  OR2X2 OR2X2_47 ( .A(_abc_55805_n240_bF_buf3), .B(sp_tms_6_), .Y(_abc_55805_n308) );
  OR2X2 OR2X2_470 ( .A(spec_req_cs_6_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n2125) );
  OR2X2 OR2X2_4700 ( .A(u5__abc_54027_n565_bF_buf4), .B(tms_s_19_), .Y(u5__abc_54027_n566_1) );
  OR2X2 OR2X2_4701 ( .A(tms_s_16_), .B(tms_s_17_), .Y(u5__abc_54027_n567) );
  OR2X2 OR2X2_4702 ( .A(u5__abc_54027_n567), .B(tms_s_18_), .Y(u5__abc_54027_n568) );
  OR2X2 OR2X2_4703 ( .A(u5__abc_54027_n566_1), .B(u5__abc_54027_n568), .Y(u5__abc_54027_n569_1) );
  OR2X2 OR2X2_4704 ( .A(u5__abc_54027_n417), .B(u5_tmr_done), .Y(u5__abc_54027_n579_1) );
  OR2X2 OR2X2_4705 ( .A(u5__abc_54027_n361), .B(u5_tmr2_done), .Y(u5__abc_54027_n580) );
  OR2X2 OR2X2_4706 ( .A(csc_s_3_), .B(csc_s_2_bF_buf1), .Y(u5__abc_54027_n593) );
  OR2X2 OR2X2_4707 ( .A(u5__abc_54027_n599), .B(u5__abc_54027_n589), .Y(u5__abc_54027_n600) );
  OR2X2 OR2X2_4708 ( .A(u5__abc_54027_n610), .B(u5__abc_54027_n609), .Y(cs_en) );
  OR2X2 OR2X2_4709 ( .A(u5__abc_54027_n614), .B(u5__abc_54027_n616), .Y(u5__abc_54027_n617) );
  OR2X2 OR2X2_471 ( .A(u0__abc_49347_n2127), .B(u0__abc_49347_n2123), .Y(u0__abc_49347_n2128) );
  OR2X2 OR2X2_4710 ( .A(u5__abc_54027_n620_1), .B(u5__abc_54027_n416), .Y(u5__abc_54027_n621) );
  OR2X2 OR2X2_4711 ( .A(u5__abc_54027_n618), .B(u5__abc_54027_n621), .Y(u5__abc_54027_n622) );
  OR2X2 OR2X2_4712 ( .A(u5__abc_54027_n622), .B(u5__abc_54027_n617), .Y(u5__abc_54027_n623) );
  OR2X2 OR2X2_4713 ( .A(u5__abc_54027_n623), .B(u5__abc_54027_n613), .Y(u5__abc_54027_n624) );
  OR2X2 OR2X2_4714 ( .A(u5__abc_54027_n570), .B(u5__abc_54027_n624), .Y(u5_data_oe_d) );
  OR2X2 OR2X2_4715 ( .A(u5__abc_54027_n627), .B(u5__abc_54027_n626), .Y(u5_data_oe_FF_INPUT) );
  OR2X2 OR2X2_4716 ( .A(u5__abc_54027_n632_1), .B(u5__abc_54027_n500), .Y(u5__abc_54027_n633) );
  OR2X2 OR2X2_4717 ( .A(u5__abc_54027_n631), .B(u5__abc_54027_n633), .Y(u5__abc_54027_n634) );
  OR2X2 OR2X2_4718 ( .A(u5__abc_54027_n640), .B(u5_ack_cnt_3_), .Y(u5__abc_54027_n641) );
  OR2X2 OR2X2_4719 ( .A(u5__abc_54027_n642), .B(u5__abc_54027_n634), .Y(u5__abc_54027_n643_1) );
  OR2X2 OR2X2_472 ( .A(u0__abc_49347_n2129), .B(u0__abc_49347_n2130), .Y(u0__abc_49347_n2131) );
  OR2X2 OR2X2_4720 ( .A(u5__abc_54027_n616), .B(u5__abc_54027_n648), .Y(u5__abc_54027_n649) );
  OR2X2 OR2X2_4721 ( .A(u5__abc_54027_n649), .B(u5__abc_54027_n645), .Y(u5__abc_54027_n650) );
  OR2X2 OR2X2_4722 ( .A(u5__abc_54027_n677), .B(u5__abc_54027_n265), .Y(u5__abc_54027_n678) );
  OR2X2 OR2X2_4723 ( .A(u5__abc_54027_n681_1), .B(u5__abc_54027_n682), .Y(u5__abc_54027_n683) );
  OR2X2 OR2X2_4724 ( .A(u5__abc_54027_n678), .B(u5__abc_54027_n685_1), .Y(u5__abc_54027_n686) );
  OR2X2 OR2X2_4725 ( .A(u5__abc_54027_n688), .B(u5_no_wb_cycle_FF_INPUT), .Y(u5__abc_54027_n689) );
  OR2X2 OR2X2_4726 ( .A(u5__abc_54027_n691), .B(u5_wb_stb_first), .Y(u5__abc_54027_n692) );
  OR2X2 OR2X2_4727 ( .A(u5__abc_54027_n696), .B(u5__abc_54027_n694_1), .Y(u5_ap_en_FF_INPUT) );
  OR2X2 OR2X2_4728 ( .A(u5__abc_54027_n687_1), .B(u5__abc_54027_n533), .Y(u5__abc_54027_n699_1) );
  OR2X2 OR2X2_4729 ( .A(u5__abc_54027_n704), .B(u5__abc_54027_n705_1), .Y(u5__abc_54027_n706) );
  OR2X2 OR2X2_473 ( .A(u0__abc_49347_n2132), .B(u0__abc_49347_n2133), .Y(u0__abc_49347_n2134) );
  OR2X2 OR2X2_4730 ( .A(u5__abc_54027_n706), .B(u5__abc_54027_n351_bF_buf0), .Y(u5__abc_54027_n707) );
  OR2X2 OR2X2_4731 ( .A(u5__abc_54027_n710), .B(u5__abc_54027_n677), .Y(u5__abc_54027_n711) );
  OR2X2 OR2X2_4732 ( .A(u5__abc_54027_n711), .B(u5__abc_54027_n414), .Y(u5__abc_54027_n712) );
  OR2X2 OR2X2_4733 ( .A(u5__abc_54027_n718), .B(u5__abc_54027_n351_bF_buf3), .Y(u5__abc_54027_n719) );
  OR2X2 OR2X2_4734 ( .A(u5__abc_54027_n719), .B(u5__abc_54027_n716), .Y(u5__abc_54027_n720) );
  OR2X2 OR2X2_4735 ( .A(u5__abc_54027_n723), .B(u5__abc_54027_n414), .Y(u5__abc_54027_n724) );
  OR2X2 OR2X2_4736 ( .A(u5__abc_54027_n724), .B(u5__abc_54027_n721), .Y(u5__abc_54027_n725) );
  OR2X2 OR2X2_4737 ( .A(u5__abc_54027_n731), .B(u5__abc_54027_n729_1), .Y(u5__abc_54027_n732) );
  OR2X2 OR2X2_4738 ( .A(u5__abc_54027_n735), .B(u5__abc_54027_n736), .Y(u5__abc_54027_n737_1) );
  OR2X2 OR2X2_4739 ( .A(u5__abc_54027_n738), .B(u5__abc_54027_n369), .Y(u5__abc_54027_n739) );
  OR2X2 OR2X2_474 ( .A(u0__abc_49347_n2135), .B(u0__abc_49347_n2136), .Y(u0__abc_49347_n2137) );
  OR2X2 OR2X2_4740 ( .A(u5__abc_54027_n733), .B(u5__abc_54027_n739), .Y(u5_burst_cnt_2__FF_INPUT) );
  OR2X2 OR2X2_4741 ( .A(u5__abc_54027_n715), .B(u5__abc_54027_n250), .Y(u5__abc_54027_n741) );
  OR2X2 OR2X2_4742 ( .A(u5__abc_54027_n743), .B(u5__abc_54027_n351_bF_buf1), .Y(u5__abc_54027_n744_1) );
  OR2X2 OR2X2_4743 ( .A(u5__abc_54027_n742), .B(u5__abc_54027_n744_1), .Y(u5__abc_54027_n745) );
  OR2X2 OR2X2_4744 ( .A(u5__abc_54027_n746), .B(u5__abc_54027_n747_1), .Y(u5__abc_54027_n748) );
  OR2X2 OR2X2_4745 ( .A(u5__abc_54027_n748), .B(u5__abc_54027_n414), .Y(u5__abc_54027_n749) );
  OR2X2 OR2X2_4746 ( .A(u5__abc_54027_n702), .B(u5__abc_54027_n252_1), .Y(u5__abc_54027_n752_1) );
  OR2X2 OR2X2_4747 ( .A(u5__abc_54027_n753), .B(u5__abc_54027_n754), .Y(u5__abc_54027_n755_1) );
  OR2X2 OR2X2_4748 ( .A(u5__abc_54027_n756), .B(u5__abc_54027_n758), .Y(u5__abc_54027_n759_1) );
  OR2X2 OR2X2_4749 ( .A(u5__abc_54027_n763_1), .B(u5__abc_54027_n351_bF_buf3), .Y(u5__abc_54027_n764) );
  OR2X2 OR2X2_475 ( .A(u0__abc_49347_n2139), .B(spec_req_cs_0_bF_buf4), .Y(u0__abc_49347_n2140) );
  OR2X2 OR2X2_4750 ( .A(u5__abc_54027_n762_1), .B(u5__abc_54027_n764), .Y(u5__abc_54027_n765) );
  OR2X2 OR2X2_4751 ( .A(u5__abc_54027_n766_1), .B(u5__abc_54027_n414), .Y(u5__abc_54027_n767_1) );
  OR2X2 OR2X2_4752 ( .A(u5__abc_54027_n771_1), .B(u5__abc_54027_n772_1), .Y(u5__abc_54027_n773) );
  OR2X2 OR2X2_4753 ( .A(u5__abc_54027_n774), .B(u5__abc_54027_n776), .Y(u5__abc_54027_n777) );
  OR2X2 OR2X2_4754 ( .A(u5__abc_54027_n781), .B(u5__abc_54027_n351_bF_buf1), .Y(u5__abc_54027_n782) );
  OR2X2 OR2X2_4755 ( .A(u5__abc_54027_n782), .B(u5__abc_54027_n780), .Y(u5__abc_54027_n783) );
  OR2X2 OR2X2_4756 ( .A(u5__abc_54027_n784), .B(u5__abc_54027_n414), .Y(u5__abc_54027_n785) );
  OR2X2 OR2X2_4757 ( .A(u5__abc_54027_n702), .B(u5__abc_54027_n790), .Y(u5__abc_54027_n791_1) );
  OR2X2 OR2X2_4758 ( .A(u5__abc_54027_n792), .B(u5__abc_54027_n351_bF_buf0), .Y(u5__abc_54027_n793) );
  OR2X2 OR2X2_4759 ( .A(u5__abc_54027_n788), .B(u5__abc_54027_n793), .Y(u5__abc_54027_n794) );
  OR2X2 OR2X2_476 ( .A(u0__abc_49347_n2138), .B(u0__abc_49347_n2140), .Y(u0__abc_49347_n2141) );
  OR2X2 OR2X2_4760 ( .A(u5__abc_54027_n795), .B(u5__abc_54027_n414), .Y(u5__abc_54027_n796) );
  OR2X2 OR2X2_4761 ( .A(u5__abc_54027_n799), .B(u5_burst_cnt_9_), .Y(u5__abc_54027_n800) );
  OR2X2 OR2X2_4762 ( .A(u5__abc_54027_n801_1), .B(u5__abc_54027_n257), .Y(u5__abc_54027_n802) );
  OR2X2 OR2X2_4763 ( .A(u5__abc_54027_n702), .B(u5__abc_54027_n803), .Y(u5__abc_54027_n804) );
  OR2X2 OR2X2_4764 ( .A(u5__abc_54027_n703), .B(u5_burst_cnt_9_), .Y(u5__abc_54027_n805) );
  OR2X2 OR2X2_4765 ( .A(u5__abc_54027_n807), .B(u5__abc_54027_n809), .Y(u5__abc_54027_n810_1) );
  OR2X2 OR2X2_4766 ( .A(u5__abc_54027_n812), .B(u5_burst_cnt_10_), .Y(u5__abc_54027_n813) );
  OR2X2 OR2X2_4767 ( .A(u5__abc_54027_n814), .B(u5__abc_54027_n256_1), .Y(u5__abc_54027_n815) );
  OR2X2 OR2X2_4768 ( .A(u5__abc_54027_n702), .B(u5__abc_54027_n816), .Y(u5__abc_54027_n817) );
  OR2X2 OR2X2_4769 ( .A(u5__abc_54027_n703), .B(u5_burst_cnt_10_), .Y(u5__abc_54027_n818) );
  OR2X2 OR2X2_477 ( .A(u0__abc_49347_n1203_bF_buf1), .B(u0_csc0_7_), .Y(u0__abc_49347_n2142) );
  OR2X2 OR2X2_4770 ( .A(u5__abc_54027_n820), .B(u5__abc_54027_n822), .Y(u5__abc_54027_n823) );
  OR2X2 OR2X2_4771 ( .A(u5__abc_54027_n827), .B(u5__abc_54027_n828), .Y(u5__abc_54027_n829) );
  OR2X2 OR2X2_4772 ( .A(u5__abc_54027_n833_1), .B(u5__abc_54027_n291), .Y(u5__abc_54027_n834) );
  OR2X2 OR2X2_4773 ( .A(u5__abc_54027_n834), .B(u5__abc_54027_n832), .Y(u5_ir_cnt_1__FF_INPUT) );
  OR2X2 OR2X2_4774 ( .A(u5__abc_54027_n837), .B(u5__abc_54027_n838), .Y(u5__abc_54027_n839) );
  OR2X2 OR2X2_4775 ( .A(u5__abc_54027_n842), .B(u5__abc_54027_n843_1), .Y(u5__abc_54027_n844) );
  OR2X2 OR2X2_4776 ( .A(u5__abc_54027_n565_bF_buf3), .B(tms_s_0_), .Y(u5__abc_54027_n846) );
  OR2X2 OR2X2_4777 ( .A(u5__abc_54027_n846), .B(u5__abc_54027_n850), .Y(u5__abc_54027_n851) );
  OR2X2 OR2X2_4778 ( .A(u5__abc_54027_n565_bF_buf2), .B(tms_s_4_), .Y(u5__abc_54027_n855_1) );
  OR2X2 OR2X2_4779 ( .A(u5__abc_54027_n461_1), .B(u5__abc_54027_n355), .Y(u5__abc_54027_n857) );
  OR2X2 OR2X2_478 ( .A(u0__abc_49347_n2144_1), .B(u0__abc_49347_n2122), .Y(u0_sp_csc_7__FF_INPUT) );
  OR2X2 OR2X2_4780 ( .A(u5__abc_54027_n857), .B(u5__abc_54027_n301_1), .Y(u5__abc_54027_n858) );
  OR2X2 OR2X2_4781 ( .A(u5__abc_54027_n565_bF_buf1), .B(tms_s_24_), .Y(u5__abc_54027_n860) );
  OR2X2 OR2X2_4782 ( .A(u5__abc_54027_n860), .B(u5__abc_54027_n859), .Y(u5__abc_54027_n861_1) );
  OR2X2 OR2X2_4783 ( .A(u5_timer_is_zero), .B(u5_mc_le), .Y(u5__abc_54027_n862) );
  OR2X2 OR2X2_4784 ( .A(u5__abc_54027_n862), .B(u5_timer_0_), .Y(u5__abc_54027_n863) );
  OR2X2 OR2X2_4785 ( .A(u5__abc_54027_n864), .B(u5__abc_54027_n865), .Y(u5__abc_54027_n866) );
  OR2X2 OR2X2_4786 ( .A(u5__abc_54027_n872), .B(u5__abc_54027_n873), .Y(u5__abc_54027_n874) );
  OR2X2 OR2X2_4787 ( .A(u5__abc_54027_n858), .B(u5__abc_54027_n874), .Y(u5__abc_54027_n875) );
  OR2X2 OR2X2_4788 ( .A(u5__abc_54027_n875), .B(u5__abc_54027_n866), .Y(u5__abc_54027_n876_1) );
  OR2X2 OR2X2_4789 ( .A(u5__abc_54027_n878), .B(u5__abc_54027_n856), .Y(u5__abc_54027_n879) );
  OR2X2 OR2X2_479 ( .A(u0__abc_49347_n1183_1_bF_buf0), .B(1'b0), .Y(u0__abc_49347_n2172) );
  OR2X2 OR2X2_4790 ( .A(u5__abc_54027_n565_bF_buf0), .B(tms_s_17_), .Y(u5__abc_54027_n884) );
  OR2X2 OR2X2_4791 ( .A(u5__abc_54027_n885), .B(u5__abc_54027_n883), .Y(u5__abc_54027_n886) );
  OR2X2 OR2X2_4792 ( .A(u5__abc_54027_n880), .B(u5__abc_54027_n886), .Y(u5__abc_54027_n887_1) );
  OR2X2 OR2X2_4793 ( .A(u5__abc_54027_n565_bF_buf4), .B(tms_s_20_), .Y(u5__abc_54027_n888) );
  OR2X2 OR2X2_4794 ( .A(u5__abc_54027_n888), .B(u5__abc_54027_n882_1), .Y(u5__abc_54027_n889) );
  OR2X2 OR2X2_4795 ( .A(u5__abc_54027_n565_bF_buf3), .B(tms_s_15_), .Y(u5__abc_54027_n893) );
  OR2X2 OR2X2_4796 ( .A(u5__abc_54027_n888), .B(tms_s_15_), .Y(u5__abc_54027_n896_1) );
  OR2X2 OR2X2_4797 ( .A(u5__abc_54027_n898_1), .B(u5__abc_54027_n892), .Y(u5__abc_54027_n899_1) );
  OR2X2 OR2X2_4798 ( .A(u5__abc_54027_n891), .B(u5__abc_54027_n899_1), .Y(u5__abc_54027_n900_1) );
  OR2X2 OR2X2_4799 ( .A(u5__abc_54027_n565_bF_buf2), .B(tms_s_8_), .Y(u5__abc_54027_n908) );
  OR2X2 OR2X2_48 ( .A(lmr_sel_bF_buf6), .B(tms_6_), .Y(_abc_55805_n309) );
  OR2X2 OR2X2_480 ( .A(spec_req_cs_6_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n2173) );
  OR2X2 OR2X2_4800 ( .A(u5__abc_54027_n909), .B(u5__abc_54027_n906_1), .Y(u5__abc_54027_n910) );
  OR2X2 OR2X2_4801 ( .A(u5__abc_54027_n902), .B(u5__abc_54027_n910), .Y(u5__abc_54027_n911) );
  OR2X2 OR2X2_4802 ( .A(u5__abc_54027_n565_bF_buf1), .B(tms_s_12_), .Y(u5__abc_54027_n912) );
  OR2X2 OR2X2_4803 ( .A(u5__abc_54027_n912), .B(u5__abc_54027_n905_1), .Y(u5__abc_54027_n913) );
  OR2X2 OR2X2_4804 ( .A(u5__abc_54027_n565_bF_buf0), .B(tms_s_13_), .Y(u5__abc_54027_n915) );
  OR2X2 OR2X2_4805 ( .A(u5__abc_54027_n565_bF_buf4), .B(tms_s_18_), .Y(u5__abc_54027_n917) );
  OR2X2 OR2X2_4806 ( .A(u5__abc_54027_n917), .B(u5__abc_54027_n583), .Y(u5__abc_54027_n918) );
  OR2X2 OR2X2_4807 ( .A(u5__abc_54027_n565_bF_buf3), .B(tms_s_25_), .Y(u5__abc_54027_n919) );
  OR2X2 OR2X2_4808 ( .A(u5__abc_54027_n919), .B(u5__abc_54027_n859), .Y(u5__abc_54027_n920) );
  OR2X2 OR2X2_4809 ( .A(u5__abc_54027_n924), .B(u5__abc_54027_n923), .Y(u5__abc_54027_n925) );
  OR2X2 OR2X2_481 ( .A(u0__abc_49347_n2175), .B(u0__abc_49347_n2171), .Y(u0__abc_49347_n2176) );
  OR2X2 OR2X2_4810 ( .A(u5__abc_54027_n925), .B(u5__abc_54027_n875), .Y(u5__abc_54027_n926) );
  OR2X2 OR2X2_4811 ( .A(u5__abc_54027_n565_bF_buf2), .B(tms_s_5_), .Y(u5__abc_54027_n929) );
  OR2X2 OR2X2_4812 ( .A(u5__abc_54027_n930), .B(u5__abc_54027_n582), .Y(u5__abc_54027_n931) );
  OR2X2 OR2X2_4813 ( .A(u5__abc_54027_n928), .B(u5__abc_54027_n931), .Y(u5__abc_54027_n932) );
  OR2X2 OR2X2_4814 ( .A(u5__abc_54027_n565_bF_buf1), .B(tms_s_21_), .Y(u5__abc_54027_n935) );
  OR2X2 OR2X2_4815 ( .A(u5__abc_54027_n936), .B(u5__abc_54027_n614), .Y(u5__abc_54027_n937) );
  OR2X2 OR2X2_4816 ( .A(u5__abc_54027_n934), .B(u5__abc_54027_n937), .Y(u5__abc_54027_n938) );
  OR2X2 OR2X2_4817 ( .A(u5__abc_54027_n565_bF_buf0), .B(tms_s_16_), .Y(u5__abc_54027_n939) );
  OR2X2 OR2X2_4818 ( .A(u5__abc_54027_n940), .B(u5__abc_54027_n944), .Y(u5__abc_54027_n945) );
  OR2X2 OR2X2_4819 ( .A(u5__abc_54027_n945), .B(u5__abc_54027_n895_1), .Y(u5__abc_54027_n946) );
  OR2X2 OR2X2_482 ( .A(u0__abc_49347_n2177), .B(u0__abc_49347_n2178), .Y(u0__abc_49347_n2179) );
  OR2X2 OR2X2_4820 ( .A(u5__abc_54027_n943), .B(u5__abc_54027_n947), .Y(u5__abc_54027_n948) );
  OR2X2 OR2X2_4821 ( .A(u5__abc_54027_n939), .B(tms_s_21_), .Y(u5__abc_54027_n949) );
  OR2X2 OR2X2_4822 ( .A(u5__abc_54027_n950), .B(u5__abc_54027_n894), .Y(u5__abc_54027_n951) );
  OR2X2 OR2X2_4823 ( .A(u5__abc_54027_n952), .B(u5__abc_54027_n424), .Y(u5__abc_54027_n953_1) );
  OR2X2 OR2X2_4824 ( .A(u5__abc_54027_n565_bF_buf4), .B(tms_s_1_), .Y(u5__abc_54027_n956) );
  OR2X2 OR2X2_4825 ( .A(u5__abc_54027_n957), .B(u5__abc_54027_n907), .Y(u5__abc_54027_n958) );
  OR2X2 OR2X2_4826 ( .A(u5__abc_54027_n955), .B(u5__abc_54027_n958), .Y(u5__abc_54027_n959) );
  OR2X2 OR2X2_4827 ( .A(u5__abc_54027_n565_bF_buf3), .B(tms_s_9_), .Y(u5__abc_54027_n961) );
  OR2X2 OR2X2_4828 ( .A(u5__abc_54027_n962), .B(u5__abc_54027_n960), .Y(u5__abc_54027_n963) );
  OR2X2 OR2X2_4829 ( .A(u5__abc_54027_n964), .B(u5__abc_54027_n916), .Y(u5_timer_1__FF_INPUT) );
  OR2X2 OR2X2_483 ( .A(u0__abc_49347_n2180_1), .B(u0__abc_49347_n2181), .Y(u0__abc_49347_n2182) );
  OR2X2 OR2X2_4830 ( .A(u5__abc_54027_n565_bF_buf2), .B(tms_s_22_), .Y(u5__abc_54027_n966) );
  OR2X2 OR2X2_4831 ( .A(u5__abc_54027_n966), .B(u5__abc_54027_n882_1), .Y(u5__abc_54027_n967) );
  OR2X2 OR2X2_4832 ( .A(u5__abc_54027_n565_bF_buf1), .B(tms_s_26_), .Y(u5__abc_54027_n969) );
  OR2X2 OR2X2_4833 ( .A(u5__abc_54027_n976), .B(u5__abc_54027_n872), .Y(u5__abc_54027_n977) );
  OR2X2 OR2X2_4834 ( .A(u5__abc_54027_n977), .B(u5__abc_54027_n974), .Y(u5__abc_54027_n978) );
  OR2X2 OR2X2_4835 ( .A(u5__abc_54027_n979), .B(u5__abc_54027_n970), .Y(u5__abc_54027_n980) );
  OR2X2 OR2X2_4836 ( .A(u5__abc_54027_n982), .B(u5__abc_54027_n883), .Y(u5__abc_54027_n983) );
  OR2X2 OR2X2_4837 ( .A(u5__abc_54027_n981), .B(u5__abc_54027_n983), .Y(u5__abc_54027_n984) );
  OR2X2 OR2X2_4838 ( .A(u5__abc_54027_n988), .B(u5__abc_54027_n987), .Y(u5__abc_54027_n989) );
  OR2X2 OR2X2_4839 ( .A(u5__abc_54027_n990), .B(u5__abc_54027_n940), .Y(u5__abc_54027_n991) );
  OR2X2 OR2X2_484 ( .A(u0__abc_49347_n2183), .B(u0__abc_49347_n2184), .Y(u0__abc_49347_n2185) );
  OR2X2 OR2X2_4840 ( .A(u5__abc_54027_n991), .B(u5__abc_54027_n966), .Y(u5__abc_54027_n992) );
  OR2X2 OR2X2_4841 ( .A(u5__abc_54027_n994), .B(u5__abc_54027_n986), .Y(u5__abc_54027_n995) );
  OR2X2 OR2X2_4842 ( .A(u5__abc_54027_n995), .B(u5__abc_54027_n892), .Y(u5__abc_54027_n996) );
  OR2X2 OR2X2_4843 ( .A(u5__abc_54027_n709_1), .B(u5__abc_54027_n850), .Y(u5__abc_54027_n997) );
  OR2X2 OR2X2_4844 ( .A(u5__abc_54027_n565_bF_buf0), .B(tms_s_10_), .Y(u5__abc_54027_n1000_1) );
  OR2X2 OR2X2_4845 ( .A(u5__abc_54027_n1001), .B(u5__abc_54027_n906_1), .Y(u5__abc_54027_n1002) );
  OR2X2 OR2X2_4846 ( .A(u5__abc_54027_n999), .B(u5__abc_54027_n1002), .Y(u5__abc_54027_n1003) );
  OR2X2 OR2X2_4847 ( .A(u5__abc_54027_n565_bF_buf4), .B(tms_s_14_), .Y(u5__abc_54027_n1004) );
  OR2X2 OR2X2_4848 ( .A(u5__abc_54027_n1004), .B(u5__abc_54027_n905_1), .Y(u5__abc_54027_n1005) );
  OR2X2 OR2X2_4849 ( .A(u5__abc_54027_n565_bF_buf3), .B(tms_s_23_), .Y(u5__abc_54027_n1009) );
  OR2X2 OR2X2_485 ( .A(u0__abc_49347_n2187), .B(spec_req_cs_0_bF_buf3), .Y(u0__abc_49347_n2188) );
  OR2X2 OR2X2_4850 ( .A(u5__abc_54027_n1012), .B(u5__abc_54027_n1011), .Y(u5__abc_54027_n1013) );
  OR2X2 OR2X2_4851 ( .A(u5__abc_54027_n1013), .B(u5__abc_54027_n424), .Y(u5__abc_54027_n1014) );
  OR2X2 OR2X2_4852 ( .A(u5__abc_54027_n565_bF_buf2), .B(tms_s_27_), .Y(u5__abc_54027_n1015) );
  OR2X2 OR2X2_4853 ( .A(u5__abc_54027_n1020), .B(u5__abc_54027_n1018), .Y(u5__abc_54027_n1021) );
  OR2X2 OR2X2_4854 ( .A(u5__abc_54027_n1022), .B(u5__abc_54027_n1016), .Y(u5__abc_54027_n1023) );
  OR2X2 OR2X2_4855 ( .A(u5__abc_54027_n1025), .B(u5__abc_54027_n1026), .Y(u5__abc_54027_n1027) );
  OR2X2 OR2X2_4856 ( .A(u5__abc_54027_n1027), .B(u5__abc_54027_n614), .Y(u5__abc_54027_n1028) );
  OR2X2 OR2X2_4857 ( .A(u5__abc_54027_n565_bF_buf1), .B(tms_s_3_), .Y(u5__abc_54027_n1031) );
  OR2X2 OR2X2_4858 ( .A(u5__abc_54027_n1032), .B(u5__abc_54027_n907), .Y(u5__abc_54027_n1033) );
  OR2X2 OR2X2_4859 ( .A(u5__abc_54027_n1030), .B(u5__abc_54027_n1033), .Y(u5__abc_54027_n1034) );
  OR2X2 OR2X2_486 ( .A(u0__abc_49347_n2186), .B(u0__abc_49347_n2188), .Y(u0__abc_49347_n2189) );
  OR2X2 OR2X2_4860 ( .A(u5__abc_54027_n565_bF_buf0), .B(tms_s_11_), .Y(u5__abc_54027_n1035) );
  OR2X2 OR2X2_4861 ( .A(u5__abc_54027_n1036), .B(u5__abc_54027_n960), .Y(u5__abc_54027_n1037) );
  OR2X2 OR2X2_4862 ( .A(u5__abc_54027_n1038), .B(u5__abc_54027_n1007), .Y(u5_timer_3__FF_INPUT) );
  OR2X2 OR2X2_4863 ( .A(u5__abc_54027_n1044), .B(u5__abc_54027_n1042), .Y(u5__abc_54027_n1045) );
  OR2X2 OR2X2_4864 ( .A(u5__abc_54027_n1053_1), .B(u5__abc_54027_n1054), .Y(u5__abc_54027_n1055) );
  OR2X2 OR2X2_4865 ( .A(u5__abc_54027_n1059), .B(u5__abc_54027_n1057), .Y(u5__abc_54027_n1060) );
  OR2X2 OR2X2_4866 ( .A(u5__abc_54027_n1061), .B(u5__abc_54027_n1062), .Y(u5__abc_54027_n1063) );
  OR2X2 OR2X2_4867 ( .A(u5__abc_54027_n565_bF_buf4), .B(tms_s_6_), .Y(u5__abc_54027_n1065) );
  OR2X2 OR2X2_4868 ( .A(u5__abc_54027_n1068), .B(u5__abc_54027_n1072), .Y(u5__abc_54027_n1073) );
  OR2X2 OR2X2_4869 ( .A(u5__abc_54027_n1074), .B(u5__abc_54027_n1066), .Y(u5__abc_54027_n1075) );
  OR2X2 OR2X2_487 ( .A(u0__abc_49347_n1203_bF_buf0), .B(u0_csc0_9_), .Y(u0__abc_49347_n2190) );
  OR2X2 OR2X2_4870 ( .A(u5__abc_54027_n565_bF_buf3), .B(tms_s_7_), .Y(u5__abc_54027_n1077) );
  OR2X2 OR2X2_4871 ( .A(u5__abc_54027_n1081), .B(u5__abc_54027_n1078), .Y(u5__abc_54027_n1082) );
  OR2X2 OR2X2_4872 ( .A(u5__abc_54027_n1087), .B(u5__abc_54027_n369), .Y(u5__abc_54027_n1088) );
  OR2X2 OR2X2_4873 ( .A(u5__abc_54027_n1088), .B(u5__abc_54027_n1084), .Y(u5__abc_54027_n1089) );
  OR2X2 OR2X2_4874 ( .A(u5__abc_54027_n431), .B(u5_cmd_asserted_bF_buf0), .Y(u5__abc_54027_n1091) );
  OR2X2 OR2X2_4875 ( .A(u5_timer2_1_), .B(u5_timer2_0_), .Y(u5__abc_54027_n1096) );
  OR2X2 OR2X2_4876 ( .A(u5__abc_54027_n1096), .B(u5_timer2_2_), .Y(u5__abc_54027_n1097) );
  OR2X2 OR2X2_4877 ( .A(u5__abc_54027_n1097), .B(u5_timer2_3_), .Y(u5__abc_54027_n1098) );
  OR2X2 OR2X2_4878 ( .A(u5__abc_54027_n1098), .B(u5_timer2_4_), .Y(u5__abc_54027_n1099) );
  OR2X2 OR2X2_4879 ( .A(u5__abc_54027_n1099), .B(u5_timer2_5_), .Y(u5__abc_54027_n1100) );
  OR2X2 OR2X2_488 ( .A(u0__abc_49347_n2192), .B(u0__abc_49347_n2170), .Y(u0_sp_csc_9__FF_INPUT) );
  OR2X2 OR2X2_4880 ( .A(u5__abc_54027_n1100), .B(u5_timer2_6_), .Y(u5__abc_54027_n1101) );
  OR2X2 OR2X2_4881 ( .A(u5__abc_54027_n1101), .B(u5_timer2_7_), .Y(u5__abc_54027_n1102) );
  OR2X2 OR2X2_4882 ( .A(u5__abc_54027_n1102), .B(u5_timer2_8_), .Y(u5__abc_54027_n1103) );
  OR2X2 OR2X2_4883 ( .A(u5__abc_54027_n1104), .B(u5__abc_54027_n1108), .Y(u5__abc_54027_n1109) );
  OR2X2 OR2X2_4884 ( .A(u5__abc_54027_n888), .B(u5__abc_54027_n658), .Y(u5__abc_54027_n1113) );
  OR2X2 OR2X2_4885 ( .A(u5__abc_54027_n1115), .B(u5__abc_54027_n1094), .Y(u5__abc_54027_n1116) );
  OR2X2 OR2X2_4886 ( .A(u5__abc_54027_n1117), .B(u5__abc_54027_n1085), .Y(u5_timer2_0__FF_INPUT) );
  OR2X2 OR2X2_4887 ( .A(u5__abc_54027_n1119), .B(u5__abc_54027_n1120), .Y(u5__abc_54027_n1121) );
  OR2X2 OR2X2_4888 ( .A(u5__abc_54027_n1125), .B(u5__abc_54027_n654_1), .Y(u5__abc_54027_n1126) );
  OR2X2 OR2X2_4889 ( .A(u5__abc_54027_n1126), .B(u5__abc_54027_n1123), .Y(u5__abc_54027_n1127) );
  OR2X2 OR2X2_489 ( .A(u0__abc_49347_n1183_1_bF_buf5), .B(1'b0), .Y(u0__abc_49347_n2196) );
  OR2X2 OR2X2_4890 ( .A(u5__abc_54027_n908), .B(u5__abc_54027_n655), .Y(u5__abc_54027_n1128) );
  OR2X2 OR2X2_4891 ( .A(u5__abc_54027_n1129), .B(u5__abc_54027_n657_1), .Y(u5__abc_54027_n1130) );
  OR2X2 OR2X2_4892 ( .A(u5__abc_54027_n935), .B(u5__abc_54027_n658), .Y(u5__abc_54027_n1131) );
  OR2X2 OR2X2_4893 ( .A(u5__abc_54027_n1132), .B(u5__abc_54027_n1110), .Y(u5__abc_54027_n1133) );
  OR2X2 OR2X2_4894 ( .A(u5__abc_54027_n939), .B(u5__abc_54027_n1111), .Y(u5__abc_54027_n1134) );
  OR2X2 OR2X2_4895 ( .A(u5__abc_54027_n1135), .B(u5__abc_54027_n1093), .Y(u5__abc_54027_n1136) );
  OR2X2 OR2X2_4896 ( .A(u5__abc_54027_n915), .B(u5__abc_54027_n1092), .Y(u5__abc_54027_n1137) );
  OR2X2 OR2X2_4897 ( .A(u5__abc_54027_n1139), .B(u5__abc_54027_n1140), .Y(u5_timer2_1__FF_INPUT) );
  OR2X2 OR2X2_4898 ( .A(u5__abc_54027_n917), .B(u5__abc_54027_n1142), .Y(u5__abc_54027_n1143) );
  OR2X2 OR2X2_4899 ( .A(u5__abc_54027_n1145), .B(u5__abc_54027_n1146), .Y(u5__abc_54027_n1147) );
  OR2X2 OR2X2_49 ( .A(_abc_55805_n240_bF_buf2), .B(sp_tms_7_), .Y(_abc_55805_n311) );
  OR2X2 OR2X2_490 ( .A(spec_req_cs_6_bF_buf2), .B(1'b0), .Y(u0__abc_49347_n2197) );
  OR2X2 OR2X2_4900 ( .A(u5__abc_54027_n1144), .B(u5__abc_54027_n1149), .Y(u5__abc_54027_n1150) );
  OR2X2 OR2X2_4901 ( .A(u5__abc_54027_n1151), .B(u5__abc_54027_n1152), .Y(u5__abc_54027_n1153) );
  OR2X2 OR2X2_4902 ( .A(u5__abc_54027_n1153), .B(u5__abc_54027_n657_1), .Y(u5__abc_54027_n1154) );
  OR2X2 OR2X2_4903 ( .A(u5__abc_54027_n966), .B(u5__abc_54027_n658), .Y(u5__abc_54027_n1155) );
  OR2X2 OR2X2_4904 ( .A(u5__abc_54027_n1157), .B(u5__abc_54027_n1158), .Y(u5__abc_54027_n1159) );
  OR2X2 OR2X2_4905 ( .A(u5__abc_54027_n1161), .B(u5__abc_54027_n1089), .Y(u5__abc_54027_n1162) );
  OR2X2 OR2X2_4906 ( .A(u5__abc_54027_n1160), .B(u5__abc_54027_n1162), .Y(u5__abc_54027_n1163) );
  OR2X2 OR2X2_4907 ( .A(u5__abc_54027_n1165), .B(u5__abc_54027_n1166), .Y(u5__abc_54027_n1167) );
  OR2X2 OR2X2_4908 ( .A(u5__abc_54027_n1170), .B(u5__abc_54027_n1169), .Y(u5__abc_54027_n1171) );
  OR2X2 OR2X2_4909 ( .A(u5__abc_54027_n1171), .B(u5__abc_54027_n654_1), .Y(u5__abc_54027_n1172) );
  OR2X2 OR2X2_491 ( .A(u0__abc_49347_n2199), .B(u0__abc_49347_n2195), .Y(u0__abc_49347_n2200) );
  OR2X2 OR2X2_4910 ( .A(u5__abc_54027_n1000_1), .B(u5__abc_54027_n655), .Y(u5__abc_54027_n1173) );
  OR2X2 OR2X2_4911 ( .A(u5__abc_54027_n1174), .B(u5__abc_54027_n657_1), .Y(u5__abc_54027_n1175) );
  OR2X2 OR2X2_4912 ( .A(u5__abc_54027_n1009), .B(u5__abc_54027_n658), .Y(u5__abc_54027_n1176) );
  OR2X2 OR2X2_4913 ( .A(u5__abc_54027_n1179), .B(u5__abc_54027_n1093), .Y(u5__abc_54027_n1180) );
  OR2X2 OR2X2_4914 ( .A(u5__abc_54027_n1178), .B(u5__abc_54027_n1180), .Y(u5__abc_54027_n1181) );
  OR2X2 OR2X2_4915 ( .A(u5__abc_54027_n893), .B(u5__abc_54027_n1092), .Y(u5__abc_54027_n1182) );
  OR2X2 OR2X2_4916 ( .A(u5__abc_54027_n1184), .B(u5__abc_54027_n1185), .Y(u5_timer2_3__FF_INPUT) );
  OR2X2 OR2X2_4917 ( .A(u5__abc_54027_n566_1), .B(u5__abc_54027_n1111), .Y(u5__abc_54027_n1189) );
  OR2X2 OR2X2_4918 ( .A(u5__abc_54027_n1191), .B(u5__abc_54027_n1192), .Y(u5__abc_54027_n1193) );
  OR2X2 OR2X2_4919 ( .A(u5__abc_54027_n1190), .B(u5__abc_54027_n1195), .Y(u5__abc_54027_n1196) );
  OR2X2 OR2X2_492 ( .A(u0__abc_49347_n2201), .B(u0__abc_49347_n2202), .Y(u0__abc_49347_n2203) );
  OR2X2 OR2X2_4920 ( .A(u5__abc_54027_n1197), .B(u5__abc_54027_n1198), .Y(u5__abc_54027_n1199) );
  OR2X2 OR2X2_4921 ( .A(u5__abc_54027_n1201), .B(u5__abc_54027_n1110), .Y(u5__abc_54027_n1202) );
  OR2X2 OR2X2_4922 ( .A(u5__abc_54027_n1200), .B(u5__abc_54027_n1202), .Y(u5__abc_54027_n1203) );
  OR2X2 OR2X2_4923 ( .A(u5__abc_54027_n1205_1), .B(u5__abc_54027_n1187), .Y(u5_timer2_4__FF_INPUT) );
  OR2X2 OR2X2_4924 ( .A(u5__abc_54027_n1209), .B(u5__abc_54027_n1210), .Y(u5__abc_54027_n1211) );
  OR2X2 OR2X2_4925 ( .A(u5__abc_54027_n1214), .B(u5__abc_54027_n1213), .Y(u5__abc_54027_n1215) );
  OR2X2 OR2X2_4926 ( .A(u5__abc_54027_n1216), .B(u5__abc_54027_n1208), .Y(u5__abc_54027_n1217) );
  OR2X2 OR2X2_4927 ( .A(u5__abc_54027_n1219), .B(u5__abc_54027_n1207), .Y(u5_timer2_5__FF_INPUT) );
  OR2X2 OR2X2_4928 ( .A(u5__abc_54027_n1222), .B(u5__abc_54027_n1223), .Y(u5__abc_54027_n1224) );
  OR2X2 OR2X2_4929 ( .A(u5__abc_54027_n1225), .B(u5__abc_54027_n1124), .Y(u5__abc_54027_n1226) );
  OR2X2 OR2X2_493 ( .A(u0__abc_49347_n2204), .B(u0__abc_49347_n2205), .Y(u0__abc_49347_n2206) );
  OR2X2 OR2X2_4930 ( .A(u5__abc_54027_n929), .B(u5__abc_54027_n1106), .Y(u5__abc_54027_n1228) );
  OR2X2 OR2X2_4931 ( .A(u5__abc_54027_n1230), .B(u5__abc_54027_n1221), .Y(u5_timer2_6__FF_INPUT) );
  OR2X2 OR2X2_4932 ( .A(u5__abc_54027_n1065), .B(u5__abc_54027_n1106), .Y(u5__abc_54027_n1233_1) );
  OR2X2 OR2X2_4933 ( .A(u5__abc_54027_n1236), .B(u5__abc_54027_n1124), .Y(u5__abc_54027_n1237) );
  OR2X2 OR2X2_4934 ( .A(u5__abc_54027_n1235_1), .B(u5__abc_54027_n1237), .Y(u5__abc_54027_n1238) );
  OR2X2 OR2X2_4935 ( .A(u5__abc_54027_n1240), .B(u5__abc_54027_n1232), .Y(u5_timer2_7__FF_INPUT) );
  OR2X2 OR2X2_4936 ( .A(u5__abc_54027_n1077), .B(u5__abc_54027_n1106), .Y(u5__abc_54027_n1243) );
  OR2X2 OR2X2_4937 ( .A(u5__abc_54027_n1244), .B(u5__abc_54027_n1124), .Y(u5__abc_54027_n1245) );
  OR2X2 OR2X2_4938 ( .A(u5__abc_54027_n1247), .B(u5__abc_54027_n1242), .Y(u5_timer2_8__FF_INPUT) );
  OR2X2 OR2X2_4939 ( .A(u5__abc_54027_n643_1), .B(dv), .Y(u5__abc_54027_n1250) );
  OR2X2 OR2X2_494 ( .A(u0__abc_49347_n2207), .B(u0__abc_49347_n2208), .Y(u0__abc_49347_n2209) );
  OR2X2 OR2X2_4940 ( .A(u5__abc_54027_n1251), .B(u5__abc_54027_n1249), .Y(u5__abc_54027_n1252) );
  OR2X2 OR2X2_4941 ( .A(u5__abc_54027_n1253), .B(u5__abc_54027_n637), .Y(u5__abc_54027_n1254) );
  OR2X2 OR2X2_4942 ( .A(u5__abc_54027_n1252), .B(u5_ack_cnt_0_), .Y(u5__abc_54027_n1256) );
  OR2X2 OR2X2_4943 ( .A(u5__abc_54027_n1259), .B(u5__abc_54027_n1260), .Y(u5__abc_54027_n1261) );
  OR2X2 OR2X2_4944 ( .A(u5__abc_54027_n1262), .B(u5__abc_54027_n636), .Y(u5__abc_54027_n1263) );
  OR2X2 OR2X2_4945 ( .A(u5__abc_54027_n1261), .B(u5_ack_cnt_1_), .Y(u5__abc_54027_n1264) );
  OR2X2 OR2X2_4946 ( .A(u5__abc_54027_n1267), .B(u5__abc_54027_n1269), .Y(u5__abc_54027_n1270) );
  OR2X2 OR2X2_4947 ( .A(u5__abc_54027_n1271), .B(u5__abc_54027_n635), .Y(u5__abc_54027_n1272) );
  OR2X2 OR2X2_4948 ( .A(u5__abc_54027_n1270), .B(u5_ack_cnt_2_), .Y(u5__abc_54027_n1273) );
  OR2X2 OR2X2_4949 ( .A(u5__abc_54027_n634), .B(u5__abc_54027_n640), .Y(u5__abc_54027_n1276) );
  OR2X2 OR2X2_495 ( .A(u0__abc_49347_n2211), .B(spec_req_cs_0_bF_buf2), .Y(u0__abc_49347_n2212) );
  OR2X2 OR2X2_4950 ( .A(dv), .B(u5__abc_54027_n1276), .Y(u5__abc_54027_n1277) );
  OR2X2 OR2X2_4951 ( .A(u5__abc_54027_n1279), .B(u5__abc_54027_n1278), .Y(u5__abc_54027_n1280) );
  OR2X2 OR2X2_4952 ( .A(u5_mc_le), .B(u5_cmd_asserted_bF_buf3), .Y(u5__abc_54027_n1285) );
  OR2X2 OR2X2_4953 ( .A(u5_mc_le_FF_INPUT), .B(u5_cmd_asserted2), .Y(u5__abc_54027_n1286) );
  OR2X2 OR2X2_4954 ( .A(u5__abc_54027_n1289), .B(u5__abc_54027_n1288), .Y(u5_cmd_asserted_FF_INPUT) );
  OR2X2 OR2X2_4955 ( .A(u5_mc_le), .B(u5_mc_adv_r1), .Y(u5__abc_54027_n1291) );
  OR2X2 OR2X2_4956 ( .A(u5_mc_le_FF_INPUT), .B(u5_mc_adv_r), .Y(u5__abc_54027_n1292) );
  OR2X2 OR2X2_4957 ( .A(u5__abc_54027_n1300), .B(u5__abc_54027_n477), .Y(u5__abc_54027_n1301) );
  OR2X2 OR2X2_4958 ( .A(mc_adv_d), .B(u5_mc_le), .Y(u5__abc_54027_n1303) );
  OR2X2 OR2X2_4959 ( .A(u5_mc_le_FF_INPUT), .B(u5_mc_adv_r1), .Y(u5__abc_54027_n1304) );
  OR2X2 OR2X2_496 ( .A(u0__abc_49347_n2210), .B(u0__abc_49347_n2212), .Y(u0__abc_49347_n2213) );
  OR2X2 OR2X2_4960 ( .A(u5__abc_54027_n678), .B(u5_wb_cycle), .Y(u5__abc_54027_n1307) );
  OR2X2 OR2X2_4961 ( .A(u5__abc_54027_n1310), .B(u5__abc_54027_n1306), .Y(u5__abc_54027_n1311) );
  OR2X2 OR2X2_4962 ( .A(u5__abc_54027_n1320), .B(u5__abc_54027_n1322), .Y(u5__abc_54027_n1323) );
  OR2X2 OR2X2_4963 ( .A(u5__abc_54027_n1329), .B(u5__abc_54027_n1332), .Y(u5__abc_54027_n1333) );
  OR2X2 OR2X2_4964 ( .A(u5__abc_54027_n678), .B(u5__abc_54027_n1340), .Y(u5__abc_54027_n1341_1) );
  OR2X2 OR2X2_4965 ( .A(u5__abc_54027_n649), .B(u5__abc_54027_n1343), .Y(u5__abc_54027_n1344) );
  OR2X2 OR2X2_4966 ( .A(u5__abc_54027_n1348), .B(u5__abc_54027_n382), .Y(u5__abc_54027_n1349) );
  OR2X2 OR2X2_4967 ( .A(u5__abc_54027_n1358), .B(u5_cmd_asserted2), .Y(u5__abc_54027_n1359) );
  OR2X2 OR2X2_4968 ( .A(u5__abc_54027_n1357), .B(u5__abc_54027_n1359), .Y(u5__abc_54027_n1360) );
  OR2X2 OR2X2_4969 ( .A(u5__abc_54027_n1355), .B(u5__abc_54027_n1360), .Y(u5__abc_54027_n1361) );
  OR2X2 OR2X2_497 ( .A(u0__abc_49347_n1203_bF_buf5), .B(u0_csc0_10_), .Y(u0__abc_49347_n2214) );
  OR2X2 OR2X2_4970 ( .A(csc_s_4_), .B(csc_s_5_bF_buf0), .Y(u5__abc_54027_n1369) );
  OR2X2 OR2X2_4971 ( .A(u5__abc_54027_n1371), .B(u5__abc_54027_n1369), .Y(u5__abc_54027_n1372) );
  OR2X2 OR2X2_4972 ( .A(u5__abc_54027_n391), .B(u5__abc_54027_n1299), .Y(u5__abc_54027_n1374) );
  OR2X2 OR2X2_4973 ( .A(u5__abc_54027_n1300), .B(u5__abc_54027_n1376), .Y(u5__abc_54027_n1377) );
  OR2X2 OR2X2_4974 ( .A(u5__abc_54027_n1391_1), .B(u5__abc_54027_n1392), .Y(u5__abc_54027_n1393) );
  OR2X2 OR2X2_4975 ( .A(u5__abc_54027_n363), .B(u5__abc_54027_n1312_1), .Y(u5__abc_54027_n1400) );
  OR2X2 OR2X2_4976 ( .A(u5__abc_54027_n545_1), .B(u1_wb_write_go), .Y(u5__abc_54027_n1402) );
  OR2X2 OR2X2_4977 ( .A(u5__abc_54027_n1401), .B(u5__abc_54027_n1403), .Y(u5__abc_54027_n1404) );
  OR2X2 OR2X2_4978 ( .A(u5__abc_54027_n1383_1), .B(u1_wb_write_go), .Y(u5__abc_54027_n1413) );
  OR2X2 OR2X2_4979 ( .A(u5__abc_54027_n1401), .B(u5__abc_54027_n1413), .Y(u5__abc_54027_n1414) );
  OR2X2 OR2X2_498 ( .A(u0__abc_49347_n2216_1), .B(u0__abc_49347_n2194), .Y(u0_sp_csc_10__FF_INPUT) );
  OR2X2 OR2X2_4980 ( .A(u5__abc_54027_n1418), .B(u5_wb_wait_r), .Y(u5__abc_54027_n1419) );
  OR2X2 OR2X2_4981 ( .A(u5__abc_54027_n644), .B(u5__abc_54027_n619), .Y(u5__abc_54027_n1421) );
  OR2X2 OR2X2_4982 ( .A(u5__abc_54027_n1425), .B(u5__abc_54027_n1424), .Y(u5__abc_54027_n1426) );
  OR2X2 OR2X2_4983 ( .A(u5__abc_54027_n1426), .B(u5__abc_54027_n1428), .Y(u5__abc_54027_n1429) );
  OR2X2 OR2X2_4984 ( .A(u5__abc_54027_n436), .B(u5__abc_54027_n1435), .Y(u5__abc_54027_n1436) );
  OR2X2 OR2X2_4985 ( .A(u5__abc_54027_n1440), .B(u5__abc_54027_n1438_1), .Y(u5__abc_54027_n1441) );
  OR2X2 OR2X2_4986 ( .A(u5__abc_54027_n1443), .B(u5__abc_54027_n1444), .Y(u5__abc_54027_n1445_1) );
  OR2X2 OR2X2_4987 ( .A(u5__abc_54027_n1448_1), .B(u5__abc_54027_n1449), .Y(u5__abc_54027_n1450_1) );
  OR2X2 OR2X2_4988 ( .A(u5__abc_54027_n1452), .B(u5__abc_54027_n366_1), .Y(u5__abc_54027_n1453) );
  OR2X2 OR2X2_4989 ( .A(u5__abc_54027_n1457), .B(u5__abc_54027_n1458), .Y(u5__abc_54027_n1459) );
  OR2X2 OR2X2_499 ( .A(u0__abc_49347_n2728_bF_buf5), .B(1'b0), .Y(u0__abc_49347_n2729) );
  OR2X2 OR2X2_4990 ( .A(u5__abc_54027_n1299), .B(mc_ack_r), .Y(u5__abc_54027_n1462) );
  OR2X2 OR2X2_4991 ( .A(u5__abc_54027_n1461), .B(u5__abc_54027_n1462), .Y(u5__abc_54027_n1463) );
  OR2X2 OR2X2_4992 ( .A(u5__abc_54027_n506), .B(u5_cs_le_r), .Y(u5__abc_54027_n1468) );
  OR2X2 OR2X2_4993 ( .A(u5__abc_54027_n1469), .B(u5__abc_54027_n1299), .Y(u5__abc_54027_n1470) );
  OR2X2 OR2X2_4994 ( .A(u5__abc_54027_n1467_1), .B(u5__abc_54027_n1475), .Y(u5__abc_54027_n1476_1) );
  OR2X2 OR2X2_4995 ( .A(u5__abc_54027_n1480), .B(u5__abc_54027_n1479), .Y(u5__abc_54027_n1481) );
  OR2X2 OR2X2_4996 ( .A(u5__abc_54027_n444), .B(u5__abc_54027_n1312_1), .Y(u5__abc_54027_n1483) );
  OR2X2 OR2X2_4997 ( .A(u5__abc_54027_n1492), .B(u3_wb_read_go), .Y(u5__abc_54027_n1493) );
  OR2X2 OR2X2_4998 ( .A(u5__abc_54027_n1495), .B(u5__abc_54027_n1494), .Y(u5__abc_54027_n1496) );
  OR2X2 OR2X2_4999 ( .A(u5__abc_54027_n1509), .B(u5__abc_54027_n1511), .Y(u5__abc_54027_n1512) );
  OR2X2 OR2X2_5 ( .A(_abc_55805_n243), .B(_abc_55805_n237_1), .Y(_abc_55805_n244_1) );
  OR2X2 OR2X2_50 ( .A(lmr_sel_bF_buf5), .B(tms_7_), .Y(_abc_55805_n312) );
  OR2X2 OR2X2_500 ( .A(1'b0), .B(1'b0), .Y(u0__abc_49347_n2731) );
  OR2X2 OR2X2_5000 ( .A(u5__abc_54027_n1512), .B(u5__abc_54027_n1506), .Y(u5__abc_54027_n1513) );
  OR2X2 OR2X2_5001 ( .A(u5__abc_54027_n1514), .B(u5_wb_wait), .Y(u5__abc_54027_n1515) );
  OR2X2 OR2X2_5002 ( .A(u5__abc_54027_n1519), .B(u5__abc_54027_n1520), .Y(u5__abc_54027_n1521) );
  OR2X2 OR2X2_5003 ( .A(u5__abc_54027_n1524), .B(u5__abc_54027_n1522), .Y(u5__abc_54027_n1525) );
  OR2X2 OR2X2_5004 ( .A(u5__abc_54027_n1525), .B(u5__abc_54027_n1521), .Y(u5__abc_54027_n1526) );
  OR2X2 OR2X2_5005 ( .A(u5__abc_54027_n1526), .B(u5__abc_54027_n1517), .Y(u5__abc_54027_n1527) );
  OR2X2 OR2X2_5006 ( .A(u5__abc_54027_n1513), .B(u5__abc_54027_n1527), .Y(u5__abc_54027_n1528) );
  OR2X2 OR2X2_5007 ( .A(u5__abc_54027_n1533_1), .B(u5__abc_54027_n457), .Y(u5__abc_54027_n1534) );
  OR2X2 OR2X2_5008 ( .A(u5__abc_54027_n1537_1), .B(u5__abc_54027_n1383_1), .Y(u5__abc_54027_n1538) );
  OR2X2 OR2X2_5009 ( .A(u5__abc_54027_n1550), .B(u5__abc_54027_n1554_1), .Y(u5__abc_54027_n1555_1) );
  OR2X2 OR2X2_501 ( .A(u0__abc_49347_n2733), .B(u0__abc_49347_n2727), .Y(u0__abc_49347_n2734) );
  OR2X2 OR2X2_5010 ( .A(u5__abc_54027_n1548), .B(u5__abc_54027_n1556), .Y(u5__abc_54027_n1557) );
  OR2X2 OR2X2_5011 ( .A(u5__abc_54027_n1547_1), .B(u5__abc_54027_n1557), .Y(u5__abc_54027_n1558_1) );
  OR2X2 OR2X2_5012 ( .A(u5__abc_54027_n1402), .B(u5__abc_54027_n519), .Y(u5__abc_54027_n1560) );
  OR2X2 OR2X2_5013 ( .A(u5__abc_54027_n1559), .B(u5__abc_54027_n1561_1), .Y(u5__abc_54027_n1562_1) );
  OR2X2 OR2X2_5014 ( .A(u5__abc_54027_n1575_1), .B(u5__abc_54027_n352), .Y(u5__abc_54027_n1576) );
  OR2X2 OR2X2_5015 ( .A(u5__abc_54027_n1576), .B(u5__abc_54027_n1572_1), .Y(u5__abc_54027_n1577) );
  OR2X2 OR2X2_5016 ( .A(u5__abc_54027_n1580), .B(u5__abc_54027_n1579), .Y(u5__abc_54027_n1581) );
  OR2X2 OR2X2_5017 ( .A(u5__abc_54027_n1589), .B(u5__abc_54027_n1590), .Y(u5__abc_54027_n1591) );
  OR2X2 OR2X2_5018 ( .A(u5__abc_54027_n1595), .B(u5__abc_54027_n1591), .Y(u5__abc_54027_n1596) );
  OR2X2 OR2X2_5019 ( .A(u5__abc_54027_n1607), .B(u5__abc_54027_n1383_1), .Y(u5__abc_54027_n1608) );
  OR2X2 OR2X2_502 ( .A(u0__abc_49347_n2735), .B(u0__abc_49347_n2736), .Y(u0__abc_49347_n2737) );
  OR2X2 OR2X2_5020 ( .A(u5__abc_54027_n1613), .B(u5__abc_54027_n1614), .Y(u5__abc_54027_n1615) );
  OR2X2 OR2X2_5021 ( .A(u5__abc_54027_n641), .B(u5__abc_54027_n1489), .Y(u5__abc_54027_n1619) );
  OR2X2 OR2X2_5022 ( .A(u5__abc_54027_n1491_1), .B(u5__abc_54027_n477), .Y(u5__abc_54027_n1620) );
  OR2X2 OR2X2_5023 ( .A(u5__abc_54027_n1621), .B(u5__abc_54027_n500), .Y(u5__abc_54027_n1622) );
  OR2X2 OR2X2_5024 ( .A(u5__abc_54027_n436), .B(u5__abc_54027_n1433), .Y(u5__abc_54027_n1624) );
  OR2X2 OR2X2_5025 ( .A(u5__abc_54027_n1629), .B(u5_pack_le1_d), .Y(u5__abc_54027_n1630) );
  OR2X2 OR2X2_5026 ( .A(u5__abc_54027_n431), .B(u5_tmr2_done), .Y(u5__abc_54027_n1632) );
  OR2X2 OR2X2_5027 ( .A(u5__abc_54027_n1644), .B(u5__abc_54027_n1333), .Y(u5__abc_54027_n1645) );
  OR2X2 OR2X2_5028 ( .A(u5__abc_54027_n1645), .B(u5__abc_54027_n1558_1), .Y(u5__abc_54027_n1646) );
  OR2X2 OR2X2_5029 ( .A(u5__abc_54027_n1656), .B(u5__abc_54027_n1655), .Y(u5__abc_54027_n1657) );
  OR2X2 OR2X2_503 ( .A(u0__abc_49347_n2738), .B(u0__abc_49347_n2739), .Y(u0__abc_49347_n2740) );
  OR2X2 OR2X2_5030 ( .A(u5__abc_54027_n1661), .B(u5__abc_54027_n1658), .Y(u5__abc_54027_n1662) );
  OR2X2 OR2X2_5031 ( .A(u5__abc_54027_n1654), .B(u5__abc_54027_n1665), .Y(u5__abc_54027_n1666) );
  OR2X2 OR2X2_5032 ( .A(u5__abc_54027_n1666), .B(u5__abc_54027_n1652), .Y(u5__abc_54027_n1667) );
  OR2X2 OR2X2_5033 ( .A(u5__abc_54027_n1646), .B(u5__abc_54027_n1670), .Y(u5__abc_41027_n1846) );
  OR2X2 OR2X2_5034 ( .A(u5__abc_54027_n421), .B(u5__abc_54027_n1676), .Y(u5__abc_54027_n1677) );
  OR2X2 OR2X2_5035 ( .A(u5__abc_54027_n1653), .B(u5__abc_54027_n1677), .Y(u5__abc_54027_n1678) );
  OR2X2 OR2X2_5036 ( .A(u5__abc_54027_n483), .B(u5__abc_54027_n421), .Y(u5__abc_54027_n1685) );
  OR2X2 OR2X2_5037 ( .A(u5__abc_54027_n1557), .B(u5__abc_54027_n1344), .Y(u5__abc_54027_n1689) );
  OR2X2 OR2X2_5038 ( .A(u5__abc_54027_n1690), .B(u5__abc_54027_n1691), .Y(u5__abc_54027_n1692) );
  OR2X2 OR2X2_5039 ( .A(u5__abc_54027_n1692), .B(u5__abc_54027_n1689), .Y(u5__abc_54027_n1693) );
  OR2X2 OR2X2_504 ( .A(u0__abc_49347_n2741), .B(u0__abc_49347_n2742), .Y(u0__abc_49347_n2743) );
  OR2X2 OR2X2_5040 ( .A(u5__abc_54027_n1703), .B(u5__abc_54027_n387_1), .Y(u5__abc_54027_n1704) );
  OR2X2 OR2X2_5041 ( .A(u5__abc_54027_n1371), .B(u5__abc_54027_n1346), .Y(u5__abc_54027_n1706) );
  OR2X2 OR2X2_5042 ( .A(u5__abc_54027_n1709), .B(u5__abc_54027_n1708), .Y(u5__abc_54027_n1710) );
  OR2X2 OR2X2_5043 ( .A(u5__abc_54027_n1713), .B(u5__abc_54027_n1714), .Y(u5__abc_54027_n1715) );
  OR2X2 OR2X2_5044 ( .A(u5__abc_54027_n1723), .B(u5__abc_54027_n1722), .Y(u5__abc_54027_n1724) );
  OR2X2 OR2X2_5045 ( .A(u5__abc_54027_n1728), .B(u5__abc_54027_n1724), .Y(u5__abc_54027_n1729) );
  OR2X2 OR2X2_5046 ( .A(u5__abc_54027_n1743), .B(u5__abc_54027_n1547_1), .Y(u5__abc_54027_n1744) );
  OR2X2 OR2X2_5047 ( .A(u5__abc_54027_n1744), .B(u5__abc_54027_n1693), .Y(u5__abc_54027_n1745) );
  OR2X2 OR2X2_5048 ( .A(u5__abc_54027_n1745), .B(u5__abc_54027_n1688), .Y(u5__abc_41027_n1847) );
  OR2X2 OR2X2_5049 ( .A(u5__abc_54027_n1750), .B(u5_tmr_done), .Y(u5__abc_54027_n1751) );
  OR2X2 OR2X2_505 ( .A(u0__abc_49347_n2745), .B(u0_cs0_bF_buf5), .Y(u0__abc_49347_n2746) );
  OR2X2 OR2X2_5050 ( .A(u5__abc_54027_n438_1), .B(u5__abc_54027_n1756), .Y(u5__abc_54027_n1757) );
  OR2X2 OR2X2_5051 ( .A(u5__abc_54027_n385), .B(u5_tmr2_done), .Y(u5__abc_54027_n1759) );
  OR2X2 OR2X2_5052 ( .A(u5__abc_54027_n1533_1), .B(u5__abc_54027_n305), .Y(u5__abc_54027_n1770) );
  OR2X2 OR2X2_5053 ( .A(u5__abc_54027_n1383_1), .B(u5_ir_cnt_done), .Y(u5__abc_54027_n1771) );
  OR2X2 OR2X2_5054 ( .A(u5__abc_54027_n1333), .B(u5__abc_54027_n1692), .Y(u5__abc_54027_n1784) );
  OR2X2 OR2X2_5055 ( .A(u5__abc_54027_n1784), .B(u5__abc_54027_n1783), .Y(u5__abc_41027_n1848) );
  OR2X2 OR2X2_5056 ( .A(u5__abc_54027_n446_1), .B(u5_cmd_asserted_bF_buf0), .Y(u5__abc_54027_n1800) );
  OR2X2 OR2X2_5057 ( .A(u5__abc_54027_n1826), .B(u5__abc_54027_n1824), .Y(u5__abc_54027_n1827) );
  OR2X2 OR2X2_5058 ( .A(u5__abc_54027_n522), .B(u5__abc_54027_n852), .Y(u5__abc_54027_n1837) );
  OR2X2 OR2X2_5059 ( .A(u5__abc_54027_n1840), .B(u5__abc_54027_n1838), .Y(u5__abc_54027_n1841) );
  OR2X2 OR2X2_506 ( .A(u0__abc_49347_n2744), .B(u0__abc_49347_n2746), .Y(u0__abc_49347_n2747) );
  OR2X2 OR2X2_5060 ( .A(u5__abc_54027_n1841), .B(u5__abc_54027_n1837), .Y(u5__abc_54027_n1842) );
  OR2X2 OR2X2_5061 ( .A(u5__abc_54027_n1836), .B(u5__abc_54027_n1842), .Y(u5__abc_54027_n1843) );
  OR2X2 OR2X2_5062 ( .A(u5__abc_54027_n1843), .B(u5__abc_54027_n1834), .Y(u5__abc_54027_n1844) );
  OR2X2 OR2X2_5063 ( .A(u5__abc_54027_n1846), .B(u5__abc_54027_n1845), .Y(u5__abc_54027_n1847) );
  OR2X2 OR2X2_5064 ( .A(u5__abc_54027_n1844), .B(u5__abc_54027_n1847), .Y(u5__abc_54027_n1848) );
  OR2X2 OR2X2_5065 ( .A(u5__abc_54027_n1848), .B(u5__abc_54027_n1528), .Y(u5__abc_54027_n1849) );
  OR2X2 OR2X2_5066 ( .A(u5__abc_54027_n1849), .B(u5__abc_54027_n1833), .Y(u5__abc_54027_n1850) );
  OR2X2 OR2X2_5067 ( .A(u5__abc_54027_n1832), .B(u5__abc_54027_n1850), .Y(u5__abc_54027_n1851) );
  OR2X2 OR2X2_5068 ( .A(u5__abc_54027_n1828), .B(u5__abc_54027_n1851), .Y(u5__abc_41027_n1851) );
  OR2X2 OR2X2_5069 ( .A(u5__abc_54027_n1853), .B(u5__abc_54027_n397), .Y(u5_pack_le0_d) );
  OR2X2 OR2X2_507 ( .A(u0__abc_49347_n2748_bF_buf5), .B(u0_tms0_0_), .Y(u0__abc_49347_n2749) );
  OR2X2 OR2X2_5070 ( .A(u5__abc_54027_n1856), .B(u5__abc_54027_n477), .Y(u5__abc_54027_n1857) );
  OR2X2 OR2X2_5071 ( .A(u5__abc_54027_n1855), .B(u5_cke_r), .Y(u5__abc_54027_n1858) );
  OR2X2 OR2X2_5072 ( .A(u5__abc_54027_n1861), .B(u5__abc_54027_n1862), .Y(u5__abc_54027_n1863) );
  OR2X2 OR2X2_5073 ( .A(u5__abc_54027_n1860), .B(u5__abc_54027_n1863), .Y(u5_cke_d) );
  OR2X2 OR2X2_5074 ( .A(u5__abc_54027_n445), .B(u5__abc_54027_n1478), .Y(u5__abc_54027_n1865) );
  OR2X2 OR2X2_5075 ( .A(u5__abc_54027_n1865), .B(u5__abc_54027_n460), .Y(u5__abc_54027_n1866) );
  OR2X2 OR2X2_5076 ( .A(u5__abc_54027_n1866), .B(u5__abc_54027_n1798), .Y(u5_lmr_ack_d) );
  OR2X2 OR2X2_5077 ( .A(u5__abc_54027_n437_1), .B(u5__abc_54027_n1520), .Y(u5__abc_54027_n1870) );
  OR2X2 OR2X2_5078 ( .A(u5__abc_54027_n1870), .B(u5__abc_54027_n369), .Y(u5__abc_54027_n1871) );
  OR2X2 OR2X2_5079 ( .A(u5__abc_54027_n1871), .B(u5__abc_54027_n1869), .Y(u5__abc_54027_n1872) );
  OR2X2 OR2X2_508 ( .A(u0__abc_49347_n2751), .B(u0__abc_49347_n2722), .Y(u0_tms_0__FF_INPUT) );
  OR2X2 OR2X2_5080 ( .A(u5__abc_54027_n1872), .B(u5__abc_54027_n1868), .Y(u5__abc_54027_n1873) );
  OR2X2 OR2X2_5081 ( .A(u5__abc_54027_n1873), .B(u5__abc_54027_n1595), .Y(mc_adsc_d) );
  OR2X2 OR2X2_5082 ( .A(u5__abc_54027_n1444), .B(u5__abc_54027_n1809), .Y(u5__abc_54027_n1875) );
  OR2X2 OR2X2_5083 ( .A(u5__abc_54027_n1875), .B(u5__abc_54027_n1881), .Y(mc_bg_d) );
  OR2X2 OR2X2_5084 ( .A(u5__abc_54027_n1884), .B(u5__abc_54027_n1883), .Y(u5__abc_54027_n1885) );
  OR2X2 OR2X2_5085 ( .A(u5__abc_54027_n1886), .B(u5_wb_stb_first), .Y(u5__abc_54027_n1887) );
  OR2X2 OR2X2_5086 ( .A(u5__abc_54027_n1890), .B(u5__abc_54027_n1891), .Y(u5__abc_54027_n1892) );
  OR2X2 OR2X2_5087 ( .A(u5__abc_54027_n1894), .B(u5__abc_54027_n1520), .Y(u5__abc_54027_n1895) );
  OR2X2 OR2X2_5088 ( .A(u5__abc_54027_n1444), .B(u5__abc_54027_n873), .Y(u5__abc_54027_n1897) );
  OR2X2 OR2X2_5089 ( .A(u5__abc_54027_n355), .B(u5__abc_54027_n1708), .Y(u5__abc_54027_n1898) );
  OR2X2 OR2X2_509 ( .A(u0__abc_49347_n2728_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n2755) );
  OR2X2 OR2X2_5090 ( .A(u5__abc_54027_n1898), .B(u5__abc_54027_n1589), .Y(u5__abc_54027_n1899) );
  OR2X2 OR2X2_5091 ( .A(u5__abc_54027_n1899), .B(u5__abc_54027_n1897), .Y(u5__abc_54027_n1900) );
  OR2X2 OR2X2_5092 ( .A(u5__abc_54027_n1900), .B(u5__abc_54027_n1896), .Y(u5__abc_54027_n1901) );
  OR2X2 OR2X2_5093 ( .A(u5__abc_54027_n1901), .B(u5__abc_54027_n1893), .Y(u5__abc_54027_n1902) );
  OR2X2 OR2X2_5094 ( .A(u5__abc_54027_n1888), .B(u5__abc_54027_n1902), .Y(cs_le_d) );
  OR2X2 OR2X2_5095 ( .A(u5__abc_54027_n1906), .B(u5__abc_54027_n1443), .Y(u5_mc_c_oe_d) );
  OR2X2 OR2X2_5096 ( .A(u5__abc_54027_n1908), .B(u5__abc_54027_n348), .Y(u5__abc_54027_n1909) );
  OR2X2 OR2X2_5097 ( .A(u5__abc_54027_n1909), .B(u5__abc_54027_n461_1), .Y(bank_clr_all) );
  OR2X2 OR2X2_5098 ( .A(u5__abc_54027_n573), .B(u5__abc_54027_n1911), .Y(bank_clr) );
  OR2X2 OR2X2_5099 ( .A(u5__abc_54027_n1913), .B(u5__abc_54027_n1914), .Y(u5__abc_54027_n1915) );
  OR2X2 OR2X2_51 ( .A(_abc_55805_n240_bF_buf1), .B(sp_tms_8_), .Y(_abc_55805_n314) );
  OR2X2 OR2X2_510 ( .A(1'b0), .B(1'b0), .Y(u0__abc_49347_n2756) );
  OR2X2 OR2X2_5100 ( .A(u5__abc_54027_n582), .B(u5__abc_54027_n646), .Y(row_sel) );
  OR2X2 OR2X2_5101 ( .A(u5__abc_54027_n1919), .B(u5_ap_en), .Y(u5__abc_54027_n1920) );
  OR2X2 OR2X2_5102 ( .A(u5__abc_54027_n1925), .B(u5__abc_54027_n1839), .Y(u5__abc_54027_n1926) );
  OR2X2 OR2X2_5103 ( .A(u5__abc_54027_n1918), .B(u5_ap_en), .Y(u5__abc_54027_n1928) );
  OR2X2 OR2X2_5104 ( .A(u5__abc_54027_n1909), .B(u5__abc_54027_n1929), .Y(u5__abc_54027_n1930) );
  OR2X2 OR2X2_5105 ( .A(u5__abc_54027_n1930), .B(u5__abc_54027_n1927), .Y(u5__abc_54027_n1931) );
  OR2X2 OR2X2_5106 ( .A(u5__abc_54027_n1931), .B(u5__abc_54027_n1924), .Y(cmd_a10) );
  OR2X2 OR2X2_5107 ( .A(u5__abc_54027_n1993), .B(u5__abc_54027_n1991), .Y(u5__abc_54027_n1994) );
  OR2X2 OR2X2_5108 ( .A(u5__abc_54027_n1994), .B(u5__abc_54027_n1306), .Y(u5__abc_54027_n1995) );
  OR2X2 OR2X2_5109 ( .A(u5__abc_54027_n614), .B(u5__abc_54027_n313_1), .Y(u5__abc_54027_n2006) );
  OR2X2 OR2X2_511 ( .A(u0__abc_49347_n2758), .B(u0__abc_49347_n2754), .Y(u0__abc_49347_n2759) );
  OR2X2 OR2X2_5110 ( .A(u5__abc_54027_n457), .B(u5__abc_54027_n1312_1), .Y(u5__abc_54027_n2009) );
  OR2X2 OR2X2_5111 ( .A(u5__abc_54027_n2010), .B(u5__abc_54027_n1440), .Y(u5_susp_sel_r_FF_INPUT) );
  OR2X2 OR2X2_5112 ( .A(u5__abc_54027_n588), .B(u5__abc_54027_n2014), .Y(u5_wb_cycle_FF_INPUT) );
  OR2X2 OR2X2_5113 ( .A(u5__abc_54027_n632_1), .B(u1_wb_write_go), .Y(u5__abc_54027_n2017) );
  OR2X2 OR2X2_5114 ( .A(u5__abc_54027_n2019), .B(u5__abc_54027_n2018), .Y(u5__abc_54027_n2020) );
  OR2X2 OR2X2_5115 ( .A(u5__abc_54027_n2021), .B(u5__abc_54027_n2016), .Y(u5_wr_cycle_FF_INPUT) );
  OR2X2 OR2X2_5116 ( .A(u6__abc_56056_n138_1), .B(u6__abc_56056_n133), .Y(u6__abc_56056_n139_1) );
  OR2X2 OR2X2_5117 ( .A(u6__abc_56056_n146_1), .B(u6__abc_56056_n151), .Y(u6_wb_ack_o_FF_INPUT) );
  OR2X2 OR2X2_5118 ( .A(u6__abc_56056_n144_bF_buf4), .B(rf_dout_0_), .Y(u6__abc_56056_n153) );
  OR2X2 OR2X2_5119 ( .A(u6__abc_56056_n154_bF_buf4), .B(mem_dout_0_), .Y(u6__abc_56056_n155_1) );
  OR2X2 OR2X2_512 ( .A(u0__abc_49347_n2760), .B(u0__abc_49347_n2761), .Y(u0__abc_49347_n2762) );
  OR2X2 OR2X2_5120 ( .A(u6__abc_56056_n144_bF_buf2), .B(rf_dout_1_), .Y(u6__abc_56056_n157_1) );
  OR2X2 OR2X2_5121 ( .A(u6__abc_56056_n154_bF_buf3), .B(mem_dout_1_), .Y(u6__abc_56056_n158) );
  OR2X2 OR2X2_5122 ( .A(u6__abc_56056_n144_bF_buf1), .B(rf_dout_2_), .Y(u6__abc_56056_n160) );
  OR2X2 OR2X2_5123 ( .A(u6__abc_56056_n154_bF_buf2), .B(mem_dout_2_), .Y(u6__abc_56056_n161) );
  OR2X2 OR2X2_5124 ( .A(u6__abc_56056_n144_bF_buf0), .B(rf_dout_3_), .Y(u6__abc_56056_n163_1) );
  OR2X2 OR2X2_5125 ( .A(u6__abc_56056_n154_bF_buf1), .B(mem_dout_3_), .Y(u6__abc_56056_n164) );
  OR2X2 OR2X2_5126 ( .A(u6__abc_56056_n144_bF_buf5), .B(rf_dout_4_), .Y(u6__abc_56056_n166_1) );
  OR2X2 OR2X2_5127 ( .A(u6__abc_56056_n154_bF_buf0), .B(mem_dout_4_), .Y(u6__abc_56056_n167_1) );
  OR2X2 OR2X2_5128 ( .A(u6__abc_56056_n144_bF_buf4), .B(rf_dout_5_), .Y(u6__abc_56056_n169) );
  OR2X2 OR2X2_5129 ( .A(u6__abc_56056_n154_bF_buf4), .B(mem_dout_5_), .Y(u6__abc_56056_n170) );
  OR2X2 OR2X2_513 ( .A(u0__abc_49347_n2763), .B(u0__abc_49347_n2764), .Y(u0__abc_49347_n2765) );
  OR2X2 OR2X2_5130 ( .A(u6__abc_56056_n144_bF_buf3), .B(rf_dout_6_), .Y(u6__abc_56056_n172) );
  OR2X2 OR2X2_5131 ( .A(u6__abc_56056_n154_bF_buf3), .B(mem_dout_6_), .Y(u6__abc_56056_n173) );
  OR2X2 OR2X2_5132 ( .A(u6__abc_56056_n144_bF_buf2), .B(rf_dout_7_), .Y(u6__abc_56056_n175) );
  OR2X2 OR2X2_5133 ( .A(u6__abc_56056_n154_bF_buf2), .B(mem_dout_7_), .Y(u6__abc_56056_n176) );
  OR2X2 OR2X2_5134 ( .A(u6__abc_56056_n144_bF_buf1), .B(rf_dout_8_), .Y(u6__abc_56056_n178) );
  OR2X2 OR2X2_5135 ( .A(u6__abc_56056_n154_bF_buf1), .B(mem_dout_8_), .Y(u6__abc_56056_n179) );
  OR2X2 OR2X2_5136 ( .A(u6__abc_56056_n144_bF_buf0), .B(rf_dout_9_), .Y(u6__abc_56056_n181) );
  OR2X2 OR2X2_5137 ( .A(u6__abc_56056_n154_bF_buf0), .B(mem_dout_9_), .Y(u6__abc_56056_n182) );
  OR2X2 OR2X2_5138 ( .A(u6__abc_56056_n144_bF_buf5), .B(rf_dout_10_), .Y(u6__abc_56056_n184) );
  OR2X2 OR2X2_5139 ( .A(u6__abc_56056_n154_bF_buf4), .B(mem_dout_10_), .Y(u6__abc_56056_n185) );
  OR2X2 OR2X2_514 ( .A(u0__abc_49347_n2766), .B(u0__abc_49347_n2767), .Y(u0__abc_49347_n2768) );
  OR2X2 OR2X2_5140 ( .A(u6__abc_56056_n144_bF_buf4), .B(rf_dout_11_), .Y(u6__abc_56056_n187) );
  OR2X2 OR2X2_5141 ( .A(u6__abc_56056_n154_bF_buf3), .B(mem_dout_11_), .Y(u6__abc_56056_n188) );
  OR2X2 OR2X2_5142 ( .A(u6__abc_56056_n144_bF_buf3), .B(rf_dout_12_), .Y(u6__abc_56056_n190) );
  OR2X2 OR2X2_5143 ( .A(u6__abc_56056_n154_bF_buf2), .B(mem_dout_12_), .Y(u6__abc_56056_n191) );
  OR2X2 OR2X2_5144 ( .A(u6__abc_56056_n144_bF_buf2), .B(rf_dout_13_), .Y(u6__abc_56056_n193) );
  OR2X2 OR2X2_5145 ( .A(u6__abc_56056_n154_bF_buf1), .B(mem_dout_13_), .Y(u6__abc_56056_n194) );
  OR2X2 OR2X2_5146 ( .A(u6__abc_56056_n144_bF_buf1), .B(rf_dout_14_), .Y(u6__abc_56056_n196) );
  OR2X2 OR2X2_5147 ( .A(u6__abc_56056_n154_bF_buf0), .B(mem_dout_14_), .Y(u6__abc_56056_n197) );
  OR2X2 OR2X2_5148 ( .A(u6__abc_56056_n144_bF_buf0), .B(rf_dout_15_), .Y(u6__abc_56056_n199) );
  OR2X2 OR2X2_5149 ( .A(u6__abc_56056_n154_bF_buf4), .B(mem_dout_15_), .Y(u6__abc_56056_n200) );
  OR2X2 OR2X2_515 ( .A(u0__abc_49347_n2770), .B(u0_cs0_bF_buf3), .Y(u0__abc_49347_n2771) );
  OR2X2 OR2X2_5150 ( .A(u6__abc_56056_n144_bF_buf5), .B(rf_dout_16_), .Y(u6__abc_56056_n202) );
  OR2X2 OR2X2_5151 ( .A(u6__abc_56056_n154_bF_buf3), .B(mem_dout_16_), .Y(u6__abc_56056_n203) );
  OR2X2 OR2X2_5152 ( .A(u6__abc_56056_n144_bF_buf4), .B(rf_dout_17_), .Y(u6__abc_56056_n205) );
  OR2X2 OR2X2_5153 ( .A(u6__abc_56056_n154_bF_buf2), .B(mem_dout_17_), .Y(u6__abc_56056_n206) );
  OR2X2 OR2X2_5154 ( .A(u6__abc_56056_n144_bF_buf3), .B(rf_dout_18_), .Y(u6__abc_56056_n208) );
  OR2X2 OR2X2_5155 ( .A(u6__abc_56056_n154_bF_buf1), .B(mem_dout_18_), .Y(u6__abc_56056_n209) );
  OR2X2 OR2X2_5156 ( .A(u6__abc_56056_n144_bF_buf2), .B(rf_dout_19_), .Y(u6__abc_56056_n211) );
  OR2X2 OR2X2_5157 ( .A(u6__abc_56056_n154_bF_buf0), .B(mem_dout_19_), .Y(u6__abc_56056_n212) );
  OR2X2 OR2X2_5158 ( .A(u6__abc_56056_n144_bF_buf1), .B(rf_dout_20_), .Y(u6__abc_56056_n214) );
  OR2X2 OR2X2_5159 ( .A(u6__abc_56056_n154_bF_buf4), .B(mem_dout_20_), .Y(u6__abc_56056_n215) );
  OR2X2 OR2X2_516 ( .A(u0__abc_49347_n2769), .B(u0__abc_49347_n2771), .Y(u0__abc_49347_n2772) );
  OR2X2 OR2X2_5160 ( .A(u6__abc_56056_n144_bF_buf0), .B(rf_dout_21_), .Y(u6__abc_56056_n217) );
  OR2X2 OR2X2_5161 ( .A(u6__abc_56056_n154_bF_buf3), .B(mem_dout_21_), .Y(u6__abc_56056_n218) );
  OR2X2 OR2X2_5162 ( .A(u6__abc_56056_n144_bF_buf5), .B(rf_dout_22_), .Y(u6__abc_56056_n220) );
  OR2X2 OR2X2_5163 ( .A(u6__abc_56056_n154_bF_buf2), .B(mem_dout_22_), .Y(u6__abc_56056_n221) );
  OR2X2 OR2X2_5164 ( .A(u6__abc_56056_n144_bF_buf4), .B(rf_dout_23_), .Y(u6__abc_56056_n223) );
  OR2X2 OR2X2_5165 ( .A(u6__abc_56056_n154_bF_buf1), .B(mem_dout_23_), .Y(u6__abc_56056_n224) );
  OR2X2 OR2X2_5166 ( .A(u6__abc_56056_n144_bF_buf3), .B(rf_dout_24_), .Y(u6__abc_56056_n226) );
  OR2X2 OR2X2_5167 ( .A(u6__abc_56056_n154_bF_buf0), .B(mem_dout_24_), .Y(u6__abc_56056_n227) );
  OR2X2 OR2X2_5168 ( .A(u6__abc_56056_n144_bF_buf2), .B(rf_dout_25_), .Y(u6__abc_56056_n229) );
  OR2X2 OR2X2_5169 ( .A(u6__abc_56056_n154_bF_buf4), .B(mem_dout_25_), .Y(u6__abc_56056_n230) );
  OR2X2 OR2X2_517 ( .A(u0__abc_49347_n2748_bF_buf4), .B(u0_tms0_1_), .Y(u0__abc_49347_n2773) );
  OR2X2 OR2X2_5170 ( .A(u6__abc_56056_n144_bF_buf1), .B(rf_dout_26_), .Y(u6__abc_56056_n232) );
  OR2X2 OR2X2_5171 ( .A(u6__abc_56056_n154_bF_buf3), .B(mem_dout_26_), .Y(u6__abc_56056_n233) );
  OR2X2 OR2X2_5172 ( .A(u6__abc_56056_n144_bF_buf0), .B(rf_dout_27_), .Y(u6__abc_56056_n235) );
  OR2X2 OR2X2_5173 ( .A(u6__abc_56056_n154_bF_buf2), .B(mem_dout_27_), .Y(u6__abc_56056_n236) );
  OR2X2 OR2X2_5174 ( .A(u6__abc_56056_n144_bF_buf5), .B(rf_dout_28_), .Y(u6__abc_56056_n238) );
  OR2X2 OR2X2_5175 ( .A(u6__abc_56056_n154_bF_buf1), .B(mem_dout_28_), .Y(u6__abc_56056_n239) );
  OR2X2 OR2X2_5176 ( .A(u6__abc_56056_n144_bF_buf4), .B(rf_dout_29_), .Y(u6__abc_56056_n241) );
  OR2X2 OR2X2_5177 ( .A(u6__abc_56056_n154_bF_buf0), .B(mem_dout_29_), .Y(u6__abc_56056_n242) );
  OR2X2 OR2X2_5178 ( .A(u6__abc_56056_n144_bF_buf3), .B(rf_dout_30_), .Y(u6__abc_56056_n244) );
  OR2X2 OR2X2_5179 ( .A(u6__abc_56056_n154_bF_buf4), .B(mem_dout_30_), .Y(u6__abc_56056_n245) );
  OR2X2 OR2X2_518 ( .A(u0__abc_49347_n2775), .B(u0__abc_49347_n2753), .Y(u0_tms_1__FF_INPUT) );
  OR2X2 OR2X2_5180 ( .A(u6__abc_56056_n144_bF_buf2), .B(rf_dout_31_), .Y(u6__abc_56056_n247) );
  OR2X2 OR2X2_5181 ( .A(u6__abc_56056_n154_bF_buf3), .B(mem_dout_31_), .Y(u6__abc_56056_n248) );
  OR2X2 OR2X2_5182 ( .A(u6__abc_56056_n251), .B(u6__abc_56056_n250), .Y(u6_wr_hold_FF_INPUT) );
  OR2X2 OR2X2_5183 ( .A(u6__abc_56056_n258), .B(u6_read_go_r), .Y(u6__abc_56056_n259) );
  OR2X2 OR2X2_5184 ( .A(u6__abc_56056_n267), .B(u6_write_go_r), .Y(u6__abc_56056_n268) );
  OR2X2 OR2X2_5185 ( .A(u6__abc_56056_n270), .B(wb_we_i), .Y(u6__abc_56056_n271) );
  OR2X2 OR2X2_5186 ( .A(u6__abc_56056_n279), .B(u6__abc_56056_n282), .Y(u5_wb_first) );
  OR2X2 OR2X2_5187 ( .A(u3_wb_read_go), .B(u1_wb_write_go), .Y(u6__abc_56056_n287) );
  OR2X2 OR2X2_5188 ( .A(u6__abc_56056_n290), .B(_auto_iopadmap_cc_313_execute_56356), .Y(u6_rmw_en_FF_INPUT) );
  OR2X2 OR2X2_5189 ( .A(u7__abc_47535_n78), .B(u1_wr_cycle), .Y(u7__abc_47535_n79_1) );
  OR2X2 OR2X2_519 ( .A(u0__abc_49347_n2728_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n2779) );
  OR2X2 OR2X2_5190 ( .A(u7__abc_47535_n80_1), .B(susp_sel), .Y(u7__abc_47535_n81_1) );
  OR2X2 OR2X2_5191 ( .A(u7__abc_47535_n81_1), .B(u7__abc_47535_n76), .Y(u7_mc_dqm_0__FF_INPUT) );
  OR2X2 OR2X2_5192 ( .A(u7__abc_47535_n81_1), .B(u7__abc_47535_n84), .Y(u7_mc_dqm_1__FF_INPUT) );
  OR2X2 OR2X2_5193 ( .A(u7__abc_47535_n81_1), .B(u7__abc_47535_n87_1), .Y(u7_mc_dqm_2__FF_INPUT) );
  OR2X2 OR2X2_5194 ( .A(u7__abc_47535_n81_1), .B(u7__abc_47535_n90_1), .Y(u7_mc_dqm_3__FF_INPUT) );
  OR2X2 OR2X2_5195 ( .A(u7__abc_47535_n95_1), .B(u7__abc_47535_n93), .Y(u7_mc_dqm_r_0__FF_INPUT) );
  OR2X2 OR2X2_5196 ( .A(u7__abc_47535_n98_1), .B(u7__abc_47535_n97_1), .Y(u7_mc_dqm_r_1__FF_INPUT) );
  OR2X2 OR2X2_5197 ( .A(u7__abc_47535_n101), .B(u7__abc_47535_n100), .Y(u7_mc_dqm_r_2__FF_INPUT) );
  OR2X2 OR2X2_5198 ( .A(u7__abc_47535_n104), .B(u7__abc_47535_n103), .Y(u7_mc_dqm_r_3__FF_INPUT) );
  OR2X2 OR2X2_5199 ( .A(susp_sel), .B(rfr_ack), .Y(u7__abc_47535_n106) );
  OR2X2 OR2X2_52 ( .A(lmr_sel_bF_buf4), .B(tms_8_), .Y(_abc_55805_n315) );
  OR2X2 OR2X2_520 ( .A(1'b0), .B(1'b0), .Y(u0__abc_49347_n2780) );
  OR2X2 OR2X2_5200 ( .A(u7__abc_47535_n108), .B(lmr_sel_bF_buf2), .Y(u7__abc_47535_n109) );
  OR2X2 OR2X2_5201 ( .A(u7__abc_47535_n116), .B(u7__abc_47535_n114), .Y(u7__abc_47535_n117) );
  OR2X2 OR2X2_5202 ( .A(u7__abc_47535_n113), .B(u7__abc_47535_n117), .Y(u7_mc_cs__FF_INPUT) );
  OR2X2 OR2X2_5203 ( .A(u7__abc_47535_n119), .B(lmr_sel_bF_buf0), .Y(u7__abc_47535_n120) );
  OR2X2 OR2X2_5204 ( .A(u7__abc_47535_n126), .B(u7__abc_47535_n114), .Y(u7__abc_47535_n127) );
  OR2X2 OR2X2_5205 ( .A(u7__abc_47535_n124), .B(u7__abc_47535_n127), .Y(u7_mc_cs__FF_INPUT) );
  OR2X2 OR2X2_5206 ( .A(u7__abc_47535_n129), .B(lmr_sel_bF_buf5), .Y(u7__abc_47535_n130) );
  OR2X2 OR2X2_5207 ( .A(u7__abc_47535_n136), .B(u7__abc_47535_n114), .Y(u7__abc_47535_n137) );
  OR2X2 OR2X2_5208 ( .A(u7__abc_47535_n134), .B(u7__abc_47535_n137), .Y(u7_mc_cs__FF_INPUT) );
  OR2X2 OR2X2_5209 ( .A(u7__abc_47535_n139), .B(lmr_sel_bF_buf3), .Y(u7__abc_47535_n140) );
  OR2X2 OR2X2_521 ( .A(u0__abc_49347_n2782), .B(u0__abc_49347_n2778), .Y(u0__abc_49347_n2783) );
  OR2X2 OR2X2_5210 ( .A(u7__abc_47535_n146), .B(u7__abc_47535_n114), .Y(u7__abc_47535_n147) );
  OR2X2 OR2X2_5211 ( .A(u7__abc_47535_n144), .B(u7__abc_47535_n147), .Y(u7_mc_cs__FF_INPUT) );
  OR2X2 OR2X2_5212 ( .A(u7__abc_47535_n149), .B(lmr_sel_bF_buf1), .Y(u7__abc_47535_n150) );
  OR2X2 OR2X2_5213 ( .A(u7__abc_47535_n156), .B(u7__abc_47535_n114), .Y(u7__abc_47535_n157) );
  OR2X2 OR2X2_5214 ( .A(u7__abc_47535_n154), .B(u7__abc_47535_n157), .Y(u7_mc_cs__FF_INPUT) );
  OR2X2 OR2X2_5215 ( .A(u7__abc_47535_n159), .B(lmr_sel_bF_buf6), .Y(u7__abc_47535_n160) );
  OR2X2 OR2X2_5216 ( .A(u7__abc_47535_n166), .B(u7__abc_47535_n114), .Y(u7__abc_47535_n167) );
  OR2X2 OR2X2_5217 ( .A(u7__abc_47535_n164), .B(u7__abc_47535_n167), .Y(u7_mc_cs__FF_INPUT) );
  OR2X2 OR2X2_5218 ( .A(u7__abc_47535_n169), .B(lmr_sel_bF_buf4), .Y(u7__abc_47535_n170) );
  OR2X2 OR2X2_5219 ( .A(u7__abc_47535_n176), .B(u7__abc_47535_n114), .Y(u7__abc_47535_n177) );
  OR2X2 OR2X2_522 ( .A(u0__abc_49347_n2784_1), .B(u0__abc_49347_n2785), .Y(u0__abc_49347_n2786) );
  OR2X2 OR2X2_5220 ( .A(u7__abc_47535_n174), .B(u7__abc_47535_n177), .Y(u7_mc_cs__FF_INPUT) );
  OR2X2 OR2X2_5221 ( .A(u7__abc_47535_n179), .B(lmr_sel_bF_buf2), .Y(u7__abc_47535_n180) );
  OR2X2 OR2X2_5222 ( .A(u7__abc_47535_n186), .B(u7__abc_47535_n114), .Y(u7__abc_47535_n187) );
  OR2X2 OR2X2_5223 ( .A(u7__abc_47535_n184), .B(u7__abc_47535_n187), .Y(u7_mc_cs__FF_INPUT) );
  OR2X2 OR2X2_5224 ( .A(susp_sel), .B(oe_), .Y(u7_mc_oe__FF_INPUT) );
  OR2X2 OR2X2_523 ( .A(u0__abc_49347_n2787), .B(u0__abc_49347_n2788), .Y(u0__abc_49347_n2789) );
  OR2X2 OR2X2_524 ( .A(u0__abc_49347_n2790), .B(u0__abc_49347_n2791), .Y(u0__abc_49347_n2792) );
  OR2X2 OR2X2_525 ( .A(u0__abc_49347_n2794), .B(u0_cs0_bF_buf2), .Y(u0__abc_49347_n2795) );
  OR2X2 OR2X2_526 ( .A(u0__abc_49347_n2793), .B(u0__abc_49347_n2795), .Y(u0__abc_49347_n2796) );
  OR2X2 OR2X2_527 ( .A(u0__abc_49347_n2748_bF_buf3), .B(u0_tms0_2_), .Y(u0__abc_49347_n2797) );
  OR2X2 OR2X2_528 ( .A(u0__abc_49347_n2799), .B(u0__abc_49347_n2777), .Y(u0_tms_2__FF_INPUT) );
  OR2X2 OR2X2_529 ( .A(u0__abc_49347_n2728_bF_buf2), .B(1'b0), .Y(u0__abc_49347_n2803) );
  OR2X2 OR2X2_53 ( .A(_abc_55805_n240_bF_buf0), .B(sp_tms_9_), .Y(_abc_55805_n317) );
  OR2X2 OR2X2_530 ( .A(1'b0), .B(1'b0), .Y(u0__abc_49347_n2804) );
  OR2X2 OR2X2_531 ( .A(u0__abc_49347_n2806), .B(u0__abc_49347_n2802), .Y(u0__abc_49347_n2807) );
  OR2X2 OR2X2_532 ( .A(u0__abc_49347_n2808), .B(u0__abc_49347_n2809), .Y(u0__abc_49347_n2810) );
  OR2X2 OR2X2_533 ( .A(u0__abc_49347_n2811), .B(u0__abc_49347_n2812), .Y(u0__abc_49347_n2813) );
  OR2X2 OR2X2_534 ( .A(u0__abc_49347_n2814), .B(u0__abc_49347_n2815), .Y(u0__abc_49347_n2816_1) );
  OR2X2 OR2X2_535 ( .A(u0__abc_49347_n2818), .B(u0_cs0_bF_buf1), .Y(u0__abc_49347_n2819) );
  OR2X2 OR2X2_536 ( .A(u0__abc_49347_n2817), .B(u0__abc_49347_n2819), .Y(u0__abc_49347_n2820) );
  OR2X2 OR2X2_537 ( .A(u0__abc_49347_n2748_bF_buf2), .B(u0_tms0_3_), .Y(u0__abc_49347_n2821) );
  OR2X2 OR2X2_538 ( .A(u0__abc_49347_n2823), .B(u0__abc_49347_n2801), .Y(u0_tms_3__FF_INPUT) );
  OR2X2 OR2X2_539 ( .A(u0__abc_49347_n2728_bF_buf1), .B(1'b0), .Y(u0__abc_49347_n2827) );
  OR2X2 OR2X2_54 ( .A(lmr_sel_bF_buf3), .B(tms_9_), .Y(_abc_55805_n318) );
  OR2X2 OR2X2_540 ( .A(1'b0), .B(1'b0), .Y(u0__abc_49347_n2828) );
  OR2X2 OR2X2_541 ( .A(u0__abc_49347_n2830), .B(u0__abc_49347_n2826), .Y(u0__abc_49347_n2831) );
  OR2X2 OR2X2_542 ( .A(u0__abc_49347_n2832), .B(u0__abc_49347_n2833), .Y(u0__abc_49347_n2834) );
  OR2X2 OR2X2_543 ( .A(u0__abc_49347_n2835), .B(u0__abc_49347_n2836), .Y(u0__abc_49347_n2837) );
  OR2X2 OR2X2_544 ( .A(u0__abc_49347_n2838), .B(u0__abc_49347_n2839), .Y(u0__abc_49347_n2840) );
  OR2X2 OR2X2_545 ( .A(u0__abc_49347_n2842), .B(u0_cs0_bF_buf0), .Y(u0__abc_49347_n2843) );
  OR2X2 OR2X2_546 ( .A(u0__abc_49347_n2841), .B(u0__abc_49347_n2843), .Y(u0__abc_49347_n2844) );
  OR2X2 OR2X2_547 ( .A(u0__abc_49347_n2748_bF_buf1), .B(u0_tms0_4_), .Y(u0__abc_49347_n2845) );
  OR2X2 OR2X2_548 ( .A(u0__abc_49347_n2847), .B(u0__abc_49347_n2825), .Y(u0_tms_4__FF_INPUT) );
  OR2X2 OR2X2_549 ( .A(u0__abc_49347_n2728_bF_buf0), .B(1'b0), .Y(u0__abc_49347_n2851) );
  OR2X2 OR2X2_55 ( .A(_abc_55805_n240_bF_buf5), .B(sp_tms_10_), .Y(_abc_55805_n320) );
  OR2X2 OR2X2_550 ( .A(1'b0), .B(1'b0), .Y(u0__abc_49347_n2852) );
  OR2X2 OR2X2_551 ( .A(u0__abc_49347_n2854), .B(u0__abc_49347_n2850), .Y(u0__abc_49347_n2855) );
  OR2X2 OR2X2_552 ( .A(u0__abc_49347_n2856), .B(u0__abc_49347_n2857), .Y(u0__abc_49347_n2858) );
  OR2X2 OR2X2_553 ( .A(u0__abc_49347_n2859), .B(u0__abc_49347_n2860), .Y(u0__abc_49347_n2861) );
  OR2X2 OR2X2_554 ( .A(u0__abc_49347_n2862), .B(u0__abc_49347_n2863), .Y(u0__abc_49347_n2864) );
  OR2X2 OR2X2_555 ( .A(u0__abc_49347_n2866), .B(u0_cs0_bF_buf5), .Y(u0__abc_49347_n2867) );
  OR2X2 OR2X2_556 ( .A(u0__abc_49347_n2865), .B(u0__abc_49347_n2867), .Y(u0__abc_49347_n2868) );
  OR2X2 OR2X2_557 ( .A(u0__abc_49347_n2748_bF_buf0), .B(u0_tms0_5_), .Y(u0__abc_49347_n2869) );
  OR2X2 OR2X2_558 ( .A(u0__abc_49347_n2871), .B(u0__abc_49347_n2849), .Y(u0_tms_5__FF_INPUT) );
  OR2X2 OR2X2_559 ( .A(u0__abc_49347_n2728_bF_buf5), .B(1'b0), .Y(u0__abc_49347_n2875) );
  OR2X2 OR2X2_56 ( .A(lmr_sel_bF_buf2), .B(tms_10_), .Y(_abc_55805_n321) );
  OR2X2 OR2X2_560 ( .A(1'b0), .B(1'b0), .Y(u0__abc_49347_n2876) );
  OR2X2 OR2X2_561 ( .A(u0__abc_49347_n2878), .B(u0__abc_49347_n2874), .Y(u0__abc_49347_n2879) );
  OR2X2 OR2X2_562 ( .A(u0__abc_49347_n2880), .B(u0__abc_49347_n2881_1), .Y(u0__abc_49347_n2882) );
  OR2X2 OR2X2_563 ( .A(u0__abc_49347_n2883), .B(u0__abc_49347_n2884), .Y(u0__abc_49347_n2885) );
  OR2X2 OR2X2_564 ( .A(u0__abc_49347_n2886), .B(u0__abc_49347_n2887), .Y(u0__abc_49347_n2888) );
  OR2X2 OR2X2_565 ( .A(u0__abc_49347_n2890), .B(u0_cs0_bF_buf4), .Y(u0__abc_49347_n2891) );
  OR2X2 OR2X2_566 ( .A(u0__abc_49347_n2889), .B(u0__abc_49347_n2891), .Y(u0__abc_49347_n2892) );
  OR2X2 OR2X2_567 ( .A(u0__abc_49347_n2748_bF_buf5), .B(u0_tms0_6_), .Y(u0__abc_49347_n2893) );
  OR2X2 OR2X2_568 ( .A(u0__abc_49347_n2895), .B(u0__abc_49347_n2873), .Y(u0_tms_6__FF_INPUT) );
  OR2X2 OR2X2_569 ( .A(u0__abc_49347_n2728_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n2899) );
  OR2X2 OR2X2_57 ( .A(_abc_55805_n240_bF_buf4), .B(sp_tms_11_), .Y(_abc_55805_n323) );
  OR2X2 OR2X2_570 ( .A(1'b0), .B(1'b0), .Y(u0__abc_49347_n2900) );
  OR2X2 OR2X2_571 ( .A(u0__abc_49347_n2902), .B(u0__abc_49347_n2898), .Y(u0__abc_49347_n2903) );
  OR2X2 OR2X2_572 ( .A(u0__abc_49347_n2904), .B(u0__abc_49347_n2905), .Y(u0__abc_49347_n2906) );
  OR2X2 OR2X2_573 ( .A(u0__abc_49347_n2907), .B(u0__abc_49347_n2908), .Y(u0__abc_49347_n2909) );
  OR2X2 OR2X2_574 ( .A(u0__abc_49347_n2910), .B(u0__abc_49347_n2911), .Y(u0__abc_49347_n2912) );
  OR2X2 OR2X2_575 ( .A(u0__abc_49347_n2914), .B(u0_cs0_bF_buf3), .Y(u0__abc_49347_n2915) );
  OR2X2 OR2X2_576 ( .A(u0__abc_49347_n2913_1), .B(u0__abc_49347_n2915), .Y(u0__abc_49347_n2916) );
  OR2X2 OR2X2_577 ( .A(u0__abc_49347_n2748_bF_buf4), .B(u0_tms0_7_), .Y(u0__abc_49347_n2917) );
  OR2X2 OR2X2_578 ( .A(u0__abc_49347_n2919), .B(u0__abc_49347_n2897), .Y(u0_tms_7__FF_INPUT) );
  OR2X2 OR2X2_579 ( .A(u0__abc_49347_n2728_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n2923) );
  OR2X2 OR2X2_58 ( .A(lmr_sel_bF_buf1), .B(tms_11_), .Y(_abc_55805_n324) );
  OR2X2 OR2X2_580 ( .A(1'b0), .B(1'b0), .Y(u0__abc_49347_n2924) );
  OR2X2 OR2X2_581 ( .A(u0__abc_49347_n2926), .B(u0__abc_49347_n2922), .Y(u0__abc_49347_n2927) );
  OR2X2 OR2X2_582 ( .A(u0__abc_49347_n2928), .B(u0__abc_49347_n2929), .Y(u0__abc_49347_n2930) );
  OR2X2 OR2X2_583 ( .A(u0__abc_49347_n2931), .B(u0__abc_49347_n2932), .Y(u0__abc_49347_n2933) );
  OR2X2 OR2X2_584 ( .A(u0__abc_49347_n2934), .B(u0__abc_49347_n2935), .Y(u0__abc_49347_n2936) );
  OR2X2 OR2X2_585 ( .A(u0__abc_49347_n2938), .B(u0_cs0_bF_buf2), .Y(u0__abc_49347_n2939) );
  OR2X2 OR2X2_586 ( .A(u0__abc_49347_n2937), .B(u0__abc_49347_n2939), .Y(u0__abc_49347_n2940) );
  OR2X2 OR2X2_587 ( .A(u0__abc_49347_n2748_bF_buf3), .B(u0_tms0_8_), .Y(u0__abc_49347_n2941) );
  OR2X2 OR2X2_588 ( .A(u0__abc_49347_n2943), .B(u0__abc_49347_n2921), .Y(u0_tms_8__FF_INPUT) );
  OR2X2 OR2X2_589 ( .A(u0__abc_49347_n2728_bF_buf2), .B(1'b0), .Y(u0__abc_49347_n2947) );
  OR2X2 OR2X2_59 ( .A(_abc_55805_n240_bF_buf3), .B(sp_tms_12_), .Y(_abc_55805_n326) );
  OR2X2 OR2X2_590 ( .A(1'b0), .B(1'b0), .Y(u0__abc_49347_n2948) );
  OR2X2 OR2X2_591 ( .A(u0__abc_49347_n2950), .B(u0__abc_49347_n2946), .Y(u0__abc_49347_n2951) );
  OR2X2 OR2X2_592 ( .A(u0__abc_49347_n2952), .B(u0__abc_49347_n2953), .Y(u0__abc_49347_n2954) );
  OR2X2 OR2X2_593 ( .A(u0__abc_49347_n2955), .B(u0__abc_49347_n2956), .Y(u0__abc_49347_n2957) );
  OR2X2 OR2X2_594 ( .A(u0__abc_49347_n2958), .B(u0__abc_49347_n2959), .Y(u0__abc_49347_n2960) );
  OR2X2 OR2X2_595 ( .A(u0__abc_49347_n2962), .B(u0_cs0_bF_buf1), .Y(u0__abc_49347_n2963) );
  OR2X2 OR2X2_596 ( .A(u0__abc_49347_n2961), .B(u0__abc_49347_n2963), .Y(u0__abc_49347_n2964) );
  OR2X2 OR2X2_597 ( .A(u0__abc_49347_n2748_bF_buf2), .B(u0_tms0_9_), .Y(u0__abc_49347_n2965) );
  OR2X2 OR2X2_598 ( .A(u0__abc_49347_n2967), .B(u0__abc_49347_n2945_1), .Y(u0_tms_9__FF_INPUT) );
  OR2X2 OR2X2_599 ( .A(u0__abc_49347_n2728_bF_buf1), .B(1'b0), .Y(u0__abc_49347_n2971) );
  OR2X2 OR2X2_6 ( .A(_abc_55805_n245_1), .B(cs_need_rfr_0_), .Y(_abc_55805_n246) );
  OR2X2 OR2X2_60 ( .A(lmr_sel_bF_buf0), .B(tms_12_), .Y(_abc_55805_n327) );
  OR2X2 OR2X2_600 ( .A(1'b0), .B(1'b0), .Y(u0__abc_49347_n2972) );
  OR2X2 OR2X2_601 ( .A(u0__abc_49347_n2974), .B(u0__abc_49347_n2970), .Y(u0__abc_49347_n2975) );
  OR2X2 OR2X2_602 ( .A(u0__abc_49347_n2976), .B(u0__abc_49347_n2977_1), .Y(u0__abc_49347_n2978) );
  OR2X2 OR2X2_603 ( .A(u0__abc_49347_n2979), .B(u0__abc_49347_n2980), .Y(u0__abc_49347_n2981) );
  OR2X2 OR2X2_604 ( .A(u0__abc_49347_n2982), .B(u0__abc_49347_n2983), .Y(u0__abc_49347_n2984) );
  OR2X2 OR2X2_605 ( .A(u0__abc_49347_n2986), .B(u0_cs0_bF_buf0), .Y(u0__abc_49347_n2987) );
  OR2X2 OR2X2_606 ( .A(u0__abc_49347_n2985), .B(u0__abc_49347_n2987), .Y(u0__abc_49347_n2988) );
  OR2X2 OR2X2_607 ( .A(u0__abc_49347_n2748_bF_buf1), .B(u0_tms0_10_), .Y(u0__abc_49347_n2989) );
  OR2X2 OR2X2_608 ( .A(u0__abc_49347_n2991), .B(u0__abc_49347_n2969), .Y(u0_tms_10__FF_INPUT) );
  OR2X2 OR2X2_609 ( .A(u0__abc_49347_n2728_bF_buf0), .B(1'b0), .Y(u0__abc_49347_n2995) );
  OR2X2 OR2X2_61 ( .A(_abc_55805_n240_bF_buf2), .B(sp_tms_13_), .Y(_abc_55805_n329) );
  OR2X2 OR2X2_610 ( .A(1'b0), .B(1'b0), .Y(u0__abc_49347_n2996) );
  OR2X2 OR2X2_611 ( .A(u0__abc_49347_n2998), .B(u0__abc_49347_n2994), .Y(u0__abc_49347_n2999) );
  OR2X2 OR2X2_612 ( .A(u0__abc_49347_n3000), .B(u0__abc_49347_n3001), .Y(u0__abc_49347_n3002) );
  OR2X2 OR2X2_613 ( .A(u0__abc_49347_n3003), .B(u0__abc_49347_n3004), .Y(u0__abc_49347_n3005) );
  OR2X2 OR2X2_614 ( .A(u0__abc_49347_n3006), .B(u0__abc_49347_n3007), .Y(u0__abc_49347_n3008) );
  OR2X2 OR2X2_615 ( .A(u0__abc_49347_n3010), .B(u0_cs0_bF_buf5), .Y(u0__abc_49347_n3011) );
  OR2X2 OR2X2_616 ( .A(u0__abc_49347_n3009_1), .B(u0__abc_49347_n3011), .Y(u0__abc_49347_n3012) );
  OR2X2 OR2X2_617 ( .A(u0__abc_49347_n2748_bF_buf0), .B(u0_tms0_11_), .Y(u0__abc_49347_n3013) );
  OR2X2 OR2X2_618 ( .A(u0__abc_49347_n3015), .B(u0__abc_49347_n2993), .Y(u0_tms_11__FF_INPUT) );
  OR2X2 OR2X2_619 ( .A(u0__abc_49347_n2728_bF_buf5), .B(1'b0), .Y(u0__abc_49347_n3019) );
  OR2X2 OR2X2_62 ( .A(lmr_sel_bF_buf6), .B(tms_13_), .Y(_abc_55805_n330) );
  OR2X2 OR2X2_620 ( .A(1'b0), .B(1'b0), .Y(u0__abc_49347_n3020) );
  OR2X2 OR2X2_621 ( .A(u0__abc_49347_n3022), .B(u0__abc_49347_n3018), .Y(u0__abc_49347_n3023) );
  OR2X2 OR2X2_622 ( .A(u0__abc_49347_n3024), .B(u0__abc_49347_n3025), .Y(u0__abc_49347_n3026) );
  OR2X2 OR2X2_623 ( .A(u0__abc_49347_n3027), .B(u0__abc_49347_n3028), .Y(u0__abc_49347_n3029) );
  OR2X2 OR2X2_624 ( .A(u0__abc_49347_n3030), .B(u0__abc_49347_n3031), .Y(u0__abc_49347_n3032) );
  OR2X2 OR2X2_625 ( .A(u0__abc_49347_n3034), .B(u0_cs0_bF_buf4), .Y(u0__abc_49347_n3035) );
  OR2X2 OR2X2_626 ( .A(u0__abc_49347_n3033), .B(u0__abc_49347_n3035), .Y(u0__abc_49347_n3036) );
  OR2X2 OR2X2_627 ( .A(u0__abc_49347_n2748_bF_buf5), .B(u0_tms0_12_), .Y(u0__abc_49347_n3037) );
  OR2X2 OR2X2_628 ( .A(u0__abc_49347_n3039), .B(u0__abc_49347_n3017), .Y(u0_tms_12__FF_INPUT) );
  OR2X2 OR2X2_629 ( .A(u0__abc_49347_n2728_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n3043) );
  OR2X2 OR2X2_63 ( .A(_abc_55805_n240_bF_buf1), .B(sp_tms_14_), .Y(_abc_55805_n332) );
  OR2X2 OR2X2_630 ( .A(1'b0), .B(1'b0), .Y(u0__abc_49347_n3044) );
  OR2X2 OR2X2_631 ( .A(u0__abc_49347_n3046), .B(u0__abc_49347_n3042), .Y(u0__abc_49347_n3047) );
  OR2X2 OR2X2_632 ( .A(u0__abc_49347_n3048), .B(u0__abc_49347_n3049), .Y(u0__abc_49347_n3050) );
  OR2X2 OR2X2_633 ( .A(u0__abc_49347_n3051), .B(u0__abc_49347_n3052), .Y(u0__abc_49347_n3053) );
  OR2X2 OR2X2_634 ( .A(u0__abc_49347_n3054), .B(u0__abc_49347_n3055), .Y(u0__abc_49347_n3056) );
  OR2X2 OR2X2_635 ( .A(u0__abc_49347_n3058), .B(u0_cs0_bF_buf3), .Y(u0__abc_49347_n3059) );
  OR2X2 OR2X2_636 ( .A(u0__abc_49347_n3057), .B(u0__abc_49347_n3059), .Y(u0__abc_49347_n3060) );
  OR2X2 OR2X2_637 ( .A(u0__abc_49347_n2748_bF_buf4), .B(u0_tms0_13_), .Y(u0__abc_49347_n3061) );
  OR2X2 OR2X2_638 ( .A(u0__abc_49347_n3063), .B(u0__abc_49347_n3041_1), .Y(u0_tms_13__FF_INPUT) );
  OR2X2 OR2X2_639 ( .A(u0__abc_49347_n2728_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n3067) );
  OR2X2 OR2X2_64 ( .A(lmr_sel_bF_buf5), .B(tms_14_), .Y(_abc_55805_n333) );
  OR2X2 OR2X2_640 ( .A(1'b0), .B(1'b0), .Y(u0__abc_49347_n3068) );
  OR2X2 OR2X2_641 ( .A(u0__abc_49347_n3070), .B(u0__abc_49347_n3066), .Y(u0__abc_49347_n3071) );
  OR2X2 OR2X2_642 ( .A(u0__abc_49347_n3072), .B(u0__abc_49347_n3073_1), .Y(u0__abc_49347_n3074) );
  OR2X2 OR2X2_643 ( .A(u0__abc_49347_n3075), .B(u0__abc_49347_n3076), .Y(u0__abc_49347_n3077) );
  OR2X2 OR2X2_644 ( .A(u0__abc_49347_n3078), .B(u0__abc_49347_n3079), .Y(u0__abc_49347_n3080) );
  OR2X2 OR2X2_645 ( .A(u0__abc_49347_n3082), .B(u0_cs0_bF_buf2), .Y(u0__abc_49347_n3083) );
  OR2X2 OR2X2_646 ( .A(u0__abc_49347_n3081), .B(u0__abc_49347_n3083), .Y(u0__abc_49347_n3084) );
  OR2X2 OR2X2_647 ( .A(u0__abc_49347_n2748_bF_buf3), .B(u0_tms0_14_), .Y(u0__abc_49347_n3085) );
  OR2X2 OR2X2_648 ( .A(u0__abc_49347_n3087), .B(u0__abc_49347_n3065), .Y(u0_tms_14__FF_INPUT) );
  OR2X2 OR2X2_649 ( .A(u0__abc_49347_n2728_bF_buf2), .B(1'b0), .Y(u0__abc_49347_n3091) );
  OR2X2 OR2X2_65 ( .A(_abc_55805_n240_bF_buf0), .B(sp_tms_15_), .Y(_abc_55805_n335) );
  OR2X2 OR2X2_650 ( .A(1'b0), .B(1'b0), .Y(u0__abc_49347_n3092) );
  OR2X2 OR2X2_651 ( .A(u0__abc_49347_n3094), .B(u0__abc_49347_n3090), .Y(u0__abc_49347_n3095) );
  OR2X2 OR2X2_652 ( .A(u0__abc_49347_n3096), .B(u0__abc_49347_n3097), .Y(u0__abc_49347_n3098) );
  OR2X2 OR2X2_653 ( .A(u0__abc_49347_n3099), .B(u0__abc_49347_n3100), .Y(u0__abc_49347_n3101) );
  OR2X2 OR2X2_654 ( .A(u0__abc_49347_n3102), .B(u0__abc_49347_n3103), .Y(u0__abc_49347_n3104) );
  OR2X2 OR2X2_655 ( .A(u0__abc_49347_n3106_1), .B(u0_cs0_bF_buf1), .Y(u0__abc_49347_n3107) );
  OR2X2 OR2X2_656 ( .A(u0__abc_49347_n3105_1), .B(u0__abc_49347_n3107), .Y(u0__abc_49347_n3108_1) );
  OR2X2 OR2X2_657 ( .A(u0__abc_49347_n2748_bF_buf2), .B(u0_tms0_15_), .Y(u0__abc_49347_n3109) );
  OR2X2 OR2X2_658 ( .A(u0__abc_49347_n3111), .B(u0__abc_49347_n3089), .Y(u0_tms_15__FF_INPUT) );
  OR2X2 OR2X2_659 ( .A(u0__abc_49347_n2728_bF_buf1), .B(1'b0), .Y(u0__abc_49347_n3115_1) );
  OR2X2 OR2X2_66 ( .A(lmr_sel_bF_buf4), .B(tms_15_), .Y(_abc_55805_n336) );
  OR2X2 OR2X2_660 ( .A(1'b0), .B(1'b0), .Y(u0__abc_49347_n3116_1) );
  OR2X2 OR2X2_661 ( .A(u0__abc_49347_n3118), .B(u0__abc_49347_n3114), .Y(u0__abc_49347_n3119) );
  OR2X2 OR2X2_662 ( .A(u0__abc_49347_n3120_1), .B(u0__abc_49347_n3121), .Y(u0__abc_49347_n3122) );
  OR2X2 OR2X2_663 ( .A(u0__abc_49347_n3123_1), .B(u0__abc_49347_n3124), .Y(u0__abc_49347_n3125) );
  OR2X2 OR2X2_664 ( .A(u0__abc_49347_n3126_1), .B(u0__abc_49347_n3127), .Y(u0__abc_49347_n3128) );
  OR2X2 OR2X2_665 ( .A(u0__abc_49347_n3130), .B(u0_cs0_bF_buf0), .Y(u0__abc_49347_n3131) );
  OR2X2 OR2X2_666 ( .A(u0__abc_49347_n3129_1), .B(u0__abc_49347_n3131), .Y(u0__abc_49347_n3132_1) );
  OR2X2 OR2X2_667 ( .A(u0__abc_49347_n2748_bF_buf1), .B(u0_tms0_16_), .Y(u0__abc_49347_n3133) );
  OR2X2 OR2X2_668 ( .A(u0__abc_49347_n3135_1), .B(u0__abc_49347_n3113), .Y(u0_tms_16__FF_INPUT) );
  OR2X2 OR2X2_669 ( .A(u0__abc_49347_n2728_bF_buf0), .B(1'b0), .Y(u0__abc_49347_n3139) );
  OR2X2 OR2X2_67 ( .A(_abc_55805_n240_bF_buf5), .B(sp_tms_16_), .Y(_abc_55805_n338) );
  OR2X2 OR2X2_670 ( .A(1'b0), .B(1'b0), .Y(u0__abc_49347_n3140) );
  OR2X2 OR2X2_671 ( .A(u0__abc_49347_n3142), .B(u0__abc_49347_n3138_1), .Y(u0__abc_49347_n3143) );
  OR2X2 OR2X2_672 ( .A(u0__abc_49347_n3144_1), .B(u0__abc_49347_n3145_1), .Y(u0__abc_49347_n3146) );
  OR2X2 OR2X2_673 ( .A(u0__abc_49347_n3147_1), .B(u0__abc_49347_n3148), .Y(u0__abc_49347_n3149_1) );
  OR2X2 OR2X2_674 ( .A(u0__abc_49347_n3150), .B(u0__abc_49347_n3151_1), .Y(u0__abc_49347_n3152) );
  OR2X2 OR2X2_675 ( .A(u0__abc_49347_n3154), .B(u0_cs0_bF_buf5), .Y(u0__abc_49347_n3155) );
  OR2X2 OR2X2_676 ( .A(u0__abc_49347_n3153_1), .B(u0__abc_49347_n3155), .Y(u0__abc_49347_n3156_1) );
  OR2X2 OR2X2_677 ( .A(u0__abc_49347_n2748_bF_buf0), .B(u0_tms0_17_), .Y(u0__abc_49347_n3157) );
  OR2X2 OR2X2_678 ( .A(u0__abc_49347_n3159), .B(u0__abc_49347_n3137), .Y(u0_tms_17__FF_INPUT) );
  OR2X2 OR2X2_679 ( .A(u0__abc_49347_n2728_bF_buf5), .B(1'b0), .Y(u0__abc_49347_n3163_1) );
  OR2X2 OR2X2_68 ( .A(lmr_sel_bF_buf3), .B(tms_16_), .Y(_abc_55805_n339) );
  OR2X2 OR2X2_680 ( .A(1'b0), .B(1'b0), .Y(u0__abc_49347_n3164) );
  OR2X2 OR2X2_681 ( .A(u0__abc_49347_n3166), .B(u0__abc_49347_n3162), .Y(u0__abc_49347_n3167) );
  OR2X2 OR2X2_682 ( .A(u0__abc_49347_n3168), .B(u0__abc_49347_n3169), .Y(u0__abc_49347_n3170_1) );
  OR2X2 OR2X2_683 ( .A(u0__abc_49347_n3171_1), .B(u0__abc_49347_n3172_1), .Y(u0__abc_49347_n3173_1) );
  OR2X2 OR2X2_684 ( .A(u0__abc_49347_n3174_1), .B(u0__abc_49347_n3175_1), .Y(u0__abc_49347_n3176_1) );
  OR2X2 OR2X2_685 ( .A(u0__abc_49347_n3178_1), .B(u0_cs0_bF_buf4), .Y(u0__abc_49347_n3179_1) );
  OR2X2 OR2X2_686 ( .A(u0__abc_49347_n3177_1), .B(u0__abc_49347_n3179_1), .Y(u0__abc_49347_n3180_1) );
  OR2X2 OR2X2_687 ( .A(u0__abc_49347_n2748_bF_buf5), .B(u0_tms0_18_), .Y(u0__abc_49347_n3181_1) );
  OR2X2 OR2X2_688 ( .A(u0__abc_49347_n3183_1), .B(u0__abc_49347_n3161), .Y(u0_tms_18__FF_INPUT) );
  OR2X2 OR2X2_689 ( .A(u0__abc_49347_n2728_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n3187_1) );
  OR2X2 OR2X2_69 ( .A(_abc_55805_n240_bF_buf4), .B(sp_tms_17_), .Y(_abc_55805_n341) );
  OR2X2 OR2X2_690 ( .A(1'b0), .B(1'b0), .Y(u0__abc_49347_n3188_1) );
  OR2X2 OR2X2_691 ( .A(u0__abc_49347_n3190), .B(u0__abc_49347_n3186_1), .Y(u0__abc_49347_n3191) );
  OR2X2 OR2X2_692 ( .A(u0__abc_49347_n3192), .B(u0__abc_49347_n3193), .Y(u0__abc_49347_n3194) );
  OR2X2 OR2X2_693 ( .A(u0__abc_49347_n3195), .B(u0__abc_49347_n3196), .Y(u0__abc_49347_n3197) );
  OR2X2 OR2X2_694 ( .A(u0__abc_49347_n3198), .B(u0__abc_49347_n3199), .Y(u0__abc_49347_n3200) );
  OR2X2 OR2X2_695 ( .A(u0__abc_49347_n3202), .B(u0_cs0_bF_buf3), .Y(u0__abc_49347_n3203) );
  OR2X2 OR2X2_696 ( .A(u0__abc_49347_n3201), .B(u0__abc_49347_n3203), .Y(u0__abc_49347_n3204) );
  OR2X2 OR2X2_697 ( .A(u0__abc_49347_n2748_bF_buf4), .B(u0_tms0_19_), .Y(u0__abc_49347_n3205) );
  OR2X2 OR2X2_698 ( .A(u0__abc_49347_n3207), .B(u0__abc_49347_n3185_1), .Y(u0_tms_19__FF_INPUT) );
  OR2X2 OR2X2_699 ( .A(u0__abc_49347_n2728_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n3211) );
  OR2X2 OR2X2_7 ( .A(_abc_55805_n240_bF_buf4), .B(spec_req_cs_1_bF_buf5), .Y(_abc_55805_n248) );
  OR2X2 OR2X2_70 ( .A(lmr_sel_bF_buf2), .B(tms_17_), .Y(_abc_55805_n342) );
  OR2X2 OR2X2_700 ( .A(1'b0), .B(1'b0), .Y(u0__abc_49347_n3212) );
  OR2X2 OR2X2_701 ( .A(u0__abc_49347_n3214), .B(u0__abc_49347_n3210), .Y(u0__abc_49347_n3215) );
  OR2X2 OR2X2_702 ( .A(u0__abc_49347_n3216), .B(u0__abc_49347_n3217), .Y(u0__abc_49347_n3218) );
  OR2X2 OR2X2_703 ( .A(u0__abc_49347_n3219), .B(u0__abc_49347_n3220), .Y(u0__abc_49347_n3221) );
  OR2X2 OR2X2_704 ( .A(u0__abc_49347_n3222), .B(u0__abc_49347_n3223), .Y(u0__abc_49347_n3224) );
  OR2X2 OR2X2_705 ( .A(u0__abc_49347_n3226), .B(u0_cs0_bF_buf2), .Y(u0__abc_49347_n3227) );
  OR2X2 OR2X2_706 ( .A(u0__abc_49347_n3225), .B(u0__abc_49347_n3227), .Y(u0__abc_49347_n3228) );
  OR2X2 OR2X2_707 ( .A(u0__abc_49347_n2748_bF_buf3), .B(u0_tms0_20_), .Y(u0__abc_49347_n3229) );
  OR2X2 OR2X2_708 ( .A(u0__abc_49347_n3231), .B(u0__abc_49347_n3209), .Y(u0_tms_20__FF_INPUT) );
  OR2X2 OR2X2_709 ( .A(u0__abc_49347_n2728_bF_buf2), .B(1'b0), .Y(u0__abc_49347_n3235) );
  OR2X2 OR2X2_71 ( .A(_abc_55805_n240_bF_buf3), .B(sp_tms_18_), .Y(_abc_55805_n344) );
  OR2X2 OR2X2_710 ( .A(1'b0), .B(1'b0), .Y(u0__abc_49347_n3236) );
  OR2X2 OR2X2_711 ( .A(u0__abc_49347_n3238), .B(u0__abc_49347_n3234), .Y(u0__abc_49347_n3239) );
  OR2X2 OR2X2_712 ( .A(u0__abc_49347_n3240), .B(u0__abc_49347_n3241), .Y(u0__abc_49347_n3242) );
  OR2X2 OR2X2_713 ( .A(u0__abc_49347_n3243), .B(u0__abc_49347_n3244), .Y(u0__abc_49347_n3245) );
  OR2X2 OR2X2_714 ( .A(u0__abc_49347_n3246), .B(u0__abc_49347_n3247), .Y(u0__abc_49347_n3248) );
  OR2X2 OR2X2_715 ( .A(u0__abc_49347_n3250), .B(u0_cs0_bF_buf1), .Y(u0__abc_49347_n3251) );
  OR2X2 OR2X2_716 ( .A(u0__abc_49347_n3249), .B(u0__abc_49347_n3251), .Y(u0__abc_49347_n3252) );
  OR2X2 OR2X2_717 ( .A(u0__abc_49347_n2748_bF_buf2), .B(u0_tms0_21_), .Y(u0__abc_49347_n3253) );
  OR2X2 OR2X2_718 ( .A(u0__abc_49347_n3255), .B(u0__abc_49347_n3233), .Y(u0_tms_21__FF_INPUT) );
  OR2X2 OR2X2_719 ( .A(u0__abc_49347_n2728_bF_buf1), .B(1'b0), .Y(u0__abc_49347_n3259) );
  OR2X2 OR2X2_72 ( .A(lmr_sel_bF_buf1), .B(tms_18_), .Y(_abc_55805_n345) );
  OR2X2 OR2X2_720 ( .A(1'b0), .B(1'b0), .Y(u0__abc_49347_n3260) );
  OR2X2 OR2X2_721 ( .A(u0__abc_49347_n3262), .B(u0__abc_49347_n3258), .Y(u0__abc_49347_n3263) );
  OR2X2 OR2X2_722 ( .A(u0__abc_49347_n3264), .B(u0__abc_49347_n3265), .Y(u0__abc_49347_n3266) );
  OR2X2 OR2X2_723 ( .A(u0__abc_49347_n3267), .B(u0__abc_49347_n3268), .Y(u0__abc_49347_n3269) );
  OR2X2 OR2X2_724 ( .A(u0__abc_49347_n3270), .B(u0__abc_49347_n3271), .Y(u0__abc_49347_n3272) );
  OR2X2 OR2X2_725 ( .A(u0__abc_49347_n3274), .B(u0_cs0_bF_buf0), .Y(u0__abc_49347_n3275) );
  OR2X2 OR2X2_726 ( .A(u0__abc_49347_n3273), .B(u0__abc_49347_n3275), .Y(u0__abc_49347_n3276) );
  OR2X2 OR2X2_727 ( .A(u0__abc_49347_n2748_bF_buf1), .B(u0_tms0_22_), .Y(u0__abc_49347_n3277) );
  OR2X2 OR2X2_728 ( .A(u0__abc_49347_n3279), .B(u0__abc_49347_n3257), .Y(u0_tms_22__FF_INPUT) );
  OR2X2 OR2X2_729 ( .A(u0__abc_49347_n2728_bF_buf0), .B(1'b0), .Y(u0__abc_49347_n3283) );
  OR2X2 OR2X2_73 ( .A(_abc_55805_n240_bF_buf2), .B(sp_tms_19_), .Y(_abc_55805_n347) );
  OR2X2 OR2X2_730 ( .A(1'b0), .B(1'b0), .Y(u0__abc_49347_n3284) );
  OR2X2 OR2X2_731 ( .A(u0__abc_49347_n3286), .B(u0__abc_49347_n3282), .Y(u0__abc_49347_n3287) );
  OR2X2 OR2X2_732 ( .A(u0__abc_49347_n3288), .B(u0__abc_49347_n3289), .Y(u0__abc_49347_n3290) );
  OR2X2 OR2X2_733 ( .A(u0__abc_49347_n3291), .B(u0__abc_49347_n3292), .Y(u0__abc_49347_n3293) );
  OR2X2 OR2X2_734 ( .A(u0__abc_49347_n3294), .B(u0__abc_49347_n3295), .Y(u0__abc_49347_n3296) );
  OR2X2 OR2X2_735 ( .A(u0__abc_49347_n3298), .B(u0_cs0_bF_buf5), .Y(u0__abc_49347_n3299) );
  OR2X2 OR2X2_736 ( .A(u0__abc_49347_n3297), .B(u0__abc_49347_n3299), .Y(u0__abc_49347_n3300) );
  OR2X2 OR2X2_737 ( .A(u0__abc_49347_n2748_bF_buf0), .B(u0_tms0_23_), .Y(u0__abc_49347_n3301) );
  OR2X2 OR2X2_738 ( .A(u0__abc_49347_n3303), .B(u0__abc_49347_n3281), .Y(u0_tms_23__FF_INPUT) );
  OR2X2 OR2X2_739 ( .A(u0__abc_49347_n2728_bF_buf5), .B(1'b0), .Y(u0__abc_49347_n3307) );
  OR2X2 OR2X2_74 ( .A(lmr_sel_bF_buf0), .B(tms_19_), .Y(_abc_55805_n348) );
  OR2X2 OR2X2_740 ( .A(1'b0), .B(1'b0), .Y(u0__abc_49347_n3308) );
  OR2X2 OR2X2_741 ( .A(u0__abc_49347_n3310), .B(u0__abc_49347_n3306), .Y(u0__abc_49347_n3311) );
  OR2X2 OR2X2_742 ( .A(u0__abc_49347_n3312), .B(u0__abc_49347_n3313), .Y(u0__abc_49347_n3314) );
  OR2X2 OR2X2_743 ( .A(u0__abc_49347_n3315), .B(u0__abc_49347_n3316), .Y(u0__abc_49347_n3317) );
  OR2X2 OR2X2_744 ( .A(u0__abc_49347_n3318), .B(u0__abc_49347_n3319), .Y(u0__abc_49347_n3320) );
  OR2X2 OR2X2_745 ( .A(u0__abc_49347_n3322), .B(u0_cs0_bF_buf4), .Y(u0__abc_49347_n3323) );
  OR2X2 OR2X2_746 ( .A(u0__abc_49347_n3321), .B(u0__abc_49347_n3323), .Y(u0__abc_49347_n3324) );
  OR2X2 OR2X2_747 ( .A(u0__abc_49347_n2748_bF_buf5), .B(u0_tms0_24_), .Y(u0__abc_49347_n3325) );
  OR2X2 OR2X2_748 ( .A(u0__abc_49347_n3327), .B(u0__abc_49347_n3305), .Y(u0_tms_24__FF_INPUT) );
  OR2X2 OR2X2_749 ( .A(u0__abc_49347_n2728_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n3331) );
  OR2X2 OR2X2_75 ( .A(_abc_55805_n240_bF_buf1), .B(sp_tms_20_), .Y(_abc_55805_n350) );
  OR2X2 OR2X2_750 ( .A(1'b0), .B(1'b0), .Y(u0__abc_49347_n3332) );
  OR2X2 OR2X2_751 ( .A(u0__abc_49347_n3334), .B(u0__abc_49347_n3330), .Y(u0__abc_49347_n3335) );
  OR2X2 OR2X2_752 ( .A(u0__abc_49347_n3336), .B(u0__abc_49347_n3337), .Y(u0__abc_49347_n3338) );
  OR2X2 OR2X2_753 ( .A(u0__abc_49347_n3339), .B(u0__abc_49347_n3340), .Y(u0__abc_49347_n3341) );
  OR2X2 OR2X2_754 ( .A(u0__abc_49347_n3342), .B(u0__abc_49347_n3343), .Y(u0__abc_49347_n3344) );
  OR2X2 OR2X2_755 ( .A(u0__abc_49347_n3346), .B(u0_cs0_bF_buf3), .Y(u0__abc_49347_n3347) );
  OR2X2 OR2X2_756 ( .A(u0__abc_49347_n3345), .B(u0__abc_49347_n3347), .Y(u0__abc_49347_n3348) );
  OR2X2 OR2X2_757 ( .A(u0__abc_49347_n2748_bF_buf4), .B(u0_tms0_25_), .Y(u0__abc_49347_n3349) );
  OR2X2 OR2X2_758 ( .A(u0__abc_49347_n3351), .B(u0__abc_49347_n3329), .Y(u0_tms_25__FF_INPUT) );
  OR2X2 OR2X2_759 ( .A(u0__abc_49347_n2728_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n3355) );
  OR2X2 OR2X2_76 ( .A(lmr_sel_bF_buf6), .B(tms_20_), .Y(_abc_55805_n351) );
  OR2X2 OR2X2_760 ( .A(1'b0), .B(1'b0), .Y(u0__abc_49347_n3356) );
  OR2X2 OR2X2_761 ( .A(u0__abc_49347_n3358), .B(u0__abc_49347_n3354), .Y(u0__abc_49347_n3359) );
  OR2X2 OR2X2_762 ( .A(u0__abc_49347_n3360), .B(u0__abc_49347_n3361), .Y(u0__abc_49347_n3362) );
  OR2X2 OR2X2_763 ( .A(u0__abc_49347_n3363), .B(u0__abc_49347_n3364), .Y(u0__abc_49347_n3365) );
  OR2X2 OR2X2_764 ( .A(u0__abc_49347_n3366), .B(u0__abc_49347_n3367), .Y(u0__abc_49347_n3368) );
  OR2X2 OR2X2_765 ( .A(u0__abc_49347_n3370), .B(u0_cs0_bF_buf2), .Y(u0__abc_49347_n3371) );
  OR2X2 OR2X2_766 ( .A(u0__abc_49347_n3369), .B(u0__abc_49347_n3371), .Y(u0__abc_49347_n3372) );
  OR2X2 OR2X2_767 ( .A(u0__abc_49347_n2748_bF_buf3), .B(u0_tms0_26_), .Y(u0__abc_49347_n3373) );
  OR2X2 OR2X2_768 ( .A(u0__abc_49347_n3375), .B(u0__abc_49347_n3353), .Y(u0_tms_26__FF_INPUT) );
  OR2X2 OR2X2_769 ( .A(u0__abc_49347_n2728_bF_buf2), .B(1'b0), .Y(u0__abc_49347_n3379) );
  OR2X2 OR2X2_77 ( .A(_abc_55805_n240_bF_buf0), .B(sp_tms_21_), .Y(_abc_55805_n353) );
  OR2X2 OR2X2_770 ( .A(1'b0), .B(1'b0), .Y(u0__abc_49347_n3380) );
  OR2X2 OR2X2_771 ( .A(u0__abc_49347_n3382), .B(u0__abc_49347_n3378), .Y(u0__abc_49347_n3383) );
  OR2X2 OR2X2_772 ( .A(u0__abc_49347_n3384), .B(u0__abc_49347_n3385), .Y(u0__abc_49347_n3386) );
  OR2X2 OR2X2_773 ( .A(u0__abc_49347_n3387), .B(u0__abc_49347_n3388), .Y(u0__abc_49347_n3389) );
  OR2X2 OR2X2_774 ( .A(u0__abc_49347_n3390), .B(u0__abc_49347_n3391), .Y(u0__abc_49347_n3392) );
  OR2X2 OR2X2_775 ( .A(u0__abc_49347_n3394), .B(u0_cs0_bF_buf1), .Y(u0__abc_49347_n3395) );
  OR2X2 OR2X2_776 ( .A(u0__abc_49347_n3393), .B(u0__abc_49347_n3395), .Y(u0__abc_49347_n3396) );
  OR2X2 OR2X2_777 ( .A(u0__abc_49347_n2748_bF_buf2), .B(u0_tms0_27_), .Y(u0__abc_49347_n3397) );
  OR2X2 OR2X2_778 ( .A(u0__abc_49347_n3399), .B(u0__abc_49347_n3377), .Y(u0_tms_27__FF_INPUT) );
  OR2X2 OR2X2_779 ( .A(u0__abc_49347_n2728_bF_buf1), .B(1'b0), .Y(u0__abc_49347_n3523) );
  OR2X2 OR2X2_78 ( .A(lmr_sel_bF_buf5), .B(tms_21_), .Y(_abc_55805_n354) );
  OR2X2 OR2X2_780 ( .A(1'b0), .B(1'b0), .Y(u0__abc_49347_n3524) );
  OR2X2 OR2X2_781 ( .A(u0__abc_49347_n3526), .B(u0__abc_49347_n3522), .Y(u0__abc_49347_n3527) );
  OR2X2 OR2X2_782 ( .A(u0__abc_49347_n3528), .B(u0__abc_49347_n3529), .Y(u0__abc_49347_n3530) );
  OR2X2 OR2X2_783 ( .A(u0__abc_49347_n3531), .B(u0__abc_49347_n3532), .Y(u0__abc_49347_n3533) );
  OR2X2 OR2X2_784 ( .A(u0__abc_49347_n3534), .B(u0__abc_49347_n3535), .Y(u0__abc_49347_n3536) );
  OR2X2 OR2X2_785 ( .A(u0__abc_49347_n3538), .B(u0_cs0_bF_buf0), .Y(u0__abc_49347_n3539) );
  OR2X2 OR2X2_786 ( .A(u0__abc_49347_n3537), .B(u0__abc_49347_n3539), .Y(u0__abc_49347_n3540) );
  OR2X2 OR2X2_787 ( .A(u0__abc_49347_n2748_bF_buf1), .B(u0_csc0_1_), .Y(u0__abc_49347_n3541) );
  OR2X2 OR2X2_788 ( .A(u0__abc_49347_n3543), .B(u0__abc_49347_n3521), .Y(u0_csc_1__FF_INPUT) );
  OR2X2 OR2X2_789 ( .A(u0__abc_49347_n2728_bF_buf0), .B(1'b0), .Y(u0__abc_49347_n3547) );
  OR2X2 OR2X2_79 ( .A(_abc_55805_n240_bF_buf5), .B(sp_tms_22_), .Y(_abc_55805_n356) );
  OR2X2 OR2X2_790 ( .A(1'b0), .B(1'b0), .Y(u0__abc_49347_n3548) );
  OR2X2 OR2X2_791 ( .A(u0__abc_49347_n3550), .B(u0__abc_49347_n3546), .Y(u0__abc_49347_n3551) );
  OR2X2 OR2X2_792 ( .A(u0__abc_49347_n3552), .B(u0__abc_49347_n3553), .Y(u0__abc_49347_n3554) );
  OR2X2 OR2X2_793 ( .A(u0__abc_49347_n3555), .B(u0__abc_49347_n3556), .Y(u0__abc_49347_n3557) );
  OR2X2 OR2X2_794 ( .A(u0__abc_49347_n3558), .B(u0__abc_49347_n3559), .Y(u0__abc_49347_n3560) );
  OR2X2 OR2X2_795 ( .A(u0__abc_49347_n3562), .B(u0_cs0_bF_buf5), .Y(u0__abc_49347_n3563) );
  OR2X2 OR2X2_796 ( .A(u0__abc_49347_n3561), .B(u0__abc_49347_n3563), .Y(u0__abc_49347_n3564) );
  OR2X2 OR2X2_797 ( .A(u0__abc_49347_n2748_bF_buf0), .B(u0_csc0_2_), .Y(u0__abc_49347_n3565) );
  OR2X2 OR2X2_798 ( .A(u0__abc_49347_n3567), .B(u0__abc_49347_n3545), .Y(u0_csc_2__FF_INPUT) );
  OR2X2 OR2X2_799 ( .A(u0__abc_49347_n2728_bF_buf5), .B(1'b0), .Y(u0__abc_49347_n3571) );
  OR2X2 OR2X2_8 ( .A(lmr_sel_bF_buf5), .B(cs_1_), .Y(_abc_55805_n249) );
  OR2X2 OR2X2_80 ( .A(lmr_sel_bF_buf4), .B(tms_22_), .Y(_abc_55805_n357) );
  OR2X2 OR2X2_800 ( .A(1'b0), .B(1'b0), .Y(u0__abc_49347_n3572) );
  OR2X2 OR2X2_801 ( .A(u0__abc_49347_n3574), .B(u0__abc_49347_n3570), .Y(u0__abc_49347_n3575) );
  OR2X2 OR2X2_802 ( .A(u0__abc_49347_n3576), .B(u0__abc_49347_n3577), .Y(u0__abc_49347_n3578) );
  OR2X2 OR2X2_803 ( .A(u0__abc_49347_n3579), .B(u0__abc_49347_n3580), .Y(u0__abc_49347_n3581) );
  OR2X2 OR2X2_804 ( .A(u0__abc_49347_n3582), .B(u0__abc_49347_n3583), .Y(u0__abc_49347_n3584) );
  OR2X2 OR2X2_805 ( .A(u0__abc_49347_n3586), .B(u0_cs0_bF_buf4), .Y(u0__abc_49347_n3587) );
  OR2X2 OR2X2_806 ( .A(u0__abc_49347_n3585), .B(u0__abc_49347_n3587), .Y(u0__abc_49347_n3588) );
  OR2X2 OR2X2_807 ( .A(u0__abc_49347_n2748_bF_buf5), .B(u0_csc0_3_), .Y(u0__abc_49347_n3589) );
  OR2X2 OR2X2_808 ( .A(u0__abc_49347_n3591), .B(u0__abc_49347_n3569), .Y(u0_csc_3__FF_INPUT) );
  OR2X2 OR2X2_809 ( .A(u0__abc_49347_n2728_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n3595) );
  OR2X2 OR2X2_81 ( .A(_abc_55805_n240_bF_buf4), .B(sp_tms_23_), .Y(_abc_55805_n359) );
  OR2X2 OR2X2_810 ( .A(1'b0), .B(1'b0), .Y(u0__abc_49347_n3596) );
  OR2X2 OR2X2_811 ( .A(u0__abc_49347_n3598), .B(u0__abc_49347_n3594), .Y(u0__abc_49347_n3599) );
  OR2X2 OR2X2_812 ( .A(u0__abc_49347_n3600), .B(u0__abc_49347_n3601), .Y(u0__abc_49347_n3602) );
  OR2X2 OR2X2_813 ( .A(u0__abc_49347_n3603), .B(u0__abc_49347_n3604), .Y(u0__abc_49347_n3605) );
  OR2X2 OR2X2_814 ( .A(u0__abc_49347_n3606), .B(u0__abc_49347_n3607), .Y(u0__abc_49347_n3608) );
  OR2X2 OR2X2_815 ( .A(u0__abc_49347_n3610), .B(u0_cs0_bF_buf3), .Y(u0__abc_49347_n3611) );
  OR2X2 OR2X2_816 ( .A(u0__abc_49347_n3609), .B(u0__abc_49347_n3611), .Y(u0__abc_49347_n3612) );
  OR2X2 OR2X2_817 ( .A(u0__abc_49347_n2748_bF_buf4), .B(u0_csc0_4_), .Y(u0__abc_49347_n3613) );
  OR2X2 OR2X2_818 ( .A(u0__abc_49347_n3615), .B(u0__abc_49347_n3593), .Y(u0_csc_4__FF_INPUT) );
  OR2X2 OR2X2_819 ( .A(u0__abc_49347_n2728_bF_buf3), .B(1'b0), .Y(u0__abc_49347_n3619) );
  OR2X2 OR2X2_82 ( .A(lmr_sel_bF_buf3), .B(tms_23_), .Y(_abc_55805_n360) );
  OR2X2 OR2X2_820 ( .A(1'b0), .B(1'b0), .Y(u0__abc_49347_n3620) );
  OR2X2 OR2X2_821 ( .A(u0__abc_49347_n3622), .B(u0__abc_49347_n3618), .Y(u0__abc_49347_n3623) );
  OR2X2 OR2X2_822 ( .A(u0__abc_49347_n3624), .B(u0__abc_49347_n3625), .Y(u0__abc_49347_n3626) );
  OR2X2 OR2X2_823 ( .A(u0__abc_49347_n3627), .B(u0__abc_49347_n3628), .Y(u0__abc_49347_n3629) );
  OR2X2 OR2X2_824 ( .A(u0__abc_49347_n3630), .B(u0__abc_49347_n3631), .Y(u0__abc_49347_n3632) );
  OR2X2 OR2X2_825 ( .A(u0__abc_49347_n3634), .B(u0_cs0_bF_buf2), .Y(u0__abc_49347_n3635) );
  OR2X2 OR2X2_826 ( .A(u0__abc_49347_n3633), .B(u0__abc_49347_n3635), .Y(u0__abc_49347_n3636) );
  OR2X2 OR2X2_827 ( .A(u0__abc_49347_n2748_bF_buf3), .B(u0_csc0_5_), .Y(u0__abc_49347_n3637) );
  OR2X2 OR2X2_828 ( .A(u0__abc_49347_n3639), .B(u0__abc_49347_n3617), .Y(u0_csc_5__FF_INPUT) );
  OR2X2 OR2X2_829 ( .A(u0__abc_49347_n2728_bF_buf2), .B(1'b0), .Y(u0__abc_49347_n3643) );
  OR2X2 OR2X2_83 ( .A(_abc_55805_n240_bF_buf3), .B(sp_tms_24_), .Y(_abc_55805_n362) );
  OR2X2 OR2X2_830 ( .A(1'b0), .B(1'b0), .Y(u0__abc_49347_n3644) );
  OR2X2 OR2X2_831 ( .A(u0__abc_49347_n3646), .B(u0__abc_49347_n3642), .Y(u0__abc_49347_n3647) );
  OR2X2 OR2X2_832 ( .A(u0__abc_49347_n3648), .B(u0__abc_49347_n3649), .Y(u0__abc_49347_n3650) );
  OR2X2 OR2X2_833 ( .A(u0__abc_49347_n3651), .B(u0__abc_49347_n3652), .Y(u0__abc_49347_n3653) );
  OR2X2 OR2X2_834 ( .A(u0__abc_49347_n3654), .B(u0__abc_49347_n3655), .Y(u0__abc_49347_n3656) );
  OR2X2 OR2X2_835 ( .A(u0__abc_49347_n3658), .B(u0_cs0_bF_buf1), .Y(u0__abc_49347_n3659) );
  OR2X2 OR2X2_836 ( .A(u0__abc_49347_n3657), .B(u0__abc_49347_n3659), .Y(u0__abc_49347_n3660) );
  OR2X2 OR2X2_837 ( .A(u0__abc_49347_n2748_bF_buf2), .B(u0_csc0_6_), .Y(u0__abc_49347_n3661) );
  OR2X2 OR2X2_838 ( .A(u0__abc_49347_n3663), .B(u0__abc_49347_n3641), .Y(u0_csc_6__FF_INPUT) );
  OR2X2 OR2X2_839 ( .A(u0__abc_49347_n2728_bF_buf1), .B(1'b0), .Y(u0__abc_49347_n3667) );
  OR2X2 OR2X2_84 ( .A(lmr_sel_bF_buf2), .B(tms_24_), .Y(_abc_55805_n363) );
  OR2X2 OR2X2_840 ( .A(1'b0), .B(1'b0), .Y(u0__abc_49347_n3668) );
  OR2X2 OR2X2_841 ( .A(u0__abc_49347_n3670), .B(u0__abc_49347_n3666), .Y(u0__abc_49347_n3671) );
  OR2X2 OR2X2_842 ( .A(u0__abc_49347_n3672), .B(u0__abc_49347_n3673), .Y(u0__abc_49347_n3674) );
  OR2X2 OR2X2_843 ( .A(u0__abc_49347_n3675), .B(u0__abc_49347_n3676), .Y(u0__abc_49347_n3677) );
  OR2X2 OR2X2_844 ( .A(u0__abc_49347_n3678), .B(u0__abc_49347_n3679), .Y(u0__abc_49347_n3680) );
  OR2X2 OR2X2_845 ( .A(u0__abc_49347_n3682), .B(u0_cs0_bF_buf0), .Y(u0__abc_49347_n3683) );
  OR2X2 OR2X2_846 ( .A(u0__abc_49347_n3681), .B(u0__abc_49347_n3683), .Y(u0__abc_49347_n3684) );
  OR2X2 OR2X2_847 ( .A(u0__abc_49347_n2748_bF_buf1), .B(u0_csc0_7_), .Y(u0__abc_49347_n3685) );
  OR2X2 OR2X2_848 ( .A(u0__abc_49347_n3687), .B(u0__abc_49347_n3665), .Y(u0_csc_7__FF_INPUT) );
  OR2X2 OR2X2_849 ( .A(u0__abc_49347_n2728_bF_buf0), .B(1'b0), .Y(u0__abc_49347_n3715) );
  OR2X2 OR2X2_85 ( .A(_abc_55805_n240_bF_buf2), .B(sp_tms_25_), .Y(_abc_55805_n365) );
  OR2X2 OR2X2_850 ( .A(1'b0), .B(1'b0), .Y(u0__abc_49347_n3716) );
  OR2X2 OR2X2_851 ( .A(u0__abc_49347_n3718), .B(u0__abc_49347_n3714), .Y(u0__abc_49347_n3719) );
  OR2X2 OR2X2_852 ( .A(u0__abc_49347_n3720), .B(u0__abc_49347_n3721), .Y(u0__abc_49347_n3722) );
  OR2X2 OR2X2_853 ( .A(u0__abc_49347_n3723), .B(u0__abc_49347_n3724), .Y(u0__abc_49347_n3725) );
  OR2X2 OR2X2_854 ( .A(u0__abc_49347_n3726), .B(u0__abc_49347_n3727), .Y(u0__abc_49347_n3728) );
  OR2X2 OR2X2_855 ( .A(u0__abc_49347_n3730), .B(u0_cs0_bF_buf5), .Y(u0__abc_49347_n3731) );
  OR2X2 OR2X2_856 ( .A(u0__abc_49347_n3729), .B(u0__abc_49347_n3731), .Y(u0__abc_49347_n3732) );
  OR2X2 OR2X2_857 ( .A(u0__abc_49347_n2748_bF_buf0), .B(u0_csc0_9_), .Y(u0__abc_49347_n3733) );
  OR2X2 OR2X2_858 ( .A(u0__abc_49347_n3735), .B(u0__abc_49347_n3713), .Y(u0_csc_9__FF_INPUT) );
  OR2X2 OR2X2_859 ( .A(u0__abc_49347_n2728_bF_buf5), .B(1'b0), .Y(u0__abc_49347_n3739) );
  OR2X2 OR2X2_86 ( .A(lmr_sel_bF_buf1), .B(tms_25_), .Y(_abc_55805_n366) );
  OR2X2 OR2X2_860 ( .A(1'b0), .B(1'b0), .Y(u0__abc_49347_n3740) );
  OR2X2 OR2X2_861 ( .A(u0__abc_49347_n3742), .B(u0__abc_49347_n3738), .Y(u0__abc_49347_n3743) );
  OR2X2 OR2X2_862 ( .A(u0__abc_49347_n3744), .B(u0__abc_49347_n3745), .Y(u0__abc_49347_n3746) );
  OR2X2 OR2X2_863 ( .A(u0__abc_49347_n3747), .B(u0__abc_49347_n3748), .Y(u0__abc_49347_n3749) );
  OR2X2 OR2X2_864 ( .A(u0__abc_49347_n3750), .B(u0__abc_49347_n3751), .Y(u0__abc_49347_n3752) );
  OR2X2 OR2X2_865 ( .A(u0__abc_49347_n3754), .B(u0_cs0_bF_buf4), .Y(u0__abc_49347_n3755) );
  OR2X2 OR2X2_866 ( .A(u0__abc_49347_n3753), .B(u0__abc_49347_n3755), .Y(u0__abc_49347_n3756) );
  OR2X2 OR2X2_867 ( .A(u0__abc_49347_n2748_bF_buf5), .B(u0_csc0_10_), .Y(u0__abc_49347_n3757) );
  OR2X2 OR2X2_868 ( .A(u0__abc_49347_n3759), .B(u0__abc_49347_n3737), .Y(u0_csc_10__FF_INPUT) );
  OR2X2 OR2X2_869 ( .A(u0__abc_49347_n2728_bF_buf4), .B(1'b0), .Y(u0__abc_49347_n3763) );
  OR2X2 OR2X2_87 ( .A(_abc_55805_n240_bF_buf1), .B(sp_tms_26_), .Y(_abc_55805_n368) );
  OR2X2 OR2X2_870 ( .A(1'b0), .B(1'b0), .Y(u0__abc_49347_n3764) );
  OR2X2 OR2X2_871 ( .A(u0__abc_49347_n3766), .B(u0__abc_49347_n3762), .Y(u0__abc_49347_n3767) );
  OR2X2 OR2X2_872 ( .A(u0__abc_49347_n3768), .B(u0__abc_49347_n3769), .Y(u0__abc_49347_n3770) );
  OR2X2 OR2X2_873 ( .A(u0__abc_49347_n3771), .B(u0__abc_49347_n3772), .Y(u0__abc_49347_n3773) );
  OR2X2 OR2X2_874 ( .A(u0__abc_49347_n3774), .B(u0__abc_49347_n3775), .Y(u0__abc_49347_n3776) );
  OR2X2 OR2X2_875 ( .A(u0__abc_49347_n3778), .B(u0_cs0_bF_buf3), .Y(u0__abc_49347_n3779) );
  OR2X2 OR2X2_876 ( .A(u0__abc_49347_n3777), .B(u0__abc_49347_n3779), .Y(u0__abc_49347_n3780) );
  OR2X2 OR2X2_877 ( .A(u0__abc_49347_n2748_bF_buf4), .B(u0_csc0_11_), .Y(u0__abc_49347_n3781) );
  OR2X2 OR2X2_878 ( .A(u0__abc_49347_n3783), .B(u0__abc_49347_n3761), .Y(u0_csc_11__FF_INPUT) );
  OR2X2 OR2X2_879 ( .A(1'b0), .B(1'b0), .Y(u0__abc_49347_n4266) );
  OR2X2 OR2X2_88 ( .A(lmr_sel_bF_buf0), .B(tms_26_), .Y(_abc_55805_n369) );
  OR2X2 OR2X2_880 ( .A(u0_u4_wp_err), .B(u0_u5_wp_err), .Y(u0__abc_49347_n4267) );
  OR2X2 OR2X2_881 ( .A(u0__abc_49347_n4266), .B(u0__abc_49347_n4267), .Y(u0__abc_49347_n4268) );
  OR2X2 OR2X2_882 ( .A(u0_u2_wp_err), .B(u0_u3_wp_err), .Y(u0__abc_49347_n4269) );
  OR2X2 OR2X2_883 ( .A(u0_u0_wp_err), .B(u0_u1_wp_err), .Y(u0__abc_49347_n4270) );
  OR2X2 OR2X2_884 ( .A(u0__abc_49347_n4269), .B(u0__abc_49347_n4270), .Y(u0__abc_49347_n4271) );
  OR2X2 OR2X2_885 ( .A(u0__abc_49347_n4268), .B(u0__abc_49347_n4271), .Y(u0__abc_49347_n4272) );
  OR2X2 OR2X2_886 ( .A(u0__abc_49347_n4273), .B(u0__abc_49347_n4276), .Y(u0_wp_err_FF_INPUT) );
  OR2X2 OR2X2_887 ( .A(cs_le_bF_buf3), .B(cs_0_), .Y(u0__abc_49347_n4278) );
  OR2X2 OR2X2_888 ( .A(u0__abc_49347_n4279), .B(u0_cs0_bF_buf2), .Y(u0__abc_49347_n4280) );
  OR2X2 OR2X2_889 ( .A(cs_le_bF_buf1), .B(cs_1_), .Y(u0__abc_49347_n4282) );
  OR2X2 OR2X2_89 ( .A(_abc_55805_n240_bF_buf0), .B(sp_tms_27_), .Y(_abc_55805_n371) );
  OR2X2 OR2X2_890 ( .A(u0__abc_49347_n4279), .B(u0_cs1_bF_buf2), .Y(u0__abc_49347_n4283) );
  OR2X2 OR2X2_891 ( .A(cs_le_bF_buf0), .B(cs_2_), .Y(u0__abc_49347_n4285) );
  OR2X2 OR2X2_892 ( .A(u0__abc_49347_n4279), .B(u0_cs2_bF_buf2), .Y(u0__abc_49347_n4286) );
  OR2X2 OR2X2_893 ( .A(cs_le_bF_buf4), .B(cs_3_), .Y(u0__abc_49347_n4288) );
  OR2X2 OR2X2_894 ( .A(u0__abc_49347_n4279), .B(u0_cs3_bF_buf2), .Y(u0__abc_49347_n4289) );
  OR2X2 OR2X2_895 ( .A(cs_le_bF_buf3), .B(cs_4_), .Y(u0__abc_49347_n4291) );
  OR2X2 OR2X2_896 ( .A(u0__abc_49347_n4279), .B(u0_cs4_bF_buf2), .Y(u0__abc_49347_n4292) );
  OR2X2 OR2X2_897 ( .A(cs_le_bF_buf2), .B(cs_5_), .Y(u0__abc_49347_n4294) );
  OR2X2 OR2X2_898 ( .A(u0__abc_49347_n4279), .B(u0_cs5_bF_buf2), .Y(u0__abc_49347_n4295) );
  OR2X2 OR2X2_899 ( .A(cs_le_bF_buf1), .B(cs_6_), .Y(u0__abc_49347_n4297) );
  OR2X2 OR2X2_9 ( .A(_abc_55805_n250), .B(_abc_55805_n237_1), .Y(_abc_55805_n251) );
  OR2X2 OR2X2_90 ( .A(lmr_sel_bF_buf6), .B(tms_27_), .Y(_abc_55805_n372) );
  OR2X2 OR2X2_900 ( .A(u0__abc_49347_n4279), .B(1'b0), .Y(u0__abc_49347_n4298) );
  OR2X2 OR2X2_901 ( .A(cs_le_bF_buf0), .B(cs_7_), .Y(u0__abc_49347_n4300) );
  OR2X2 OR2X2_902 ( .A(u0__abc_49347_n4279), .B(1'b0), .Y(u0__abc_49347_n4301) );
  OR2X2 OR2X2_903 ( .A(_auto_iopadmap_cc_313_execute_56321_0_), .B(u0_rst_r3_bF_buf4), .Y(u0__abc_49347_n4303) );
  OR2X2 OR2X2_904 ( .A(u0__abc_49347_n4304_bF_buf4), .B(mc_data_ir_0_), .Y(u0__abc_49347_n4305) );
  OR2X2 OR2X2_905 ( .A(u0_rst_r3_bF_buf2), .B(_auto_iopadmap_cc_313_execute_56321_1_), .Y(u0__abc_49347_n4307) );
  OR2X2 OR2X2_906 ( .A(u0__abc_49347_n4304_bF_buf3), .B(mc_data_ir_1_), .Y(u0__abc_49347_n4308) );
  OR2X2 OR2X2_907 ( .A(u0_rst_r3_bF_buf1), .B(_auto_iopadmap_cc_313_execute_56321_2_), .Y(u0__abc_49347_n4310) );
  OR2X2 OR2X2_908 ( .A(u0__abc_49347_n4304_bF_buf2), .B(mc_data_ir_2_), .Y(u0__abc_49347_n4311) );
  OR2X2 OR2X2_909 ( .A(u0_rst_r3_bF_buf0), .B(_auto_iopadmap_cc_313_execute_56321_3_), .Y(u0__abc_49347_n4313) );
  OR2X2 OR2X2_91 ( .A(_abc_55805_n240_bF_buf5), .B(sp_csc_1_), .Y(_abc_55805_n389) );
  OR2X2 OR2X2_910 ( .A(u0__abc_49347_n4304_bF_buf1), .B(mc_data_ir_3_), .Y(u0__abc_49347_n4314) );
  OR2X2 OR2X2_911 ( .A(u0_rst_r3_bF_buf4), .B(_auto_iopadmap_cc_313_execute_56321_4_), .Y(u0__abc_49347_n4316) );
  OR2X2 OR2X2_912 ( .A(u0__abc_49347_n4304_bF_buf0), .B(mc_data_ir_4_), .Y(u0__abc_49347_n4317) );
  OR2X2 OR2X2_913 ( .A(u0_rst_r3_bF_buf3), .B(_auto_iopadmap_cc_313_execute_56321_5_), .Y(u0__abc_49347_n4319) );
  OR2X2 OR2X2_914 ( .A(u0__abc_49347_n4304_bF_buf4), .B(mc_data_ir_5_), .Y(u0__abc_49347_n4320) );
  OR2X2 OR2X2_915 ( .A(u0_rst_r3_bF_buf2), .B(_auto_iopadmap_cc_313_execute_56321_6_), .Y(u0__abc_49347_n4322) );
  OR2X2 OR2X2_916 ( .A(u0__abc_49347_n4304_bF_buf3), .B(mc_data_ir_6_), .Y(u0__abc_49347_n4323) );
  OR2X2 OR2X2_917 ( .A(u0_rst_r3_bF_buf1), .B(_auto_iopadmap_cc_313_execute_56321_7_), .Y(u0__abc_49347_n4325) );
  OR2X2 OR2X2_918 ( .A(u0__abc_49347_n4304_bF_buf2), .B(mc_data_ir_7_), .Y(u0__abc_49347_n4326) );
  OR2X2 OR2X2_919 ( .A(u0_rst_r3_bF_buf0), .B(_auto_iopadmap_cc_313_execute_56321_8_), .Y(u0__abc_49347_n4328) );
  OR2X2 OR2X2_92 ( .A(lmr_sel_bF_buf5), .B(csc_1_), .Y(_abc_55805_n390) );
  OR2X2 OR2X2_920 ( .A(u0__abc_49347_n4304_bF_buf1), .B(mc_data_ir_8_), .Y(u0__abc_49347_n4329) );
  OR2X2 OR2X2_921 ( .A(u0_rst_r3_bF_buf4), .B(_auto_iopadmap_cc_313_execute_56321_9_), .Y(u0__abc_49347_n4331) );
  OR2X2 OR2X2_922 ( .A(u0__abc_49347_n4304_bF_buf0), .B(mc_data_ir_9_), .Y(u0__abc_49347_n4332) );
  OR2X2 OR2X2_923 ( .A(u0_rst_r3_bF_buf3), .B(_auto_iopadmap_cc_313_execute_56321_10_), .Y(u0__abc_49347_n4334) );
  OR2X2 OR2X2_924 ( .A(u0__abc_49347_n4304_bF_buf4), .B(mc_data_ir_10_), .Y(u0__abc_49347_n4335) );
  OR2X2 OR2X2_925 ( .A(u0_rst_r3_bF_buf2), .B(_auto_iopadmap_cc_313_execute_56321_11_), .Y(u0__abc_49347_n4337) );
  OR2X2 OR2X2_926 ( .A(u0__abc_49347_n4304_bF_buf3), .B(mc_data_ir_11_), .Y(u0__abc_49347_n4338) );
  OR2X2 OR2X2_927 ( .A(u0_rst_r3_bF_buf1), .B(_auto_iopadmap_cc_313_execute_56321_12_), .Y(u0__abc_49347_n4340) );
  OR2X2 OR2X2_928 ( .A(u0__abc_49347_n4304_bF_buf2), .B(mc_data_ir_12_), .Y(u0__abc_49347_n4341) );
  OR2X2 OR2X2_929 ( .A(u0_rst_r3_bF_buf0), .B(_auto_iopadmap_cc_313_execute_56321_13_), .Y(u0__abc_49347_n4343) );
  OR2X2 OR2X2_93 ( .A(_abc_55805_n240_bF_buf4), .B(sp_csc_2_), .Y(_abc_55805_n392) );
  OR2X2 OR2X2_930 ( .A(u0__abc_49347_n4304_bF_buf1), .B(mc_data_ir_13_), .Y(u0__abc_49347_n4344) );
  OR2X2 OR2X2_931 ( .A(u0_rst_r3_bF_buf4), .B(_auto_iopadmap_cc_313_execute_56321_14_), .Y(u0__abc_49347_n4346) );
  OR2X2 OR2X2_932 ( .A(u0__abc_49347_n4304_bF_buf0), .B(mc_data_ir_14_), .Y(u0__abc_49347_n4347) );
  OR2X2 OR2X2_933 ( .A(u0_rst_r3_bF_buf3), .B(_auto_iopadmap_cc_313_execute_56321_15_), .Y(u0__abc_49347_n4349) );
  OR2X2 OR2X2_934 ( .A(u0__abc_49347_n4304_bF_buf4), .B(mc_data_ir_15_), .Y(u0__abc_49347_n4350) );
  OR2X2 OR2X2_935 ( .A(u0_rst_r3_bF_buf2), .B(_auto_iopadmap_cc_313_execute_56321_16_), .Y(u0__abc_49347_n4352) );
  OR2X2 OR2X2_936 ( .A(u0__abc_49347_n4304_bF_buf3), .B(mc_data_ir_16_), .Y(u0__abc_49347_n4353) );
  OR2X2 OR2X2_937 ( .A(u0_rst_r3_bF_buf1), .B(_auto_iopadmap_cc_313_execute_56321_17_), .Y(u0__abc_49347_n4355) );
  OR2X2 OR2X2_938 ( .A(u0__abc_49347_n4304_bF_buf2), .B(mc_data_ir_17_), .Y(u0__abc_49347_n4356) );
  OR2X2 OR2X2_939 ( .A(u0_rst_r3_bF_buf0), .B(_auto_iopadmap_cc_313_execute_56321_18_), .Y(u0__abc_49347_n4358) );
  OR2X2 OR2X2_94 ( .A(lmr_sel_bF_buf4), .B(csc_2_), .Y(_abc_55805_n393) );
  OR2X2 OR2X2_940 ( .A(u0__abc_49347_n4304_bF_buf1), .B(mc_data_ir_18_), .Y(u0__abc_49347_n4359) );
  OR2X2 OR2X2_941 ( .A(u0_rst_r3_bF_buf4), .B(_auto_iopadmap_cc_313_execute_56321_19_), .Y(u0__abc_49347_n4361) );
  OR2X2 OR2X2_942 ( .A(u0__abc_49347_n4304_bF_buf0), .B(mc_data_ir_19_), .Y(u0__abc_49347_n4362) );
  OR2X2 OR2X2_943 ( .A(u0_rst_r3_bF_buf3), .B(_auto_iopadmap_cc_313_execute_56321_20_), .Y(u0__abc_49347_n4364) );
  OR2X2 OR2X2_944 ( .A(u0__abc_49347_n4304_bF_buf4), .B(mc_data_ir_20_), .Y(u0__abc_49347_n4365) );
  OR2X2 OR2X2_945 ( .A(u0_rst_r3_bF_buf2), .B(_auto_iopadmap_cc_313_execute_56321_21_), .Y(u0__abc_49347_n4367) );
  OR2X2 OR2X2_946 ( .A(u0__abc_49347_n4304_bF_buf3), .B(mc_data_ir_21_), .Y(u0__abc_49347_n4368) );
  OR2X2 OR2X2_947 ( .A(u0_rst_r3_bF_buf1), .B(_auto_iopadmap_cc_313_execute_56321_22_), .Y(u0__abc_49347_n4370) );
  OR2X2 OR2X2_948 ( .A(u0__abc_49347_n4304_bF_buf2), .B(mc_data_ir_22_), .Y(u0__abc_49347_n4371) );
  OR2X2 OR2X2_949 ( .A(u0_rst_r3_bF_buf0), .B(_auto_iopadmap_cc_313_execute_56321_23_), .Y(u0__abc_49347_n4373) );
  OR2X2 OR2X2_95 ( .A(_abc_55805_n240_bF_buf3), .B(sp_csc_3_), .Y(_abc_55805_n395) );
  OR2X2 OR2X2_950 ( .A(u0__abc_49347_n4304_bF_buf1), .B(mc_data_ir_23_), .Y(u0__abc_49347_n4374) );
  OR2X2 OR2X2_951 ( .A(u0_rst_r3_bF_buf4), .B(_auto_iopadmap_cc_313_execute_56321_24_), .Y(u0__abc_49347_n4376) );
  OR2X2 OR2X2_952 ( .A(u0__abc_49347_n4304_bF_buf0), .B(mc_data_ir_24_), .Y(u0__abc_49347_n4377) );
  OR2X2 OR2X2_953 ( .A(u0_rst_r3_bF_buf3), .B(_auto_iopadmap_cc_313_execute_56321_25_), .Y(u0__abc_49347_n4379) );
  OR2X2 OR2X2_954 ( .A(u0__abc_49347_n4304_bF_buf4), .B(mc_data_ir_25_), .Y(u0__abc_49347_n4380) );
  OR2X2 OR2X2_955 ( .A(u0_rst_r3_bF_buf2), .B(_auto_iopadmap_cc_313_execute_56321_26_), .Y(u0__abc_49347_n4382) );
  OR2X2 OR2X2_956 ( .A(u0__abc_49347_n4304_bF_buf3), .B(mc_data_ir_26_), .Y(u0__abc_49347_n4383) );
  OR2X2 OR2X2_957 ( .A(u0_rst_r3_bF_buf1), .B(_auto_iopadmap_cc_313_execute_56321_27_), .Y(u0__abc_49347_n4385) );
  OR2X2 OR2X2_958 ( .A(u0__abc_49347_n4304_bF_buf2), .B(mc_data_ir_27_), .Y(u0__abc_49347_n4386) );
  OR2X2 OR2X2_959 ( .A(u0_rst_r3_bF_buf0), .B(_auto_iopadmap_cc_313_execute_56321_28_), .Y(u0__abc_49347_n4388) );
  OR2X2 OR2X2_96 ( .A(lmr_sel_bF_buf3), .B(csc_3_), .Y(_abc_55805_n396) );
  OR2X2 OR2X2_960 ( .A(u0__abc_49347_n4304_bF_buf1), .B(mc_data_ir_28_), .Y(u0__abc_49347_n4389) );
  OR2X2 OR2X2_961 ( .A(u0_rst_r3_bF_buf4), .B(_auto_iopadmap_cc_313_execute_56321_29_), .Y(u0__abc_49347_n4391) );
  OR2X2 OR2X2_962 ( .A(u0__abc_49347_n4304_bF_buf0), .B(mc_data_ir_29_), .Y(u0__abc_49347_n4392) );
  OR2X2 OR2X2_963 ( .A(u0_rst_r3_bF_buf3), .B(_auto_iopadmap_cc_313_execute_56321_30_), .Y(u0__abc_49347_n4394) );
  OR2X2 OR2X2_964 ( .A(u0__abc_49347_n4304_bF_buf4), .B(mc_data_ir_30_), .Y(u0__abc_49347_n4395) );
  OR2X2 OR2X2_965 ( .A(u0_rst_r3_bF_buf2), .B(_auto_iopadmap_cc_313_execute_56321_31_), .Y(u0__abc_49347_n4397) );
  OR2X2 OR2X2_966 ( .A(u0__abc_49347_n4304_bF_buf3), .B(mc_data_ir_31_), .Y(u0__abc_49347_n4398) );
  OR2X2 OR2X2_967 ( .A(u0_wb_addr_r_6_), .B(u0_wb_addr_r_2_), .Y(u0__abc_49347_n4401) );
  OR2X2 OR2X2_968 ( .A(u0__abc_49347_n4401), .B(u0__abc_49347_n4400), .Y(u0__abc_49347_n4402) );
  OR2X2 OR2X2_969 ( .A(u0_wb_addr_r_5_), .B(u0_wb_addr_r_4_), .Y(u0__abc_49347_n4404) );
  OR2X2 OR2X2_97 ( .A(_abc_55805_n240_bF_buf2), .B(sp_csc_4_), .Y(_abc_55805_n398) );
  OR2X2 OR2X2_970 ( .A(u0__abc_49347_n4407), .B(u0_csc_mask_0_), .Y(u0__abc_49347_n4408) );
  OR2X2 OR2X2_971 ( .A(u0__abc_49347_n4409), .B(\wb_data_i[0] ), .Y(u0__abc_49347_n4410) );
  OR2X2 OR2X2_972 ( .A(u0__abc_49347_n4407), .B(u0_csc_mask_1_), .Y(u0__abc_49347_n4412) );
  OR2X2 OR2X2_973 ( .A(u0__abc_49347_n4409), .B(\wb_data_i[1] ), .Y(u0__abc_49347_n4413) );
  OR2X2 OR2X2_974 ( .A(u0__abc_49347_n4407), .B(u0_csc_mask_2_), .Y(u0__abc_49347_n4415) );
  OR2X2 OR2X2_975 ( .A(u0__abc_49347_n4409), .B(\wb_data_i[2] ), .Y(u0__abc_49347_n4416) );
  OR2X2 OR2X2_976 ( .A(u0__abc_49347_n4407), .B(u0_csc_mask_3_), .Y(u0__abc_49347_n4418) );
  OR2X2 OR2X2_977 ( .A(u0__abc_49347_n4409), .B(\wb_data_i[3] ), .Y(u0__abc_49347_n4419) );
  OR2X2 OR2X2_978 ( .A(u0__abc_49347_n4407), .B(u0_csc_mask_4_), .Y(u0__abc_49347_n4421) );
  OR2X2 OR2X2_979 ( .A(u0__abc_49347_n4409), .B(\wb_data_i[4] ), .Y(u0__abc_49347_n4422) );
  OR2X2 OR2X2_98 ( .A(lmr_sel_bF_buf2), .B(csc_4_), .Y(_abc_55805_n399) );
  OR2X2 OR2X2_980 ( .A(u0__abc_49347_n4407), .B(u0_csc_mask_5_), .Y(u0__abc_49347_n4424) );
  OR2X2 OR2X2_981 ( .A(u0__abc_49347_n4409), .B(\wb_data_i[5] ), .Y(u0__abc_49347_n4425) );
  OR2X2 OR2X2_982 ( .A(u0__abc_49347_n4407), .B(u0_csc_mask_6_), .Y(u0__abc_49347_n4427) );
  OR2X2 OR2X2_983 ( .A(u0__abc_49347_n4409), .B(\wb_data_i[6] ), .Y(u0__abc_49347_n4428) );
  OR2X2 OR2X2_984 ( .A(u0__abc_49347_n4407), .B(u0_csc_mask_7_), .Y(u0__abc_49347_n4430) );
  OR2X2 OR2X2_985 ( .A(u0__abc_49347_n4409), .B(\wb_data_i[7] ), .Y(u0__abc_49347_n4431) );
  OR2X2 OR2X2_986 ( .A(u0__abc_49347_n4407), .B(u0_csc_mask_8_), .Y(u0__abc_49347_n4433) );
  OR2X2 OR2X2_987 ( .A(u0__abc_49347_n4409), .B(\wb_data_i[8] ), .Y(u0__abc_49347_n4434) );
  OR2X2 OR2X2_988 ( .A(u0__abc_49347_n4407), .B(u0_csc_mask_9_), .Y(u0__abc_49347_n4436) );
  OR2X2 OR2X2_989 ( .A(u0__abc_49347_n4409), .B(\wb_data_i[9] ), .Y(u0__abc_49347_n4437) );
  OR2X2 OR2X2_99 ( .A(_abc_55805_n240_bF_buf1), .B(sp_csc_5_), .Y(_abc_55805_n401) );
  OR2X2 OR2X2_990 ( .A(u0__abc_49347_n4407), .B(u0_csc_mask_10_), .Y(u0__abc_49347_n4439) );
  OR2X2 OR2X2_991 ( .A(u0__abc_49347_n4409), .B(\wb_data_i[10] ), .Y(u0__abc_49347_n4440) );
  OR2X2 OR2X2_992 ( .A(u0__abc_49347_n4404), .B(u0_wb_addr_r_3_), .Y(u0__abc_49347_n4442) );
  OR2X2 OR2X2_993 ( .A(u0__abc_49347_n4402), .B(u0__abc_49347_n4442), .Y(u0__abc_49347_n4443) );
  OR2X2 OR2X2_994 ( .A(u0__abc_49347_n4444_bF_buf3), .B(_auto_iopadmap_cc_313_execute_56315), .Y(u0__abc_49347_n4445) );
  OR2X2 OR2X2_995 ( .A(u0__abc_49347_n4443_bF_buf2), .B(\wb_data_i[1] ), .Y(u0__abc_49347_n4446) );
  OR2X2 OR2X2_996 ( .A(u0__abc_49347_n4444_bF_buf2), .B(fs), .Y(u0__abc_49347_n4448) );
  OR2X2 OR2X2_997 ( .A(u0__abc_49347_n4443_bF_buf1), .B(\wb_data_i[2] ), .Y(u0__abc_49347_n4449) );
  OR2X2 OR2X2_998 ( .A(u0__abc_49347_n4444_bF_buf1), .B(u0_csr_3_), .Y(u0__abc_49347_n4451) );
  OR2X2 OR2X2_999 ( .A(u0__abc_49347_n4443_bF_buf0), .B(\wb_data_i[3] ), .Y(u0__abc_49347_n4452) );
endmodule
