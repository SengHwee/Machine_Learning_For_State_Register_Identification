module uart(clk, rst, rx, transmit, \tx_byte[0] , \tx_byte[1] , \tx_byte[2] , \tx_byte[3] , \tx_byte[4] , \tx_byte[5] , \tx_byte[6] , \tx_byte[7] , tx, received, \rx_byte[0] , \rx_byte[1] , \rx_byte[2] , \rx_byte[3] , \rx_byte[4] , \rx_byte[5] , \rx_byte[6] , \rx_byte[7] , is_receiving, is_transmitting, recv_error);
  wire _abc_2290_n144;
  wire _abc_2290_n145;
  wire _abc_2290_n146;
  wire _abc_2290_n147_1;
  wire _abc_2290_n150;
  wire _abc_2290_n152_1;
  wire _abc_2290_n153;
  wire _abc_2290_n155;
  wire _abc_2290_n156_1;
  wire _abc_2290_n157_1;
  wire _abc_2290_n158;
  wire _abc_2290_n159;
  wire _abc_2290_n160;
  wire _abc_2290_n161_1;
  wire _abc_2290_n162;
  wire _abc_2290_n163;
  wire _abc_2290_n164;
  wire _abc_2290_n165_1;
  wire _abc_2290_n166_1;
  wire _abc_2290_n167;
  wire _abc_2290_n168;
  wire _abc_2290_n169;
  wire _abc_2290_n170_1;
  wire _abc_2290_n171;
  wire _abc_2290_n172;
  wire _abc_2290_n173;
  wire _abc_2290_n174_1;
  wire _abc_2290_n175_1;
  wire _abc_2290_n176;
  wire _abc_2290_n177;
  wire _abc_2290_n178;
  wire _abc_2290_n179_1;
  wire _abc_2290_n180;
  wire _abc_2290_n181;
  wire _abc_2290_n182;
  wire _abc_2290_n183_1;
  wire _abc_2290_n184;
  wire _abc_2290_n185_1;
  wire _abc_2290_n186;
  wire _abc_2290_n187;
  wire _abc_2290_n188;
  wire _abc_2290_n189_1;
  wire _abc_2290_n190;
  wire _abc_2290_n191;
  wire _abc_2290_n192;
  wire _abc_2290_n193;
  wire _abc_2290_n194;
  wire _abc_2290_n195_1;
  wire _abc_2290_n196;
  wire _abc_2290_n197;
  wire _abc_2290_n198;
  wire _abc_2290_n199;
  wire _abc_2290_n200;
  wire _abc_2290_n201;
  wire _abc_2290_n202_1;
  wire _abc_2290_n203;
  wire _abc_2290_n204;
  wire _abc_2290_n205;
  wire _abc_2290_n206;
  wire _abc_2290_n207;
  wire _abc_2290_n208;
  wire _abc_2290_n209_1;
  wire _abc_2290_n210;
  wire _abc_2290_n211;
  wire _abc_2290_n212;
  wire _abc_2290_n213;
  wire _abc_2290_n214;
  wire _abc_2290_n215;
  wire _abc_2290_n216;
  wire _abc_2290_n217_1;
  wire _abc_2290_n218;
  wire _abc_2290_n219;
  wire _abc_2290_n220;
  wire _abc_2290_n221;
  wire _abc_2290_n222_1;
  wire _abc_2290_n223;
  wire _abc_2290_n224;
  wire _abc_2290_n225;
  wire _abc_2290_n226;
  wire _abc_2290_n227_1;
  wire _abc_2290_n228;
  wire _abc_2290_n229;
  wire _abc_2290_n230;
  wire _abc_2290_n231;
  wire _abc_2290_n232_1;
  wire _abc_2290_n233;
  wire _abc_2290_n234;
  wire _abc_2290_n235;
  wire _abc_2290_n236;
  wire _abc_2290_n237_1;
  wire _abc_2290_n238;
  wire _abc_2290_n239;
  wire _abc_2290_n240;
  wire _abc_2290_n241_1;
  wire _abc_2290_n242;
  wire _abc_2290_n243;
  wire _abc_2290_n244;
  wire _abc_2290_n245_1;
  wire _abc_2290_n246;
  wire _abc_2290_n247;
  wire _abc_2290_n248;
  wire _abc_2290_n249;
  wire _abc_2290_n250_1;
  wire _abc_2290_n251;
  wire _abc_2290_n252;
  wire _abc_2290_n253;
  wire _abc_2290_n254;
  wire _abc_2290_n255;
  wire _abc_2290_n256;
  wire _abc_2290_n257_1;
  wire _abc_2290_n258_1;
  wire _abc_2290_n259;
  wire _abc_2290_n260;
  wire _abc_2290_n261;
  wire _abc_2290_n262;
  wire _abc_2290_n263;
  wire _abc_2290_n264_1;
  wire _abc_2290_n265_1;
  wire _abc_2290_n266;
  wire _abc_2290_n267_1;
  wire _abc_2290_n268_1;
  wire _abc_2290_n269;
  wire _abc_2290_n270_1;
  wire _abc_2290_n271_1;
  wire _abc_2290_n272;
  wire _abc_2290_n273_1;
  wire _abc_2290_n274_1;
  wire _abc_2290_n275;
  wire _abc_2290_n276;
  wire _abc_2290_n277;
  wire _abc_2290_n278;
  wire _abc_2290_n279;
  wire _abc_2290_n280;
  wire _abc_2290_n281_1;
  wire _abc_2290_n282;
  wire _abc_2290_n283;
  wire _abc_2290_n284;
  wire _abc_2290_n285;
  wire _abc_2290_n287;
  wire _abc_2290_n288;
  wire _abc_2290_n289;
  wire _abc_2290_n290;
  wire _abc_2290_n291;
  wire _abc_2290_n292;
  wire _abc_2290_n294;
  wire _abc_2290_n295;
  wire _abc_2290_n296;
  wire _abc_2290_n297;
  wire _abc_2290_n298;
  wire _abc_2290_n299_1;
  wire _abc_2290_n301;
  wire _abc_2290_n302;
  wire _abc_2290_n303;
  wire _abc_2290_n304;
  wire _abc_2290_n305;
  wire _abc_2290_n306;
  wire _abc_2290_n308;
  wire _abc_2290_n309;
  wire _abc_2290_n310;
  wire _abc_2290_n311;
  wire _abc_2290_n312_1;
  wire _abc_2290_n313;
  wire _abc_2290_n315;
  wire _abc_2290_n316;
  wire _abc_2290_n317;
  wire _abc_2290_n318;
  wire _abc_2290_n319_1;
  wire _abc_2290_n320;
  wire _abc_2290_n322;
  wire _abc_2290_n323_1;
  wire _abc_2290_n324;
  wire _abc_2290_n325;
  wire _abc_2290_n326;
  wire _abc_2290_n327;
  wire _abc_2290_n328;
  wire _abc_2290_n330;
  wire _abc_2290_n331;
  wire _abc_2290_n332;
  wire _abc_2290_n334;
  wire _abc_2290_n335;
  wire _abc_2290_n336;
  wire _abc_2290_n337;
  wire _abc_2290_n338;
  wire _abc_2290_n340;
  wire _abc_2290_n341;
  wire _abc_2290_n342;
  wire _abc_2290_n343;
  wire _abc_2290_n344_1;
  wire _abc_2290_n345;
  wire _abc_2290_n346;
  wire _abc_2290_n347;
  wire _abc_2290_n348;
  wire _abc_2290_n349;
  wire _abc_2290_n351;
  wire _abc_2290_n352_1;
  wire _abc_2290_n353;
  wire _abc_2290_n354;
  wire _abc_2290_n355;
  wire _abc_2290_n356;
  wire _abc_2290_n357_1;
  wire _abc_2290_n358;
  wire _abc_2290_n360;
  wire _abc_2290_n361;
  wire _abc_2290_n362;
  wire _abc_2290_n364;
  wire _abc_2290_n367;
  wire _abc_2290_n369;
  wire _abc_2290_n370;
  wire _abc_2290_n372;
  wire _abc_2290_n373;
  wire _abc_2290_n374_1;
  wire _abc_2290_n375;
  wire _abc_2290_n376;
  wire _abc_2290_n377;
  wire _abc_2290_n378;
  wire _abc_2290_n379;
  wire _abc_2290_n382_1;
  wire _abc_2290_n383;
  wire _abc_2290_n384;
  wire _abc_2290_n385;
  wire _abc_2290_n387;
  wire _abc_2290_n388;
  wire _abc_2290_n390;
  wire _abc_2290_n391;
  wire _abc_2290_n392;
  wire _abc_2290_n393;
  wire _abc_2290_n394;
  wire _abc_2290_n396;
  wire _abc_2290_n397;
  wire _abc_2290_n398_1;
  wire _abc_2290_n399;
  wire _abc_2290_n400;
  wire _abc_2290_n401;
  wire _abc_2290_n402;
  wire _abc_2290_n403;
  wire _abc_2290_n404_1;
  wire _abc_2290_n405;
  wire _abc_2290_n406;
  wire _abc_2290_n407;
  wire _abc_2290_n408;
  wire _abc_2290_n409;
  wire _abc_2290_n410_1;
  wire _abc_2290_n411;
  wire _abc_2290_n412;
  wire _abc_2290_n413;
  wire _abc_2290_n414;
  wire _abc_2290_n415;
  wire _abc_2290_n416;
  wire _abc_2290_n417;
  wire _abc_2290_n418;
  wire _abc_2290_n419;
  wire _abc_2290_n420;
  wire _abc_2290_n421;
  wire _abc_2290_n422;
  wire _abc_2290_n423_1;
  wire _abc_2290_n424;
  wire _abc_2290_n425_1;
  wire _abc_2290_n426;
  wire _abc_2290_n427_1;
  wire _abc_2290_n428_1;
  wire _abc_2290_n429;
  wire _abc_2290_n430;
  wire _abc_2290_n431;
  wire _abc_2290_n432;
  wire _abc_2290_n433;
  wire _abc_2290_n434;
  wire _abc_2290_n435;
  wire _abc_2290_n436;
  wire _abc_2290_n437;
  wire _abc_2290_n438;
  wire _abc_2290_n439;
  wire _abc_2290_n440;
  wire _abc_2290_n441_1;
  wire _abc_2290_n442;
  wire _abc_2290_n443;
  wire _abc_2290_n444;
  wire _abc_2290_n445;
  wire _abc_2290_n446;
  wire _abc_2290_n447;
  wire _abc_2290_n448;
  wire _abc_2290_n449_1;
  wire _abc_2290_n450;
  wire _abc_2290_n451;
  wire _abc_2290_n452;
  wire _abc_2290_n453;
  wire _abc_2290_n454;
  wire _abc_2290_n455;
  wire _abc_2290_n456;
  wire _abc_2290_n457;
  wire _abc_2290_n458;
  wire _abc_2290_n459_1;
  wire _abc_2290_n460;
  wire _abc_2290_n461;
  wire _abc_2290_n462;
  wire _abc_2290_n463;
  wire _abc_2290_n464_1;
  wire _abc_2290_n465;
  wire _abc_2290_n466;
  wire _abc_2290_n467;
  wire _abc_2290_n468;
  wire _abc_2290_n469_1;
  wire _abc_2290_n470;
  wire _abc_2290_n471;
  wire _abc_2290_n473_1;
  wire _abc_2290_n474;
  wire _abc_2290_n475;
  wire _abc_2290_n476;
  wire _abc_2290_n477_1;
  wire _abc_2290_n478;
  wire _abc_2290_n479_1;
  wire _abc_2290_n480;
  wire _abc_2290_n481;
  wire _abc_2290_n483;
  wire _abc_2290_n484_1;
  wire _abc_2290_n485;
  wire _abc_2290_n486;
  wire _abc_2290_n487_1;
  wire _abc_2290_n488;
  wire _abc_2290_n489_1;
  wire _abc_2290_n490;
  wire _abc_2290_n491_1;
  wire _abc_2290_n492;
  wire _abc_2290_n493_1;
  wire _abc_2290_n494_1;
  wire _abc_2290_n495;
  wire _abc_2290_n496_1;
  wire _abc_2290_n497;
  wire _abc_2290_n498_1;
  wire _abc_2290_n499;
  wire _abc_2290_n500_1;
  wire _abc_2290_n501;
  wire _abc_2290_n502_1;
  wire _abc_2290_n503;
  wire _abc_2290_n504;
  wire _abc_2290_n505_1;
  wire _abc_2290_n506;
  wire _abc_2290_n507_1;
  wire _abc_2290_n508;
  wire _abc_2290_n509;
  wire _abc_2290_n510_1;
  wire _abc_2290_n511;
  wire _abc_2290_n512_1;
  wire _abc_2290_n513;
  wire _abc_2290_n514_1;
  wire _abc_2290_n515;
  wire _abc_2290_n516_1;
  wire _abc_2290_n517;
  wire _abc_2290_n518_1;
  wire _abc_2290_n519;
  wire _abc_2290_n520_1;
  wire _abc_2290_n521;
  wire _abc_2290_n522_1;
  wire _abc_2290_n523;
  wire _abc_2290_n524_1;
  wire _abc_2290_n525_1;
  wire _abc_2290_n526_1;
  wire _abc_2290_n527;
  wire _abc_2290_n528_1;
  wire _abc_2290_n529_1;
  wire _abc_2290_n530;
  wire _abc_2290_n531_1;
  wire _abc_2290_n532_1;
  wire _abc_2290_n533;
  wire _abc_2290_n534_1;
  wire _abc_2290_n535_1;
  wire _abc_2290_n536;
  wire _abc_2290_n537_1;
  wire _abc_2290_n538_1;
  wire _abc_2290_n539;
  wire _abc_2290_n540_1;
  wire _abc_2290_n541_1;
  wire _abc_2290_n542;
  wire _abc_2290_n543_1;
  wire _abc_2290_n544_1;
  wire _abc_2290_n545;
  wire _abc_2290_n546_1;
  wire _abc_2290_n547;
  wire _abc_2290_n548_1;
  wire _abc_2290_n548_1_bF_buf0;
  wire _abc_2290_n548_1_bF_buf1;
  wire _abc_2290_n548_1_bF_buf2;
  wire _abc_2290_n548_1_bF_buf3;
  wire _abc_2290_n549;
  wire _abc_2290_n551;
  wire _abc_2290_n552;
  wire _abc_2290_n553;
  wire _abc_2290_n555;
  wire _abc_2290_n557;
  wire _abc_2290_n559;
  wire _abc_2290_n560;
  wire _abc_2290_n561;
  wire _abc_2290_n562;
  wire _abc_2290_n563;
  wire _abc_2290_n564;
  wire _abc_2290_n565;
  wire _abc_2290_n566;
  wire _abc_2290_n567;
  wire _abc_2290_n568;
  wire _abc_2290_n569;
  wire _abc_2290_n570;
  wire _abc_2290_n571;
  wire _abc_2290_n572;
  wire _abc_2290_n573;
  wire _abc_2290_n574;
  wire _abc_2290_n575;
  wire _abc_2290_n576;
  wire _abc_2290_n577;
  wire _abc_2290_n578;
  wire _abc_2290_n579;
  wire _abc_2290_n580;
  wire _abc_2290_n582;
  wire _abc_2290_n583;
  wire _abc_2290_n584;
  wire _abc_2290_n585;
  wire _abc_2290_n586;
  wire _abc_2290_n587;
  wire _abc_2290_n588;
  wire _abc_2290_n589;
  wire _abc_2290_n591;
  wire _abc_2290_n592;
  wire _abc_2290_n593;
  wire _abc_2290_n594;
  wire _abc_2290_n595;
  wire _abc_2290_n597;
  wire _abc_2290_n598;
  wire _abc_2290_n599;
  wire _abc_2290_n600;
  wire _abc_2290_n601;
  wire _abc_2290_n603;
  wire _abc_2290_n604;
  wire _abc_2290_n605;
  wire _abc_2290_n606;
  wire _abc_2290_n607;
  wire _abc_2290_n608;
  wire _abc_2290_n609;
  wire _abc_2290_n610;
  wire _abc_2290_n611;
  wire _abc_2290_n613;
  wire _abc_2290_n614;
  wire _abc_2290_n615;
  wire _abc_2290_n616;
  wire _abc_2290_n617;
  wire _abc_2290_n618;
  wire _abc_2290_n619;
  wire _abc_2290_n620;
  wire _abc_2290_n621;
  wire _abc_2290_n623;
  wire _abc_2290_n624;
  wire _abc_2290_n625;
  wire _abc_2290_n626;
  wire _abc_2290_n627;
  wire _abc_2290_n630;
  wire _abc_2290_n631;
  wire _abc_2290_n632;
  wire _abc_2290_n634;
  wire _abc_2290_n635;
  wire _abc_2290_n636;
  wire _abc_2290_n637;
  wire _abc_2290_n638;
  wire _abc_2290_n640;
  wire _abc_2290_n641;
  wire _abc_2290_n643;
  wire _abc_2290_n644;
  wire _abc_2290_n645;
  wire _abc_2290_n647;
  wire _abc_2290_n649;
  wire _abc_2290_n650;
  wire _abc_2290_n652;
  wire _abc_2290_n654;
  wire _abc_2290_n656;
  wire _abc_2290_n658;
  wire _abc_2290_n661;
  wire _abc_2290_n662;
  wire _abc_2290_n663;
  wire _abc_2290_n665;
  wire _abc_2290_n666;
  wire _abc_2290_n667;
  wire _abc_2290_n668;
  wire _abc_2290_n670;
  wire _abc_2290_n671;
  wire _abc_2290_n672;
  wire _abc_2290_n674;
  wire _abc_2290_n675;
  wire _abc_2290_n677;
  wire _abc_2290_n679;
  wire _abc_2290_n681;
  wire _abc_2290_n683;
  wire _abc_2290_n684;
  wire _abc_2290_n686;
  wire _abc_2290_n688;
  wire _abc_2290_n689;
  wire _abc_2290_n691;
  wire _abc_2290_n692;
  wire _abc_2290_n693;
  wire _abc_2290_n694;
  wire _abc_2290_n696;
  wire _abc_2290_n697;
  wire _abc_2290_n698;
  wire _abc_2290_n699;
  wire _abc_2290_n701;
  wire _abc_2290_n702;
  wire _abc_2290_n703;
  wire _abc_2290_n704;
  wire _abc_2290_n706;
  wire _abc_2290_n707;
  wire _abc_2290_n708;
  wire _abc_2290_n709;
  wire _abc_2290_n711;
  wire _abc_2290_n712;
  wire _abc_2290_n713;
  wire _abc_2290_n714;
  wire _abc_2290_n716;
  wire _abc_2290_n717;
  wire _abc_2290_n718;
  wire _abc_2290_n719;
  wire _abc_2290_n721;
  wire _abc_2290_n722;
  wire _abc_2290_n723;
  wire _abc_2290_n724;
  wire _abc_2290_n726;
  wire _abc_2290_n727;
  wire _abc_2290_n728;
  input clk;
  wire clk_bF_buf0;
  wire clk_bF_buf1;
  wire clk_bF_buf2;
  wire clk_bF_buf3;
  wire clk_bF_buf4;
  wire clk_bF_buf5;
  wire clk_bF_buf6;
  wire clk_bF_buf7;
  output is_receiving;
  output is_transmitting;
  output received;
  output recv_error;
  wire recv_state_0_;
  wire recv_state_0__FF_INPUT;
  wire recv_state_1_;
  wire recv_state_1__FF_INPUT;
  wire recv_state_2_;
  wire recv_state_2__FF_INPUT;
  input rst;
  input rx;
  wire rx_bits_remaining_0_;
  wire rx_bits_remaining_0__FF_INPUT;
  wire rx_bits_remaining_1_;
  wire rx_bits_remaining_1__FF_INPUT;
  wire rx_bits_remaining_2_;
  wire rx_bits_remaining_2__FF_INPUT;
  wire rx_bits_remaining_3_;
  wire rx_bits_remaining_3__FF_INPUT;
  output \rx_byte[0] ;
  output \rx_byte[1] ;
  output \rx_byte[2] ;
  output \rx_byte[3] ;
  output \rx_byte[4] ;
  output \rx_byte[5] ;
  output \rx_byte[6] ;
  output \rx_byte[7] ;
  wire rx_clk_divider_0_;
  wire rx_clk_divider_0__FF_INPUT;
  wire rx_clk_divider_10_;
  wire rx_clk_divider_10__FF_INPUT;
  wire rx_clk_divider_1_;
  wire rx_clk_divider_1__FF_INPUT;
  wire rx_clk_divider_2_;
  wire rx_clk_divider_2__FF_INPUT;
  wire rx_clk_divider_3_;
  wire rx_clk_divider_3__FF_INPUT;
  wire rx_clk_divider_4_;
  wire rx_clk_divider_4__FF_INPUT;
  wire rx_clk_divider_5_;
  wire rx_clk_divider_5__FF_INPUT;
  wire rx_clk_divider_6_;
  wire rx_clk_divider_6__FF_INPUT;
  wire rx_clk_divider_7_;
  wire rx_clk_divider_7__FF_INPUT;
  wire rx_clk_divider_8_;
  wire rx_clk_divider_8__FF_INPUT;
  wire rx_clk_divider_9_;
  wire rx_clk_divider_9__FF_INPUT;
  wire rx_countdown_0_;
  wire rx_countdown_0__FF_INPUT;
  wire rx_countdown_1_;
  wire rx_countdown_1__FF_INPUT;
  wire rx_countdown_2_;
  wire rx_countdown_2__FF_INPUT;
  wire rx_countdown_3_;
  wire rx_countdown_3__FF_INPUT;
  wire rx_countdown_4_;
  wire rx_countdown_4__FF_INPUT;
  wire rx_countdown_5_;
  wire rx_countdown_5__FF_INPUT;
  wire rx_data_0__FF_INPUT;
  wire rx_data_1__FF_INPUT;
  wire rx_data_2__FF_INPUT;
  wire rx_data_3__FF_INPUT;
  wire rx_data_4__FF_INPUT;
  wire rx_data_5__FF_INPUT;
  wire rx_data_6__FF_INPUT;
  wire rx_data_7__FF_INPUT;
  input transmit;
  output tx;
  wire tx_bits_remaining_0_;
  wire tx_bits_remaining_0__FF_INPUT;
  wire tx_bits_remaining_1_;
  wire tx_bits_remaining_1__FF_INPUT;
  wire tx_bits_remaining_2_;
  wire tx_bits_remaining_2__FF_INPUT;
  wire tx_bits_remaining_3_;
  wire tx_bits_remaining_3__FF_INPUT;
  input \tx_byte[0] ;
  input \tx_byte[1] ;
  input \tx_byte[2] ;
  input \tx_byte[3] ;
  input \tx_byte[4] ;
  input \tx_byte[5] ;
  input \tx_byte[6] ;
  input \tx_byte[7] ;
  wire tx_clk_divider_0_;
  wire tx_clk_divider_0__FF_INPUT;
  wire tx_clk_divider_10_;
  wire tx_clk_divider_10__FF_INPUT;
  wire tx_clk_divider_1_;
  wire tx_clk_divider_1__FF_INPUT;
  wire tx_clk_divider_2_;
  wire tx_clk_divider_2__FF_INPUT;
  wire tx_clk_divider_3_;
  wire tx_clk_divider_3__FF_INPUT;
  wire tx_clk_divider_4_;
  wire tx_clk_divider_4__FF_INPUT;
  wire tx_clk_divider_5_;
  wire tx_clk_divider_5__FF_INPUT;
  wire tx_clk_divider_6_;
  wire tx_clk_divider_6__FF_INPUT;
  wire tx_clk_divider_7_;
  wire tx_clk_divider_7__FF_INPUT;
  wire tx_clk_divider_8_;
  wire tx_clk_divider_8__FF_INPUT;
  wire tx_clk_divider_9_;
  wire tx_clk_divider_9__FF_INPUT;
  wire tx_countdown_0_;
  wire tx_countdown_0__FF_INPUT;
  wire tx_countdown_1_;
  wire tx_countdown_1__FF_INPUT;
  wire tx_countdown_2_;
  wire tx_countdown_2__FF_INPUT;
  wire tx_countdown_3_;
  wire tx_countdown_3__FF_INPUT;
  wire tx_countdown_4_;
  wire tx_countdown_4__FF_INPUT;
  wire tx_countdown_5_;
  wire tx_countdown_5__FF_INPUT;
  wire tx_data_0_;
  wire tx_data_0__FF_INPUT;
  wire tx_data_1_;
  wire tx_data_1__FF_INPUT;
  wire tx_data_2_;
  wire tx_data_2__FF_INPUT;
  wire tx_data_3_;
  wire tx_data_3__FF_INPUT;
  wire tx_data_4_;
  wire tx_data_4__FF_INPUT;
  wire tx_data_5_;
  wire tx_data_5__FF_INPUT;
  wire tx_data_6_;
  wire tx_data_6__FF_INPUT;
  wire tx_data_7_;
  wire tx_data_7__FF_INPUT;
  wire tx_out;
  wire tx_out_FF_INPUT;
  wire tx_state_0_;
  wire tx_state_0__FF_INPUT;
  wire tx_state_1_;
  wire tx_state_1__FF_INPUT;
  AND2X2 AND2X2_1 ( .A(_abc_2290_n144), .B(_abc_2290_n145), .Y(_abc_2290_n146) );
  AND2X2 AND2X2_10 ( .A(_abc_2290_n162), .B(_abc_2290_n165_1), .Y(_abc_2290_n166_1) );
  AND2X2 AND2X2_100 ( .A(_abc_2290_n158), .B(tx_bits_remaining_3_), .Y(_abc_2290_n353) );
  AND2X2 AND2X2_101 ( .A(_abc_2290_n352_1), .B(_abc_2290_n353), .Y(_abc_2290_n354) );
  AND2X2 AND2X2_102 ( .A(_abc_2290_n355), .B(_abc_2290_n158), .Y(_abc_2290_n356) );
  AND2X2 AND2X2_103 ( .A(_abc_2290_n357_1), .B(tx_bits_remaining_2_), .Y(_abc_2290_n358) );
  AND2X2 AND2X2_104 ( .A(_abc_2290_n352_1), .B(_abc_2290_n158), .Y(_abc_2290_n360) );
  AND2X2 AND2X2_105 ( .A(_abc_2290_n361), .B(tx_bits_remaining_3_), .Y(_abc_2290_n362) );
  AND2X2 AND2X2_106 ( .A(_abc_2290_n243), .B(_abc_2290_n364), .Y(tx_countdown_0__FF_INPUT) );
  AND2X2 AND2X2_107 ( .A(_abc_2290_n258_1), .B(_abc_2290_n364), .Y(tx_countdown_1__FF_INPUT) );
  AND2X2 AND2X2_108 ( .A(_abc_2290_n283), .B(_abc_2290_n345), .Y(_abc_2290_n369) );
  AND2X2 AND2X2_109 ( .A(_abc_2290_n370), .B(_abc_2290_n331), .Y(tx_countdown_3__FF_INPUT) );
  AND2X2 AND2X2_11 ( .A(_abc_2290_n167), .B(_abc_2290_n168), .Y(_abc_2290_n169) );
  AND2X2 AND2X2_110 ( .A(_abc_2290_n197), .B(_abc_2290_n208), .Y(_abc_2290_n372) );
  AND2X2 AND2X2_111 ( .A(_abc_2290_n372), .B(_abc_2290_n206), .Y(_abc_2290_n373) );
  AND2X2 AND2X2_112 ( .A(_abc_2290_n373), .B(_abc_2290_n218), .Y(_abc_2290_n374_1) );
  AND2X2 AND2X2_113 ( .A(_abc_2290_n374_1), .B(_abc_2290_n213), .Y(_abc_2290_n375) );
  AND2X2 AND2X2_114 ( .A(_abc_2290_n375), .B(_abc_2290_n212), .Y(_abc_2290_n376) );
  AND2X2 AND2X2_115 ( .A(_abc_2290_n377), .B(tx_countdown_4_), .Y(_abc_2290_n378) );
  AND2X2 AND2X2_116 ( .A(_abc_2290_n379), .B(_abc_2290_n364), .Y(tx_countdown_4__FF_INPUT) );
  AND2X2 AND2X2_117 ( .A(_abc_2290_n228), .B(_abc_2290_n364), .Y(tx_countdown_5__FF_INPUT) );
  AND2X2 AND2X2_118 ( .A(_abc_2290_n345), .B(_abc_2290_n268_1), .Y(_abc_2290_n382_1) );
  AND2X2 AND2X2_119 ( .A(_abc_2290_n382_1), .B(_abc_2290_n155), .Y(_abc_2290_n383) );
  AND2X2 AND2X2_12 ( .A(_abc_2290_n166_1), .B(_abc_2290_n169), .Y(_abc_2290_n170_1) );
  AND2X2 AND2X2_120 ( .A(_abc_2290_n384), .B(_abc_2290_n157_1), .Y(_abc_2290_n385) );
  AND2X2 AND2X2_121 ( .A(_abc_2290_n387), .B(_abc_2290_n388), .Y(tx_state_1__FF_INPUT) );
  AND2X2 AND2X2_122 ( .A(_abc_2290_n391), .B(_abc_2290_n158), .Y(_abc_2290_n392) );
  AND2X2 AND2X2_123 ( .A(_abc_2290_n392), .B(_abc_2290_n390), .Y(_abc_2290_n393) );
  AND2X2 AND2X2_124 ( .A(_abc_2290_n280), .B(tx), .Y(_abc_2290_n394) );
  AND2X2 AND2X2_125 ( .A(_abc_2290_n397), .B(_abc_2290_n398_1), .Y(_abc_2290_n399) );
  AND2X2 AND2X2_126 ( .A(_abc_2290_n400), .B(_abc_2290_n401), .Y(_abc_2290_n402) );
  AND2X2 AND2X2_127 ( .A(_abc_2290_n399), .B(_abc_2290_n402), .Y(_abc_2290_n403) );
  AND2X2 AND2X2_128 ( .A(_abc_2290_n404_1), .B(_abc_2290_n405), .Y(_abc_2290_n406) );
  AND2X2 AND2X2_129 ( .A(_abc_2290_n407), .B(_abc_2290_n408), .Y(_abc_2290_n409) );
  AND2X2 AND2X2_13 ( .A(_abc_2290_n170_1), .B(_abc_2290_n172), .Y(_abc_2290_n173) );
  AND2X2 AND2X2_130 ( .A(_abc_2290_n406), .B(_abc_2290_n409), .Y(_abc_2290_n410_1) );
  AND2X2 AND2X2_131 ( .A(_abc_2290_n403), .B(_abc_2290_n410_1), .Y(_abc_2290_n411) );
  AND2X2 AND2X2_132 ( .A(_abc_2290_n412), .B(_abc_2290_n413), .Y(_abc_2290_n414) );
  AND2X2 AND2X2_133 ( .A(_abc_2290_n411), .B(_abc_2290_n414), .Y(_abc_2290_n415) );
  AND2X2 AND2X2_134 ( .A(_abc_2290_n426), .B(_abc_2290_n416), .Y(_abc_2290_n427_1) );
  AND2X2 AND2X2_135 ( .A(_abc_2290_n431), .B(_abc_2290_n423_1), .Y(_abc_2290_n432) );
  AND2X2 AND2X2_136 ( .A(_abc_2290_n403), .B(_abc_2290_n406), .Y(_abc_2290_n433) );
  AND2X2 AND2X2_137 ( .A(_abc_2290_n434), .B(_abc_2290_n429), .Y(_abc_2290_n435) );
  AND2X2 AND2X2_138 ( .A(_abc_2290_n403), .B(_abc_2290_n405), .Y(_abc_2290_n436) );
  AND2X2 AND2X2_139 ( .A(_abc_2290_n437), .B(_abc_2290_n428_1), .Y(_abc_2290_n438) );
  AND2X2 AND2X2_14 ( .A(_abc_2290_n173), .B(_abc_2290_n159), .Y(_abc_2290_n174_1) );
  AND2X2 AND2X2_140 ( .A(_abc_2290_n401), .B(_abc_2290_n412), .Y(_abc_2290_n440) );
  AND2X2 AND2X2_141 ( .A(_abc_2290_n440), .B(_abc_2290_n439), .Y(_abc_2290_n441_1) );
  AND2X2 AND2X2_142 ( .A(_abc_2290_n405), .B(rx_clk_divider_0_), .Y(_abc_2290_n442) );
  AND2X2 AND2X2_143 ( .A(_abc_2290_n399), .B(_abc_2290_n442), .Y(_abc_2290_n443) );
  AND2X2 AND2X2_144 ( .A(_abc_2290_n441_1), .B(_abc_2290_n443), .Y(_abc_2290_n444) );
  AND2X2 AND2X2_145 ( .A(_abc_2290_n438), .B(_abc_2290_n444), .Y(_abc_2290_n445) );
  AND2X2 AND2X2_146 ( .A(_abc_2290_n445), .B(_abc_2290_n435), .Y(_abc_2290_n446) );
  AND2X2 AND2X2_147 ( .A(_abc_2290_n446), .B(_abc_2290_n432), .Y(_abc_2290_n447) );
  AND2X2 AND2X2_148 ( .A(_abc_2290_n447), .B(_abc_2290_n427_1), .Y(_abc_2290_n448) );
  AND2X2 AND2X2_149 ( .A(_abc_2290_n448), .B(_abc_2290_n396), .Y(_abc_2290_n450) );
  AND2X2 AND2X2_15 ( .A(_abc_2290_n178), .B(tx_clk_divider_8_), .Y(_abc_2290_n179_1) );
  AND2X2 AND2X2_150 ( .A(_abc_2290_n451), .B(_abc_2290_n449_1), .Y(_abc_2290_n452) );
  AND2X2 AND2X2_151 ( .A(_abc_2290_n156_1), .B(recv_state_2_), .Y(_abc_2290_n454) );
  AND2X2 AND2X2_152 ( .A(_abc_2290_n454), .B(_abc_2290_n144), .Y(_abc_2290_n455) );
  AND2X2 AND2X2_153 ( .A(_abc_2290_n156_1), .B(recv_state_0_), .Y(_abc_2290_n456) );
  AND2X2 AND2X2_154 ( .A(_abc_2290_n456), .B(recv_state_1_), .Y(_abc_2290_n457) );
  AND2X2 AND2X2_155 ( .A(is_receiving), .B(_abc_2290_n156_1), .Y(_abc_2290_n459_1) );
  AND2X2 AND2X2_156 ( .A(_abc_2290_n460), .B(rx), .Y(_abc_2290_n461) );
  AND2X2 AND2X2_157 ( .A(_abc_2290_n156_1), .B(recv_state_1_), .Y(_abc_2290_n462) );
  AND2X2 AND2X2_158 ( .A(_abc_2290_n146), .B(_abc_2290_n462), .Y(_abc_2290_n463) );
  AND2X2 AND2X2_159 ( .A(_abc_2290_n456), .B(_abc_2290_n152_1), .Y(_abc_2290_n465) );
  AND2X2 AND2X2_16 ( .A(_abc_2290_n170_1), .B(_abc_2290_n183_1), .Y(_abc_2290_n184) );
  AND2X2 AND2X2_160 ( .A(_abc_2290_n465), .B(_abc_2290_n145), .Y(_abc_2290_n466) );
  AND2X2 AND2X2_161 ( .A(_abc_2290_n467), .B(_abc_2290_n464_1), .Y(_abc_2290_n468) );
  AND2X2 AND2X2_162 ( .A(_abc_2290_n453), .B(_abc_2290_n471), .Y(rx_countdown_0__FF_INPUT) );
  AND2X2 AND2X2_163 ( .A(_abc_2290_n460), .B(_abc_2290_n473_1), .Y(_abc_2290_n474) );
  AND2X2 AND2X2_164 ( .A(_abc_2290_n451), .B(rx_countdown_1_), .Y(_abc_2290_n475) );
  AND2X2 AND2X2_165 ( .A(_abc_2290_n450), .B(_abc_2290_n476), .Y(_abc_2290_n477_1) );
  AND2X2 AND2X2_166 ( .A(recv_error), .B(_abc_2290_n156_1), .Y(_abc_2290_n479_1) );
  AND2X2 AND2X2_167 ( .A(_abc_2290_n478), .B(_abc_2290_n480), .Y(_abc_2290_n481) );
  AND2X2 AND2X2_168 ( .A(_abc_2290_n484_1), .B(_abc_2290_n483), .Y(_abc_2290_n485) );
  AND2X2 AND2X2_169 ( .A(_abc_2290_n427_1), .B(_abc_2290_n485), .Y(_abc_2290_n486) );
  AND2X2 AND2X2_17 ( .A(_abc_2290_n185_1), .B(_abc_2290_n178), .Y(_abc_2290_n186) );
  AND2X2 AND2X2_170 ( .A(_abc_2290_n488), .B(_abc_2290_n487_1), .Y(_abc_2290_n489_1) );
  AND2X2 AND2X2_171 ( .A(_abc_2290_n401), .B(rx_clk_divider_0_), .Y(_abc_2290_n490) );
  AND2X2 AND2X2_172 ( .A(_abc_2290_n490), .B(_abc_2290_n398_1), .Y(_abc_2290_n491_1) );
  AND2X2 AND2X2_173 ( .A(_abc_2290_n491_1), .B(_abc_2290_n397), .Y(_abc_2290_n492) );
  AND2X2 AND2X2_174 ( .A(_abc_2290_n489_1), .B(_abc_2290_n492), .Y(_abc_2290_n493_1) );
  AND2X2 AND2X2_175 ( .A(_abc_2290_n438), .B(_abc_2290_n493_1), .Y(_abc_2290_n494_1) );
  AND2X2 AND2X2_176 ( .A(_abc_2290_n495), .B(_abc_2290_n424), .Y(_abc_2290_n496_1) );
  AND2X2 AND2X2_177 ( .A(_abc_2290_n496_1), .B(_abc_2290_n435), .Y(_abc_2290_n497) );
  AND2X2 AND2X2_178 ( .A(_abc_2290_n497), .B(_abc_2290_n494_1), .Y(_abc_2290_n498_1) );
  AND2X2 AND2X2_179 ( .A(_abc_2290_n498_1), .B(_abc_2290_n432), .Y(_abc_2290_n499) );
  AND2X2 AND2X2_18 ( .A(_abc_2290_n166_1), .B(_abc_2290_n168), .Y(_abc_2290_n188) );
  AND2X2 AND2X2_180 ( .A(_abc_2290_n499), .B(_abc_2290_n486), .Y(_abc_2290_n500_1) );
  AND2X2 AND2X2_181 ( .A(_abc_2290_n396), .B(_abc_2290_n476), .Y(_abc_2290_n502_1) );
  AND2X2 AND2X2_182 ( .A(_abc_2290_n502_1), .B(_abc_2290_n501), .Y(_abc_2290_n503) );
  AND2X2 AND2X2_183 ( .A(_abc_2290_n504), .B(rx_countdown_2_), .Y(_abc_2290_n505_1) );
  AND2X2 AND2X2_184 ( .A(_abc_2290_n500_1), .B(_abc_2290_n506), .Y(_abc_2290_n507_1) );
  AND2X2 AND2X2_185 ( .A(_abc_2290_n508), .B(_abc_2290_n509), .Y(_abc_2290_n510_1) );
  AND2X2 AND2X2_186 ( .A(_abc_2290_n511), .B(_abc_2290_n471), .Y(_abc_2290_n512_1) );
  AND2X2 AND2X2_187 ( .A(_abc_2290_n452), .B(_abc_2290_n476), .Y(_abc_2290_n513) );
  AND2X2 AND2X2_188 ( .A(_abc_2290_n503), .B(_abc_2290_n515), .Y(_abc_2290_n516_1) );
  AND2X2 AND2X2_189 ( .A(_abc_2290_n516_1), .B(_abc_2290_n514_1), .Y(_abc_2290_n517) );
  AND2X2 AND2X2_19 ( .A(_abc_2290_n189_1), .B(_abc_2290_n187), .Y(_abc_2290_n190) );
  AND2X2 AND2X2_190 ( .A(_abc_2290_n518_1), .B(rx_countdown_5_), .Y(_abc_2290_n519) );
  AND2X2 AND2X2_191 ( .A(_abc_2290_n517), .B(_abc_2290_n520_1), .Y(_abc_2290_n521) );
  AND2X2 AND2X2_192 ( .A(_abc_2290_n500_1), .B(_abc_2290_n522_1), .Y(_abc_2290_n523) );
  AND2X2 AND2X2_193 ( .A(_abc_2290_n524_1), .B(_abc_2290_n525_1), .Y(_abc_2290_n526_1) );
  AND2X2 AND2X2_194 ( .A(_abc_2290_n527), .B(rx_countdown_4_), .Y(_abc_2290_n528_1) );
  AND2X2 AND2X2_195 ( .A(_abc_2290_n500_1), .B(_abc_2290_n529_1), .Y(_abc_2290_n530) );
  AND2X2 AND2X2_196 ( .A(_abc_2290_n531_1), .B(_abc_2290_n532_1), .Y(_abc_2290_n533) );
  AND2X2 AND2X2_197 ( .A(_abc_2290_n526_1), .B(_abc_2290_n533), .Y(_abc_2290_n534_1) );
  AND2X2 AND2X2_198 ( .A(_abc_2290_n536), .B(_abc_2290_n537_1), .Y(_abc_2290_n538_1) );
  AND2X2 AND2X2_199 ( .A(_abc_2290_n500_1), .B(_abc_2290_n538_1), .Y(_abc_2290_n539) );
  AND2X2 AND2X2_2 ( .A(recv_state_1_), .B(recv_state_2_), .Y(_abc_2290_n150) );
  AND2X2 AND2X2_20 ( .A(_abc_2290_n164), .B(tx_clk_divider_0_), .Y(_abc_2290_n191) );
  AND2X2 AND2X2_200 ( .A(_abc_2290_n540_1), .B(_abc_2290_n541_1), .Y(_abc_2290_n542) );
  AND2X2 AND2X2_201 ( .A(_abc_2290_n510_1), .B(_abc_2290_n542), .Y(_abc_2290_n543_1) );
  AND2X2 AND2X2_202 ( .A(_abc_2290_n534_1), .B(_abc_2290_n543_1), .Y(_abc_2290_n544_1) );
  AND2X2 AND2X2_203 ( .A(_abc_2290_n544_1), .B(_abc_2290_n513), .Y(_abc_2290_n545) );
  AND2X2 AND2X2_204 ( .A(_abc_2290_n545), .B(_abc_2290_n473_1), .Y(_abc_2290_n546_1) );
  AND2X2 AND2X2_205 ( .A(_abc_2290_n546_1), .B(_abc_2290_n466), .Y(_abc_2290_n547) );
  AND2X2 AND2X2_206 ( .A(_abc_2290_n545), .B(_abc_2290_n463), .Y(_abc_2290_n548_1) );
  AND2X2 AND2X2_207 ( .A(_abc_2290_n552), .B(_abc_2290_n551), .Y(_abc_2290_n553) );
  AND2X2 AND2X2_208 ( .A(_abc_2290_n555), .B(_abc_2290_n471), .Y(rx_countdown_4__FF_INPUT) );
  AND2X2 AND2X2_209 ( .A(_abc_2290_n557), .B(_abc_2290_n471), .Y(rx_countdown_5__FF_INPUT) );
  AND2X2 AND2X2_21 ( .A(_abc_2290_n183_1), .B(_abc_2290_n168), .Y(_abc_2290_n192) );
  AND2X2 AND2X2_210 ( .A(_abc_2290_n466), .B(rx), .Y(_abc_2290_n560) );
  AND2X2 AND2X2_211 ( .A(_abc_2290_n545), .B(_abc_2290_n561), .Y(_abc_2290_n562) );
  AND2X2 AND2X2_212 ( .A(_abc_2290_n563), .B(_abc_2290_n469_1), .Y(_abc_2290_n564) );
  AND2X2 AND2X2_213 ( .A(_abc_2290_n565), .B(_abc_2290_n566), .Y(_abc_2290_n567) );
  AND2X2 AND2X2_214 ( .A(_abc_2290_n568), .B(rx_bits_remaining_0_), .Y(_abc_2290_n569) );
  AND2X2 AND2X2_215 ( .A(_abc_2290_n567), .B(_abc_2290_n569), .Y(_abc_2290_n570) );
  AND2X2 AND2X2_216 ( .A(_abc_2290_n570), .B(_abc_2290_n463), .Y(_abc_2290_n571) );
  AND2X2 AND2X2_217 ( .A(_abc_2290_n572), .B(_abc_2290_n559), .Y(_abc_2290_n573) );
  AND2X2 AND2X2_218 ( .A(_abc_2290_n457), .B(_abc_2290_n145), .Y(_abc_2290_n574) );
  AND2X2 AND2X2_219 ( .A(_abc_2290_n545), .B(rx), .Y(_abc_2290_n575) );
  AND2X2 AND2X2_22 ( .A(_abc_2290_n192), .B(_abc_2290_n191), .Y(_abc_2290_n193) );
  AND2X2 AND2X2_220 ( .A(_abc_2290_n576), .B(_abc_2290_n574), .Y(_abc_2290_n577) );
  AND2X2 AND2X2_221 ( .A(_abc_2290_n456), .B(_abc_2290_n150), .Y(_abc_2290_n578) );
  AND2X2 AND2X2_222 ( .A(_abc_2290_n584), .B(_abc_2290_n585), .Y(_abc_2290_n586) );
  AND2X2 AND2X2_223 ( .A(_abc_2290_n587), .B(_abc_2290_n582), .Y(_abc_2290_n588) );
  AND2X2 AND2X2_224 ( .A(_abc_2290_n592), .B(_abc_2290_n454), .Y(_abc_2290_n593) );
  AND2X2 AND2X2_225 ( .A(_abc_2290_n545), .B(_abc_2290_n594), .Y(_abc_2290_n595) );
  AND2X2 AND2X2_226 ( .A(_abc_2290_n548_1), .B(_abc_2290_n597), .Y(_abc_2290_n598) );
  AND2X2 AND2X2_227 ( .A(_abc_2290_n562), .B(_abc_2290_n469_1), .Y(_abc_2290_n599) );
  AND2X2 AND2X2_228 ( .A(_abc_2290_n600), .B(rx_bits_remaining_0_), .Y(_abc_2290_n601) );
  AND2X2 AND2X2_229 ( .A(_abc_2290_n468), .B(rx_bits_remaining_1_), .Y(_abc_2290_n604) );
  AND2X2 AND2X2_23 ( .A(_abc_2290_n193), .B(_abc_2290_n162), .Y(_abc_2290_n194) );
  AND2X2 AND2X2_230 ( .A(_abc_2290_n597), .B(rx_bits_remaining_1_), .Y(_abc_2290_n606) );
  AND2X2 AND2X2_231 ( .A(_abc_2290_n545), .B(_abc_2290_n606), .Y(_abc_2290_n607) );
  AND2X2 AND2X2_232 ( .A(_abc_2290_n605), .B(_abc_2290_n608), .Y(_abc_2290_n609) );
  AND2X2 AND2X2_233 ( .A(_abc_2290_n611), .B(_abc_2290_n603), .Y(rx_bits_remaining_1__FF_INPUT) );
  AND2X2 AND2X2_234 ( .A(_abc_2290_n564), .B(rx_bits_remaining_2_), .Y(_abc_2290_n613) );
  AND2X2 AND2X2_235 ( .A(_abc_2290_n468), .B(rx_bits_remaining_2_), .Y(_abc_2290_n614) );
  AND2X2 AND2X2_236 ( .A(_abc_2290_n566), .B(_abc_2290_n597), .Y(_abc_2290_n615) );
  AND2X2 AND2X2_237 ( .A(_abc_2290_n615), .B(_abc_2290_n565), .Y(_abc_2290_n616) );
  AND2X2 AND2X2_238 ( .A(_abc_2290_n617), .B(rx_bits_remaining_2_), .Y(_abc_2290_n618) );
  AND2X2 AND2X2_239 ( .A(_abc_2290_n548_1), .B(_abc_2290_n619), .Y(_abc_2290_n620) );
  AND2X2 AND2X2_24 ( .A(_abc_2290_n190), .B(_abc_2290_n194), .Y(_abc_2290_n195_1) );
  AND2X2 AND2X2_240 ( .A(_abc_2290_n548_1), .B(_abc_2290_n616), .Y(_abc_2290_n623) );
  AND2X2 AND2X2_241 ( .A(_abc_2290_n624), .B(rx_bits_remaining_3_), .Y(_abc_2290_n625) );
  AND2X2 AND2X2_242 ( .A(_abc_2290_n623), .B(_abc_2290_n568), .Y(_abc_2290_n626) );
  AND2X2 AND2X2_243 ( .A(_abc_2290_n364), .B(_abc_2290_n163), .Y(tx_clk_divider_0__FF_INPUT) );
  AND2X2 AND2X2_244 ( .A(tx_clk_divider_0_), .B(tx_clk_divider_1_), .Y(_abc_2290_n630) );
  AND2X2 AND2X2_245 ( .A(_abc_2290_n634), .B(tx_clk_divider_2_), .Y(_abc_2290_n637) );
  AND2X2 AND2X2_246 ( .A(_abc_2290_n635), .B(tx_clk_divider_3_), .Y(_abc_2290_n640) );
  AND2X2 AND2X2_247 ( .A(_abc_2290_n641), .B(_abc_2290_n364), .Y(tx_clk_divider_3__FF_INPUT) );
  AND2X2 AND2X2_248 ( .A(_abc_2290_n175_1), .B(tx_clk_divider_4_), .Y(_abc_2290_n643) );
  AND2X2 AND2X2_249 ( .A(_abc_2290_n647), .B(_abc_2290_n364), .Y(tx_clk_divider_5__FF_INPUT) );
  AND2X2 AND2X2_25 ( .A(_abc_2290_n186), .B(_abc_2290_n195_1), .Y(_abc_2290_n196) );
  AND2X2 AND2X2_250 ( .A(_abc_2290_n187), .B(tx_clk_divider_6_), .Y(_abc_2290_n649) );
  AND2X2 AND2X2_251 ( .A(_abc_2290_n650), .B(_abc_2290_n364), .Y(tx_clk_divider_6__FF_INPUT) );
  AND2X2 AND2X2_252 ( .A(_abc_2290_n652), .B(_abc_2290_n364), .Y(tx_clk_divider_7__FF_INPUT) );
  AND2X2 AND2X2_253 ( .A(_abc_2290_n656), .B(_abc_2290_n364), .Y(tx_clk_divider_9__FF_INPUT) );
  AND2X2 AND2X2_254 ( .A(_abc_2290_n551), .B(_abc_2290_n400), .Y(rx_clk_divider_0__FF_INPUT) );
  AND2X2 AND2X2_255 ( .A(rx_clk_divider_0_), .B(rx_clk_divider_1_), .Y(_abc_2290_n661) );
  AND2X2 AND2X2_256 ( .A(_abc_2290_n402), .B(_abc_2290_n398_1), .Y(_abc_2290_n665) );
  AND2X2 AND2X2_257 ( .A(_abc_2290_n418), .B(rx_clk_divider_2_), .Y(_abc_2290_n666) );
  AND2X2 AND2X2_258 ( .A(_abc_2290_n670), .B(rx_clk_divider_3_), .Y(_abc_2290_n671) );
  AND2X2 AND2X2_259 ( .A(_abc_2290_n551), .B(_abc_2290_n672), .Y(rx_clk_divider_3__FF_INPUT) );
  AND2X2 AND2X2_26 ( .A(_abc_2290_n196), .B(_abc_2290_n181), .Y(_abc_2290_n197) );
  AND2X2 AND2X2_260 ( .A(_abc_2290_n551), .B(_abc_2290_n677), .Y(rx_clk_divider_5__FF_INPUT) );
  AND2X2 AND2X2_261 ( .A(_abc_2290_n551), .B(_abc_2290_n679), .Y(rx_clk_divider_6__FF_INPUT) );
  AND2X2 AND2X2_262 ( .A(_abc_2290_n681), .B(_abc_2290_n551), .Y(rx_clk_divider_7__FF_INPUT) );
  AND2X2 AND2X2_263 ( .A(_abc_2290_n686), .B(_abc_2290_n551), .Y(rx_clk_divider_9__FF_INPUT) );
  AND2X2 AND2X2_264 ( .A(_abc_2290_n548_1), .B(_abc_2290_n692), .Y(_abc_2290_n693) );
  AND2X2 AND2X2_265 ( .A(_abc_2290_n694), .B(_abc_2290_n691), .Y(rx_data_0__FF_INPUT) );
  AND2X2 AND2X2_266 ( .A(_abc_2290_n548_1), .B(_abc_2290_n697), .Y(_abc_2290_n698) );
  AND2X2 AND2X2_267 ( .A(_abc_2290_n699), .B(_abc_2290_n696), .Y(rx_data_1__FF_INPUT) );
  AND2X2 AND2X2_268 ( .A(_abc_2290_n548_1), .B(_abc_2290_n702), .Y(_abc_2290_n703) );
  AND2X2 AND2X2_269 ( .A(_abc_2290_n704), .B(_abc_2290_n701), .Y(rx_data_2__FF_INPUT) );
  AND2X2 AND2X2_27 ( .A(_abc_2290_n159), .B(_abc_2290_n199), .Y(_abc_2290_n200) );
  AND2X2 AND2X2_270 ( .A(_abc_2290_n548_1), .B(_abc_2290_n707), .Y(_abc_2290_n708) );
  AND2X2 AND2X2_271 ( .A(_abc_2290_n709), .B(_abc_2290_n706), .Y(rx_data_3__FF_INPUT) );
  AND2X2 AND2X2_272 ( .A(_abc_2290_n548_1), .B(_abc_2290_n712), .Y(_abc_2290_n713) );
  AND2X2 AND2X2_273 ( .A(_abc_2290_n714), .B(_abc_2290_n711), .Y(rx_data_4__FF_INPUT) );
  AND2X2 AND2X2_274 ( .A(_abc_2290_n548_1), .B(_abc_2290_n717), .Y(_abc_2290_n718) );
  AND2X2 AND2X2_275 ( .A(_abc_2290_n719), .B(_abc_2290_n716), .Y(rx_data_5__FF_INPUT) );
  AND2X2 AND2X2_276 ( .A(_abc_2290_n548_1), .B(_abc_2290_n722), .Y(_abc_2290_n723) );
  AND2X2 AND2X2_277 ( .A(_abc_2290_n724), .B(_abc_2290_n721), .Y(rx_data_6__FF_INPUT) );
  AND2X2 AND2X2_278 ( .A(_abc_2290_n548_1), .B(_abc_2290_n473_1), .Y(_abc_2290_n726) );
  AND2X2 AND2X2_279 ( .A(_abc_2290_n727), .B(_abc_2290_n728), .Y(rx_data_7__FF_INPUT) );
  AND2X2 AND2X2_28 ( .A(_abc_2290_n173), .B(_abc_2290_n200), .Y(_abc_2290_n201) );
  AND2X2 AND2X2_29 ( .A(_abc_2290_n202_1), .B(_abc_2290_n205), .Y(_abc_2290_n206) );
  AND2X2 AND2X2_3 ( .A(_abc_2290_n150), .B(_abc_2290_n144), .Y(received) );
  AND2X2 AND2X2_30 ( .A(_abc_2290_n207), .B(_abc_2290_n204), .Y(_abc_2290_n208) );
  AND2X2 AND2X2_31 ( .A(_abc_2290_n206), .B(_abc_2290_n208), .Y(_abc_2290_n209_1) );
  AND2X2 AND2X2_32 ( .A(_abc_2290_n209_1), .B(_abc_2290_n197), .Y(_abc_2290_n210) );
  AND2X2 AND2X2_33 ( .A(_abc_2290_n215), .B(_abc_2290_n216), .Y(_abc_2290_n217_1) );
  AND2X2 AND2X2_34 ( .A(_abc_2290_n217_1), .B(_abc_2290_n214), .Y(_abc_2290_n218) );
  AND2X2 AND2X2_35 ( .A(_abc_2290_n218), .B(_abc_2290_n213), .Y(_abc_2290_n219) );
  AND2X2 AND2X2_36 ( .A(_abc_2290_n219), .B(_abc_2290_n212), .Y(_abc_2290_n220) );
  AND2X2 AND2X2_37 ( .A(_abc_2290_n221), .B(_abc_2290_n211), .Y(_abc_2290_n222_1) );
  AND2X2 AND2X2_38 ( .A(_abc_2290_n220), .B(tx_countdown_5_), .Y(_abc_2290_n223) );
  AND2X2 AND2X2_39 ( .A(_abc_2290_n210), .B(_abc_2290_n224), .Y(_abc_2290_n225) );
  AND2X2 AND2X2_4 ( .A(recv_state_0_), .B(recv_state_2_), .Y(_abc_2290_n153) );
  AND2X2 AND2X2_40 ( .A(_abc_2290_n226), .B(_abc_2290_n227_1), .Y(_abc_2290_n228) );
  AND2X2 AND2X2_41 ( .A(_abc_2290_n229), .B(_abc_2290_n214), .Y(_abc_2290_n230) );
  AND2X2 AND2X2_42 ( .A(_abc_2290_n217_1), .B(tx_countdown_2_), .Y(_abc_2290_n231) );
  AND2X2 AND2X2_43 ( .A(_abc_2290_n210), .B(_abc_2290_n232_1), .Y(_abc_2290_n233) );
  AND2X2 AND2X2_44 ( .A(_abc_2290_n234), .B(_abc_2290_n235), .Y(_abc_2290_n236) );
  AND2X2 AND2X2_45 ( .A(_abc_2290_n210), .B(tx_countdown_0_), .Y(_abc_2290_n239) );
  AND2X2 AND2X2_46 ( .A(_abc_2290_n244), .B(_abc_2290_n213), .Y(_abc_2290_n245_1) );
  AND2X2 AND2X2_47 ( .A(_abc_2290_n218), .B(tx_countdown_3_), .Y(_abc_2290_n246) );
  AND2X2 AND2X2_48 ( .A(_abc_2290_n210), .B(_abc_2290_n247), .Y(_abc_2290_n248) );
  AND2X2 AND2X2_49 ( .A(_abc_2290_n249), .B(_abc_2290_n250_1), .Y(_abc_2290_n251) );
  AND2X2 AND2X2_5 ( .A(_abc_2290_n153), .B(_abc_2290_n152_1), .Y(recv_error) );
  AND2X2 AND2X2_50 ( .A(_abc_2290_n216), .B(tx_countdown_0_), .Y(_abc_2290_n252) );
  AND2X2 AND2X2_51 ( .A(_abc_2290_n215), .B(tx_countdown_1_), .Y(_abc_2290_n253) );
  AND2X2 AND2X2_52 ( .A(_abc_2290_n210), .B(_abc_2290_n254), .Y(_abc_2290_n255) );
  AND2X2 AND2X2_53 ( .A(_abc_2290_n256), .B(_abc_2290_n257_1), .Y(_abc_2290_n258_1) );
  AND2X2 AND2X2_54 ( .A(_abc_2290_n262), .B(_abc_2290_n263), .Y(_abc_2290_n264_1) );
  AND2X2 AND2X2_55 ( .A(_abc_2290_n270_1), .B(_abc_2290_n158), .Y(_abc_2290_n271_1) );
  AND2X2 AND2X2_56 ( .A(_abc_2290_n271_1), .B(tx_data_1_), .Y(_abc_2290_n272) );
  AND2X2 AND2X2_57 ( .A(is_transmitting), .B(_abc_2290_n156_1), .Y(_abc_2290_n273_1) );
  AND2X2 AND2X2_58 ( .A(_abc_2290_n274_1), .B(transmit), .Y(_abc_2290_n275) );
  AND2X2 AND2X2_59 ( .A(_abc_2290_n275), .B(\tx_byte[0] ), .Y(_abc_2290_n276) );
  AND2X2 AND2X2_6 ( .A(_abc_2290_n156_1), .B(tx_state_0_), .Y(_abc_2290_n157_1) );
  AND2X2 AND2X2_60 ( .A(_abc_2290_n156_1), .B(tx_state_1_), .Y(_abc_2290_n277) );
  AND2X2 AND2X2_61 ( .A(_abc_2290_n274_1), .B(_abc_2290_n278), .Y(_abc_2290_n279) );
  AND2X2 AND2X2_62 ( .A(_abc_2290_n280), .B(tx_data_0_), .Y(_abc_2290_n281_1) );
  AND2X2 AND2X2_63 ( .A(_abc_2290_n269), .B(_abc_2290_n158), .Y(_abc_2290_n283) );
  AND2X2 AND2X2_64 ( .A(_abc_2290_n283), .B(tx_data_0_), .Y(_abc_2290_n284) );
  AND2X2 AND2X2_65 ( .A(_abc_2290_n271_1), .B(tx_data_2_), .Y(_abc_2290_n287) );
  AND2X2 AND2X2_66 ( .A(_abc_2290_n275), .B(\tx_byte[1] ), .Y(_abc_2290_n288) );
  AND2X2 AND2X2_67 ( .A(_abc_2290_n280), .B(tx_data_1_), .Y(_abc_2290_n289) );
  AND2X2 AND2X2_68 ( .A(_abc_2290_n283), .B(tx_data_1_), .Y(_abc_2290_n291) );
  AND2X2 AND2X2_69 ( .A(_abc_2290_n271_1), .B(tx_data_3_), .Y(_abc_2290_n294) );
  AND2X2 AND2X2_7 ( .A(_abc_2290_n157_1), .B(_abc_2290_n155), .Y(_abc_2290_n158) );
  AND2X2 AND2X2_70 ( .A(_abc_2290_n275), .B(\tx_byte[2] ), .Y(_abc_2290_n295) );
  AND2X2 AND2X2_71 ( .A(_abc_2290_n280), .B(tx_data_2_), .Y(_abc_2290_n296) );
  AND2X2 AND2X2_72 ( .A(_abc_2290_n283), .B(tx_data_2_), .Y(_abc_2290_n298) );
  AND2X2 AND2X2_73 ( .A(_abc_2290_n271_1), .B(tx_data_4_), .Y(_abc_2290_n301) );
  AND2X2 AND2X2_74 ( .A(_abc_2290_n275), .B(\tx_byte[3] ), .Y(_abc_2290_n302) );
  AND2X2 AND2X2_75 ( .A(_abc_2290_n280), .B(tx_data_3_), .Y(_abc_2290_n303) );
  AND2X2 AND2X2_76 ( .A(_abc_2290_n283), .B(tx_data_3_), .Y(_abc_2290_n305) );
  AND2X2 AND2X2_77 ( .A(_abc_2290_n271_1), .B(tx_data_5_), .Y(_abc_2290_n308) );
  AND2X2 AND2X2_78 ( .A(_abc_2290_n275), .B(\tx_byte[4] ), .Y(_abc_2290_n309) );
  AND2X2 AND2X2_79 ( .A(_abc_2290_n280), .B(tx_data_4_), .Y(_abc_2290_n310) );
  AND2X2 AND2X2_8 ( .A(_abc_2290_n160), .B(_abc_2290_n161_1), .Y(_abc_2290_n162) );
  AND2X2 AND2X2_80 ( .A(_abc_2290_n283), .B(tx_data_4_), .Y(_abc_2290_n312_1) );
  AND2X2 AND2X2_81 ( .A(_abc_2290_n271_1), .B(tx_data_6_), .Y(_abc_2290_n315) );
  AND2X2 AND2X2_82 ( .A(_abc_2290_n275), .B(\tx_byte[5] ), .Y(_abc_2290_n316) );
  AND2X2 AND2X2_83 ( .A(_abc_2290_n280), .B(tx_data_5_), .Y(_abc_2290_n317) );
  AND2X2 AND2X2_84 ( .A(_abc_2290_n283), .B(tx_data_5_), .Y(_abc_2290_n319_1) );
  AND2X2 AND2X2_85 ( .A(_abc_2290_n275), .B(\tx_byte[6] ), .Y(_abc_2290_n322) );
  AND2X2 AND2X2_86 ( .A(_abc_2290_n280), .B(tx_data_6_), .Y(_abc_2290_n323_1) );
  AND2X2 AND2X2_87 ( .A(_abc_2290_n158), .B(tx_data_7_), .Y(_abc_2290_n326) );
  AND2X2 AND2X2_88 ( .A(_abc_2290_n327), .B(_abc_2290_n325), .Y(_abc_2290_n328) );
  AND2X2 AND2X2_89 ( .A(_abc_2290_n275), .B(\tx_byte[7] ), .Y(_abc_2290_n330) );
  AND2X2 AND2X2_9 ( .A(_abc_2290_n163), .B(_abc_2290_n164), .Y(_abc_2290_n165_1) );
  AND2X2 AND2X2_90 ( .A(_abc_2290_n331), .B(tx_data_7_), .Y(_abc_2290_n332) );
  AND2X2 AND2X2_91 ( .A(_abc_2290_n335), .B(_abc_2290_n158), .Y(_abc_2290_n336) );
  AND2X2 AND2X2_92 ( .A(_abc_2290_n280), .B(tx_bits_remaining_0_), .Y(_abc_2290_n337) );
  AND2X2 AND2X2_93 ( .A(_abc_2290_n338), .B(_abc_2290_n334), .Y(tx_bits_remaining_0__FF_INPUT) );
  AND2X2 AND2X2_94 ( .A(_abc_2290_n340), .B(_abc_2290_n341), .Y(_abc_2290_n342) );
  AND2X2 AND2X2_95 ( .A(_abc_2290_n267_1), .B(_abc_2290_n342), .Y(_abc_2290_n343) );
  AND2X2 AND2X2_96 ( .A(_abc_2290_n346), .B(_abc_2290_n344_1), .Y(_abc_2290_n347) );
  AND2X2 AND2X2_97 ( .A(_abc_2290_n347), .B(_abc_2290_n158), .Y(_abc_2290_n348) );
  AND2X2 AND2X2_98 ( .A(_abc_2290_n280), .B(tx_bits_remaining_1_), .Y(_abc_2290_n349) );
  AND2X2 AND2X2_99 ( .A(_abc_2290_n345), .B(_abc_2290_n351), .Y(_abc_2290_n352_1) );
  DFFPOSX1 DFFPOSX1_1 ( .CLK(clk), .D(rx_clk_divider_2__FF_INPUT), .Q(rx_clk_divider_2_) );
  DFFPOSX1 DFFPOSX1_10 ( .CLK(clk), .D(tx_clk_divider_0__FF_INPUT), .Q(tx_clk_divider_0_) );
  DFFPOSX1 DFFPOSX1_11 ( .CLK(clk), .D(tx_clk_divider_1__FF_INPUT), .Q(tx_clk_divider_1_) );
  DFFPOSX1 DFFPOSX1_12 ( .CLK(clk), .D(tx_clk_divider_2__FF_INPUT), .Q(tx_clk_divider_2_) );
  DFFPOSX1 DFFPOSX1_13 ( .CLK(clk), .D(tx_clk_divider_3__FF_INPUT), .Q(tx_clk_divider_3_) );
  DFFPOSX1 DFFPOSX1_14 ( .CLK(clk), .D(tx_clk_divider_4__FF_INPUT), .Q(tx_clk_divider_4_) );
  DFFPOSX1 DFFPOSX1_15 ( .CLK(clk), .D(tx_clk_divider_5__FF_INPUT), .Q(tx_clk_divider_5_) );
  DFFPOSX1 DFFPOSX1_16 ( .CLK(clk), .D(tx_clk_divider_6__FF_INPUT), .Q(tx_clk_divider_6_) );
  DFFPOSX1 DFFPOSX1_17 ( .CLK(clk), .D(tx_clk_divider_7__FF_INPUT), .Q(tx_clk_divider_7_) );
  DFFPOSX1 DFFPOSX1_18 ( .CLK(clk), .D(tx_clk_divider_8__FF_INPUT), .Q(tx_clk_divider_8_) );
  DFFPOSX1 DFFPOSX1_19 ( .CLK(clk), .D(tx_clk_divider_9__FF_INPUT), .Q(tx_clk_divider_9_) );
  DFFPOSX1 DFFPOSX1_2 ( .CLK(clk), .D(rx_clk_divider_3__FF_INPUT), .Q(rx_clk_divider_3_) );
  DFFPOSX1 DFFPOSX1_20 ( .CLK(clk), .D(tx_clk_divider_10__FF_INPUT), .Q(tx_clk_divider_10_) );
  DFFPOSX1 DFFPOSX1_21 ( .CLK(clk), .D(recv_state_0__FF_INPUT), .Q(recv_state_0_) );
  DFFPOSX1 DFFPOSX1_22 ( .CLK(clk), .D(recv_state_1__FF_INPUT), .Q(recv_state_1_) );
  DFFPOSX1 DFFPOSX1_23 ( .CLK(clk), .D(recv_state_2__FF_INPUT), .Q(recv_state_2_) );
  DFFPOSX1 DFFPOSX1_24 ( .CLK(clk), .D(rx_countdown_0__FF_INPUT), .Q(rx_countdown_0_) );
  DFFPOSX1 DFFPOSX1_25 ( .CLK(clk), .D(rx_countdown_1__FF_INPUT), .Q(rx_countdown_1_) );
  DFFPOSX1 DFFPOSX1_26 ( .CLK(clk), .D(rx_countdown_2__FF_INPUT), .Q(rx_countdown_2_) );
  DFFPOSX1 DFFPOSX1_27 ( .CLK(clk), .D(rx_countdown_3__FF_INPUT), .Q(rx_countdown_3_) );
  DFFPOSX1 DFFPOSX1_28 ( .CLK(clk), .D(rx_countdown_4__FF_INPUT), .Q(rx_countdown_4_) );
  DFFPOSX1 DFFPOSX1_29 ( .CLK(clk), .D(rx_countdown_5__FF_INPUT), .Q(rx_countdown_5_) );
  DFFPOSX1 DFFPOSX1_3 ( .CLK(clk), .D(rx_clk_divider_4__FF_INPUT), .Q(rx_clk_divider_4_) );
  DFFPOSX1 DFFPOSX1_30 ( .CLK(clk), .D(rx_bits_remaining_0__FF_INPUT), .Q(rx_bits_remaining_0_) );
  DFFPOSX1 DFFPOSX1_31 ( .CLK(clk), .D(rx_bits_remaining_1__FF_INPUT), .Q(rx_bits_remaining_1_) );
  DFFPOSX1 DFFPOSX1_32 ( .CLK(clk), .D(rx_bits_remaining_2__FF_INPUT), .Q(rx_bits_remaining_2_) );
  DFFPOSX1 DFFPOSX1_33 ( .CLK(clk), .D(rx_bits_remaining_3__FF_INPUT), .Q(rx_bits_remaining_3_) );
  DFFPOSX1 DFFPOSX1_34 ( .CLK(clk), .D(rx_data_0__FF_INPUT), .Q(\rx_byte[0] ) );
  DFFPOSX1 DFFPOSX1_35 ( .CLK(clk), .D(rx_data_1__FF_INPUT), .Q(\rx_byte[1] ) );
  DFFPOSX1 DFFPOSX1_36 ( .CLK(clk), .D(rx_data_2__FF_INPUT), .Q(\rx_byte[2] ) );
  DFFPOSX1 DFFPOSX1_37 ( .CLK(clk), .D(rx_data_3__FF_INPUT), .Q(\rx_byte[3] ) );
  DFFPOSX1 DFFPOSX1_38 ( .CLK(clk), .D(rx_data_4__FF_INPUT), .Q(\rx_byte[4] ) );
  DFFPOSX1 DFFPOSX1_39 ( .CLK(clk), .D(rx_data_5__FF_INPUT), .Q(\rx_byte[5] ) );
  DFFPOSX1 DFFPOSX1_4 ( .CLK(clk), .D(rx_clk_divider_5__FF_INPUT), .Q(rx_clk_divider_5_) );
  DFFPOSX1 DFFPOSX1_40 ( .CLK(clk), .D(rx_data_6__FF_INPUT), .Q(\rx_byte[6] ) );
  DFFPOSX1 DFFPOSX1_41 ( .CLK(clk), .D(rx_data_7__FF_INPUT), .Q(\rx_byte[7] ) );
  DFFPOSX1 DFFPOSX1_42 ( .CLK(clk), .D(tx_out_FF_INPUT), .Q(tx) );
  DFFPOSX1 DFFPOSX1_43 ( .CLK(clk), .D(tx_state_0__FF_INPUT), .Q(tx_state_0_) );
  DFFPOSX1 DFFPOSX1_44 ( .CLK(clk), .D(tx_state_1__FF_INPUT), .Q(tx_state_1_) );
  DFFPOSX1 DFFPOSX1_45 ( .CLK(clk), .D(tx_countdown_0__FF_INPUT), .Q(tx_countdown_0_) );
  DFFPOSX1 DFFPOSX1_46 ( .CLK(clk), .D(tx_countdown_1__FF_INPUT), .Q(tx_countdown_1_) );
  DFFPOSX1 DFFPOSX1_47 ( .CLK(clk), .D(tx_countdown_2__FF_INPUT), .Q(tx_countdown_2_) );
  DFFPOSX1 DFFPOSX1_48 ( .CLK(clk), .D(tx_countdown_3__FF_INPUT), .Q(tx_countdown_3_) );
  DFFPOSX1 DFFPOSX1_49 ( .CLK(clk), .D(tx_countdown_4__FF_INPUT), .Q(tx_countdown_4_) );
  DFFPOSX1 DFFPOSX1_5 ( .CLK(clk), .D(rx_clk_divider_6__FF_INPUT), .Q(rx_clk_divider_6_) );
  DFFPOSX1 DFFPOSX1_50 ( .CLK(clk), .D(tx_countdown_5__FF_INPUT), .Q(tx_countdown_5_) );
  DFFPOSX1 DFFPOSX1_51 ( .CLK(clk), .D(tx_bits_remaining_0__FF_INPUT), .Q(tx_bits_remaining_0_) );
  DFFPOSX1 DFFPOSX1_52 ( .CLK(clk), .D(tx_bits_remaining_1__FF_INPUT), .Q(tx_bits_remaining_1_) );
  DFFPOSX1 DFFPOSX1_53 ( .CLK(clk), .D(tx_bits_remaining_2__FF_INPUT), .Q(tx_bits_remaining_2_) );
  DFFPOSX1 DFFPOSX1_54 ( .CLK(clk), .D(tx_bits_remaining_3__FF_INPUT), .Q(tx_bits_remaining_3_) );
  DFFPOSX1 DFFPOSX1_55 ( .CLK(clk), .D(tx_data_0__FF_INPUT), .Q(tx_data_0_) );
  DFFPOSX1 DFFPOSX1_56 ( .CLK(clk), .D(tx_data_1__FF_INPUT), .Q(tx_data_1_) );
  DFFPOSX1 DFFPOSX1_57 ( .CLK(clk), .D(tx_data_2__FF_INPUT), .Q(tx_data_2_) );
  DFFPOSX1 DFFPOSX1_58 ( .CLK(clk), .D(tx_data_3__FF_INPUT), .Q(tx_data_3_) );
  DFFPOSX1 DFFPOSX1_59 ( .CLK(clk), .D(tx_data_4__FF_INPUT), .Q(tx_data_4_) );
  DFFPOSX1 DFFPOSX1_6 ( .CLK(clk), .D(rx_clk_divider_7__FF_INPUT), .Q(rx_clk_divider_7_) );
  DFFPOSX1 DFFPOSX1_60 ( .CLK(clk), .D(tx_data_5__FF_INPUT), .Q(tx_data_5_) );
  DFFPOSX1 DFFPOSX1_61 ( .CLK(clk), .D(tx_data_6__FF_INPUT), .Q(tx_data_6_) );
  DFFPOSX1 DFFPOSX1_62 ( .CLK(clk), .D(tx_data_7__FF_INPUT), .Q(tx_data_7_) );
  DFFPOSX1 DFFPOSX1_63 ( .CLK(clk), .D(rx_clk_divider_0__FF_INPUT), .Q(rx_clk_divider_0_) );
  DFFPOSX1 DFFPOSX1_64 ( .CLK(clk), .D(rx_clk_divider_1__FF_INPUT), .Q(rx_clk_divider_1_) );
  DFFPOSX1 DFFPOSX1_7 ( .CLK(clk), .D(rx_clk_divider_8__FF_INPUT), .Q(rx_clk_divider_8_) );
  DFFPOSX1 DFFPOSX1_8 ( .CLK(clk), .D(rx_clk_divider_9__FF_INPUT), .Q(rx_clk_divider_9_) );
  DFFPOSX1 DFFPOSX1_9 ( .CLK(clk), .D(rx_clk_divider_10__FF_INPUT), .Q(rx_clk_divider_10_) );
  INVX1 INVX1_1 ( .A(recv_state_0_), .Y(_abc_2290_n144) );
  INVX1 INVX1_10 ( .A(tx_clk_divider_1_), .Y(_abc_2290_n164) );
  INVX1 INVX1_100 ( .A(_abc_2290_n609), .Y(_abc_2290_n610) );
  INVX1 INVX1_101 ( .A(_abc_2290_n615), .Y(_abc_2290_n617) );
  INVX1 INVX1_102 ( .A(_abc_2290_n623), .Y(_abc_2290_n624) );
  INVX1 INVX1_103 ( .A(_abc_2290_n165_1), .Y(_abc_2290_n634) );
  INVX1 INVX1_104 ( .A(_abc_2290_n635), .Y(_abc_2290_n636) );
  INVX1 INVX1_105 ( .A(_abc_2290_n190), .Y(_abc_2290_n647) );
  INVX1 INVX1_106 ( .A(_abc_2290_n186), .Y(_abc_2290_n652) );
  INVX1 INVX1_107 ( .A(_abc_2290_n208), .Y(_abc_2290_n656) );
  INVX1 INVX1_108 ( .A(_abc_2290_n206), .Y(_abc_2290_n658) );
  INVX1 INVX1_109 ( .A(_abc_2290_n665), .Y(_abc_2290_n670) );
  INVX1 INVX1_11 ( .A(tx_clk_divider_5_), .Y(_abc_2290_n167) );
  INVX1 INVX1_110 ( .A(_abc_2290_n489_1), .Y(_abc_2290_n674) );
  INVX1 INVX1_111 ( .A(_abc_2290_n438), .Y(_abc_2290_n677) );
  INVX1 INVX1_112 ( .A(_abc_2290_n435), .Y(_abc_2290_n679) );
  INVX1 INVX1_113 ( .A(_abc_2290_n432), .Y(_abc_2290_n681) );
  INVX1 INVX1_114 ( .A(_abc_2290_n496_1), .Y(_abc_2290_n683) );
  INVX1 INVX1_115 ( .A(_abc_2290_n427_1), .Y(_abc_2290_n686) );
  INVX1 INVX1_116 ( .A(_abc_2290_n485), .Y(_abc_2290_n688) );
  INVX1 INVX1_117 ( .A(\rx_byte[1] ), .Y(_abc_2290_n692) );
  INVX1 INVX1_118 ( .A(_abc_2290_n693), .Y(_abc_2290_n694) );
  INVX1 INVX1_119 ( .A(\rx_byte[2] ), .Y(_abc_2290_n697) );
  INVX1 INVX1_12 ( .A(tx_clk_divider_4_), .Y(_abc_2290_n168) );
  INVX1 INVX1_120 ( .A(_abc_2290_n698), .Y(_abc_2290_n699) );
  INVX1 INVX1_121 ( .A(\rx_byte[3] ), .Y(_abc_2290_n702) );
  INVX1 INVX1_122 ( .A(_abc_2290_n703), .Y(_abc_2290_n704) );
  INVX1 INVX1_123 ( .A(\rx_byte[4] ), .Y(_abc_2290_n707) );
  INVX1 INVX1_124 ( .A(_abc_2290_n708), .Y(_abc_2290_n709) );
  INVX1 INVX1_125 ( .A(\rx_byte[5] ), .Y(_abc_2290_n712) );
  INVX1 INVX1_126 ( .A(_abc_2290_n713), .Y(_abc_2290_n714) );
  INVX1 INVX1_127 ( .A(\rx_byte[6] ), .Y(_abc_2290_n717) );
  INVX1 INVX1_128 ( .A(_abc_2290_n718), .Y(_abc_2290_n719) );
  INVX1 INVX1_129 ( .A(\rx_byte[7] ), .Y(_abc_2290_n722) );
  INVX1 INVX1_13 ( .A(_abc_2290_n171), .Y(_abc_2290_n172) );
  INVX1 INVX1_130 ( .A(_abc_2290_n723), .Y(_abc_2290_n724) );
  INVX1 INVX1_131 ( .A(_abc_2290_n726), .Y(_abc_2290_n727) );
  INVX1 INVX1_14 ( .A(_abc_2290_n166_1), .Y(_abc_2290_n175_1) );
  INVX1 INVX1_15 ( .A(_abc_2290_n169), .Y(_abc_2290_n176) );
  INVX1 INVX1_16 ( .A(_abc_2290_n180), .Y(_abc_2290_n181) );
  INVX1 INVX1_17 ( .A(tx_clk_divider_7_), .Y(_abc_2290_n182) );
  INVX1 INVX1_18 ( .A(tx_clk_divider_6_), .Y(_abc_2290_n183_1) );
  INVX1 INVX1_19 ( .A(_abc_2290_n170_1), .Y(_abc_2290_n187) );
  INVX1 INVX1_2 ( .A(recv_state_2_), .Y(_abc_2290_n145) );
  INVX1 INVX1_20 ( .A(tx_clk_divider_10_), .Y(_abc_2290_n198) );
  INVX1 INVX1_21 ( .A(tx_clk_divider_9_), .Y(_abc_2290_n199) );
  INVX1 INVX1_22 ( .A(_abc_2290_n200), .Y(_abc_2290_n203) );
  INVX1 INVX1_23 ( .A(tx_countdown_5_), .Y(_abc_2290_n211) );
  INVX1 INVX1_24 ( .A(tx_countdown_4_), .Y(_abc_2290_n212) );
  INVX1 INVX1_25 ( .A(tx_countdown_3_), .Y(_abc_2290_n213) );
  INVX1 INVX1_26 ( .A(tx_countdown_2_), .Y(_abc_2290_n214) );
  INVX1 INVX1_27 ( .A(tx_countdown_0_), .Y(_abc_2290_n215) );
  INVX1 INVX1_28 ( .A(tx_countdown_1_), .Y(_abc_2290_n216) );
  INVX1 INVX1_29 ( .A(_abc_2290_n220), .Y(_abc_2290_n221) );
  INVX1 INVX1_3 ( .A(_abc_2290_n146), .Y(_abc_2290_n147_1) );
  INVX1 INVX1_30 ( .A(_abc_2290_n225), .Y(_abc_2290_n226) );
  INVX1 INVX1_31 ( .A(_abc_2290_n217_1), .Y(_abc_2290_n229) );
  INVX1 INVX1_32 ( .A(_abc_2290_n233), .Y(_abc_2290_n234) );
  INVX1 INVX1_33 ( .A(_abc_2290_n240), .Y(_abc_2290_n241_1) );
  INVX1 INVX1_34 ( .A(_abc_2290_n242), .Y(_abc_2290_n243) );
  INVX1 INVX1_35 ( .A(_abc_2290_n218), .Y(_abc_2290_n244) );
  INVX1 INVX1_36 ( .A(_abc_2290_n248), .Y(_abc_2290_n249) );
  INVX1 INVX1_37 ( .A(_abc_2290_n255), .Y(_abc_2290_n256) );
  INVX1 INVX1_38 ( .A(tx_bits_remaining_1_), .Y(_abc_2290_n262) );
  INVX1 INVX1_39 ( .A(tx_bits_remaining_0_), .Y(_abc_2290_n263) );
  INVX1 INVX1_4 ( .A(recv_state_1_), .Y(_abc_2290_n152_1) );
  INVX1 INVX1_40 ( .A(_abc_2290_n264_1), .Y(_abc_2290_n265_1) );
  INVX1 INVX1_41 ( .A(_abc_2290_n267_1), .Y(_abc_2290_n268_1) );
  INVX1 INVX1_42 ( .A(_abc_2290_n269), .Y(_abc_2290_n270_1) );
  INVX1 INVX1_43 ( .A(_abc_2290_n273_1), .Y(_abc_2290_n274_1) );
  INVX1 INVX1_44 ( .A(transmit), .Y(_abc_2290_n278) );
  INVX1 INVX1_45 ( .A(_abc_2290_n266), .Y(_abc_2290_n351) );
  INVX1 INVX1_46 ( .A(_abc_2290_n360), .Y(_abc_2290_n361) );
  INVX1 INVX1_47 ( .A(_abc_2290_n375), .Y(_abc_2290_n377) );
  INVX1 INVX1_48 ( .A(_abc_2290_n383), .Y(_abc_2290_n384) );
  INVX1 INVX1_49 ( .A(rx_countdown_0_), .Y(_abc_2290_n396) );
  INVX1 INVX1_5 ( .A(tx_state_1_), .Y(_abc_2290_n155) );
  INVX1 INVX1_50 ( .A(rx_clk_divider_3_), .Y(_abc_2290_n397) );
  INVX1 INVX1_51 ( .A(rx_clk_divider_2_), .Y(_abc_2290_n398_1) );
  INVX1 INVX1_52 ( .A(rx_clk_divider_0_), .Y(_abc_2290_n400) );
  INVX1 INVX1_53 ( .A(rx_clk_divider_1_), .Y(_abc_2290_n401) );
  INVX1 INVX1_54 ( .A(rx_clk_divider_5_), .Y(_abc_2290_n404_1) );
  INVX1 INVX1_55 ( .A(rx_clk_divider_4_), .Y(_abc_2290_n405) );
  INVX1 INVX1_56 ( .A(rx_clk_divider_6_), .Y(_abc_2290_n407) );
  INVX1 INVX1_57 ( .A(rx_clk_divider_7_), .Y(_abc_2290_n408) );
  INVX1 INVX1_58 ( .A(rx_clk_divider_8_), .Y(_abc_2290_n412) );
  INVX1 INVX1_59 ( .A(rx_clk_divider_9_), .Y(_abc_2290_n413) );
  INVX1 INVX1_6 ( .A(tx_clk_divider_8_), .Y(_abc_2290_n159) );
  INVX1 INVX1_60 ( .A(_abc_2290_n415), .Y(_abc_2290_n416) );
  INVX1 INVX1_61 ( .A(_abc_2290_n424), .Y(_abc_2290_n425_1) );
  INVX1 INVX1_62 ( .A(_abc_2290_n429), .Y(_abc_2290_n430) );
  INVX1 INVX1_63 ( .A(rx_clk_divider_10_), .Y(_abc_2290_n439) );
  INVX1 INVX1_64 ( .A(_abc_2290_n450), .Y(_abc_2290_n451) );
  INVX1 INVX1_65 ( .A(_abc_2290_n452), .Y(_abc_2290_n453) );
  INVX1 INVX1_66 ( .A(_abc_2290_n459_1), .Y(_abc_2290_n460) );
  INVX1 INVX1_67 ( .A(_abc_2290_n463), .Y(_abc_2290_n464_1) );
  INVX1 INVX1_68 ( .A(_abc_2290_n466), .Y(_abc_2290_n467) );
  INVX1 INVX1_69 ( .A(_abc_2290_n468), .Y(_abc_2290_n469_1) );
  INVX1 INVX1_7 ( .A(tx_clk_divider_3_), .Y(_abc_2290_n160) );
  INVX1 INVX1_70 ( .A(rx), .Y(_abc_2290_n473_1) );
  INVX1 INVX1_71 ( .A(rx_countdown_1_), .Y(_abc_2290_n476) );
  INVX1 INVX1_72 ( .A(_abc_2290_n479_1), .Y(_abc_2290_n480) );
  INVX1 INVX1_73 ( .A(rx_countdown_2_), .Y(_abc_2290_n501) );
  INVX1 INVX1_74 ( .A(_abc_2290_n502_1), .Y(_abc_2290_n504) );
  INVX1 INVX1_75 ( .A(_abc_2290_n507_1), .Y(_abc_2290_n508) );
  INVX1 INVX1_76 ( .A(_abc_2290_n510_1), .Y(_abc_2290_n511) );
  INVX1 INVX1_77 ( .A(rx_countdown_4_), .Y(_abc_2290_n514_1) );
  INVX1 INVX1_78 ( .A(rx_countdown_3_), .Y(_abc_2290_n515) );
  INVX1 INVX1_79 ( .A(_abc_2290_n517), .Y(_abc_2290_n518_1) );
  INVX1 INVX1_8 ( .A(tx_clk_divider_2_), .Y(_abc_2290_n161_1) );
  INVX1 INVX1_80 ( .A(rx_countdown_5_), .Y(_abc_2290_n520_1) );
  INVX1 INVX1_81 ( .A(_abc_2290_n523), .Y(_abc_2290_n524_1) );
  INVX1 INVX1_82 ( .A(_abc_2290_n516_1), .Y(_abc_2290_n527) );
  INVX1 INVX1_83 ( .A(_abc_2290_n530), .Y(_abc_2290_n531_1) );
  INVX1 INVX1_84 ( .A(_abc_2290_n503), .Y(_abc_2290_n535_1) );
  INVX1 INVX1_85 ( .A(_abc_2290_n539), .Y(_abc_2290_n540_1) );
  INVX1 INVX1_86 ( .A(_abc_2290_n542), .Y(_abc_2290_n552) );
  INVX1 INVX1_87 ( .A(_abc_2290_n533), .Y(_abc_2290_n555) );
  INVX1 INVX1_88 ( .A(_abc_2290_n526_1), .Y(_abc_2290_n557) );
  INVX1 INVX1_89 ( .A(_abc_2290_n560), .Y(_abc_2290_n561) );
  INVX1 INVX1_9 ( .A(tx_clk_divider_0_), .Y(_abc_2290_n163) );
  INVX1 INVX1_90 ( .A(_abc_2290_n562), .Y(_abc_2290_n563) );
  INVX1 INVX1_91 ( .A(rx_bits_remaining_2_), .Y(_abc_2290_n565) );
  INVX1 INVX1_92 ( .A(rx_bits_remaining_1_), .Y(_abc_2290_n566) );
  INVX1 INVX1_93 ( .A(rx_bits_remaining_3_), .Y(_abc_2290_n568) );
  INVX1 INVX1_94 ( .A(_abc_2290_n575), .Y(_abc_2290_n576) );
  INVX1 INVX1_95 ( .A(_abc_2290_n574), .Y(_abc_2290_n583) );
  INVX1 INVX1_96 ( .A(_abc_2290_n586), .Y(_abc_2290_n587) );
  INVX1 INVX1_97 ( .A(_abc_2290_n582), .Y(_abc_2290_n591) );
  INVX1 INVX1_98 ( .A(rx_bits_remaining_0_), .Y(_abc_2290_n597) );
  INVX1 INVX1_99 ( .A(_abc_2290_n599), .Y(_abc_2290_n600) );
  INVX2 INVX2_1 ( .A(rst), .Y(_abc_2290_n156_1) );
  INVX2 INVX2_2 ( .A(_abc_2290_n261), .Y(_abc_2290_n345) );
  INVX2 INVX2_3 ( .A(_abc_2290_n275), .Y(_abc_2290_n364) );
  INVX2 INVX2_4 ( .A(_abc_2290_n474), .Y(_abc_2290_n551) );
  OR2X2 OR2X2_1 ( .A(_abc_2290_n147_1), .B(recv_state_1_), .Y(is_receiving) );
  OR2X2 OR2X2_10 ( .A(_abc_2290_n178), .B(_abc_2290_n203), .Y(_abc_2290_n204) );
  OR2X2 OR2X2_100 ( .A(_abc_2290_n419), .B(rx_clk_divider_4_), .Y(_abc_2290_n487_1) );
  OR2X2 OR2X2_101 ( .A(_abc_2290_n403), .B(_abc_2290_n405), .Y(_abc_2290_n488) );
  OR2X2 OR2X2_102 ( .A(_abc_2290_n411), .B(_abc_2290_n412), .Y(_abc_2290_n495) );
  OR2X2 OR2X2_103 ( .A(_abc_2290_n505_1), .B(_abc_2290_n503), .Y(_abc_2290_n506) );
  OR2X2 OR2X2_104 ( .A(_abc_2290_n500_1), .B(_abc_2290_n501), .Y(_abc_2290_n509) );
  OR2X2 OR2X2_105 ( .A(_abc_2290_n519), .B(_abc_2290_n521), .Y(_abc_2290_n522_1) );
  OR2X2 OR2X2_106 ( .A(_abc_2290_n500_1), .B(_abc_2290_n520_1), .Y(_abc_2290_n525_1) );
  OR2X2 OR2X2_107 ( .A(_abc_2290_n528_1), .B(_abc_2290_n517), .Y(_abc_2290_n529_1) );
  OR2X2 OR2X2_108 ( .A(_abc_2290_n500_1), .B(_abc_2290_n514_1), .Y(_abc_2290_n532_1) );
  OR2X2 OR2X2_109 ( .A(_abc_2290_n535_1), .B(_abc_2290_n515), .Y(_abc_2290_n536) );
  OR2X2 OR2X2_11 ( .A(_abc_2290_n204), .B(tx_clk_divider_10_), .Y(_abc_2290_n205) );
  OR2X2 OR2X2_110 ( .A(_abc_2290_n503), .B(rx_countdown_3_), .Y(_abc_2290_n537_1) );
  OR2X2 OR2X2_111 ( .A(_abc_2290_n500_1), .B(_abc_2290_n515), .Y(_abc_2290_n541_1) );
  OR2X2 OR2X2_112 ( .A(_abc_2290_n547), .B(_abc_2290_n548_1), .Y(_abc_2290_n549) );
  OR2X2 OR2X2_113 ( .A(_abc_2290_n549), .B(_abc_2290_n512_1), .Y(rx_countdown_2__FF_INPUT) );
  OR2X2 OR2X2_114 ( .A(_abc_2290_n553), .B(_abc_2290_n479_1), .Y(rx_countdown_3__FF_INPUT) );
  OR2X2 OR2X2_115 ( .A(_abc_2290_n545), .B(_abc_2290_n456), .Y(_abc_2290_n559) );
  OR2X2 OR2X2_116 ( .A(_abc_2290_n564), .B(_abc_2290_n571), .Y(_abc_2290_n572) );
  OR2X2 OR2X2_117 ( .A(_abc_2290_n474), .B(_abc_2290_n578), .Y(_abc_2290_n579) );
  OR2X2 OR2X2_118 ( .A(_abc_2290_n577), .B(_abc_2290_n579), .Y(_abc_2290_n580) );
  OR2X2 OR2X2_119 ( .A(_abc_2290_n573), .B(_abc_2290_n580), .Y(recv_state_0__FF_INPUT) );
  OR2X2 OR2X2_12 ( .A(_abc_2290_n174_1), .B(_abc_2290_n199), .Y(_abc_2290_n207) );
  OR2X2 OR2X2_120 ( .A(_abc_2290_n545), .B(_abc_2290_n462), .Y(_abc_2290_n582) );
  OR2X2 OR2X2_121 ( .A(_abc_2290_n546_1), .B(_abc_2290_n583), .Y(_abc_2290_n584) );
  OR2X2 OR2X2_122 ( .A(_abc_2290_n575), .B(_abc_2290_n467), .Y(_abc_2290_n585) );
  OR2X2 OR2X2_123 ( .A(_abc_2290_n463), .B(_abc_2290_n578), .Y(_abc_2290_n589) );
  OR2X2 OR2X2_124 ( .A(_abc_2290_n588), .B(_abc_2290_n589), .Y(recv_state_1__FF_INPUT) );
  OR2X2 OR2X2_125 ( .A(_abc_2290_n591), .B(recv_state_0_), .Y(_abc_2290_n592) );
  OR2X2 OR2X2_126 ( .A(_abc_2290_n560), .B(_abc_2290_n574), .Y(_abc_2290_n594) );
  OR2X2 OR2X2_127 ( .A(_abc_2290_n593), .B(_abc_2290_n595), .Y(recv_state_2__FF_INPUT) );
  OR2X2 OR2X2_128 ( .A(_abc_2290_n601), .B(_abc_2290_n598), .Y(rx_bits_remaining_0__FF_INPUT) );
  OR2X2 OR2X2_129 ( .A(_abc_2290_n598), .B(rx_bits_remaining_1_), .Y(_abc_2290_n603) );
  OR2X2 OR2X2_13 ( .A(_abc_2290_n222_1), .B(_abc_2290_n223), .Y(_abc_2290_n224) );
  OR2X2 OR2X2_130 ( .A(_abc_2290_n546_1), .B(_abc_2290_n467), .Y(_abc_2290_n605) );
  OR2X2 OR2X2_131 ( .A(_abc_2290_n607), .B(_abc_2290_n464_1), .Y(_abc_2290_n608) );
  OR2X2 OR2X2_132 ( .A(_abc_2290_n610), .B(_abc_2290_n604), .Y(_abc_2290_n611) );
  OR2X2 OR2X2_133 ( .A(_abc_2290_n618), .B(_abc_2290_n616), .Y(_abc_2290_n619) );
  OR2X2 OR2X2_134 ( .A(_abc_2290_n620), .B(_abc_2290_n614), .Y(_abc_2290_n621) );
  OR2X2 OR2X2_135 ( .A(_abc_2290_n613), .B(_abc_2290_n621), .Y(rx_bits_remaining_2__FF_INPUT) );
  OR2X2 OR2X2_136 ( .A(_abc_2290_n626), .B(_abc_2290_n547), .Y(_abc_2290_n627) );
  OR2X2 OR2X2_137 ( .A(_abc_2290_n627), .B(_abc_2290_n625), .Y(rx_bits_remaining_3__FF_INPUT) );
  OR2X2 OR2X2_138 ( .A(_abc_2290_n165_1), .B(_abc_2290_n630), .Y(_abc_2290_n631) );
  OR2X2 OR2X2_139 ( .A(_abc_2290_n373), .B(_abc_2290_n275), .Y(_abc_2290_n632) );
  OR2X2 OR2X2_14 ( .A(_abc_2290_n210), .B(tx_countdown_5_), .Y(_abc_2290_n227_1) );
  OR2X2 OR2X2_140 ( .A(_abc_2290_n632), .B(_abc_2290_n631), .Y(tx_clk_divider_1__FF_INPUT) );
  OR2X2 OR2X2_141 ( .A(_abc_2290_n634), .B(tx_clk_divider_2_), .Y(_abc_2290_n635) );
  OR2X2 OR2X2_142 ( .A(_abc_2290_n636), .B(_abc_2290_n637), .Y(_abc_2290_n638) );
  OR2X2 OR2X2_143 ( .A(_abc_2290_n632), .B(_abc_2290_n638), .Y(tx_clk_divider_2__FF_INPUT) );
  OR2X2 OR2X2_144 ( .A(_abc_2290_n640), .B(_abc_2290_n166_1), .Y(_abc_2290_n641) );
  OR2X2 OR2X2_145 ( .A(_abc_2290_n275), .B(_abc_2290_n188), .Y(_abc_2290_n644) );
  OR2X2 OR2X2_146 ( .A(_abc_2290_n644), .B(_abc_2290_n643), .Y(_abc_2290_n645) );
  OR2X2 OR2X2_147 ( .A(_abc_2290_n373), .B(_abc_2290_n645), .Y(tx_clk_divider_4__FF_INPUT) );
  OR2X2 OR2X2_148 ( .A(_abc_2290_n649), .B(_abc_2290_n184), .Y(_abc_2290_n650) );
  OR2X2 OR2X2_149 ( .A(_abc_2290_n180), .B(_abc_2290_n275), .Y(_abc_2290_n654) );
  OR2X2 OR2X2_15 ( .A(_abc_2290_n230), .B(_abc_2290_n231), .Y(_abc_2290_n232_1) );
  OR2X2 OR2X2_150 ( .A(_abc_2290_n373), .B(_abc_2290_n654), .Y(tx_clk_divider_8__FF_INPUT) );
  OR2X2 OR2X2_151 ( .A(_abc_2290_n632), .B(_abc_2290_n658), .Y(tx_clk_divider_10__FF_INPUT) );
  OR2X2 OR2X2_152 ( .A(_abc_2290_n402), .B(_abc_2290_n661), .Y(_abc_2290_n662) );
  OR2X2 OR2X2_153 ( .A(_abc_2290_n474), .B(_abc_2290_n662), .Y(_abc_2290_n663) );
  OR2X2 OR2X2_154 ( .A(_abc_2290_n448), .B(_abc_2290_n663), .Y(rx_clk_divider_1__FF_INPUT) );
  OR2X2 OR2X2_155 ( .A(_abc_2290_n665), .B(_abc_2290_n666), .Y(_abc_2290_n667) );
  OR2X2 OR2X2_156 ( .A(_abc_2290_n474), .B(_abc_2290_n667), .Y(_abc_2290_n668) );
  OR2X2 OR2X2_157 ( .A(_abc_2290_n448), .B(_abc_2290_n668), .Y(rx_clk_divider_2__FF_INPUT) );
  OR2X2 OR2X2_158 ( .A(_abc_2290_n671), .B(_abc_2290_n403), .Y(_abc_2290_n672) );
  OR2X2 OR2X2_159 ( .A(_abc_2290_n474), .B(_abc_2290_n674), .Y(_abc_2290_n675) );
  OR2X2 OR2X2_16 ( .A(_abc_2290_n210), .B(tx_countdown_2_), .Y(_abc_2290_n235) );
  OR2X2 OR2X2_160 ( .A(_abc_2290_n448), .B(_abc_2290_n675), .Y(rx_clk_divider_4__FF_INPUT) );
  OR2X2 OR2X2_161 ( .A(_abc_2290_n500_1), .B(_abc_2290_n683), .Y(_abc_2290_n684) );
  OR2X2 OR2X2_162 ( .A(_abc_2290_n684), .B(_abc_2290_n474), .Y(rx_clk_divider_8__FF_INPUT) );
  OR2X2 OR2X2_163 ( .A(_abc_2290_n500_1), .B(_abc_2290_n688), .Y(_abc_2290_n689) );
  OR2X2 OR2X2_164 ( .A(_abc_2290_n689), .B(_abc_2290_n474), .Y(rx_clk_divider_10__FF_INPUT) );
  OR2X2 OR2X2_165 ( .A(_abc_2290_n548_1), .B(\rx_byte[0] ), .Y(_abc_2290_n691) );
  OR2X2 OR2X2_166 ( .A(_abc_2290_n548_1), .B(\rx_byte[1] ), .Y(_abc_2290_n696) );
  OR2X2 OR2X2_167 ( .A(_abc_2290_n548_1), .B(\rx_byte[2] ), .Y(_abc_2290_n701) );
  OR2X2 OR2X2_168 ( .A(_abc_2290_n548_1), .B(\rx_byte[3] ), .Y(_abc_2290_n706) );
  OR2X2 OR2X2_169 ( .A(_abc_2290_n548_1), .B(\rx_byte[4] ), .Y(_abc_2290_n711) );
  OR2X2 OR2X2_17 ( .A(_abc_2290_n236), .B(tx_countdown_4_), .Y(_abc_2290_n237_1) );
  OR2X2 OR2X2_170 ( .A(_abc_2290_n548_1), .B(\rx_byte[5] ), .Y(_abc_2290_n716) );
  OR2X2 OR2X2_171 ( .A(_abc_2290_n548_1), .B(\rx_byte[6] ), .Y(_abc_2290_n721) );
  OR2X2 OR2X2_172 ( .A(_abc_2290_n548_1), .B(\rx_byte[7] ), .Y(_abc_2290_n728) );
  OR2X2 OR2X2_18 ( .A(_abc_2290_n237_1), .B(_abc_2290_n228), .Y(_abc_2290_n238) );
  OR2X2 OR2X2_19 ( .A(_abc_2290_n210), .B(tx_countdown_0_), .Y(_abc_2290_n240) );
  OR2X2 OR2X2_2 ( .A(tx_state_1_), .B(tx_state_0_), .Y(is_transmitting) );
  OR2X2 OR2X2_20 ( .A(_abc_2290_n241_1), .B(_abc_2290_n239), .Y(_abc_2290_n242) );
  OR2X2 OR2X2_21 ( .A(_abc_2290_n245_1), .B(_abc_2290_n246), .Y(_abc_2290_n247) );
  OR2X2 OR2X2_22 ( .A(_abc_2290_n210), .B(tx_countdown_3_), .Y(_abc_2290_n250_1) );
  OR2X2 OR2X2_23 ( .A(_abc_2290_n252), .B(_abc_2290_n253), .Y(_abc_2290_n254) );
  OR2X2 OR2X2_24 ( .A(_abc_2290_n210), .B(tx_countdown_1_), .Y(_abc_2290_n257_1) );
  OR2X2 OR2X2_25 ( .A(_abc_2290_n251), .B(_abc_2290_n258_1), .Y(_abc_2290_n259) );
  OR2X2 OR2X2_26 ( .A(_abc_2290_n259), .B(_abc_2290_n243), .Y(_abc_2290_n260) );
  OR2X2 OR2X2_27 ( .A(_abc_2290_n260), .B(_abc_2290_n238), .Y(_abc_2290_n261) );
  OR2X2 OR2X2_28 ( .A(_abc_2290_n265_1), .B(tx_bits_remaining_2_), .Y(_abc_2290_n266) );
  OR2X2 OR2X2_29 ( .A(_abc_2290_n266), .B(tx_bits_remaining_3_), .Y(_abc_2290_n267_1) );
  OR2X2 OR2X2_3 ( .A(tx_clk_divider_6_), .B(tx_clk_divider_7_), .Y(_abc_2290_n171) );
  OR2X2 OR2X2_30 ( .A(_abc_2290_n261), .B(_abc_2290_n268_1), .Y(_abc_2290_n269) );
  OR2X2 OR2X2_31 ( .A(_abc_2290_n279), .B(_abc_2290_n277), .Y(_abc_2290_n280) );
  OR2X2 OR2X2_32 ( .A(_abc_2290_n281_1), .B(_abc_2290_n276), .Y(_abc_2290_n282) );
  OR2X2 OR2X2_33 ( .A(_abc_2290_n284), .B(_abc_2290_n282), .Y(_abc_2290_n285) );
  OR2X2 OR2X2_34 ( .A(_abc_2290_n285), .B(_abc_2290_n272), .Y(tx_data_0__FF_INPUT) );
  OR2X2 OR2X2_35 ( .A(_abc_2290_n289), .B(_abc_2290_n288), .Y(_abc_2290_n290) );
  OR2X2 OR2X2_36 ( .A(_abc_2290_n291), .B(_abc_2290_n290), .Y(_abc_2290_n292) );
  OR2X2 OR2X2_37 ( .A(_abc_2290_n292), .B(_abc_2290_n287), .Y(tx_data_1__FF_INPUT) );
  OR2X2 OR2X2_38 ( .A(_abc_2290_n296), .B(_abc_2290_n295), .Y(_abc_2290_n297) );
  OR2X2 OR2X2_39 ( .A(_abc_2290_n298), .B(_abc_2290_n297), .Y(_abc_2290_n299_1) );
  OR2X2 OR2X2_4 ( .A(_abc_2290_n176), .B(_abc_2290_n171), .Y(_abc_2290_n177) );
  OR2X2 OR2X2_40 ( .A(_abc_2290_n299_1), .B(_abc_2290_n294), .Y(tx_data_2__FF_INPUT) );
  OR2X2 OR2X2_41 ( .A(_abc_2290_n303), .B(_abc_2290_n302), .Y(_abc_2290_n304) );
  OR2X2 OR2X2_42 ( .A(_abc_2290_n305), .B(_abc_2290_n304), .Y(_abc_2290_n306) );
  OR2X2 OR2X2_43 ( .A(_abc_2290_n306), .B(_abc_2290_n301), .Y(tx_data_3__FF_INPUT) );
  OR2X2 OR2X2_44 ( .A(_abc_2290_n310), .B(_abc_2290_n309), .Y(_abc_2290_n311) );
  OR2X2 OR2X2_45 ( .A(_abc_2290_n312_1), .B(_abc_2290_n311), .Y(_abc_2290_n313) );
  OR2X2 OR2X2_46 ( .A(_abc_2290_n313), .B(_abc_2290_n308), .Y(tx_data_4__FF_INPUT) );
  OR2X2 OR2X2_47 ( .A(_abc_2290_n317), .B(_abc_2290_n316), .Y(_abc_2290_n318) );
  OR2X2 OR2X2_48 ( .A(_abc_2290_n319_1), .B(_abc_2290_n318), .Y(_abc_2290_n320) );
  OR2X2 OR2X2_49 ( .A(_abc_2290_n320), .B(_abc_2290_n315), .Y(tx_data_5__FF_INPUT) );
  OR2X2 OR2X2_5 ( .A(_abc_2290_n177), .B(_abc_2290_n175_1), .Y(_abc_2290_n178) );
  OR2X2 OR2X2_50 ( .A(_abc_2290_n323_1), .B(_abc_2290_n322), .Y(_abc_2290_n324) );
  OR2X2 OR2X2_51 ( .A(_abc_2290_n270_1), .B(tx_data_6_), .Y(_abc_2290_n325) );
  OR2X2 OR2X2_52 ( .A(_abc_2290_n283), .B(_abc_2290_n326), .Y(_abc_2290_n327) );
  OR2X2 OR2X2_53 ( .A(_abc_2290_n328), .B(_abc_2290_n324), .Y(tx_data_6__FF_INPUT) );
  OR2X2 OR2X2_54 ( .A(_abc_2290_n283), .B(_abc_2290_n280), .Y(_abc_2290_n331) );
  OR2X2 OR2X2_55 ( .A(_abc_2290_n332), .B(_abc_2290_n330), .Y(tx_data_7__FF_INPUT) );
  OR2X2 OR2X2_56 ( .A(_abc_2290_n270_1), .B(tx_bits_remaining_0_), .Y(_abc_2290_n334) );
  OR2X2 OR2X2_57 ( .A(_abc_2290_n261), .B(_abc_2290_n263), .Y(_abc_2290_n335) );
  OR2X2 OR2X2_58 ( .A(_abc_2290_n336), .B(_abc_2290_n337), .Y(_abc_2290_n338) );
  OR2X2 OR2X2_59 ( .A(_abc_2290_n263), .B(tx_bits_remaining_1_), .Y(_abc_2290_n340) );
  OR2X2 OR2X2_6 ( .A(_abc_2290_n174_1), .B(_abc_2290_n179_1), .Y(_abc_2290_n180) );
  OR2X2 OR2X2_60 ( .A(_abc_2290_n262), .B(tx_bits_remaining_0_), .Y(_abc_2290_n341) );
  OR2X2 OR2X2_61 ( .A(_abc_2290_n261), .B(_abc_2290_n343), .Y(_abc_2290_n344_1) );
  OR2X2 OR2X2_62 ( .A(_abc_2290_n345), .B(tx_bits_remaining_1_), .Y(_abc_2290_n346) );
  OR2X2 OR2X2_63 ( .A(_abc_2290_n348), .B(_abc_2290_n349), .Y(tx_bits_remaining_1__FF_INPUT) );
  OR2X2 OR2X2_64 ( .A(_abc_2290_n261), .B(_abc_2290_n265_1), .Y(_abc_2290_n355) );
  OR2X2 OR2X2_65 ( .A(_abc_2290_n356), .B(_abc_2290_n280), .Y(_abc_2290_n357_1) );
  OR2X2 OR2X2_66 ( .A(_abc_2290_n358), .B(_abc_2290_n354), .Y(tx_bits_remaining_2__FF_INPUT) );
  OR2X2 OR2X2_67 ( .A(_abc_2290_n362), .B(_abc_2290_n275), .Y(tx_bits_remaining_3__FF_INPUT) );
  OR2X2 OR2X2_68 ( .A(_abc_2290_n236), .B(_abc_2290_n275), .Y(_abc_2290_n367) );
  OR2X2 OR2X2_69 ( .A(_abc_2290_n271_1), .B(_abc_2290_n367), .Y(tx_countdown_2__FF_INPUT) );
  OR2X2 OR2X2_7 ( .A(_abc_2290_n184), .B(_abc_2290_n182), .Y(_abc_2290_n185_1) );
  OR2X2 OR2X2_70 ( .A(_abc_2290_n369), .B(_abc_2290_n251), .Y(_abc_2290_n370) );
  OR2X2 OR2X2_71 ( .A(_abc_2290_n378), .B(_abc_2290_n376), .Y(_abc_2290_n379) );
  OR2X2 OR2X2_72 ( .A(_abc_2290_n385), .B(_abc_2290_n275), .Y(tx_state_0__FF_INPUT) );
  OR2X2 OR2X2_73 ( .A(_abc_2290_n382_1), .B(_abc_2290_n277), .Y(_abc_2290_n387) );
  OR2X2 OR2X2_74 ( .A(_abc_2290_n261), .B(_abc_2290_n157_1), .Y(_abc_2290_n388) );
  OR2X2 OR2X2_75 ( .A(_abc_2290_n269), .B(tx_data_0_), .Y(_abc_2290_n390) );
  OR2X2 OR2X2_76 ( .A(_abc_2290_n345), .B(tx), .Y(_abc_2290_n391) );
  OR2X2 OR2X2_77 ( .A(_abc_2290_n393), .B(_abc_2290_n394), .Y(tx_out_FF_INPUT) );
  OR2X2 OR2X2_78 ( .A(rx_clk_divider_3_), .B(rx_clk_divider_2_), .Y(_abc_2290_n417) );
  OR2X2 OR2X2_79 ( .A(rx_clk_divider_0_), .B(rx_clk_divider_1_), .Y(_abc_2290_n418) );
  OR2X2 OR2X2_8 ( .A(_abc_2290_n188), .B(_abc_2290_n167), .Y(_abc_2290_n189_1) );
  OR2X2 OR2X2_80 ( .A(_abc_2290_n417), .B(_abc_2290_n418), .Y(_abc_2290_n419) );
  OR2X2 OR2X2_81 ( .A(rx_clk_divider_5_), .B(rx_clk_divider_4_), .Y(_abc_2290_n420) );
  OR2X2 OR2X2_82 ( .A(rx_clk_divider_6_), .B(rx_clk_divider_7_), .Y(_abc_2290_n421) );
  OR2X2 OR2X2_83 ( .A(_abc_2290_n420), .B(_abc_2290_n421), .Y(_abc_2290_n422) );
  OR2X2 OR2X2_84 ( .A(_abc_2290_n419), .B(_abc_2290_n422), .Y(_abc_2290_n423_1) );
  OR2X2 OR2X2_85 ( .A(_abc_2290_n423_1), .B(rx_clk_divider_8_), .Y(_abc_2290_n424) );
  OR2X2 OR2X2_86 ( .A(_abc_2290_n425_1), .B(_abc_2290_n413), .Y(_abc_2290_n426) );
  OR2X2 OR2X2_87 ( .A(_abc_2290_n419), .B(_abc_2290_n420), .Y(_abc_2290_n428_1) );
  OR2X2 OR2X2_88 ( .A(_abc_2290_n428_1), .B(rx_clk_divider_6_), .Y(_abc_2290_n429) );
  OR2X2 OR2X2_89 ( .A(_abc_2290_n430), .B(_abc_2290_n408), .Y(_abc_2290_n431) );
  OR2X2 OR2X2_9 ( .A(_abc_2290_n201), .B(_abc_2290_n198), .Y(_abc_2290_n202_1) );
  OR2X2 OR2X2_90 ( .A(_abc_2290_n433), .B(_abc_2290_n407), .Y(_abc_2290_n434) );
  OR2X2 OR2X2_91 ( .A(_abc_2290_n436), .B(_abc_2290_n404_1), .Y(_abc_2290_n437) );
  OR2X2 OR2X2_92 ( .A(_abc_2290_n448), .B(_abc_2290_n396), .Y(_abc_2290_n449_1) );
  OR2X2 OR2X2_93 ( .A(_abc_2290_n455), .B(_abc_2290_n457), .Y(_abc_2290_n458) );
  OR2X2 OR2X2_94 ( .A(_abc_2290_n461), .B(_abc_2290_n469_1), .Y(_abc_2290_n470) );
  OR2X2 OR2X2_95 ( .A(_abc_2290_n470), .B(_abc_2290_n458), .Y(_abc_2290_n471) );
  OR2X2 OR2X2_96 ( .A(_abc_2290_n475), .B(_abc_2290_n477_1), .Y(_abc_2290_n478) );
  OR2X2 OR2X2_97 ( .A(_abc_2290_n481), .B(_abc_2290_n474), .Y(rx_countdown_1__FF_INPUT) );
  OR2X2 OR2X2_98 ( .A(_abc_2290_n415), .B(_abc_2290_n439), .Y(_abc_2290_n483) );
  OR2X2 OR2X2_99 ( .A(_abc_2290_n416), .B(rx_clk_divider_10_), .Y(_abc_2290_n484_1) );
endmodule