
module cpu8080(\data[0] , \data[1] , \data[2] , \data[3] , \data[4] , \data[5] , \data[6] , \data[7] , intr, waitr, reset, clock, \addr[0] , \addr[1] , \addr[2] , \addr[3] , \addr[4] , \addr[5] , \addr[6] , \addr[7] , \addr[8] , \addr[9] , \addr[10] , \addr[11] , \addr[12] , \addr[13] , \addr[14] , \addr[15] , readmem, writemem, readio, writeio, inta);
  wire _abc_36783_n3361;
  wire _abc_36783_n3364;
  wire _abc_36783_n3367;
  wire _abc_36783_n3370;
  wire _abc_36783_n3373;
  wire _abc_36783_n3376;
  wire _abc_36783_n3379;
  wire _abc_36783_n3382;
  wire _abc_36783_n3435;
  wire _abc_36783_n3438;
  wire _abc_36783_n3441;
  wire _abc_36783_n3444;
  wire _abc_36783_n3447;
  wire _abc_36783_n3450;
  wire _abc_36783_n3453;
  wire _abc_36783_n3456;
  wire _abc_36783_n3520;
  wire _abc_36783_n3523;
  wire _abc_36783_n3526;
  wire _abc_36783_n3529;
  wire _abc_36783_n3532;
  wire _abc_36783_n3535;
  wire _abc_36783_n3538;
  wire _abc_36783_n3541;
  wire _abc_36783_n3554;
  wire _abc_36783_n3557;
  wire _abc_36783_n3560;
  wire _abc_36783_n3563;
  wire _abc_36783_n3566;
  wire _abc_36783_n3569;
  wire _abc_36783_n3572;
  wire _abc_36783_n3575;
  wire _abc_36783_n3638;
  wire _abc_36783_n3640;
  wire _abc_36783_n3642;
  wire _abc_36783_n3644;
  wire _abc_36783_n3646;
  wire _abc_36783_n3648;
  wire _abc_36783_n3650;
  wire _abc_36783_n3652;
  wire _abc_36783_n3731;
  wire _abc_36783_n3732;
  wire _abc_36783_n3733;
  wire _abc_36783_n3734;
  wire _abc_36783_n3735;
  wire _abc_36783_n3736;
  wire _abc_36783_n3737;
  wire _abc_36783_n3738;
  wire _abc_36783_n4531;
  wire _abc_36783_n4532;
  wire _abc_36783_n4533;
  wire _abc_36783_n4534;
  wire _abc_36783_n4535;
  wire _abc_36783_n4536;
  wire _abc_36783_n4537;
  wire _abc_36783_n4538;
  wire _abc_36783_n4579;
  wire _abc_36783_n4580;
  wire _abc_36783_n4581;
  wire _abc_36783_n4582;
  wire _abc_36783_n4583;
  wire _abc_36783_n4584;
  wire _abc_36783_n4585;
  wire _abc_36783_n4586;
  wire _abc_36783_n4644;
  wire _abc_36783_n4645;
  wire _abc_36783_n4646;
  wire _abc_36783_n4647;
  wire _abc_36783_n4648;
  wire _abc_36783_n4649;
  wire _abc_42016_n1000;
  wire _abc_42016_n1001_1;
  wire _abc_42016_n1002;
  wire _abc_42016_n1003;
  wire _abc_42016_n1004;
  wire _abc_42016_n1005;
  wire _abc_42016_n1006;
  wire _abc_42016_n1007;
  wire _abc_42016_n1008;
  wire _abc_42016_n1009;
  wire _abc_42016_n1010;
  wire _abc_42016_n1011;
  wire _abc_42016_n1012;
  wire _abc_42016_n1013;
  wire _abc_42016_n1014;
  wire _abc_42016_n1015;
  wire _abc_42016_n1016;
  wire _abc_42016_n1017;
  wire _abc_42016_n1018;
  wire _abc_42016_n1019;
  wire _abc_42016_n1020;
  wire _abc_42016_n1021;
  wire _abc_42016_n1022;
  wire _abc_42016_n1023;
  wire _abc_42016_n1024;
  wire _abc_42016_n1025;
  wire _abc_42016_n1026;
  wire _abc_42016_n1027;
  wire _abc_42016_n1028;
  wire _abc_42016_n1029;
  wire _abc_42016_n1030;
  wire _abc_42016_n1031_1;
  wire _abc_42016_n1032;
  wire _abc_42016_n1033;
  wire _abc_42016_n1034;
  wire _abc_42016_n1035;
  wire _abc_42016_n1036;
  wire _abc_42016_n1037;
  wire _abc_42016_n1038;
  wire _abc_42016_n1039;
  wire _abc_42016_n1040;
  wire _abc_42016_n1041;
  wire _abc_42016_n1042;
  wire _abc_42016_n1043;
  wire _abc_42016_n1044;
  wire _abc_42016_n1045;
  wire _abc_42016_n1046;
  wire _abc_42016_n1047_1;
  wire _abc_42016_n1048;
  wire _abc_42016_n1049;
  wire _abc_42016_n1050;
  wire _abc_42016_n1051;
  wire _abc_42016_n1052;
  wire _abc_42016_n1053;
  wire _abc_42016_n1055;
  wire _abc_42016_n1056;
  wire _abc_42016_n1057;
  wire _abc_42016_n1058;
  wire _abc_42016_n1059;
  wire _abc_42016_n1060;
  wire _abc_42016_n1061;
  wire _abc_42016_n1062;
  wire _abc_42016_n1063;
  wire _abc_42016_n1064;
  wire _abc_42016_n1065;
  wire _abc_42016_n1066;
  wire _abc_42016_n1067;
  wire _abc_42016_n1068;
  wire _abc_42016_n1069;
  wire _abc_42016_n1070_1;
  wire _abc_42016_n1071;
  wire _abc_42016_n1072;
  wire _abc_42016_n1073_1;
  wire _abc_42016_n1074;
  wire _abc_42016_n1075;
  wire _abc_42016_n1076;
  wire _abc_42016_n1077;
  wire _abc_42016_n1078;
  wire _abc_42016_n1079;
  wire _abc_42016_n1080;
  wire _abc_42016_n1081;
  wire _abc_42016_n1082;
  wire _abc_42016_n1083;
  wire _abc_42016_n1084;
  wire _abc_42016_n1085;
  wire _abc_42016_n1086;
  wire _abc_42016_n1087;
  wire _abc_42016_n1088;
  wire _abc_42016_n1089;
  wire _abc_42016_n1090;
  wire _abc_42016_n1091;
  wire _abc_42016_n1092;
  wire _abc_42016_n1094;
  wire _abc_42016_n1095;
  wire _abc_42016_n1096;
  wire _abc_42016_n1097;
  wire _abc_42016_n1098;
  wire _abc_42016_n1099;
  wire _abc_42016_n1100;
  wire _abc_42016_n1101_1;
  wire _abc_42016_n1102;
  wire _abc_42016_n1103_1;
  wire _abc_42016_n1104_1;
  wire _abc_42016_n1105;
  wire _abc_42016_n1106_1;
  wire _abc_42016_n1107_1;
  wire _abc_42016_n1108;
  wire _abc_42016_n1109;
  wire _abc_42016_n1110_1;
  wire _abc_42016_n1111_1;
  wire _abc_42016_n1112;
  wire _abc_42016_n1113_1;
  wire _abc_42016_n1114_1;
  wire _abc_42016_n1115;
  wire _abc_42016_n1116;
  wire _abc_42016_n1117;
  wire _abc_42016_n1118;
  wire _abc_42016_n1119;
  wire _abc_42016_n1120;
  wire _abc_42016_n1121_1;
  wire _abc_42016_n1122;
  wire _abc_42016_n1123;
  wire _abc_42016_n1124;
  wire _abc_42016_n1125;
  wire _abc_42016_n1126;
  wire _abc_42016_n1127;
  wire _abc_42016_n1128;
  wire _abc_42016_n1129;
  wire _abc_42016_n1130;
  wire _abc_42016_n1131;
  wire _abc_42016_n1132;
  wire _abc_42016_n1133;
  wire _abc_42016_n1134;
  wire _abc_42016_n1136;
  wire _abc_42016_n1137;
  wire _abc_42016_n1138;
  wire _abc_42016_n1139;
  wire _abc_42016_n1140;
  wire _abc_42016_n1141;
  wire _abc_42016_n1142;
  wire _abc_42016_n1143;
  wire _abc_42016_n1144;
  wire _abc_42016_n1145;
  wire _abc_42016_n1146_1;
  wire _abc_42016_n1147_1;
  wire _abc_42016_n1148;
  wire _abc_42016_n1149_1;
  wire _abc_42016_n1150;
  wire _abc_42016_n1151;
  wire _abc_42016_n1152;
  wire _abc_42016_n1153;
  wire _abc_42016_n1154;
  wire _abc_42016_n1155;
  wire _abc_42016_n1156;
  wire _abc_42016_n1157;
  wire _abc_42016_n1158;
  wire _abc_42016_n1159;
  wire _abc_42016_n1160;
  wire _abc_42016_n1161;
  wire _abc_42016_n1162;
  wire _abc_42016_n1163;
  wire _abc_42016_n1164;
  wire _abc_42016_n1165;
  wire _abc_42016_n1166;
  wire _abc_42016_n1167;
  wire _abc_42016_n1168;
  wire _abc_42016_n1169;
  wire _abc_42016_n1170;
  wire _abc_42016_n1171_1;
  wire _abc_42016_n1172_1;
  wire _abc_42016_n1173;
  wire _abc_42016_n1174_1;
  wire _abc_42016_n1175;
  wire _abc_42016_n1176;
  wire _abc_42016_n1177;
  wire _abc_42016_n1179;
  wire _abc_42016_n1180;
  wire _abc_42016_n1181;
  wire _abc_42016_n1182;
  wire _abc_42016_n1183;
  wire _abc_42016_n1184;
  wire _abc_42016_n1185;
  wire _abc_42016_n1186;
  wire _abc_42016_n1187;
  wire _abc_42016_n1188;
  wire _abc_42016_n1189;
  wire _abc_42016_n1190;
  wire _abc_42016_n1191;
  wire _abc_42016_n1192;
  wire _abc_42016_n1193;
  wire _abc_42016_n1194;
  wire _abc_42016_n1195;
  wire _abc_42016_n1196_1;
  wire _abc_42016_n1197_1;
  wire _abc_42016_n1198;
  wire _abc_42016_n1199_1;
  wire _abc_42016_n1200;
  wire _abc_42016_n1201;
  wire _abc_42016_n1202;
  wire _abc_42016_n1203;
  wire _abc_42016_n1204;
  wire _abc_42016_n1205;
  wire _abc_42016_n1206;
  wire _abc_42016_n1207;
  wire _abc_42016_n1208;
  wire _abc_42016_n1209;
  wire _abc_42016_n1210;
  wire _abc_42016_n1211;
  wire _abc_42016_n1212;
  wire _abc_42016_n1213;
  wire _abc_42016_n1214;
  wire _abc_42016_n1215;
  wire _abc_42016_n1216;
  wire _abc_42016_n1217;
  wire _abc_42016_n1218;
  wire _abc_42016_n1219;
  wire _abc_42016_n1220;
  wire _abc_42016_n1221_1;
  wire _abc_42016_n1223;
  wire _abc_42016_n1224_1;
  wire _abc_42016_n1225;
  wire _abc_42016_n1226;
  wire _abc_42016_n1227;
  wire _abc_42016_n1228;
  wire _abc_42016_n1229;
  wire _abc_42016_n1230;
  wire _abc_42016_n1231;
  wire _abc_42016_n1232;
  wire _abc_42016_n1233;
  wire _abc_42016_n1234;
  wire _abc_42016_n1235;
  wire _abc_42016_n1236;
  wire _abc_42016_n1237;
  wire _abc_42016_n1238;
  wire _abc_42016_n1239;
  wire _abc_42016_n1240;
  wire _abc_42016_n1241;
  wire _abc_42016_n1242;
  wire _abc_42016_n1243;
  wire _abc_42016_n1244;
  wire _abc_42016_n1245;
  wire _abc_42016_n1246;
  wire _abc_42016_n1247_1;
  wire _abc_42016_n1248_1;
  wire _abc_42016_n1249;
  wire _abc_42016_n1250_1;
  wire _abc_42016_n1251;
  wire _abc_42016_n1252;
  wire _abc_42016_n1253;
  wire _abc_42016_n1254;
  wire _abc_42016_n1255;
  wire _abc_42016_n1256;
  wire _abc_42016_n1257;
  wire _abc_42016_n1259;
  wire _abc_42016_n1260;
  wire _abc_42016_n1261;
  wire _abc_42016_n1262;
  wire _abc_42016_n1263;
  wire _abc_42016_n1264;
  wire _abc_42016_n1265;
  wire _abc_42016_n1266;
  wire _abc_42016_n1267;
  wire _abc_42016_n1268;
  wire _abc_42016_n1269;
  wire _abc_42016_n1270;
  wire _abc_42016_n1271_1;
  wire _abc_42016_n1272_1;
  wire _abc_42016_n1273;
  wire _abc_42016_n1274_1;
  wire _abc_42016_n1275;
  wire _abc_42016_n1276;
  wire _abc_42016_n1277;
  wire _abc_42016_n1278;
  wire _abc_42016_n1279;
  wire _abc_42016_n1280;
  wire _abc_42016_n1281;
  wire _abc_42016_n1282;
  wire _abc_42016_n1283;
  wire _abc_42016_n1284;
  wire _abc_42016_n1285;
  wire _abc_42016_n1286;
  wire _abc_42016_n1287;
  wire _abc_42016_n1288;
  wire _abc_42016_n1289;
  wire _abc_42016_n1290;
  wire _abc_42016_n1291;
  wire _abc_42016_n1292;
  wire _abc_42016_n1293;
  wire _abc_42016_n1294;
  wire _abc_42016_n1295;
  wire _abc_42016_n1296_1;
  wire _abc_42016_n1297_1;
  wire _abc_42016_n1298;
  wire _abc_42016_n1299_1;
  wire _abc_42016_n1300;
  wire _abc_42016_n1302;
  wire _abc_42016_n1303;
  wire _abc_42016_n1304;
  wire _abc_42016_n1305;
  wire _abc_42016_n1306;
  wire _abc_42016_n1307;
  wire _abc_42016_n1308;
  wire _abc_42016_n1309;
  wire _abc_42016_n1310;
  wire _abc_42016_n1311;
  wire _abc_42016_n1312;
  wire _abc_42016_n1313;
  wire _abc_42016_n1314;
  wire _abc_42016_n1315;
  wire _abc_42016_n1316;
  wire _abc_42016_n1317;
  wire _abc_42016_n1318;
  wire _abc_42016_n1319;
  wire _abc_42016_n1320;
  wire _abc_42016_n1321_1;
  wire _abc_42016_n1322;
  wire _abc_42016_n1323;
  wire _abc_42016_n1324;
  wire _abc_42016_n1325;
  wire _abc_42016_n1326;
  wire _abc_42016_n1327_1;
  wire _abc_42016_n1328;
  wire _abc_42016_n1329_1;
  wire _abc_42016_n1330;
  wire _abc_42016_n1331_1;
  wire _abc_42016_n1332;
  wire _abc_42016_n1333_1;
  wire _abc_42016_n1334;
  wire _abc_42016_n1335_1;
  wire _abc_42016_n1336;
  wire _abc_42016_n1337_1;
  wire _abc_42016_n1338;
  wire _abc_42016_n1339_1;
  wire _abc_42016_n1340;
  wire _abc_42016_n1341_1;
  wire _abc_42016_n1342;
  wire _abc_42016_n1344;
  wire _abc_42016_n1345;
  wire _abc_42016_n1346;
  wire _abc_42016_n1347;
  wire _abc_42016_n1348;
  wire _abc_42016_n1349;
  wire _abc_42016_n1350;
  wire _abc_42016_n1351;
  wire _abc_42016_n1352;
  wire _abc_42016_n1353;
  wire _abc_42016_n1354;
  wire _abc_42016_n1355;
  wire _abc_42016_n1356;
  wire _abc_42016_n1357;
  wire _abc_42016_n1358;
  wire _abc_42016_n1359;
  wire _abc_42016_n1360;
  wire _abc_42016_n1361;
  wire _abc_42016_n1362;
  wire _abc_42016_n1363;
  wire _abc_42016_n1364;
  wire _abc_42016_n1365;
  wire _abc_42016_n1366;
  wire _abc_42016_n1367;
  wire _abc_42016_n1368;
  wire _abc_42016_n1369;
  wire _abc_42016_n1370;
  wire _abc_42016_n1371;
  wire _abc_42016_n1372;
  wire _abc_42016_n1373;
  wire _abc_42016_n1374;
  wire _abc_42016_n1375;
  wire _abc_42016_n1376;
  wire _abc_42016_n1377;
  wire _abc_42016_n1378;
  wire _abc_42016_n1379;
  wire _abc_42016_n1380;
  wire _abc_42016_n1381;
  wire _abc_42016_n1382;
  wire _abc_42016_n1383;
  wire _abc_42016_n1384;
  wire _abc_42016_n1385;
  wire _abc_42016_n1386_1;
  wire _abc_42016_n1387;
  wire _abc_42016_n1388;
  wire _abc_42016_n1389;
  wire _abc_42016_n1390;
  wire _abc_42016_n1391;
  wire _abc_42016_n1392;
  wire _abc_42016_n1393;
  wire _abc_42016_n1394;
  wire _abc_42016_n1395;
  wire _abc_42016_n1396;
  wire _abc_42016_n1397;
  wire _abc_42016_n1398;
  wire _abc_42016_n1399;
  wire _abc_42016_n1400;
  wire _abc_42016_n1401;
  wire _abc_42016_n1402;
  wire _abc_42016_n1403;
  wire _abc_42016_n1404;
  wire _abc_42016_n1405;
  wire _abc_42016_n1406;
  wire _abc_42016_n1407;
  wire _abc_42016_n1408;
  wire _abc_42016_n1409;
  wire _abc_42016_n1410_1;
  wire _abc_42016_n1411;
  wire _abc_42016_n1412;
  wire _abc_42016_n1413;
  wire _abc_42016_n1414;
  wire _abc_42016_n1415;
  wire _abc_42016_n1416;
  wire _abc_42016_n1417;
  wire _abc_42016_n1419;
  wire _abc_42016_n1420;
  wire _abc_42016_n1421;
  wire _abc_42016_n1422;
  wire _abc_42016_n1423;
  wire _abc_42016_n1424;
  wire _abc_42016_n1425;
  wire _abc_42016_n1426;
  wire _abc_42016_n1427;
  wire _abc_42016_n1428;
  wire _abc_42016_n1429;
  wire _abc_42016_n1430;
  wire _abc_42016_n1431;
  wire _abc_42016_n1432;
  wire _abc_42016_n1433;
  wire _abc_42016_n1434;
  wire _abc_42016_n1435;
  wire _abc_42016_n1436;
  wire _abc_42016_n1437;
  wire _abc_42016_n1438;
  wire _abc_42016_n1439_1;
  wire _abc_42016_n1440;
  wire _abc_42016_n1441;
  wire _abc_42016_n1442;
  wire _abc_42016_n1443;
  wire _abc_42016_n1445;
  wire _abc_42016_n1446;
  wire _abc_42016_n1447;
  wire _abc_42016_n1448;
  wire _abc_42016_n1449;
  wire _abc_42016_n1450;
  wire _abc_42016_n1451;
  wire _abc_42016_n1452;
  wire _abc_42016_n1453;
  wire _abc_42016_n1454;
  wire _abc_42016_n1455;
  wire _abc_42016_n1456;
  wire _abc_42016_n1457;
  wire _abc_42016_n1458;
  wire _abc_42016_n1459;
  wire _abc_42016_n1460;
  wire _abc_42016_n1461;
  wire _abc_42016_n1462;
  wire _abc_42016_n1463;
  wire _abc_42016_n1464;
  wire _abc_42016_n1465_1;
  wire _abc_42016_n1466;
  wire _abc_42016_n1467;
  wire _abc_42016_n1468;
  wire _abc_42016_n1469;
  wire _abc_42016_n1470;
  wire _abc_42016_n1471;
  wire _abc_42016_n1472;
  wire _abc_42016_n1474;
  wire _abc_42016_n1475;
  wire _abc_42016_n1476;
  wire _abc_42016_n1477;
  wire _abc_42016_n1478;
  wire _abc_42016_n1479;
  wire _abc_42016_n1480;
  wire _abc_42016_n1481;
  wire _abc_42016_n1482;
  wire _abc_42016_n1483;
  wire _abc_42016_n1484;
  wire _abc_42016_n1485;
  wire _abc_42016_n1486;
  wire _abc_42016_n1487;
  wire _abc_42016_n1488;
  wire _abc_42016_n1489;
  wire _abc_42016_n1490;
  wire _abc_42016_n1491;
  wire _abc_42016_n1492;
  wire _abc_42016_n1493;
  wire _abc_42016_n1494;
  wire _abc_42016_n1495;
  wire _abc_42016_n1496_1;
  wire _abc_42016_n1497;
  wire _abc_42016_n1498;
  wire _abc_42016_n1500;
  wire _abc_42016_n1501;
  wire _abc_42016_n1502;
  wire _abc_42016_n1503;
  wire _abc_42016_n1504;
  wire _abc_42016_n1505;
  wire _abc_42016_n1506;
  wire _abc_42016_n1507;
  wire _abc_42016_n1508;
  wire _abc_42016_n1509;
  wire _abc_42016_n1510;
  wire _abc_42016_n1511;
  wire _abc_42016_n1512;
  wire _abc_42016_n1513;
  wire _abc_42016_n1514;
  wire _abc_42016_n1515;
  wire _abc_42016_n1516;
  wire _abc_42016_n1517;
  wire _abc_42016_n1518;
  wire _abc_42016_n1519;
  wire _abc_42016_n1520;
  wire _abc_42016_n1521;
  wire _abc_42016_n1522_1;
  wire _abc_42016_n1523;
  wire _abc_42016_n1524;
  wire _abc_42016_n1526;
  wire _abc_42016_n1527;
  wire _abc_42016_n1528;
  wire _abc_42016_n1529;
  wire _abc_42016_n1530;
  wire _abc_42016_n1531;
  wire _abc_42016_n1532;
  wire _abc_42016_n1533;
  wire _abc_42016_n1534;
  wire _abc_42016_n1535;
  wire _abc_42016_n1536;
  wire _abc_42016_n1537;
  wire _abc_42016_n1538;
  wire _abc_42016_n1539;
  wire _abc_42016_n1540;
  wire _abc_42016_n1541;
  wire _abc_42016_n1542;
  wire _abc_42016_n1543;
  wire _abc_42016_n1544;
  wire _abc_42016_n1545;
  wire _abc_42016_n1546;
  wire _abc_42016_n1547;
  wire _abc_42016_n1548;
  wire _abc_42016_n1549;
  wire _abc_42016_n1550;
  wire _abc_42016_n1551;
  wire _abc_42016_n1553;
  wire _abc_42016_n1554;
  wire _abc_42016_n1555;
  wire _abc_42016_n1556;
  wire _abc_42016_n1557;
  wire _abc_42016_n1558;
  wire _abc_42016_n1559;
  wire _abc_42016_n1560;
  wire _abc_42016_n1561;
  wire _abc_42016_n1562;
  wire _abc_42016_n1563;
  wire _abc_42016_n1564;
  wire _abc_42016_n1565;
  wire _abc_42016_n1566;
  wire _abc_42016_n1567;
  wire _abc_42016_n1568;
  wire _abc_42016_n1569;
  wire _abc_42016_n1570;
  wire _abc_42016_n1571;
  wire _abc_42016_n1572;
  wire _abc_42016_n1573;
  wire _abc_42016_n1574;
  wire _abc_42016_n1575;
  wire _abc_42016_n1576;
  wire _abc_42016_n1577;
  wire _abc_42016_n1578_1;
  wire _abc_42016_n1579;
  wire _abc_42016_n1580;
  wire _abc_42016_n1581;
  wire _abc_42016_n1583;
  wire _abc_42016_n1584_1;
  wire _abc_42016_n1585;
  wire _abc_42016_n1586_1;
  wire _abc_42016_n1587;
  wire _abc_42016_n1588_1;
  wire _abc_42016_n1589;
  wire _abc_42016_n1590_1;
  wire _abc_42016_n1591;
  wire _abc_42016_n1592_1;
  wire _abc_42016_n1593;
  wire _abc_42016_n1594_1;
  wire _abc_42016_n1595;
  wire _abc_42016_n1596_1;
  wire _abc_42016_n1597;
  wire _abc_42016_n1598;
  wire _abc_42016_n1599_1;
  wire _abc_42016_n1600_1;
  wire _abc_42016_n1601_1;
  wire _abc_42016_n1603_1;
  wire _abc_42016_n1604_1;
  wire _abc_42016_n1605_1;
  wire _abc_42016_n1606_1;
  wire _abc_42016_n1607_1;
  wire _abc_42016_n1609;
  wire _abc_42016_n1611;
  wire _abc_42016_n1613;
  wire _abc_42016_n1615;
  wire _abc_42016_n1617;
  wire _abc_42016_n1619;
  wire _abc_42016_n1621;
  wire _abc_42016_n1623;
  wire _abc_42016_n1624;
  wire _abc_42016_n1625;
  wire _abc_42016_n1626;
  wire _abc_42016_n1627;
  wire _abc_42016_n1628;
  wire _abc_42016_n1629_1;
  wire _abc_42016_n1630_1;
  wire _abc_42016_n1631;
  wire _abc_42016_n1632;
  wire _abc_42016_n1633;
  wire _abc_42016_n1634;
  wire _abc_42016_n1635;
  wire _abc_42016_n1636;
  wire _abc_42016_n1637;
  wire _abc_42016_n1638_1;
  wire _abc_42016_n1639_1;
  wire _abc_42016_n1640;
  wire _abc_42016_n1641;
  wire _abc_42016_n1642;
  wire _abc_42016_n1643;
  wire _abc_42016_n1645;
  wire _abc_42016_n1646;
  wire _abc_42016_n1647_1;
  wire _abc_42016_n1648;
  wire _abc_42016_n1649_1;
  wire _abc_42016_n1650;
  wire _abc_42016_n1651;
  wire _abc_42016_n1652_1;
  wire _abc_42016_n1653;
  wire _abc_42016_n1654;
  wire _abc_42016_n1655;
  wire _abc_42016_n1656;
  wire _abc_42016_n1657;
  wire _abc_42016_n1658_1;
  wire _abc_42016_n1659;
  wire _abc_42016_n1660;
  wire _abc_42016_n1661;
  wire _abc_42016_n1663;
  wire _abc_42016_n1664_1;
  wire _abc_42016_n1665;
  wire _abc_42016_n1666;
  wire _abc_42016_n1667;
  wire _abc_42016_n1668;
  wire _abc_42016_n1669;
  wire _abc_42016_n1670;
  wire _abc_42016_n1671;
  wire _abc_42016_n1672;
  wire _abc_42016_n1673_1;
  wire _abc_42016_n1674_1;
  wire _abc_42016_n1675;
  wire _abc_42016_n1676;
  wire _abc_42016_n1677;
  wire _abc_42016_n1678;
  wire _abc_42016_n1679;
  wire _abc_42016_n1680;
  wire _abc_42016_n1681_1;
  wire _abc_42016_n1682_1;
  wire _abc_42016_n1683;
  wire _abc_42016_n1684;
  wire _abc_42016_n1686;
  wire _abc_42016_n1687;
  wire _abc_42016_n1688;
  wire _abc_42016_n1689_1;
  wire _abc_42016_n1690_1;
  wire _abc_42016_n1691;
  wire _abc_42016_n1692;
  wire _abc_42016_n1693;
  wire _abc_42016_n1694;
  wire _abc_42016_n1695;
  wire _abc_42016_n1696;
  wire _abc_42016_n1697_1;
  wire _abc_42016_n1698_1;
  wire _abc_42016_n1699;
  wire _abc_42016_n1700;
  wire _abc_42016_n1701;
  wire _abc_42016_n1702;
  wire _abc_42016_n1703;
  wire _abc_42016_n1704;
  wire _abc_42016_n1706_1;
  wire _abc_42016_n1707;
  wire _abc_42016_n1708;
  wire _abc_42016_n1709;
  wire _abc_42016_n1710;
  wire _abc_42016_n1711;
  wire _abc_42016_n1712;
  wire _abc_42016_n1713_1;
  wire _abc_42016_n1714_1;
  wire _abc_42016_n1715;
  wire _abc_42016_n1716;
  wire _abc_42016_n1717;
  wire _abc_42016_n1718;
  wire _abc_42016_n1719;
  wire _abc_42016_n1720;
  wire _abc_42016_n1721_1;
  wire _abc_42016_n1722_1;
  wire _abc_42016_n1723;
  wire _abc_42016_n1724;
  wire _abc_42016_n1725;
  wire _abc_42016_n1727;
  wire _abc_42016_n1728;
  wire _abc_42016_n1729_1;
  wire _abc_42016_n1730;
  wire _abc_42016_n1731;
  wire _abc_42016_n1732_1;
  wire _abc_42016_n1733;
  wire _abc_42016_n1734;
  wire _abc_42016_n1735;
  wire _abc_42016_n1736;
  wire _abc_42016_n1737;
  wire _abc_42016_n1738;
  wire _abc_42016_n1739;
  wire _abc_42016_n1740;
  wire _abc_42016_n1741;
  wire _abc_42016_n1742;
  wire _abc_42016_n1743;
  wire _abc_42016_n1744;
  wire _abc_42016_n1745;
  wire _abc_42016_n1746;
  wire _abc_42016_n1747;
  wire _abc_42016_n1749_1;
  wire _abc_42016_n1750_1;
  wire _abc_42016_n1751;
  wire _abc_42016_n1752;
  wire _abc_42016_n1753;
  wire _abc_42016_n1754;
  wire _abc_42016_n1755;
  wire _abc_42016_n1756;
  wire _abc_42016_n1758;
  wire _abc_42016_n1759;
  wire _abc_42016_n1760;
  wire _abc_42016_n1761;
  wire _abc_42016_n1762;
  wire _abc_42016_n1763;
  wire _abc_42016_n1764;
  wire _abc_42016_n1765;
  wire _abc_42016_n1767_1;
  wire _abc_42016_n1768;
  wire _abc_42016_n1769;
  wire _abc_42016_n1771;
  wire _abc_42016_n1772;
  wire _abc_42016_n1774;
  wire _abc_42016_n1775;
  wire _abc_42016_n1777;
  wire _abc_42016_n1778;
  wire _abc_42016_n1780;
  wire _abc_42016_n1781;
  wire _abc_42016_n1783_1;
  wire _abc_42016_n1784_1;
  wire _abc_42016_n1785;
  wire _abc_42016_n1787;
  wire _abc_42016_n1788;
  wire _abc_42016_n1789;
  wire _abc_42016_n1790;
  wire _abc_42016_n1791;
  wire _abc_42016_n1792;
  wire _abc_42016_n1793;
  wire _abc_42016_n1794;
  wire _abc_42016_n1795;
  wire _abc_42016_n1796;
  wire _abc_42016_n1797;
  wire _abc_42016_n1798;
  wire _abc_42016_n1800;
  wire _abc_42016_n1801_1;
  wire _abc_42016_n1802_1;
  wire _abc_42016_n1803;
  wire _abc_42016_n1804;
  wire _abc_42016_n1805;
  wire _abc_42016_n1806;
  wire _abc_42016_n1807;
  wire _abc_42016_n1808;
  wire _abc_42016_n1809;
  wire _abc_42016_n1810;
  wire _abc_42016_n1811;
  wire _abc_42016_n1813;
  wire _abc_42016_n1814;
  wire _abc_42016_n1815;
  wire _abc_42016_n1816;
  wire _abc_42016_n1818;
  wire _abc_42016_n1820_1;
  wire _abc_42016_n1822;
  wire _abc_42016_n1824;
  wire _abc_42016_n1826;
  wire _abc_42016_n1827;
  wire _abc_42016_n1829;
  wire _abc_42016_n1830;
  wire _abc_42016_n1832;
  wire _abc_42016_n1833;
  wire _abc_42016_n1835;
  wire _abc_42016_n1836;
  wire _abc_42016_n1837_1;
  wire _abc_42016_n1838_1;
  wire _abc_42016_n1839;
  wire _abc_42016_n1840;
  wire _abc_42016_n1841;
  wire _abc_42016_n1842;
  wire _abc_42016_n1843;
  wire _abc_42016_n1844;
  wire _abc_42016_n1846;
  wire _abc_42016_n1847;
  wire _abc_42016_n1848;
  wire _abc_42016_n1849;
  wire _abc_42016_n1850;
  wire _abc_42016_n1851;
  wire _abc_42016_n1852;
  wire _abc_42016_n1853;
  wire _abc_42016_n1854;
  wire _abc_42016_n1856_1;
  wire _abc_42016_n1857;
  wire _abc_42016_n1858;
  wire _abc_42016_n1860;
  wire _abc_42016_n1861;
  wire _abc_42016_n1863;
  wire _abc_42016_n1864;
  wire _abc_42016_n1865;
  wire _abc_42016_n1866;
  wire _abc_42016_n1867;
  wire _abc_42016_n1868;
  wire _abc_42016_n1869;
  wire _abc_42016_n1870;
  wire _abc_42016_n1871;
  wire _abc_42016_n1872;
  wire _abc_42016_n1873_1;
  wire _abc_42016_n1874_1;
  wire _abc_42016_n1875_1;
  wire _abc_42016_n1876;
  wire _abc_42016_n1878;
  wire _abc_42016_n1879_1;
  wire _abc_42016_n1880;
  wire _abc_42016_n1881;
  wire _abc_42016_n1882;
  wire _abc_42016_n1883;
  wire _abc_42016_n1885;
  wire _abc_42016_n1886_1;
  wire _abc_42016_n1888_1;
  wire _abc_42016_n1889;
  wire _abc_42016_n1891;
  wire _abc_42016_n1892;
  wire _abc_42016_n1894_1;
  wire _abc_42016_n1895;
  wire _abc_42016_n1897;
  wire _abc_42016_n1898;
  wire _abc_42016_n1900;
  wire _abc_42016_n1901_1;
  wire _abc_42016_n1903_1;
  wire _abc_42016_n1904;
  wire _abc_42016_n1905_1;
  wire _abc_42016_n1906;
  wire _abc_42016_n1907;
  wire _abc_42016_n1908;
  wire _abc_42016_n1909_1;
  wire _abc_42016_n1910;
  wire _abc_42016_n1911;
  wire _abc_42016_n1912;
  wire _abc_42016_n1913;
  wire _abc_42016_n1914;
  wire _abc_42016_n1915;
  wire _abc_42016_n1916;
  wire _abc_42016_n1917;
  wire _abc_42016_n1918;
  wire _abc_42016_n1919;
  wire _abc_42016_n1920;
  wire _abc_42016_n1921;
  wire _abc_42016_n1922_1;
  wire _abc_42016_n1923;
  wire _abc_42016_n1924;
  wire _abc_42016_n1925;
  wire _abc_42016_n1926_1;
  wire _abc_42016_n1927;
  wire _abc_42016_n1928;
  wire _abc_42016_n1929;
  wire _abc_42016_n1930;
  wire _abc_42016_n1931;
  wire _abc_42016_n1933;
  wire _abc_42016_n1934;
  wire _abc_42016_n1935;
  wire _abc_42016_n1936;
  wire _abc_42016_n1937;
  wire _abc_42016_n1938;
  wire _abc_42016_n1939;
  wire _abc_42016_n1940;
  wire _abc_42016_n1941;
  wire _abc_42016_n1942;
  wire _abc_42016_n1943;
  wire _abc_42016_n1944;
  wire _abc_42016_n1945;
  wire _abc_42016_n1946;
  wire _abc_42016_n1948;
  wire _abc_42016_n1949;
  wire _abc_42016_n1950_1;
  wire _abc_42016_n1951;
  wire _abc_42016_n1952_1;
  wire _abc_42016_n1953;
  wire _abc_42016_n1954;
  wire _abc_42016_n1955_1;
  wire _abc_42016_n1956;
  wire _abc_42016_n1957_1;
  wire _abc_42016_n1958;
  wire _abc_42016_n1959;
  wire _abc_42016_n1961_1;
  wire _abc_42016_n1962;
  wire _abc_42016_n1963_1;
  wire _abc_42016_n1964;
  wire _abc_42016_n1965;
  wire _abc_42016_n1966_1;
  wire _abc_42016_n1967;
  wire _abc_42016_n1968_1;
  wire _abc_42016_n1969;
  wire _abc_42016_n1970;
  wire _abc_42016_n1971;
  wire _abc_42016_n1972;
  wire _abc_42016_n1974;
  wire _abc_42016_n1975;
  wire _abc_42016_n1976;
  wire _abc_42016_n1977;
  wire _abc_42016_n1978;
  wire _abc_42016_n1979;
  wire _abc_42016_n1980;
  wire _abc_42016_n1981;
  wire _abc_42016_n1982;
  wire _abc_42016_n1983;
  wire _abc_42016_n1984;
  wire _abc_42016_n1985;
  wire _abc_42016_n1987;
  wire _abc_42016_n1988;
  wire _abc_42016_n1989;
  wire _abc_42016_n1990;
  wire _abc_42016_n1991;
  wire _abc_42016_n1992;
  wire _abc_42016_n1993;
  wire _abc_42016_n1994;
  wire _abc_42016_n1995;
  wire _abc_42016_n1996;
  wire _abc_42016_n1997;
  wire _abc_42016_n1998;
  wire _abc_42016_n2000;
  wire _abc_42016_n2001;
  wire _abc_42016_n2002;
  wire _abc_42016_n2003;
  wire _abc_42016_n2004;
  wire _abc_42016_n2005;
  wire _abc_42016_n2006;
  wire _abc_42016_n2007;
  wire _abc_42016_n2008;
  wire _abc_42016_n2009;
  wire _abc_42016_n2011;
  wire _abc_42016_n2012;
  wire _abc_42016_n2013;
  wire _abc_42016_n2014;
  wire _abc_42016_n2015;
  wire _abc_42016_n2016;
  wire _abc_42016_n2017;
  wire _abc_42016_n2018;
  wire _abc_42016_n2019;
  wire _abc_42016_n2020;
  wire _abc_42016_n2021;
  wire _abc_42016_n2022;
  wire _abc_42016_n2024;
  wire _abc_42016_n2025;
  wire _abc_42016_n2026;
  wire _abc_42016_n2027;
  wire _abc_42016_n2029;
  wire _abc_42016_n2030;
  wire _abc_42016_n2031;
  wire _abc_42016_n2032;
  wire _abc_42016_n2033;
  wire _abc_42016_n2034;
  wire _abc_42016_n2035;
  wire _abc_42016_n2036;
  wire _abc_42016_n2037;
  wire _abc_42016_n2038;
  wire _abc_42016_n2039;
  wire _abc_42016_n2040;
  wire _abc_42016_n2041;
  wire _abc_42016_n2042;
  wire _abc_42016_n2043;
  wire _abc_42016_n2044;
  wire _abc_42016_n2045;
  wire _abc_42016_n2046;
  wire _abc_42016_n2047;
  wire _abc_42016_n2048;
  wire _abc_42016_n2050;
  wire _abc_42016_n2051;
  wire _abc_42016_n2052;
  wire _abc_42016_n2053;
  wire _abc_42016_n2054;
  wire _abc_42016_n2056;
  wire _abc_42016_n2057;
  wire _abc_42016_n2058;
  wire _abc_42016_n2059;
  wire _abc_42016_n2060;
  wire _abc_42016_n2061;
  wire _abc_42016_n2062;
  wire _abc_42016_n2064;
  wire _abc_42016_n2065;
  wire _abc_42016_n2066;
  wire _abc_42016_n2067;
  wire _abc_42016_n2068;
  wire _abc_42016_n2069;
  wire _abc_42016_n2070;
  wire _abc_42016_n2071;
  wire _abc_42016_n2072;
  wire _abc_42016_n2073;
  wire _abc_42016_n2074;
  wire _abc_42016_n2075;
  wire _abc_42016_n2076;
  wire _abc_42016_n2078;
  wire _abc_42016_n2079;
  wire _abc_42016_n2080;
  wire _abc_42016_n2081;
  wire _abc_42016_n2082;
  wire _abc_42016_n2083;
  wire _abc_42016_n2084;
  wire _abc_42016_n2085;
  wire _abc_42016_n2086;
  wire _abc_42016_n2087;
  wire _abc_42016_n2088;
  wire _abc_42016_n2089;
  wire _abc_42016_n2090;
  wire _abc_42016_n2091;
  wire _abc_42016_n2092;
  wire _abc_42016_n2093;
  wire _abc_42016_n2094;
  wire _abc_42016_n2095;
  wire _abc_42016_n2096;
  wire _abc_42016_n2097;
  wire _abc_42016_n2098;
  wire _abc_42016_n2099;
  wire _abc_42016_n2100;
  wire _abc_42016_n2101;
  wire _abc_42016_n2102_1;
  wire _abc_42016_n2103;
  wire _abc_42016_n2104;
  wire _abc_42016_n2105;
  wire _abc_42016_n2106;
  wire _abc_42016_n2107;
  wire _abc_42016_n2108;
  wire _abc_42016_n2109_1;
  wire _abc_42016_n2110_1;
  wire _abc_42016_n2111;
  wire _abc_42016_n2112;
  wire _abc_42016_n2113;
  wire _abc_42016_n2114;
  wire _abc_42016_n2115_1;
  wire _abc_42016_n2116_1;
  wire _abc_42016_n2117;
  wire _abc_42016_n2118;
  wire _abc_42016_n2119_1;
  wire _abc_42016_n2120_1;
  wire _abc_42016_n2121;
  wire _abc_42016_n2122;
  wire _abc_42016_n2123_1;
  wire _abc_42016_n2124_1;
  wire _abc_42016_n2125;
  wire _abc_42016_n2126;
  wire _abc_42016_n2127_1;
  wire _abc_42016_n2128_1;
  wire _abc_42016_n2129;
  wire _abc_42016_n2130;
  wire _abc_42016_n2131_1;
  wire _abc_42016_n2132_1;
  wire _abc_42016_n2133;
  wire _abc_42016_n2134;
  wire _abc_42016_n2135_1;
  wire _abc_42016_n2136_1;
  wire _abc_42016_n2137;
  wire _abc_42016_n2138;
  wire _abc_42016_n2139_1;
  wire _abc_42016_n2140_1;
  wire _abc_42016_n2141;
  wire _abc_42016_n2142;
  wire _abc_42016_n2143_1;
  wire _abc_42016_n2144_1;
  wire _abc_42016_n2145;
  wire _abc_42016_n2146;
  wire _abc_42016_n2147;
  wire _abc_42016_n2148;
  wire _abc_42016_n2149;
  wire _abc_42016_n2150;
  wire _abc_42016_n2151_1;
  wire _abc_42016_n2152;
  wire _abc_42016_n2153;
  wire _abc_42016_n2154;
  wire _abc_42016_n2155;
  wire _abc_42016_n2156;
  wire _abc_42016_n2157;
  wire _abc_42016_n2158;
  wire _abc_42016_n2159;
  wire _abc_42016_n2160;
  wire _abc_42016_n2161;
  wire _abc_42016_n2162;
  wire _abc_42016_n2163;
  wire _abc_42016_n2164;
  wire _abc_42016_n2165;
  wire _abc_42016_n2166;
  wire _abc_42016_n2167;
  wire _abc_42016_n2168;
  wire _abc_42016_n2169;
  wire _abc_42016_n2170;
  wire _abc_42016_n2171;
  wire _abc_42016_n2172_1;
  wire _abc_42016_n2173;
  wire _abc_42016_n2174;
  wire _abc_42016_n2175;
  wire _abc_42016_n2176;
  wire _abc_42016_n2177;
  wire _abc_42016_n2178;
  wire _abc_42016_n2179;
  wire _abc_42016_n2180;
  wire _abc_42016_n2181;
  wire _abc_42016_n2182;
  wire _abc_42016_n2183;
  wire _abc_42016_n2184;
  wire _abc_42016_n2185;
  wire _abc_42016_n2186;
  wire _abc_42016_n2187;
  wire _abc_42016_n2188;
  wire _abc_42016_n2189;
  wire _abc_42016_n2190;
  wire _abc_42016_n2191;
  wire _abc_42016_n2192;
  wire _abc_42016_n2193;
  wire _abc_42016_n2194;
  wire _abc_42016_n2195;
  wire _abc_42016_n2196;
  wire _abc_42016_n2197;
  wire _abc_42016_n2198;
  wire _abc_42016_n2199;
  wire _abc_42016_n2200;
  wire _abc_42016_n2201;
  wire _abc_42016_n2202;
  wire _abc_42016_n2203;
  wire _abc_42016_n2204;
  wire _abc_42016_n2205;
  wire _abc_42016_n2206;
  wire _abc_42016_n2207;
  wire _abc_42016_n2208;
  wire _abc_42016_n2209;
  wire _abc_42016_n2210;
  wire _abc_42016_n2211;
  wire _abc_42016_n2212;
  wire _abc_42016_n2213;
  wire _abc_42016_n2214;
  wire _abc_42016_n2215;
  wire _abc_42016_n2216;
  wire _abc_42016_n2217;
  wire _abc_42016_n2218;
  wire _abc_42016_n2219;
  wire _abc_42016_n2220;
  wire _abc_42016_n2221;
  wire _abc_42016_n2222;
  wire _abc_42016_n2223;
  wire _abc_42016_n2225;
  wire _abc_42016_n2226;
  wire _abc_42016_n2227;
  wire _abc_42016_n2228;
  wire _abc_42016_n2229;
  wire _abc_42016_n2230;
  wire _abc_42016_n2231;
  wire _abc_42016_n2232;
  wire _abc_42016_n2234;
  wire _abc_42016_n2235;
  wire _abc_42016_n2237;
  wire _abc_42016_n2238;
  wire _abc_42016_n2240;
  wire _abc_42016_n2241;
  wire _abc_42016_n2243;
  wire _abc_42016_n2244;
  wire _abc_42016_n2246;
  wire _abc_42016_n2248;
  wire _abc_42016_n2250;
  wire _abc_42016_n2251;
  wire _abc_42016_n2253;
  wire _abc_42016_n2254;
  wire _abc_42016_n2255;
  wire _abc_42016_n2256;
  wire _abc_42016_n2257;
  wire _abc_42016_n2259;
  wire _abc_42016_n2260;
  wire _abc_42016_n2261;
  wire _abc_42016_n2262;
  wire _abc_42016_n2263;
  wire _abc_42016_n2264;
  wire _abc_42016_n2265;
  wire _abc_42016_n2266;
  wire _abc_42016_n2267;
  wire _abc_42016_n2268;
  wire _abc_42016_n2269;
  wire _abc_42016_n2270_1;
  wire _abc_42016_n2271_1;
  wire _abc_42016_n2272;
  wire _abc_42016_n2273;
  wire _abc_42016_n2274;
  wire _abc_42016_n2275;
  wire _abc_42016_n2276;
  wire _abc_42016_n2277;
  wire _abc_42016_n2278;
  wire _abc_42016_n2279;
  wire _abc_42016_n2280;
  wire _abc_42016_n2281;
  wire _abc_42016_n2282;
  wire _abc_42016_n2283;
  wire _abc_42016_n2284;
  wire _abc_42016_n2285;
  wire _abc_42016_n2286;
  wire _abc_42016_n2287;
  wire _abc_42016_n2288;
  wire _abc_42016_n2289;
  wire _abc_42016_n2290;
  wire _abc_42016_n2291;
  wire _abc_42016_n2292;
  wire _abc_42016_n2293;
  wire _abc_42016_n2294;
  wire _abc_42016_n2295;
  wire _abc_42016_n2296_1;
  wire _abc_42016_n2297_1;
  wire _abc_42016_n2298;
  wire _abc_42016_n2299;
  wire _abc_42016_n2300;
  wire _abc_42016_n2301;
  wire _abc_42016_n2302;
  wire _abc_42016_n2303;
  wire _abc_42016_n2304;
  wire _abc_42016_n2305;
  wire _abc_42016_n2306;
  wire _abc_42016_n2307;
  wire _abc_42016_n2308;
  wire _abc_42016_n2309;
  wire _abc_42016_n2310;
  wire _abc_42016_n2311;
  wire _abc_42016_n2312;
  wire _abc_42016_n2313;
  wire _abc_42016_n2314;
  wire _abc_42016_n2315;
  wire _abc_42016_n2316;
  wire _abc_42016_n2317;
  wire _abc_42016_n2318;
  wire _abc_42016_n2319;
  wire _abc_42016_n2320;
  wire _abc_42016_n2321;
  wire _abc_42016_n2322;
  wire _abc_42016_n2323_1;
  wire _abc_42016_n2324_1;
  wire _abc_42016_n2325;
  wire _abc_42016_n2326;
  wire _abc_42016_n2327;
  wire _abc_42016_n2328;
  wire _abc_42016_n2329;
  wire _abc_42016_n2330;
  wire _abc_42016_n2331;
  wire _abc_42016_n2332;
  wire _abc_42016_n2333;
  wire _abc_42016_n2334;
  wire _abc_42016_n2335;
  wire _abc_42016_n2336;
  wire _abc_42016_n2337;
  wire _abc_42016_n2338;
  wire _abc_42016_n2339;
  wire _abc_42016_n2340;
  wire _abc_42016_n2341;
  wire _abc_42016_n2342;
  wire _abc_42016_n2344;
  wire _abc_42016_n2345;
  wire _abc_42016_n2346;
  wire _abc_42016_n2347_1;
  wire _abc_42016_n2348_1;
  wire _abc_42016_n2349;
  wire _abc_42016_n2350;
  wire _abc_42016_n2351;
  wire _abc_42016_n2352;
  wire _abc_42016_n2353;
  wire _abc_42016_n2354;
  wire _abc_42016_n2355;
  wire _abc_42016_n2356;
  wire _abc_42016_n2357;
  wire _abc_42016_n2358;
  wire _abc_42016_n2359;
  wire _abc_42016_n2360;
  wire _abc_42016_n2361;
  wire _abc_42016_n2362;
  wire _abc_42016_n2363;
  wire _abc_42016_n2364;
  wire _abc_42016_n2365;
  wire _abc_42016_n2366;
  wire _abc_42016_n2367;
  wire _abc_42016_n2369;
  wire _abc_42016_n2370;
  wire _abc_42016_n2371;
  wire _abc_42016_n2372_1;
  wire _abc_42016_n2373_1;
  wire _abc_42016_n2374;
  wire _abc_42016_n2375;
  wire _abc_42016_n2376;
  wire _abc_42016_n2377;
  wire _abc_42016_n2378;
  wire _abc_42016_n2379;
  wire _abc_42016_n2380;
  wire _abc_42016_n2381;
  wire _abc_42016_n2382;
  wire _abc_42016_n2383;
  wire _abc_42016_n2384;
  wire _abc_42016_n2385;
  wire _abc_42016_n2386;
  wire _abc_42016_n2387;
  wire _abc_42016_n2388;
  wire _abc_42016_n2389;
  wire _abc_42016_n2390;
  wire _abc_42016_n2391;
  wire _abc_42016_n2392;
  wire _abc_42016_n2394_1;
  wire _abc_42016_n2395;
  wire _abc_42016_n2396;
  wire _abc_42016_n2397;
  wire _abc_42016_n2398_1;
  wire _abc_42016_n2399;
  wire _abc_42016_n2400;
  wire _abc_42016_n2401;
  wire _abc_42016_n2402_1;
  wire _abc_42016_n2403;
  wire _abc_42016_n2404;
  wire _abc_42016_n2405_1;
  wire _abc_42016_n2406;
  wire _abc_42016_n2407;
  wire _abc_42016_n2408_1;
  wire _abc_42016_n2409;
  wire _abc_42016_n2410;
  wire _abc_42016_n2411_1;
  wire _abc_42016_n2412;
  wire _abc_42016_n2413;
  wire _abc_42016_n2414_1;
  wire _abc_42016_n2415;
  wire _abc_42016_n2417_1;
  wire _abc_42016_n2418;
  wire _abc_42016_n2419;
  wire _abc_42016_n2420_1;
  wire _abc_42016_n2421;
  wire _abc_42016_n2422;
  wire _abc_42016_n2423_1;
  wire _abc_42016_n2424;
  wire _abc_42016_n2425;
  wire _abc_42016_n2426_1;
  wire _abc_42016_n2427;
  wire _abc_42016_n2428;
  wire _abc_42016_n2429_1;
  wire _abc_42016_n2430;
  wire _abc_42016_n2431;
  wire _abc_42016_n2432_1;
  wire _abc_42016_n2433;
  wire _abc_42016_n2434;
  wire _abc_42016_n2435_1;
  wire _abc_42016_n2436;
  wire _abc_42016_n2437;
  wire _abc_42016_n2438_1;
  wire _abc_42016_n2439;
  wire _abc_42016_n2440;
  wire _abc_42016_n2441_1;
  wire _abc_42016_n2442;
  wire _abc_42016_n2443;
  wire _abc_42016_n2444_1;
  wire _abc_42016_n2446;
  wire _abc_42016_n2447_1;
  wire _abc_42016_n2448;
  wire _abc_42016_n2449;
  wire _abc_42016_n2450_1;
  wire _abc_42016_n2451;
  wire _abc_42016_n2452;
  wire _abc_42016_n2453;
  wire _abc_42016_n2454;
  wire _abc_42016_n2455_1;
  wire _abc_42016_n2457;
  wire _abc_42016_n2458;
  wire _abc_42016_n2460;
  wire _abc_42016_n2462;
  wire _abc_42016_n2463;
  wire _abc_42016_n2465;
  wire _abc_42016_n2467;
  wire _abc_42016_n2469;
  wire _abc_42016_n2471;
  wire _abc_42016_n2472;
  wire _abc_42016_n2474;
  wire _abc_42016_n2476;
  wire _abc_42016_n2478;
  wire _abc_42016_n2479;
  wire _abc_42016_n2481;
  wire _abc_42016_n2483;
  wire _abc_42016_n2485;
  wire _abc_42016_n2487_1;
  wire _abc_42016_n2489;
  wire _abc_42016_n2492;
  wire _abc_42016_n2494;
  wire _abc_42016_n2496;
  wire _abc_42016_n2497;
  wire _abc_42016_n2498;
  wire _abc_42016_n2499;
  wire _abc_42016_n2500;
  wire _abc_42016_n2501;
  wire _abc_42016_n2502;
  wire _abc_42016_n2503;
  wire _abc_42016_n2504;
  wire _abc_42016_n2505;
  wire _abc_42016_n2506;
  wire _abc_42016_n2507;
  wire _abc_42016_n2508;
  wire _abc_42016_n2509;
  wire _abc_42016_n2510;
  wire _abc_42016_n2511;
  wire _abc_42016_n2512;
  wire _abc_42016_n2513;
  wire _abc_42016_n2514;
  wire _abc_42016_n2515;
  wire _abc_42016_n2516;
  wire _abc_42016_n2517_1;
  wire _abc_42016_n2518_1;
  wire _abc_42016_n2519;
  wire _abc_42016_n2520;
  wire _abc_42016_n2521;
  wire _abc_42016_n2522;
  wire _abc_42016_n2524;
  wire _abc_42016_n2525;
  wire _abc_42016_n2526;
  wire _abc_42016_n2527;
  wire _abc_42016_n2528;
  wire _abc_42016_n2529;
  wire _abc_42016_n2530;
  wire _abc_42016_n2531;
  wire _abc_42016_n2532;
  wire _abc_42016_n2533;
  wire _abc_42016_n2534;
  wire _abc_42016_n2535;
  wire _abc_42016_n2536;
  wire _abc_42016_n2537;
  wire _abc_42016_n2538;
  wire _abc_42016_n2539;
  wire _abc_42016_n2540;
  wire _abc_42016_n2541;
  wire _abc_42016_n2542;
  wire _abc_42016_n2543;
  wire _abc_42016_n2544;
  wire _abc_42016_n2545;
  wire _abc_42016_n2546;
  wire _abc_42016_n2547_1;
  wire _abc_42016_n2548_1;
  wire _abc_42016_n2549;
  wire _abc_42016_n2550;
  wire _abc_42016_n2551;
  wire _abc_42016_n2552;
  wire _abc_42016_n2553;
  wire _abc_42016_n2555;
  wire _abc_42016_n2556;
  wire _abc_42016_n2557;
  wire _abc_42016_n2558;
  wire _abc_42016_n2559;
  wire _abc_42016_n2560;
  wire _abc_42016_n2561;
  wire _abc_42016_n2562;
  wire _abc_42016_n2563;
  wire _abc_42016_n2564;
  wire _abc_42016_n2565;
  wire _abc_42016_n2566;
  wire _abc_42016_n2567;
  wire _abc_42016_n2568;
  wire _abc_42016_n2569;
  wire _abc_42016_n2570;
  wire _abc_42016_n2571;
  wire _abc_42016_n2572;
  wire _abc_42016_n2573;
  wire _abc_42016_n2574;
  wire _abc_42016_n2575;
  wire _abc_42016_n2576;
  wire _abc_42016_n2577;
  wire _abc_42016_n2578_1;
  wire _abc_42016_n2579_1;
  wire _abc_42016_n2580;
  wire _abc_42016_n2581;
  wire _abc_42016_n2582;
  wire _abc_42016_n2583;
  wire _abc_42016_n2584;
  wire _abc_42016_n2585;
  wire _abc_42016_n2587;
  wire _abc_42016_n2588;
  wire _abc_42016_n2589;
  wire _abc_42016_n2590;
  wire _abc_42016_n2591;
  wire _abc_42016_n2592;
  wire _abc_42016_n2593;
  wire _abc_42016_n2594;
  wire _abc_42016_n2595;
  wire _abc_42016_n2596;
  wire _abc_42016_n2597;
  wire _abc_42016_n2598;
  wire _abc_42016_n2599;
  wire _abc_42016_n2600;
  wire _abc_42016_n2601;
  wire _abc_42016_n2602;
  wire _abc_42016_n2603;
  wire _abc_42016_n2604;
  wire _abc_42016_n2605;
  wire _abc_42016_n2606;
  wire _abc_42016_n2607;
  wire _abc_42016_n2608_1;
  wire _abc_42016_n2609_1;
  wire _abc_42016_n2610;
  wire _abc_42016_n2611;
  wire _abc_42016_n2612;
  wire _abc_42016_n2613;
  wire _abc_42016_n2614;
  wire _abc_42016_n2615;
  wire _abc_42016_n2616;
  wire _abc_42016_n2617;
  wire _abc_42016_n2619;
  wire _abc_42016_n2620;
  wire _abc_42016_n2621;
  wire _abc_42016_n2622;
  wire _abc_42016_n2623;
  wire _abc_42016_n2624;
  wire _abc_42016_n2625;
  wire _abc_42016_n2626;
  wire _abc_42016_n2627;
  wire _abc_42016_n2628;
  wire _abc_42016_n2629;
  wire _abc_42016_n2630;
  wire _abc_42016_n2631;
  wire _abc_42016_n2632;
  wire _abc_42016_n2633;
  wire _abc_42016_n2634;
  wire _abc_42016_n2635;
  wire _abc_42016_n2636;
  wire _abc_42016_n2637;
  wire _abc_42016_n2638;
  wire _abc_42016_n2639_1;
  wire _abc_42016_n2640_1;
  wire _abc_42016_n2641;
  wire _abc_42016_n2642;
  wire _abc_42016_n2643;
  wire _abc_42016_n2644;
  wire _abc_42016_n2645;
  wire _abc_42016_n2646;
  wire _abc_42016_n2648;
  wire _abc_42016_n2649;
  wire _abc_42016_n2650;
  wire _abc_42016_n2651;
  wire _abc_42016_n2652;
  wire _abc_42016_n2653;
  wire _abc_42016_n2654;
  wire _abc_42016_n2655;
  wire _abc_42016_n2656;
  wire _abc_42016_n2657;
  wire _abc_42016_n2658;
  wire _abc_42016_n2659;
  wire _abc_42016_n2660;
  wire _abc_42016_n2661;
  wire _abc_42016_n2662;
  wire _abc_42016_n2663;
  wire _abc_42016_n2664;
  wire _abc_42016_n2665;
  wire _abc_42016_n2666;
  wire _abc_42016_n2667;
  wire _abc_42016_n2668;
  wire _abc_42016_n2669;
  wire _abc_42016_n2670;
  wire _abc_42016_n2671;
  wire _abc_42016_n2672_1;
  wire _abc_42016_n2674;
  wire _abc_42016_n2675;
  wire _abc_42016_n2676;
  wire _abc_42016_n2677;
  wire _abc_42016_n2678;
  wire _abc_42016_n2679;
  wire _abc_42016_n2680;
  wire _abc_42016_n2681;
  wire _abc_42016_n2682;
  wire _abc_42016_n2683;
  wire _abc_42016_n2684;
  wire _abc_42016_n2685;
  wire _abc_42016_n2686;
  wire _abc_42016_n2687;
  wire _abc_42016_n2688;
  wire _abc_42016_n2689;
  wire _abc_42016_n2690;
  wire _abc_42016_n2691;
  wire _abc_42016_n2692;
  wire _abc_42016_n2693;
  wire _abc_42016_n2694;
  wire _abc_42016_n2695;
  wire _abc_42016_n2696;
  wire _abc_42016_n2697;
  wire _abc_42016_n2698;
  wire _abc_42016_n2700;
  wire _abc_42016_n2701;
  wire _abc_42016_n2702;
  wire _abc_42016_n2703;
  wire _abc_42016_n2704;
  wire _abc_42016_n2705;
  wire _abc_42016_n2706_1;
  wire _abc_42016_n2707;
  wire _abc_42016_n2708;
  wire _abc_42016_n2709;
  wire _abc_42016_n2710;
  wire _abc_42016_n2711_1;
  wire _abc_42016_n2712;
  wire _abc_42016_n2713;
  wire _abc_42016_n2714;
  wire _abc_42016_n2715;
  wire _abc_42016_n2716;
  wire _abc_42016_n2717;
  wire _abc_42016_n2718;
  wire _abc_42016_n2719;
  wire _abc_42016_n2720;
  wire _abc_42016_n2721;
  wire _abc_42016_n2722;
  wire _abc_42016_n2723;
  wire _abc_42016_n2724;
  wire _abc_42016_n2725;
  wire _abc_42016_n2726;
  wire _abc_42016_n2727;
  wire _abc_42016_n2728;
  wire _abc_42016_n2729;
  wire _abc_42016_n2731;
  wire _abc_42016_n2732;
  wire _abc_42016_n2733;
  wire _abc_42016_n2734;
  wire _abc_42016_n2735;
  wire _abc_42016_n2736;
  wire _abc_42016_n2737;
  wire _abc_42016_n2738;
  wire _abc_42016_n2739;
  wire _abc_42016_n2740;
  wire _abc_42016_n2741;
  wire _abc_42016_n2742;
  wire _abc_42016_n2743;
  wire _abc_42016_n2744;
  wire _abc_42016_n2745;
  wire _abc_42016_n2746;
  wire _abc_42016_n2747_1;
  wire _abc_42016_n2748_1;
  wire _abc_42016_n2749;
  wire _abc_42016_n2750;
  wire _abc_42016_n2751;
  wire _abc_42016_n2752;
  wire _abc_42016_n2753;
  wire _abc_42016_n2754;
  wire _abc_42016_n2755;
  wire _abc_42016_n2756;
  wire _abc_42016_n2757;
  wire _abc_42016_n2758;
  wire _abc_42016_n2759;
  wire _abc_42016_n2760;
  wire _abc_42016_n2761;
  wire _abc_42016_n2762;
  wire _abc_42016_n2763;
  wire _abc_42016_n2765;
  wire _abc_42016_n2766;
  wire _abc_42016_n2767_1;
  wire _abc_42016_n2768_1;
  wire _abc_42016_n2769;
  wire _abc_42016_n2770;
  wire _abc_42016_n2771;
  wire _abc_42016_n2772;
  wire _abc_42016_n2773;
  wire _abc_42016_n2774;
  wire _abc_42016_n2775;
  wire _abc_42016_n2776;
  wire _abc_42016_n2777;
  wire _abc_42016_n2778;
  wire _abc_42016_n2779;
  wire _abc_42016_n2780;
  wire _abc_42016_n2781;
  wire _abc_42016_n2782;
  wire _abc_42016_n2783;
  wire _abc_42016_n2784;
  wire _abc_42016_n2786;
  wire _abc_42016_n2787;
  wire _abc_42016_n2788_1;
  wire _abc_42016_n2789_1;
  wire _abc_42016_n2790;
  wire _abc_42016_n2791;
  wire _abc_42016_n2792;
  wire _abc_42016_n2793;
  wire _abc_42016_n2794;
  wire _abc_42016_n2795;
  wire _abc_42016_n2796;
  wire _abc_42016_n2797;
  wire _abc_42016_n2798;
  wire _abc_42016_n2799;
  wire _abc_42016_n2800;
  wire _abc_42016_n2801;
  wire _abc_42016_n2803;
  wire _abc_42016_n2804;
  wire _abc_42016_n2805;
  wire _abc_42016_n2806;
  wire _abc_42016_n2807;
  wire _abc_42016_n2808;
  wire _abc_42016_n2809;
  wire _abc_42016_n2810_1;
  wire _abc_42016_n2811_1;
  wire _abc_42016_n2812;
  wire _abc_42016_n2813;
  wire _abc_42016_n2814;
  wire _abc_42016_n2815;
  wire _abc_42016_n2816;
  wire _abc_42016_n2817;
  wire _abc_42016_n2818;
  wire _abc_42016_n2820;
  wire _abc_42016_n2821;
  wire _abc_42016_n2822;
  wire _abc_42016_n2823;
  wire _abc_42016_n2824;
  wire _abc_42016_n2825;
  wire _abc_42016_n2826;
  wire _abc_42016_n2827;
  wire _abc_42016_n2828;
  wire _abc_42016_n2829;
  wire _abc_42016_n2830;
  wire _abc_42016_n2831;
  wire _abc_42016_n2832;
  wire _abc_42016_n2833_1;
  wire _abc_42016_n2834_1;
  wire _abc_42016_n2836;
  wire _abc_42016_n2837;
  wire _abc_42016_n2838;
  wire _abc_42016_n2839;
  wire _abc_42016_n2840;
  wire _abc_42016_n2841;
  wire _abc_42016_n2842;
  wire _abc_42016_n2843;
  wire _abc_42016_n2844;
  wire _abc_42016_n2845;
  wire _abc_42016_n2846;
  wire _abc_42016_n2847;
  wire _abc_42016_n2848;
  wire _abc_42016_n2849;
  wire _abc_42016_n2850;
  wire _abc_42016_n2852;
  wire _abc_42016_n2853;
  wire _abc_42016_n2854;
  wire _abc_42016_n2855_1;
  wire _abc_42016_n2856_1;
  wire _abc_42016_n2857;
  wire _abc_42016_n2858;
  wire _abc_42016_n2859;
  wire _abc_42016_n2860;
  wire _abc_42016_n2861;
  wire _abc_42016_n2862;
  wire _abc_42016_n2863;
  wire _abc_42016_n2864;
  wire _abc_42016_n2865;
  wire _abc_42016_n2866;
  wire _abc_42016_n2867;
  wire _abc_42016_n2869;
  wire _abc_42016_n2870;
  wire _abc_42016_n2871;
  wire _abc_42016_n2872;
  wire _abc_42016_n2873;
  wire _abc_42016_n2874;
  wire _abc_42016_n2875;
  wire _abc_42016_n2876;
  wire _abc_42016_n2877;
  wire _abc_42016_n2878_1;
  wire _abc_42016_n2879_1;
  wire _abc_42016_n2880;
  wire _abc_42016_n2881;
  wire _abc_42016_n2882;
  wire _abc_42016_n2883;
  wire _abc_42016_n2884;
  wire _abc_42016_n2885;
  wire _abc_42016_n2887;
  wire _abc_42016_n2888;
  wire _abc_42016_n2889;
  wire _abc_42016_n2890;
  wire _abc_42016_n2891;
  wire _abc_42016_n2892;
  wire _abc_42016_n2893;
  wire _abc_42016_n2894;
  wire _abc_42016_n2895;
  wire _abc_42016_n2896;
  wire _abc_42016_n2897;
  wire _abc_42016_n2898;
  wire _abc_42016_n2899;
  wire _abc_42016_n2900_1;
  wire _abc_42016_n2902;
  wire _abc_42016_n2903;
  wire _abc_42016_n2904;
  wire _abc_42016_n2905;
  wire _abc_42016_n2906;
  wire _abc_42016_n2907;
  wire _abc_42016_n2908;
  wire _abc_42016_n2909;
  wire _abc_42016_n2910;
  wire _abc_42016_n2911;
  wire _abc_42016_n2912;
  wire _abc_42016_n2913;
  wire _abc_42016_n2914;
  wire _abc_42016_n2915;
  wire _abc_42016_n2916;
  wire _abc_42016_n2917;
  wire _abc_42016_n2918;
  wire _abc_42016_n2920;
  wire _abc_42016_n2921;
  wire _abc_42016_n2922;
  wire _abc_42016_n2923;
  wire _abc_42016_n2924_1;
  wire _abc_42016_n2925_1;
  wire _abc_42016_n2926;
  wire _abc_42016_n2927;
  wire _abc_42016_n2928;
  wire _abc_42016_n2929;
  wire _abc_42016_n2930;
  wire _abc_42016_n2931;
  wire _abc_42016_n2932;
  wire _abc_42016_n2933;
  wire _abc_42016_n2934;
  wire _abc_42016_n2935;
  wire _abc_42016_n2936;
  wire _abc_42016_n2937;
  wire _abc_42016_n2938;
  wire _abc_42016_n2940;
  wire _abc_42016_n2941;
  wire _abc_42016_n2942;
  wire _abc_42016_n2943;
  wire _abc_42016_n2944;
  wire _abc_42016_n2945;
  wire _abc_42016_n2946_1;
  wire _abc_42016_n2947_1;
  wire _abc_42016_n2948;
  wire _abc_42016_n2949;
  wire _abc_42016_n2950;
  wire _abc_42016_n2951;
  wire _abc_42016_n2952;
  wire _abc_42016_n2953;
  wire _abc_42016_n2954;
  wire _abc_42016_n2956;
  wire _abc_42016_n2957;
  wire _abc_42016_n2958;
  wire _abc_42016_n2959;
  wire _abc_42016_n2960;
  wire _abc_42016_n2961;
  wire _abc_42016_n2962;
  wire _abc_42016_n2963;
  wire _abc_42016_n2964;
  wire _abc_42016_n2965;
  wire _abc_42016_n2966;
  wire _abc_42016_n2967;
  wire _abc_42016_n2968;
  wire _abc_42016_n2969_1;
  wire _abc_42016_n2970_1;
  wire _abc_42016_n2972;
  wire _abc_42016_n2973;
  wire _abc_42016_n2974;
  wire _abc_42016_n2975;
  wire _abc_42016_n2976;
  wire _abc_42016_n2977;
  wire _abc_42016_n2978;
  wire _abc_42016_n2979;
  wire _abc_42016_n2980;
  wire _abc_42016_n2981;
  wire _abc_42016_n2982;
  wire _abc_42016_n2983;
  wire _abc_42016_n2984;
  wire _abc_42016_n2985;
  wire _abc_42016_n2986;
  wire _abc_42016_n2987;
  wire _abc_42016_n2988;
  wire _abc_42016_n2990_1;
  wire _abc_42016_n2991_1;
  wire _abc_42016_n2992;
  wire _abc_42016_n2993;
  wire _abc_42016_n2994;
  wire _abc_42016_n2995;
  wire _abc_42016_n2996;
  wire _abc_42016_n2997;
  wire _abc_42016_n2998;
  wire _abc_42016_n2999;
  wire _abc_42016_n3000;
  wire _abc_42016_n3001;
  wire _abc_42016_n3002;
  wire _abc_42016_n3003;
  wire _abc_42016_n3004;
  wire _abc_42016_n3005;
  wire _abc_42016_n3006;
  wire _abc_42016_n3007;
  wire _abc_42016_n3009;
  wire _abc_42016_n3010;
  wire _abc_42016_n3011;
  wire _abc_42016_n3012;
  wire _abc_42016_n3013;
  wire _abc_42016_n3014_1;
  wire _abc_42016_n3015_1;
  wire _abc_42016_n3016;
  wire _abc_42016_n3017;
  wire _abc_42016_n3018;
  wire _abc_42016_n3019;
  wire _abc_42016_n3020;
  wire _abc_42016_n3021;
  wire _abc_42016_n3022;
  wire _abc_42016_n3023;
  wire _abc_42016_n3024;
  wire _abc_42016_n3025;
  wire _abc_42016_n3026;
  wire _abc_42016_n3028;
  wire _abc_42016_n3029;
  wire _abc_42016_n3030;
  wire _abc_42016_n3031;
  wire _abc_42016_n3032;
  wire _abc_42016_n3033;
  wire _abc_42016_n3034;
  wire _abc_42016_n3035_1;
  wire _abc_42016_n3036_1;
  wire _abc_42016_n3037;
  wire _abc_42016_n3038;
  wire _abc_42016_n3039;
  wire _abc_42016_n3040;
  wire _abc_42016_n3041;
  wire _abc_42016_n3042;
  wire _abc_42016_n3043;
  wire _abc_42016_n3044;
  wire _abc_42016_n3045;
  wire _abc_42016_n3046;
  wire _abc_42016_n3047;
  wire _abc_42016_n3048;
  wire _abc_42016_n3050;
  wire _abc_42016_n3051;
  wire _abc_42016_n3052;
  wire _abc_42016_n3053;
  wire _abc_42016_n3054;
  wire _abc_42016_n3055;
  wire _abc_42016_n3056;
  wire _abc_42016_n3057_1;
  wire _abc_42016_n3058_1;
  wire _abc_42016_n3059;
  wire _abc_42016_n3060;
  wire _abc_42016_n3061;
  wire _abc_42016_n3062;
  wire _abc_42016_n3063;
  wire _abc_42016_n3064;
  wire _abc_42016_n3065;
  wire _abc_42016_n3066;
  wire _abc_42016_n3067;
  wire _abc_42016_n3068;
  wire _abc_42016_n3069;
  wire _abc_42016_n3070;
  wire _abc_42016_n3071;
  wire _abc_42016_n3072;
  wire _abc_42016_n3073;
  wire _abc_42016_n3074;
  wire _abc_42016_n3075;
  wire _abc_42016_n3076;
  wire _abc_42016_n3078_1;
  wire _abc_42016_n3079;
  wire _abc_42016_n3080_1;
  wire _abc_42016_n3081;
  wire _abc_42016_n3082;
  wire _abc_42016_n3083;
  wire _abc_42016_n3084;
  wire _abc_42016_n3085;
  wire _abc_42016_n3086;
  wire _abc_42016_n3087;
  wire _abc_42016_n3088;
  wire _abc_42016_n3089;
  wire _abc_42016_n3090;
  wire _abc_42016_n3091;
  wire _abc_42016_n3092;
  wire _abc_42016_n3093;
  wire _abc_42016_n3094;
  wire _abc_42016_n3095;
  wire _abc_42016_n3096;
  wire _abc_42016_n3097;
  wire _abc_42016_n3098;
  wire _abc_42016_n3099;
  wire _abc_42016_n3100;
  wire _abc_42016_n3101;
  wire _abc_42016_n3102;
  wire _abc_42016_n3103;
  wire _abc_42016_n3105_1;
  wire _abc_42016_n3106_1;
  wire _abc_42016_n3107;
  wire _abc_42016_n3108;
  wire _abc_42016_n3109;
  wire _abc_42016_n3110;
  wire _abc_42016_n3111;
  wire _abc_42016_n3112;
  wire _abc_42016_n3113;
  wire _abc_42016_n3114;
  wire _abc_42016_n3115;
  wire _abc_42016_n3116;
  wire _abc_42016_n3117;
  wire _abc_42016_n3118;
  wire _abc_42016_n3119;
  wire _abc_42016_n3120;
  wire _abc_42016_n3121;
  wire _abc_42016_n3122;
  wire _abc_42016_n3123;
  wire _abc_42016_n3124;
  wire _abc_42016_n3125_1;
  wire _abc_42016_n3126_1;
  wire _abc_42016_n3128;
  wire _abc_42016_n3129;
  wire _abc_42016_n3130;
  wire _abc_42016_n3131;
  wire _abc_42016_n3132;
  wire _abc_42016_n3133;
  wire _abc_42016_n3134;
  wire _abc_42016_n3135;
  wire _abc_42016_n3136;
  wire _abc_42016_n3137;
  wire _abc_42016_n3138;
  wire _abc_42016_n3139;
  wire _abc_42016_n3140;
  wire _abc_42016_n3141;
  wire _abc_42016_n3142;
  wire _abc_42016_n3143;
  wire _abc_42016_n3144;
  wire _abc_42016_n3145;
  wire _abc_42016_n3146;
  wire _abc_42016_n3147_1;
  wire _abc_42016_n3148_1;
  wire _abc_42016_n3149;
  wire _abc_42016_n3150;
  wire _abc_42016_n3151;
  wire _abc_42016_n3153;
  wire _abc_42016_n3154;
  wire _abc_42016_n3155;
  wire _abc_42016_n3156;
  wire _abc_42016_n3157;
  wire _abc_42016_n3158;
  wire _abc_42016_n3159;
  wire _abc_42016_n3160;
  wire _abc_42016_n3161;
  wire _abc_42016_n3162;
  wire _abc_42016_n3163;
  wire _abc_42016_n3164;
  wire _abc_42016_n3165;
  wire _abc_42016_n3166;
  wire _abc_42016_n3167;
  wire _abc_42016_n3168;
  wire _abc_42016_n3169_1;
  wire _abc_42016_n3170_1;
  wire _abc_42016_n3171;
  wire _abc_42016_n3172;
  wire _abc_42016_n3173;
  wire _abc_42016_n3175;
  wire _abc_42016_n3176;
  wire _abc_42016_n3177;
  wire _abc_42016_n3178;
  wire _abc_42016_n3179;
  wire _abc_42016_n3180;
  wire _abc_42016_n3181;
  wire _abc_42016_n3182;
  wire _abc_42016_n3183;
  wire _abc_42016_n3184;
  wire _abc_42016_n3185;
  wire _abc_42016_n3186;
  wire _abc_42016_n3187;
  wire _abc_42016_n3188;
  wire _abc_42016_n3189;
  wire _abc_42016_n3190;
  wire _abc_42016_n3191;
  wire _abc_42016_n3192;
  wire _abc_42016_n3193;
  wire _abc_42016_n3194;
  wire _abc_42016_n3195_1;
  wire _abc_42016_n3196_1;
  wire _abc_42016_n3197;
  wire _abc_42016_n3198;
  wire _abc_42016_n3199;
  wire _abc_42016_n3201;
  wire _abc_42016_n3202;
  wire _abc_42016_n3203;
  wire _abc_42016_n3204;
  wire _abc_42016_n3205;
  wire _abc_42016_n3206;
  wire _abc_42016_n3207;
  wire _abc_42016_n3208;
  wire _abc_42016_n3209;
  wire _abc_42016_n3210;
  wire _abc_42016_n3211;
  wire _abc_42016_n3212;
  wire _abc_42016_n3213;
  wire _abc_42016_n3214;
  wire _abc_42016_n3215;
  wire _abc_42016_n3216;
  wire _abc_42016_n3217_1;
  wire _abc_42016_n3218_1;
  wire _abc_42016_n3219;
  wire _abc_42016_n3220;
  wire _abc_42016_n3221;
  wire _abc_42016_n3223;
  wire _abc_42016_n3224;
  wire _abc_42016_n3225;
  wire _abc_42016_n3226;
  wire _abc_42016_n3227;
  wire _abc_42016_n3228;
  wire _abc_42016_n3229;
  wire _abc_42016_n3230;
  wire _abc_42016_n3231;
  wire _abc_42016_n3232;
  wire _abc_42016_n3233;
  wire _abc_42016_n3234;
  wire _abc_42016_n3235;
  wire _abc_42016_n3236;
  wire _abc_42016_n3237;
  wire _abc_42016_n3238;
  wire _abc_42016_n3239;
  wire _abc_42016_n3240;
  wire _abc_42016_n3241;
  wire _abc_42016_n3242;
  wire _abc_42016_n3243;
  wire _abc_42016_n3245_1;
  wire _abc_42016_n3246;
  wire _abc_42016_n3247;
  wire _abc_42016_n3248;
  wire _abc_42016_n3249;
  wire _abc_42016_n3250;
  wire _abc_42016_n3251;
  wire _abc_42016_n3252;
  wire _abc_42016_n3253;
  wire _abc_42016_n3254;
  wire _abc_42016_n3255;
  wire _abc_42016_n3256;
  wire _abc_42016_n3257;
  wire _abc_42016_n3258;
  wire _abc_42016_n3259;
  wire _abc_42016_n3260;
  wire _abc_42016_n3261;
  wire _abc_42016_n3262;
  wire _abc_42016_n3263;
  wire _abc_42016_n3264;
  wire _abc_42016_n3265;
  wire _abc_42016_n3266_1;
  wire _abc_42016_n3268;
  wire _abc_42016_n3269;
  wire _abc_42016_n3270;
  wire _abc_42016_n3271;
  wire _abc_42016_n3272;
  wire _abc_42016_n3273;
  wire _abc_42016_n3274;
  wire _abc_42016_n3275;
  wire _abc_42016_n3276;
  wire _abc_42016_n3277;
  wire _abc_42016_n3278;
  wire _abc_42016_n3279;
  wire _abc_42016_n3280;
  wire _abc_42016_n3281;
  wire _abc_42016_n3282;
  wire _abc_42016_n3283;
  wire _abc_42016_n3284;
  wire _abc_42016_n3285;
  wire _abc_42016_n3286;
  wire _abc_42016_n3287;
  wire _abc_42016_n3288;
  wire _abc_42016_n3289;
  wire _abc_42016_n3291;
  wire _abc_42016_n3292;
  wire _abc_42016_n3293;
  wire _abc_42016_n3294;
  wire _abc_42016_n3295_1;
  wire _abc_42016_n3296_1;
  wire _abc_42016_n3297;
  wire _abc_42016_n3298;
  wire _abc_42016_n3299;
  wire _abc_42016_n3300;
  wire _abc_42016_n3301;
  wire _abc_42016_n3302;
  wire _abc_42016_n3303;
  wire _abc_42016_n3304;
  wire _abc_42016_n3305;
  wire _abc_42016_n3306;
  wire _abc_42016_n3307;
  wire _abc_42016_n3308;
  wire _abc_42016_n3309;
  wire _abc_42016_n3310;
  wire _abc_42016_n3311;
  wire _abc_42016_n3312;
  wire _abc_42016_n3313;
  wire _abc_42016_n3314;
  wire _abc_42016_n3316;
  wire _abc_42016_n3317;
  wire _abc_42016_n3318_1;
  wire _abc_42016_n3319_1;
  wire _abc_42016_n3320;
  wire _abc_42016_n3321;
  wire _abc_42016_n3322;
  wire _abc_42016_n3323;
  wire _abc_42016_n3324;
  wire _abc_42016_n3325;
  wire _abc_42016_n3326;
  wire _abc_42016_n3327;
  wire _abc_42016_n3328;
  wire _abc_42016_n3329;
  wire _abc_42016_n3330;
  wire _abc_42016_n3331;
  wire _abc_42016_n3332;
  wire _abc_42016_n3333;
  wire _abc_42016_n3334;
  wire _abc_42016_n3335;
  wire _abc_42016_n3337;
  wire _abc_42016_n3338;
  wire _abc_42016_n3339;
  wire _abc_42016_n3340;
  wire _abc_42016_n3341;
  wire _abc_42016_n3342;
  wire _abc_42016_n3343;
  wire _abc_42016_n3344;
  wire _abc_42016_n3345_1;
  wire _abc_42016_n3346_1;
  wire _abc_42016_n3347;
  wire _abc_42016_n3348;
  wire _abc_42016_n3349;
  wire _abc_42016_n3350;
  wire _abc_42016_n3351;
  wire _abc_42016_n3352;
  wire _abc_42016_n3353;
  wire _abc_42016_n3354;
  wire _abc_42016_n3355;
  wire _abc_42016_n3356;
  wire _abc_42016_n3357;
  wire _abc_42016_n3358;
  wire _abc_42016_n3359;
  wire _abc_42016_n3361;
  wire _abc_42016_n3362;
  wire _abc_42016_n3363;
  wire _abc_42016_n3364;
  wire _abc_42016_n3365;
  wire _abc_42016_n3366;
  wire _abc_42016_n3367;
  wire _abc_42016_n3368_1;
  wire _abc_42016_n3369_1;
  wire _abc_42016_n3370;
  wire _abc_42016_n3371;
  wire _abc_42016_n3372;
  wire _abc_42016_n3373;
  wire _abc_42016_n3374;
  wire _abc_42016_n3375;
  wire _abc_42016_n3376;
  wire _abc_42016_n3377;
  wire _abc_42016_n3378;
  wire _abc_42016_n3379;
  wire _abc_42016_n3380;
  wire _abc_42016_n3381;
  wire _abc_42016_n3382;
  wire _abc_42016_n3383;
  wire _abc_42016_n3384;
  wire _abc_42016_n3385;
  wire _abc_42016_n3386;
  wire _abc_42016_n3388;
  wire _abc_42016_n3389;
  wire _abc_42016_n3390;
  wire _abc_42016_n3391;
  wire _abc_42016_n3392;
  wire _abc_42016_n3393;
  wire _abc_42016_n3394;
  wire _abc_42016_n3395;
  wire _abc_42016_n3396;
  wire _abc_42016_n3397_1;
  wire _abc_42016_n3398_1;
  wire _abc_42016_n3399;
  wire _abc_42016_n3400;
  wire _abc_42016_n3401;
  wire _abc_42016_n3402;
  wire _abc_42016_n3403;
  wire _abc_42016_n3404;
  wire _abc_42016_n3405;
  wire _abc_42016_n3407;
  wire _abc_42016_n3408;
  wire _abc_42016_n3409;
  wire _abc_42016_n3410;
  wire _abc_42016_n3411;
  wire _abc_42016_n3412;
  wire _abc_42016_n3414;
  wire _abc_42016_n3416;
  wire _abc_42016_n3418;
  wire _abc_42016_n3419;
  wire _abc_42016_n3421_1;
  wire _abc_42016_n3423;
  wire _abc_42016_n3425;
  wire _abc_42016_n3427;
  wire _abc_42016_n3429;
  wire _abc_42016_n3430;
  wire _abc_42016_n3431;
  wire _abc_42016_n3432;
  wire _abc_42016_n3433;
  wire _abc_42016_n3434;
  wire _abc_42016_n3435;
  wire _abc_42016_n3436;
  wire _abc_42016_n3437;
  wire _abc_42016_n3438;
  wire _abc_42016_n3440;
  wire _abc_42016_n3441;
  wire _abc_42016_n3442;
  wire _abc_42016_n3443;
  wire _abc_42016_n3444;
  wire _abc_42016_n3446;
  wire _abc_42016_n3447_1;
  wire _abc_42016_n3448_1;
  wire _abc_42016_n3449;
  wire _abc_42016_n3450;
  wire _abc_42016_n3452;
  wire _abc_42016_n3453;
  wire _abc_42016_n3454;
  wire _abc_42016_n3455;
  wire _abc_42016_n3456;
  wire _abc_42016_n3457;
  wire _abc_42016_n3458;
  wire _abc_42016_n3459;
  wire _abc_42016_n3460;
  wire _abc_42016_n3461;
  wire _abc_42016_n3462;
  wire _abc_42016_n3463;
  wire _abc_42016_n3464;
  wire _abc_42016_n3465;
  wire _abc_42016_n3466;
  wire _abc_42016_n3467;
  wire _abc_42016_n3469;
  wire _abc_42016_n3470_1;
  wire _abc_42016_n3471;
  wire _abc_42016_n3472;
  wire _abc_42016_n3473;
  wire _abc_42016_n3474;
  wire _abc_42016_n3475;
  wire _abc_42016_n3476_1;
  wire _abc_42016_n3477;
  wire _abc_42016_n3478;
  wire _abc_42016_n3479_1;
  wire _abc_42016_n3480;
  wire _abc_42016_n3481;
  wire _abc_42016_n3482_1;
  wire _abc_42016_n3483;
  wire _abc_42016_n3484;
  wire _abc_42016_n3486;
  wire _abc_42016_n3487;
  wire _abc_42016_n3488_1;
  wire _abc_42016_n3489;
  wire _abc_42016_n3490;
  wire _abc_42016_n3491_1;
  wire _abc_42016_n3492;
  wire _abc_42016_n3493;
  wire _abc_42016_n3494_1;
  wire _abc_42016_n3495;
  wire _abc_42016_n3496;
  wire _abc_42016_n3497_1;
  wire _abc_42016_n3498;
  wire _abc_42016_n3499;
  wire _abc_42016_n3500;
  wire _abc_42016_n3501;
  wire _abc_42016_n3502;
  wire _abc_42016_n3503;
  wire _abc_42016_n3504;
  wire _abc_42016_n3505;
  wire _abc_42016_n3506;
  wire _abc_42016_n3508;
  wire _abc_42016_n3509;
  wire _abc_42016_n3510_1;
  wire _abc_42016_n3511;
  wire _abc_42016_n3512;
  wire _abc_42016_n3513;
  wire _abc_42016_n3514;
  wire _abc_42016_n3515;
  wire _abc_42016_n3516;
  wire _abc_42016_n3517;
  wire _abc_42016_n3518_1;
  wire _abc_42016_n3519;
  wire _abc_42016_n3520;
  wire _abc_42016_n3521;
  wire _abc_42016_n3522;
  wire _abc_42016_n3523;
  wire _abc_42016_n3524;
  wire _abc_42016_n3525;
  wire _abc_42016_n3526_1;
  wire _abc_42016_n3527;
  wire _abc_42016_n3528;
  wire _abc_42016_n3529;
  wire _abc_42016_n3530;
  wire _abc_42016_n3532;
  wire _abc_42016_n3533;
  wire _abc_42016_n3534;
  wire _abc_42016_n3535;
  wire _abc_42016_n3536;
  wire _abc_42016_n3537;
  wire _abc_42016_n3538;
  wire _abc_42016_n3539;
  wire _abc_42016_n3540;
  wire _abc_42016_n3541;
  wire _abc_42016_n3542;
  wire _abc_42016_n3543;
  wire _abc_42016_n3544;
  wire _abc_42016_n3545;
  wire _abc_42016_n3546;
  wire _abc_42016_n3547;
  wire _abc_42016_n3548;
  wire _abc_42016_n3549;
  wire _abc_42016_n3550;
  wire _abc_42016_n3551;
  wire _abc_42016_n3552_1;
  wire _abc_42016_n3554;
  wire _abc_42016_n3555;
  wire _abc_42016_n3556;
  wire _abc_42016_n3557;
  wire _abc_42016_n3558;
  wire _abc_42016_n3559;
  wire _abc_42016_n3560;
  wire _abc_42016_n3561;
  wire _abc_42016_n3562;
  wire _abc_42016_n3563;
  wire _abc_42016_n3564;
  wire _abc_42016_n3565;
  wire _abc_42016_n3566;
  wire _abc_42016_n3567_1;
  wire _abc_42016_n3568;
  wire _abc_42016_n3569;
  wire _abc_42016_n3570;
  wire _abc_42016_n3571;
  wire _abc_42016_n3572;
  wire _abc_42016_n3573;
  wire _abc_42016_n3574;
  wire _abc_42016_n3575;
  wire _abc_42016_n3576;
  wire _abc_42016_n3577;
  wire _abc_42016_n3578;
  wire _abc_42016_n3579;
  wire _abc_42016_n3581;
  wire _abc_42016_n3582;
  wire _abc_42016_n3583;
  wire _abc_42016_n3584;
  wire _abc_42016_n3585;
  wire _abc_42016_n3586_1;
  wire _abc_42016_n3587;
  wire _abc_42016_n3588;
  wire _abc_42016_n3589;
  wire _abc_42016_n3590;
  wire _abc_42016_n3591;
  wire _abc_42016_n3592;
  wire _abc_42016_n3593;
  wire _abc_42016_n3594;
  wire _abc_42016_n3595;
  wire _abc_42016_n3596;
  wire _abc_42016_n3597;
  wire _abc_42016_n3598;
  wire _abc_42016_n3599;
  wire _abc_42016_n3600;
  wire _abc_42016_n3601;
  wire _abc_42016_n3602;
  wire _abc_42016_n3603;
  wire _abc_42016_n3605;
  wire _abc_42016_n3606_1;
  wire _abc_42016_n3607;
  wire _abc_42016_n3608;
  wire _abc_42016_n3609;
  wire _abc_42016_n3610;
  wire _abc_42016_n3611;
  wire _abc_42016_n3612;
  wire _abc_42016_n3613;
  wire _abc_42016_n3614;
  wire _abc_42016_n3615;
  wire _abc_42016_n3616;
  wire _abc_42016_n3617;
  wire _abc_42016_n3618;
  wire _abc_42016_n3619;
  wire _abc_42016_n3620;
  wire _abc_42016_n3621;
  wire _abc_42016_n3622;
  wire _abc_42016_n3623;
  wire _abc_42016_n3624;
  wire _abc_42016_n3626;
  wire _abc_42016_n3627;
  wire _abc_42016_n3628_1;
  wire _abc_42016_n3629;
  wire _abc_42016_n3630;
  wire _abc_42016_n3631;
  wire _abc_42016_n3632;
  wire _abc_42016_n3633;
  wire _abc_42016_n3634;
  wire _abc_42016_n3635;
  wire _abc_42016_n3636;
  wire _abc_42016_n3637;
  wire _abc_42016_n3638;
  wire _abc_42016_n3639;
  wire _abc_42016_n3640;
  wire _abc_42016_n3641;
  wire _abc_42016_n3642;
  wire _abc_42016_n3643;
  wire _abc_42016_n3644;
  wire _abc_42016_n3645;
  wire _abc_42016_n3646;
  wire _abc_42016_n3647;
  wire _abc_42016_n3649;
  wire _abc_42016_n3650;
  wire _abc_42016_n3651;
  wire _abc_42016_n3652;
  wire _abc_42016_n3653;
  wire _abc_42016_n3654;
  wire _abc_42016_n3655;
  wire _abc_42016_n3656;
  wire _abc_42016_n3657;
  wire _abc_42016_n3658;
  wire _abc_42016_n3659;
  wire _abc_42016_n3660;
  wire _abc_42016_n3661;
  wire _abc_42016_n3662;
  wire _abc_42016_n3663;
  wire _abc_42016_n3664;
  wire _abc_42016_n3665;
  wire _abc_42016_n3666;
  wire _abc_42016_n3667;
  wire _abc_42016_n3669;
  wire _abc_42016_n3670_1;
  wire _abc_42016_n3671;
  wire _abc_42016_n3672;
  wire _abc_42016_n3673;
  wire _abc_42016_n3674;
  wire _abc_42016_n3675;
  wire _abc_42016_n3676;
  wire _abc_42016_n3677;
  wire _abc_42016_n3678;
  wire _abc_42016_n3679;
  wire _abc_42016_n3680;
  wire _abc_42016_n3681;
  wire _abc_42016_n3682;
  wire _abc_42016_n3683;
  wire _abc_42016_n3684;
  wire _abc_42016_n3685;
  wire _abc_42016_n3686;
  wire _abc_42016_n3687;
  wire _abc_42016_n3688;
  wire _abc_42016_n3690_1;
  wire _abc_42016_n3691;
  wire _abc_42016_n3692;
  wire _abc_42016_n3693;
  wire _abc_42016_n3694;
  wire _abc_42016_n3695;
  wire _abc_42016_n3696;
  wire _abc_42016_n3697;
  wire _abc_42016_n3698;
  wire _abc_42016_n3699;
  wire _abc_42016_n3700;
  wire _abc_42016_n3701;
  wire _abc_42016_n3702;
  wire _abc_42016_n3703;
  wire _abc_42016_n3704;
  wire _abc_42016_n3705;
  wire _abc_42016_n3706;
  wire _abc_42016_n3707;
  wire _abc_42016_n3708;
  wire _abc_42016_n3709;
  wire _abc_42016_n3710;
  wire _abc_42016_n3711;
  wire _abc_42016_n3713_1;
  wire _abc_42016_n3714;
  wire _abc_42016_n3715;
  wire _abc_42016_n3716;
  wire _abc_42016_n3717;
  wire _abc_42016_n3718;
  wire _abc_42016_n3719;
  wire _abc_42016_n3720;
  wire _abc_42016_n3721;
  wire _abc_42016_n3722;
  wire _abc_42016_n3723;
  wire _abc_42016_n3724;
  wire _abc_42016_n3725;
  wire _abc_42016_n3726;
  wire _abc_42016_n3727;
  wire _abc_42016_n3728;
  wire _abc_42016_n3729;
  wire _abc_42016_n3730;
  wire _abc_42016_n3731;
  wire _abc_42016_n3732;
  wire _abc_42016_n3733_1;
  wire _abc_42016_n3734;
  wire _abc_42016_n3735;
  wire _abc_42016_n3737;
  wire _abc_42016_n3738;
  wire _abc_42016_n3739;
  wire _abc_42016_n3740;
  wire _abc_42016_n3741;
  wire _abc_42016_n3742;
  wire _abc_42016_n3743;
  wire _abc_42016_n3744;
  wire _abc_42016_n3745;
  wire _abc_42016_n3746;
  wire _abc_42016_n3747;
  wire _abc_42016_n3748;
  wire _abc_42016_n3749;
  wire _abc_42016_n3750;
  wire _abc_42016_n3751;
  wire _abc_42016_n3752;
  wire _abc_42016_n3753;
  wire _abc_42016_n3754;
  wire _abc_42016_n3755_1;
  wire _abc_42016_n3756;
  wire _abc_42016_n3758;
  wire _abc_42016_n3759;
  wire _abc_42016_n3760;
  wire _abc_42016_n3761;
  wire _abc_42016_n3762;
  wire _abc_42016_n3763;
  wire _abc_42016_n3764;
  wire _abc_42016_n3765;
  wire _abc_42016_n3766;
  wire _abc_42016_n3767;
  wire _abc_42016_n3768;
  wire _abc_42016_n3769;
  wire _abc_42016_n3770;
  wire _abc_42016_n3771;
  wire _abc_42016_n3772;
  wire _abc_42016_n3773;
  wire _abc_42016_n3774;
  wire _abc_42016_n3775_1;
  wire _abc_42016_n3776;
  wire _abc_42016_n3777;
  wire _abc_42016_n3779;
  wire _abc_42016_n3780;
  wire _abc_42016_n3781;
  wire _abc_42016_n3782;
  wire _abc_42016_n3783;
  wire _abc_42016_n3784;
  wire _abc_42016_n3785;
  wire _abc_42016_n3786;
  wire _abc_42016_n3787;
  wire _abc_42016_n3788;
  wire _abc_42016_n3789;
  wire _abc_42016_n3790;
  wire _abc_42016_n3791;
  wire _abc_42016_n3792;
  wire _abc_42016_n3793;
  wire _abc_42016_n3794;
  wire _abc_42016_n3795;
  wire _abc_42016_n3796;
  wire _abc_42016_n3797_1;
  wire _abc_42016_n3799;
  wire _abc_42016_n3800;
  wire _abc_42016_n3801;
  wire _abc_42016_n3802;
  wire _abc_42016_n3803;
  wire _abc_42016_n3804;
  wire _abc_42016_n3805;
  wire _abc_42016_n3806;
  wire _abc_42016_n3807;
  wire _abc_42016_n3808;
  wire _abc_42016_n3809;
  wire _abc_42016_n3810;
  wire _abc_42016_n3811;
  wire _abc_42016_n3812;
  wire _abc_42016_n3813;
  wire _abc_42016_n3814;
  wire _abc_42016_n3815;
  wire _abc_42016_n3816;
  wire _abc_42016_n3817_1;
  wire _abc_42016_n3818;
  wire _abc_42016_n3819;
  wire _abc_42016_n3820;
  wire _abc_42016_n3821;
  wire _abc_42016_n3822;
  wire _abc_42016_n3823;
  wire _abc_42016_n3824;
  wire _abc_42016_n3825;
  wire _abc_42016_n3826;
  wire _abc_42016_n3827;
  wire _abc_42016_n3828;
  wire _abc_42016_n3829;
  wire _abc_42016_n3830;
  wire _abc_42016_n3831;
  wire _abc_42016_n3833;
  wire _abc_42016_n3834;
  wire _abc_42016_n3835;
  wire _abc_42016_n3836;
  wire _abc_42016_n3837;
  wire _abc_42016_n3838;
  wire _abc_42016_n3839_1;
  wire _abc_42016_n3840;
  wire _abc_42016_n3841;
  wire _abc_42016_n3842;
  wire _abc_42016_n3843;
  wire _abc_42016_n3844;
  wire _abc_42016_n3845;
  wire _abc_42016_n3846;
  wire _abc_42016_n3847;
  wire _abc_42016_n3848;
  wire _abc_42016_n3849;
  wire _abc_42016_n3850;
  wire _abc_42016_n3851;
  wire _abc_42016_n3852;
  wire _abc_42016_n3853;
  wire _abc_42016_n3854;
  wire _abc_42016_n3855;
  wire _abc_42016_n3856;
  wire _abc_42016_n3857;
  wire _abc_42016_n3858;
  wire _abc_42016_n3859_1;
  wire _abc_42016_n3860;
  wire _abc_42016_n3861;
  wire _abc_42016_n3862;
  wire _abc_42016_n3864;
  wire _abc_42016_n3865;
  wire _abc_42016_n3866;
  wire _abc_42016_n3867;
  wire _abc_42016_n3868;
  wire _abc_42016_n3869;
  wire _abc_42016_n3870;
  wire _abc_42016_n3871;
  wire _abc_42016_n3872;
  wire _abc_42016_n3873;
  wire _abc_42016_n3874;
  wire _abc_42016_n3875;
  wire _abc_42016_n3876;
  wire _abc_42016_n3877;
  wire _abc_42016_n3878;
  wire _abc_42016_n3879;
  wire _abc_42016_n3880;
  wire _abc_42016_n3881;
  wire _abc_42016_n3882;
  wire _abc_42016_n3883;
  wire _abc_42016_n3884;
  wire _abc_42016_n3885;
  wire _abc_42016_n3886;
  wire _abc_42016_n3887;
  wire _abc_42016_n3888;
  wire _abc_42016_n3889;
  wire _abc_42016_n3890;
  wire _abc_42016_n3891;
  wire _abc_42016_n3892;
  wire _abc_42016_n3893;
  wire _abc_42016_n3894;
  wire _abc_42016_n3896;
  wire _abc_42016_n3897;
  wire _abc_42016_n3898;
  wire _abc_42016_n3899;
  wire _abc_42016_n3900;
  wire _abc_42016_n3901;
  wire _abc_42016_n3902;
  wire _abc_42016_n3903;
  wire _abc_42016_n3904;
  wire _abc_42016_n3905;
  wire _abc_42016_n3906;
  wire _abc_42016_n3907;
  wire _abc_42016_n3908;
  wire _abc_42016_n3909;
  wire _abc_42016_n3910;
  wire _abc_42016_n3911;
  wire _abc_42016_n3912;
  wire _abc_42016_n3913;
  wire _abc_42016_n3914;
  wire _abc_42016_n3915;
  wire _abc_42016_n3916;
  wire _abc_42016_n3917;
  wire _abc_42016_n3918;
  wire _abc_42016_n3919;
  wire _abc_42016_n3920;
  wire _abc_42016_n3921;
  wire _abc_42016_n3922;
  wire _abc_42016_n3923;
  wire _abc_42016_n3924;
  wire _abc_42016_n3926;
  wire _abc_42016_n3927;
  wire _abc_42016_n3928;
  wire _abc_42016_n3929;
  wire _abc_42016_n3930;
  wire _abc_42016_n3931;
  wire _abc_42016_n3932;
  wire _abc_42016_n3933;
  wire _abc_42016_n3934;
  wire _abc_42016_n3935_1;
  wire _abc_42016_n3936;
  wire _abc_42016_n3937;
  wire _abc_42016_n3938;
  wire _abc_42016_n3939;
  wire _abc_42016_n3940;
  wire _abc_42016_n3941;
  wire _abc_42016_n3942;
  wire _abc_42016_n3943;
  wire _abc_42016_n3944;
  wire _abc_42016_n3945;
  wire _abc_42016_n3946;
  wire _abc_42016_n3947;
  wire _abc_42016_n3948;
  wire _abc_42016_n3949;
  wire _abc_42016_n3950;
  wire _abc_42016_n3951;
  wire _abc_42016_n3952;
  wire _abc_42016_n3953;
  wire _abc_42016_n3955;
  wire _abc_42016_n3956;
  wire _abc_42016_n3957;
  wire _abc_42016_n3958;
  wire _abc_42016_n3959;
  wire _abc_42016_n3960;
  wire _abc_42016_n3961;
  wire _abc_42016_n3962;
  wire _abc_42016_n3963;
  wire _abc_42016_n3964;
  wire _abc_42016_n3965;
  wire _abc_42016_n3966;
  wire _abc_42016_n3967;
  wire _abc_42016_n3968;
  wire _abc_42016_n3969;
  wire _abc_42016_n3970;
  wire _abc_42016_n3971;
  wire _abc_42016_n3972;
  wire _abc_42016_n3973;
  wire _abc_42016_n3974;
  wire _abc_42016_n3975;
  wire _abc_42016_n3976;
  wire _abc_42016_n3977;
  wire _abc_42016_n3978;
  wire _abc_42016_n3979;
  wire _abc_42016_n3980;
  wire _abc_42016_n3981;
  wire _abc_42016_n3982;
  wire _abc_42016_n3983_1;
  wire _abc_42016_n3985;
  wire _abc_42016_n3986;
  wire _abc_42016_n3987;
  wire _abc_42016_n3988;
  wire _abc_42016_n3989;
  wire _abc_42016_n3990;
  wire _abc_42016_n3991;
  wire _abc_42016_n3992;
  wire _abc_42016_n3993;
  wire _abc_42016_n3994;
  wire _abc_42016_n3995;
  wire _abc_42016_n3996;
  wire _abc_42016_n3997;
  wire _abc_42016_n3998;
  wire _abc_42016_n3999;
  wire _abc_42016_n4000;
  wire _abc_42016_n4001;
  wire _abc_42016_n4002;
  wire _abc_42016_n4003;
  wire _abc_42016_n4004;
  wire _abc_42016_n4005;
  wire _abc_42016_n4006;
  wire _abc_42016_n4007;
  wire _abc_42016_n4008;
  wire _abc_42016_n4009;
  wire _abc_42016_n4011;
  wire _abc_42016_n4012;
  wire _abc_42016_n4013;
  wire _abc_42016_n4014;
  wire _abc_42016_n4015;
  wire _abc_42016_n4016;
  wire _abc_42016_n4017;
  wire _abc_42016_n4018;
  wire _abc_42016_n4019;
  wire _abc_42016_n4020;
  wire _abc_42016_n4021;
  wire _abc_42016_n4022;
  wire _abc_42016_n4023;
  wire _abc_42016_n4024;
  wire _abc_42016_n4025;
  wire _abc_42016_n4026;
  wire _abc_42016_n4027;
  wire _abc_42016_n4028;
  wire _abc_42016_n4029;
  wire _abc_42016_n4030;
  wire _abc_42016_n4031;
  wire _abc_42016_n4032;
  wire _abc_42016_n4033;
  wire _abc_42016_n4034;
  wire _abc_42016_n4035;
  wire _abc_42016_n4036;
  wire _abc_42016_n4037;
  wire _abc_42016_n4038;
  wire _abc_42016_n4039;
  wire _abc_42016_n4040;
  wire _abc_42016_n4041_1;
  wire _abc_42016_n4042;
  wire _abc_42016_n4043;
  wire _abc_42016_n4044;
  wire _abc_42016_n4045;
  wire _abc_42016_n4046;
  wire _abc_42016_n4047;
  wire _abc_42016_n4048;
  wire _abc_42016_n4049;
  wire _abc_42016_n4050;
  wire _abc_42016_n4051;
  wire _abc_42016_n4052;
  wire _abc_42016_n4053;
  wire _abc_42016_n4054;
  wire _abc_42016_n4055;
  wire _abc_42016_n4056;
  wire _abc_42016_n4057;
  wire _abc_42016_n4058;
  wire _abc_42016_n4059;
  wire _abc_42016_n4060;
  wire _abc_42016_n4061;
  wire _abc_42016_n4062;
  wire _abc_42016_n4063;
  wire _abc_42016_n4064;
  wire _abc_42016_n4065;
  wire _abc_42016_n4066;
  wire _abc_42016_n4067;
  wire _abc_42016_n4068;
  wire _abc_42016_n4069;
  wire _abc_42016_n4070;
  wire _abc_42016_n4071;
  wire _abc_42016_n4072;
  wire _abc_42016_n4073;
  wire _abc_42016_n4075;
  wire _abc_42016_n4076;
  wire _abc_42016_n4077;
  wire _abc_42016_n4078;
  wire _abc_42016_n4079;
  wire _abc_42016_n4080;
  wire _abc_42016_n4081;
  wire _abc_42016_n4082;
  wire _abc_42016_n4083;
  wire _abc_42016_n4084;
  wire _abc_42016_n4085;
  wire _abc_42016_n4086;
  wire _abc_42016_n4087;
  wire _abc_42016_n4088;
  wire _abc_42016_n4089;
  wire _abc_42016_n4090;
  wire _abc_42016_n4091;
  wire _abc_42016_n4092_1;
  wire _abc_42016_n4093;
  wire _abc_42016_n4094;
  wire _abc_42016_n4095;
  wire _abc_42016_n4096;
  wire _abc_42016_n4097;
  wire _abc_42016_n4098;
  wire _abc_42016_n4099;
  wire _abc_42016_n4100;
  wire _abc_42016_n4101;
  wire _abc_42016_n4102;
  wire _abc_42016_n4103;
  wire _abc_42016_n4104;
  wire _abc_42016_n4105;
  wire _abc_42016_n4106;
  wire _abc_42016_n4107;
  wire _abc_42016_n4108;
  wire _abc_42016_n4109;
  wire _abc_42016_n4110;
  wire _abc_42016_n4111;
  wire _abc_42016_n4112;
  wire _abc_42016_n4113;
  wire _abc_42016_n4114;
  wire _abc_42016_n4115;
  wire _abc_42016_n4116;
  wire _abc_42016_n4117;
  wire _abc_42016_n4118;
  wire _abc_42016_n4119;
  wire _abc_42016_n4120;
  wire _abc_42016_n4121;
  wire _abc_42016_n4122;
  wire _abc_42016_n4124;
  wire _abc_42016_n4125;
  wire _abc_42016_n4126;
  wire _abc_42016_n4127;
  wire _abc_42016_n4128;
  wire _abc_42016_n4129;
  wire _abc_42016_n4130;
  wire _abc_42016_n4131;
  wire _abc_42016_n4132;
  wire _abc_42016_n4133;
  wire _abc_42016_n4134;
  wire _abc_42016_n4135;
  wire _abc_42016_n4136;
  wire _abc_42016_n4137;
  wire _abc_42016_n4138;
  wire _abc_42016_n4139;
  wire _abc_42016_n4141;
  wire _abc_42016_n4142;
  wire _abc_42016_n4143;
  wire _abc_42016_n4144;
  wire _abc_42016_n4145;
  wire _abc_42016_n4146;
  wire _abc_42016_n4147;
  wire _abc_42016_n4148;
  wire _abc_42016_n4149;
  wire _abc_42016_n4150_1;
  wire _abc_42016_n4151;
  wire _abc_42016_n4152;
  wire _abc_42016_n4153;
  wire _abc_42016_n4154;
  wire _abc_42016_n4156;
  wire _abc_42016_n4157;
  wire _abc_42016_n4158;
  wire _abc_42016_n4159;
  wire _abc_42016_n4160;
  wire _abc_42016_n4161;
  wire _abc_42016_n4162;
  wire _abc_42016_n4163;
  wire _abc_42016_n4164;
  wire _abc_42016_n4165;
  wire _abc_42016_n4166;
  wire _abc_42016_n4167;
  wire _abc_42016_n4168;
  wire _abc_42016_n4169;
  wire _abc_42016_n4170;
  wire _abc_42016_n4172;
  wire _abc_42016_n4173;
  wire _abc_42016_n4174;
  wire _abc_42016_n4175;
  wire _abc_42016_n4176;
  wire _abc_42016_n4177;
  wire _abc_42016_n4178;
  wire _abc_42016_n4179;
  wire _abc_42016_n4180;
  wire _abc_42016_n4181;
  wire _abc_42016_n4182;
  wire _abc_42016_n4184;
  wire _abc_42016_n4185;
  wire _abc_42016_n4186;
  wire _abc_42016_n4187;
  wire _abc_42016_n4188;
  wire _abc_42016_n4189;
  wire _abc_42016_n4190;
  wire _abc_42016_n4191;
  wire _abc_42016_n4192;
  wire _abc_42016_n4193;
  wire _abc_42016_n4194;
  wire _abc_42016_n4195;
  wire _abc_42016_n4196;
  wire _abc_42016_n4198;
  wire _abc_42016_n4199;
  wire _abc_42016_n4200;
  wire _abc_42016_n4201;
  wire _abc_42016_n4202;
  wire _abc_42016_n4203;
  wire _abc_42016_n4204_1;
  wire _abc_42016_n4205;
  wire _abc_42016_n4206;
  wire _abc_42016_n4207;
  wire _abc_42016_n4208;
  wire _abc_42016_n4210;
  wire _abc_42016_n4211;
  wire _abc_42016_n4212;
  wire _abc_42016_n4213;
  wire _abc_42016_n4214;
  wire _abc_42016_n4215;
  wire _abc_42016_n4216;
  wire _abc_42016_n4217;
  wire _abc_42016_n4218;
  wire _abc_42016_n4219;
  wire _abc_42016_n4220;
  wire _abc_42016_n4221;
  wire _abc_42016_n4223;
  wire _abc_42016_n4224;
  wire _abc_42016_n4225;
  wire _abc_42016_n4226;
  wire _abc_42016_n4227;
  wire _abc_42016_n4228;
  wire _abc_42016_n4229;
  wire _abc_42016_n4230;
  wire _abc_42016_n4231;
  wire _abc_42016_n4232;
  wire _abc_42016_n4233;
  wire _abc_42016_n4234;
  wire _abc_42016_n4236;
  wire _abc_42016_n4237;
  wire _abc_42016_n4238;
  wire _abc_42016_n4239;
  wire _abc_42016_n4240;
  wire _abc_42016_n4241;
  wire _abc_42016_n4242;
  wire _abc_42016_n4243;
  wire _abc_42016_n4244;
  wire _abc_42016_n4245;
  wire _abc_42016_n4246;
  wire _abc_42016_n4247;
  wire _abc_42016_n4249;
  wire _abc_42016_n4250;
  wire _abc_42016_n4251;
  wire _abc_42016_n4252;
  wire _abc_42016_n4253;
  wire _abc_42016_n4254;
  wire _abc_42016_n4255;
  wire _abc_42016_n4256;
  wire _abc_42016_n4257;
  wire _abc_42016_n4258;
  wire _abc_42016_n4259;
  wire _abc_42016_n4261;
  wire _abc_42016_n4262;
  wire _abc_42016_n4263;
  wire _abc_42016_n4264;
  wire _abc_42016_n4265;
  wire _abc_42016_n4266_1;
  wire _abc_42016_n4267;
  wire _abc_42016_n4268;
  wire _abc_42016_n4269;
  wire _abc_42016_n4270;
  wire _abc_42016_n4271;
  wire _abc_42016_n4272;
  wire _abc_42016_n4273;
  wire _abc_42016_n4275;
  wire _abc_42016_n4276;
  wire _abc_42016_n4277;
  wire _abc_42016_n4278;
  wire _abc_42016_n4279;
  wire _abc_42016_n4280;
  wire _abc_42016_n4281;
  wire _abc_42016_n4282;
  wire _abc_42016_n4283;
  wire _abc_42016_n4284;
  wire _abc_42016_n4285;
  wire _abc_42016_n4287;
  wire _abc_42016_n4288;
  wire _abc_42016_n4289;
  wire _abc_42016_n4290;
  wire _abc_42016_n4291;
  wire _abc_42016_n4292;
  wire _abc_42016_n4293;
  wire _abc_42016_n4294;
  wire _abc_42016_n4295;
  wire _abc_42016_n4296;
  wire _abc_42016_n4297;
  wire _abc_42016_n4299;
  wire _abc_42016_n4300;
  wire _abc_42016_n4301;
  wire _abc_42016_n4302;
  wire _abc_42016_n4303;
  wire _abc_42016_n4304;
  wire _abc_42016_n4305;
  wire _abc_42016_n4306;
  wire _abc_42016_n4307;
  wire _abc_42016_n4308;
  wire _abc_42016_n4309;
  wire _abc_42016_n4310;
  wire _abc_42016_n4311;
  wire _abc_42016_n4312;
  wire _abc_42016_n4314;
  wire _abc_42016_n4315;
  wire _abc_42016_n4316;
  wire _abc_42016_n4317;
  wire _abc_42016_n4318;
  wire _abc_42016_n4319;
  wire _abc_42016_n4320_1;
  wire _abc_42016_n4321;
  wire _abc_42016_n4323;
  wire _abc_42016_n4324;
  wire _abc_42016_n4325;
  wire _abc_42016_n4326;
  wire _abc_42016_n4327;
  wire _abc_42016_n4328;
  wire _abc_42016_n4329;
  wire _abc_42016_n4330;
  wire _abc_42016_n4332;
  wire _abc_42016_n4333;
  wire _abc_42016_n4334;
  wire _abc_42016_n4335;
  wire _abc_42016_n4337;
  wire _abc_42016_n4338;
  wire _abc_42016_n4340;
  wire _abc_42016_n4341;
  wire _abc_42016_n4342;
  wire _abc_42016_n4343;
  wire _abc_42016_n4344;
  wire _abc_42016_n4345;
  wire _abc_42016_n4346;
  wire _abc_42016_n4347;
  wire _abc_42016_n4348;
  wire _abc_42016_n4349;
  wire _abc_42016_n4350;
  wire _abc_42016_n4351;
  wire _abc_42016_n4352;
  wire _abc_42016_n4353;
  wire _abc_42016_n4354;
  wire _abc_42016_n4355;
  wire _abc_42016_n4356;
  wire _abc_42016_n4357;
  wire _abc_42016_n4359;
  wire _abc_42016_n4360;
  wire _abc_42016_n4361;
  wire _abc_42016_n4362;
  wire _abc_42016_n4363;
  wire _abc_42016_n4364;
  wire _abc_42016_n4365;
  wire _abc_42016_n4366;
  wire _abc_42016_n4367;
  wire _abc_42016_n4368;
  wire _abc_42016_n4369;
  wire _abc_42016_n4370;
  wire _abc_42016_n4372;
  wire _abc_42016_n4373;
  wire _abc_42016_n4374;
  wire _abc_42016_n4375;
  wire _abc_42016_n4376;
  wire _abc_42016_n4377;
  wire _abc_42016_n4378;
  wire _abc_42016_n4379;
  wire _abc_42016_n4380;
  wire _abc_42016_n4381;
  wire _abc_42016_n4382;
  wire _abc_42016_n4383;
  wire _abc_42016_n4384;
  wire _abc_42016_n4385;
  wire _abc_42016_n4387;
  wire _abc_42016_n4388;
  wire _abc_42016_n4389;
  wire _abc_42016_n4390;
  wire _abc_42016_n4391;
  wire _abc_42016_n4392;
  wire _abc_42016_n4393;
  wire _abc_42016_n4394;
  wire _abc_42016_n4395;
  wire _abc_42016_n4396;
  wire _abc_42016_n4397;
  wire _abc_42016_n4398;
  wire _abc_42016_n4399;
  wire _abc_42016_n4400;
  wire _abc_42016_n4402;
  wire _abc_42016_n4403_1;
  wire _abc_42016_n4404;
  wire _abc_42016_n4405;
  wire _abc_42016_n4406;
  wire _abc_42016_n4407;
  wire _abc_42016_n4408;
  wire _abc_42016_n4409;
  wire _abc_42016_n4410;
  wire _abc_42016_n4411;
  wire _abc_42016_n4412;
  wire _abc_42016_n4414;
  wire _abc_42016_n4415;
  wire _abc_42016_n4416_1;
  wire _abc_42016_n4417;
  wire _abc_42016_n4418;
  wire _abc_42016_n4419;
  wire _abc_42016_n4420;
  wire _abc_42016_n4421;
  wire _abc_42016_n4422;
  wire _abc_42016_n4423;
  wire _abc_42016_n4424;
  wire _abc_42016_n4426;
  wire _abc_42016_n4427;
  wire _abc_42016_n4428;
  wire _abc_42016_n4429;
  wire _abc_42016_n4430;
  wire _abc_42016_n4431_1;
  wire _abc_42016_n4432;
  wire _abc_42016_n4433;
  wire _abc_42016_n4434;
  wire _abc_42016_n4435;
  wire _abc_42016_n4436;
  wire _abc_42016_n4437;
  wire _abc_42016_n4438;
  wire _abc_42016_n4439;
  wire _abc_42016_n4441;
  wire _abc_42016_n4442;
  wire _abc_42016_n4443;
  wire _abc_42016_n4444;
  wire _abc_42016_n4445;
  wire _abc_42016_n4446;
  wire _abc_42016_n4447_1;
  wire _abc_42016_n4448;
  wire _abc_42016_n4449;
  wire _abc_42016_n4450;
  wire _abc_42016_n4451;
  wire _abc_42016_n4452;
  wire _abc_42016_n4453;
  wire _abc_42016_n4454;
  wire _abc_42016_n4455;
  wire _abc_42016_n4456;
  wire _abc_42016_n4458;
  wire _abc_42016_n4459;
  wire _abc_42016_n4460;
  wire _abc_42016_n4461;
  wire _abc_42016_n4463_1;
  wire _abc_42016_n4464;
  wire _abc_42016_n4466;
  wire _abc_42016_n4467;
  wire _abc_42016_n4468;
  wire _abc_42016_n4469;
  wire _abc_42016_n4470;
  wire _abc_42016_n4471;
  wire _abc_42016_n4472;
  wire _abc_42016_n4473;
  wire _abc_42016_n4474;
  wire _abc_42016_n4475;
  wire _abc_42016_n4476;
  wire _abc_42016_n4478;
  wire _abc_42016_n4479_1;
  wire _abc_42016_n4480;
  wire _abc_42016_n4481;
  wire _abc_42016_n4482;
  wire _abc_42016_n4484;
  wire _abc_42016_n4485;
  wire _abc_42016_n4486;
  wire _abc_42016_n4487;
  wire _abc_42016_n4489;
  wire _abc_42016_n4490;
  wire _abc_42016_n4491;
  wire _abc_42016_n4492;
  wire _abc_42016_n4494_1;
  wire _abc_42016_n4495;
  wire _abc_42016_n4496;
  wire _abc_42016_n4497;
  wire _abc_42016_n4499;
  wire _abc_42016_n4500;
  wire _abc_42016_n4501;
  wire _abc_42016_n4502;
  wire _abc_42016_n4504;
  wire _abc_42016_n4505;
  wire _abc_42016_n4506;
  wire _abc_42016_n4507;
  wire _abc_42016_n4509_1;
  wire _abc_42016_n4510;
  wire _abc_42016_n4511;
  wire _abc_42016_n4512;
  wire _abc_42016_n4514;
  wire _abc_42016_n4515;
  wire _abc_42016_n4516;
  wire _abc_42016_n4517;
  wire _abc_42016_n4519;
  wire _abc_42016_n4520;
  wire _abc_42016_n4521;
  wire _abc_42016_n4523;
  wire _abc_42016_n4524_1;
  wire _abc_42016_n4525;
  wire _abc_42016_n4527;
  wire _abc_42016_n4528;
  wire _abc_42016_n4529;
  wire _abc_42016_n4531;
  wire _abc_42016_n4532;
  wire _abc_42016_n4533;
  wire _abc_42016_n4535;
  wire _abc_42016_n4536;
  wire _abc_42016_n4537;
  wire _abc_42016_n4538;
  wire _abc_42016_n4540;
  wire _abc_42016_n4541;
  wire _abc_42016_n4542;
  wire _abc_42016_n4544;
  wire _abc_42016_n4545;
  wire _abc_42016_n4546;
  wire _abc_42016_n4548;
  wire _abc_42016_n4549;
  wire _abc_42016_n4550;
  wire _abc_42016_n4551;
  wire _abc_42016_n4552;
  wire _abc_42016_n4553;
  wire _abc_42016_n4554_1;
  wire _abc_42016_n4555;
  wire _abc_42016_n4556;
  wire _abc_42016_n4557;
  wire _abc_42016_n4558;
  wire _abc_42016_n4559;
  wire _abc_42016_n4560;
  wire _abc_42016_n4561;
  wire _abc_42016_n4562;
  wire _abc_42016_n4563;
  wire _abc_42016_n4564;
  wire _abc_42016_n4565;
  wire _abc_42016_n4566;
  wire _abc_42016_n4567;
  wire _abc_42016_n4568;
  wire _abc_42016_n4569;
  wire _abc_42016_n4570_1;
  wire _abc_42016_n4571;
  wire _abc_42016_n4572;
  wire _abc_42016_n4573;
  wire _abc_42016_n4574;
  wire _abc_42016_n4575;
  wire _abc_42016_n4576;
  wire _abc_42016_n4577;
  wire _abc_42016_n4578;
  wire _abc_42016_n4579;
  wire _abc_42016_n4580;
  wire _abc_42016_n4581;
  wire _abc_42016_n4582;
  wire _abc_42016_n4583;
  wire _abc_42016_n4584;
  wire _abc_42016_n4585_1;
  wire _abc_42016_n4586;
  wire _abc_42016_n4587;
  wire _abc_42016_n4588;
  wire _abc_42016_n4589;
  wire _abc_42016_n4590;
  wire _abc_42016_n4591;
  wire _abc_42016_n4592;
  wire _abc_42016_n4593;
  wire _abc_42016_n4594;
  wire _abc_42016_n4595;
  wire _abc_42016_n4596;
  wire _abc_42016_n4597;
  wire _abc_42016_n4598;
  wire _abc_42016_n4599;
  wire _abc_42016_n4600_1;
  wire _abc_42016_n4601;
  wire _abc_42016_n4602;
  wire _abc_42016_n4603;
  wire _abc_42016_n4604;
  wire _abc_42016_n4605;
  wire _abc_42016_n4606;
  wire _abc_42016_n4607;
  wire _abc_42016_n4608;
  wire _abc_42016_n4609;
  wire _abc_42016_n4610;
  wire _abc_42016_n4611;
  wire _abc_42016_n4612;
  wire _abc_42016_n4613;
  wire _abc_42016_n4614;
  wire _abc_42016_n4615_1;
  wire _abc_42016_n4616;
  wire _abc_42016_n4617;
  wire _abc_42016_n4618;
  wire _abc_42016_n4619;
  wire _abc_42016_n4620;
  wire _abc_42016_n4621;
  wire _abc_42016_n4622;
  wire _abc_42016_n4623;
  wire _abc_42016_n4624;
  wire _abc_42016_n4625;
  wire _abc_42016_n4626;
  wire _abc_42016_n4627;
  wire _abc_42016_n4628;
  wire _abc_42016_n4629;
  wire _abc_42016_n4630;
  wire _abc_42016_n4631_1;
  wire _abc_42016_n4632_1;
  wire _abc_42016_n4633;
  wire _abc_42016_n4634;
  wire _abc_42016_n4635;
  wire _abc_42016_n4636;
  wire _abc_42016_n4637;
  wire _abc_42016_n4638;
  wire _abc_42016_n4639;
  wire _abc_42016_n4640;
  wire _abc_42016_n4641;
  wire _abc_42016_n4642;
  wire _abc_42016_n4643;
  wire _abc_42016_n4644;
  wire _abc_42016_n4645;
  wire _abc_42016_n4646_1;
  wire _abc_42016_n4647;
  wire _abc_42016_n4648;
  wire _abc_42016_n4649;
  wire _abc_42016_n4650_1;
  wire _abc_42016_n4651;
  wire _abc_42016_n4652;
  wire _abc_42016_n4653;
  wire _abc_42016_n4654_1;
  wire _abc_42016_n4655;
  wire _abc_42016_n4656;
  wire _abc_42016_n4657_1;
  wire _abc_42016_n4658;
  wire _abc_42016_n4659;
  wire _abc_42016_n4660;
  wire _abc_42016_n4661_1;
  wire _abc_42016_n4662;
  wire _abc_42016_n4663;
  wire _abc_42016_n4664;
  wire _abc_42016_n4665;
  wire _abc_42016_n4666_1;
  wire _abc_42016_n4667;
  wire _abc_42016_n4668_1;
  wire _abc_42016_n4669;
  wire _abc_42016_n4670_1;
  wire _abc_42016_n4671;
  wire _abc_42016_n4672_1;
  wire _abc_42016_n4673;
  wire _abc_42016_n4674_1;
  wire _abc_42016_n4675;
  wire _abc_42016_n4676_1;
  wire _abc_42016_n4677;
  wire _abc_42016_n4678_1;
  wire _abc_42016_n4679;
  wire _abc_42016_n4680_1;
  wire _abc_42016_n4681;
  wire _abc_42016_n4682;
  wire _abc_42016_n4683;
  wire _abc_42016_n4684_1;
  wire _abc_42016_n4685;
  wire _abc_42016_n4686;
  wire _abc_42016_n4687;
  wire _abc_42016_n4688_1;
  wire _abc_42016_n4689_1;
  wire _abc_42016_n4690;
  wire _abc_42016_n4691;
  wire _abc_42016_n4692;
  wire _abc_42016_n4693;
  wire _abc_42016_n4694;
  wire _abc_42016_n4696;
  wire _abc_42016_n4697;
  wire _abc_42016_n4698_1;
  wire _abc_42016_n4699;
  wire _abc_42016_n4701;
  wire _abc_42016_n4702;
  wire _abc_42016_n4703;
  wire _abc_42016_n4704;
  wire _abc_42016_n4705_1;
  wire _abc_42016_n4706;
  wire _abc_42016_n4708;
  wire _abc_42016_n4709;
  wire _abc_42016_n4710;
  wire _abc_42016_n4711_1;
  wire _abc_42016_n4712;
  wire _abc_42016_n4713_1;
  wire _abc_42016_n4714;
  wire _abc_42016_n4715;
  wire _abc_42016_n4716;
  wire _abc_42016_n4717_1;
  wire _abc_42016_n4719_1;
  wire _abc_42016_n4720;
  wire _abc_42016_n4721;
  wire _abc_42016_n4722;
  wire _abc_42016_n4723_1;
  wire _abc_42016_n4724;
  wire _abc_42016_n4725_1;
  wire _abc_42016_n4726;
  wire _abc_42016_n4727;
  wire _abc_42016_n4728;
  wire _abc_42016_n4730;
  wire _abc_42016_n4731_1;
  wire _abc_42016_n4732;
  wire _abc_42016_n4733;
  wire _abc_42016_n4735_1;
  wire _abc_42016_n4736;
  wire _abc_42016_n4737_1;
  wire _abc_42016_n4738;
  wire _abc_42016_n4739;
  wire _abc_42016_n501;
  wire _abc_42016_n502;
  wire _abc_42016_n503;
  wire _abc_42016_n504;
  wire _abc_42016_n505;
  wire _abc_42016_n506;
  wire _abc_42016_n507;
  wire _abc_42016_n508;
  wire _abc_42016_n509;
  wire _abc_42016_n510;
  wire _abc_42016_n511;
  wire _abc_42016_n512;
  wire _abc_42016_n513;
  wire _abc_42016_n514;
  wire _abc_42016_n515;
  wire _abc_42016_n516;
  wire _abc_42016_n517;
  wire _abc_42016_n518_1;
  wire _abc_42016_n519;
  wire _abc_42016_n520;
  wire _abc_42016_n521;
  wire _abc_42016_n522;
  wire _abc_42016_n523_1;
  wire _abc_42016_n524_1;
  wire _abc_42016_n525;
  wire _abc_42016_n526_1;
  wire _abc_42016_n527;
  wire _abc_42016_n528_1;
  wire _abc_42016_n529;
  wire _abc_42016_n530;
  wire _abc_42016_n531;
  wire _abc_42016_n532_1;
  wire _abc_42016_n533;
  wire _abc_42016_n534_1;
  wire _abc_42016_n535;
  wire _abc_42016_n536;
  wire _abc_42016_n537_1;
  wire _abc_42016_n538_1;
  wire _abc_42016_n539;
  wire _abc_42016_n540;
  wire _abc_42016_n541;
  wire _abc_42016_n542;
  wire _abc_42016_n543;
  wire _abc_42016_n544_1;
  wire _abc_42016_n545_1;
  wire _abc_42016_n546;
  wire _abc_42016_n547;
  wire _abc_42016_n548;
  wire _abc_42016_n549;
  wire _abc_42016_n550;
  wire _abc_42016_n551;
  wire _abc_42016_n552;
  wire _abc_42016_n553;
  wire _abc_42016_n554;
  wire _abc_42016_n555;
  wire _abc_42016_n556;
  wire _abc_42016_n557;
  wire _abc_42016_n558;
  wire _abc_42016_n559;
  wire _abc_42016_n560;
  wire _abc_42016_n561;
  wire _abc_42016_n562;
  wire _abc_42016_n563;
  wire _abc_42016_n564;
  wire _abc_42016_n565;
  wire _abc_42016_n566;
  wire _abc_42016_n567;
  wire _abc_42016_n568;
  wire _abc_42016_n569;
  wire _abc_42016_n570;
  wire _abc_42016_n571;
  wire _abc_42016_n572;
  wire _abc_42016_n573;
  wire _abc_42016_n574;
  wire _abc_42016_n575;
  wire _abc_42016_n576_1;
  wire _abc_42016_n577;
  wire _abc_42016_n578;
  wire _abc_42016_n579;
  wire _abc_42016_n580;
  wire _abc_42016_n581_1;
  wire _abc_42016_n582_1;
  wire _abc_42016_n583;
  wire _abc_42016_n584_1;
  wire _abc_42016_n585;
  wire _abc_42016_n586;
  wire _abc_42016_n587;
  wire _abc_42016_n588_1;
  wire _abc_42016_n589;
  wire _abc_42016_n590;
  wire _abc_42016_n591;
  wire _abc_42016_n592_1;
  wire _abc_42016_n593;
  wire _abc_42016_n594_1;
  wire _abc_42016_n595;
  wire _abc_42016_n596;
  wire _abc_42016_n597_1;
  wire _abc_42016_n598_1;
  wire _abc_42016_n599;
  wire _abc_42016_n600;
  wire _abc_42016_n601;
  wire _abc_42016_n602;
  wire _abc_42016_n603;
  wire _abc_42016_n604_1;
  wire _abc_42016_n605_1;
  wire _abc_42016_n606;
  wire _abc_42016_n607;
  wire _abc_42016_n608;
  wire _abc_42016_n609;
  wire _abc_42016_n610;
  wire _abc_42016_n611;
  wire _abc_42016_n612;
  wire _abc_42016_n613;
  wire _abc_42016_n614;
  wire _abc_42016_n615;
  wire _abc_42016_n616;
  wire _abc_42016_n617;
  wire _abc_42016_n618;
  wire _abc_42016_n619;
  wire _abc_42016_n620;
  wire _abc_42016_n621;
  wire _abc_42016_n622;
  wire _abc_42016_n623;
  wire _abc_42016_n624;
  wire _abc_42016_n625;
  wire _abc_42016_n626;
  wire _abc_42016_n627;
  wire _abc_42016_n628;
  wire _abc_42016_n629;
  wire _abc_42016_n630;
  wire _abc_42016_n631;
  wire _abc_42016_n632;
  wire _abc_42016_n633;
  wire _abc_42016_n634;
  wire _abc_42016_n635;
  wire _abc_42016_n636;
  wire _abc_42016_n637;
  wire _abc_42016_n638;
  wire _abc_42016_n639;
  wire _abc_42016_n640;
  wire _abc_42016_n641;
  wire _abc_42016_n642;
  wire _abc_42016_n643_1;
  wire _abc_42016_n644;
  wire _abc_42016_n645;
  wire _abc_42016_n646;
  wire _abc_42016_n647;
  wire _abc_42016_n648_1;
  wire _abc_42016_n649_1;
  wire _abc_42016_n650;
  wire _abc_42016_n651_1;
  wire _abc_42016_n652;
  wire _abc_42016_n653;
  wire _abc_42016_n654;
  wire _abc_42016_n655_1;
  wire _abc_42016_n656;
  wire _abc_42016_n657;
  wire _abc_42016_n658;
  wire _abc_42016_n659_1;
  wire _abc_42016_n660;
  wire _abc_42016_n661_1;
  wire _abc_42016_n662;
  wire _abc_42016_n663;
  wire _abc_42016_n664_1;
  wire _abc_42016_n665_1;
  wire _abc_42016_n666;
  wire _abc_42016_n667;
  wire _abc_42016_n668;
  wire _abc_42016_n669;
  wire _abc_42016_n670;
  wire _abc_42016_n671_1;
  wire _abc_42016_n672_1;
  wire _abc_42016_n673;
  wire _abc_42016_n674;
  wire _abc_42016_n675;
  wire _abc_42016_n676;
  wire _abc_42016_n677;
  wire _abc_42016_n678;
  wire _abc_42016_n679;
  wire _abc_42016_n680;
  wire _abc_42016_n681;
  wire _abc_42016_n682;
  wire _abc_42016_n683;
  wire _abc_42016_n684;
  wire _abc_42016_n685;
  wire _abc_42016_n686;
  wire _abc_42016_n687;
  wire _abc_42016_n688;
  wire _abc_42016_n689;
  wire _abc_42016_n690;
  wire _abc_42016_n691;
  wire _abc_42016_n692;
  wire _abc_42016_n693;
  wire _abc_42016_n694;
  wire _abc_42016_n695;
  wire _abc_42016_n696;
  wire _abc_42016_n697;
  wire _abc_42016_n698;
  wire _abc_42016_n699;
  wire _abc_42016_n701;
  wire _abc_42016_n702_1;
  wire _abc_42016_n703;
  wire _abc_42016_n704;
  wire _abc_42016_n705;
  wire _abc_42016_n706;
  wire _abc_42016_n707_1;
  wire _abc_42016_n708;
  wire _abc_42016_n709;
  wire _abc_42016_n710;
  wire _abc_42016_n711;
  wire _abc_42016_n712;
  wire _abc_42016_n713;
  wire _abc_42016_n714;
  wire _abc_42016_n715;
  wire _abc_42016_n716;
  wire _abc_42016_n717;
  wire _abc_42016_n718;
  wire _abc_42016_n719;
  wire _abc_42016_n720;
  wire _abc_42016_n721;
  wire _abc_42016_n722;
  wire _abc_42016_n723;
  wire _abc_42016_n724;
  wire _abc_42016_n725;
  wire _abc_42016_n726;
  wire _abc_42016_n727;
  wire _abc_42016_n728;
  wire _abc_42016_n729;
  wire _abc_42016_n730;
  wire _abc_42016_n731;
  wire _abc_42016_n732;
  wire _abc_42016_n733;
  wire _abc_42016_n734;
  wire _abc_42016_n735;
  wire _abc_42016_n736;
  wire _abc_42016_n737;
  wire _abc_42016_n738;
  wire _abc_42016_n739;
  wire _abc_42016_n740;
  wire _abc_42016_n741;
  wire _abc_42016_n743;
  wire _abc_42016_n744;
  wire _abc_42016_n745;
  wire _abc_42016_n746;
  wire _abc_42016_n747;
  wire _abc_42016_n748;
  wire _abc_42016_n749;
  wire _abc_42016_n750;
  wire _abc_42016_n751;
  wire _abc_42016_n752;
  wire _abc_42016_n753;
  wire _abc_42016_n754;
  wire _abc_42016_n755;
  wire _abc_42016_n756;
  wire _abc_42016_n757;
  wire _abc_42016_n758;
  wire _abc_42016_n759;
  wire _abc_42016_n760;
  wire _abc_42016_n761;
  wire _abc_42016_n762;
  wire _abc_42016_n763_1;
  wire _abc_42016_n764;
  wire _abc_42016_n765;
  wire _abc_42016_n766;
  wire _abc_42016_n767;
  wire _abc_42016_n768;
  wire _abc_42016_n769;
  wire _abc_42016_n770;
  wire _abc_42016_n771;
  wire _abc_42016_n772;
  wire _abc_42016_n773;
  wire _abc_42016_n774;
  wire _abc_42016_n775;
  wire _abc_42016_n776;
  wire _abc_42016_n777;
  wire _abc_42016_n778_1;
  wire _abc_42016_n779;
  wire _abc_42016_n780;
  wire _abc_42016_n781;
  wire _abc_42016_n782;
  wire _abc_42016_n783;
  wire _abc_42016_n784;
  wire _abc_42016_n785;
  wire _abc_42016_n786;
  wire _abc_42016_n787;
  wire _abc_42016_n789;
  wire _abc_42016_n790;
  wire _abc_42016_n791_1;
  wire _abc_42016_n792;
  wire _abc_42016_n793;
  wire _abc_42016_n794;
  wire _abc_42016_n795;
  wire _abc_42016_n796;
  wire _abc_42016_n797;
  wire _abc_42016_n798;
  wire _abc_42016_n799;
  wire _abc_42016_n800;
  wire _abc_42016_n801;
  wire _abc_42016_n802;
  wire _abc_42016_n803;
  wire _abc_42016_n804;
  wire _abc_42016_n805;
  wire _abc_42016_n806;
  wire _abc_42016_n807;
  wire _abc_42016_n808;
  wire _abc_42016_n809;
  wire _abc_42016_n810_1;
  wire _abc_42016_n811;
  wire _abc_42016_n812;
  wire _abc_42016_n813;
  wire _abc_42016_n814;
  wire _abc_42016_n815;
  wire _abc_42016_n816;
  wire _abc_42016_n817;
  wire _abc_42016_n818;
  wire _abc_42016_n819;
  wire _abc_42016_n820;
  wire _abc_42016_n821;
  wire _abc_42016_n822;
  wire _abc_42016_n823;
  wire _abc_42016_n824;
  wire _abc_42016_n825;
  wire _abc_42016_n826_1;
  wire _abc_42016_n827;
  wire _abc_42016_n828;
  wire _abc_42016_n829;
  wire _abc_42016_n830;
  wire _abc_42016_n831;
  wire _abc_42016_n832;
  wire _abc_42016_n834;
  wire _abc_42016_n835;
  wire _abc_42016_n836;
  wire _abc_42016_n837;
  wire _abc_42016_n838;
  wire _abc_42016_n839;
  wire _abc_42016_n840;
  wire _abc_42016_n841;
  wire _abc_42016_n842;
  wire _abc_42016_n843;
  wire _abc_42016_n844;
  wire _abc_42016_n845;
  wire _abc_42016_n846;
  wire _abc_42016_n847;
  wire _abc_42016_n848;
  wire _abc_42016_n849;
  wire _abc_42016_n850;
  wire _abc_42016_n851_1;
  wire _abc_42016_n852;
  wire _abc_42016_n853;
  wire _abc_42016_n854;
  wire _abc_42016_n855;
  wire _abc_42016_n856;
  wire _abc_42016_n857;
  wire _abc_42016_n858;
  wire _abc_42016_n859;
  wire _abc_42016_n860;
  wire _abc_42016_n861;
  wire _abc_42016_n862;
  wire _abc_42016_n863;
  wire _abc_42016_n864;
  wire _abc_42016_n865;
  wire _abc_42016_n866;
  wire _abc_42016_n867_1;
  wire _abc_42016_n868;
  wire _abc_42016_n869;
  wire _abc_42016_n870;
  wire _abc_42016_n872;
  wire _abc_42016_n873;
  wire _abc_42016_n874;
  wire _abc_42016_n875;
  wire _abc_42016_n876;
  wire _abc_42016_n877;
  wire _abc_42016_n878;
  wire _abc_42016_n879;
  wire _abc_42016_n880;
  wire _abc_42016_n881;
  wire _abc_42016_n882;
  wire _abc_42016_n883;
  wire _abc_42016_n884;
  wire _abc_42016_n885;
  wire _abc_42016_n886;
  wire _abc_42016_n887;
  wire _abc_42016_n888;
  wire _abc_42016_n889_1;
  wire _abc_42016_n890;
  wire _abc_42016_n891;
  wire _abc_42016_n892;
  wire _abc_42016_n893;
  wire _abc_42016_n894;
  wire _abc_42016_n895;
  wire _abc_42016_n896;
  wire _abc_42016_n897;
  wire _abc_42016_n898;
  wire _abc_42016_n899;
  wire _abc_42016_n900;
  wire _abc_42016_n901;
  wire _abc_42016_n902;
  wire _abc_42016_n903;
  wire _abc_42016_n904;
  wire _abc_42016_n905;
  wire _abc_42016_n906;
  wire _abc_42016_n907;
  wire _abc_42016_n908;
  wire _abc_42016_n909;
  wire _abc_42016_n910_1;
  wire _abc_42016_n911;
  wire _abc_42016_n913;
  wire _abc_42016_n914;
  wire _abc_42016_n915;
  wire _abc_42016_n916;
  wire _abc_42016_n917;
  wire _abc_42016_n918;
  wire _abc_42016_n919;
  wire _abc_42016_n920;
  wire _abc_42016_n921;
  wire _abc_42016_n922;
  wire _abc_42016_n923;
  wire _abc_42016_n924;
  wire _abc_42016_n925;
  wire _abc_42016_n926;
  wire _abc_42016_n927;
  wire _abc_42016_n928;
  wire _abc_42016_n929;
  wire _abc_42016_n930;
  wire _abc_42016_n931;
  wire _abc_42016_n932;
  wire _abc_42016_n933;
  wire _abc_42016_n934;
  wire _abc_42016_n935;
  wire _abc_42016_n936;
  wire _abc_42016_n937;
  wire _abc_42016_n938;
  wire _abc_42016_n939;
  wire _abc_42016_n940;
  wire _abc_42016_n941_1;
  wire _abc_42016_n942;
  wire _abc_42016_n943;
  wire _abc_42016_n944;
  wire _abc_42016_n945;
  wire _abc_42016_n946;
  wire _abc_42016_n947;
  wire _abc_42016_n949;
  wire _abc_42016_n950;
  wire _abc_42016_n951;
  wire _abc_42016_n952;
  wire _abc_42016_n953;
  wire _abc_42016_n954;
  wire _abc_42016_n955;
  wire _abc_42016_n956;
  wire _abc_42016_n957_1;
  wire _abc_42016_n958;
  wire _abc_42016_n959;
  wire _abc_42016_n960;
  wire _abc_42016_n961;
  wire _abc_42016_n962;
  wire _abc_42016_n963;
  wire _abc_42016_n964;
  wire _abc_42016_n965;
  wire _abc_42016_n966;
  wire _abc_42016_n967;
  wire _abc_42016_n968;
  wire _abc_42016_n969;
  wire _abc_42016_n970;
  wire _abc_42016_n971;
  wire _abc_42016_n972;
  wire _abc_42016_n973;
  wire _abc_42016_n974;
  wire _abc_42016_n975;
  wire _abc_42016_n976;
  wire _abc_42016_n977;
  wire _abc_42016_n978;
  wire _abc_42016_n979_1;
  wire _abc_42016_n980;
  wire _abc_42016_n981;
  wire _abc_42016_n982;
  wire _abc_42016_n983;
  wire _abc_42016_n984;
  wire _abc_42016_n985;
  wire _abc_42016_n987;
  wire _abc_42016_n988;
  wire _abc_42016_n989;
  wire _abc_42016_n990;
  wire _abc_42016_n991;
  wire _abc_42016_n992;
  wire _abc_42016_n993;
  wire _abc_42016_n994;
  wire _abc_42016_n995;
  wire _abc_42016_n996;
  wire _abc_42016_n997;
  wire _abc_42016_n998;
  wire _abc_42016_n999;
  wire _auto_iopadmap_cc_313_execute_46257_0_;
  wire _auto_iopadmap_cc_313_execute_46257_10_;
  wire _auto_iopadmap_cc_313_execute_46257_11_;
  wire _auto_iopadmap_cc_313_execute_46257_12_;
  wire _auto_iopadmap_cc_313_execute_46257_13_;
  wire _auto_iopadmap_cc_313_execute_46257_14_;
  wire _auto_iopadmap_cc_313_execute_46257_15_;
  wire _auto_iopadmap_cc_313_execute_46257_1_;
  wire _auto_iopadmap_cc_313_execute_46257_2_;
  wire _auto_iopadmap_cc_313_execute_46257_3_;
  wire _auto_iopadmap_cc_313_execute_46257_4_;
  wire _auto_iopadmap_cc_313_execute_46257_5_;
  wire _auto_iopadmap_cc_313_execute_46257_6_;
  wire _auto_iopadmap_cc_313_execute_46257_7_;
  wire _auto_iopadmap_cc_313_execute_46257_8_;
  wire _auto_iopadmap_cc_313_execute_46257_9_;
  wire _auto_iopadmap_cc_313_execute_46274;
  wire _auto_iopadmap_cc_313_execute_46276;
  wire _auto_iopadmap_cc_313_execute_46278;
  wire _auto_iopadmap_cc_313_execute_46280;
  wire _auto_iopadmap_cc_313_execute_46282;
  output \addr[0] ;
  output \addr[10] ;
  output \addr[11] ;
  output \addr[12] ;
  output \addr[13] ;
  output \addr[14] ;
  output \addr[15] ;
  output \addr[1] ;
  output \addr[2] ;
  output \addr[3] ;
  output \addr[4] ;
  output \addr[5] ;
  output \addr[6] ;
  output \addr[7] ;
  output \addr[8] ;
  output \addr[9] ;
  wire addr_0__FF_INPUT;
  wire addr_10__FF_INPUT;
  wire addr_11__FF_INPUT;
  wire addr_12__FF_INPUT;
  wire addr_13__FF_INPUT;
  wire addr_14__FF_INPUT;
  wire addr_15__FF_INPUT;
  wire addr_1__FF_INPUT;
  wire addr_2__FF_INPUT;
  wire addr_3__FF_INPUT;
  wire addr_4__FF_INPUT;
  wire addr_5__FF_INPUT;
  wire addr_6__FF_INPUT;
  wire addr_7__FF_INPUT;
  wire addr_8__FF_INPUT;
  wire addr_9__FF_INPUT;
  wire alu__abc_41682_n100;
  wire alu__abc_41682_n101;
  wire alu__abc_41682_n102;
  wire alu__abc_41682_n103;
  wire alu__abc_41682_n104;
  wire alu__abc_41682_n105;
  wire alu__abc_41682_n106;
  wire alu__abc_41682_n107;
  wire alu__abc_41682_n108;
  wire alu__abc_41682_n109;
  wire alu__abc_41682_n110;
  wire alu__abc_41682_n111;
  wire alu__abc_41682_n112;
  wire alu__abc_41682_n113;
  wire alu__abc_41682_n114;
  wire alu__abc_41682_n115;
  wire alu__abc_41682_n116;
  wire alu__abc_41682_n117;
  wire alu__abc_41682_n118;
  wire alu__abc_41682_n119;
  wire alu__abc_41682_n120;
  wire alu__abc_41682_n121;
  wire alu__abc_41682_n122;
  wire alu__abc_41682_n123;
  wire alu__abc_41682_n124_1;
  wire alu__abc_41682_n125;
  wire alu__abc_41682_n126;
  wire alu__abc_41682_n127;
  wire alu__abc_41682_n128;
  wire alu__abc_41682_n129;
  wire alu__abc_41682_n130;
  wire alu__abc_41682_n131;
  wire alu__abc_41682_n132;
  wire alu__abc_41682_n133;
  wire alu__abc_41682_n134;
  wire alu__abc_41682_n135;
  wire alu__abc_41682_n136;
  wire alu__abc_41682_n137;
  wire alu__abc_41682_n138;
  wire alu__abc_41682_n139;
  wire alu__abc_41682_n140;
  wire alu__abc_41682_n141;
  wire alu__abc_41682_n142;
  wire alu__abc_41682_n143;
  wire alu__abc_41682_n144;
  wire alu__abc_41682_n145;
  wire alu__abc_41682_n146;
  wire alu__abc_41682_n147;
  wire alu__abc_41682_n148;
  wire alu__abc_41682_n149;
  wire alu__abc_41682_n150;
  wire alu__abc_41682_n151;
  wire alu__abc_41682_n152;
  wire alu__abc_41682_n153;
  wire alu__abc_41682_n154;
  wire alu__abc_41682_n155;
  wire alu__abc_41682_n156;
  wire alu__abc_41682_n157;
  wire alu__abc_41682_n158;
  wire alu__abc_41682_n159;
  wire alu__abc_41682_n160;
  wire alu__abc_41682_n161;
  wire alu__abc_41682_n162;
  wire alu__abc_41682_n163;
  wire alu__abc_41682_n164;
  wire alu__abc_41682_n165;
  wire alu__abc_41682_n166;
  wire alu__abc_41682_n167;
  wire alu__abc_41682_n168;
  wire alu__abc_41682_n169_1;
  wire alu__abc_41682_n170;
  wire alu__abc_41682_n171;
  wire alu__abc_41682_n172;
  wire alu__abc_41682_n173;
  wire alu__abc_41682_n174;
  wire alu__abc_41682_n175;
  wire alu__abc_41682_n176;
  wire alu__abc_41682_n177;
  wire alu__abc_41682_n178;
  wire alu__abc_41682_n179;
  wire alu__abc_41682_n180;
  wire alu__abc_41682_n181;
  wire alu__abc_41682_n182;
  wire alu__abc_41682_n183;
  wire alu__abc_41682_n184;
  wire alu__abc_41682_n185;
  wire alu__abc_41682_n186;
  wire alu__abc_41682_n187;
  wire alu__abc_41682_n188;
  wire alu__abc_41682_n189;
  wire alu__abc_41682_n190;
  wire alu__abc_41682_n191;
  wire alu__abc_41682_n192;
  wire alu__abc_41682_n193;
  wire alu__abc_41682_n194;
  wire alu__abc_41682_n195;
  wire alu__abc_41682_n196;
  wire alu__abc_41682_n198;
  wire alu__abc_41682_n199;
  wire alu__abc_41682_n200;
  wire alu__abc_41682_n201;
  wire alu__abc_41682_n202;
  wire alu__abc_41682_n203;
  wire alu__abc_41682_n204;
  wire alu__abc_41682_n205;
  wire alu__abc_41682_n206;
  wire alu__abc_41682_n207;
  wire alu__abc_41682_n208;
  wire alu__abc_41682_n209;
  wire alu__abc_41682_n210;
  wire alu__abc_41682_n211;
  wire alu__abc_41682_n212;
  wire alu__abc_41682_n213;
  wire alu__abc_41682_n214;
  wire alu__abc_41682_n215;
  wire alu__abc_41682_n216;
  wire alu__abc_41682_n217;
  wire alu__abc_41682_n218;
  wire alu__abc_41682_n219;
  wire alu__abc_41682_n220;
  wire alu__abc_41682_n221;
  wire alu__abc_41682_n222;
  wire alu__abc_41682_n223;
  wire alu__abc_41682_n224;
  wire alu__abc_41682_n225;
  wire alu__abc_41682_n226;
  wire alu__abc_41682_n227;
  wire alu__abc_41682_n228;
  wire alu__abc_41682_n229;
  wire alu__abc_41682_n230;
  wire alu__abc_41682_n231;
  wire alu__abc_41682_n232;
  wire alu__abc_41682_n233;
  wire alu__abc_41682_n234;
  wire alu__abc_41682_n235;
  wire alu__abc_41682_n236;
  wire alu__abc_41682_n237;
  wire alu__abc_41682_n238;
  wire alu__abc_41682_n239;
  wire alu__abc_41682_n240;
  wire alu__abc_41682_n241;
  wire alu__abc_41682_n242;
  wire alu__abc_41682_n243;
  wire alu__abc_41682_n244;
  wire alu__abc_41682_n245;
  wire alu__abc_41682_n246;
  wire alu__abc_41682_n247;
  wire alu__abc_41682_n248;
  wire alu__abc_41682_n249;
  wire alu__abc_41682_n250;
  wire alu__abc_41682_n251;
  wire alu__abc_41682_n252;
  wire alu__abc_41682_n253;
  wire alu__abc_41682_n254;
  wire alu__abc_41682_n255;
  wire alu__abc_41682_n256;
  wire alu__abc_41682_n257;
  wire alu__abc_41682_n258;
  wire alu__abc_41682_n259_1;
  wire alu__abc_41682_n260;
  wire alu__abc_41682_n261;
  wire alu__abc_41682_n262;
  wire alu__abc_41682_n263;
  wire alu__abc_41682_n264;
  wire alu__abc_41682_n265;
  wire alu__abc_41682_n266_1;
  wire alu__abc_41682_n267;
  wire alu__abc_41682_n268_1;
  wire alu__abc_41682_n269;
  wire alu__abc_41682_n270_1;
  wire alu__abc_41682_n271_1;
  wire alu__abc_41682_n272;
  wire alu__abc_41682_n273_1;
  wire alu__abc_41682_n274;
  wire alu__abc_41682_n275_1;
  wire alu__abc_41682_n276;
  wire alu__abc_41682_n277_1;
  wire alu__abc_41682_n278;
  wire alu__abc_41682_n279_1;
  wire alu__abc_41682_n280_1;
  wire alu__abc_41682_n281;
  wire alu__abc_41682_n282;
  wire alu__abc_41682_n283;
  wire alu__abc_41682_n284;
  wire alu__abc_41682_n285;
  wire alu__abc_41682_n286_1;
  wire alu__abc_41682_n287;
  wire alu__abc_41682_n288;
  wire alu__abc_41682_n289;
  wire alu__abc_41682_n290;
  wire alu__abc_41682_n291;
  wire alu__abc_41682_n292;
  wire alu__abc_41682_n293;
  wire alu__abc_41682_n294;
  wire alu__abc_41682_n295;
  wire alu__abc_41682_n296;
  wire alu__abc_41682_n297;
  wire alu__abc_41682_n298;
  wire alu__abc_41682_n299;
  wire alu__abc_41682_n300;
  wire alu__abc_41682_n301;
  wire alu__abc_41682_n302;
  wire alu__abc_41682_n303;
  wire alu__abc_41682_n304;
  wire alu__abc_41682_n305;
  wire alu__abc_41682_n306;
  wire alu__abc_41682_n307;
  wire alu__abc_41682_n308;
  wire alu__abc_41682_n309;
  wire alu__abc_41682_n310;
  wire alu__abc_41682_n311;
  wire alu__abc_41682_n312;
  wire alu__abc_41682_n313;
  wire alu__abc_41682_n314_1;
  wire alu__abc_41682_n315;
  wire alu__abc_41682_n316;
  wire alu__abc_41682_n317;
  wire alu__abc_41682_n318;
  wire alu__abc_41682_n319;
  wire alu__abc_41682_n320;
  wire alu__abc_41682_n321;
  wire alu__abc_41682_n322;
  wire alu__abc_41682_n323;
  wire alu__abc_41682_n324;
  wire alu__abc_41682_n325;
  wire alu__abc_41682_n326;
  wire alu__abc_41682_n327;
  wire alu__abc_41682_n328;
  wire alu__abc_41682_n329;
  wire alu__abc_41682_n330;
  wire alu__abc_41682_n331;
  wire alu__abc_41682_n332;
  wire alu__abc_41682_n333;
  wire alu__abc_41682_n334;
  wire alu__abc_41682_n336;
  wire alu__abc_41682_n337;
  wire alu__abc_41682_n339;
  wire alu__abc_41682_n34;
  wire alu__abc_41682_n342;
  wire alu__abc_41682_n344;
  wire alu__abc_41682_n346;
  wire alu__abc_41682_n349;
  wire alu__abc_41682_n35;
  wire alu__abc_41682_n351;
  wire alu__abc_41682_n353;
  wire alu__abc_41682_n354;
  wire alu__abc_41682_n355;
  wire alu__abc_41682_n356;
  wire alu__abc_41682_n357;
  wire alu__abc_41682_n359;
  wire alu__abc_41682_n36;
  wire alu__abc_41682_n360;
  wire alu__abc_41682_n361;
  wire alu__abc_41682_n362;
  wire alu__abc_41682_n363;
  wire alu__abc_41682_n364;
  wire alu__abc_41682_n365;
  wire alu__abc_41682_n37;
  wire alu__abc_41682_n38;
  wire alu__abc_41682_n39;
  wire alu__abc_41682_n40;
  wire alu__abc_41682_n41;
  wire alu__abc_41682_n42;
  wire alu__abc_41682_n43;
  wire alu__abc_41682_n44;
  wire alu__abc_41682_n45_1;
  wire alu__abc_41682_n46_1;
  wire alu__abc_41682_n47;
  wire alu__abc_41682_n48;
  wire alu__abc_41682_n49;
  wire alu__abc_41682_n50_1;
  wire alu__abc_41682_n51;
  wire alu__abc_41682_n52;
  wire alu__abc_41682_n53;
  wire alu__abc_41682_n54;
  wire alu__abc_41682_n55;
  wire alu__abc_41682_n56;
  wire alu__abc_41682_n57;
  wire alu__abc_41682_n58;
  wire alu__abc_41682_n59;
  wire alu__abc_41682_n60;
  wire alu__abc_41682_n61;
  wire alu__abc_41682_n62;
  wire alu__abc_41682_n63;
  wire alu__abc_41682_n64;
  wire alu__abc_41682_n65;
  wire alu__abc_41682_n66;
  wire alu__abc_41682_n67;
  wire alu__abc_41682_n68;
  wire alu__abc_41682_n69;
  wire alu__abc_41682_n70;
  wire alu__abc_41682_n71;
  wire alu__abc_41682_n72;
  wire alu__abc_41682_n73;
  wire alu__abc_41682_n74;
  wire alu__abc_41682_n75;
  wire alu__abc_41682_n76;
  wire alu__abc_41682_n77;
  wire alu__abc_41682_n78;
  wire alu__abc_41682_n79;
  wire alu__abc_41682_n80;
  wire alu__abc_41682_n81;
  wire alu__abc_41682_n82;
  wire alu__abc_41682_n83;
  wire alu__abc_41682_n84;
  wire alu__abc_41682_n85;
  wire alu__abc_41682_n86;
  wire alu__abc_41682_n87;
  wire alu__abc_41682_n88;
  wire alu__abc_41682_n89;
  wire alu__abc_41682_n90;
  wire alu__abc_41682_n91;
  wire alu__abc_41682_n92;
  wire alu__abc_41682_n93;
  wire alu__abc_41682_n94;
  wire alu__abc_41682_n95;
  wire alu__abc_41682_n96;
  wire alu__abc_41682_n97;
  wire alu__abc_41682_n98;
  wire alu__abc_41682_n99;
  wire alu_auxcar;
  wire alu_cin;
  wire alu_cout;
  wire alu_opra_0_;
  wire alu_opra_1_;
  wire alu_opra_2_;
  wire alu_opra_3_;
  wire alu_opra_4_;
  wire alu_opra_5_;
  wire alu_opra_6_;
  wire alu_opra_7_;
  wire alu_oprb_0_;
  wire alu_oprb_1_;
  wire alu_oprb_2_;
  wire alu_oprb_3_;
  wire alu_oprb_4_;
  wire alu_oprb_5_;
  wire alu_oprb_6_;
  wire alu_oprb_7_;
  wire alu_parity;
  wire alu_res_0_;
  wire alu_res_1_;
  wire alu_res_2_;
  wire alu_res_3_;
  wire alu_res_4_;
  wire alu_res_5_;
  wire alu_res_6_;
  wire alu_res_7_;
  wire alu_sel_0_;
  wire alu_sel_1_;
  wire alu_sel_2_;
  wire alu_sout;
  wire alu_zout;
  wire alucin_FF_INPUT;
  wire aluopra_0__FF_INPUT;
  wire aluopra_1__FF_INPUT;
  wire aluopra_2__FF_INPUT;
  wire aluopra_3__FF_INPUT;
  wire aluopra_4__FF_INPUT;
  wire aluopra_5__FF_INPUT;
  wire aluopra_6__FF_INPUT;
  wire aluopra_7__FF_INPUT;
  wire aluoprb_0__FF_INPUT;
  wire aluoprb_1__FF_INPUT;
  wire aluoprb_2__FF_INPUT;
  wire aluoprb_3__FF_INPUT;
  wire aluoprb_4__FF_INPUT;
  wire aluoprb_5__FF_INPUT;
  wire aluoprb_6__FF_INPUT;
  wire aluoprb_7__FF_INPUT;
  wire alusel_0__FF_INPUT;
  wire alusel_1__FF_INPUT;
  wire alusel_2__FF_INPUT;
  wire auxcar;
  wire auxcar_FF_INPUT;
  wire carry;
  wire carry_FF_INPUT;
  input clock;
  input \data[0] ;
  input \data[1] ;
  input \data[2] ;
  input \data[3] ;
  input \data[4] ;
  input \data[5] ;
  input \data[6] ;
  input \data[7] ;
  wire datao_0__FF_INPUT;
  wire datao_1__FF_INPUT;
  wire datao_2__FF_INPUT;
  wire datao_3__FF_INPUT;
  wire datao_4__FF_INPUT;
  wire datao_5__FF_INPUT;
  wire datao_6__FF_INPUT;
  wire datao_7__FF_INPUT;
  wire ei;
  wire ei_FF_INPUT;
  wire eienb;
  wire eienb_FF_INPUT;
  output inta;
  wire inta_FF_INPUT;
  wire intcyc;
  wire intcyc_FF_INPUT;
  input intr;
  wire opcode_0_;
  wire opcode_0__FF_INPUT;
  wire opcode_1_;
  wire opcode_1__FF_INPUT;
  wire opcode_2_;
  wire opcode_2__FF_INPUT;
  wire opcode_3_;
  wire opcode_3__FF_INPUT;
  wire opcode_4_;
  wire opcode_4__FF_INPUT;
  wire opcode_5_;
  wire opcode_5__FF_INPUT;
  wire opcode_6_;
  wire opcode_6__FF_INPUT;
  wire opcode_7_;
  wire opcode_7__FF_INPUT;
  wire parity;
  wire parity_FF_INPUT;
  wire pc_0_;
  wire pc_0__FF_INPUT;
  wire pc_10_;
  wire pc_10__FF_INPUT;
  wire pc_11_;
  wire pc_11__FF_INPUT;
  wire pc_12_;
  wire pc_12__FF_INPUT;
  wire pc_13_;
  wire pc_13__FF_INPUT;
  wire pc_14_;
  wire pc_14__FF_INPUT;
  wire pc_15_;
  wire pc_15__FF_INPUT;
  wire pc_1_;
  wire pc_1__FF_INPUT;
  wire pc_2_;
  wire pc_2__FF_INPUT;
  wire pc_3_;
  wire pc_3__FF_INPUT;
  wire pc_4_;
  wire pc_4__FF_INPUT;
  wire pc_5_;
  wire pc_5__FF_INPUT;
  wire pc_6_;
  wire pc_6__FF_INPUT;
  wire pc_7_;
  wire pc_7__FF_INPUT;
  wire pc_8_;
  wire pc_8__FF_INPUT;
  wire pc_9_;
  wire pc_9__FF_INPUT;
  wire popdes_0_;
  wire popdes_0__FF_INPUT;
  wire popdes_1_;
  wire popdes_1__FF_INPUT;
  wire raddrhold_0_;
  wire raddrhold_0__FF_INPUT;
  wire raddrhold_10_;
  wire raddrhold_10__FF_INPUT;
  wire raddrhold_11_;
  wire raddrhold_11__FF_INPUT;
  wire raddrhold_12_;
  wire raddrhold_12__FF_INPUT;
  wire raddrhold_13_;
  wire raddrhold_13__FF_INPUT;
  wire raddrhold_14_;
  wire raddrhold_14__FF_INPUT;
  wire raddrhold_15_;
  wire raddrhold_15__FF_INPUT;
  wire raddrhold_1_;
  wire raddrhold_1__FF_INPUT;
  wire raddrhold_2_;
  wire raddrhold_2__FF_INPUT;
  wire raddrhold_3_;
  wire raddrhold_3__FF_INPUT;
  wire raddrhold_4_;
  wire raddrhold_4__FF_INPUT;
  wire raddrhold_5_;
  wire raddrhold_5__FF_INPUT;
  wire raddrhold_6_;
  wire raddrhold_6__FF_INPUT;
  wire raddrhold_7_;
  wire raddrhold_7__FF_INPUT;
  wire raddrhold_8_;
  wire raddrhold_8__FF_INPUT;
  wire raddrhold_9_;
  wire raddrhold_9__FF_INPUT;
  wire rdatahold2_0_;
  wire rdatahold2_0__FF_INPUT;
  wire rdatahold2_1_;
  wire rdatahold2_1__FF_INPUT;
  wire rdatahold2_2_;
  wire rdatahold2_2__FF_INPUT;
  wire rdatahold2_3_;
  wire rdatahold2_3__FF_INPUT;
  wire rdatahold2_4_;
  wire rdatahold2_4__FF_INPUT;
  wire rdatahold2_5_;
  wire rdatahold2_5__FF_INPUT;
  wire rdatahold2_6_;
  wire rdatahold2_6__FF_INPUT;
  wire rdatahold2_7_;
  wire rdatahold2_7__FF_INPUT;
  wire rdatahold_0_;
  wire rdatahold_0__FF_INPUT;
  wire rdatahold_1_;
  wire rdatahold_1__FF_INPUT;
  wire rdatahold_2_;
  wire rdatahold_2__FF_INPUT;
  wire rdatahold_3_;
  wire rdatahold_3__FF_INPUT;
  wire rdatahold_4_;
  wire rdatahold_4__FF_INPUT;
  wire rdatahold_5_;
  wire rdatahold_5__FF_INPUT;
  wire rdatahold_6_;
  wire rdatahold_6__FF_INPUT;
  wire rdatahold_7_;
  wire rdatahold_7__FF_INPUT;
  output readio;
  wire readio_FF_INPUT;
  output readmem;
  wire readmem_FF_INPUT;
  wire regd_0_;
  wire regd_0__FF_INPUT;
  wire regd_1_;
  wire regd_1__FF_INPUT;
  wire regd_2_;
  wire regd_2__FF_INPUT;
  wire regfil_0__0_;
  wire regfil_0__1_;
  wire regfil_0__2_;
  wire regfil_0__3_;
  wire regfil_0__4_;
  wire regfil_0__5_;
  wire regfil_0__6_;
  wire regfil_0__7_;
  wire regfil_1__0_;
  wire regfil_1__1_;
  wire regfil_1__2_;
  wire regfil_1__3_;
  wire regfil_1__4_;
  wire regfil_1__5_;
  wire regfil_1__6_;
  wire regfil_1__7_;
  wire regfil_2__0_;
  wire regfil_2__1_;
  wire regfil_2__2_;
  wire regfil_2__3_;
  wire regfil_2__4_;
  wire regfil_2__5_;
  wire regfil_2__6_;
  wire regfil_2__7_;
  wire regfil_3__0_;
  wire regfil_3__1_;
  wire regfil_3__2_;
  wire regfil_3__3_;
  wire regfil_3__4_;
  wire regfil_3__5_;
  wire regfil_3__6_;
  wire regfil_3__7_;
  wire regfil_4__0_;
  wire regfil_4__1_;
  wire regfil_4__2_;
  wire regfil_4__3_;
  wire regfil_4__4_;
  wire regfil_4__5_;
  wire regfil_4__6_;
  wire regfil_4__7_;
  wire regfil_5__0_;
  wire regfil_5__1_;
  wire regfil_5__2_;
  wire regfil_5__3_;
  wire regfil_5__4_;
  wire regfil_5__5_;
  wire regfil_5__6_;
  wire regfil_5__7_;
  wire regfil_6__0_;
  wire regfil_6__1_;
  wire regfil_6__2_;
  wire regfil_6__3_;
  wire regfil_6__4_;
  wire regfil_6__5_;
  wire regfil_6__6_;
  wire regfil_6__7_;
  wire regfil_7__0_;
  wire regfil_7__1_;
  wire regfil_7__2_;
  wire regfil_7__3_;
  wire regfil_7__4_;
  wire regfil_7__5_;
  wire regfil_7__6_;
  wire regfil_7__7_;
  input reset;
  wire sign;
  wire sign_FF_INPUT;
  wire sp_0_;
  wire sp_0__FF_INPUT;
  wire sp_10_;
  wire sp_10__FF_INPUT;
  wire sp_11_;
  wire sp_11__FF_INPUT;
  wire sp_12_;
  wire sp_12__FF_INPUT;
  wire sp_13_;
  wire sp_13__FF_INPUT;
  wire sp_14_;
  wire sp_14__FF_INPUT;
  wire sp_15_;
  wire sp_15__FF_INPUT;
  wire sp_1_;
  wire sp_1__FF_INPUT;
  wire sp_2_;
  wire sp_2__FF_INPUT;
  wire sp_3_;
  wire sp_3__FF_INPUT;
  wire sp_4_;
  wire sp_4__FF_INPUT;
  wire sp_5_;
  wire sp_5__FF_INPUT;
  wire sp_6_;
  wire sp_6__FF_INPUT;
  wire sp_7_;
  wire sp_7__FF_INPUT;
  wire sp_8_;
  wire sp_8__FF_INPUT;
  wire sp_9_;
  wire sp_9__FF_INPUT;
  wire state_0_;
  wire state_1_;
  wire state_2_;
  wire state_3_;
  wire state_4_;
  wire state_5_;
  wire statesel_0_;
  wire statesel_0__FF_INPUT;
  wire statesel_1_;
  wire statesel_1__FF_INPUT;
  wire statesel_2_;
  wire statesel_2__FF_INPUT;
  wire statesel_3_;
  wire statesel_3__FF_INPUT;
  wire statesel_4_;
  wire statesel_4__FF_INPUT;
  wire statesel_5_;
  wire statesel_5__FF_INPUT;
  wire waddrhold_0_;
  wire waddrhold_0__FF_INPUT;
  wire waddrhold_10_;
  wire waddrhold_10__FF_INPUT;
  wire waddrhold_11_;
  wire waddrhold_11__FF_INPUT;
  wire waddrhold_12_;
  wire waddrhold_12__FF_INPUT;
  wire waddrhold_13_;
  wire waddrhold_13__FF_INPUT;
  wire waddrhold_14_;
  wire waddrhold_14__FF_INPUT;
  wire waddrhold_15_;
  wire waddrhold_15__FF_INPUT;
  wire waddrhold_1_;
  wire waddrhold_1__FF_INPUT;
  wire waddrhold_2_;
  wire waddrhold_2__FF_INPUT;
  wire waddrhold_3_;
  wire waddrhold_3__FF_INPUT;
  wire waddrhold_4_;
  wire waddrhold_4__FF_INPUT;
  wire waddrhold_5_;
  wire waddrhold_5__FF_INPUT;
  wire waddrhold_6_;
  wire waddrhold_6__FF_INPUT;
  wire waddrhold_7_;
  wire waddrhold_7__FF_INPUT;
  wire waddrhold_8_;
  wire waddrhold_8__FF_INPUT;
  wire waddrhold_9_;
  wire waddrhold_9__FF_INPUT;
  input waitr;
  wire wdatahold2_0_;
  wire wdatahold2_0__FF_INPUT;
  wire wdatahold2_1_;
  wire wdatahold2_1__FF_INPUT;
  wire wdatahold2_2_;
  wire wdatahold2_2__FF_INPUT;
  wire wdatahold2_3_;
  wire wdatahold2_3__FF_INPUT;
  wire wdatahold2_4_;
  wire wdatahold2_4__FF_INPUT;
  wire wdatahold2_5_;
  wire wdatahold2_5__FF_INPUT;
  wire wdatahold2_6_;
  wire wdatahold2_6__FF_INPUT;
  wire wdatahold2_7_;
  wire wdatahold2_7__FF_INPUT;
  wire wdatahold_0_;
  wire wdatahold_0__FF_INPUT;
  wire wdatahold_1_;
  wire wdatahold_1__FF_INPUT;
  wire wdatahold_2_;
  wire wdatahold_2__FF_INPUT;
  wire wdatahold_3_;
  wire wdatahold_3__FF_INPUT;
  wire wdatahold_4_;
  wire wdatahold_4__FF_INPUT;
  wire wdatahold_5_;
  wire wdatahold_5__FF_INPUT;
  wire wdatahold_6_;
  wire wdatahold_6__FF_INPUT;
  wire wdatahold_7_;
  wire wdatahold_7__FF_INPUT;
  output writeio;
  wire writeio_FF_INPUT;
  output writemem;
  wire writemem_FF_INPUT;
  wire zero;
  wire zero_FF_INPUT;
  AND2X2 AND2X2_1 ( .A(_abc_42016_n624), .B(_abc_42016_n731), .Y(_abc_42016_n732) );
  AND2X2 AND2X2_10 ( .A(_abc_42016_n1048), .B(_abc_42016_n1002), .Y(_abc_42016_n1049) );
  AND2X2 AND2X2_100 ( .A(_abc_42016_n4464), .B(_abc_42016_n4328), .Y(readmem_FF_INPUT) );
  AND2X2 AND2X2_101 ( .A(_abc_42016_n4592), .B(_abc_42016_n4599), .Y(_abc_42016_n4600_1) );
  AND2X2 AND2X2_102 ( .A(_abc_42016_n4621), .B(_abc_42016_n4611), .Y(_abc_42016_n4622) );
  AND2X2 AND2X2_103 ( .A(_abc_42016_n4633), .B(_abc_42016_n4078), .Y(_abc_42016_n4634) );
  AND2X2 AND2X2_104 ( .A(_abc_42016_n4641), .B(_abc_42016_n4645), .Y(_abc_42016_n4646_1) );
  AND2X2 AND2X2_105 ( .A(_abc_42016_n4665), .B(_abc_42016_n4663), .Y(_abc_42016_n4666_1) );
  AND2X2 AND2X2_106 ( .A(_abc_42016_n4684_1), .B(_abc_42016_n4685), .Y(_abc_42016_n4686) );
  AND2X2 AND2X2_107 ( .A(_abc_42016_n4698_1), .B(_abc_42016_n4674_1), .Y(_abc_42016_n4699) );
  AND2X2 AND2X2_108 ( .A(_abc_42016_n4623), .B(_abc_42016_n4337), .Y(_abc_42016_n4720) );
  AND2X2 AND2X2_109 ( .A(alu_oprb_1_), .B(alu_opra_1_), .Y(alu__abc_41682_n35) );
  AND2X2 AND2X2_11 ( .A(_abc_42016_n1103_1), .B(_abc_42016_n1100), .Y(_abc_42016_n1104_1) );
  AND2X2 AND2X2_110 ( .A(alu_oprb_0_), .B(alu_opra_0_), .Y(alu__abc_41682_n37) );
  AND2X2 AND2X2_111 ( .A(alu__abc_41682_n41), .B(alu__abc_41682_n44), .Y(alu__abc_41682_n45_1) );
  AND2X2 AND2X2_112 ( .A(alu__abc_41682_n55), .B(alu__abc_41682_n52), .Y(alu__abc_41682_n57) );
  AND2X2 AND2X2_113 ( .A(alu__abc_41682_n183), .B(alu__abc_41682_n185), .Y(alu__abc_41682_n186) );
  AND2X2 AND2X2_114 ( .A(alu__abc_41682_n222), .B(alu__abc_41682_n213), .Y(alu__abc_41682_n223) );
  AND2X2 AND2X2_115 ( .A(alu__abc_41682_n252), .B(alu__abc_41682_n253), .Y(alu__abc_41682_n254) );
  AND2X2 AND2X2_116 ( .A(alu__abc_41682_n283), .B(alu__abc_41682_n161), .Y(alu__abc_41682_n293) );
  AND2X2 AND2X2_117 ( .A(alu__abc_41682_n330), .B(alu__abc_41682_n337), .Y(alu_zout) );
  AND2X2 AND2X2_118 ( .A(alu__abc_41682_n177), .B(alu__abc_41682_n190), .Y(alu__abc_41682_n361) );
  AND2X2 AND2X2_12 ( .A(_abc_42016_n1125), .B(_abc_42016_n1126), .Y(_abc_42016_n1127) );
  AND2X2 AND2X2_13 ( .A(_abc_42016_n1144), .B(_abc_42016_n1143), .Y(_abc_42016_n1145) );
  AND2X2 AND2X2_14 ( .A(_abc_42016_n1192), .B(_abc_42016_n1193), .Y(_abc_42016_n1194) );
  AND2X2 AND2X2_15 ( .A(_abc_42016_n1188), .B(_abc_42016_n872), .Y(_abc_42016_n1227) );
  AND2X2 AND2X2_16 ( .A(_abc_42016_n1204), .B(_abc_42016_n1241), .Y(_abc_42016_n1242) );
  AND2X2 AND2X2_17 ( .A(_abc_42016_n1275), .B(_abc_42016_n1277), .Y(_abc_42016_n1278) );
  AND2X2 AND2X2_18 ( .A(_abc_42016_n971), .B(_abc_42016_n989), .Y(_abc_42016_n1303) );
  AND2X2 AND2X2_19 ( .A(_abc_42016_n1314), .B(_abc_42016_n1313), .Y(_abc_42016_n1315) );
  AND2X2 AND2X2_2 ( .A(_abc_42016_n767), .B(_abc_42016_n747), .Y(_abc_42016_n768) );
  AND2X2 AND2X2_20 ( .A(_abc_42016_n1468), .B(_abc_42016_n1460), .Y(_abc_42016_n1469) );
  AND2X2 AND2X2_21 ( .A(_abc_42016_n649_1), .B(_abc_42016_n1709), .Y(_abc_42016_n1710) );
  AND2X2 AND2X2_22 ( .A(_abc_42016_n1729_1), .B(_abc_42016_n1730), .Y(_abc_42016_n1731) );
  AND2X2 AND2X2_23 ( .A(_abc_42016_n1924), .B(_abc_42016_n529), .Y(_abc_42016_n1930) );
  AND2X2 AND2X2_24 ( .A(_abc_42016_n1980), .B(_abc_42016_n1910), .Y(_abc_42016_n1981) );
  AND2X2 AND2X2_25 ( .A(_abc_42016_n1993), .B(_abc_42016_n1910), .Y(_abc_42016_n1994) );
  AND2X2 AND2X2_26 ( .A(_abc_42016_n2036), .B(alu_parity), .Y(_abc_42016_n2039) );
  AND2X2 AND2X2_27 ( .A(_abc_42016_n2036), .B(_abc_42016_n529), .Y(_abc_42016_n2051) );
  AND2X2 AND2X2_28 ( .A(_abc_42016_n2105), .B(_abc_42016_n2104), .Y(_abc_42016_n2106) );
  AND2X2 AND2X2_29 ( .A(_abc_42016_n2114), .B(_abc_42016_n2112), .Y(_abc_42016_n2115_1) );
  AND2X2 AND2X2_3 ( .A(_abc_42016_n784), .B(_abc_42016_n701), .Y(_abc_42016_n785) );
  AND2X2 AND2X2_30 ( .A(_abc_42016_n2123_1), .B(_abc_42016_n2121), .Y(_abc_42016_n2124_1) );
  AND2X2 AND2X2_31 ( .A(_abc_42016_n2132_1), .B(_abc_42016_n2130), .Y(_abc_42016_n2133) );
  AND2X2 AND2X2_32 ( .A(_abc_42016_n2160), .B(_abc_42016_n2159), .Y(_abc_42016_n2161) );
  AND2X2 AND2X2_33 ( .A(_abc_42016_n2181), .B(_abc_42016_n2180), .Y(_abc_42016_n2182) );
  AND2X2 AND2X2_34 ( .A(_abc_42016_n2192), .B(_abc_42016_n2191), .Y(_abc_42016_n2193) );
  AND2X2 AND2X2_35 ( .A(_abc_42016_n2199), .B(_abc_42016_n2197), .Y(_abc_42016_n2200) );
  AND2X2 AND2X2_36 ( .A(_abc_42016_n2295), .B(_abc_42016_n559), .Y(_abc_42016_n2296_1) );
  AND2X2 AND2X2_37 ( .A(_abc_42016_n2431), .B(_abc_42016_n2432_1), .Y(_abc_42016_n2433) );
  AND2X2 AND2X2_38 ( .A(_abc_42016_n2337), .B(_abc_42016_n2454), .Y(_abc_42016_n2455_1) );
  AND2X2 AND2X2_39 ( .A(_abc_42016_n2559), .B(_abc_42016_n2560), .Y(_abc_42016_n2561) );
  AND2X2 AND2X2_4 ( .A(_abc_42016_n790), .B(_abc_42016_n791_1), .Y(_abc_42016_n792) );
  AND2X2 AND2X2_40 ( .A(_abc_42016_n2564), .B(_abc_42016_n530), .Y(_abc_42016_n2565) );
  AND2X2 AND2X2_41 ( .A(_abc_42016_n1438), .B(_abc_42016_n2573), .Y(_abc_42016_n2574) );
  AND2X2 AND2X2_42 ( .A(_abc_42016_n2602), .B(_abc_42016_n2537), .Y(_abc_42016_n2603) );
  AND2X2 AND2X2_43 ( .A(_abc_42016_n1362), .B(_abc_42016_n2650), .Y(_abc_42016_n2651) );
  AND2X2 AND2X2_44 ( .A(_abc_42016_n1364), .B(_abc_42016_n2686), .Y(_abc_42016_n2687) );
  AND2X2 AND2X2_45 ( .A(_abc_42016_n2299), .B(_abc_42016_n967), .Y(_abc_42016_n2708) );
  AND2X2 AND2X2_46 ( .A(_abc_42016_n1366), .B(_abc_42016_n2723), .Y(_abc_42016_n2724) );
  AND2X2 AND2X2_47 ( .A(_abc_42016_n2747_1), .B(_abc_42016_n2766), .Y(_abc_42016_n2767_1) );
  AND2X2 AND2X2_48 ( .A(_abc_42016_n2977), .B(_abc_42016_n2428), .Y(_abc_42016_n2978) );
  AND2X2 AND2X2_49 ( .A(_abc_42016_n3058_1), .B(_abc_42016_n673), .Y(_abc_42016_n3059) );
  AND2X2 AND2X2_5 ( .A(_abc_42016_n830), .B(_abc_42016_n826_1), .Y(_abc_42016_n831) );
  AND2X2 AND2X2_50 ( .A(_abc_42016_n3112), .B(_abc_42016_n1848), .Y(_abc_42016_n3115) );
  AND2X2 AND2X2_51 ( .A(_abc_42016_n3147_1), .B(waddrhold_5_), .Y(_abc_42016_n3170_1) );
  AND2X2 AND2X2_52 ( .A(_abc_42016_n3180), .B(_abc_42016_n3181), .Y(_abc_42016_n3182) );
  AND2X2 AND2X2_53 ( .A(_abc_42016_n3256), .B(_abc_42016_n3258), .Y(_abc_42016_n3259) );
  AND2X2 AND2X2_54 ( .A(_abc_42016_n3269), .B(_abc_42016_n3270), .Y(_abc_42016_n3271) );
  AND2X2 AND2X2_55 ( .A(_abc_42016_n3273), .B(_abc_42016_n673), .Y(_abc_42016_n3274) );
  AND2X2 AND2X2_56 ( .A(_abc_42016_n3319_1), .B(_abc_42016_n3320), .Y(_abc_42016_n3321) );
  AND2X2 AND2X2_57 ( .A(_abc_42016_n3343), .B(_abc_42016_n673), .Y(_abc_42016_n3344) );
  AND2X2 AND2X2_58 ( .A(_abc_42016_n3368_1), .B(_abc_42016_n673), .Y(_abc_42016_n3369_1) );
  AND2X2 AND2X2_59 ( .A(_abc_42016_n1346), .B(_abc_42016_n1574), .Y(_abc_42016_n3371) );
  AND2X2 AND2X2_6 ( .A(_abc_42016_n837), .B(_abc_42016_n856), .Y(_abc_42016_n857) );
  AND2X2 AND2X2_60 ( .A(_abc_42016_n3501), .B(_abc_42016_n3505), .Y(_abc_42016_n3506) );
  AND2X2 AND2X2_61 ( .A(_abc_42016_n3509), .B(_abc_42016_n3508), .Y(_abc_42016_n3510_1) );
  AND2X2 AND2X2_62 ( .A(_abc_42016_n3522), .B(_abc_42016_n3521), .Y(_abc_42016_n3523) );
  AND2X2 AND2X2_63 ( .A(_abc_42016_n3534), .B(_abc_42016_n3532), .Y(_abc_42016_n3535) );
  AND2X2 AND2X2_64 ( .A(_abc_42016_n3545), .B(_abc_42016_n2256), .Y(_abc_42016_n3546) );
  AND2X2 AND2X2_65 ( .A(_abc_42016_n3607), .B(_abc_42016_n3608), .Y(_abc_42016_n3609) );
  AND2X2 AND2X2_66 ( .A(_abc_42016_n3642), .B(_abc_42016_n3643), .Y(_abc_42016_n3644) );
  AND2X2 AND2X2_67 ( .A(_abc_42016_n3653), .B(_abc_42016_n3657), .Y(_abc_42016_n3658) );
  AND2X2 AND2X2_68 ( .A(_abc_42016_n3672), .B(_abc_42016_n3678), .Y(_abc_42016_n3679) );
  AND2X2 AND2X2_69 ( .A(_abc_42016_n3679), .B(_abc_42016_n2347_1), .Y(_abc_42016_n3680) );
  AND2X2 AND2X2_7 ( .A(_abc_42016_n879), .B(_abc_42016_n701), .Y(_abc_42016_n880) );
  AND2X2 AND2X2_70 ( .A(_abc_42016_n3710), .B(_abc_42016_n3708), .Y(_abc_42016_n3711) );
  AND2X2 AND2X2_71 ( .A(_abc_42016_n3729), .B(_abc_42016_n3722), .Y(_abc_42016_n3730) );
  AND2X2 AND2X2_72 ( .A(_abc_42016_n3758), .B(_abc_42016_n2101), .Y(_abc_42016_n3780) );
  AND2X2 AND2X2_73 ( .A(_abc_42016_n3763), .B(_abc_42016_n2101), .Y(_abc_42016_n3783) );
  AND2X2 AND2X2_74 ( .A(_abc_42016_n3810), .B(_abc_42016_n3811), .Y(_abc_42016_n3812) );
  AND2X2 AND2X2_75 ( .A(_abc_42016_n2170), .B(_abc_42016_n2165), .Y(_abc_42016_n3849) );
  AND2X2 AND2X2_76 ( .A(_abc_42016_n3876), .B(_abc_42016_n2138), .Y(_abc_42016_n3877) );
  AND2X2 AND2X2_77 ( .A(_abc_42016_n3883), .B(_abc_42016_n2172_1), .Y(_abc_42016_n3884) );
  AND2X2 AND2X2_78 ( .A(_abc_42016_n2140_1), .B(_abc_42016_n1023), .Y(_abc_42016_n3932) );
  AND2X2 AND2X2_79 ( .A(_abc_42016_n3907), .B(regfil_4__4_), .Y(_abc_42016_n3933) );
  AND2X2 AND2X2_8 ( .A(_abc_42016_n624), .B(_abc_42016_n902), .Y(_abc_42016_n903) );
  AND2X2 AND2X2_80 ( .A(_abc_42016_n2206), .B(_abc_42016_n2188), .Y(_abc_42016_n3939) );
  AND2X2 AND2X2_81 ( .A(_abc_42016_n2207), .B(_abc_42016_n1036), .Y(_abc_42016_n3940) );
  AND2X2 AND2X2_82 ( .A(_abc_42016_n2173), .B(_abc_42016_n2156), .Y(_abc_42016_n3942) );
  AND2X2 AND2X2_83 ( .A(_abc_42016_n2174), .B(_abc_42016_n1031_1), .Y(_abc_42016_n3943) );
  AND2X2 AND2X2_84 ( .A(_abc_42016_n2207), .B(_abc_42016_n2186), .Y(_abc_42016_n3965) );
  AND2X2 AND2X2_85 ( .A(_abc_42016_n2175), .B(_abc_42016_n2150), .Y(_abc_42016_n3997) );
  AND2X2 AND2X2_86 ( .A(_abc_42016_n4041_1), .B(_abc_42016_n1010), .Y(_abc_42016_n4042) );
  AND2X2 AND2X2_87 ( .A(_abc_42016_n4099), .B(_abc_42016_n2090), .Y(_abc_42016_n4100) );
  AND2X2 AND2X2_88 ( .A(_abc_42016_n4111), .B(_abc_42016_n4105), .Y(_abc_42016_n4112) );
  AND2X2 AND2X2_89 ( .A(_abc_42016_n4118), .B(_abc_42016_n4121), .Y(_abc_42016_n4122) );
  AND2X2 AND2X2_9 ( .A(_abc_42016_n597_1), .B(_abc_42016_n591), .Y(_abc_42016_n987) );
  AND2X2 AND2X2_90 ( .A(_abc_42016_n4093), .B(_abc_42016_n673), .Y(_abc_42016_n4127) );
  AND2X2 AND2X2_91 ( .A(_abc_42016_n2674), .B(_abc_42016_n4199), .Y(_abc_42016_n4200) );
  AND2X2 AND2X2_92 ( .A(_abc_42016_n1389), .B(_abc_42016_n4211), .Y(_abc_42016_n4212) );
  AND2X2 AND2X2_93 ( .A(_abc_42016_n4279), .B(_abc_42016_n4132), .Y(_abc_42016_n4280) );
  AND2X2 AND2X2_94 ( .A(_abc_42016_n4289), .B(_abc_42016_n559), .Y(_abc_42016_n4290) );
  AND2X2 AND2X2_95 ( .A(_abc_42016_n4303), .B(_abc_42016_n4132), .Y(_abc_42016_n4304) );
  AND2X2 AND2X2_96 ( .A(_abc_42016_n4347), .B(_abc_42016_n557), .Y(_abc_42016_n4348) );
  AND2X2 AND2X2_97 ( .A(_abc_42016_n4365), .B(_abc_42016_n4361), .Y(_abc_42016_n4366) );
  AND2X2 AND2X2_98 ( .A(_abc_42016_n4435), .B(_abc_42016_n4436), .Y(_abc_42016_n4437) );
  AND2X2 AND2X2_99 ( .A(_abc_42016_n4445), .B(_abc_42016_n4444), .Y(_abc_42016_n4446) );
  AOI21X1 AOI21X1_1 ( .A(_abc_42016_n549), .B(_abc_42016_n535), .C(_abc_42016_n528_1), .Y(_abc_42016_n550) );
  AOI21X1 AOI21X1_10 ( .A(_abc_42016_n799), .B(_abc_42016_n538_1), .C(_abc_42016_n802), .Y(_abc_42016_n803) );
  AOI21X1 AOI21X1_100 ( .A(_abc_42016_n609), .B(_abc_42016_n1729_1), .C(_abc_42016_n659_1), .Y(_abc_42016_n1755) );
  AOI21X1 AOI21X1_101 ( .A(_abc_42016_n651_1), .B(_abc_42016_n1755), .C(_abc_42016_n1754), .Y(_abc_42016_n1756) );
  AOI21X1 AOI21X1_102 ( .A(_abc_42016_n641), .B(_abc_42016_n651_1), .C(_abc_42016_n1758), .Y(_abc_42016_n1759) );
  AOI21X1 AOI21X1_103 ( .A(_abc_42016_n664_1), .B(_abc_42016_n1767_1), .C(_abc_42016_n1768), .Y(_abc_42016_n1769) );
  AOI21X1 AOI21X1_104 ( .A(_abc_42016_n691), .B(_abc_42016_n1643), .C(_abc_42016_n1769), .Y(_abc_36783_n3638) );
  AOI21X1 AOI21X1_105 ( .A(_abc_42016_n769), .B(_abc_42016_n1767_1), .C(_abc_42016_n1774), .Y(_abc_42016_n1775) );
  AOI21X1 AOI21X1_106 ( .A(_abc_42016_n691), .B(_abc_42016_n1684), .C(_abc_42016_n1775), .Y(_abc_36783_n3642) );
  AOI21X1 AOI21X1_107 ( .A(_abc_42016_n858), .B(_abc_42016_n1767_1), .C(_abc_42016_n1780), .Y(_abc_42016_n1781) );
  AOI21X1 AOI21X1_108 ( .A(_abc_42016_n691), .B(_abc_42016_n1725), .C(_abc_42016_n1781), .Y(_abc_36783_n3646) );
  AOI21X1 AOI21X1_109 ( .A(_abc_42016_n1783_1), .B(_abc_42016_n895), .C(_abc_42016_n691), .Y(_abc_42016_n1784_1) );
  AOI21X1 AOI21X1_11 ( .A(_abc_42016_n601), .B(_abc_42016_n795), .C(_abc_42016_n691), .Y(_abc_42016_n820) );
  AOI21X1 AOI21X1_110 ( .A(_abc_42016_n919), .B(_abc_42016_n1738), .C(_abc_42016_n1787), .Y(_abc_42016_n1788) );
  AOI21X1 AOI21X1_111 ( .A(_abc_42016_n696), .B(regfil_4__6_), .C(_abc_42016_n689), .Y(_abc_42016_n1791) );
  AOI21X1 AOI21X1_112 ( .A(_abc_42016_n1793), .B(_abc_42016_n689), .C(_abc_42016_n690), .Y(_abc_42016_n1794) );
  AOI21X1 AOI21X1_113 ( .A(rdatahold_6_), .B(_abc_42016_n1639_1), .C(_abc_42016_n692), .Y(_abc_42016_n1796) );
  AOI21X1 AOI21X1_114 ( .A(rdatahold_7_), .B(_abc_42016_n1639_1), .C(_abc_42016_n692), .Y(_abc_42016_n1800) );
  AOI21X1 AOI21X1_115 ( .A(_abc_42016_n1787), .B(_abc_42016_n1803), .C(_abc_42016_n964), .Y(_abc_42016_n1804) );
  AOI21X1 AOI21X1_116 ( .A(_abc_42016_n964), .B(_abc_42016_n1806), .C(_abc_42016_n1804), .Y(_abc_42016_n1807) );
  AOI21X1 AOI21X1_117 ( .A(_abc_42016_n663), .B(_abc_42016_n1815), .C(_abc_42016_n1816), .Y(_abc_36783_n3731) );
  AOI21X1 AOI21X1_118 ( .A(_abc_42016_n857), .B(_abc_42016_n1815), .C(_abc_42016_n1824), .Y(_abc_36783_n3735) );
  AOI21X1 AOI21X1_119 ( .A(_abc_42016_n559), .B(_abc_42016_n1837_1), .C(_abc_42016_n1836), .Y(_abc_42016_n1838_1) );
  AOI21X1 AOI21X1_12 ( .A(_abc_42016_n834), .B(_abc_42016_n815), .C(_abc_42016_n835), .Y(_abc_42016_n836) );
  AOI21X1 AOI21X1_120 ( .A(opcode_4_), .B(_abc_42016_n1851), .C(_abc_42016_n1836), .Y(_abc_42016_n1852) );
  AOI21X1 AOI21X1_121 ( .A(_abc_42016_n559), .B(_abc_42016_n1847), .C(_abc_42016_n1853), .Y(_abc_42016_n1854) );
  AOI21X1 AOI21X1_122 ( .A(_abc_42016_n1846), .B(_abc_42016_n1836), .C(_abc_42016_n1854), .Y(alusel_1__FF_INPUT) );
  AOI21X1 AOI21X1_123 ( .A(alu_oprb_0_), .B(_abc_42016_n1863), .C(_abc_42016_n1865), .Y(_abc_42016_n1866) );
  AOI21X1 AOI21X1_124 ( .A(_abc_42016_n557), .B(_abc_42016_n1880), .C(_abc_42016_n1875_1), .Y(_abc_42016_n1881) );
  AOI21X1 AOI21X1_125 ( .A(_abc_42016_n1905_1), .B(_abc_42016_n1906), .C(_abc_42016_n1907), .Y(_abc_42016_n1908) );
  AOI21X1 AOI21X1_126 ( .A(_abc_42016_n1917), .B(regfil_7__0_), .C(_abc_42016_n530), .Y(_abc_42016_n1918) );
  AOI21X1 AOI21X1_127 ( .A(alu_opra_1_), .B(_abc_42016_n1933), .C(_abc_42016_n1944), .Y(_abc_42016_n1945) );
  AOI21X1 AOI21X1_128 ( .A(alu_opra_3_), .B(_abc_42016_n1933), .C(_abc_42016_n1970), .Y(_abc_42016_n1971) );
  AOI21X1 AOI21X1_129 ( .A(regfil_1__4_), .B(_abc_42016_n1915), .C(_abc_42016_n1978), .Y(_abc_42016_n1979) );
  AOI21X1 AOI21X1_13 ( .A(_abc_42016_n607), .B(_abc_42016_n840), .C(_abc_42016_n855), .Y(_abc_42016_n856) );
  AOI21X1 AOI21X1_130 ( .A(alu_opra_4_), .B(_abc_42016_n1933), .C(_abc_42016_n1983), .Y(_abc_42016_n1984) );
  AOI21X1 AOI21X1_131 ( .A(_abc_42016_n1911), .B(regfil_4__5_), .C(_abc_42016_n530), .Y(_abc_42016_n1990) );
  AOI21X1 AOI21X1_132 ( .A(regfil_6__5_), .B(_abc_42016_n532_1), .C(_abc_42016_n1991), .Y(_abc_42016_n1992) );
  AOI21X1 AOI21X1_133 ( .A(alu_opra_5_), .B(_abc_42016_n1933), .C(_abc_42016_n1996), .Y(_abc_42016_n1997) );
  AOI21X1 AOI21X1_134 ( .A(_abc_42016_n1917), .B(regfil_3__6_), .C(opcode_5_), .Y(_abc_42016_n2000) );
  AOI21X1 AOI21X1_135 ( .A(regfil_1__6_), .B(_abc_42016_n1915), .C(_abc_42016_n2001), .Y(_abc_42016_n2002) );
  AOI21X1 AOI21X1_136 ( .A(alu_opra_6_), .B(_abc_42016_n1933), .C(_abc_42016_n2007), .Y(_abc_42016_n2008) );
  AOI21X1 AOI21X1_137 ( .A(regfil_2__7_), .B(_abc_42016_n532_1), .C(_abc_42016_n2016), .Y(_abc_42016_n2017) );
  AOI21X1 AOI21X1_138 ( .A(_abc_42016_n2017), .B(_abc_42016_n2015), .C(_abc_42016_n1909_1), .Y(_abc_42016_n2018) );
  AOI21X1 AOI21X1_139 ( .A(alu_opra_7_), .B(_abc_42016_n1933), .C(_abc_42016_n2020), .Y(_abc_42016_n2021) );
  AOI21X1 AOI21X1_14 ( .A(_abc_42016_n783), .B(_abc_42016_n795), .C(_abc_42016_n861), .Y(_abc_42016_n865) );
  AOI21X1 AOI21X1_140 ( .A(ei), .B(intr), .C(_abc_42016_n2024), .Y(_abc_42016_n2025) );
  AOI21X1 AOI21X1_141 ( .A(regfil_7__7_), .B(_abc_42016_n2069), .C(_abc_42016_n2070), .Y(_abc_42016_n2071) );
  AOI21X1 AOI21X1_142 ( .A(rdatahold2_4_), .B(_abc_42016_n2043), .C(_abc_42016_n2075), .Y(_abc_42016_n2076) );
  AOI21X1 AOI21X1_143 ( .A(_abc_42016_n2092), .B(_abc_42016_n1860), .C(_abc_42016_n548), .Y(_abc_42016_n2215) );
  AOI21X1 AOI21X1_144 ( .A(_abc_42016_n2047), .B(carry), .C(_abc_42016_n2220), .Y(_abc_42016_n2221) );
  AOI21X1 AOI21X1_145 ( .A(_abc_42016_n2293), .B(_abc_42016_n2280), .C(_abc_42016_n2292), .Y(_abc_42016_n2294) );
  AOI21X1 AOI21X1_146 ( .A(_abc_42016_n2259), .B(_abc_42016_n2336), .C(_abc_42016_n2341), .Y(_abc_42016_n2342) );
  AOI21X1 AOI21X1_147 ( .A(_abc_42016_n1848), .B(_abc_42016_n2344), .C(_abc_42016_n1863), .Y(_abc_42016_n2345) );
  AOI21X1 AOI21X1_148 ( .A(opcode_4_), .B(_abc_42016_n2347_1), .C(_abc_42016_n2309), .Y(_abc_42016_n2348_1) );
  AOI21X1 AOI21X1_149 ( .A(_abc_42016_n2373_1), .B(_abc_42016_n2301), .C(_abc_42016_n2369), .Y(_abc_42016_n2374) );
  AOI21X1 AOI21X1_15 ( .A(rdatahold2_4_), .B(_abc_42016_n694), .C(_abc_42016_n869), .Y(_abc_42016_n870) );
  AOI21X1 AOI21X1_150 ( .A(_abc_42016_n2281), .B(opcode_5_), .C(_abc_42016_n1841), .Y(_abc_42016_n2377) );
  AOI21X1 AOI21X1_151 ( .A(_abc_42016_n2375), .B(_abc_42016_n2379), .C(_abc_42016_n560), .Y(_abc_42016_n2380) );
  AOI21X1 AOI21X1_152 ( .A(_abc_42016_n2288), .B(_abc_42016_n2369), .C(_abc_42016_n548), .Y(_abc_42016_n2381) );
  AOI21X1 AOI21X1_153 ( .A(statesel_2_), .B(_abc_42016_n2339), .C(_abc_42016_n2278), .Y(_abc_42016_n2390) );
  AOI21X1 AOI21X1_154 ( .A(_abc_42016_n2384), .B(_abc_42016_n675), .C(_abc_42016_n2391), .Y(_abc_42016_n2392) );
  AOI21X1 AOI21X1_155 ( .A(_abc_42016_n2394_1), .B(_abc_42016_n2280), .C(_abc_42016_n2395), .Y(_abc_42016_n2396) );
  AOI21X1 AOI21X1_156 ( .A(_abc_42016_n2347_1), .B(opcode_5_), .C(_abc_42016_n1841), .Y(_abc_42016_n2397) );
  AOI21X1 AOI21X1_157 ( .A(_abc_42016_n2394_1), .B(_abc_42016_n2288), .C(_abc_42016_n2399), .Y(_abc_42016_n2400) );
  AOI21X1 AOI21X1_158 ( .A(statesel_3_), .B(_abc_42016_n2326), .C(_abc_42016_n2321), .Y(_abc_42016_n2401) );
  AOI21X1 AOI21X1_159 ( .A(_abc_42016_n2336), .B(_abc_42016_n2410), .C(_abc_42016_n2414_1), .Y(_abc_42016_n2415) );
  AOI21X1 AOI21X1_16 ( .A(_abc_42016_n898), .B(_abc_42016_n564), .C(_abc_42016_n899), .Y(_abc_42016_n900) );
  AOI21X1 AOI21X1_160 ( .A(_abc_42016_n2329), .B(_abc_42016_n2419), .C(_abc_42016_n2420_1), .Y(_abc_42016_n2421) );
  AOI21X1 AOI21X1_161 ( .A(_abc_42016_n2289), .B(_abc_42016_n559), .C(_abc_42016_n2402_1), .Y(_abc_42016_n2422) );
  AOI21X1 AOI21X1_162 ( .A(_abc_42016_n2283), .B(_abc_42016_n559), .C(_abc_42016_n2403), .Y(_abc_42016_n2432_1) );
  AOI21X1 AOI21X1_163 ( .A(_abc_42016_n2336), .B(_abc_42016_n2442), .C(_abc_42016_n2443), .Y(_abc_42016_n2444_1) );
  AOI21X1 AOI21X1_164 ( .A(_abc_42016_n2340), .B(_abc_42016_n2441_1), .C(_abc_42016_n2446), .Y(_abc_42016_n2453) );
  AOI21X1 AOI21X1_165 ( .A(carry), .B(_abc_42016_n1003), .C(_abc_42016_n2502), .Y(_abc_42016_n2503) );
  AOI21X1 AOI21X1_166 ( .A(regfil_5__0_), .B(_abc_42016_n1426), .C(_abc_42016_n2504), .Y(_abc_42016_n2505) );
  AOI21X1 AOI21X1_167 ( .A(_abc_42016_n559), .B(_abc_42016_n1347), .C(_abc_42016_n2359), .Y(_abc_42016_n2509) );
  AOI21X1 AOI21X1_168 ( .A(_abc_42016_n2512), .B(_abc_42016_n2511), .C(_abc_42016_n1851), .Y(_abc_42016_n2513) );
  AOI21X1 AOI21X1_169 ( .A(_abc_42016_n637), .B(_abc_42016_n2299), .C(_abc_42016_n2514), .Y(_abc_42016_n2515) );
  AOI21X1 AOI21X1_17 ( .A(_abc_42016_n890), .B(_abc_42016_n607), .C(_abc_42016_n907), .Y(_abc_42016_n908) );
  AOI21X1 AOI21X1_170 ( .A(_abc_42016_n2508), .B(_abc_42016_n2515), .C(_abc_42016_n2516), .Y(_abc_42016_n2517_1) );
  AOI21X1 AOI21X1_171 ( .A(_abc_42016_n1508), .B(_abc_42016_n2526), .C(_abc_42016_n2532), .Y(_abc_42016_n2533) );
  AOI21X1 AOI21X1_172 ( .A(_abc_42016_n731), .B(_abc_42016_n2299), .C(_abc_42016_n2545), .Y(_abc_42016_n2546) );
  AOI21X1 AOI21X1_173 ( .A(_abc_42016_n2548_1), .B(_abc_42016_n1851), .C(_abc_42016_n548), .Y(_abc_42016_n2549) );
  AOI21X1 AOI21X1_174 ( .A(_abc_42016_n2547_1), .B(_abc_42016_n2549), .C(_abc_42016_n2551), .Y(_abc_42016_n2552) );
  AOI21X1 AOI21X1_175 ( .A(_abc_42016_n1381), .B(_abc_42016_n2572), .C(_abc_42016_n2571), .Y(_abc_42016_n2573) );
  AOI21X1 AOI21X1_176 ( .A(_abc_42016_n761), .B(_abc_42016_n2299), .C(_abc_42016_n2578_1), .Y(_abc_42016_n2579_1) );
  AOI21X1 AOI21X1_177 ( .A(_abc_42016_n2575), .B(_abc_42016_n2579_1), .C(_abc_42016_n2558), .Y(_abc_42016_n2580) );
  AOI21X1 AOI21X1_178 ( .A(_abc_42016_n2583), .B(_abc_42016_n1851), .C(_abc_42016_n548), .Y(_abc_42016_n2584) );
  AOI21X1 AOI21X1_179 ( .A(_abc_42016_n2582), .B(_abc_42016_n2584), .C(_abc_42016_n2499), .Y(_abc_42016_n2585) );
  AOI21X1 AOI21X1_18 ( .A(_abc_42016_n913), .B(_abc_42016_n885), .C(_abc_42016_n931), .Y(_abc_42016_n932) );
  AOI21X1 AOI21X1_180 ( .A(_abc_42016_n2512), .B(_abc_42016_n2607), .C(_abc_42016_n1851), .Y(_abc_42016_n2608_1) );
  AOI21X1 AOI21X1_181 ( .A(_abc_42016_n2587), .B(_abc_42016_n1851), .C(_abc_42016_n548), .Y(_abc_42016_n2610) );
  AOI21X1 AOI21X1_182 ( .A(regfil_7__4_), .B(_abc_42016_n669), .C(_abc_42016_n1245), .Y(_abc_42016_n2640_1) );
  AOI21X1 AOI21X1_183 ( .A(_abc_42016_n2299), .B(_abc_42016_n850), .C(_abc_42016_n2641), .Y(_abc_42016_n2642) );
  AOI21X1 AOI21X1_184 ( .A(_abc_42016_n2619), .B(_abc_42016_n1851), .C(_abc_42016_n548), .Y(_abc_42016_n2644) );
  AOI21X1 AOI21X1_185 ( .A(_abc_42016_n2643), .B(_abc_42016_n2644), .C(_abc_42016_n2645), .Y(_abc_42016_n2646) );
  AOI21X1 AOI21X1_186 ( .A(regfil_5__5_), .B(_abc_42016_n1426), .C(_abc_42016_n2657), .Y(_abc_42016_n2658) );
  AOI21X1 AOI21X1_187 ( .A(_abc_42016_n1438), .B(_abc_42016_n2651), .C(_abc_42016_n2659), .Y(_abc_42016_n2660) );
  AOI21X1 AOI21X1_188 ( .A(_abc_42016_n902), .B(_abc_42016_n2299), .C(_abc_42016_n2665), .Y(_abc_42016_n2666) );
  AOI21X1 AOI21X1_189 ( .A(_abc_42016_n2648), .B(_abc_42016_n1851), .C(_abc_42016_n548), .Y(_abc_42016_n2668) );
  AOI21X1 AOI21X1_19 ( .A(rdatahold_6_), .B(_abc_42016_n751), .C(_abc_42016_n932), .Y(_abc_42016_n933) );
  AOI21X1 AOI21X1_190 ( .A(_abc_42016_n2512), .B(_abc_42016_n2692), .C(_abc_42016_n1851), .Y(_abc_42016_n2693) );
  AOI21X1 AOI21X1_191 ( .A(_abc_42016_n2694), .B(_abc_42016_n2584), .C(_abc_42016_n2697), .Y(_abc_42016_n2698) );
  AOI21X1 AOI21X1_192 ( .A(alu_res_7_), .B(_abc_42016_n2518_1), .C(_abc_42016_n2706_1), .Y(_abc_42016_n2707) );
  AOI21X1 AOI21X1_193 ( .A(_abc_42016_n2512), .B(_abc_42016_n2711_1), .C(_abc_42016_n1851), .Y(_abc_42016_n2712) );
  AOI21X1 AOI21X1_194 ( .A(_abc_42016_n2724), .B(_abc_42016_n1438), .C(_abc_42016_n2722), .Y(_abc_42016_n2725) );
  AOI21X1 AOI21X1_195 ( .A(_abc_42016_n2726), .B(_abc_42016_n2537), .C(_abc_42016_n2714), .Y(_abc_42016_n2727) );
  AOI21X1 AOI21X1_196 ( .A(_abc_42016_n2744), .B(_abc_42016_n673), .C(_abc_42016_n2304), .Y(_abc_42016_n2745) );
  AOI21X1 AOI21X1_197 ( .A(_abc_42016_n2749), .B(raddrhold_0_), .C(_abc_42016_n2755), .Y(_abc_42016_n2756) );
  AOI21X1 AOI21X1_198 ( .A(_abc_42016_n2760), .B(_abc_42016_n675), .C(_abc_42016_n2757), .Y(_abc_42016_n2761) );
  AOI21X1 AOI21X1_199 ( .A(rdatahold2_1_), .B(_abc_42016_n2271_1), .C(_abc_42016_n2735), .Y(_abc_42016_n2782) );
  AOI21X1 AOI21X1_2 ( .A(_abc_42016_n624), .B(_abc_42016_n637), .C(_abc_42016_n639), .Y(_abc_42016_n640) );
  AOI21X1 AOI21X1_20 ( .A(rdatahold2_6_), .B(_abc_42016_n694), .C(_abc_42016_n946), .Y(_abc_42016_n947) );
  AOI21X1 AOI21X1_200 ( .A(_abc_42016_n2776), .B(_abc_42016_n675), .C(_abc_42016_n2783), .Y(_abc_42016_n2784) );
  AOI21X1 AOI21X1_201 ( .A(rdatahold2_2_), .B(_abc_42016_n2271_1), .C(_abc_42016_n2790), .Y(_abc_42016_n2791) );
  AOI21X1 AOI21X1_202 ( .A(_abc_42016_n2747_1), .B(_abc_42016_n2792), .C(_abc_42016_n2786), .Y(_abc_42016_n2793) );
  AOI21X1 AOI21X1_203 ( .A(_abc_42016_n2431), .B(_abc_42016_n2754), .C(_abc_42016_n1139), .Y(_abc_42016_n2809) );
  AOI21X1 AOI21X1_204 ( .A(_abc_42016_n1910), .B(_abc_42016_n2811_1), .C(_abc_42016_n2746), .Y(_abc_42016_n2812) );
  AOI21X1 AOI21X1_205 ( .A(_abc_42016_n2747_1), .B(_abc_42016_n2821), .C(_abc_42016_n2820), .Y(_abc_42016_n2822) );
  AOI21X1 AOI21X1_206 ( .A(_abc_42016_n2833_1), .B(_abc_42016_n675), .C(_abc_42016_n2832), .Y(_abc_42016_n2834_1) );
  AOI21X1 AOI21X1_207 ( .A(_abc_42016_n2431), .B(_abc_42016_n2754), .C(_abc_42016_n872), .Y(_abc_42016_n2837) );
  AOI21X1 AOI21X1_208 ( .A(rdatahold2_5_), .B(_abc_42016_n2271_1), .C(_abc_42016_n2849), .Y(_abc_42016_n2850) );
  AOI21X1 AOI21X1_209 ( .A(raddrhold_6_), .B(_abc_42016_n2847), .C(_abc_42016_n2733), .Y(_abc_42016_n2862) );
  AOI21X1 AOI21X1_21 ( .A(_abc_42016_n950), .B(_abc_42016_n949), .C(_abc_42016_n606), .Y(_abc_42016_n951) );
  AOI21X1 AOI21X1_210 ( .A(_abc_42016_n2866), .B(_abc_42016_n675), .C(_abc_42016_n2865), .Y(_abc_42016_n2867) );
  AOI21X1 AOI21X1_211 ( .A(_abc_42016_n2279), .B(_abc_42016_n959), .C(_abc_42016_n1837_1), .Y(_abc_42016_n2870) );
  AOI21X1 AOI21X1_212 ( .A(_abc_42016_n2872), .B(_abc_42016_n2424), .C(_abc_42016_n2873), .Y(_abc_42016_n2874) );
  AOI21X1 AOI21X1_213 ( .A(_abc_42016_n2871), .B(_abc_42016_n2874), .C(_abc_42016_n560), .Y(_abc_42016_n2875) );
  AOI21X1 AOI21X1_214 ( .A(_abc_42016_n2880), .B(_abc_42016_n2869), .C(_abc_42016_n2733), .Y(_abc_42016_n2883) );
  AOI21X1 AOI21X1_215 ( .A(_abc_42016_n2882), .B(_abc_42016_n2883), .C(_abc_42016_n2884), .Y(_abc_42016_n2885) );
  AOI21X1 AOI21X1_216 ( .A(rdatahold_0_), .B(_abc_42016_n2271_1), .C(_abc_42016_n2890), .Y(_abc_42016_n2891) );
  AOI21X1 AOI21X1_217 ( .A(_abc_42016_n2280), .B(_abc_42016_n2887), .C(_abc_42016_n1837_1), .Y(_abc_42016_n2894) );
  AOI21X1 AOI21X1_218 ( .A(_abc_42016_n2911), .B(_abc_42016_n547), .C(_abc_42016_n2915), .Y(_abc_42016_n2916) );
  AOI21X1 AOI21X1_219 ( .A(_abc_42016_n2921), .B(_abc_42016_n2925_1), .C(_abc_42016_n2926), .Y(_abc_42016_n2927) );
  AOI21X1 AOI21X1_22 ( .A(rdatahold2_7_), .B(_abc_42016_n694), .C(_abc_42016_n984), .Y(_abc_42016_n985) );
  AOI21X1 AOI21X1_220 ( .A(_abc_42016_n2929), .B(raddrhold_10_), .C(_abc_42016_n2930), .Y(_abc_42016_n2931) );
  AOI21X1 AOI21X1_221 ( .A(_abc_42016_n2912), .B(_abc_42016_n2920), .C(_abc_42016_n2733), .Y(_abc_42016_n2936) );
  AOI21X1 AOI21X1_222 ( .A(_abc_42016_n2935), .B(_abc_42016_n2936), .C(_abc_42016_n2937), .Y(_abc_42016_n2938) );
  AOI21X1 AOI21X1_223 ( .A(_abc_42016_n2942), .B(_abc_42016_n2280), .C(_abc_42016_n2943), .Y(_abc_42016_n2944) );
  AOI21X1 AOI21X1_224 ( .A(_abc_42016_n2949), .B(_abc_42016_n2947_1), .C(_abc_42016_n548), .Y(_abc_42016_n2950) );
  AOI21X1 AOI21X1_225 ( .A(_abc_42016_n1513), .B(_abc_42016_n2424), .C(_abc_42016_n2960), .Y(_abc_42016_n2961) );
  AOI21X1 AOI21X1_226 ( .A(raddrhold_12_), .B(_abc_42016_n2951), .C(_abc_42016_n2967), .Y(_abc_42016_n2968) );
  AOI21X1 AOI21X1_227 ( .A(_abc_42016_n1527), .B(_abc_42016_n2279), .C(_abc_42016_n2974), .Y(_abc_42016_n2975) );
  AOI21X1 AOI21X1_228 ( .A(_abc_42016_n2973), .B(_abc_42016_n2424), .C(_abc_42016_n2975), .Y(_abc_42016_n2976) );
  AOI21X1 AOI21X1_229 ( .A(_abc_42016_n2983), .B(_abc_42016_n2972), .C(_abc_42016_n2733), .Y(_abc_42016_n2986) );
  AOI21X1 AOI21X1_23 ( .A(_abc_42016_n696), .B(regfil_3__0_), .C(_abc_42016_n1041), .Y(_abc_42016_n1042) );
  AOI21X1 AOI21X1_230 ( .A(_abc_42016_n2985), .B(_abc_42016_n2986), .C(_abc_42016_n2987), .Y(_abc_42016_n2988) );
  AOI21X1 AOI21X1_231 ( .A(_abc_42016_n2279), .B(_abc_42016_n1554), .C(_abc_42016_n1837_1), .Y(_abc_42016_n2993) );
  AOI21X1 AOI21X1_232 ( .A(_abc_42016_n2985), .B(_abc_42016_n2990_1), .C(_abc_42016_n2733), .Y(_abc_42016_n3005) );
  AOI21X1 AOI21X1_233 ( .A(_abc_42016_n3004), .B(_abc_42016_n3005), .C(_abc_42016_n3006), .Y(_abc_42016_n3007) );
  AOI21X1 AOI21X1_234 ( .A(_abc_42016_n1801_1), .B(_abc_42016_n2279), .C(_abc_42016_n3011), .Y(_abc_42016_n3012) );
  AOI21X1 AOI21X1_235 ( .A(_abc_42016_n1593), .B(_abc_42016_n2309), .C(_abc_42016_n2737), .Y(_abc_42016_n3013) );
  AOI21X1 AOI21X1_236 ( .A(rdatahold_7_), .B(_abc_42016_n2271_1), .C(_abc_42016_n2735), .Y(_abc_42016_n3024) );
  AOI21X1 AOI21X1_237 ( .A(_abc_42016_n3022), .B(_abc_42016_n547), .C(_abc_42016_n3025), .Y(_abc_42016_n3026) );
  AOI21X1 AOI21X1_238 ( .A(_abc_42016_n2700), .B(_abc_42016_n2358), .C(_abc_42016_n3028), .Y(_abc_42016_n3032) );
  AOI21X1 AOI21X1_239 ( .A(_abc_42016_n2293), .B(_abc_42016_n2300), .C(_abc_42016_n3028), .Y(_abc_42016_n3036_1) );
  AOI21X1 AOI21X1_24 ( .A(_abc_42016_n1044), .B(_abc_42016_n993), .C(_abc_42016_n1051), .Y(_abc_42016_n1052) );
  AOI21X1 AOI21X1_240 ( .A(_abc_42016_n3040), .B(_abc_42016_n3039), .C(_abc_42016_n1851), .Y(_abc_42016_n3041) );
  AOI21X1 AOI21X1_241 ( .A(_abc_42016_n3028), .B(_abc_42016_n1851), .C(_abc_42016_n548), .Y(_abc_42016_n3043) );
  AOI21X1 AOI21X1_242 ( .A(_abc_42016_n1399), .B(_abc_42016_n3052), .C(_abc_42016_n1373), .Y(_abc_42016_n3053) );
  AOI21X1 AOI21X1_243 ( .A(_abc_42016_n3050), .B(_abc_42016_n2280), .C(_abc_42016_n3060), .Y(_abc_42016_n3061) );
  AOI21X1 AOI21X1_244 ( .A(_abc_42016_n3050), .B(_abc_42016_n1851), .C(_abc_42016_n548), .Y(_abc_42016_n3068) );
  AOI21X1 AOI21X1_245 ( .A(_abc_42016_n3078_1), .B(_abc_42016_n1851), .C(_abc_42016_n548), .Y(_abc_42016_n3081) );
  AOI21X1 AOI21X1_246 ( .A(_abc_42016_n3092), .B(_abc_42016_n559), .C(_abc_42016_n3095), .Y(_abc_42016_n3096) );
  AOI21X1 AOI21X1_247 ( .A(_abc_42016_n3102), .B(_abc_42016_n3081), .C(_abc_42016_n3086), .Y(_abc_42016_n3103) );
  AOI21X1 AOI21X1_248 ( .A(_abc_42016_n3105_1), .B(_abc_42016_n1851), .C(_abc_42016_n548), .Y(_abc_42016_n3106_1) );
  AOI21X1 AOI21X1_249 ( .A(_abc_42016_n3125_1), .B(_abc_42016_n3106_1), .C(_abc_42016_n3110), .Y(_abc_42016_n3126_1) );
  AOI21X1 AOI21X1_25 ( .A(_abc_42016_n1025), .B(_abc_42016_n1072), .C(_abc_42016_n1022), .Y(_abc_42016_n1073_1) );
  AOI21X1 AOI21X1_250 ( .A(_abc_42016_n2359), .B(waddrhold_4_), .C(_abc_42016_n1851), .Y(_abc_42016_n3141) );
  AOI21X1 AOI21X1_251 ( .A(_abc_42016_n3140), .B(_abc_42016_n559), .C(_abc_42016_n3142), .Y(_abc_42016_n3143) );
  AOI21X1 AOI21X1_252 ( .A(_abc_42016_n3136), .B(_abc_42016_n3143), .C(_abc_42016_n3144), .Y(_abc_42016_n3145) );
  AOI21X1 AOI21X1_253 ( .A(_abc_42016_n3153), .B(_abc_42016_n2280), .C(_abc_42016_n2838), .Y(_abc_42016_n3154) );
  AOI21X1 AOI21X1_254 ( .A(_abc_42016_n3120), .B(_abc_42016_n1210), .C(_abc_42016_n1279), .Y(_abc_42016_n3162) );
  AOI21X1 AOI21X1_255 ( .A(_abc_42016_n3161), .B(_abc_42016_n3167), .C(_abc_42016_n2701), .Y(_abc_42016_n3168) );
  AOI21X1 AOI21X1_256 ( .A(_abc_42016_n3090), .B(waddrhold_6_), .C(_abc_42016_n3186), .Y(_abc_42016_n3187) );
  AOI21X1 AOI21X1_257 ( .A(_abc_42016_n2359), .B(waddrhold_6_), .C(_abc_42016_n1851), .Y(_abc_42016_n3189) );
  AOI21X1 AOI21X1_258 ( .A(_abc_42016_n3188), .B(_abc_42016_n559), .C(_abc_42016_n3190), .Y(_abc_42016_n3191) );
  AOI21X1 AOI21X1_259 ( .A(_abc_42016_n3184), .B(_abc_42016_n3191), .C(_abc_42016_n3192), .Y(_abc_42016_n3193) );
  AOI21X1 AOI21X1_26 ( .A(_abc_42016_n1078), .B(_abc_42016_n1081), .C(_abc_42016_n1082), .Y(_abc_42016_n1083) );
  AOI21X1 AOI21X1_260 ( .A(_abc_42016_n3205), .B(_abc_42016_n3204), .C(_abc_42016_n674), .Y(_abc_42016_n3206) );
  AOI21X1 AOI21X1_261 ( .A(_abc_42016_n959), .B(_abc_42016_n2279), .C(_abc_42016_n1848), .Y(_abc_42016_n3208) );
  AOI21X1 AOI21X1_262 ( .A(_abc_42016_n3201), .B(_abc_42016_n1851), .C(_abc_42016_n548), .Y(_abc_42016_n3214) );
  AOI21X1 AOI21X1_263 ( .A(_abc_42016_n3194), .B(_abc_42016_n3201), .C(_abc_42016_n2497), .Y(_abc_42016_n3218_1) );
  AOI21X1 AOI21X1_264 ( .A(regfil_5__7_), .B(_abc_42016_n2518_1), .C(_abc_42016_n3031), .Y(_abc_42016_n3219) );
  AOI21X1 AOI21X1_265 ( .A(_abc_42016_n3217_1), .B(_abc_42016_n3218_1), .C(_abc_42016_n3220), .Y(_abc_42016_n3221) );
  AOI21X1 AOI21X1_266 ( .A(_abc_42016_n3227), .B(_abc_42016_n3228), .C(_abc_42016_n674), .Y(_abc_42016_n3229) );
  AOI21X1 AOI21X1_267 ( .A(_abc_42016_n3223), .B(_abc_42016_n1851), .C(_abc_42016_n548), .Y(_abc_42016_n3236) );
  AOI21X1 AOI21X1_268 ( .A(_abc_42016_n3217_1), .B(_abc_42016_n3223), .C(_abc_42016_n2497), .Y(_abc_42016_n3240) );
  AOI21X1 AOI21X1_269 ( .A(_abc_42016_n3239), .B(_abc_42016_n3240), .C(_abc_42016_n3242), .Y(_abc_42016_n3243) );
  AOI21X1 AOI21X1_27 ( .A(_abc_42016_n1071), .B(_abc_42016_n1073_1), .C(_abc_42016_n1085), .Y(_abc_42016_n1086) );
  AOI21X1 AOI21X1_270 ( .A(_abc_42016_n3245_1), .B(_abc_42016_n1851), .C(_abc_42016_n548), .Y(_abc_42016_n3246) );
  AOI21X1 AOI21X1_271 ( .A(waddrhold_9_), .B(_abc_42016_n1410_1), .C(_abc_42016_n3250), .Y(_abc_42016_n3251) );
  AOI21X1 AOI21X1_272 ( .A(_abc_42016_n3245_1), .B(_abc_42016_n2280), .C(_abc_42016_n2903), .Y(_abc_42016_n3252) );
  AOI21X1 AOI21X1_273 ( .A(_abc_42016_n1841), .B(_abc_42016_n3245_1), .C(_abc_42016_n2355), .Y(_abc_42016_n3257) );
  AOI21X1 AOI21X1_274 ( .A(regfil_4__1_), .B(_abc_42016_n2518_1), .C(_abc_42016_n3031), .Y(_abc_42016_n3262) );
  AOI21X1 AOI21X1_275 ( .A(_abc_42016_n3239), .B(_abc_42016_n3245_1), .C(_abc_42016_n2497), .Y(_abc_42016_n3265) );
  AOI21X1 AOI21X1_276 ( .A(_abc_42016_n3265), .B(_abc_42016_n3264), .C(_abc_42016_n3263), .Y(_abc_42016_n3266_1) );
  AOI21X1 AOI21X1_277 ( .A(_abc_42016_n3268), .B(_abc_42016_n1851), .C(_abc_42016_n548), .Y(_abc_42016_n3282) );
  AOI21X1 AOI21X1_278 ( .A(regfil_4__2_), .B(_abc_42016_n2518_1), .C(_abc_42016_n3031), .Y(_abc_42016_n3287) );
  AOI21X1 AOI21X1_279 ( .A(_abc_42016_n3286), .B(_abc_42016_n3284), .C(_abc_42016_n3288), .Y(_abc_42016_n3289) );
  AOI21X1 AOI21X1_28 ( .A(_abc_42016_n1086), .B(_abc_42016_n1067), .C(_abc_42016_n1087), .Y(_abc_42016_n1088) );
  AOI21X1 AOI21X1_280 ( .A(_abc_42016_n3300), .B(_abc_42016_n673), .C(_abc_42016_n3306), .Y(_abc_42016_n3307) );
  AOI21X1 AOI21X1_281 ( .A(_abc_42016_n3307), .B(_abc_42016_n1863), .C(_abc_42016_n548), .Y(_abc_42016_n3308) );
  AOI21X1 AOI21X1_282 ( .A(_abc_42016_n3308), .B(_abc_42016_n3292), .C(_abc_42016_n3313), .Y(_abc_42016_n3314) );
  AOI21X1 AOI21X1_283 ( .A(_abc_42016_n3309), .B(_abc_42016_n3316), .C(_abc_42016_n2497), .Y(_abc_42016_n3317) );
  AOI21X1 AOI21X1_284 ( .A(_abc_42016_n3328), .B(_abc_42016_n559), .C(_abc_42016_n3329), .Y(_abc_42016_n3330) );
  AOI21X1 AOI21X1_285 ( .A(_abc_42016_n3316), .B(_abc_42016_n1851), .C(_abc_42016_n548), .Y(_abc_42016_n3332) );
  AOI21X1 AOI21X1_286 ( .A(rdatahold_4_), .B(_abc_42016_n3045), .C(_abc_42016_n3031), .Y(_abc_42016_n3333) );
  AOI21X1 AOI21X1_287 ( .A(_abc_42016_n3331), .B(_abc_42016_n3332), .C(_abc_42016_n3334), .Y(_abc_42016_n3335) );
  AOI21X1 AOI21X1_288 ( .A(_abc_42016_n1346), .B(_abc_42016_n1536), .C(_abc_42016_n3347), .Y(_abc_42016_n3348) );
  AOI21X1 AOI21X1_289 ( .A(waddrhold_13_), .B(_abc_42016_n2359), .C(_abc_42016_n3349), .Y(_abc_42016_n3350) );
  AOI21X1 AOI21X1_29 ( .A(rdatahold2_1_), .B(_abc_42016_n1057), .C(_abc_42016_n1090), .Y(_abc_42016_n1091) );
  AOI21X1 AOI21X1_290 ( .A(_abc_42016_n3337), .B(_abc_42016_n1851), .C(_abc_42016_n548), .Y(_abc_42016_n3352) );
  AOI21X1 AOI21X1_291 ( .A(waddrhold_13_), .B(_abc_42016_n3354), .C(_abc_42016_n3355), .Y(_abc_42016_n3356) );
  AOI21X1 AOI21X1_292 ( .A(regfil_4__5_), .B(_abc_42016_n2518_1), .C(_abc_42016_n3031), .Y(_abc_42016_n3357) );
  AOI21X1 AOI21X1_293 ( .A(waddrhold_14_), .B(_abc_42016_n2359), .C(_abc_42016_n3375), .Y(_abc_42016_n3376) );
  AOI21X1 AOI21X1_294 ( .A(_abc_42016_n3361), .B(_abc_42016_n1851), .C(_abc_42016_n548), .Y(_abc_42016_n3378) );
  AOI21X1 AOI21X1_295 ( .A(_abc_42016_n3380), .B(_abc_42016_n3361), .C(_abc_42016_n2497), .Y(_abc_42016_n3383) );
  AOI21X1 AOI21X1_296 ( .A(regfil_4__6_), .B(_abc_42016_n2518_1), .C(_abc_42016_n3031), .Y(_abc_42016_n3384) );
  AOI21X1 AOI21X1_297 ( .A(_abc_42016_n3382), .B(_abc_42016_n3383), .C(_abc_42016_n3385), .Y(_abc_42016_n3386) );
  AOI21X1 AOI21X1_298 ( .A(_abc_42016_n3390), .B(_abc_42016_n3391), .C(_abc_42016_n674), .Y(_abc_42016_n3392) );
  AOI21X1 AOI21X1_299 ( .A(_abc_42016_n3388), .B(_abc_42016_n1851), .C(_abc_42016_n548), .Y(_abc_42016_n3400) );
  AOI21X1 AOI21X1_3 ( .A(rdatahold2_0_), .B(_abc_42016_n694), .C(_abc_42016_n698), .Y(_abc_42016_n699) );
  AOI21X1 AOI21X1_30 ( .A(_abc_42016_n769), .B(_abc_42016_n989), .C(_abc_42016_n1055), .Y(_abc_42016_n1095) );
  AOI21X1 AOI21X1_300 ( .A(rdatahold_7_), .B(_abc_42016_n3045), .C(_abc_42016_n3031), .Y(_abc_42016_n3402) );
  AOI21X1 AOI21X1_301 ( .A(_abc_42016_n3404), .B(_abc_42016_n2519), .C(_abc_42016_n3403), .Y(_abc_42016_n3405) );
  AOI21X1 AOI21X1_302 ( .A(_abc_42016_n3433), .B(_abc_42016_n566), .C(_abc_42016_n560), .Y(_abc_42016_n3434) );
  AOI21X1 AOI21X1_303 ( .A(_abc_42016_n531), .B(_abc_42016_n3433), .C(_abc_42016_n3440), .Y(_abc_42016_n3441) );
  AOI21X1 AOI21X1_304 ( .A(_abc_42016_n530), .B(_abc_42016_n3433), .C(_abc_42016_n3446), .Y(_abc_42016_n3447_1) );
  AOI21X1 AOI21X1_305 ( .A(_abc_42016_n530), .B(_abc_42016_n1841), .C(_abc_42016_n3448_1), .Y(_abc_42016_n3449) );
  AOI21X1 AOI21X1_306 ( .A(_abc_42016_n2775), .B(_abc_42016_n2306), .C(_abc_42016_n3471), .Y(_abc_42016_n3472) );
  AOI21X1 AOI21X1_307 ( .A(sp_1_), .B(_abc_42016_n3453), .C(_abc_42016_n3478), .Y(_abc_42016_n3479_1) );
  AOI21X1 AOI21X1_308 ( .A(_abc_42016_n2775), .B(_abc_42016_n1344), .C(_abc_42016_n548), .Y(_abc_42016_n3481) );
  AOI21X1 AOI21X1_309 ( .A(_abc_42016_n1005), .B(regfil_5__2_), .C(_abc_42016_n674), .Y(_abc_42016_n3488_1) );
  AOI21X1 AOI21X1_31 ( .A(_abc_42016_n1005), .B(_abc_42016_n1118), .C(_abc_42016_n996), .Y(_abc_42016_n1119) );
  AOI21X1 AOI21X1_310 ( .A(sp_0_), .B(_abc_42016_n3098), .C(_abc_42016_n3475), .Y(_abc_42016_n3495) );
  AOI21X1 AOI21X1_311 ( .A(_abc_42016_n3495), .B(_abc_42016_n3494_1), .C(_abc_42016_n560), .Y(_abc_42016_n3496) );
  AOI21X1 AOI21X1_312 ( .A(_abc_42016_n3496), .B(_abc_42016_n3493), .C(_abc_42016_n3498), .Y(_abc_42016_n3499) );
  AOI21X1 AOI21X1_313 ( .A(_abc_42016_n3099), .B(_abc_42016_n3502), .C(_abc_42016_n3504), .Y(_abc_42016_n3505) );
  AOI21X1 AOI21X1_314 ( .A(_abc_42016_n3097), .B(_abc_42016_n2758), .C(_abc_42016_n2813), .Y(_abc_42016_n3515) );
  AOI21X1 AOI21X1_315 ( .A(_abc_42016_n3453), .B(sp_3_), .C(_abc_42016_n560), .Y(_abc_42016_n3522) );
  AOI21X1 AOI21X1_316 ( .A(_abc_42016_n3523), .B(_abc_42016_n3516), .C(_abc_42016_n3524), .Y(_abc_42016_n3525) );
  AOI21X1 AOI21X1_317 ( .A(_abc_42016_n2347_1), .B(_abc_42016_n3535), .C(_abc_42016_n3536), .Y(_abc_42016_n3537) );
  AOI21X1 AOI21X1_318 ( .A(_abc_42016_n3546), .B(_abc_42016_n3544), .C(_abc_42016_n560), .Y(_abc_42016_n3547) );
  AOI21X1 AOI21X1_319 ( .A(_abc_42016_n3547), .B(_abc_42016_n3543), .C(_abc_42016_n548), .Y(_abc_42016_n3548) );
  AOI21X1 AOI21X1_32 ( .A(_abc_42016_n1113_1), .B(_abc_42016_n1119), .C(_abc_42016_n1123), .Y(_abc_42016_n1124) );
  AOI21X1 AOI21X1_320 ( .A(_abc_42016_n3133), .B(_abc_42016_n3527), .C(_abc_42016_n3551), .Y(_abc_42016_n3552_1) );
  AOI21X1 AOI21X1_321 ( .A(_abc_42016_n3519), .B(sp_4_), .C(sp_5_), .Y(_abc_42016_n3564) );
  AOI21X1 AOI21X1_322 ( .A(_abc_42016_n3566), .B(_abc_42016_n1279), .C(_abc_42016_n560), .Y(_abc_42016_n3567_1) );
  AOI21X1 AOI21X1_323 ( .A(_abc_42016_n3572), .B(_abc_42016_n1279), .C(_abc_42016_n548), .Y(_abc_42016_n3573) );
  AOI21X1 AOI21X1_324 ( .A(_abc_42016_n3595), .B(_abc_42016_n3593), .C(_abc_42016_n3596), .Y(_abc_42016_n3597) );
  AOI21X1 AOI21X1_325 ( .A(_abc_42016_n3597), .B(_abc_42016_n3592), .C(_abc_42016_n548), .Y(_abc_42016_n3598) );
  AOI21X1 AOI21X1_326 ( .A(rdatahold2_6_), .B(_abc_42016_n3459), .C(_abc_42016_n3462), .Y(_abc_42016_n3601) );
  AOI21X1 AOI21X1_327 ( .A(_abc_42016_n3609), .B(_abc_42016_n3502), .C(_abc_42016_n3462), .Y(_abc_42016_n3610) );
  AOI21X1 AOI21X1_328 ( .A(rdatahold2_7_), .B(_abc_42016_n3459), .C(_abc_42016_n3611), .Y(_abc_42016_n3612) );
  AOI21X1 AOI21X1_329 ( .A(_abc_42016_n3594), .B(sp_7_), .C(_abc_42016_n3475), .Y(_abc_42016_n3616) );
  AOI21X1 AOI21X1_33 ( .A(_abc_42016_n696), .B(regfil_3__2_), .C(_abc_42016_n1131), .Y(_abc_42016_n1132) );
  AOI21X1 AOI21X1_330 ( .A(_abc_42016_n3617), .B(_abc_42016_n3615), .C(_abc_42016_n560), .Y(_abc_42016_n3618) );
  AOI21X1 AOI21X1_331 ( .A(_abc_42016_n3627), .B(_abc_42016_n3490), .C(_abc_42016_n560), .Y(_abc_42016_n3628_1) );
  AOI21X1 AOI21X1_332 ( .A(_abc_42016_n3572), .B(_abc_42016_n2131_1), .C(_abc_42016_n548), .Y(_abc_42016_n3643) );
  AOI21X1 AOI21X1_333 ( .A(rdatahold_0_), .B(_abc_42016_n3459), .C(_abc_42016_n3462), .Y(_abc_42016_n3645) );
  AOI21X1 AOI21X1_334 ( .A(_abc_42016_n3644), .B(_abc_42016_n3636), .C(_abc_42016_n3646), .Y(_abc_42016_n3647) );
  AOI21X1 AOI21X1_335 ( .A(_abc_42016_n3630), .B(_abc_42016_n2127_1), .C(_abc_42016_n3475), .Y(_abc_42016_n3654) );
  AOI21X1 AOI21X1_336 ( .A(_abc_42016_n3655), .B(_abc_42016_n3651), .C(_abc_42016_n560), .Y(_abc_42016_n3656) );
  AOI21X1 AOI21X1_337 ( .A(rdatahold_1_), .B(_abc_42016_n3459), .C(_abc_42016_n3462), .Y(_abc_42016_n3665) );
  AOI21X1 AOI21X1_338 ( .A(_abc_42016_n3502), .B(_abc_42016_n3658), .C(_abc_42016_n3666), .Y(_abc_42016_n3667) );
  AOI21X1 AOI21X1_339 ( .A(_abc_42016_n3652), .B(sp_0_), .C(sp_10_), .Y(_abc_42016_n3674) );
  AOI21X1 AOI21X1_34 ( .A(_abc_42016_n819), .B(_abc_42016_n989), .C(_abc_42016_n1055), .Y(_abc_42016_n1137) );
  AOI21X1 AOI21X1_340 ( .A(_abc_42016_n3490), .B(_abc_42016_n3671), .C(_abc_42016_n3675), .Y(_abc_42016_n3676) );
  AOI21X1 AOI21X1_341 ( .A(regfil_4__2_), .B(_abc_42016_n1005), .C(_abc_42016_n3554), .Y(_abc_42016_n3681) );
  AOI21X1 AOI21X1_342 ( .A(_abc_42016_n3679), .B(_abc_42016_n3502), .C(_abc_42016_n3687), .Y(_abc_42016_n3688) );
  AOI21X1 AOI21X1_343 ( .A(_abc_42016_n1005), .B(regfil_4__3_), .C(_abc_42016_n674), .Y(_abc_42016_n3690_1) );
  AOI21X1 AOI21X1_344 ( .A(_abc_42016_n3703), .B(_abc_42016_n3701), .C(_abc_42016_n560), .Y(_abc_42016_n3704) );
  AOI21X1 AOI21X1_345 ( .A(_abc_42016_n3704), .B(_abc_42016_n3700), .C(_abc_42016_n3705), .Y(_abc_42016_n3706) );
  AOI21X1 AOI21X1_346 ( .A(_abc_42016_n3297), .B(_abc_42016_n3527), .C(_abc_42016_n3709), .Y(_abc_42016_n3710) );
  AOI21X1 AOI21X1_347 ( .A(_abc_42016_n3714), .B(_abc_42016_n3715), .C(_abc_42016_n2256), .Y(_abc_42016_n3716) );
  AOI21X1 AOI21X1_348 ( .A(_abc_42016_n3730), .B(_abc_42016_n3721), .C(_abc_42016_n548), .Y(_abc_42016_n3731) );
  AOI21X1 AOI21X1_349 ( .A(_abc_42016_n3341), .B(_abc_42016_n1407), .C(_abc_42016_n3554), .Y(_abc_42016_n3749) );
  AOI21X1 AOI21X1_35 ( .A(_abc_42016_n1100), .B(_abc_42016_n1147_1), .C(_abc_42016_n1101_1), .Y(_abc_42016_n1148) );
  AOI21X1 AOI21X1_350 ( .A(_abc_42016_n3572), .B(_abc_42016_n2109_1), .C(_abc_42016_n548), .Y(_abc_42016_n3751) );
  AOI21X1 AOI21X1_351 ( .A(_abc_42016_n3365), .B(_abc_42016_n1407), .C(_abc_42016_n3770), .Y(_abc_42016_n3771) );
  AOI21X1 AOI21X1_352 ( .A(_abc_42016_n3572), .B(_abc_42016_n2103), .C(_abc_42016_n548), .Y(_abc_42016_n3773) );
  AOI21X1 AOI21X1_353 ( .A(_abc_42016_n3469), .B(sp_15_), .C(_abc_42016_n3787), .Y(_abc_42016_n3788) );
  AOI21X1 AOI21X1_354 ( .A(_abc_42016_n3790), .B(_abc_42016_n3788), .C(_abc_42016_n3791), .Y(_abc_42016_n3792) );
  AOI21X1 AOI21X1_355 ( .A(rdatahold_7_), .B(_abc_42016_n3459), .C(_abc_42016_n3462), .Y(_abc_42016_n3795) );
  AOI21X1 AOI21X1_356 ( .A(_abc_42016_n3502), .B(_abc_42016_n3789), .C(_abc_42016_n3796), .Y(_abc_42016_n3797_1) );
  AOI21X1 AOI21X1_357 ( .A(_abc_42016_n3800), .B(_abc_42016_n664_1), .C(_abc_42016_n1055), .Y(_abc_42016_n3801) );
  AOI21X1 AOI21X1_358 ( .A(regfil_5__7_), .B(_abc_42016_n1047_1), .C(_abc_42016_n3824), .Y(_abc_42016_n3825) );
  AOI21X1 AOI21X1_359 ( .A(_abc_42016_n1138), .B(_abc_42016_n3812), .C(_abc_42016_n3826), .Y(_abc_42016_n3827) );
  AOI21X1 AOI21X1_36 ( .A(_abc_42016_n1148), .B(_abc_42016_n1149_1), .C(_abc_42016_n1030), .Y(_abc_42016_n1150) );
  AOI21X1 AOI21X1_360 ( .A(_abc_42016_n3827), .B(_abc_42016_n1170), .C(_abc_42016_n3809), .Y(_abc_42016_n3828) );
  AOI21X1 AOI21X1_361 ( .A(_abc_42016_n602), .B(_abc_42016_n993), .C(_abc_42016_n1011), .Y(_abc_42016_n3829) );
  AOI21X1 AOI21X1_362 ( .A(rdatahold_0_), .B(_abc_42016_n1019), .C(_abc_42016_n1020), .Y(_abc_42016_n3831) );
  AOI21X1 AOI21X1_363 ( .A(_abc_42016_n3834), .B(regfil_4__1_), .C(_abc_42016_n1055), .Y(_abc_42016_n3835) );
  AOI21X1 AOI21X1_364 ( .A(_abc_42016_n1337_1), .B(regfil_4__0_), .C(regfil_4__1_), .Y(_abc_42016_n3837) );
  AOI21X1 AOI21X1_365 ( .A(_abc_42016_n3849), .B(_abc_42016_n3850), .C(_abc_42016_n1030), .Y(_abc_42016_n3851) );
  AOI21X1 AOI21X1_366 ( .A(_abc_42016_n3855), .B(_abc_42016_n3840), .C(_abc_42016_n3858), .Y(_abc_42016_n3859_1) );
  AOI21X1 AOI21X1_367 ( .A(_abc_42016_n3834), .B(_abc_42016_n1446), .C(_abc_42016_n1055), .Y(_abc_42016_n3864) );
  AOI21X1 AOI21X1_368 ( .A(_abc_42016_n2204), .B(_abc_42016_n2194), .C(_abc_42016_n2193), .Y(_abc_42016_n3879) );
  AOI21X1 AOI21X1_369 ( .A(_abc_42016_n1023), .B(_abc_42016_n3877), .C(_abc_42016_n3886), .Y(_abc_42016_n3887) );
  AOI21X1 AOI21X1_37 ( .A(_abc_42016_n1146_1), .B(_abc_42016_n1150), .C(_abc_42016_n1157), .Y(_abc_42016_n1158) );
  AOI21X1 AOI21X1_370 ( .A(_abc_42016_n3891), .B(regfil_2__2_), .C(_abc_42016_n993), .Y(_abc_42016_n3892) );
  AOI21X1 AOI21X1_371 ( .A(rdatahold_2_), .B(_abc_42016_n1019), .C(_abc_42016_n3893), .Y(_abc_42016_n3894) );
  AOI21X1 AOI21X1_372 ( .A(_abc_42016_n3902), .B(_abc_42016_n3903), .C(_abc_42016_n1151), .Y(_abc_42016_n3904) );
  AOI21X1 AOI21X1_373 ( .A(_abc_42016_n3838), .B(regfil_4__2_), .C(regfil_4__3_), .Y(_abc_42016_n3908) );
  AOI21X1 AOI21X1_374 ( .A(_abc_42016_n1225), .B(_abc_42016_n3909), .C(_abc_42016_n3918), .Y(_abc_42016_n3919) );
  AOI21X1 AOI21X1_375 ( .A(_abc_42016_n3920), .B(_abc_42016_n3900), .C(_abc_42016_n3921), .Y(_abc_42016_n3922) );
  AOI21X1 AOI21X1_376 ( .A(_abc_42016_n3834), .B(_abc_42016_n842), .C(_abc_42016_n1055), .Y(_abc_42016_n3926) );
  AOI21X1 AOI21X1_377 ( .A(_abc_42016_n3932), .B(_abc_42016_n3931), .C(_abc_42016_n3937), .Y(_abc_42016_n3938) );
  AOI21X1 AOI21X1_378 ( .A(_abc_42016_n3949), .B(_abc_42016_n3946), .C(_abc_42016_n1293), .Y(_abc_42016_n3950) );
  AOI21X1 AOI21X1_379 ( .A(rdatahold_4_), .B(_abc_42016_n1019), .C(_abc_42016_n993), .Y(_abc_42016_n3951) );
  AOI21X1 AOI21X1_38 ( .A(_abc_42016_n1162), .B(_abc_42016_n1163), .C(_abc_42016_n1160), .Y(_abc_42016_n1164) );
  AOI21X1 AOI21X1_380 ( .A(_abc_42016_n3945), .B(_abc_42016_n3950), .C(_abc_42016_n3952), .Y(_abc_42016_n3953) );
  AOI21X1 AOI21X1_381 ( .A(_abc_42016_n3834), .B(regfil_4__5_), .C(_abc_42016_n1055), .Y(_abc_42016_n3956) );
  AOI21X1 AOI21X1_382 ( .A(_abc_42016_n3965), .B(_abc_42016_n3966), .C(_abc_42016_n1151), .Y(_abc_42016_n3967) );
  AOI21X1 AOI21X1_383 ( .A(_abc_42016_n3973), .B(_abc_42016_n1023), .C(_abc_42016_n3804), .Y(_abc_42016_n3974) );
  AOI21X1 AOI21X1_384 ( .A(_abc_42016_n3978), .B(_abc_42016_n3976), .C(_abc_42016_n1125), .Y(_abc_42016_n3979) );
  AOI21X1 AOI21X1_385 ( .A(_abc_42016_n3975), .B(_abc_42016_n3979), .C(_abc_42016_n3960), .Y(_abc_42016_n3980) );
  AOI21X1 AOI21X1_386 ( .A(_abc_42016_n891), .B(_abc_42016_n993), .C(_abc_42016_n1011), .Y(_abc_42016_n3981) );
  AOI21X1 AOI21X1_387 ( .A(rdatahold_5_), .B(_abc_42016_n1019), .C(_abc_42016_n1020), .Y(_abc_42016_n3983_1) );
  AOI21X1 AOI21X1_388 ( .A(_abc_42016_n3834), .B(_abc_42016_n1554), .C(_abc_42016_n1055), .Y(_abc_42016_n3985) );
  AOI21X1 AOI21X1_389 ( .A(_abc_42016_n3958), .B(_abc_42016_n1554), .C(_abc_42016_n1170), .Y(_abc_42016_n3989) );
  AOI21X1 AOI21X1_39 ( .A(_abc_42016_n696), .B(regfil_3__3_), .C(_abc_42016_n993), .Y(_abc_42016_n1171_1) );
  AOI21X1 AOI21X1_390 ( .A(_abc_42016_n2141), .B(_abc_42016_n2108), .C(_abc_42016_n2106), .Y(_abc_42016_n3995) );
  AOI21X1 AOI21X1_391 ( .A(_abc_42016_n3933), .B(regfil_4__5_), .C(regfil_4__6_), .Y(_abc_42016_n4001) );
  AOI21X1 AOI21X1_392 ( .A(_abc_42016_n1023), .B(_abc_42016_n3996), .C(_abc_42016_n4004), .Y(_abc_42016_n4005) );
  AOI21X1 AOI21X1_393 ( .A(_abc_42016_n1793), .B(_abc_42016_n993), .C(_abc_42016_n1051), .Y(_abc_42016_n4008) );
  AOI21X1 AOI21X1_394 ( .A(_abc_42016_n3834), .B(_abc_42016_n1801_1), .C(_abc_42016_n1055), .Y(_abc_42016_n4011) );
  AOI21X1 AOI21X1_395 ( .A(_abc_42016_n4036), .B(_abc_42016_n4034), .C(_abc_42016_n1125), .Y(_abc_42016_n4037) );
  AOI21X1 AOI21X1_396 ( .A(_abc_42016_n4039), .B(regfil_4__7_), .C(_abc_42016_n1170), .Y(_abc_42016_n4040) );
  AOI21X1 AOI21X1_397 ( .A(_abc_42016_n2478), .B(_abc_42016_n1096), .C(_abc_42016_n4071), .Y(_abc_42016_n4072) );
  AOI21X1 AOI21X1_398 ( .A(_abc_42016_n1381), .B(_abc_42016_n4114), .C(_abc_42016_n4116), .Y(_abc_42016_n4117) );
  AOI21X1 AOI21X1_399 ( .A(_abc_42016_n4122), .B(_abc_42016_n4096), .C(reset), .Y(pc_0__FF_INPUT) );
  AOI21X1 AOI21X1_4 ( .A(_abc_42016_n705), .B(_abc_42016_n707_1), .C(_abc_42016_n684), .Y(_abc_42016_n708) );
  AOI21X1 AOI21X1_40 ( .A(_abc_42016_n1174_1), .B(_abc_42016_n993), .C(_abc_42016_n1011), .Y(_abc_42016_n1175) );
  AOI21X1 AOI21X1_400 ( .A(_abc_42016_n4124), .B(_abc_42016_n4125), .C(_abc_42016_n560), .Y(_abc_42016_n4126) );
  AOI21X1 AOI21X1_401 ( .A(_abc_42016_n4129), .B(_abc_42016_n559), .C(_abc_42016_n4127), .Y(_abc_42016_n4130) );
  AOI21X1 AOI21X1_402 ( .A(_abc_42016_n4087), .B(_abc_42016_n2526), .C(_abc_42016_n4133), .Y(_abc_42016_n4134) );
  AOI21X1 AOI21X1_403 ( .A(_abc_42016_n4138), .B(_abc_42016_n4139), .C(reset), .Y(pc_1__FF_INPUT) );
  AOI21X1 AOI21X1_404 ( .A(_abc_42016_n4141), .B(_abc_42016_n4143), .C(_abc_42016_n560), .Y(_abc_42016_n4144) );
  AOI21X1 AOI21X1_405 ( .A(_abc_42016_n4153), .B(_abc_42016_n4154), .C(reset), .Y(pc_2__FF_INPUT) );
  AOI21X1 AOI21X1_406 ( .A(_abc_42016_n4169), .B(_abc_42016_n4170), .C(reset), .Y(pc_3__FF_INPUT) );
  AOI21X1 AOI21X1_407 ( .A(_abc_42016_n4089), .B(_abc_42016_n4173), .C(_abc_42016_n4176), .Y(_abc_42016_n4177) );
  AOI21X1 AOI21X1_408 ( .A(_abc_42016_n4181), .B(_abc_42016_n4182), .C(reset), .Y(pc_4__FF_INPUT) );
  AOI21X1 AOI21X1_409 ( .A(_abc_42016_n4195), .B(_abc_42016_n4196), .C(reset), .Y(pc_5__FF_INPUT) );
  AOI21X1 AOI21X1_41 ( .A(rdatahold2_3_), .B(_abc_42016_n1019), .C(_abc_42016_n1020), .Y(_abc_42016_n1177) );
  AOI21X1 AOI21X1_410 ( .A(_abc_42016_n4207), .B(_abc_42016_n4208), .C(reset), .Y(pc_6__FF_INPUT) );
  AOI21X1 AOI21X1_411 ( .A(_abc_42016_n2724), .B(_abc_42016_n4077), .C(_abc_42016_n4215), .Y(_abc_42016_n4216) );
  AOI21X1 AOI21X1_412 ( .A(_abc_42016_n4210), .B(pc_7_), .C(_abc_42016_n4217), .Y(_abc_42016_n4218) );
  AOI21X1 AOI21X1_413 ( .A(_abc_42016_n4220), .B(_abc_42016_n4221), .C(reset), .Y(pc_7__FF_INPUT) );
  AOI21X1 AOI21X1_414 ( .A(_abc_42016_n4233), .B(_abc_42016_n4234), .C(reset), .Y(pc_8__FF_INPUT) );
  AOI21X1 AOI21X1_415 ( .A(_abc_42016_n4246), .B(_abc_42016_n4247), .C(reset), .Y(pc_9__FF_INPUT) );
  AOI21X1 AOI21X1_416 ( .A(_abc_42016_n4253), .B(_abc_42016_n4252), .C(_abc_42016_n4131), .Y(_abc_42016_n4254) );
  AOI21X1 AOI21X1_417 ( .A(_abc_42016_n4258), .B(_abc_42016_n4259), .C(reset), .Y(pc_10__FF_INPUT) );
  AOI21X1 AOI21X1_418 ( .A(_abc_42016_n4264), .B(_abc_42016_n4089), .C(_abc_42016_n3935_1), .Y(_abc_42016_n4265) );
  AOI21X1 AOI21X1_419 ( .A(_abc_42016_n4261), .B(_abc_42016_n4087), .C(_abc_42016_n4266_1), .Y(_abc_42016_n4267) );
  AOI21X1 AOI21X1_42 ( .A(_abc_42016_n1047_1), .B(regfil_5__3_), .C(_abc_42016_n1023), .Y(_abc_42016_n1207) );
  AOI21X1 AOI21X1_420 ( .A(_abc_42016_n4272), .B(_abc_42016_n4273), .C(reset), .Y(pc_11__FF_INPUT) );
  AOI21X1 AOI21X1_421 ( .A(_abc_42016_n1513), .B(_abc_42016_n4087), .C(_abc_42016_n4277), .Y(_abc_42016_n4278) );
  AOI21X1 AOI21X1_422 ( .A(_abc_42016_n4284), .B(_abc_42016_n4285), .C(reset), .Y(pc_12__FF_INPUT) );
  AOI21X1 AOI21X1_423 ( .A(_abc_42016_n4296), .B(_abc_42016_n4297), .C(reset), .Y(pc_13__FF_INPUT) );
  AOI21X1 AOI21X1_424 ( .A(_abc_42016_n4301), .B(_abc_42016_n4077), .C(_abc_42016_n4026), .Y(_abc_42016_n4302) );
  AOI21X1 AOI21X1_425 ( .A(_abc_42016_n2285), .B(_abc_42016_n4301), .C(_abc_42016_n4306), .Y(_abc_42016_n4307) );
  AOI21X1 AOI21X1_426 ( .A(_abc_42016_n4309), .B(_abc_42016_n4312), .C(reset), .Y(pc_14__FF_INPUT) );
  AOI21X1 AOI21X1_427 ( .A(_abc_42016_n4314), .B(_abc_42016_n4315), .C(_abc_42016_n4131), .Y(_abc_42016_n4316) );
  AOI21X1 AOI21X1_428 ( .A(_abc_42016_n4320_1), .B(_abc_42016_n4321), .C(reset), .Y(pc_15__FF_INPUT) );
  AOI21X1 AOI21X1_429 ( .A(_abc_42016_n4340), .B(_abc_42016_n663), .C(_abc_42016_n4071), .Y(_abc_42016_n4341) );
  AOI21X1 AOI21X1_43 ( .A(_abc_42016_n1023), .B(_abc_42016_n1216), .C(_abc_42016_n1009), .Y(_abc_42016_n1217) );
  AOI21X1 AOI21X1_430 ( .A(_abc_42016_n4065), .B(_abc_42016_n4351), .C(_abc_42016_n4353), .Y(_abc_42016_n4354) );
  AOI21X1 AOI21X1_431 ( .A(regfil_7__1_), .B(_abc_42016_n4056), .C(_abc_42016_n4360), .Y(_abc_42016_n4361) );
  AOI21X1 AOI21X1_432 ( .A(rdatahold_1_), .B(_abc_42016_n4362), .C(_abc_42016_n4364), .Y(_abc_42016_n4365) );
  AOI21X1 AOI21X1_433 ( .A(_abc_42016_n768), .B(_abc_42016_n4340), .C(_abc_42016_n4071), .Y(_abc_42016_n4372) );
  AOI21X1 AOI21X1_434 ( .A(regfil_7__2_), .B(_abc_42016_n4056), .C(_abc_42016_n4375), .Y(_abc_42016_n4376) );
  AOI21X1 AOI21X1_435 ( .A(regfil_7__1_), .B(_abc_42016_n4377), .C(_abc_42016_n4384), .Y(_abc_42016_n4385) );
  AOI21X1 AOI21X1_436 ( .A(_abc_42016_n4340), .B(_abc_42016_n818), .C(_abc_42016_n4071), .Y(_abc_42016_n4387) );
  AOI21X1 AOI21X1_437 ( .A(regfil_7__3_), .B(_abc_42016_n4056), .C(_abc_42016_n4390), .Y(_abc_42016_n4391) );
  AOI21X1 AOI21X1_438 ( .A(regfil_7__5_), .B(_abc_42016_n4381), .C(_abc_42016_n4407), .Y(_abc_42016_n4408) );
  AOI21X1 AOI21X1_439 ( .A(regfil_7__6_), .B(_abc_42016_n4381), .C(_abc_42016_n4417), .Y(_abc_42016_n4418) );
  AOI21X1 AOI21X1_44 ( .A(_abc_42016_n1208), .B(_abc_42016_n1217), .C(_abc_42016_n1191), .Y(_abc_42016_n1218) );
  AOI21X1 AOI21X1_440 ( .A(_abc_42016_n4428), .B(_abc_42016_n924), .C(_abc_42016_n4379), .Y(_abc_42016_n4429) );
  AOI21X1 AOI21X1_441 ( .A(_abc_42016_n4381), .B(regfil_7__7_), .C(_abc_42016_n4432), .Y(_abc_42016_n4433) );
  AOI21X1 AOI21X1_442 ( .A(\data[7] ), .B(_abc_42016_n4047), .C(_abc_42016_n4443), .Y(_abc_42016_n4444) );
  AOI21X1 AOI21X1_443 ( .A(alu_res_7_), .B(_abc_42016_n4057), .C(_abc_42016_n4369), .Y(_abc_42016_n4445) );
  AOI21X1 AOI21X1_444 ( .A(pc_0_), .B(_abc_42016_n2026), .C(_abc_42016_n4473), .Y(_abc_42016_n4474) );
  AOI21X1 AOI21X1_445 ( .A(raddrhold_9_), .B(_abc_42016_n2732), .C(_abc_42016_n4519), .Y(_abc_42016_n4520) );
  AOI21X1 AOI21X1_446 ( .A(_abc_42016_n4471), .B(_abc_42016_n4520), .C(_abc_42016_n4521), .Y(addr_9__FF_INPUT) );
  AOI21X1 AOI21X1_447 ( .A(raddrhold_10_), .B(_abc_42016_n2732), .C(_abc_42016_n4523), .Y(_abc_42016_n4524_1) );
  AOI21X1 AOI21X1_448 ( .A(_abc_42016_n4471), .B(_abc_42016_n4524_1), .C(_abc_42016_n4525), .Y(addr_10__FF_INPUT) );
  AOI21X1 AOI21X1_449 ( .A(raddrhold_11_), .B(_abc_42016_n2732), .C(_abc_42016_n4527), .Y(_abc_42016_n4528) );
  AOI21X1 AOI21X1_45 ( .A(_abc_42016_n1230), .B(_abc_42016_n1229), .C(_abc_42016_n1231), .Y(_abc_42016_n1233) );
  AOI21X1 AOI21X1_450 ( .A(_abc_42016_n4471), .B(_abc_42016_n4528), .C(_abc_42016_n4529), .Y(addr_11__FF_INPUT) );
  AOI21X1 AOI21X1_451 ( .A(raddrhold_12_), .B(_abc_42016_n2732), .C(_abc_42016_n4531), .Y(_abc_42016_n4532) );
  AOI21X1 AOI21X1_452 ( .A(_abc_42016_n4471), .B(_abc_42016_n4532), .C(_abc_42016_n4533), .Y(addr_12__FF_INPUT) );
  AOI21X1 AOI21X1_453 ( .A(raddrhold_14_), .B(_abc_42016_n2732), .C(_abc_42016_n4540), .Y(_abc_42016_n4541) );
  AOI21X1 AOI21X1_454 ( .A(_abc_42016_n4471), .B(_abc_42016_n4541), .C(_abc_42016_n4542), .Y(addr_14__FF_INPUT) );
  AOI21X1 AOI21X1_455 ( .A(pc_15_), .B(_abc_42016_n2026), .C(_abc_42016_n4544), .Y(_abc_42016_n4545) );
  AOI21X1 AOI21X1_456 ( .A(_abc_42016_n4471), .B(_abc_42016_n4545), .C(_abc_42016_n4546), .Y(addr_15__FF_INPUT) );
  AOI21X1 AOI21X1_457 ( .A(_abc_42016_n4570_1), .B(_abc_42016_n4594), .C(_abc_42016_n4598), .Y(_abc_42016_n4599) );
  AOI21X1 AOI21X1_458 ( .A(_abc_42016_n2226), .B(_abc_42016_n4459), .C(_abc_42016_n4605), .Y(_abc_42016_n4606) );
  AOI21X1 AOI21X1_459 ( .A(_abc_42016_n4549), .B(_abc_42016_n4553), .C(_abc_42016_n4609), .Y(_abc_42016_n4610) );
  AOI21X1 AOI21X1_46 ( .A(_abc_42016_n1197_1), .B(_abc_42016_n1193), .C(_abc_42016_n1236), .Y(_abc_42016_n1237) );
  AOI21X1 AOI21X1_460 ( .A(_abc_42016_n677), .B(_abc_42016_n4653), .C(_abc_42016_n4671), .Y(_abc_42016_n4672_1) );
  AOI21X1 AOI21X1_461 ( .A(_abc_42016_n4550), .B(_abc_42016_n4681), .C(_abc_42016_n4683), .Y(_abc_42016_n4684_1) );
  AOI21X1 AOI21X1_462 ( .A(_abc_42016_n4550), .B(_abc_42016_n4615_1), .C(_abc_42016_n4348), .Y(_abc_42016_n4730) );
  AOI21X1 AOI21X1_463 ( .A(_abc_42016_n2026), .B(_abc_42016_n4738), .C(reset), .Y(_abc_42016_n4739) );
  AOI21X1 AOI21X1_464 ( .A(alu__abc_41682_n41), .B(alu__abc_41682_n44), .C(alu__abc_41682_n54), .Y(alu__abc_41682_n55) );
  AOI21X1 AOI21X1_465 ( .A(alu__abc_41682_n68), .B(alu__abc_41682_n60), .C(alu__abc_41682_n76), .Y(alu__abc_41682_n83) );
  AOI21X1 AOI21X1_466 ( .A(alu__abc_41682_n89), .B(alu__abc_41682_n94), .C(alu__abc_41682_n99), .Y(alu__abc_41682_n100) );
  AOI21X1 AOI21X1_467 ( .A(alu__abc_41682_n89), .B(alu__abc_41682_n94), .C(alu__abc_41682_n108), .Y(alu__abc_41682_n111) );
  AOI21X1 AOI21X1_468 ( .A(alu__abc_41682_n126), .B(alu__abc_41682_n124_1), .C(alu__abc_41682_n41), .Y(alu__abc_41682_n127) );
  AOI21X1 AOI21X1_469 ( .A(alu__abc_41682_n142), .B(alu__abc_41682_n166), .C(alu__abc_41682_n165), .Y(alu__abc_41682_n167) );
  AOI21X1 AOI21X1_47 ( .A(_abc_42016_n1031_1), .B(_abc_42016_n1244), .C(_abc_42016_n1247_1), .Y(_abc_42016_n1248_1) );
  AOI21X1 AOI21X1_470 ( .A(alu__abc_41682_n144), .B(alu__abc_41682_n160), .C(alu__abc_41682_n171), .Y(alu__abc_41682_n172) );
  AOI21X1 AOI21X1_471 ( .A(alu__abc_41682_n146), .B(alu__abc_41682_n151), .C(alu__abc_41682_n189), .Y(alu__abc_41682_n190) );
  AOI21X1 AOI21X1_472 ( .A(alu__abc_41682_n177), .B(alu__abc_41682_n190), .C(alu__abc_41682_n187), .Y(alu__abc_41682_n191) );
  AOI21X1 AOI21X1_473 ( .A(alu__abc_41682_n92), .B(alu__abc_41682_n81), .C(alu__abc_41682_n198), .Y(alu__abc_41682_n199) );
  AOI21X1 AOI21X1_474 ( .A(alu__abc_41682_n143), .B(alu__abc_41682_n49), .C(alu__abc_41682_n135), .Y(alu__abc_41682_n201) );
  AOI21X1 AOI21X1_475 ( .A(alu__abc_41682_n203), .B(alu__abc_41682_n126), .C(alu__abc_41682_n161), .Y(alu__abc_41682_n204) );
  AOI21X1 AOI21X1_476 ( .A(alu__abc_41682_n207), .B(alu__abc_41682_n208), .C(alu__abc_41682_n206), .Y(alu__abc_41682_n209) );
  AOI21X1 AOI21X1_477 ( .A(alu__abc_41682_n130), .B(alu__abc_41682_n156), .C(alu__abc_41682_n216), .Y(alu__abc_41682_n217) );
  AOI21X1 AOI21X1_478 ( .A(alu__abc_41682_n214), .B(alu__abc_41682_n217), .C(alu__abc_41682_n221), .Y(alu__abc_41682_n222) );
  AOI21X1 AOI21X1_479 ( .A(alu__abc_41682_n235), .B(alu__abc_41682_n236), .C(alu__abc_41682_n234), .Y(alu__abc_41682_n237) );
  AOI21X1 AOI21X1_48 ( .A(_abc_42016_n1225), .B(_abc_42016_n1228), .C(_abc_42016_n1249), .Y(_abc_42016_n1250_1) );
  AOI21X1 AOI21X1_480 ( .A(alu__abc_41682_n229), .B(alu__abc_41682_n58), .C(alu__abc_41682_n198), .Y(alu__abc_41682_n239) );
  AOI21X1 AOI21X1_481 ( .A(alu__abc_41682_n62), .B(alu__abc_41682_n240), .C(alu__abc_41682_n242), .Y(alu__abc_41682_n243) );
  AOI21X1 AOI21X1_482 ( .A(alu__abc_41682_n239), .B(alu__abc_41682_n238), .C(alu__abc_41682_n244), .Y(alu__abc_41682_n245) );
  AOI21X1 AOI21X1_483 ( .A(alu__abc_41682_n257), .B(alu__abc_41682_n248), .C(alu__abc_41682_n246), .Y(alu__abc_41682_n258) );
  AOI21X1 AOI21X1_484 ( .A(alu__abc_41682_n168), .B(alu__abc_41682_n170), .C(alu__abc_41682_n154), .Y(alu__abc_41682_n266_1) );
  AOI21X1 AOI21X1_485 ( .A(alu__abc_41682_n58), .B(alu__abc_41682_n107), .C(alu__abc_41682_n194), .Y(alu__abc_41682_n269) );
  AOI21X1 AOI21X1_486 ( .A(alu__abc_41682_n279_1), .B(alu__abc_41682_n265), .C(alu__abc_41682_n280_1), .Y(alu__abc_41682_n281) );
  AOI21X1 AOI21X1_487 ( .A(alu__abc_41682_n285), .B(alu__abc_41682_n150), .C(alu__abc_41682_n282), .Y(alu__abc_41682_n286_1) );
  AOI21X1 AOI21X1_488 ( .A(alu__abc_41682_n291), .B(alu__abc_41682_n299), .C(alu__abc_41682_n198), .Y(alu__abc_41682_n300) );
  AOI21X1 AOI21X1_489 ( .A(alu__abc_41682_n193), .B(alu__abc_41682_n305), .C(alu__abc_41682_n310), .Y(alu__abc_41682_n311) );
  AOI21X1 AOI21X1_49 ( .A(_abc_42016_n933), .B(_abc_42016_n930), .C(_abc_42016_n990), .Y(_abc_42016_n1259) );
  AOI21X1 AOI21X1_490 ( .A(alu__abc_41682_n192), .B(alu__abc_41682_n195), .C(alu__abc_41682_n224), .Y(alu__abc_41682_n330) );
  AOI21X1 AOI21X1_491 ( .A(alu__abc_41682_n237), .B(alu__abc_41682_n107), .C(alu__abc_41682_n356), .Y(alu__abc_41682_n357) );
  AOI21X1 AOI21X1_492 ( .A(alu__abc_41682_n89), .B(alu__abc_41682_n94), .C(alu__abc_41682_n95), .Y(alu__abc_41682_n359) );
  AOI21X1 AOI21X1_493 ( .A(alu__abc_41682_n96), .B(alu_opra_7_), .C(alu__abc_41682_n362), .Y(alu__abc_41682_n363) );
  AOI21X1 AOI21X1_5 ( .A(_abc_42016_n712), .B(_abc_42016_n655_1), .C(_abc_42016_n713), .Y(_abc_42016_n714) );
  AOI21X1 AOI21X1_50 ( .A(_abc_42016_n1204), .B(_abc_42016_n1241), .C(_abc_42016_n1243), .Y(_abc_42016_n1271_1) );
  AOI21X1 AOI21X1_51 ( .A(_abc_42016_n1272_1), .B(_abc_42016_n1273), .C(_abc_42016_n1030), .Y(_abc_42016_n1274_1) );
  AOI21X1 AOI21X1_52 ( .A(_abc_42016_n1278), .B(_abc_42016_n1269), .C(_abc_42016_n1287), .Y(_abc_42016_n1288) );
  AOI21X1 AOI21X1_53 ( .A(_abc_42016_n1294), .B(_abc_42016_n1297_1), .C(_abc_42016_n1293), .Y(_abc_42016_n1298) );
  AOI21X1 AOI21X1_54 ( .A(regfil_3__6_), .B(_abc_42016_n696), .C(_abc_42016_n1058), .Y(_abc_42016_n1300) );
  AOI21X1 AOI21X1_55 ( .A(_abc_42016_n1299_1), .B(_abc_42016_n1300), .C(_abc_42016_n1263), .Y(_abc_36783_n3453) );
  AOI21X1 AOI21X1_56 ( .A(_abc_42016_n1266), .B(_abc_42016_n1305), .C(_abc_42016_n1308), .Y(_abc_42016_n1309) );
  AOI21X1 AOI21X1_57 ( .A(_abc_42016_n1319), .B(_abc_42016_n1031_1), .C(_abc_42016_n1321_1), .Y(_abc_42016_n1322) );
  AOI21X1 AOI21X1_58 ( .A(_abc_42016_n1324), .B(_abc_42016_n1330), .C(_abc_42016_n1045), .Y(_abc_42016_n1332) );
  AOI21X1 AOI21X1_59 ( .A(_abc_42016_n1290), .B(_abc_42016_n959), .C(_abc_42016_n1187), .Y(_abc_42016_n1339_1) );
  AOI21X1 AOI21X1_6 ( .A(_abc_42016_n716), .B(_abc_42016_n717), .C(_abc_42016_n606), .Y(_abc_42016_n718) );
  AOI21X1 AOI21X1_60 ( .A(opcode_4_), .B(regfil_2__0_), .C(_abc_42016_n1394), .Y(_abc_42016_n1395) );
  AOI21X1 AOI21X1_61 ( .A(_abc_42016_n1370), .B(_abc_42016_n1379), .C(_abc_42016_n1415), .Y(_abc_42016_n1416) );
  AOI21X1 AOI21X1_62 ( .A(regfil_4__1_), .B(_abc_42016_n1426), .C(_abc_42016_n1431), .Y(_abc_42016_n1432) );
  AOI21X1 AOI21X1_63 ( .A(pc_9_), .B(_abc_42016_n1437), .C(_abc_42016_n1438), .Y(_abc_42016_n1439_1) );
  AOI21X1 AOI21X1_64 ( .A(_abc_42016_n1410_1), .B(_abc_42016_n1419), .C(_abc_42016_n674), .Y(_abc_42016_n1442) );
  AOI21X1 AOI21X1_65 ( .A(pc_10_), .B(_abc_42016_n1437), .C(_abc_42016_n1438), .Y(_abc_42016_n1453) );
  AOI21X1 AOI21X1_66 ( .A(_abc_42016_n1464), .B(pc_0_), .C(pc_10_), .Y(_abc_42016_n1465_1) );
  AOI21X1 AOI21X1_67 ( .A(pc_0_), .B(_abc_42016_n1466), .C(_abc_42016_n1465_1), .Y(_abc_42016_n1467) );
  AOI21X1 AOI21X1_68 ( .A(_abc_42016_n1410_1), .B(_abc_42016_n1445), .C(_abc_42016_n674), .Y(_abc_42016_n1471) );
  AOI21X1 AOI21X1_69 ( .A(_abc_42016_n1486), .B(_abc_42016_n1487), .C(_abc_42016_n1494), .Y(_abc_42016_n1495) );
  AOI21X1 AOI21X1_7 ( .A(_abc_42016_n743), .B(_abc_42016_n744), .C(_abc_42016_n745), .Y(_abc_42016_n746) );
  AOI21X1 AOI21X1_70 ( .A(_abc_42016_n1410_1), .B(_abc_42016_n1474), .C(_abc_42016_n674), .Y(_abc_42016_n1497) );
  AOI21X1 AOI21X1_71 ( .A(_abc_42016_n1506), .B(_abc_42016_n1437), .C(_abc_42016_n1438), .Y(_abc_42016_n1507) );
  AOI21X1 AOI21X1_72 ( .A(_abc_42016_n1513), .B(_abc_42016_n1508), .C(_abc_42016_n1520), .Y(_abc_42016_n1521) );
  AOI21X1 AOI21X1_73 ( .A(_abc_42016_n1410_1), .B(_abc_42016_n1500), .C(_abc_42016_n674), .Y(_abc_42016_n1523) );
  AOI21X1 AOI21X1_74 ( .A(_abc_42016_n1546), .B(_abc_42016_n1547), .C(_abc_42016_n1541), .Y(_abc_42016_n1548) );
  AOI21X1 AOI21X1_75 ( .A(_abc_42016_n1410_1), .B(_abc_42016_n1526), .C(_abc_42016_n674), .Y(_abc_42016_n1550) );
  AOI21X1 AOI21X1_76 ( .A(regfil_7__6_), .B(_abc_42016_n1003), .C(_abc_42016_n1574), .Y(_abc_42016_n1575) );
  AOI21X1 AOI21X1_77 ( .A(regfil_4__6_), .B(_abc_42016_n1426), .C(_abc_42016_n1410_1), .Y(_abc_42016_n1576) );
  AOI21X1 AOI21X1_78 ( .A(_abc_42016_n1569), .B(_abc_42016_n1571), .C(_abc_42016_n1577), .Y(_abc_42016_n1578_1) );
  AOI21X1 AOI21X1_79 ( .A(_abc_42016_n1410_1), .B(_abc_42016_n1553), .C(_abc_42016_n674), .Y(_abc_42016_n1580) );
  AOI21X1 AOI21X1_8 ( .A(_abc_42016_n607), .B(_abc_42016_n750), .C(_abc_42016_n766), .Y(_abc_42016_n767) );
  AOI21X1 AOI21X1_80 ( .A(pc_15_), .B(_abc_42016_n1437), .C(_abc_42016_n1438), .Y(_abc_42016_n1591) );
  AOI21X1 AOI21X1_81 ( .A(_abc_42016_n1588_1), .B(_abc_42016_n1508), .C(_abc_42016_n1599_1), .Y(_abc_42016_n1600_1) );
  AOI21X1 AOI21X1_82 ( .A(_abc_42016_n720), .B(_abc_42016_n1604_1), .C(_abc_42016_n1605_1), .Y(_abc_42016_n1606_1) );
  AOI21X1 AOI21X1_83 ( .A(_abc_42016_n1636), .B(_abc_42016_n685), .C(_abc_42016_n1642), .Y(_abc_42016_n1643) );
  AOI21X1 AOI21X1_84 ( .A(_abc_42016_n751), .B(rdatahold2_1_), .C(_abc_42016_n1658_1), .Y(_abc_42016_n1659) );
  AOI21X1 AOI21X1_85 ( .A(_abc_42016_n696), .B(regfil_4__2_), .C(_abc_42016_n689), .Y(_abc_42016_n1670) );
  AOI21X1 AOI21X1_86 ( .A(_abc_42016_n1675), .B(_abc_42016_n689), .C(_abc_42016_n690), .Y(_abc_42016_n1676) );
  AOI21X1 AOI21X1_87 ( .A(_abc_42016_n1674_1), .B(_abc_42016_n1676), .C(_abc_42016_n1683), .Y(_abc_42016_n1684) );
  AOI21X1 AOI21X1_88 ( .A(_abc_42016_n1690_1), .B(_abc_42016_n1691), .C(_abc_42016_n606), .Y(_abc_42016_n1692) );
  AOI21X1 AOI21X1_89 ( .A(rdatahold_3_), .B(_abc_42016_n694), .C(_abc_42016_n1692), .Y(_abc_42016_n1693) );
  AOI21X1 AOI21X1_9 ( .A(_abc_42016_n630), .B(_abc_42016_n800), .C(_abc_42016_n536), .Y(_abc_42016_n801) );
  AOI21X1 AOI21X1_90 ( .A(rdatahold2_3_), .B(_abc_42016_n751), .C(_abc_42016_n1694), .Y(_abc_42016_n1695) );
  AOI21X1 AOI21X1_91 ( .A(_abc_42016_n1700), .B(_abc_42016_n1699), .C(_abc_42016_n778_1), .Y(_abc_42016_n1701) );
  AOI21X1 AOI21X1_92 ( .A(regfil_4__3_), .B(_abc_42016_n696), .C(_abc_42016_n1701), .Y(_abc_42016_n1702) );
  AOI21X1 AOI21X1_93 ( .A(_abc_42016_n1711), .B(regfil_2__4_), .C(_abc_42016_n772), .Y(_abc_42016_n1712) );
  AOI21X1 AOI21X1_94 ( .A(_abc_42016_n1672), .B(_abc_42016_n796), .C(_abc_42016_n847), .Y(_abc_42016_n1714_1) );
  AOI21X1 AOI21X1_95 ( .A(_abc_42016_n696), .B(regfil_4__4_), .C(_abc_42016_n689), .Y(_abc_42016_n1717) );
  AOI21X1 AOI21X1_96 ( .A(_abc_42016_n660), .B(_abc_42016_n1710), .C(_abc_42016_n1724), .Y(_abc_42016_n1725) );
  AOI21X1 AOI21X1_97 ( .A(_abc_42016_n1624), .B(_abc_42016_n642), .C(_abc_42016_n588_1), .Y(_abc_42016_n1727) );
  AOI21X1 AOI21X1_98 ( .A(_abc_42016_n1736), .B(_abc_42016_n895), .C(_abc_42016_n772), .Y(_abc_42016_n1739) );
  AOI21X1 AOI21X1_99 ( .A(_abc_42016_n660), .B(_abc_42016_n1731), .C(_abc_42016_n1746), .Y(_abc_42016_n1747) );
  AOI22X1 AOI22X1_1 ( .A(_abc_42016_n629), .B(_abc_42016_n630), .C(_abc_42016_n628), .D(_abc_42016_n564), .Y(_abc_42016_n631) );
  AOI22X1 AOI22X1_10 ( .A(_abc_42016_n552), .B(alu_res_3_), .C(rdatahold_3_), .D(_abc_42016_n526_1), .Y(_abc_42016_n807) );
  AOI22X1 AOI22X1_100 ( .A(_abc_42016_n668), .B(regfil_5__7_), .C(sign), .D(_abc_42016_n1003), .Y(_abc_42016_n2719) );
  AOI22X1 AOI22X1_101 ( .A(_abc_42016_n1399), .B(_abc_42016_n2720), .C(regfil_5__7_), .D(_abc_42016_n996), .Y(_abc_42016_n2721) );
  AOI22X1 AOI22X1_102 ( .A(_abc_42016_n2309), .B(_abc_42016_n2528), .C(regfil_5__1_), .D(_abc_42016_n2430), .Y(_abc_42016_n2770) );
  AOI22X1 AOI22X1_103 ( .A(regfil_5__1_), .B(_abc_42016_n2768_1), .C(_abc_42016_n2771), .D(_abc_42016_n2428), .Y(_abc_42016_n2772) );
  AOI22X1 AOI22X1_104 ( .A(_abc_42016_n2765), .B(_abc_42016_n2735), .C(_abc_42016_n2784), .D(_abc_42016_n2774), .Y(raddrhold_1__FF_INPUT) );
  AOI22X1 AOI22X1_105 ( .A(regfil_5__2_), .B(_abc_42016_n2768_1), .C(_abc_42016_n673), .D(_abc_42016_n2798), .Y(_abc_42016_n2799) );
  AOI22X1 AOI22X1_106 ( .A(_abc_42016_n2786), .B(_abc_42016_n2735), .C(_abc_42016_n2791), .D(_abc_42016_n2801), .Y(raddrhold_2__FF_INPUT) );
  AOI22X1 AOI22X1_107 ( .A(_abc_42016_n673), .B(_abc_42016_n2814), .C(_abc_42016_n2815), .D(_abc_42016_n2428), .Y(_abc_42016_n2816) );
  AOI22X1 AOI22X1_108 ( .A(_abc_42016_n2803), .B(_abc_42016_n2735), .C(_abc_42016_n2808), .D(_abc_42016_n2818), .Y(raddrhold_3__FF_INPUT) );
  AOI22X1 AOI22X1_109 ( .A(_abc_42016_n2820), .B(_abc_42016_n2735), .C(_abc_42016_n2834_1), .D(_abc_42016_n2827), .Y(raddrhold_4__FF_INPUT) );
  AOI22X1 AOI22X1_11 ( .A(_abc_42016_n779), .B(_abc_42016_n829), .C(regfil_5__3_), .D(_abc_42016_n696), .Y(_abc_42016_n830) );
  AOI22X1 AOI22X1_110 ( .A(_abc_42016_n673), .B(_abc_42016_n2841), .C(_abc_42016_n2843), .D(_abc_42016_n2428), .Y(_abc_42016_n2844) );
  AOI22X1 AOI22X1_111 ( .A(_abc_42016_n2836), .B(_abc_42016_n2735), .C(_abc_42016_n2850), .D(_abc_42016_n2846), .Y(raddrhold_5__FF_INPUT) );
  AOI22X1 AOI22X1_112 ( .A(_abc_42016_n2852), .B(_abc_42016_n2735), .C(_abc_42016_n2867), .D(_abc_42016_n2861), .Y(raddrhold_6__FF_INPUT) );
  AOI22X1 AOI22X1_113 ( .A(regfil_5__7_), .B(_abc_42016_n2768_1), .C(_abc_42016_n673), .D(_abc_42016_n2876), .Y(_abc_42016_n2877) );
  AOI22X1 AOI22X1_114 ( .A(_abc_42016_n2869), .B(_abc_42016_n2735), .C(_abc_42016_n2885), .D(_abc_42016_n2879_1), .Y(raddrhold_7__FF_INPUT) );
  AOI22X1 AOI22X1_115 ( .A(_abc_42016_n2309), .B(_abc_42016_n1396), .C(_abc_42016_n2893), .D(_abc_42016_n2894), .Y(_abc_42016_n2895) );
  AOI22X1 AOI22X1_116 ( .A(_abc_42016_n673), .B(_abc_42016_n2897), .C(_abc_42016_n2896), .D(_abc_42016_n2428), .Y(_abc_42016_n2898) );
  AOI22X1 AOI22X1_117 ( .A(_abc_42016_n2887), .B(_abc_42016_n2735), .C(_abc_42016_n2891), .D(_abc_42016_n2900_1), .Y(raddrhold_8__FF_INPUT) );
  AOI22X1 AOI22X1_118 ( .A(regfil_4__1_), .B(_abc_42016_n2768_1), .C(_abc_42016_n2909), .D(_abc_42016_n2907), .Y(_abc_42016_n2910) );
  AOI22X1 AOI22X1_119 ( .A(sp_10_), .B(_abc_42016_n2740), .C(_abc_42016_n2743), .D(_abc_42016_n1467), .Y(_abc_42016_n2928) );
  AOI22X1 AOI22X1_12 ( .A(_abc_42016_n842), .B(_abc_42016_n630), .C(_abc_42016_n843), .D(_abc_42016_n625), .Y(_abc_42016_n844) );
  AOI22X1 AOI22X1_120 ( .A(_abc_42016_n2920), .B(_abc_42016_n2735), .C(_abc_42016_n2938), .D(_abc_42016_n2933), .Y(raddrhold_10__FF_INPUT) );
  AOI22X1 AOI22X1_121 ( .A(regfil_4__3_), .B(_abc_42016_n2768_1), .C(_abc_42016_n2909), .D(_abc_42016_n2948), .Y(_abc_42016_n2949) );
  AOI22X1 AOI22X1_122 ( .A(sp_12_), .B(_abc_42016_n2740), .C(_abc_42016_n2743), .D(_abc_42016_n1513), .Y(_abc_42016_n2963) );
  AOI22X1 AOI22X1_123 ( .A(regfil_4__4_), .B(_abc_42016_n2768_1), .C(raddrhold_12_), .D(_abc_42016_n2746), .Y(_abc_42016_n2964) );
  AOI22X1 AOI22X1_124 ( .A(_abc_42016_n2956), .B(_abc_42016_n2735), .C(_abc_42016_n2970_1), .D(_abc_42016_n2966), .Y(raddrhold_12__FF_INPUT) );
  AOI22X1 AOI22X1_125 ( .A(sp_13_), .B(_abc_42016_n2740), .C(_abc_42016_n2743), .D(_abc_42016_n2973), .Y(_abc_42016_n2979) );
  AOI22X1 AOI22X1_126 ( .A(regfil_4__5_), .B(_abc_42016_n2768_1), .C(raddrhold_13_), .D(_abc_42016_n2746), .Y(_abc_42016_n2980) );
  AOI22X1 AOI22X1_127 ( .A(_abc_42016_n2972), .B(_abc_42016_n2735), .C(_abc_42016_n2988), .D(_abc_42016_n2982), .Y(raddrhold_13__FF_INPUT) );
  AOI22X1 AOI22X1_128 ( .A(sp_14_), .B(_abc_42016_n2740), .C(_abc_42016_n2743), .D(_abc_42016_n1563), .Y(_abc_42016_n2992) );
  AOI22X1 AOI22X1_129 ( .A(raddrhold_14_), .B(_abc_42016_n2929), .C(_abc_42016_n2999), .D(_abc_42016_n2997), .Y(_abc_42016_n3000) );
  AOI22X1 AOI22X1_13 ( .A(_abc_42016_n834), .B(_abc_42016_n630), .C(_abc_42016_n847), .D(_abc_42016_n538_1), .Y(_abc_42016_n848) );
  AOI22X1 AOI22X1_130 ( .A(_abc_42016_n2990_1), .B(_abc_42016_n2735), .C(_abc_42016_n3007), .D(_abc_42016_n3002), .Y(raddrhold_14__FF_INPUT) );
  AOI22X1 AOI22X1_131 ( .A(regfil_4__7_), .B(_abc_42016_n2768_1), .C(raddrhold_15_), .D(_abc_42016_n2929), .Y(_abc_42016_n3021) );
  AOI22X1 AOI22X1_132 ( .A(_abc_42016_n3009), .B(_abc_42016_n2735), .C(_abc_42016_n3010), .D(_abc_42016_n3026), .Y(raddrhold_15__FF_INPUT) );
  AOI22X1 AOI22X1_133 ( .A(_abc_42016_n2519), .B(_abc_42016_n3028), .C(rdatahold2_0_), .D(_abc_42016_n3045), .Y(_abc_42016_n3046) );
  AOI22X1 AOI22X1_134 ( .A(_abc_42016_n3028), .B(_abc_42016_n3031), .C(_abc_42016_n3048), .D(_abc_42016_n3044), .Y(waddrhold_0__FF_INPUT) );
  AOI22X1 AOI22X1_135 ( .A(_abc_42016_n3050), .B(_abc_42016_n3031), .C(_abc_42016_n3076), .D(_abc_42016_n3069), .Y(waddrhold_1__FF_INPUT) );
  AOI22X1 AOI22X1_136 ( .A(_abc_42016_n3045), .B(rdatahold2_2_), .C(regfil_5__2_), .D(_abc_42016_n2518_1), .Y(_abc_42016_n3085) );
  AOI22X1 AOI22X1_137 ( .A(sp_2_), .B(_abc_42016_n996), .C(_abc_42016_n3100), .D(_abc_42016_n3056), .Y(_abc_42016_n3101) );
  AOI22X1 AOI22X1_138 ( .A(_abc_42016_n3045), .B(rdatahold2_3_), .C(regfil_5__3_), .D(_abc_42016_n2518_1), .Y(_abc_42016_n3109) );
  AOI22X1 AOI22X1_139 ( .A(sp_3_), .B(_abc_42016_n996), .C(_abc_42016_n3123), .D(_abc_42016_n3056), .Y(_abc_42016_n3124) );
  AOI22X1 AOI22X1_14 ( .A(_abc_42016_n552), .B(alu_res_4_), .C(rdatahold_4_), .D(_abc_42016_n526_1), .Y(_abc_42016_n852) );
  AOI22X1 AOI22X1_140 ( .A(_abc_42016_n1841), .B(_abc_42016_n3138), .C(waddrhold_4_), .D(_abc_42016_n3090), .Y(_abc_42016_n3139) );
  AOI22X1 AOI22X1_141 ( .A(_abc_42016_n3045), .B(rdatahold2_4_), .C(regfil_5__4_), .D(_abc_42016_n2518_1), .Y(_abc_42016_n3149) );
  AOI22X1 AOI22X1_142 ( .A(_abc_42016_n3033), .B(_abc_42016_n2655), .C(_abc_42016_n1841), .D(_abc_42016_n3154), .Y(_abc_42016_n3155) );
  AOI22X1 AOI22X1_143 ( .A(_abc_42016_n3045), .B(rdatahold2_5_), .C(regfil_5__5_), .D(_abc_42016_n2518_1), .Y(_abc_42016_n3169_1) );
  AOI22X1 AOI22X1_144 ( .A(_abc_42016_n3045), .B(rdatahold2_6_), .C(regfil_5__6_), .D(_abc_42016_n2518_1), .Y(_abc_42016_n3197) );
  AOI22X1 AOI22X1_145 ( .A(sp_7_), .B(_abc_42016_n996), .C(waddrhold_7_), .D(_abc_42016_n1410_1), .Y(_abc_42016_n3205) );
  AOI22X1 AOI22X1_146 ( .A(regfil_5__7_), .B(_abc_42016_n2299), .C(waddrhold_7_), .D(_abc_42016_n2359), .Y(_abc_42016_n3212) );
  AOI22X1 AOI22X1_147 ( .A(_abc_42016_n3201), .B(_abc_42016_n3031), .C(_abc_42016_n3221), .D(_abc_42016_n3215), .Y(waddrhold_7__FF_INPUT) );
  AOI22X1 AOI22X1_148 ( .A(sp_8_), .B(_abc_42016_n996), .C(waddrhold_8_), .D(_abc_42016_n1410_1), .Y(_abc_42016_n3228) );
  AOI22X1 AOI22X1_149 ( .A(regfil_4__0_), .B(_abc_42016_n2299), .C(waddrhold_8_), .D(_abc_42016_n2359), .Y(_abc_42016_n3234) );
  AOI22X1 AOI22X1_15 ( .A(rdatahold_4_), .B(_abc_42016_n751), .C(_abc_42016_n853), .D(_abc_42016_n720), .Y(_abc_42016_n854) );
  AOI22X1 AOI22X1_150 ( .A(_abc_42016_n3045), .B(rdatahold_0_), .C(regfil_4__0_), .D(_abc_42016_n2518_1), .Y(_abc_42016_n3241) );
  AOI22X1 AOI22X1_151 ( .A(_abc_42016_n3223), .B(_abc_42016_n3031), .C(_abc_42016_n3237), .D(_abc_42016_n3243), .Y(waddrhold_8__FF_INPUT) );
  AOI22X1 AOI22X1_152 ( .A(_abc_42016_n3245_1), .B(_abc_42016_n3031), .C(_abc_42016_n3266_1), .D(_abc_42016_n3261), .Y(waddrhold_9__FF_INPUT) );
  AOI22X1 AOI22X1_153 ( .A(sp_10_), .B(_abc_42016_n996), .C(waddrhold_10_), .D(_abc_42016_n1410_1), .Y(_abc_42016_n3272) );
  AOI22X1 AOI22X1_154 ( .A(regfil_4__2_), .B(_abc_42016_n2299), .C(waddrhold_10_), .D(_abc_42016_n2359), .Y(_abc_42016_n3280) );
  AOI22X1 AOI22X1_155 ( .A(_abc_42016_n3268), .B(_abc_42016_n3031), .C(_abc_42016_n3283), .D(_abc_42016_n3289), .Y(waddrhold_10__FF_INPUT) );
  AOI22X1 AOI22X1_156 ( .A(sp_11_), .B(_abc_42016_n996), .C(waddrhold_11_), .D(_abc_42016_n1410_1), .Y(_abc_42016_n3299) );
  AOI22X1 AOI22X1_157 ( .A(regfil_4__3_), .B(_abc_42016_n2299), .C(waddrhold_11_), .D(_abc_42016_n2359), .Y(_abc_42016_n3305) );
  AOI22X1 AOI22X1_158 ( .A(_abc_42016_n3045), .B(rdatahold_3_), .C(regfil_4__3_), .D(_abc_42016_n2518_1), .Y(_abc_42016_n3312) );
  AOI22X1 AOI22X1_159 ( .A(sp_12_), .B(_abc_42016_n996), .C(waddrhold_12_), .D(_abc_42016_n1410_1), .Y(_abc_42016_n3322) );
  AOI22X1 AOI22X1_16 ( .A(_abc_42016_n538_1), .B(_abc_42016_n919), .C(_abc_42016_n609), .D(_abc_42016_n625), .Y(_abc_42016_n920) );
  AOI22X1 AOI22X1_160 ( .A(_abc_42016_n1841), .B(_abc_42016_n2957), .C(waddrhold_12_), .D(_abc_42016_n3090), .Y(_abc_42016_n3327) );
  AOI22X1 AOI22X1_161 ( .A(_abc_42016_n3316), .B(_abc_42016_n3031), .C(_abc_42016_n3318_1), .D(_abc_42016_n3335), .Y(waddrhold_12__FF_INPUT) );
  AOI22X1 AOI22X1_162 ( .A(sp_13_), .B(_abc_42016_n996), .C(_abc_42016_n3056), .D(_abc_42016_n3341), .Y(_abc_42016_n3342) );
  AOI22X1 AOI22X1_163 ( .A(_abc_42016_n3337), .B(_abc_42016_n2280), .C(_abc_42016_n2293), .D(_abc_42016_n3346_1), .Y(_abc_42016_n3347) );
  AOI22X1 AOI22X1_164 ( .A(_abc_42016_n3337), .B(_abc_42016_n3031), .C(_abc_42016_n3359), .D(_abc_42016_n3353), .Y(waddrhold_13__FF_INPUT) );
  AOI22X1 AOI22X1_165 ( .A(sp_14_), .B(_abc_42016_n996), .C(waddrhold_14_), .D(_abc_42016_n1410_1), .Y(_abc_42016_n3367) );
  AOI22X1 AOI22X1_166 ( .A(_abc_42016_n3361), .B(_abc_42016_n2280), .C(_abc_42016_n2293), .D(_abc_42016_n3372), .Y(_abc_42016_n3373) );
  AOI22X1 AOI22X1_167 ( .A(_abc_42016_n3361), .B(_abc_42016_n3031), .C(_abc_42016_n3386), .D(_abc_42016_n3379), .Y(waddrhold_14__FF_INPUT) );
  AOI22X1 AOI22X1_168 ( .A(sp_15_), .B(_abc_42016_n996), .C(waddrhold_15_), .D(_abc_42016_n1410_1), .Y(_abc_42016_n3391) );
  AOI22X1 AOI22X1_169 ( .A(regfil_4__7_), .B(_abc_42016_n2299), .C(waddrhold_15_), .D(_abc_42016_n2359), .Y(_abc_42016_n3393) );
  AOI22X1 AOI22X1_17 ( .A(_abc_42016_n625), .B(_abc_42016_n923), .C(_abc_42016_n924), .D(_abc_42016_n564), .Y(_abc_42016_n925) );
  AOI22X1 AOI22X1_170 ( .A(_abc_42016_n1841), .B(_abc_42016_n3395), .C(waddrhold_15_), .D(_abc_42016_n3090), .Y(_abc_42016_n3396) );
  AOI22X1 AOI22X1_171 ( .A(_abc_42016_n3388), .B(_abc_42016_n3031), .C(_abc_42016_n3405), .D(_abc_42016_n3401), .Y(waddrhold_15__FF_INPUT) );
  AOI22X1 AOI22X1_172 ( .A(regfil_7__0_), .B(_abc_42016_n3409), .C(\data[0] ), .D(_abc_42016_n3411), .Y(_abc_42016_n3412) );
  AOI22X1 AOI22X1_173 ( .A(regfil_7__1_), .B(_abc_42016_n3409), .C(\data[1] ), .D(_abc_42016_n3411), .Y(_abc_42016_n3414) );
  AOI22X1 AOI22X1_174 ( .A(regfil_7__2_), .B(_abc_42016_n3409), .C(\data[2] ), .D(_abc_42016_n3411), .Y(_abc_42016_n3416) );
  AOI22X1 AOI22X1_175 ( .A(wdatahold_3_), .B(_abc_42016_n3407), .C(\data[3] ), .D(_abc_42016_n3411), .Y(_abc_42016_n3419) );
  AOI22X1 AOI22X1_176 ( .A(regfil_7__4_), .B(_abc_42016_n3409), .C(\data[4] ), .D(_abc_42016_n3411), .Y(_abc_42016_n3421_1) );
  AOI22X1 AOI22X1_177 ( .A(regfil_7__5_), .B(_abc_42016_n3409), .C(\data[5] ), .D(_abc_42016_n3411), .Y(_abc_42016_n3423) );
  AOI22X1 AOI22X1_178 ( .A(wdatahold_6_), .B(_abc_42016_n3407), .C(\data[6] ), .D(_abc_42016_n3411), .Y(_abc_42016_n3425) );
  AOI22X1 AOI22X1_179 ( .A(regfil_7__7_), .B(_abc_42016_n3409), .C(\data[7] ), .D(_abc_42016_n3411), .Y(_abc_42016_n3427) );
  AOI22X1 AOI22X1_18 ( .A(rdatahold_6_), .B(_abc_42016_n526_1), .C(_abc_42016_n927), .D(_abc_42016_n624), .Y(_abc_42016_n928) );
  AOI22X1 AOI22X1_180 ( .A(_abc_42016_n551), .B(_abc_42016_n3430), .C(_abc_42016_n3435), .D(_abc_42016_n3438), .Y(regd_0__FF_INPUT) );
  AOI22X1 AOI22X1_181 ( .A(_abc_42016_n3455), .B(_abc_42016_n2758), .C(regfil_5__0_), .D(_abc_42016_n3452), .Y(_abc_42016_n3456) );
  AOI22X1 AOI22X1_182 ( .A(_abc_42016_n2775), .B(_abc_42016_n3462), .C(_abc_42016_n3484), .D(_abc_42016_n3482_1), .Y(sp_1__FF_INPUT) );
  AOI22X1 AOI22X1_183 ( .A(sp_2_), .B(_abc_42016_n3453), .C(_abc_42016_n3492), .D(_abc_42016_n3490), .Y(_abc_42016_n3493) );
  AOI22X1 AOI22X1_184 ( .A(_abc_42016_n1159), .B(_abc_42016_n3462), .C(_abc_42016_n3506), .D(_abc_42016_n3500), .Y(sp_2__FF_INPUT) );
  AOI22X1 AOI22X1_185 ( .A(_abc_42016_n2347_1), .B(_abc_42016_n3510_1), .C(_abc_42016_n1407), .D(_abc_42016_n3123), .Y(_abc_42016_n3511) );
  AOI22X1 AOI22X1_186 ( .A(_abc_42016_n3527), .B(_abc_42016_n3123), .C(_abc_42016_n3502), .D(_abc_42016_n3510_1), .Y(_abc_42016_n3528) );
  AOI22X1 AOI22X1_187 ( .A(_abc_42016_n2813), .B(_abc_42016_n3462), .C(_abc_42016_n3530), .D(_abc_42016_n3526_1), .Y(sp_3__FF_INPUT) );
  AOI22X1 AOI22X1_188 ( .A(rdatahold2_4_), .B(_abc_42016_n3459), .C(_abc_42016_n3502), .D(_abc_42016_n3535), .Y(_abc_42016_n3550) );
  AOI22X1 AOI22X1_189 ( .A(_abc_42016_n1210), .B(_abc_42016_n3462), .C(_abc_42016_n3552_1), .D(_abc_42016_n3549), .Y(sp_4__FF_INPUT) );
  AOI22X1 AOI22X1_19 ( .A(_abc_42016_n720), .B(_abc_42016_n929), .C(_abc_42016_n607), .D(_abc_42016_n916), .Y(_abc_42016_n930) );
  AOI22X1 AOI22X1_190 ( .A(_abc_42016_n1279), .B(_abc_42016_n3462), .C(_abc_42016_n3579), .D(_abc_42016_n3574), .Y(sp_5__FF_INPUT) );
  AOI22X1 AOI22X1_191 ( .A(_abc_42016_n1323), .B(_abc_42016_n3462), .C(_abc_42016_n3603), .D(_abc_42016_n3599), .Y(sp_6__FF_INPUT) );
  AOI22X1 AOI22X1_192 ( .A(regfil_5__7_), .B(_abc_42016_n1005), .C(_abc_42016_n2347_1), .D(_abc_42016_n3609), .Y(_abc_42016_n3620) );
  AOI22X1 AOI22X1_193 ( .A(_abc_42016_n1327_1), .B(_abc_42016_n3462), .C(_abc_42016_n3612), .D(_abc_42016_n3624), .Y(sp_7__FF_INPUT) );
  AOI22X1 AOI22X1_194 ( .A(_abc_42016_n2131_1), .B(_abc_42016_n3462), .C(_abc_42016_n3626), .D(_abc_42016_n3647), .Y(sp_8__FF_INPUT) );
  AOI22X1 AOI22X1_195 ( .A(_abc_42016_n2127_1), .B(_abc_42016_n3462), .C(_abc_42016_n3667), .D(_abc_42016_n3664), .Y(sp_9__FF_INPUT) );
  AOI22X1 AOI22X1_196 ( .A(_abc_42016_n2122), .B(_abc_42016_n3462), .C(_abc_42016_n3688), .D(_abc_42016_n3686), .Y(sp_10__FF_INPUT) );
  AOI22X1 AOI22X1_197 ( .A(_abc_42016_n2118), .B(_abc_42016_n3462), .C(_abc_42016_n3711), .D(_abc_42016_n3707), .Y(sp_11__FF_INPUT) );
  AOI22X1 AOI22X1_198 ( .A(rdatahold_4_), .B(_abc_42016_n3459), .C(_abc_42016_n3527), .D(_abc_42016_n3732), .Y(_abc_42016_n3733_1) );
  AOI22X1 AOI22X1_199 ( .A(regfil_4__5_), .B(_abc_42016_n1005), .C(_abc_42016_n2347_1), .D(_abc_42016_n3747), .Y(_abc_42016_n3748) );
  AOI22X1 AOI22X1_2 ( .A(_abc_42016_n608), .B(_abc_42016_n630), .C(_abc_42016_n634), .D(_abc_42016_n564), .Y(_abc_42016_n635) );
  AOI22X1 AOI22X1_20 ( .A(_abc_42016_n779), .B(_abc_42016_n944), .C(regfil_5__6_), .D(_abc_42016_n696), .Y(_abc_42016_n945) );
  AOI22X1 AOI22X1_200 ( .A(rdatahold_5_), .B(_abc_42016_n3459), .C(_abc_42016_n3527), .D(_abc_42016_n3341), .Y(_abc_42016_n3754) );
  AOI22X1 AOI22X1_201 ( .A(_abc_42016_n2103), .B(_abc_42016_n3462), .C(_abc_42016_n3777), .D(_abc_42016_n3774), .Y(sp_14__FF_INPUT) );
  AOI22X1 AOI22X1_202 ( .A(_abc_42016_n2347_1), .B(_abc_42016_n3789), .C(_abc_42016_n1407), .D(_abc_42016_n3389), .Y(_abc_42016_n3790) );
  AOI22X1 AOI22X1_203 ( .A(_abc_42016_n2101), .B(_abc_42016_n3462), .C(_abc_42016_n3797_1), .D(_abc_42016_n3793), .Y(sp_15__FF_INPUT) );
  AOI22X1 AOI22X1_204 ( .A(_abc_42016_n3799), .B(_abc_42016_n3801), .C(_abc_42016_n3831), .D(_abc_42016_n3830), .Y(_abc_36783_n4531) );
  AOI22X1 AOI22X1_205 ( .A(_abc_42016_n3833), .B(_abc_42016_n3835), .C(_abc_42016_n1055), .D(_abc_42016_n3862), .Y(_abc_36783_n4532) );
  AOI22X1 AOI22X1_206 ( .A(_abc_42016_n1036), .B(_abc_42016_n3880), .C(_abc_42016_n1031_1), .D(_abc_42016_n3884), .Y(_abc_42016_n3885) );
  AOI22X1 AOI22X1_207 ( .A(_abc_42016_n3955), .B(_abc_42016_n3956), .C(_abc_42016_n3983_1), .D(_abc_42016_n3982), .Y(_abc_36783_n4536) );
  AOI22X1 AOI22X1_208 ( .A(regfil_4__5_), .B(_abc_42016_n1047_1), .C(_abc_42016_n1225), .D(_abc_42016_n4002), .Y(_abc_42016_n4003) );
  AOI22X1 AOI22X1_209 ( .A(_abc_42016_n3988), .B(_abc_42016_n3989), .C(_abc_42016_n3993), .D(_abc_42016_n4005), .Y(_abc_42016_n4006) );
  AOI22X1 AOI22X1_21 ( .A(_abc_42016_n625), .B(_abc_42016_n959), .C(_abc_42016_n960), .D(_abc_42016_n564), .Y(_abc_42016_n961) );
  AOI22X1 AOI22X1_210 ( .A(_abc_42016_n2478), .B(_abc_42016_n993), .C(_abc_42016_n4015), .D(_abc_42016_n4043), .Y(_abc_42016_n4044) );
  AOI22X1 AOI22X1_211 ( .A(_abc_42016_n1371), .B(_abc_42016_n604_1), .C(_abc_42016_n531), .D(_abc_42016_n569), .Y(_abc_42016_n4083) );
  AOI22X1 AOI22X1_212 ( .A(_abc_42016_n1371), .B(_abc_42016_n1003), .C(_abc_42016_n3052), .D(_abc_42016_n4108), .Y(_abc_42016_n4109) );
  AOI22X1 AOI22X1_213 ( .A(rdatahold2_0_), .B(_abc_42016_n4119), .C(pc_0_), .D(_abc_42016_n4120), .Y(_abc_42016_n4121) );
  AOI22X1 AOI22X1_214 ( .A(_abc_42016_n1383), .B(_abc_42016_n1841), .C(_abc_42016_n2769), .D(_abc_42016_n2285), .Y(_abc_42016_n4125) );
  AOI22X1 AOI22X1_215 ( .A(_abc_42016_n1344), .B(_abc_42016_n2526), .C(_abc_42016_n4135), .D(_abc_42016_n4132), .Y(_abc_42016_n4136) );
  AOI22X1 AOI22X1_216 ( .A(rdatahold2_1_), .B(_abc_42016_n4119), .C(pc_1_), .D(_abc_42016_n4120), .Y(_abc_42016_n4139) );
  AOI22X1 AOI22X1_217 ( .A(regfil_5__2_), .B(_abc_42016_n1006), .C(_abc_42016_n2561), .D(_abc_42016_n4087), .Y(_abc_42016_n4149) );
  AOI22X1 AOI22X1_218 ( .A(_abc_42016_n2561), .B(_abc_42016_n4146), .C(_abc_42016_n4150_1), .D(_abc_42016_n4132), .Y(_abc_42016_n4151) );
  AOI22X1 AOI22X1_219 ( .A(rdatahold2_2_), .B(_abc_42016_n4119), .C(pc_2_), .D(_abc_42016_n4120), .Y(_abc_42016_n4154) );
  AOI22X1 AOI22X1_22 ( .A(_abc_42016_n954), .B(_abc_42016_n630), .C(_abc_42016_n964), .D(_abc_42016_n538_1), .Y(_abc_42016_n965) );
  AOI22X1 AOI22X1_220 ( .A(_abc_42016_n559), .B(_abc_42016_n4162), .C(_abc_42016_n4166), .D(_abc_42016_n4132), .Y(_abc_42016_n4167) );
  AOI22X1 AOI22X1_221 ( .A(rdatahold2_3_), .B(_abc_42016_n4119), .C(pc_3_), .D(_abc_42016_n4120), .Y(_abc_42016_n4170) );
  AOI22X1 AOI22X1_222 ( .A(_abc_42016_n559), .B(_abc_42016_n4175), .C(_abc_42016_n4178), .D(_abc_42016_n4132), .Y(_abc_42016_n4179) );
  AOI22X1 AOI22X1_223 ( .A(rdatahold2_4_), .B(_abc_42016_n4119), .C(pc_4_), .D(_abc_42016_n4120), .Y(_abc_42016_n4182) );
  AOI22X1 AOI22X1_224 ( .A(_abc_42016_n559), .B(_abc_42016_n4188), .C(_abc_42016_n4192), .D(_abc_42016_n4132), .Y(_abc_42016_n4193) );
  AOI22X1 AOI22X1_225 ( .A(rdatahold2_5_), .B(_abc_42016_n4119), .C(pc_5_), .D(_abc_42016_n4120), .Y(_abc_42016_n4196) );
  AOI22X1 AOI22X1_226 ( .A(regfil_5__6_), .B(_abc_42016_n1006), .C(_abc_42016_n4089), .D(_abc_42016_n4200), .Y(_abc_42016_n4203) );
  AOI22X1 AOI22X1_227 ( .A(_abc_42016_n559), .B(_abc_42016_n4202), .C(_abc_42016_n4204_1), .D(_abc_42016_n4132), .Y(_abc_42016_n4205) );
  AOI22X1 AOI22X1_228 ( .A(rdatahold2_6_), .B(_abc_42016_n4119), .C(pc_6_), .D(_abc_42016_n4120), .Y(_abc_42016_n4208) );
  AOI22X1 AOI22X1_229 ( .A(_abc_42016_n1841), .B(_abc_42016_n4212), .C(_abc_42016_n2285), .D(_abc_42016_n2724), .Y(_abc_42016_n4213) );
  AOI22X1 AOI22X1_23 ( .A(alu_res_7_), .B(_abc_42016_n552), .C(_abc_42016_n967), .D(_abc_42016_n624), .Y(_abc_42016_n968) );
  AOI22X1 AOI22X1_230 ( .A(rdatahold2_7_), .B(_abc_42016_n4119), .C(pc_7_), .D(_abc_42016_n4120), .Y(_abc_42016_n4221) );
  AOI22X1 AOI22X1_231 ( .A(_abc_42016_n559), .B(_abc_42016_n4230), .C(_abc_42016_n4229), .D(_abc_42016_n4146), .Y(_abc_42016_n4231) );
  AOI22X1 AOI22X1_232 ( .A(rdatahold_0_), .B(_abc_42016_n4119), .C(pc_8_), .D(_abc_42016_n4120), .Y(_abc_42016_n4234) );
  AOI22X1 AOI22X1_233 ( .A(_abc_42016_n559), .B(_abc_42016_n4243), .C(_abc_42016_n4242), .D(_abc_42016_n4146), .Y(_abc_42016_n4244) );
  AOI22X1 AOI22X1_234 ( .A(rdatahold_1_), .B(_abc_42016_n4119), .C(pc_9_), .D(_abc_42016_n4120), .Y(_abc_42016_n4247) );
  AOI22X1 AOI22X1_235 ( .A(_abc_42016_n4251), .B(_abc_42016_n4089), .C(_abc_42016_n4077), .D(_abc_42016_n4249), .Y(_abc_42016_n4252) );
  AOI22X1 AOI22X1_236 ( .A(regfil_4__2_), .B(_abc_42016_n1006), .C(_abc_42016_n4087), .D(_abc_42016_n1467), .Y(_abc_42016_n4253) );
  AOI22X1 AOI22X1_237 ( .A(_abc_42016_n4251), .B(_abc_42016_n1841), .C(_abc_42016_n2285), .D(_abc_42016_n4249), .Y(_abc_42016_n4255) );
  AOI22X1 AOI22X1_238 ( .A(_abc_42016_n1467), .B(_abc_42016_n4146), .C(pc_10_), .D(_abc_42016_n4210), .Y(_abc_42016_n4256) );
  AOI22X1 AOI22X1_239 ( .A(rdatahold_2_), .B(_abc_42016_n4119), .C(pc_10_), .D(_abc_42016_n4120), .Y(_abc_42016_n4259) );
  AOI22X1 AOI22X1_24 ( .A(rdatahold2_0_), .B(_abc_42016_n1019), .C(_abc_42016_n1043), .D(_abc_42016_n1052), .Y(_abc_42016_n1053) );
  AOI22X1 AOI22X1_240 ( .A(_abc_42016_n559), .B(_abc_42016_n4269), .C(pc_11_), .D(_abc_42016_n4210), .Y(_abc_42016_n4270) );
  AOI22X1 AOI22X1_241 ( .A(rdatahold_3_), .B(_abc_42016_n4119), .C(pc_11_), .D(_abc_42016_n4120), .Y(_abc_42016_n4273) );
  AOI22X1 AOI22X1_242 ( .A(_abc_42016_n1513), .B(_abc_42016_n4146), .C(_abc_42016_n559), .D(_abc_42016_n4281), .Y(_abc_42016_n4282) );
  AOI22X1 AOI22X1_243 ( .A(rdatahold_4_), .B(_abc_42016_n4119), .C(pc_12_), .D(_abc_42016_n4120), .Y(_abc_42016_n4285) );
  AOI22X1 AOI22X1_244 ( .A(_abc_42016_n2973), .B(_abc_42016_n4157), .C(pc_13_), .D(_abc_42016_n4210), .Y(_abc_42016_n4294) );
  AOI22X1 AOI22X1_245 ( .A(rdatahold_5_), .B(_abc_42016_n4119), .C(pc_13_), .D(_abc_42016_n4120), .Y(_abc_42016_n4297) );
  AOI22X1 AOI22X1_246 ( .A(rdatahold_6_), .B(_abc_42016_n4119), .C(pc_14_), .D(_abc_42016_n4311), .Y(_abc_42016_n4312) );
  AOI22X1 AOI22X1_247 ( .A(regfil_4__7_), .B(_abc_42016_n1006), .C(_abc_42016_n4089), .D(_abc_42016_n1586_1), .Y(_abc_42016_n4315) );
  AOI22X1 AOI22X1_248 ( .A(_abc_42016_n1841), .B(_abc_42016_n1586_1), .C(_abc_42016_n2285), .D(_abc_42016_n1589), .Y(_abc_42016_n4317) );
  AOI22X1 AOI22X1_249 ( .A(pc_15_), .B(_abc_42016_n4210), .C(_abc_42016_n4157), .D(_abc_42016_n1588_1), .Y(_abc_42016_n4318) );
  AOI22X1 AOI22X1_25 ( .A(_abc_42016_n1055), .B(_abc_42016_n1134), .C(_abc_42016_n1094), .D(_abc_42016_n1095), .Y(_abc_36783_n3441) );
  AOI22X1 AOI22X1_250 ( .A(rdatahold_7_), .B(_abc_42016_n4119), .C(pc_15_), .D(_abc_42016_n4120), .Y(_abc_42016_n4321) );
  AOI22X1 AOI22X1_251 ( .A(alu_res_0_), .B(_abc_42016_n4057), .C(regfil_7__0_), .D(_abc_42016_n4056), .Y(_abc_42016_n4357) );
  AOI22X1 AOI22X1_252 ( .A(_abc_42016_n4050), .B(regfil_7__0_), .C(regfil_7__2_), .D(_abc_42016_n4059), .Y(_abc_42016_n4363) );
  AOI22X1 AOI22X1_253 ( .A(rdatahold_2_), .B(_abc_42016_n4382), .C(regfil_7__3_), .D(_abc_42016_n4381), .Y(_abc_42016_n4383) );
  AOI22X1 AOI22X1_254 ( .A(_abc_42016_n4050), .B(regfil_7__3_), .C(rdatahold_4_), .D(_abc_42016_n4382), .Y(_abc_42016_n4406) );
  AOI22X1 AOI22X1_255 ( .A(alu_res_4_), .B(_abc_42016_n4057), .C(\data[4] ), .D(_abc_42016_n4047), .Y(_abc_42016_n4410) );
  AOI22X1 AOI22X1_256 ( .A(_abc_42016_n4050), .B(regfil_7__4_), .C(rdatahold_5_), .D(_abc_42016_n4382), .Y(_abc_42016_n4416_1) );
  AOI22X1 AOI22X1_257 ( .A(alu_res_5_), .B(_abc_42016_n4057), .C(\data[5] ), .D(_abc_42016_n4047), .Y(_abc_42016_n4420) );
  AOI22X1 AOI22X1_258 ( .A(alu_res_6_), .B(_abc_42016_n4057), .C(\data[6] ), .D(_abc_42016_n4047), .Y(_abc_42016_n4436) );
  AOI22X1 AOI22X1_259 ( .A(_abc_42016_n4050), .B(regfil_7__6_), .C(_abc_42016_n4059), .D(_abc_42016_n4449), .Y(_abc_42016_n4450) );
  AOI22X1 AOI22X1_26 ( .A(_abc_42016_n1176), .B(_abc_42016_n1177), .C(_abc_42016_n1136), .D(_abc_42016_n1137), .Y(_abc_36783_n3444) );
  AOI22X1 AOI22X1_260 ( .A(_abc_42016_n4446), .B(_abc_42016_n4454), .C(_abc_42016_n4369), .D(_abc_42016_n4456), .Y(_abc_36783_n4586) );
  AOI22X1 AOI22X1_261 ( .A(_abc_42016_n517), .B(_abc_42016_n1872), .C(_abc_42016_n535), .D(_abc_42016_n4561), .Y(_abc_42016_n4562) );
  AOI22X1 AOI22X1_262 ( .A(_abc_42016_n4550), .B(_abc_42016_n4584), .C(_abc_42016_n2438_1), .D(_abc_42016_n4553), .Y(_abc_42016_n4585_1) );
  AOI22X1 AOI22X1_263 ( .A(_abc_42016_n515), .B(_abc_42016_n2078), .C(_abc_42016_n4325), .D(_abc_42016_n2229), .Y(_abc_42016_n4597) );
  AOI22X1 AOI22X1_264 ( .A(_abc_42016_n508), .B(_abc_42016_n517), .C(_abc_42016_n4325), .D(_abc_42016_n4045), .Y(_abc_42016_n4623) );
  AOI22X1 AOI22X1_265 ( .A(_abc_42016_n517), .B(_abc_42016_n2227), .C(_abc_42016_n4325), .D(_abc_42016_n2334), .Y(_abc_42016_n4628) );
  AOI22X1 AOI22X1_266 ( .A(_abc_42016_n1911), .B(_abc_42016_n2050), .C(carry), .D(_abc_42016_n1917), .Y(_abc_42016_n4639) );
  AOI22X1 AOI22X1_267 ( .A(_abc_42016_n4642), .B(_abc_42016_n668), .C(_abc_42016_n532_1), .D(_abc_42016_n4644), .Y(_abc_42016_n4645) );
  AOI22X1 AOI22X1_268 ( .A(_abc_42016_n2408_1), .B(statesel_0_), .C(_abc_42016_n2363), .D(_abc_42016_n4568), .Y(_abc_42016_n4660) );
  AOI22X1 AOI22X1_269 ( .A(_abc_42016_n2768_1), .B(_abc_42016_n557), .C(_abc_42016_n4561), .D(_abc_42016_n4669), .Y(_abc_42016_n4670_1) );
  AOI22X1 AOI22X1_27 ( .A(rdatahold2_4_), .B(_abc_42016_n1019), .C(_abc_42016_n1180), .D(_abc_42016_n1219), .Y(_abc_42016_n1220) );
  AOI22X1 AOI22X1_270 ( .A(_abc_42016_n2446), .B(_abc_42016_n4549), .C(_abc_42016_n2450_1), .D(_abc_42016_n4675), .Y(_abc_42016_n4676_1) );
  AOI22X1 AOI22X1_271 ( .A(_abc_42016_n549), .B(_abc_42016_n4669), .C(_abc_42016_n3033), .D(_abc_42016_n561), .Y(_abc_42016_n4682) );
  AOI22X1 AOI22X1_272 ( .A(_abc_42016_n1871), .B(_abc_42016_n4688_1), .C(_abc_42016_n2302), .D(_abc_42016_n557), .Y(_abc_42016_n4689_1) );
  AOI22X1 AOI22X1_273 ( .A(_abc_42016_n4587), .B(_abc_42016_n4551), .C(_abc_42016_n4578), .D(_abc_42016_n4626), .Y(_abc_42016_n4691) );
  AOI22X1 AOI22X1_274 ( .A(alu__abc_41682_n120), .B(alu__abc_41682_n60), .C(alu__abc_41682_n51), .D(alu__abc_41682_n128), .Y(alu__abc_41682_n129) );
  AOI22X1 AOI22X1_275 ( .A(alu__abc_41682_n114), .B(alu__abc_41682_n94), .C(alu__abc_41682_n117), .D(alu__abc_41682_n130), .Y(alu__abc_41682_n131) );
  AOI22X1 AOI22X1_276 ( .A(alu_oprb_0_), .B(alu__abc_41682_n139), .C(alu__abc_41682_n42), .D(alu__abc_41682_n140), .Y(alu__abc_41682_n141) );
  AOI22X1 AOI22X1_277 ( .A(alu__abc_41682_n74), .B(alu__abc_41682_n75), .C(alu__abc_41682_n134), .D(alu__abc_41682_n144), .Y(alu__abc_41682_n145) );
  AOI22X1 AOI22X1_278 ( .A(alu__abc_41682_n92), .B(alu__abc_41682_n194), .C(alu__abc_41682_n200), .D(alu__abc_41682_n223), .Y(alu__abc_41682_n224) );
  AOI22X1 AOI22X1_279 ( .A(alu__abc_41682_n229), .B(alu__abc_41682_n194), .C(alu__abc_41682_n231), .D(alu__abc_41682_n245), .Y(alu__abc_41682_n246) );
  AOI22X1 AOI22X1_28 ( .A(_abc_42016_n1023), .B(_abc_42016_n1235), .C(_abc_42016_n1240), .D(_abc_42016_n1248_1), .Y(_abc_42016_n1249) );
  AOI22X1 AOI22X1_280 ( .A(alu__abc_41682_n52), .B(alu__abc_41682_n240), .C(alu__abc_41682_n150), .D(alu__abc_41682_n209), .Y(alu__abc_41682_n270_1) );
  AOI22X1 AOI22X1_281 ( .A(alu__abc_41682_n265), .B(alu__abc_41682_n283), .C(alu__abc_41682_n40), .D(alu__abc_41682_n300), .Y(alu__abc_41682_n301) );
  AOI22X1 AOI22X1_29 ( .A(_abc_42016_n1331_1), .B(_abc_42016_n1332), .C(_abc_42016_n1312), .D(_abc_42016_n1322), .Y(_abc_42016_n1333_1) );
  AOI22X1 AOI22X1_3 ( .A(_abc_42016_n722), .B(_abc_42016_n630), .C(_abc_42016_n723), .D(_abc_42016_n538_1), .Y(_abc_42016_n724) );
  AOI22X1 AOI22X1_30 ( .A(_abc_42016_n1339_1), .B(_abc_42016_n1338), .C(regfil_3__7_), .D(_abc_42016_n696), .Y(_abc_42016_n1340) );
  AOI22X1 AOI22X1_31 ( .A(_abc_42016_n1302), .B(_abc_42016_n1057), .C(_abc_42016_n1056), .D(_abc_42016_n1342), .Y(_abc_36783_n3456) );
  AOI22X1 AOI22X1_32 ( .A(_abc_42016_n1351), .B(regfil_4__0_), .C(wdatahold2_0_), .D(_abc_42016_n1349), .Y(_abc_42016_n1352) );
  AOI22X1 AOI22X1_33 ( .A(_abc_42016_n1401), .B(_abc_42016_n1396), .C(regfil_7__0_), .D(_abc_42016_n1402), .Y(_abc_42016_n1403) );
  AOI22X1 AOI22X1_34 ( .A(regfil_0__1_), .B(_abc_42016_n570), .C(regfil_2__1_), .D(_abc_42016_n679), .Y(_abc_42016_n1428) );
  AOI22X1 AOI22X1_35 ( .A(_abc_42016_n559), .B(_abc_42016_n1421), .C(_abc_42016_n1442), .D(_abc_42016_n1441), .Y(_abc_42016_n1443) );
  AOI22X1 AOI22X1_36 ( .A(_abc_42016_n1399), .B(_abc_42016_n1457), .C(regfil_4__2_), .D(_abc_42016_n1426), .Y(_abc_42016_n1458) );
  AOI22X1 AOI22X1_37 ( .A(_abc_42016_n559), .B(_abc_42016_n1448), .C(_abc_42016_n1471), .D(_abc_42016_n1470), .Y(_abc_42016_n1472) );
  AOI22X1 AOI22X1_38 ( .A(regfil_0__3_), .B(_abc_42016_n570), .C(regfil_2__3_), .D(_abc_42016_n679), .Y(_abc_42016_n1489) );
  AOI22X1 AOI22X1_39 ( .A(_abc_42016_n559), .B(_abc_42016_n1476), .C(_abc_42016_n1497), .D(_abc_42016_n1496_1), .Y(_abc_42016_n1498) );
  AOI22X1 AOI22X1_4 ( .A(_abc_42016_n538_1), .B(_abc_42016_n728), .C(_abc_42016_n645), .D(_abc_42016_n625), .Y(_abc_42016_n729) );
  AOI22X1 AOI22X1_40 ( .A(_abc_42016_n1399), .B(_abc_42016_n1516), .C(regfil_7__4_), .D(_abc_42016_n1402), .Y(_abc_42016_n1517) );
  AOI22X1 AOI22X1_41 ( .A(_abc_42016_n559), .B(_abc_42016_n1502), .C(_abc_42016_n1523), .D(_abc_42016_n1522_1), .Y(_abc_42016_n1524) );
  AOI22X1 AOI22X1_42 ( .A(_abc_42016_n1399), .B(_abc_42016_n1538), .C(regfil_4__5_), .D(_abc_42016_n1426), .Y(_abc_42016_n1539) );
  AOI22X1 AOI22X1_43 ( .A(_abc_42016_n559), .B(_abc_42016_n1529), .C(_abc_42016_n1550), .D(_abc_42016_n1549), .Y(_abc_42016_n1551) );
  AOI22X1 AOI22X1_44 ( .A(_abc_42016_n559), .B(_abc_42016_n1556), .C(_abc_42016_n1580), .D(_abc_42016_n1579), .Y(_abc_42016_n1581) );
  AOI22X1 AOI22X1_45 ( .A(_abc_42016_n1351), .B(regfil_4__7_), .C(wdatahold2_7_), .D(_abc_42016_n1349), .Y(_abc_42016_n1583) );
  AOI22X1 AOI22X1_46 ( .A(_abc_42016_n1399), .B(_abc_42016_n1595), .C(regfil_4__7_), .D(_abc_42016_n1426), .Y(_abc_42016_n1596_1) );
  AOI22X1 AOI22X1_47 ( .A(rdatahold_2_), .B(_abc_42016_n1639_1), .C(_abc_42016_n1681_1), .D(_abc_42016_n607), .Y(_abc_42016_n1682_1) );
  AOI22X1 AOI22X1_48 ( .A(rdatahold_4_), .B(_abc_42016_n1639_1), .C(_abc_42016_n1722_1), .D(_abc_42016_n607), .Y(_abc_42016_n1723) );
  AOI22X1 AOI22X1_49 ( .A(regfil_4__5_), .B(_abc_42016_n696), .C(_abc_42016_n1739), .D(_abc_42016_n1738), .Y(_abc_42016_n1740) );
  AOI22X1 AOI22X1_5 ( .A(_abc_42016_n743), .B(_abc_42016_n630), .C(_abc_42016_n753), .D(_abc_42016_n538_1), .Y(_abc_42016_n754) );
  AOI22X1 AOI22X1_50 ( .A(rdatahold_5_), .B(_abc_42016_n1639_1), .C(_abc_42016_n1744), .D(_abc_42016_n607), .Y(_abc_42016_n1745) );
  AOI22X1 AOI22X1_51 ( .A(_abc_42016_n1795), .B(_abc_42016_n1796), .C(_abc_42016_n692), .D(_abc_42016_n1798), .Y(_abc_36783_n3650) );
  AOI22X1 AOI22X1_52 ( .A(_abc_42016_n1809), .B(_abc_42016_n1800), .C(_abc_42016_n692), .D(_abc_42016_n1811), .Y(_abc_36783_n3652) );
  AOI22X1 AOI22X1_53 ( .A(rdatahold_0_), .B(_abc_42016_n1874_1), .C(alu_oprb_0_), .D(_abc_42016_n1875_1), .Y(_abc_42016_n1876) );
  AOI22X1 AOI22X1_54 ( .A(rdatahold_1_), .B(_abc_42016_n1874_1), .C(_abc_42016_n731), .D(_abc_42016_n1882), .Y(_abc_42016_n1883) );
  AOI22X1 AOI22X1_55 ( .A(rdatahold_2_), .B(_abc_42016_n1874_1), .C(_abc_42016_n761), .D(_abc_42016_n1882), .Y(_abc_42016_n1886_1) );
  AOI22X1 AOI22X1_56 ( .A(rdatahold_3_), .B(_abc_42016_n1874_1), .C(_abc_42016_n805), .D(_abc_42016_n1882), .Y(_abc_42016_n1889) );
  AOI22X1 AOI22X1_57 ( .A(rdatahold_4_), .B(_abc_42016_n1874_1), .C(_abc_42016_n850), .D(_abc_42016_n1882), .Y(_abc_42016_n1892) );
  AOI22X1 AOI22X1_58 ( .A(rdatahold_5_), .B(_abc_42016_n1874_1), .C(_abc_42016_n902), .D(_abc_42016_n1882), .Y(_abc_42016_n1895) );
  AOI22X1 AOI22X1_59 ( .A(rdatahold_6_), .B(_abc_42016_n1874_1), .C(_abc_42016_n927), .D(_abc_42016_n1882), .Y(_abc_42016_n1898) );
  AOI22X1 AOI22X1_6 ( .A(_abc_42016_n538_1), .B(_abc_42016_n758), .C(_abc_42016_n757), .D(_abc_42016_n625), .Y(_abc_42016_n759) );
  AOI22X1 AOI22X1_60 ( .A(alu_oprb_7_), .B(_abc_42016_n1880), .C(_abc_42016_n1851), .D(_abc_42016_n967), .Y(_abc_42016_n1900) );
  AOI22X1 AOI22X1_61 ( .A(rdatahold_7_), .B(_abc_42016_n1874_1), .C(alu_oprb_7_), .D(_abc_42016_n1875_1), .Y(_abc_42016_n1901_1) );
  AOI22X1 AOI22X1_62 ( .A(regfil_4__1_), .B(_abc_42016_n1911), .C(regfil_6__1_), .D(_abc_42016_n532_1), .Y(_abc_42016_n1936) );
  AOI22X1 AOI22X1_63 ( .A(_abc_42016_n532_1), .B(regfil_2__1_), .C(regfil_1__1_), .D(_abc_42016_n1915), .Y(_abc_42016_n1939) );
  AOI22X1 AOI22X1_64 ( .A(_abc_42016_n1930), .B(rdatahold_1_), .C(alu_opra_1_), .D(_abc_42016_n1925), .Y(_abc_42016_n1946) );
  AOI22X1 AOI22X1_65 ( .A(_abc_42016_n1911), .B(regfil_4__2_), .C(regfil_7__2_), .D(_abc_42016_n1917), .Y(_abc_42016_n1953) );
  AOI22X1 AOI22X1_66 ( .A(regfil_4__3_), .B(_abc_42016_n1911), .C(regfil_5__3_), .D(_abc_42016_n1915), .Y(_abc_42016_n1962) );
  AOI22X1 AOI22X1_67 ( .A(_abc_42016_n532_1), .B(regfil_2__3_), .C(regfil_1__3_), .D(_abc_42016_n1915), .Y(_abc_42016_n1965) );
  AOI22X1 AOI22X1_68 ( .A(_abc_42016_n1930), .B(rdatahold_3_), .C(alu_opra_3_), .D(_abc_42016_n1925), .Y(_abc_42016_n1972) );
  AOI22X1 AOI22X1_69 ( .A(_abc_42016_n532_1), .B(regfil_6__4_), .C(regfil_5__4_), .D(_abc_42016_n1915), .Y(_abc_42016_n1976) );
  AOI22X1 AOI22X1_7 ( .A(_abc_42016_n552), .B(alu_res_2_), .C(rdatahold_2_), .D(_abc_42016_n526_1), .Y(_abc_42016_n763_1) );
  AOI22X1 AOI22X1_70 ( .A(_abc_42016_n1930), .B(rdatahold_4_), .C(alu_opra_4_), .D(_abc_42016_n1925), .Y(_abc_42016_n1985) );
  AOI22X1 AOI22X1_71 ( .A(regfil_0__5_), .B(_abc_42016_n1911), .C(regfil_1__5_), .D(_abc_42016_n1915), .Y(_abc_42016_n1988) );
  AOI22X1 AOI22X1_72 ( .A(_abc_42016_n1930), .B(rdatahold_5_), .C(alu_opra_5_), .D(_abc_42016_n1925), .Y(_abc_42016_n1998) );
  AOI22X1 AOI22X1_73 ( .A(_abc_42016_n1915), .B(regfil_5__6_), .C(regfil_7__6_), .D(_abc_42016_n1917), .Y(_abc_42016_n2004) );
  AOI22X1 AOI22X1_74 ( .A(_abc_42016_n1930), .B(rdatahold_6_), .C(alu_opra_6_), .D(_abc_42016_n1925), .Y(_abc_42016_n2009) );
  AOI22X1 AOI22X1_75 ( .A(regfil_0__7_), .B(_abc_42016_n1911), .C(regfil_1__7_), .D(_abc_42016_n1915), .Y(_abc_42016_n2015) );
  AOI22X1 AOI22X1_76 ( .A(_abc_42016_n1930), .B(rdatahold_7_), .C(alu_opra_7_), .D(_abc_42016_n1925), .Y(_abc_42016_n2022) );
  AOI22X1 AOI22X1_77 ( .A(_abc_42016_n582_1), .B(_abc_42016_n2053), .C(alu_zout), .D(_abc_42016_n2051), .Y(_abc_42016_n2054) );
  AOI22X1 AOI22X1_78 ( .A(_abc_42016_n2036), .B(alu_auxcar), .C(auxcar), .D(_abc_42016_n2047), .Y(_abc_42016_n2074) );
  AOI22X1 AOI22X1_79 ( .A(_abc_42016_n1860), .B(_abc_42016_n2082), .C(_abc_42016_n2223), .D(_abc_42016_n2216), .Y(carry_FF_INPUT) );
  AOI22X1 AOI22X1_8 ( .A(rdatahold_2_), .B(_abc_42016_n751), .C(_abc_42016_n764), .D(_abc_42016_n720), .Y(_abc_42016_n765) );
  AOI22X1 AOI22X1_80 ( .A(_abc_42016_n2259), .B(_abc_42016_n2278), .C(_abc_42016_n2342), .D(_abc_42016_n2333), .Y(statesel_0__FF_INPUT) );
  AOI22X1 AOI22X1_81 ( .A(_abc_42016_n2344), .B(_abc_42016_n2278), .C(_abc_42016_n2367), .D(_abc_42016_n2362), .Y(statesel_1__FF_INPUT) );
  AOI22X1 AOI22X1_82 ( .A(_abc_42016_n2369), .B(_abc_42016_n2278), .C(_abc_42016_n2382), .D(_abc_42016_n2392), .Y(statesel_2__FF_INPUT) );
  AOI22X1 AOI22X1_83 ( .A(_abc_42016_n2394_1), .B(_abc_42016_n2278), .C(_abc_42016_n2415), .D(_abc_42016_n2406), .Y(statesel_3__FF_INPUT) );
  AOI22X1 AOI22X1_84 ( .A(_abc_42016_n2417_1), .B(_abc_42016_n2278), .C(_abc_42016_n2444_1), .D(_abc_42016_n2435_1), .Y(statesel_4__FF_INPUT) );
  AOI22X1 AOI22X1_85 ( .A(_abc_42016_n674), .B(_abc_42016_n2422), .C(_abc_42016_n2446), .D(_abc_42016_n2431), .Y(_abc_42016_n2447_1) );
  AOI22X1 AOI22X1_86 ( .A(_abc_42016_n2411_1), .B(_abc_42016_n2453), .C(_abc_42016_n2336), .D(_abc_42016_n2452), .Y(_abc_42016_n2454) );
  AOI22X1 AOI22X1_87 ( .A(_abc_42016_n2446), .B(_abc_42016_n2278), .C(_abc_42016_n2455_1), .D(_abc_42016_n2449), .Y(statesel_5__FF_INPUT) );
  AOI22X1 AOI22X1_88 ( .A(wdatahold2_0_), .B(_abc_42016_n2519), .C(alu_res_0_), .D(_abc_42016_n2518_1), .Y(_abc_42016_n2520) );
  AOI22X1 AOI22X1_89 ( .A(wdatahold2_1_), .B(_abc_42016_n2519), .C(alu_res_1_), .D(_abc_42016_n2518_1), .Y(_abc_42016_n2550) );
  AOI22X1 AOI22X1_9 ( .A(regfil_0__3_), .B(_abc_42016_n630), .C(regfil_1__3_), .D(_abc_42016_n625), .Y(_abc_42016_n793) );
  AOI22X1 AOI22X1_90 ( .A(wdatahold2_2_), .B(_abc_42016_n2519), .C(alu_res_2_), .D(_abc_42016_n2518_1), .Y(_abc_42016_n2556) );
  AOI22X1 AOI22X1_91 ( .A(_abc_42016_n2614), .B(rdatahold_3_), .C(wdatahold2_3_), .D(_abc_42016_n2519), .Y(_abc_42016_n2615) );
  AOI22X1 AOI22X1_92 ( .A(_abc_42016_n2587), .B(_abc_42016_n2499), .C(_abc_42016_n2617), .D(_abc_42016_n2611), .Y(wdatahold_3__FF_INPUT) );
  AOI22X1 AOI22X1_93 ( .A(wdatahold2_4_), .B(_abc_42016_n2519), .C(alu_res_4_), .D(_abc_42016_n2518_1), .Y(_abc_42016_n2620) );
  AOI22X1 AOI22X1_94 ( .A(_abc_42016_n2619), .B(_abc_42016_n2499), .C(_abc_42016_n2620), .D(_abc_42016_n2646), .Y(wdatahold_4__FF_INPUT) );
  AOI22X1 AOI22X1_95 ( .A(rdatahold_5_), .B(_abc_42016_n2614), .C(alu_res_5_), .D(_abc_42016_n2518_1), .Y(_abc_42016_n2670) );
  AOI22X1 AOI22X1_96 ( .A(_abc_42016_n2648), .B(_abc_42016_n2499), .C(_abc_42016_n2672_1), .D(_abc_42016_n2669), .Y(wdatahold_5__FF_INPUT) );
  AOI22X1 AOI22X1_97 ( .A(regfil_1__6_), .B(_abc_42016_n570), .C(regfil_3__6_), .D(_abc_42016_n679), .Y(_abc_42016_n2678) );
  AOI22X1 AOI22X1_98 ( .A(_abc_42016_n1399), .B(_abc_42016_n2682), .C(regfil_5__6_), .D(_abc_42016_n996), .Y(_abc_42016_n2683) );
  AOI22X1 AOI22X1_99 ( .A(_abc_42016_n2614), .B(rdatahold_6_), .C(wdatahold2_6_), .D(_abc_42016_n2519), .Y(_abc_42016_n2696) );
  BUFX2 BUFX2_1 ( .A(_auto_iopadmap_cc_313_execute_46257_0_), .Y(\addr[0] ) );
  BUFX2 BUFX2_10 ( .A(_auto_iopadmap_cc_313_execute_46257_9_), .Y(\addr[9] ) );
  BUFX2 BUFX2_11 ( .A(_auto_iopadmap_cc_313_execute_46257_10_), .Y(\addr[10] ) );
  BUFX2 BUFX2_12 ( .A(_auto_iopadmap_cc_313_execute_46257_11_), .Y(\addr[11] ) );
  BUFX2 BUFX2_13 ( .A(_auto_iopadmap_cc_313_execute_46257_12_), .Y(\addr[12] ) );
  BUFX2 BUFX2_14 ( .A(_auto_iopadmap_cc_313_execute_46257_13_), .Y(\addr[13] ) );
  BUFX2 BUFX2_15 ( .A(_auto_iopadmap_cc_313_execute_46257_14_), .Y(\addr[14] ) );
  BUFX2 BUFX2_16 ( .A(_auto_iopadmap_cc_313_execute_46257_15_), .Y(\addr[15] ) );
  BUFX2 BUFX2_17 ( .A(_auto_iopadmap_cc_313_execute_46274), .Y(inta) );
  BUFX2 BUFX2_18 ( .A(_auto_iopadmap_cc_313_execute_46276), .Y(readio) );
  BUFX2 BUFX2_19 ( .A(_auto_iopadmap_cc_313_execute_46278), .Y(readmem) );
  BUFX2 BUFX2_2 ( .A(_auto_iopadmap_cc_313_execute_46257_1_), .Y(\addr[1] ) );
  BUFX2 BUFX2_20 ( .A(_auto_iopadmap_cc_313_execute_46280), .Y(writeio) );
  BUFX2 BUFX2_21 ( .A(_auto_iopadmap_cc_313_execute_46282), .Y(writemem) );
  BUFX2 BUFX2_3 ( .A(_auto_iopadmap_cc_313_execute_46257_2_), .Y(\addr[2] ) );
  BUFX2 BUFX2_4 ( .A(_auto_iopadmap_cc_313_execute_46257_3_), .Y(\addr[3] ) );
  BUFX2 BUFX2_5 ( .A(_auto_iopadmap_cc_313_execute_46257_4_), .Y(\addr[4] ) );
  BUFX2 BUFX2_6 ( .A(_auto_iopadmap_cc_313_execute_46257_5_), .Y(\addr[5] ) );
  BUFX2 BUFX2_7 ( .A(_auto_iopadmap_cc_313_execute_46257_6_), .Y(\addr[6] ) );
  BUFX2 BUFX2_8 ( .A(_auto_iopadmap_cc_313_execute_46257_7_), .Y(\addr[7] ) );
  BUFX2 BUFX2_9 ( .A(_auto_iopadmap_cc_313_execute_46257_8_), .Y(\addr[8] ) );
  DFFPOSX1 DFFPOSX1_1 ( .CLK(clock), .D(_abc_36783_n4644), .Q(state_0_) );
  DFFPOSX1 DFFPOSX1_10 ( .CLK(clock), .D(_abc_36783_n3644), .Q(regfil_2__3_) );
  DFFPOSX1 DFFPOSX1_100 ( .CLK(clock), .D(sp_8__FF_INPUT), .Q(sp_8_) );
  DFFPOSX1 DFFPOSX1_101 ( .CLK(clock), .D(sp_9__FF_INPUT), .Q(sp_9_) );
  DFFPOSX1 DFFPOSX1_102 ( .CLK(clock), .D(sp_10__FF_INPUT), .Q(sp_10_) );
  DFFPOSX1 DFFPOSX1_103 ( .CLK(clock), .D(sp_11__FF_INPUT), .Q(sp_11_) );
  DFFPOSX1 DFFPOSX1_104 ( .CLK(clock), .D(sp_12__FF_INPUT), .Q(sp_12_) );
  DFFPOSX1 DFFPOSX1_105 ( .CLK(clock), .D(sp_13__FF_INPUT), .Q(sp_13_) );
  DFFPOSX1 DFFPOSX1_106 ( .CLK(clock), .D(sp_14__FF_INPUT), .Q(sp_14_) );
  DFFPOSX1 DFFPOSX1_107 ( .CLK(clock), .D(sp_15__FF_INPUT), .Q(sp_15_) );
  DFFPOSX1 DFFPOSX1_108 ( .CLK(clock), .D(regd_0__FF_INPUT), .Q(regd_0_) );
  DFFPOSX1 DFFPOSX1_109 ( .CLK(clock), .D(regd_1__FF_INPUT), .Q(regd_1_) );
  DFFPOSX1 DFFPOSX1_11 ( .CLK(clock), .D(_abc_36783_n3646), .Q(regfil_2__4_) );
  DFFPOSX1 DFFPOSX1_110 ( .CLK(clock), .D(regd_2__FF_INPUT), .Q(regd_2_) );
  DFFPOSX1 DFFPOSX1_111 ( .CLK(clock), .D(datao_0__FF_INPUT), .Q(\data[0] ) );
  DFFPOSX1 DFFPOSX1_112 ( .CLK(clock), .D(datao_1__FF_INPUT), .Q(\data[1] ) );
  DFFPOSX1 DFFPOSX1_113 ( .CLK(clock), .D(datao_2__FF_INPUT), .Q(\data[2] ) );
  DFFPOSX1 DFFPOSX1_114 ( .CLK(clock), .D(datao_3__FF_INPUT), .Q(\data[3] ) );
  DFFPOSX1 DFFPOSX1_115 ( .CLK(clock), .D(datao_4__FF_INPUT), .Q(\data[4] ) );
  DFFPOSX1 DFFPOSX1_116 ( .CLK(clock), .D(datao_5__FF_INPUT), .Q(\data[5] ) );
  DFFPOSX1 DFFPOSX1_117 ( .CLK(clock), .D(datao_6__FF_INPUT), .Q(\data[6] ) );
  DFFPOSX1 DFFPOSX1_118 ( .CLK(clock), .D(datao_7__FF_INPUT), .Q(\data[7] ) );
  DFFPOSX1 DFFPOSX1_119 ( .CLK(clock), .D(waddrhold_0__FF_INPUT), .Q(waddrhold_0_) );
  DFFPOSX1 DFFPOSX1_12 ( .CLK(clock), .D(_abc_36783_n3648), .Q(regfil_2__5_) );
  DFFPOSX1 DFFPOSX1_120 ( .CLK(clock), .D(waddrhold_1__FF_INPUT), .Q(waddrhold_1_) );
  DFFPOSX1 DFFPOSX1_121 ( .CLK(clock), .D(waddrhold_2__FF_INPUT), .Q(waddrhold_2_) );
  DFFPOSX1 DFFPOSX1_122 ( .CLK(clock), .D(waddrhold_3__FF_INPUT), .Q(waddrhold_3_) );
  DFFPOSX1 DFFPOSX1_123 ( .CLK(clock), .D(waddrhold_4__FF_INPUT), .Q(waddrhold_4_) );
  DFFPOSX1 DFFPOSX1_124 ( .CLK(clock), .D(waddrhold_5__FF_INPUT), .Q(waddrhold_5_) );
  DFFPOSX1 DFFPOSX1_125 ( .CLK(clock), .D(waddrhold_6__FF_INPUT), .Q(waddrhold_6_) );
  DFFPOSX1 DFFPOSX1_126 ( .CLK(clock), .D(waddrhold_7__FF_INPUT), .Q(waddrhold_7_) );
  DFFPOSX1 DFFPOSX1_127 ( .CLK(clock), .D(waddrhold_8__FF_INPUT), .Q(waddrhold_8_) );
  DFFPOSX1 DFFPOSX1_128 ( .CLK(clock), .D(waddrhold_9__FF_INPUT), .Q(waddrhold_9_) );
  DFFPOSX1 DFFPOSX1_129 ( .CLK(clock), .D(waddrhold_10__FF_INPUT), .Q(waddrhold_10_) );
  DFFPOSX1 DFFPOSX1_13 ( .CLK(clock), .D(_abc_36783_n3650), .Q(regfil_2__6_) );
  DFFPOSX1 DFFPOSX1_130 ( .CLK(clock), .D(waddrhold_11__FF_INPUT), .Q(waddrhold_11_) );
  DFFPOSX1 DFFPOSX1_131 ( .CLK(clock), .D(waddrhold_12__FF_INPUT), .Q(waddrhold_12_) );
  DFFPOSX1 DFFPOSX1_132 ( .CLK(clock), .D(waddrhold_13__FF_INPUT), .Q(waddrhold_13_) );
  DFFPOSX1 DFFPOSX1_133 ( .CLK(clock), .D(waddrhold_14__FF_INPUT), .Q(waddrhold_14_) );
  DFFPOSX1 DFFPOSX1_134 ( .CLK(clock), .D(waddrhold_15__FF_INPUT), .Q(waddrhold_15_) );
  DFFPOSX1 DFFPOSX1_135 ( .CLK(clock), .D(raddrhold_0__FF_INPUT), .Q(raddrhold_0_) );
  DFFPOSX1 DFFPOSX1_136 ( .CLK(clock), .D(raddrhold_1__FF_INPUT), .Q(raddrhold_1_) );
  DFFPOSX1 DFFPOSX1_137 ( .CLK(clock), .D(raddrhold_2__FF_INPUT), .Q(raddrhold_2_) );
  DFFPOSX1 DFFPOSX1_138 ( .CLK(clock), .D(raddrhold_3__FF_INPUT), .Q(raddrhold_3_) );
  DFFPOSX1 DFFPOSX1_139 ( .CLK(clock), .D(raddrhold_4__FF_INPUT), .Q(raddrhold_4_) );
  DFFPOSX1 DFFPOSX1_14 ( .CLK(clock), .D(_abc_36783_n3652), .Q(regfil_2__7_) );
  DFFPOSX1 DFFPOSX1_140 ( .CLK(clock), .D(raddrhold_5__FF_INPUT), .Q(raddrhold_5_) );
  DFFPOSX1 DFFPOSX1_141 ( .CLK(clock), .D(raddrhold_6__FF_INPUT), .Q(raddrhold_6_) );
  DFFPOSX1 DFFPOSX1_142 ( .CLK(clock), .D(raddrhold_7__FF_INPUT), .Q(raddrhold_7_) );
  DFFPOSX1 DFFPOSX1_143 ( .CLK(clock), .D(raddrhold_8__FF_INPUT), .Q(raddrhold_8_) );
  DFFPOSX1 DFFPOSX1_144 ( .CLK(clock), .D(raddrhold_9__FF_INPUT), .Q(raddrhold_9_) );
  DFFPOSX1 DFFPOSX1_145 ( .CLK(clock), .D(raddrhold_10__FF_INPUT), .Q(raddrhold_10_) );
  DFFPOSX1 DFFPOSX1_146 ( .CLK(clock), .D(raddrhold_11__FF_INPUT), .Q(raddrhold_11_) );
  DFFPOSX1 DFFPOSX1_147 ( .CLK(clock), .D(raddrhold_12__FF_INPUT), .Q(raddrhold_12_) );
  DFFPOSX1 DFFPOSX1_148 ( .CLK(clock), .D(raddrhold_13__FF_INPUT), .Q(raddrhold_13_) );
  DFFPOSX1 DFFPOSX1_149 ( .CLK(clock), .D(raddrhold_14__FF_INPUT), .Q(raddrhold_14_) );
  DFFPOSX1 DFFPOSX1_15 ( .CLK(clock), .D(_abc_36783_n3520), .Q(regfil_0__0_) );
  DFFPOSX1 DFFPOSX1_150 ( .CLK(clock), .D(raddrhold_15__FF_INPUT), .Q(raddrhold_15_) );
  DFFPOSX1 DFFPOSX1_151 ( .CLK(clock), .D(wdatahold_0__FF_INPUT), .Q(wdatahold_0_) );
  DFFPOSX1 DFFPOSX1_152 ( .CLK(clock), .D(wdatahold_1__FF_INPUT), .Q(wdatahold_1_) );
  DFFPOSX1 DFFPOSX1_153 ( .CLK(clock), .D(wdatahold_2__FF_INPUT), .Q(wdatahold_2_) );
  DFFPOSX1 DFFPOSX1_154 ( .CLK(clock), .D(wdatahold_3__FF_INPUT), .Q(wdatahold_3_) );
  DFFPOSX1 DFFPOSX1_155 ( .CLK(clock), .D(wdatahold_4__FF_INPUT), .Q(wdatahold_4_) );
  DFFPOSX1 DFFPOSX1_156 ( .CLK(clock), .D(wdatahold_5__FF_INPUT), .Q(wdatahold_5_) );
  DFFPOSX1 DFFPOSX1_157 ( .CLK(clock), .D(wdatahold_6__FF_INPUT), .Q(wdatahold_6_) );
  DFFPOSX1 DFFPOSX1_158 ( .CLK(clock), .D(wdatahold_7__FF_INPUT), .Q(wdatahold_7_) );
  DFFPOSX1 DFFPOSX1_159 ( .CLK(clock), .D(wdatahold2_0__FF_INPUT), .Q(wdatahold2_0_) );
  DFFPOSX1 DFFPOSX1_16 ( .CLK(clock), .D(_abc_36783_n3523), .Q(regfil_0__1_) );
  DFFPOSX1 DFFPOSX1_160 ( .CLK(clock), .D(wdatahold2_1__FF_INPUT), .Q(wdatahold2_1_) );
  DFFPOSX1 DFFPOSX1_161 ( .CLK(clock), .D(wdatahold2_2__FF_INPUT), .Q(wdatahold2_2_) );
  DFFPOSX1 DFFPOSX1_162 ( .CLK(clock), .D(wdatahold2_3__FF_INPUT), .Q(wdatahold2_3_) );
  DFFPOSX1 DFFPOSX1_163 ( .CLK(clock), .D(wdatahold2_4__FF_INPUT), .Q(wdatahold2_4_) );
  DFFPOSX1 DFFPOSX1_164 ( .CLK(clock), .D(wdatahold2_5__FF_INPUT), .Q(wdatahold2_5_) );
  DFFPOSX1 DFFPOSX1_165 ( .CLK(clock), .D(wdatahold2_6__FF_INPUT), .Q(wdatahold2_6_) );
  DFFPOSX1 DFFPOSX1_166 ( .CLK(clock), .D(wdatahold2_7__FF_INPUT), .Q(wdatahold2_7_) );
  DFFPOSX1 DFFPOSX1_167 ( .CLK(clock), .D(rdatahold_0__FF_INPUT), .Q(rdatahold_0_) );
  DFFPOSX1 DFFPOSX1_168 ( .CLK(clock), .D(rdatahold_1__FF_INPUT), .Q(rdatahold_1_) );
  DFFPOSX1 DFFPOSX1_169 ( .CLK(clock), .D(rdatahold_2__FF_INPUT), .Q(rdatahold_2_) );
  DFFPOSX1 DFFPOSX1_17 ( .CLK(clock), .D(_abc_36783_n3526), .Q(regfil_0__2_) );
  DFFPOSX1 DFFPOSX1_170 ( .CLK(clock), .D(rdatahold_3__FF_INPUT), .Q(rdatahold_3_) );
  DFFPOSX1 DFFPOSX1_171 ( .CLK(clock), .D(rdatahold_4__FF_INPUT), .Q(rdatahold_4_) );
  DFFPOSX1 DFFPOSX1_172 ( .CLK(clock), .D(rdatahold_5__FF_INPUT), .Q(rdatahold_5_) );
  DFFPOSX1 DFFPOSX1_173 ( .CLK(clock), .D(rdatahold_6__FF_INPUT), .Q(rdatahold_6_) );
  DFFPOSX1 DFFPOSX1_174 ( .CLK(clock), .D(rdatahold_7__FF_INPUT), .Q(rdatahold_7_) );
  DFFPOSX1 DFFPOSX1_175 ( .CLK(clock), .D(rdatahold2_0__FF_INPUT), .Q(rdatahold2_0_) );
  DFFPOSX1 DFFPOSX1_176 ( .CLK(clock), .D(rdatahold2_1__FF_INPUT), .Q(rdatahold2_1_) );
  DFFPOSX1 DFFPOSX1_177 ( .CLK(clock), .D(rdatahold2_2__FF_INPUT), .Q(rdatahold2_2_) );
  DFFPOSX1 DFFPOSX1_178 ( .CLK(clock), .D(rdatahold2_3__FF_INPUT), .Q(rdatahold2_3_) );
  DFFPOSX1 DFFPOSX1_179 ( .CLK(clock), .D(rdatahold2_4__FF_INPUT), .Q(rdatahold2_4_) );
  DFFPOSX1 DFFPOSX1_18 ( .CLK(clock), .D(_abc_36783_n3529), .Q(regfil_0__3_) );
  DFFPOSX1 DFFPOSX1_180 ( .CLK(clock), .D(rdatahold2_5__FF_INPUT), .Q(rdatahold2_5_) );
  DFFPOSX1 DFFPOSX1_181 ( .CLK(clock), .D(rdatahold2_6__FF_INPUT), .Q(rdatahold2_6_) );
  DFFPOSX1 DFFPOSX1_182 ( .CLK(clock), .D(rdatahold2_7__FF_INPUT), .Q(rdatahold2_7_) );
  DFFPOSX1 DFFPOSX1_183 ( .CLK(clock), .D(popdes_0__FF_INPUT), .Q(popdes_0_) );
  DFFPOSX1 DFFPOSX1_184 ( .CLK(clock), .D(popdes_1__FF_INPUT), .Q(popdes_1_) );
  DFFPOSX1 DFFPOSX1_185 ( .CLK(clock), .D(statesel_0__FF_INPUT), .Q(statesel_0_) );
  DFFPOSX1 DFFPOSX1_186 ( .CLK(clock), .D(statesel_1__FF_INPUT), .Q(statesel_1_) );
  DFFPOSX1 DFFPOSX1_187 ( .CLK(clock), .D(statesel_2__FF_INPUT), .Q(statesel_2_) );
  DFFPOSX1 DFFPOSX1_188 ( .CLK(clock), .D(statesel_3__FF_INPUT), .Q(statesel_3_) );
  DFFPOSX1 DFFPOSX1_189 ( .CLK(clock), .D(statesel_4__FF_INPUT), .Q(statesel_4_) );
  DFFPOSX1 DFFPOSX1_19 ( .CLK(clock), .D(_abc_36783_n3532), .Q(regfil_0__4_) );
  DFFPOSX1 DFFPOSX1_190 ( .CLK(clock), .D(statesel_5__FF_INPUT), .Q(statesel_5_) );
  DFFPOSX1 DFFPOSX1_191 ( .CLK(clock), .D(eienb_FF_INPUT), .Q(eienb) );
  DFFPOSX1 DFFPOSX1_192 ( .CLK(clock), .D(opcode_0__FF_INPUT), .Q(opcode_0_) );
  DFFPOSX1 DFFPOSX1_193 ( .CLK(clock), .D(opcode_1__FF_INPUT), .Q(opcode_1_) );
  DFFPOSX1 DFFPOSX1_194 ( .CLK(clock), .D(opcode_2__FF_INPUT), .Q(opcode_2_) );
  DFFPOSX1 DFFPOSX1_195 ( .CLK(clock), .D(opcode_3__FF_INPUT), .Q(opcode_3_) );
  DFFPOSX1 DFFPOSX1_196 ( .CLK(clock), .D(opcode_4__FF_INPUT), .Q(opcode_4_) );
  DFFPOSX1 DFFPOSX1_197 ( .CLK(clock), .D(opcode_5__FF_INPUT), .Q(opcode_5_) );
  DFFPOSX1 DFFPOSX1_198 ( .CLK(clock), .D(opcode_6__FF_INPUT), .Q(opcode_6_) );
  DFFPOSX1 DFFPOSX1_199 ( .CLK(clock), .D(opcode_7__FF_INPUT), .Q(opcode_7_) );
  DFFPOSX1 DFFPOSX1_2 ( .CLK(clock), .D(_abc_36783_n4645), .Q(state_1_) );
  DFFPOSX1 DFFPOSX1_20 ( .CLK(clock), .D(_abc_36783_n3535), .Q(regfil_0__5_) );
  DFFPOSX1 DFFPOSX1_200 ( .CLK(clock), .D(carry_FF_INPUT), .Q(carry) );
  DFFPOSX1 DFFPOSX1_201 ( .CLK(clock), .D(auxcar_FF_INPUT), .Q(auxcar) );
  DFFPOSX1 DFFPOSX1_202 ( .CLK(clock), .D(sign_FF_INPUT), .Q(sign) );
  DFFPOSX1 DFFPOSX1_203 ( .CLK(clock), .D(zero_FF_INPUT), .Q(zero) );
  DFFPOSX1 DFFPOSX1_204 ( .CLK(clock), .D(parity_FF_INPUT), .Q(parity) );
  DFFPOSX1 DFFPOSX1_205 ( .CLK(clock), .D(ei_FF_INPUT), .Q(ei) );
  DFFPOSX1 DFFPOSX1_206 ( .CLK(clock), .D(intcyc_FF_INPUT), .Q(intcyc) );
  DFFPOSX1 DFFPOSX1_207 ( .CLK(clock), .D(aluopra_0__FF_INPUT), .Q(alu_opra_0_) );
  DFFPOSX1 DFFPOSX1_208 ( .CLK(clock), .D(aluopra_1__FF_INPUT), .Q(alu_opra_1_) );
  DFFPOSX1 DFFPOSX1_209 ( .CLK(clock), .D(aluopra_2__FF_INPUT), .Q(alu_opra_2_) );
  DFFPOSX1 DFFPOSX1_21 ( .CLK(clock), .D(_abc_36783_n3538), .Q(regfil_0__6_) );
  DFFPOSX1 DFFPOSX1_210 ( .CLK(clock), .D(aluopra_3__FF_INPUT), .Q(alu_opra_3_) );
  DFFPOSX1 DFFPOSX1_211 ( .CLK(clock), .D(aluopra_4__FF_INPUT), .Q(alu_opra_4_) );
  DFFPOSX1 DFFPOSX1_212 ( .CLK(clock), .D(aluopra_5__FF_INPUT), .Q(alu_opra_5_) );
  DFFPOSX1 DFFPOSX1_213 ( .CLK(clock), .D(aluopra_6__FF_INPUT), .Q(alu_opra_6_) );
  DFFPOSX1 DFFPOSX1_214 ( .CLK(clock), .D(aluopra_7__FF_INPUT), .Q(alu_opra_7_) );
  DFFPOSX1 DFFPOSX1_215 ( .CLK(clock), .D(aluoprb_0__FF_INPUT), .Q(alu_oprb_0_) );
  DFFPOSX1 DFFPOSX1_216 ( .CLK(clock), .D(aluoprb_1__FF_INPUT), .Q(alu_oprb_1_) );
  DFFPOSX1 DFFPOSX1_217 ( .CLK(clock), .D(aluoprb_2__FF_INPUT), .Q(alu_oprb_2_) );
  DFFPOSX1 DFFPOSX1_218 ( .CLK(clock), .D(aluoprb_3__FF_INPUT), .Q(alu_oprb_3_) );
  DFFPOSX1 DFFPOSX1_219 ( .CLK(clock), .D(aluoprb_4__FF_INPUT), .Q(alu_oprb_4_) );
  DFFPOSX1 DFFPOSX1_22 ( .CLK(clock), .D(_abc_36783_n3541), .Q(regfil_0__7_) );
  DFFPOSX1 DFFPOSX1_220 ( .CLK(clock), .D(aluoprb_5__FF_INPUT), .Q(alu_oprb_5_) );
  DFFPOSX1 DFFPOSX1_221 ( .CLK(clock), .D(aluoprb_6__FF_INPUT), .Q(alu_oprb_6_) );
  DFFPOSX1 DFFPOSX1_222 ( .CLK(clock), .D(aluoprb_7__FF_INPUT), .Q(alu_oprb_7_) );
  DFFPOSX1 DFFPOSX1_223 ( .CLK(clock), .D(alucin_FF_INPUT), .Q(alu_cin) );
  DFFPOSX1 DFFPOSX1_224 ( .CLK(clock), .D(alusel_0__FF_INPUT), .Q(alu_sel_0_) );
  DFFPOSX1 DFFPOSX1_225 ( .CLK(clock), .D(alusel_1__FF_INPUT), .Q(alu_sel_1_) );
  DFFPOSX1 DFFPOSX1_226 ( .CLK(clock), .D(alusel_2__FF_INPUT), .Q(alu_sel_2_) );
  DFFPOSX1 DFFPOSX1_227 ( .CLK(clock), .D(_abc_36783_n4531), .Q(regfil_4__0_) );
  DFFPOSX1 DFFPOSX1_228 ( .CLK(clock), .D(_abc_36783_n4532), .Q(regfil_4__1_) );
  DFFPOSX1 DFFPOSX1_229 ( .CLK(clock), .D(_abc_36783_n4533), .Q(regfil_4__2_) );
  DFFPOSX1 DFFPOSX1_23 ( .CLK(clock), .D(_abc_36783_n3731), .Q(regfil_6__0_) );
  DFFPOSX1 DFFPOSX1_230 ( .CLK(clock), .D(_abc_36783_n4534), .Q(regfil_4__3_) );
  DFFPOSX1 DFFPOSX1_231 ( .CLK(clock), .D(_abc_36783_n4535), .Q(regfil_4__4_) );
  DFFPOSX1 DFFPOSX1_232 ( .CLK(clock), .D(_abc_36783_n4536), .Q(regfil_4__5_) );
  DFFPOSX1 DFFPOSX1_233 ( .CLK(clock), .D(_abc_36783_n4537), .Q(regfil_4__6_) );
  DFFPOSX1 DFFPOSX1_234 ( .CLK(clock), .D(_abc_36783_n4538), .Q(regfil_4__7_) );
  DFFPOSX1 DFFPOSX1_235 ( .CLK(clock), .D(_abc_36783_n4579), .Q(regfil_7__0_) );
  DFFPOSX1 DFFPOSX1_236 ( .CLK(clock), .D(_abc_36783_n4580), .Q(regfil_7__1_) );
  DFFPOSX1 DFFPOSX1_237 ( .CLK(clock), .D(_abc_36783_n4581), .Q(regfil_7__2_) );
  DFFPOSX1 DFFPOSX1_238 ( .CLK(clock), .D(_abc_36783_n4582), .Q(regfil_7__3_) );
  DFFPOSX1 DFFPOSX1_239 ( .CLK(clock), .D(_abc_36783_n4583), .Q(regfil_7__4_) );
  DFFPOSX1 DFFPOSX1_24 ( .CLK(clock), .D(_abc_36783_n3732), .Q(regfil_6__1_) );
  DFFPOSX1 DFFPOSX1_240 ( .CLK(clock), .D(_abc_36783_n4584), .Q(regfil_7__5_) );
  DFFPOSX1 DFFPOSX1_241 ( .CLK(clock), .D(_abc_36783_n4585), .Q(regfil_7__6_) );
  DFFPOSX1 DFFPOSX1_242 ( .CLK(clock), .D(_abc_36783_n4586), .Q(regfil_7__7_) );
  DFFPOSX1 DFFPOSX1_25 ( .CLK(clock), .D(_abc_36783_n3733), .Q(regfil_6__2_) );
  DFFPOSX1 DFFPOSX1_26 ( .CLK(clock), .D(_abc_36783_n3734), .Q(regfil_6__3_) );
  DFFPOSX1 DFFPOSX1_27 ( .CLK(clock), .D(_abc_36783_n3735), .Q(regfil_6__4_) );
  DFFPOSX1 DFFPOSX1_28 ( .CLK(clock), .D(_abc_36783_n3736), .Q(regfil_6__5_) );
  DFFPOSX1 DFFPOSX1_29 ( .CLK(clock), .D(_abc_36783_n3737), .Q(regfil_6__6_) );
  DFFPOSX1 DFFPOSX1_3 ( .CLK(clock), .D(_abc_36783_n4646), .Q(state_2_) );
  DFFPOSX1 DFFPOSX1_30 ( .CLK(clock), .D(_abc_36783_n3738), .Q(regfil_6__7_) );
  DFFPOSX1 DFFPOSX1_31 ( .CLK(clock), .D(_abc_36783_n3361), .Q(regfil_3__0_) );
  DFFPOSX1 DFFPOSX1_32 ( .CLK(clock), .D(_abc_36783_n3364), .Q(regfil_3__1_) );
  DFFPOSX1 DFFPOSX1_33 ( .CLK(clock), .D(_abc_36783_n3367), .Q(regfil_3__2_) );
  DFFPOSX1 DFFPOSX1_34 ( .CLK(clock), .D(_abc_36783_n3370), .Q(regfil_3__3_) );
  DFFPOSX1 DFFPOSX1_35 ( .CLK(clock), .D(_abc_36783_n3373), .Q(regfil_3__4_) );
  DFFPOSX1 DFFPOSX1_36 ( .CLK(clock), .D(_abc_36783_n3376), .Q(regfil_3__5_) );
  DFFPOSX1 DFFPOSX1_37 ( .CLK(clock), .D(_abc_36783_n3379), .Q(regfil_3__6_) );
  DFFPOSX1 DFFPOSX1_38 ( .CLK(clock), .D(_abc_36783_n3382), .Q(regfil_3__7_) );
  DFFPOSX1 DFFPOSX1_39 ( .CLK(clock), .D(_abc_36783_n3554), .Q(regfil_1__0_) );
  DFFPOSX1 DFFPOSX1_4 ( .CLK(clock), .D(_abc_36783_n4647), .Q(state_3_) );
  DFFPOSX1 DFFPOSX1_40 ( .CLK(clock), .D(_abc_36783_n3557), .Q(regfil_1__1_) );
  DFFPOSX1 DFFPOSX1_41 ( .CLK(clock), .D(_abc_36783_n3560), .Q(regfil_1__2_) );
  DFFPOSX1 DFFPOSX1_42 ( .CLK(clock), .D(_abc_36783_n3563), .Q(regfil_1__3_) );
  DFFPOSX1 DFFPOSX1_43 ( .CLK(clock), .D(_abc_36783_n3566), .Q(regfil_1__4_) );
  DFFPOSX1 DFFPOSX1_44 ( .CLK(clock), .D(_abc_36783_n3569), .Q(regfil_1__5_) );
  DFFPOSX1 DFFPOSX1_45 ( .CLK(clock), .D(_abc_36783_n3572), .Q(regfil_1__6_) );
  DFFPOSX1 DFFPOSX1_46 ( .CLK(clock), .D(_abc_36783_n3575), .Q(regfil_1__7_) );
  DFFPOSX1 DFFPOSX1_47 ( .CLK(clock), .D(_abc_36783_n3435), .Q(regfil_5__0_) );
  DFFPOSX1 DFFPOSX1_48 ( .CLK(clock), .D(_abc_36783_n3438), .Q(regfil_5__1_) );
  DFFPOSX1 DFFPOSX1_49 ( .CLK(clock), .D(_abc_36783_n3441), .Q(regfil_5__2_) );
  DFFPOSX1 DFFPOSX1_5 ( .CLK(clock), .D(_abc_36783_n4648), .Q(state_4_) );
  DFFPOSX1 DFFPOSX1_50 ( .CLK(clock), .D(_abc_36783_n3444), .Q(regfil_5__3_) );
  DFFPOSX1 DFFPOSX1_51 ( .CLK(clock), .D(_abc_36783_n3447), .Q(regfil_5__4_) );
  DFFPOSX1 DFFPOSX1_52 ( .CLK(clock), .D(_abc_36783_n3450), .Q(regfil_5__5_) );
  DFFPOSX1 DFFPOSX1_53 ( .CLK(clock), .D(_abc_36783_n3453), .Q(regfil_5__6_) );
  DFFPOSX1 DFFPOSX1_54 ( .CLK(clock), .D(_abc_36783_n3456), .Q(regfil_5__7_) );
  DFFPOSX1 DFFPOSX1_55 ( .CLK(clock), .D(addr_0__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_46257_0_) );
  DFFPOSX1 DFFPOSX1_56 ( .CLK(clock), .D(addr_1__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_46257_1_) );
  DFFPOSX1 DFFPOSX1_57 ( .CLK(clock), .D(addr_2__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_46257_2_) );
  DFFPOSX1 DFFPOSX1_58 ( .CLK(clock), .D(addr_3__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_46257_3_) );
  DFFPOSX1 DFFPOSX1_59 ( .CLK(clock), .D(addr_4__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_46257_4_) );
  DFFPOSX1 DFFPOSX1_6 ( .CLK(clock), .D(_abc_36783_n4649), .Q(state_5_) );
  DFFPOSX1 DFFPOSX1_60 ( .CLK(clock), .D(addr_5__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_46257_5_) );
  DFFPOSX1 DFFPOSX1_61 ( .CLK(clock), .D(addr_6__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_46257_6_) );
  DFFPOSX1 DFFPOSX1_62 ( .CLK(clock), .D(addr_7__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_46257_7_) );
  DFFPOSX1 DFFPOSX1_63 ( .CLK(clock), .D(addr_8__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_46257_8_) );
  DFFPOSX1 DFFPOSX1_64 ( .CLK(clock), .D(addr_9__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_46257_9_) );
  DFFPOSX1 DFFPOSX1_65 ( .CLK(clock), .D(addr_10__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_46257_10_) );
  DFFPOSX1 DFFPOSX1_66 ( .CLK(clock), .D(addr_11__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_46257_11_) );
  DFFPOSX1 DFFPOSX1_67 ( .CLK(clock), .D(addr_12__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_46257_12_) );
  DFFPOSX1 DFFPOSX1_68 ( .CLK(clock), .D(addr_13__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_46257_13_) );
  DFFPOSX1 DFFPOSX1_69 ( .CLK(clock), .D(addr_14__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_46257_14_) );
  DFFPOSX1 DFFPOSX1_7 ( .CLK(clock), .D(_abc_36783_n3638), .Q(regfil_2__0_) );
  DFFPOSX1 DFFPOSX1_70 ( .CLK(clock), .D(addr_15__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_46257_15_) );
  DFFPOSX1 DFFPOSX1_71 ( .CLK(clock), .D(readmem_FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_46278) );
  DFFPOSX1 DFFPOSX1_72 ( .CLK(clock), .D(writemem_FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_46282) );
  DFFPOSX1 DFFPOSX1_73 ( .CLK(clock), .D(readio_FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_46276) );
  DFFPOSX1 DFFPOSX1_74 ( .CLK(clock), .D(writeio_FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_46280) );
  DFFPOSX1 DFFPOSX1_75 ( .CLK(clock), .D(inta_FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_46274) );
  DFFPOSX1 DFFPOSX1_76 ( .CLK(clock), .D(pc_0__FF_INPUT), .Q(pc_0_) );
  DFFPOSX1 DFFPOSX1_77 ( .CLK(clock), .D(pc_1__FF_INPUT), .Q(pc_1_) );
  DFFPOSX1 DFFPOSX1_78 ( .CLK(clock), .D(pc_2__FF_INPUT), .Q(pc_2_) );
  DFFPOSX1 DFFPOSX1_79 ( .CLK(clock), .D(pc_3__FF_INPUT), .Q(pc_3_) );
  DFFPOSX1 DFFPOSX1_8 ( .CLK(clock), .D(_abc_36783_n3640), .Q(regfil_2__1_) );
  DFFPOSX1 DFFPOSX1_80 ( .CLK(clock), .D(pc_4__FF_INPUT), .Q(pc_4_) );
  DFFPOSX1 DFFPOSX1_81 ( .CLK(clock), .D(pc_5__FF_INPUT), .Q(pc_5_) );
  DFFPOSX1 DFFPOSX1_82 ( .CLK(clock), .D(pc_6__FF_INPUT), .Q(pc_6_) );
  DFFPOSX1 DFFPOSX1_83 ( .CLK(clock), .D(pc_7__FF_INPUT), .Q(pc_7_) );
  DFFPOSX1 DFFPOSX1_84 ( .CLK(clock), .D(pc_8__FF_INPUT), .Q(pc_8_) );
  DFFPOSX1 DFFPOSX1_85 ( .CLK(clock), .D(pc_9__FF_INPUT), .Q(pc_9_) );
  DFFPOSX1 DFFPOSX1_86 ( .CLK(clock), .D(pc_10__FF_INPUT), .Q(pc_10_) );
  DFFPOSX1 DFFPOSX1_87 ( .CLK(clock), .D(pc_11__FF_INPUT), .Q(pc_11_) );
  DFFPOSX1 DFFPOSX1_88 ( .CLK(clock), .D(pc_12__FF_INPUT), .Q(pc_12_) );
  DFFPOSX1 DFFPOSX1_89 ( .CLK(clock), .D(pc_13__FF_INPUT), .Q(pc_13_) );
  DFFPOSX1 DFFPOSX1_9 ( .CLK(clock), .D(_abc_36783_n3642), .Q(regfil_2__2_) );
  DFFPOSX1 DFFPOSX1_90 ( .CLK(clock), .D(pc_14__FF_INPUT), .Q(pc_14_) );
  DFFPOSX1 DFFPOSX1_91 ( .CLK(clock), .D(pc_15__FF_INPUT), .Q(pc_15_) );
  DFFPOSX1 DFFPOSX1_92 ( .CLK(clock), .D(sp_0__FF_INPUT), .Q(sp_0_) );
  DFFPOSX1 DFFPOSX1_93 ( .CLK(clock), .D(sp_1__FF_INPUT), .Q(sp_1_) );
  DFFPOSX1 DFFPOSX1_94 ( .CLK(clock), .D(sp_2__FF_INPUT), .Q(sp_2_) );
  DFFPOSX1 DFFPOSX1_95 ( .CLK(clock), .D(sp_3__FF_INPUT), .Q(sp_3_) );
  DFFPOSX1 DFFPOSX1_96 ( .CLK(clock), .D(sp_4__FF_INPUT), .Q(sp_4_) );
  DFFPOSX1 DFFPOSX1_97 ( .CLK(clock), .D(sp_5__FF_INPUT), .Q(sp_5_) );
  DFFPOSX1 DFFPOSX1_98 ( .CLK(clock), .D(sp_6__FF_INPUT), .Q(sp_6_) );
  DFFPOSX1 DFFPOSX1_99 ( .CLK(clock), .D(sp_7__FF_INPUT), .Q(sp_7_) );
  INVX1 INVX1_1 ( .A(state_2_), .Y(_abc_42016_n501) );
  INVX1 INVX1_10 ( .A(_abc_42016_n515), .Y(_abc_42016_n516) );
  INVX1 INVX1_100 ( .A(_abc_42016_n587), .Y(_abc_42016_n751) );
  INVX1 INVX1_101 ( .A(regfil_2__2_), .Y(_abc_42016_n753) );
  INVX1 INVX1_102 ( .A(regfil_5__2_), .Y(_abc_42016_n757) );
  INVX1 INVX1_103 ( .A(regfil_6__2_), .Y(_abc_42016_n758) );
  INVX1 INVX1_104 ( .A(_abc_42016_n765), .Y(_abc_42016_n766) );
  INVX1 INVX1_105 ( .A(_abc_42016_n768), .Y(_abc_42016_n769) );
  INVX1 INVX1_106 ( .A(regfil_3__2_), .Y(_abc_42016_n773) );
  INVX1 INVX1_107 ( .A(_abc_42016_n778_1), .Y(_abc_42016_n779) );
  INVX1 INVX1_108 ( .A(_abc_42016_n780), .Y(_abc_42016_n781) );
  INVX1 INVX1_109 ( .A(_abc_42016_n702_1), .Y(_abc_42016_n782) );
  INVX1 INVX1_11 ( .A(_abc_42016_n517), .Y(_abc_42016_n518_1) );
  INVX1 INVX1_110 ( .A(_abc_42016_n789), .Y(_abc_42016_n790) );
  INVX1 INVX1_111 ( .A(_abc_42016_n793), .Y(_abc_42016_n794) );
  INVX1 INVX1_112 ( .A(regfil_3__3_), .Y(_abc_42016_n795) );
  INVX1 INVX1_113 ( .A(regfil_2__3_), .Y(_abc_42016_n796) );
  INVX1 INVX1_114 ( .A(regfil_6__3_), .Y(_abc_42016_n799) );
  INVX1 INVX1_115 ( .A(regfil_4__3_), .Y(_abc_42016_n800) );
  INVX1 INVX1_116 ( .A(_abc_42016_n805), .Y(_abc_42016_n806) );
  INVX1 INVX1_117 ( .A(rdatahold_3_), .Y(_abc_42016_n811) );
  INVX1 INVX1_118 ( .A(regfil_0__3_), .Y(_abc_42016_n812) );
  INVX1 INVX1_119 ( .A(_abc_42016_n818), .Y(_abc_42016_n819) );
  INVX1 INVX1_12 ( .A(_abc_42016_n519), .Y(_abc_42016_n520) );
  INVX1 INVX1_120 ( .A(_abc_42016_n772), .Y(_abc_42016_n822) );
  INVX1 INVX1_121 ( .A(_abc_42016_n824), .Y(_abc_42016_n825) );
  INVX1 INVX1_122 ( .A(regfil_0__4_), .Y(_abc_42016_n834) );
  INVX1 INVX1_123 ( .A(_abc_42016_n836), .Y(_abc_42016_n837) );
  INVX1 INVX1_124 ( .A(regfil_4__4_), .Y(_abc_42016_n842) );
  INVX1 INVX1_125 ( .A(regfil_5__4_), .Y(_abc_42016_n843) );
  INVX1 INVX1_126 ( .A(regfil_2__4_), .Y(_abc_42016_n847) );
  INVX1 INVX1_127 ( .A(_abc_42016_n854), .Y(_abc_42016_n855) );
  INVX1 INVX1_128 ( .A(_abc_42016_n857), .Y(_abc_42016_n858) );
  INVX1 INVX1_129 ( .A(regfil_3__4_), .Y(_abc_42016_n861) );
  INVX1 INVX1_13 ( .A(state_3_), .Y(_abc_42016_n521) );
  INVX1 INVX1_130 ( .A(regfil_5__5_), .Y(_abc_42016_n872) );
  INVX1 INVX1_131 ( .A(regfil_3__5_), .Y(_abc_42016_n874) );
  INVX1 INVX1_132 ( .A(_abc_42016_n877), .Y(_abc_42016_n878) );
  INVX1 INVX1_133 ( .A(_abc_42016_n887), .Y(_abc_42016_n888) );
  INVX1 INVX1_134 ( .A(rdatahold_5_), .Y(_abc_42016_n891) );
  INVX1 INVX1_135 ( .A(regfil_0__5_), .Y(_abc_42016_n893) );
  INVX1 INVX1_136 ( .A(regfil_2__5_), .Y(_abc_42016_n895) );
  INVX1 INVX1_137 ( .A(regfil_7__5_), .Y(_abc_42016_n898) );
  INVX1 INVX1_138 ( .A(regfil_0__6_), .Y(_abc_42016_n913) );
  INVX1 INVX1_139 ( .A(regfil_2__6_), .Y(_abc_42016_n919) );
  INVX1 INVX1_14 ( .A(_abc_42016_n522), .Y(_abc_42016_n523_1) );
  INVX1 INVX1_140 ( .A(regfil_5__6_), .Y(_abc_42016_n923) );
  INVX1 INVX1_141 ( .A(regfil_7__6_), .Y(_abc_42016_n924) );
  INVX1 INVX1_142 ( .A(regfil_3__6_), .Y(_abc_42016_n939) );
  INVX1 INVX1_143 ( .A(regfil_0__7_), .Y(_abc_42016_n954) );
  INVX1 INVX1_144 ( .A(regfil_5__7_), .Y(_abc_42016_n959) );
  INVX1 INVX1_145 ( .A(regfil_7__7_), .Y(_abc_42016_n960) );
  INVX1 INVX1_146 ( .A(regfil_2__7_), .Y(_abc_42016_n964) );
  INVX1 INVX1_147 ( .A(regfil_3__7_), .Y(_abc_42016_n974) );
  INVX1 INVX1_148 ( .A(_abc_42016_n976), .Y(_abc_42016_n977) );
  INVX1 INVX1_149 ( .A(_abc_42016_n938), .Y(_abc_42016_n979_1) );
  INVX1 INVX1_15 ( .A(_abc_42016_n524_1), .Y(_abc_42016_n525) );
  INVX1 INVX1_150 ( .A(_abc_42016_n987), .Y(_abc_42016_n988) );
  INVX1 INVX1_151 ( .A(_abc_42016_n989), .Y(_abc_42016_n990) );
  INVX1 INVX1_152 ( .A(popdes_1_), .Y(_abc_42016_n992) );
  INVX1 INVX1_153 ( .A(_abc_42016_n993), .Y(_abc_42016_n994) );
  INVX1 INVX1_154 ( .A(_abc_42016_n998), .Y(_abc_42016_n999) );
  INVX1 INVX1_155 ( .A(_abc_42016_n1003), .Y(_abc_42016_n1004) );
  INVX1 INVX1_156 ( .A(_abc_42016_n1008), .Y(_abc_42016_n1009) );
  INVX1 INVX1_157 ( .A(_abc_42016_n1011), .Y(_abc_42016_n1012) );
  INVX1 INVX1_158 ( .A(_abc_42016_n1015), .Y(_abc_42016_n1016) );
  INVX1 INVX1_159 ( .A(_abc_42016_n1005), .Y(_abc_42016_n1022) );
  INVX1 INVX1_16 ( .A(_abc_42016_n526_1), .Y(_abc_42016_n527) );
  INVX1 INVX1_160 ( .A(_abc_42016_n1024), .Y(_abc_42016_n1025) );
  INVX1 INVX1_161 ( .A(_abc_42016_n1028), .Y(_abc_42016_n1029) );
  INVX1 INVX1_162 ( .A(_abc_42016_n1030), .Y(_abc_42016_n1031_1) );
  INVX1 INVX1_163 ( .A(_abc_42016_n1001_1), .Y(_abc_42016_n1035) );
  INVX1 INVX1_164 ( .A(rdatahold2_0_), .Y(_abc_42016_n1044) );
  INVX1 INVX1_165 ( .A(_abc_42016_n1023), .Y(_abc_42016_n1045) );
  INVX1 INVX1_166 ( .A(_abc_42016_n1006), .Y(_abc_42016_n1046) );
  INVX1 INVX1_167 ( .A(_abc_42016_n1047_1), .Y(_abc_42016_n1048) );
  INVX1 INVX1_168 ( .A(_abc_42016_n1020), .Y(_abc_42016_n1055) );
  INVX1 INVX1_169 ( .A(_abc_42016_n1019), .Y(_abc_42016_n1056) );
  INVX1 INVX1_17 ( .A(reset), .Y(_abc_42016_n529) );
  INVX1 INVX1_170 ( .A(_abc_42016_n1058), .Y(_abc_42016_n1059) );
  INVX1 INVX1_171 ( .A(_abc_42016_n996), .Y(_abc_42016_n1061) );
  INVX1 INVX1_172 ( .A(_abc_42016_n1064), .Y(_abc_42016_n1065) );
  INVX1 INVX1_173 ( .A(_abc_42016_n1069), .Y(_abc_42016_n1070_1) );
  INVX1 INVX1_174 ( .A(_abc_42016_n1033), .Y(_abc_42016_n1078) );
  INVX1 INVX1_175 ( .A(_abc_42016_n1000), .Y(_abc_42016_n1082) );
  INVX1 INVX1_176 ( .A(rdatahold2_2_), .Y(_abc_42016_n1130) );
  INVX1 INVX1_177 ( .A(regfil_5__3_), .Y(_abc_42016_n1139) );
  INVX1 INVX1_178 ( .A(_abc_42016_n1102), .Y(_abc_42016_n1147_1) );
  INVX1 INVX1_179 ( .A(_abc_42016_n1145), .Y(_abc_42016_n1149_1) );
  INVX1 INVX1_18 ( .A(opcode_5_), .Y(_abc_42016_n530) );
  INVX1 INVX1_180 ( .A(_abc_42016_n1036), .Y(_abc_42016_n1151) );
  INVX1 INVX1_181 ( .A(sp_2_), .Y(_abc_42016_n1159) );
  INVX1 INVX1_182 ( .A(_abc_42016_n1161), .Y(_abc_42016_n1162) );
  INVX1 INVX1_183 ( .A(_abc_42016_n1160), .Y(_abc_42016_n1165) );
  INVX1 INVX1_184 ( .A(_abc_42016_n1125), .Y(_abc_42016_n1170) );
  INVX1 INVX1_185 ( .A(rdatahold2_3_), .Y(_abc_42016_n1174_1) );
  INVX1 INVX1_186 ( .A(rdatahold2_4_), .Y(_abc_42016_n1179) );
  INVX1 INVX1_187 ( .A(_abc_42016_n1138), .Y(_abc_42016_n1187) );
  INVX1 INVX1_188 ( .A(_abc_42016_n1194), .Y(_abc_42016_n1198) );
  INVX1 INVX1_189 ( .A(sp_4_), .Y(_abc_42016_n1210) );
  INVX1 INVX1_19 ( .A(opcode_4_), .Y(_abc_42016_n531) );
  INVX1 INVX1_190 ( .A(_abc_42016_n1040), .Y(_abc_42016_n1225) );
  INVX1 INVX1_191 ( .A(_abc_42016_n1211), .Y(_abc_42016_n1229) );
  INVX1 INVX1_192 ( .A(_abc_42016_n1233), .Y(_abc_42016_n1234) );
  INVX1 INVX1_193 ( .A(_abc_42016_n1237), .Y(_abc_42016_n1238) );
  INVX1 INVX1_194 ( .A(_abc_42016_n1184), .Y(_abc_42016_n1252) );
  INVX1 INVX1_195 ( .A(rdatahold2_6_), .Y(_abc_42016_n1261) );
  INVX1 INVX1_196 ( .A(sp_5_), .Y(_abc_42016_n1279) );
  INVX1 INVX1_197 ( .A(_abc_42016_n1284), .Y(_abc_42016_n1285) );
  INVX1 INVX1_198 ( .A(_abc_42016_n1010), .Y(_abc_42016_n1293) );
  INVX1 INVX1_199 ( .A(_abc_42016_n1295), .Y(_abc_42016_n1296_1) );
  INVX1 INVX1_2 ( .A(_abc_42016_n502), .Y(_abc_42016_n503) );
  INVX1 INVX1_20 ( .A(_abc_42016_n532_1), .Y(_abc_42016_n533) );
  INVX1 INVX1_200 ( .A(rdatahold2_7_), .Y(_abc_42016_n1302) );
  INVX1 INVX1_201 ( .A(_abc_42016_n1310), .Y(_abc_42016_n1311) );
  INVX1 INVX1_202 ( .A(sp_6_), .Y(_abc_42016_n1323) );
  INVX1 INVX1_203 ( .A(_abc_42016_n1325), .Y(_abc_42016_n1326) );
  INVX1 INVX1_204 ( .A(sp_7_), .Y(_abc_42016_n1327_1) );
  INVX1 INVX1_205 ( .A(_abc_42016_n1328), .Y(_abc_42016_n1329_1) );
  INVX1 INVX1_206 ( .A(_abc_42016_n1337_1), .Y(_abc_42016_n1338) );
  INVX1 INVX1_207 ( .A(_abc_42016_n1346), .Y(_abc_42016_n1347) );
  INVX1 INVX1_208 ( .A(_abc_42016_n1348), .Y(_abc_42016_n1350) );
  INVX1 INVX1_209 ( .A(pc_8_), .Y(_abc_42016_n1353) );
  INVX1 INVX1_21 ( .A(_abc_42016_n534_1), .Y(_abc_42016_n535) );
  INVX1 INVX1_210 ( .A(pc_7_), .Y(_abc_42016_n1354) );
  INVX1 INVX1_211 ( .A(pc_6_), .Y(_abc_42016_n1355) );
  INVX1 INVX1_212 ( .A(pc_4_), .Y(_abc_42016_n1356) );
  INVX1 INVX1_213 ( .A(pc_3_), .Y(_abc_42016_n1357) );
  INVX1 INVX1_214 ( .A(_abc_42016_n1359), .Y(_abc_42016_n1360) );
  INVX1 INVX1_215 ( .A(_abc_42016_n1363), .Y(_abc_42016_n1364) );
  INVX1 INVX1_216 ( .A(_abc_42016_n1367), .Y(_abc_42016_n1368) );
  INVX1 INVX1_217 ( .A(_abc_42016_n1369), .Y(_abc_42016_n1370) );
  INVX1 INVX1_218 ( .A(_abc_42016_n1371), .Y(_abc_42016_n1372) );
  INVX1 INVX1_219 ( .A(intcyc), .Y(_abc_42016_n1375) );
  INVX1 INVX1_22 ( .A(opcode_2_), .Y(_abc_42016_n536) );
  INVX1 INVX1_220 ( .A(pc_0_), .Y(_abc_42016_n1381) );
  INVX1 INVX1_221 ( .A(pc_2_), .Y(_abc_42016_n1382) );
  INVX1 INVX1_222 ( .A(pc_1_), .Y(_abc_42016_n1383) );
  INVX1 INVX1_223 ( .A(_abc_42016_n1391), .Y(_abc_42016_n1392) );
  INVX1 INVX1_224 ( .A(_abc_42016_n1395), .Y(_abc_42016_n1396) );
  INVX1 INVX1_225 ( .A(_abc_42016_n1397), .Y(_abc_42016_n1398) );
  INVX1 INVX1_226 ( .A(_abc_42016_n1399), .Y(_abc_42016_n1400) );
  INVX1 INVX1_227 ( .A(_abc_42016_n1404), .Y(_abc_42016_n1405) );
  INVX1 INVX1_228 ( .A(_abc_42016_n1407), .Y(_abc_42016_n1408) );
  INVX1 INVX1_229 ( .A(_abc_42016_n1410_1), .Y(_abc_42016_n1411) );
  INVX1 INVX1_23 ( .A(opcode_1_), .Y(_abc_42016_n537_1) );
  INVX1 INVX1_230 ( .A(wdatahold2_1_), .Y(_abc_42016_n1419) );
  INVX1 INVX1_231 ( .A(pc_9_), .Y(_abc_42016_n1422) );
  INVX1 INVX1_232 ( .A(_abc_42016_n1412), .Y(_abc_42016_n1426) );
  INVX1 INVX1_233 ( .A(regfil_7__1_), .Y(_abc_42016_n1427) );
  INVX1 INVX1_234 ( .A(_abc_42016_n1374), .Y(_abc_42016_n1437) );
  INVX1 INVX1_235 ( .A(_abc_42016_n1378), .Y(_abc_42016_n1438) );
  INVX1 INVX1_236 ( .A(wdatahold2_2_), .Y(_abc_42016_n1445) );
  INVX1 INVX1_237 ( .A(regfil_4__2_), .Y(_abc_42016_n1446) );
  INVX1 INVX1_238 ( .A(pc_10_), .Y(_abc_42016_n1449) );
  INVX1 INVX1_239 ( .A(regfil_7__2_), .Y(_abc_42016_n1454) );
  INVX1 INVX1_24 ( .A(_abc_42016_n538_1), .Y(_abc_42016_n539) );
  INVX1 INVX1_240 ( .A(_abc_42016_n1424), .Y(_abc_42016_n1464) );
  INVX1 INVX1_241 ( .A(wdatahold2_3_), .Y(_abc_42016_n1474) );
  INVX1 INVX1_242 ( .A(pc_11_), .Y(_abc_42016_n1477) );
  INVX1 INVX1_243 ( .A(_abc_42016_n1466), .Y(_abc_42016_n1478) );
  INVX1 INVX1_244 ( .A(_abc_42016_n1485), .Y(_abc_42016_n1486) );
  INVX1 INVX1_245 ( .A(regfil_7__3_), .Y(_abc_42016_n1488) );
  INVX1 INVX1_246 ( .A(wdatahold2_4_), .Y(_abc_42016_n1500) );
  INVX1 INVX1_247 ( .A(pc_12_), .Y(_abc_42016_n1503) );
  INVX1 INVX1_248 ( .A(_abc_42016_n1380), .Y(_abc_42016_n1508) );
  INVX1 INVX1_249 ( .A(_abc_42016_n1510), .Y(_abc_42016_n1511) );
  INVX1 INVX1_25 ( .A(opcode_6_), .Y(_abc_42016_n540) );
  INVX1 INVX1_250 ( .A(_abc_42016_n1512), .Y(_abc_42016_n1513) );
  INVX1 INVX1_251 ( .A(wdatahold2_5_), .Y(_abc_42016_n1526) );
  INVX1 INVX1_252 ( .A(regfil_4__5_), .Y(_abc_42016_n1527) );
  INVX1 INVX1_253 ( .A(pc_13_), .Y(_abc_42016_n1530) );
  INVX1 INVX1_254 ( .A(_abc_42016_n1536), .Y(_abc_42016_n1537) );
  INVX1 INVX1_255 ( .A(_abc_42016_n1545), .Y(_abc_42016_n1546) );
  INVX1 INVX1_256 ( .A(wdatahold2_6_), .Y(_abc_42016_n1553) );
  INVX1 INVX1_257 ( .A(regfil_4__6_), .Y(_abc_42016_n1554) );
  INVX1 INVX1_258 ( .A(pc_14_), .Y(_abc_42016_n1557) );
  INVX1 INVX1_259 ( .A(_abc_42016_n1561), .Y(_abc_42016_n1562) );
  INVX1 INVX1_26 ( .A(_abc_42016_n543), .Y(_abc_42016_n544_1) );
  INVX1 INVX1_260 ( .A(_abc_42016_n1563), .Y(_abc_42016_n1564) );
  INVX1 INVX1_261 ( .A(_abc_42016_n1566), .Y(_abc_42016_n1567) );
  INVX1 INVX1_262 ( .A(pc_15_), .Y(_abc_42016_n1584_1) );
  INVX1 INVX1_263 ( .A(_abc_42016_n1587), .Y(_abc_42016_n1588_1) );
  INVX1 INVX1_264 ( .A(_abc_42016_n1589), .Y(_abc_42016_n1590_1) );
  INVX1 INVX1_265 ( .A(_abc_42016_n550), .Y(_abc_42016_n1603_1) );
  INVX1 INVX1_266 ( .A(_abc_42016_n1623), .Y(_abc_42016_n1624) );
  INVX1 INVX1_267 ( .A(_abc_42016_n1627), .Y(_abc_42016_n1628) );
  INVX1 INVX1_268 ( .A(regfil_2__0_), .Y(_abc_42016_n1631) );
  INVX1 INVX1_269 ( .A(_abc_42016_n1651), .Y(_abc_42016_n1652_1) );
  INVX1 INVX1_27 ( .A(_abc_42016_n545_1), .Y(_abc_42016_n546) );
  INVX1 INVX1_270 ( .A(_abc_42016_n1656), .Y(_abc_42016_n1657) );
  INVX1 INVX1_271 ( .A(_abc_42016_n1666), .Y(_abc_42016_n1667) );
  INVX1 INVX1_272 ( .A(rdatahold_2_), .Y(_abc_42016_n1675) );
  INVX1 INVX1_273 ( .A(_abc_42016_n614), .Y(_abc_42016_n1690_1) );
  INVX1 INVX1_274 ( .A(_abc_42016_n1695), .Y(_abc_42016_n1696) );
  INVX1 INVX1_275 ( .A(_abc_42016_n650), .Y(_abc_42016_n1729_1) );
  INVX1 INVX1_276 ( .A(_abc_42016_n1733), .Y(_abc_42016_n1734) );
  INVX1 INVX1_277 ( .A(_abc_42016_n1737), .Y(_abc_42016_n1738) );
  INVX1 INVX1_278 ( .A(_abc_42016_n617), .Y(_abc_42016_n1751) );
  INVX1 INVX1_279 ( .A(_abc_42016_n1767_1), .Y(_abc_42016_n1783_1) );
  INVX1 INVX1_28 ( .A(_abc_42016_n547), .Y(_abc_42016_n548) );
  INVX1 INVX1_280 ( .A(rdatahold_6_), .Y(_abc_42016_n1793) );
  INVX1 INVX1_281 ( .A(regfil_4__7_), .Y(_abc_42016_n1801_1) );
  INVX1 INVX1_282 ( .A(_abc_42016_n1813), .Y(_abc_42016_n1814) );
  INVX1 INVX1_283 ( .A(regfil_6__5_), .Y(_abc_42016_n1826) );
  INVX1 INVX1_284 ( .A(regfil_6__6_), .Y(_abc_42016_n1829) );
  INVX1 INVX1_285 ( .A(regfil_6__7_), .Y(_abc_42016_n1832) );
  INVX1 INVX1_286 ( .A(_abc_42016_n1843), .Y(_abc_42016_n1844) );
  INVX1 INVX1_287 ( .A(alu_sel_1_), .Y(_abc_42016_n1846) );
  INVX1 INVX1_288 ( .A(_abc_42016_n1841), .Y(_abc_42016_n1848) );
  INVX1 INVX1_289 ( .A(carry), .Y(_abc_42016_n1860) );
  INVX1 INVX1_29 ( .A(regd_0_), .Y(_abc_42016_n551) );
  INVX1 INVX1_290 ( .A(_abc_42016_n1851), .Y(_abc_42016_n1863) );
  INVX1 INVX1_291 ( .A(state_5_), .Y(_abc_42016_n1867) );
  INVX1 INVX1_292 ( .A(_abc_42016_n1869), .Y(_abc_42016_n1870) );
  INVX1 INVX1_293 ( .A(alu_oprb_1_), .Y(_abc_42016_n1878) );
  INVX1 INVX1_294 ( .A(_abc_42016_n1837_1), .Y(_abc_42016_n1879_1) );
  INVX1 INVX1_295 ( .A(alu_oprb_2_), .Y(_abc_42016_n1885) );
  INVX1 INVX1_296 ( .A(alu_oprb_3_), .Y(_abc_42016_n1888_1) );
  INVX1 INVX1_297 ( .A(alu_oprb_4_), .Y(_abc_42016_n1891) );
  INVX1 INVX1_298 ( .A(alu_oprb_5_), .Y(_abc_42016_n1894_1) );
  INVX1 INVX1_299 ( .A(alu_oprb_6_), .Y(_abc_42016_n1897) );
  INVX1 INVX1_3 ( .A(state_1_), .Y(_abc_42016_n504) );
  INVX1 INVX1_30 ( .A(_abc_42016_n555), .Y(_abc_42016_n556) );
  INVX1 INVX1_300 ( .A(_abc_42016_n1909_1), .Y(_abc_42016_n1910) );
  INVX1 INVX1_301 ( .A(_abc_42016_n1911), .Y(_abc_42016_n1912) );
  INVX1 INVX1_302 ( .A(_abc_42016_n1915), .Y(_abc_42016_n1916) );
  INVX1 INVX1_303 ( .A(_abc_42016_n1868), .Y(_abc_42016_n1923) );
  INVX1 INVX1_304 ( .A(_abc_42016_n1925), .Y(_abc_42016_n1926_1) );
  INVX1 INVX1_305 ( .A(_abc_42016_n1927), .Y(_abc_42016_n1933) );
  INVX1 INVX1_306 ( .A(_abc_42016_n1917), .Y(_abc_42016_n1935) );
  INVX1 INVX1_307 ( .A(_abc_42016_n1941), .Y(_abc_42016_n1942) );
  INVX1 INVX1_308 ( .A(_abc_42016_n1967), .Y(_abc_42016_n1968_1) );
  INVX1 INVX1_309 ( .A(regfil_7__4_), .Y(_abc_42016_n1974) );
  INVX1 INVX1_31 ( .A(_abc_42016_n557), .Y(_abc_42016_n558) );
  INVX1 INVX1_310 ( .A(_abc_42016_n2024), .Y(_abc_42016_n2026) );
  INVX1 INVX1_311 ( .A(parity), .Y(_abc_42016_n2029) );
  INVX1 INVX1_312 ( .A(_abc_42016_n2030), .Y(_abc_42016_n2031) );
  INVX1 INVX1_313 ( .A(_abc_42016_n1872), .Y(_abc_42016_n2033) );
  INVX1 INVX1_314 ( .A(_abc_42016_n2034), .Y(_abc_42016_n2035) );
  INVX1 INVX1_315 ( .A(_abc_42016_n2037), .Y(_abc_42016_n2038) );
  INVX1 INVX1_316 ( .A(_abc_42016_n2032), .Y(_abc_42016_n2040) );
  INVX1 INVX1_317 ( .A(_abc_42016_n2041), .Y(_abc_42016_n2042) );
  INVX1 INVX1_318 ( .A(_abc_42016_n2043), .Y(_abc_42016_n2044) );
  INVX1 INVX1_319 ( .A(zero), .Y(_abc_42016_n2050) );
  INVX1 INVX1_32 ( .A(_abc_42016_n559), .Y(_abc_42016_n560) );
  INVX1 INVX1_320 ( .A(sign), .Y(_abc_42016_n2056) );
  INVX1 INVX1_321 ( .A(alu_sout), .Y(_abc_42016_n2058) );
  INVX1 INVX1_322 ( .A(auxcar), .Y(_abc_42016_n2064) );
  INVX1 INVX1_323 ( .A(_abc_42016_n2070), .Y(_abc_42016_n2072) );
  INVX1 INVX1_324 ( .A(_abc_42016_n2078), .Y(_abc_42016_n2079) );
  INVX1 INVX1_325 ( .A(_abc_42016_n1463), .Y(_abc_42016_n2084) );
  INVX1 INVX1_326 ( .A(_abc_42016_n1462), .Y(_abc_42016_n2085) );
  INVX1 INVX1_327 ( .A(_abc_42016_n2086), .Y(_abc_42016_n2087) );
  INVX1 INVX1_328 ( .A(_abc_42016_n2093), .Y(_abc_42016_n2094) );
  INVX1 INVX1_329 ( .A(sp_15_), .Y(_abc_42016_n2101) );
  INVX1 INVX1_33 ( .A(_abc_42016_n561), .Y(_abc_42016_n562) );
  INVX1 INVX1_330 ( .A(sp_14_), .Y(_abc_42016_n2103) );
  INVX1 INVX1_331 ( .A(_abc_42016_n2107), .Y(_abc_42016_n2108) );
  INVX1 INVX1_332 ( .A(sp_13_), .Y(_abc_42016_n2109_1) );
  INVX1 INVX1_333 ( .A(_abc_42016_n2110_1), .Y(_abc_42016_n2111) );
  INVX1 INVX1_334 ( .A(sp_12_), .Y(_abc_42016_n2113) );
  INVX1 INVX1_335 ( .A(_abc_42016_n2116_1), .Y(_abc_42016_n2117) );
  INVX1 INVX1_336 ( .A(sp_11_), .Y(_abc_42016_n2118) );
  INVX1 INVX1_337 ( .A(_abc_42016_n2119_1), .Y(_abc_42016_n2120_1) );
  INVX1 INVX1_338 ( .A(sp_10_), .Y(_abc_42016_n2122) );
  INVX1 INVX1_339 ( .A(_abc_42016_n2125), .Y(_abc_42016_n2126) );
  INVX1 INVX1_34 ( .A(opcode_0_), .Y(_abc_42016_n563) );
  INVX1 INVX1_340 ( .A(sp_9_), .Y(_abc_42016_n2127_1) );
  INVX1 INVX1_341 ( .A(_abc_42016_n2128_1), .Y(_abc_42016_n2129) );
  INVX1 INVX1_342 ( .A(sp_8_), .Y(_abc_42016_n2131_1) );
  INVX1 INVX1_343 ( .A(_abc_42016_n2151_1), .Y(_abc_42016_n2152) );
  INVX1 INVX1_344 ( .A(_abc_42016_n2155), .Y(_abc_42016_n2156) );
  INVX1 INVX1_345 ( .A(_abc_42016_n2157), .Y(_abc_42016_n2158) );
  INVX1 INVX1_346 ( .A(_abc_42016_n2163), .Y(_abc_42016_n2164) );
  INVX1 INVX1_347 ( .A(_abc_42016_n1317), .Y(_abc_42016_n2166) );
  INVX1 INVX1_348 ( .A(_abc_42016_n1316), .Y(_abc_42016_n2168) );
  INVX1 INVX1_349 ( .A(_abc_42016_n2184), .Y(_abc_42016_n2185) );
  INVX1 INVX1_35 ( .A(_abc_42016_n564), .Y(_abc_42016_n565) );
  INVX1 INVX1_350 ( .A(_abc_42016_n2189), .Y(_abc_42016_n2190) );
  INVX1 INVX1_351 ( .A(_abc_42016_n2195), .Y(_abc_42016_n2196) );
  INVX1 INVX1_352 ( .A(_abc_42016_n1306), .Y(_abc_42016_n2198) );
  INVX1 INVX1_353 ( .A(_abc_42016_n1307), .Y(_abc_42016_n2201) );
  INVX1 INVX1_354 ( .A(_abc_42016_n2080), .Y(_abc_42016_n2217) );
  INVX1 INVX1_355 ( .A(\data[0] ), .Y(_abc_42016_n2225) );
  INVX1 INVX1_356 ( .A(_abc_42016_n2228), .Y(_abc_42016_n2229) );
  INVX1 INVX1_357 ( .A(_abc_42016_n2226), .Y(_abc_42016_n2231) );
  INVX1 INVX1_358 ( .A(\data[1] ), .Y(_abc_42016_n2234) );
  INVX1 INVX1_359 ( .A(\data[2] ), .Y(_abc_42016_n2237) );
  INVX1 INVX1_36 ( .A(opcode_3_), .Y(_abc_42016_n566) );
  INVX1 INVX1_360 ( .A(\data[3] ), .Y(_abc_42016_n2240) );
  INVX1 INVX1_361 ( .A(\data[4] ), .Y(_abc_42016_n2243) );
  INVX1 INVX1_362 ( .A(\data[5] ), .Y(_abc_42016_n2246) );
  INVX1 INVX1_363 ( .A(\data[6] ), .Y(_abc_42016_n2248) );
  INVX1 INVX1_364 ( .A(\data[7] ), .Y(_abc_42016_n2250) );
  INVX1 INVX1_365 ( .A(_abc_42016_n2253), .Y(_abc_42016_n2254) );
  INVX1 INVX1_366 ( .A(statesel_0_), .Y(_abc_42016_n2259) );
  INVX1 INVX1_367 ( .A(_abc_42016_n2269), .Y(_abc_42016_n2270_1) );
  INVX1 INVX1_368 ( .A(_abc_42016_n2271_1), .Y(_abc_42016_n2272) );
  INVX1 INVX1_369 ( .A(_abc_42016_n2275), .Y(_abc_42016_n2276) );
  INVX1 INVX1_37 ( .A(_abc_42016_n567), .Y(_abc_42016_n568) );
  INVX1 INVX1_370 ( .A(_abc_42016_n2279), .Y(_abc_42016_n2280) );
  INVX1 INVX1_371 ( .A(_abc_42016_n2283), .Y(_abc_42016_n2284) );
  INVX1 INVX1_372 ( .A(_abc_42016_n2281), .Y(_abc_42016_n2291) );
  INVX1 INVX1_373 ( .A(_abc_42016_n542), .Y(_abc_42016_n2297_1) );
  INVX1 INVX1_374 ( .A(_abc_42016_n2298), .Y(_abc_42016_n2299) );
  INVX1 INVX1_375 ( .A(_abc_42016_n2301), .Y(_abc_42016_n2302) );
  INVX1 INVX1_376 ( .A(_abc_42016_n2303), .Y(_abc_42016_n2304) );
  INVX1 INVX1_377 ( .A(_abc_42016_n2309), .Y(_abc_42016_n2310) );
  INVX1 INVX1_378 ( .A(_abc_42016_n2311), .Y(_abc_42016_n2312) );
  INVX1 INVX1_379 ( .A(_abc_42016_n2314), .Y(_abc_42016_n2315) );
  INVX1 INVX1_38 ( .A(_abc_42016_n571), .Y(_abc_42016_n572) );
  INVX1 INVX1_380 ( .A(_abc_42016_n2320), .Y(_abc_42016_n2321) );
  INVX1 INVX1_381 ( .A(_abc_42016_n2322), .Y(_abc_42016_n2323_1) );
  INVX1 INVX1_382 ( .A(_abc_42016_n2324_1), .Y(_abc_42016_n2325) );
  INVX1 INVX1_383 ( .A(_abc_42016_n2326), .Y(_abc_42016_n2327) );
  INVX1 INVX1_384 ( .A(_abc_42016_n2328), .Y(_abc_42016_n2329) );
  INVX1 INVX1_385 ( .A(_abc_42016_n2334), .Y(_abc_42016_n2335) );
  INVX1 INVX1_386 ( .A(_abc_42016_n2278), .Y(_abc_42016_n2337) );
  INVX1 INVX1_387 ( .A(waitr), .Y(_abc_42016_n2338) );
  INVX1 INVX1_388 ( .A(_abc_42016_n2339), .Y(_abc_42016_n2340) );
  INVX1 INVX1_389 ( .A(statesel_1_), .Y(_abc_42016_n2344) );
  INVX1 INVX1_39 ( .A(_abc_42016_n575), .Y(_abc_42016_n576_1) );
  INVX1 INVX1_390 ( .A(_abc_42016_n541), .Y(_abc_42016_n2355) );
  INVX1 INVX1_391 ( .A(_abc_42016_n2358), .Y(_abc_42016_n2359) );
  INVX1 INVX1_392 ( .A(statesel_2_), .Y(_abc_42016_n2369) );
  INVX1 INVX1_393 ( .A(_abc_42016_n2372_1), .Y(_abc_42016_n2373_1) );
  INVX1 INVX1_394 ( .A(_abc_42016_n2347_1), .Y(_abc_42016_n2376) );
  INVX1 INVX1_395 ( .A(_abc_42016_n2378), .Y(_abc_42016_n2379) );
  INVX1 INVX1_396 ( .A(_abc_42016_n2336), .Y(_abc_42016_n2385) );
  INVX1 INVX1_397 ( .A(statesel_3_), .Y(_abc_42016_n2394_1) );
  INVX1 INVX1_398 ( .A(_abc_42016_n2289), .Y(_abc_42016_n2395) );
  INVX1 INVX1_399 ( .A(_abc_42016_n2387), .Y(_abc_42016_n2407) );
  INVX1 INVX1_4 ( .A(state_0_), .Y(_abc_42016_n505) );
  INVX1 INVX1_40 ( .A(_abc_42016_n577), .Y(_abc_42016_n578) );
  INVX1 INVX1_400 ( .A(_abc_42016_n2408_1), .Y(_abc_42016_n2409) );
  INVX1 INVX1_401 ( .A(_abc_42016_n2411_1), .Y(_abc_42016_n2412) );
  INVX1 INVX1_402 ( .A(statesel_4_), .Y(_abc_42016_n2417_1) );
  INVX1 INVX1_403 ( .A(_abc_42016_n2285), .Y(_abc_42016_n2423_1) );
  INVX1 INVX1_404 ( .A(_abc_42016_n2424), .Y(_abc_42016_n2425) );
  INVX1 INVX1_405 ( .A(_abc_42016_n2427), .Y(_abc_42016_n2428) );
  INVX1 INVX1_406 ( .A(_abc_42016_n2429_1), .Y(_abc_42016_n2430) );
  INVX1 INVX1_407 ( .A(_abc_42016_n2436), .Y(_abc_42016_n2437) );
  INVX1 INVX1_408 ( .A(_abc_42016_n2438_1), .Y(_abc_42016_n2440) );
  INVX1 INVX1_409 ( .A(statesel_5_), .Y(_abc_42016_n2446) );
  INVX1 INVX1_41 ( .A(_abc_42016_n580), .Y(_abc_42016_n581_1) );
  INVX1 INVX1_410 ( .A(_abc_42016_n2450_1), .Y(_abc_42016_n2451) );
  INVX1 INVX1_411 ( .A(rdatahold_4_), .Y(_abc_42016_n2471) );
  INVX1 INVX1_412 ( .A(rdatahold_7_), .Y(_abc_42016_n2478) );
  INVX1 INVX1_413 ( .A(wdatahold_0_), .Y(_abc_42016_n2496) );
  INVX1 INVX1_414 ( .A(_abc_42016_n2499), .Y(_abc_42016_n2500) );
  INVX1 INVX1_415 ( .A(_abc_42016_n2497), .Y(_abc_42016_n2519) );
  INVX1 INVX1_416 ( .A(_abc_42016_n2536), .Y(_abc_42016_n2537) );
  INVX1 INVX1_417 ( .A(_abc_42016_n2529), .Y(_abc_42016_n2543) );
  INVX1 INVX1_418 ( .A(wdatahold_1_), .Y(_abc_42016_n2548_1) );
  INVX1 INVX1_419 ( .A(wdatahold_2_), .Y(_abc_42016_n2555) );
  INVX1 INVX1_42 ( .A(_abc_42016_n582_1), .Y(_abc_42016_n583) );
  INVX1 INVX1_420 ( .A(_abc_42016_n2561), .Y(_abc_42016_n2562) );
  INVX1 INVX1_421 ( .A(_abc_42016_n1358), .Y(_abc_42016_n2571) );
  INVX1 INVX1_422 ( .A(wdatahold_6_), .Y(_abc_42016_n2583) );
  INVX1 INVX1_423 ( .A(wdatahold_3_), .Y(_abc_42016_n2587) );
  INVX1 INVX1_424 ( .A(_abc_42016_n2589), .Y(_abc_42016_n2590) );
  INVX1 INVX1_425 ( .A(_abc_42016_n2597), .Y(_abc_42016_n2598) );
  INVX1 INVX1_426 ( .A(_abc_42016_n2593), .Y(_abc_42016_n2606) );
  INVX1 INVX1_427 ( .A(alu_res_3_), .Y(_abc_42016_n2612) );
  INVX1 INVX1_428 ( .A(_abc_42016_n2518_1), .Y(_abc_42016_n2613) );
  INVX1 INVX1_429 ( .A(_abc_42016_n2267), .Y(_abc_42016_n2614) );
  INVX1 INVX1_43 ( .A(_abc_42016_n584_1), .Y(_abc_42016_n585) );
  INVX1 INVX1_430 ( .A(wdatahold_4_), .Y(_abc_42016_n2619) );
  INVX1 INVX1_431 ( .A(_abc_42016_n1245), .Y(_abc_42016_n2624) );
  INVX1 INVX1_432 ( .A(_abc_42016_n1386_1), .Y(_abc_42016_n2630) );
  INVX1 INVX1_433 ( .A(_abc_42016_n1361), .Y(_abc_42016_n2633) );
  INVX1 INVX1_434 ( .A(_abc_42016_n2512), .Y(_abc_42016_n2639_1) );
  INVX1 INVX1_435 ( .A(wdatahold_5_), .Y(_abc_42016_n2648) );
  INVX1 INVX1_436 ( .A(pc_5_), .Y(_abc_42016_n2649) );
  INVX1 INVX1_437 ( .A(_abc_42016_n1388), .Y(_abc_42016_n2674) );
  INVX1 INVX1_438 ( .A(_abc_42016_n2678), .Y(_abc_42016_n2679) );
  INVX1 INVX1_439 ( .A(_abc_42016_n2684), .Y(_abc_42016_n2685) );
  INVX1 INVX1_44 ( .A(regd_1_), .Y(_abc_42016_n589) );
  INVX1 INVX1_440 ( .A(_abc_42016_n2687), .Y(_abc_42016_n2688) );
  INVX1 INVX1_441 ( .A(alu_res_6_), .Y(_abc_42016_n2695) );
  INVX1 INVX1_442 ( .A(_abc_42016_n2539), .Y(_abc_42016_n2700) );
  INVX1 INVX1_443 ( .A(wdatahold_7_), .Y(_abc_42016_n2709) );
  INVX1 INVX1_444 ( .A(raddrhold_0_), .Y(_abc_42016_n2731) );
  INVX1 INVX1_445 ( .A(_abc_42016_n2732), .Y(_abc_42016_n2733) );
  INVX1 INVX1_446 ( .A(_abc_42016_n2735), .Y(_abc_42016_n2736) );
  INVX1 INVX1_447 ( .A(_abc_42016_n2737), .Y(_abc_42016_n2738) );
  INVX1 INVX1_448 ( .A(_abc_42016_n2739), .Y(_abc_42016_n2740) );
  INVX1 INVX1_449 ( .A(_abc_42016_n2746), .Y(_abc_42016_n2747_1) );
  INVX1 INVX1_45 ( .A(_abc_42016_n592_1), .Y(_abc_42016_n593) );
  INVX1 INVX1_450 ( .A(sp_0_), .Y(_abc_42016_n2758) );
  INVX1 INVX1_451 ( .A(_abc_42016_n2743), .Y(_abc_42016_n2759) );
  INVX1 INVX1_452 ( .A(raddrhold_1_), .Y(_abc_42016_n2765) );
  INVX1 INVX1_453 ( .A(_abc_42016_n2754), .Y(_abc_42016_n2768_1) );
  INVX1 INVX1_454 ( .A(_abc_42016_n2526), .Y(_abc_42016_n2769) );
  INVX1 INVX1_455 ( .A(sp_1_), .Y(_abc_42016_n2775) );
  INVX1 INVX1_456 ( .A(_abc_42016_n2777), .Y(_abc_42016_n2778) );
  INVX1 INVX1_457 ( .A(raddrhold_2_), .Y(_abc_42016_n2786) );
  INVX1 INVX1_458 ( .A(_abc_42016_n2787), .Y(_abc_42016_n2788_1) );
  INVX1 INVX1_459 ( .A(raddrhold_3_), .Y(_abc_42016_n2803) );
  INVX1 INVX1_46 ( .A(regd_2_), .Y(_abc_42016_n594_1) );
  INVX1 INVX1_460 ( .A(_abc_42016_n2810_1), .Y(_abc_42016_n2811_1) );
  INVX1 INVX1_461 ( .A(sp_3_), .Y(_abc_42016_n2813) );
  INVX1 INVX1_462 ( .A(raddrhold_4_), .Y(_abc_42016_n2820) );
  INVX1 INVX1_463 ( .A(_abc_42016_n2828), .Y(_abc_42016_n2829) );
  INVX1 INVX1_464 ( .A(raddrhold_5_), .Y(_abc_42016_n2836) );
  INVX1 INVX1_465 ( .A(raddrhold_6_), .Y(_abc_42016_n2852) );
  INVX1 INVX1_466 ( .A(raddrhold_7_), .Y(_abc_42016_n2869) );
  INVX1 INVX1_467 ( .A(_abc_42016_n2716), .Y(_abc_42016_n2872) );
  INVX1 INVX1_468 ( .A(_abc_42016_n2881), .Y(_abc_42016_n2882) );
  INVX1 INVX1_469 ( .A(raddrhold_8_), .Y(_abc_42016_n2887) );
  INVX1 INVX1_47 ( .A(_abc_42016_n598_1), .Y(_abc_42016_n599) );
  INVX1 INVX1_470 ( .A(_abc_42016_n2908), .Y(_abc_42016_n2909) );
  INVX1 INVX1_471 ( .A(_abc_42016_n2912), .Y(_abc_42016_n2913) );
  INVX1 INVX1_472 ( .A(raddrhold_10_), .Y(_abc_42016_n2920) );
  INVX1 INVX1_473 ( .A(_abc_42016_n2745), .Y(_abc_42016_n2929) );
  INVX1 INVX1_474 ( .A(_abc_42016_n2934), .Y(_abc_42016_n2935) );
  INVX1 INVX1_475 ( .A(raddrhold_11_), .Y(_abc_42016_n2942) );
  INVX1 INVX1_476 ( .A(raddrhold_12_), .Y(_abc_42016_n2956) );
  INVX1 INVX1_477 ( .A(raddrhold_13_), .Y(_abc_42016_n2972) );
  INVX1 INVX1_478 ( .A(_abc_42016_n1533), .Y(_abc_42016_n2973) );
  INVX1 INVX1_479 ( .A(_abc_42016_n2984), .Y(_abc_42016_n2985) );
  INVX1 INVX1_48 ( .A(_abc_42016_n600), .Y(_abc_42016_n601) );
  INVX1 INVX1_480 ( .A(raddrhold_14_), .Y(_abc_42016_n2990_1) );
  INVX1 INVX1_481 ( .A(_abc_42016_n2998), .Y(_abc_42016_n2999) );
  INVX1 INVX1_482 ( .A(_abc_42016_n3003), .Y(_abc_42016_n3004) );
  INVX1 INVX1_483 ( .A(raddrhold_15_), .Y(_abc_42016_n3009) );
  INVX1 INVX1_484 ( .A(_abc_42016_n3015_1), .Y(_abc_42016_n3016) );
  INVX1 INVX1_485 ( .A(waddrhold_0_), .Y(_abc_42016_n3028) );
  INVX1 INVX1_486 ( .A(_abc_42016_n3033), .Y(_abc_42016_n3034) );
  INVX1 INVX1_487 ( .A(_abc_42016_n2261), .Y(_abc_42016_n3045) );
  INVX1 INVX1_488 ( .A(waddrhold_1_), .Y(_abc_42016_n3050) );
  INVX1 INVX1_489 ( .A(_abc_42016_n2089), .Y(_abc_42016_n3052) );
  INVX1 INVX1_49 ( .A(rdatahold_0_), .Y(_abc_42016_n602) );
  INVX1 INVX1_490 ( .A(rdatahold2_1_), .Y(_abc_42016_n3070) );
  INVX1 INVX1_491 ( .A(_abc_42016_n3031), .Y(_abc_42016_n3072) );
  INVX1 INVX1_492 ( .A(waddrhold_2_), .Y(_abc_42016_n3078_1) );
  INVX1 INVX1_493 ( .A(_abc_42016_n3079), .Y(_abc_42016_n3080_1) );
  INVX1 INVX1_494 ( .A(_abc_42016_n3082), .Y(_abc_42016_n3083) );
  INVX1 INVX1_495 ( .A(_abc_42016_n2293), .Y(_abc_42016_n3090) );
  INVX1 INVX1_496 ( .A(_abc_42016_n3099), .Y(_abc_42016_n3100) );
  INVX1 INVX1_497 ( .A(waddrhold_3_), .Y(_abc_42016_n3105_1) );
  INVX1 INVX1_498 ( .A(_abc_42016_n3097), .Y(_abc_42016_n3119) );
  INVX1 INVX1_499 ( .A(_abc_42016_n3120), .Y(_abc_42016_n3121) );
  INVX1 INVX1_5 ( .A(_abc_42016_n506), .Y(_abc_42016_n507) );
  INVX1 INVX1_50 ( .A(_abc_42016_n569), .Y(_abc_42016_n603) );
  INVX1 INVX1_500 ( .A(waddrhold_4_), .Y(_abc_42016_n3128) );
  INVX1 INVX1_501 ( .A(_abc_42016_n3056), .Y(_abc_42016_n3130) );
  INVX1 INVX1_502 ( .A(_abc_42016_n3133), .Y(_abc_42016_n3134) );
  INVX1 INVX1_503 ( .A(_abc_42016_n3107), .Y(_abc_42016_n3146) );
  INVX1 INVX1_504 ( .A(waddrhold_5_), .Y(_abc_42016_n3153) );
  INVX1 INVX1_505 ( .A(waddrhold_6_), .Y(_abc_42016_n3175) );
  INVX1 INVX1_506 ( .A(_abc_42016_n3177), .Y(_abc_42016_n3178) );
  INVX1 INVX1_507 ( .A(_abc_42016_n3179), .Y(_abc_42016_n3180) );
  INVX1 INVX1_508 ( .A(_abc_42016_n3194), .Y(_abc_42016_n3195_1) );
  INVX1 INVX1_509 ( .A(waddrhold_7_), .Y(_abc_42016_n3201) );
  INVX1 INVX1_51 ( .A(_abc_42016_n570), .Y(_abc_42016_n604_1) );
  INVX1 INVX1_510 ( .A(_abc_42016_n3216), .Y(_abc_42016_n3217_1) );
  INVX1 INVX1_511 ( .A(waddrhold_8_), .Y(_abc_42016_n3223) );
  INVX1 INVX1_512 ( .A(_abc_42016_n3224), .Y(_abc_42016_n3225) );
  INVX1 INVX1_513 ( .A(_abc_42016_n3238), .Y(_abc_42016_n3239) );
  INVX1 INVX1_514 ( .A(waddrhold_9_), .Y(_abc_42016_n3245_1) );
  INVX1 INVX1_515 ( .A(waddrhold_10_), .Y(_abc_42016_n3268) );
  INVX1 INVX1_516 ( .A(waddrhold_11_), .Y(_abc_42016_n3291) );
  INVX1 INVX1_517 ( .A(_abc_42016_n3248), .Y(_abc_42016_n3293) );
  INVX1 INVX1_518 ( .A(_abc_42016_n3295_1), .Y(_abc_42016_n3296_1) );
  INVX1 INVX1_519 ( .A(_abc_42016_n3297), .Y(_abc_42016_n3298) );
  INVX1 INVX1_52 ( .A(_abc_42016_n606), .Y(_abc_42016_n607) );
  INVX1 INVX1_520 ( .A(_abc_42016_n3309), .Y(_abc_42016_n3310) );
  INVX1 INVX1_521 ( .A(waddrhold_12_), .Y(_abc_42016_n3316) );
  INVX1 INVX1_522 ( .A(waddrhold_13_), .Y(_abc_42016_n3337) );
  INVX1 INVX1_523 ( .A(_abc_42016_n3339), .Y(_abc_42016_n3340) );
  INVX1 INVX1_524 ( .A(waddrhold_14_), .Y(_abc_42016_n3361) );
  INVX1 INVX1_525 ( .A(_abc_42016_n3362), .Y(_abc_42016_n3363) );
  INVX1 INVX1_526 ( .A(_abc_42016_n3365), .Y(_abc_42016_n3366) );
  INVX1 INVX1_527 ( .A(_abc_42016_n3381), .Y(_abc_42016_n3382) );
  INVX1 INVX1_528 ( .A(waddrhold_15_), .Y(_abc_42016_n3388) );
  INVX1 INVX1_529 ( .A(_abc_42016_n3407), .Y(_abc_42016_n3408) );
  INVX1 INVX1_53 ( .A(regfil_0__0_), .Y(_abc_42016_n608) );
  INVX1 INVX1_530 ( .A(_abc_42016_n3409), .Y(_abc_42016_n3418) );
  INVX1 INVX1_531 ( .A(_abc_42016_n3429), .Y(_abc_42016_n3430) );
  INVX1 INVX1_532 ( .A(_abc_42016_n3431), .Y(_abc_42016_n3433) );
  INVX1 INVX1_533 ( .A(_abc_42016_n2255), .Y(_abc_42016_n3453) );
  INVX1 INVX1_534 ( .A(_abc_42016_n3458), .Y(_abc_42016_n3459) );
  INVX1 INVX1_535 ( .A(_abc_42016_n3460), .Y(_abc_42016_n3466) );
  INVX1 INVX1_536 ( .A(_abc_42016_n3469), .Y(_abc_42016_n3470_1) );
  INVX1 INVX1_537 ( .A(_abc_42016_n3474), .Y(_abc_42016_n3475) );
  INVX1 INVX1_538 ( .A(_abc_42016_n3476_1), .Y(_abc_42016_n3477) );
  INVX1 INVX1_539 ( .A(_abc_42016_n2256), .Y(_abc_42016_n3490) );
  INVX1 INVX1_54 ( .A(regfil_1__6_), .Y(_abc_42016_n609) );
  INVX1 INVX1_540 ( .A(_abc_42016_n1344), .Y(_abc_42016_n3497_1) );
  INVX1 INVX1_541 ( .A(_abc_42016_n3462), .Y(_abc_42016_n3501) );
  INVX1 INVX1_542 ( .A(_abc_42016_n3098), .Y(_abc_42016_n3517) );
  INVX1 INVX1_543 ( .A(_abc_42016_n3519), .Y(_abc_42016_n3520) );
  INVX1 INVX1_544 ( .A(_abc_42016_n3503), .Y(_abc_42016_n3527) );
  INVX1 INVX1_545 ( .A(_abc_42016_n3533), .Y(_abc_42016_n3534) );
  INVX1 INVX1_546 ( .A(_abc_42016_n3555), .Y(_abc_42016_n3556) );
  INVX1 INVX1_547 ( .A(_abc_42016_n3568), .Y(_abc_42016_n3569) );
  INVX1 INVX1_548 ( .A(_abc_42016_n3571), .Y(_abc_42016_n3572) );
  INVX1 INVX1_549 ( .A(_abc_42016_n3502), .Y(_abc_42016_n3575) );
  INVX1 INVX1_55 ( .A(regfil_1__4_), .Y(_abc_42016_n610) );
  INVX1 INVX1_550 ( .A(rdatahold2_5_), .Y(_abc_42016_n3577) );
  INVX1 INVX1_551 ( .A(_abc_42016_n3554), .Y(_abc_42016_n3581) );
  INVX1 INVX1_552 ( .A(_abc_42016_n3589), .Y(_abc_42016_n3590) );
  INVX1 INVX1_553 ( .A(_abc_42016_n3606_1), .Y(_abc_42016_n3607) );
  INVX1 INVX1_554 ( .A(_abc_42016_n3614), .Y(_abc_42016_n3632) );
  INVX1 INVX1_555 ( .A(_abc_42016_n3652), .Y(_abc_42016_n3653) );
  INVX1 INVX1_556 ( .A(_abc_42016_n3658), .Y(_abc_42016_n3659) );
  INVX1 INVX1_557 ( .A(_abc_42016_n3693), .Y(_abc_42016_n3694) );
  INVX1 INVX1_558 ( .A(_abc_42016_n3713_1), .Y(_abc_42016_n3714) );
  INVX1 INVX1_559 ( .A(_abc_42016_n3725), .Y(_abc_42016_n3726) );
  INVX1 INVX1_56 ( .A(regfil_1__2_), .Y(_abc_42016_n611) );
  INVX1 INVX1_560 ( .A(_abc_42016_n3321), .Y(_abc_42016_n3732) );
  INVX1 INVX1_561 ( .A(_abc_42016_n3806), .Y(_abc_42016_n3807) );
  INVX1 INVX1_562 ( .A(_abc_42016_n2133), .Y(_abc_42016_n3813) );
  INVX1 INVX1_563 ( .A(_abc_42016_n2135_1), .Y(_abc_42016_n3814) );
  INVX1 INVX1_564 ( .A(_abc_42016_n2170), .Y(_abc_42016_n3817_1) );
  INVX1 INVX1_565 ( .A(_abc_42016_n2200), .Y(_abc_42016_n3818) );
  INVX1 INVX1_566 ( .A(_abc_42016_n2202), .Y(_abc_42016_n3819) );
  INVX1 INVX1_567 ( .A(_abc_42016_n3800), .Y(_abc_42016_n3834) );
  INVX1 INVX1_568 ( .A(_abc_42016_n3841), .Y(_abc_42016_n3842) );
  INVX1 INVX1_569 ( .A(_abc_42016_n3867), .Y(_abc_42016_n3868) );
  INVX1 INVX1_57 ( .A(_abc_42016_n619), .Y(_abc_42016_n620) );
  INVX1 INVX1_570 ( .A(_abc_42016_n2124_1), .Y(_abc_42016_n3874) );
  INVX1 INVX1_571 ( .A(_abc_42016_n2137), .Y(_abc_42016_n3875) );
  INVX1 INVX1_572 ( .A(_abc_42016_n2205), .Y(_abc_42016_n3878) );
  INVX1 INVX1_573 ( .A(_abc_42016_n2161), .Y(_abc_42016_n3881) );
  INVX1 INVX1_574 ( .A(_abc_42016_n3901), .Y(_abc_42016_n3902) );
  INVX1 INVX1_575 ( .A(_abc_42016_n3910), .Y(_abc_42016_n3912) );
  INVX1 INVX1_576 ( .A(_abc_42016_n2115_1), .Y(_abc_42016_n3929) );
  INVX1 INVX1_577 ( .A(_abc_42016_n2139_1), .Y(_abc_42016_n3930) );
  INVX1 INVX1_578 ( .A(_abc_42016_n3947), .Y(_abc_42016_n3948) );
  INVX1 INVX1_579 ( .A(_abc_42016_n2182), .Y(_abc_42016_n3990) );
  INVX1 INVX1_58 ( .A(_abc_42016_n528_1), .Y(_abc_42016_n624) );
  INVX1 INVX1_580 ( .A(_abc_42016_n2142), .Y(_abc_42016_n3994) );
  INVX1 INVX1_581 ( .A(_abc_42016_n1096), .Y(_abc_42016_n4013) );
  INVX1 INVX1_582 ( .A(_abc_42016_n4016), .Y(_abc_42016_n4017) );
  INVX1 INVX1_583 ( .A(_abc_42016_n4021), .Y(_abc_42016_n4023) );
  INVX1 INVX1_584 ( .A(_abc_42016_n4029), .Y(_abc_42016_n4030) );
  INVX1 INVX1_585 ( .A(_abc_42016_n4045), .Y(_abc_42016_n4046) );
  INVX1 INVX1_586 ( .A(_abc_42016_n4047), .Y(_abc_42016_n4048) );
  INVX1 INVX1_587 ( .A(_abc_42016_n4050), .Y(_abc_42016_n4051) );
  INVX1 INVX1_588 ( .A(_abc_42016_n4055), .Y(_abc_42016_n4056) );
  INVX1 INVX1_589 ( .A(_abc_42016_n4059), .Y(_abc_42016_n4060) );
  INVX1 INVX1_59 ( .A(_abc_42016_n625), .Y(_abc_42016_n626) );
  INVX1 INVX1_590 ( .A(_abc_42016_n4063), .Y(_abc_42016_n4064) );
  INVX1 INVX1_591 ( .A(_abc_42016_n2066), .Y(_abc_42016_n4066) );
  INVX1 INVX1_592 ( .A(_abc_42016_n4068), .Y(_abc_42016_n4069) );
  INVX1 INVX1_593 ( .A(_abc_42016_n4076), .Y(_abc_42016_n4077) );
  INVX1 INVX1_594 ( .A(_abc_42016_n4078), .Y(_abc_42016_n4079) );
  INVX1 INVX1_595 ( .A(_abc_42016_n4086), .Y(_abc_42016_n4087) );
  INVX1 INVX1_596 ( .A(_abc_42016_n4088), .Y(_abc_42016_n4090) );
  INVX1 INVX1_597 ( .A(_abc_42016_n4089), .Y(_abc_42016_n4091) );
  INVX1 INVX1_598 ( .A(_abc_42016_n4128), .Y(_abc_42016_n4129) );
  INVX1 INVX1_599 ( .A(_abc_42016_n4131), .Y(_abc_42016_n4132) );
  INVX1 INVX1_6 ( .A(_abc_42016_n508), .Y(_abc_42016_n509) );
  INVX1 INVX1_60 ( .A(regfil_7__0_), .Y(_abc_42016_n628) );
  INVX1 INVX1_600 ( .A(_abc_42016_n4113), .Y(_abc_42016_n4145) );
  INVX1 INVX1_601 ( .A(_abc_42016_n4146), .Y(_abc_42016_n4156) );
  INVX1 INVX1_602 ( .A(_abc_42016_n4157), .Y(_abc_42016_n4158) );
  INVX1 INVX1_603 ( .A(_abc_42016_n2651), .Y(_abc_42016_n4185) );
  INVX1 INVX1_604 ( .A(_abc_42016_n4130), .Y(_abc_42016_n4210) );
  INVX1 INVX1_605 ( .A(_abc_42016_n1393), .Y(_abc_42016_n4229) );
  INVX1 INVX1_606 ( .A(_abc_42016_n1425), .Y(_abc_42016_n4242) );
  INVX1 INVX1_607 ( .A(_abc_42016_n1452), .Y(_abc_42016_n4249) );
  INVX1 INVX1_608 ( .A(_abc_42016_n1481), .Y(_abc_42016_n4261) );
  INVX1 INVX1_609 ( .A(_abc_42016_n4263), .Y(_abc_42016_n4264) );
  INVX1 INVX1_61 ( .A(regfil_4__0_), .Y(_abc_42016_n629) );
  INVX1 INVX1_610 ( .A(_abc_42016_n1585), .Y(_abc_42016_n4299) );
  INVX1 INVX1_611 ( .A(_abc_42016_n4325), .Y(_abc_42016_n4326) );
  INVX1 INVX1_612 ( .A(_abc_42016_n4349), .Y(_abc_42016_n4350) );
  INVX1 INVX1_613 ( .A(_abc_42016_n4340), .Y(_abc_42016_n4367) );
  INVX1 INVX1_614 ( .A(_abc_42016_n4071), .Y(_abc_42016_n4369) );
  INVX1 INVX1_615 ( .A(_abc_42016_n4378), .Y(_abc_42016_n4379) );
  INVX1 INVX1_616 ( .A(_abc_42016_n4362), .Y(_abc_42016_n4392) );
  INVX1 INVX1_617 ( .A(_abc_42016_n4399), .Y(_abc_42016_n4400) );
  INVX1 INVX1_618 ( .A(_abc_42016_n4438), .Y(_abc_42016_n4439) );
  INVX1 INVX1_619 ( .A(_abc_42016_n4459), .Y(_abc_42016_n4460) );
  INVX1 INVX1_62 ( .A(regfil_3__0_), .Y(_abc_42016_n634) );
  INVX1 INVX1_620 ( .A(_auto_iopadmap_cc_313_execute_46257_0_), .Y(_abc_42016_n4466) );
  INVX1 INVX1_621 ( .A(_abc_42016_n3410), .Y(_abc_42016_n4468) );
  INVX1 INVX1_622 ( .A(_abc_42016_n4469), .Y(_abc_42016_n4472) );
  INVX1 INVX1_623 ( .A(_auto_iopadmap_cc_313_execute_46257_1_), .Y(_abc_42016_n4478) );
  INVX1 INVX1_624 ( .A(_abc_42016_n2780), .Y(_abc_42016_n4479_1) );
  INVX1 INVX1_625 ( .A(_auto_iopadmap_cc_313_execute_46257_2_), .Y(_abc_42016_n4484) );
  INVX1 INVX1_626 ( .A(_auto_iopadmap_cc_313_execute_46257_3_), .Y(_abc_42016_n4489) );
  INVX1 INVX1_627 ( .A(_auto_iopadmap_cc_313_execute_46257_4_), .Y(_abc_42016_n4494_1) );
  INVX1 INVX1_628 ( .A(_auto_iopadmap_cc_313_execute_46257_5_), .Y(_abc_42016_n4499) );
  INVX1 INVX1_629 ( .A(_auto_iopadmap_cc_313_execute_46257_6_), .Y(_abc_42016_n4504) );
  INVX1 INVX1_63 ( .A(regfil_1__7_), .Y(_abc_42016_n641) );
  INVX1 INVX1_630 ( .A(_auto_iopadmap_cc_313_execute_46257_7_), .Y(_abc_42016_n4509_1) );
  INVX1 INVX1_631 ( .A(_auto_iopadmap_cc_313_execute_46257_8_), .Y(_abc_42016_n4514) );
  INVX1 INVX1_632 ( .A(_auto_iopadmap_cc_313_execute_46257_13_), .Y(_abc_42016_n4535) );
  INVX1 INVX1_633 ( .A(_abc_42016_n2364), .Y(_abc_42016_n4548) );
  INVX1 INVX1_634 ( .A(_abc_42016_n4552), .Y(_abc_42016_n4553) );
  INVX1 INVX1_635 ( .A(_abc_42016_n4549), .Y(_abc_42016_n4555) );
  INVX1 INVX1_636 ( .A(_abc_42016_n4550), .Y(_abc_42016_n4556) );
  INVX1 INVX1_637 ( .A(_abc_42016_n4557), .Y(_abc_42016_n4558) );
  INVX1 INVX1_638 ( .A(_abc_42016_n4559), .Y(_abc_42016_n4560) );
  INVX1 INVX1_639 ( .A(_abc_42016_n2363), .Y(_abc_42016_n4564) );
  INVX1 INVX1_64 ( .A(regfil_1__5_), .Y(_abc_42016_n642) );
  INVX1 INVX1_640 ( .A(_abc_42016_n4565), .Y(_abc_42016_n4566) );
  INVX1 INVX1_641 ( .A(_abc_42016_n4568), .Y(_abc_42016_n4569) );
  INVX1 INVX1_642 ( .A(_abc_42016_n4574), .Y(_abc_42016_n4575) );
  INVX1 INVX1_643 ( .A(_abc_42016_n2410), .Y(_abc_42016_n4577) );
  INVX1 INVX1_644 ( .A(_abc_42016_n4580), .Y(_abc_42016_n4581) );
  INVX1 INVX1_645 ( .A(_abc_42016_n4582), .Y(_abc_42016_n4583) );
  INVX1 INVX1_646 ( .A(_abc_42016_n4587), .Y(_abc_42016_n4588) );
  INVX1 INVX1_647 ( .A(_abc_42016_n4589), .Y(_abc_42016_n4590) );
  INVX1 INVX1_648 ( .A(_abc_42016_n4593), .Y(_abc_42016_n4594) );
  INVX1 INVX1_649 ( .A(_abc_42016_n4595), .Y(_abc_42016_n4596) );
  INVX1 INVX1_65 ( .A(regfil_1__3_), .Y(_abc_42016_n643_1) );
  INVX1 INVX1_650 ( .A(_abc_42016_n4601), .Y(_abc_42016_n4602) );
  INVX1 INVX1_651 ( .A(_abc_42016_n4617), .Y(_abc_42016_n4618) );
  INVX1 INVX1_652 ( .A(_abc_42016_n4624), .Y(_abc_42016_n4625) );
  INVX1 INVX1_653 ( .A(_abc_42016_n4630), .Y(_abc_42016_n4631_1) );
  INVX1 INVX1_654 ( .A(_abc_42016_n4673), .Y(_abc_42016_n4674_1) );
  INVX1 INVX1_655 ( .A(_abc_42016_n4637), .Y(_abc_42016_n4701) );
  INVX1 INVX1_656 ( .A(_abc_42016_n4675), .Y(_abc_42016_n4731_1) );
  INVX1 INVX1_657 ( .A(ei), .Y(_abc_42016_n4736) );
  INVX1 INVX1_658 ( .A(eienb), .Y(_abc_42016_n4737_1) );
  INVX1 INVX1_659 ( .A(alu_opra_3_), .Y(alu__abc_41682_n48) );
  INVX1 INVX1_66 ( .A(regfil_1__0_), .Y(_abc_42016_n644) );
  INVX1 INVX1_660 ( .A(alu_oprb_3_), .Y(alu__abc_41682_n50_1) );
  INVX1 INVX1_661 ( .A(alu__abc_41682_n53), .Y(alu__abc_41682_n54) );
  INVX1 INVX1_662 ( .A(alu__abc_41682_n60), .Y(alu__abc_41682_n61) );
  INVX1 INVX1_663 ( .A(alu__abc_41682_n63), .Y(alu__abc_41682_n64) );
  INVX1 INVX1_664 ( .A(alu__abc_41682_n68), .Y(alu__abc_41682_n69) );
  INVX1 INVX1_665 ( .A(alu__abc_41682_n73), .Y(alu__abc_41682_n74) );
  INVX1 INVX1_666 ( .A(alu__abc_41682_n76), .Y(alu__abc_41682_n77) );
  INVX1 INVX1_667 ( .A(alu__abc_41682_n75), .Y(alu__abc_41682_n82) );
  INVX1 INVX1_668 ( .A(alu_oprb_6_), .Y(alu__abc_41682_n85) );
  INVX1 INVX1_669 ( .A(alu_opra_6_), .Y(alu__abc_41682_n86) );
  INVX1 INVX1_67 ( .A(regfil_1__1_), .Y(_abc_42016_n645) );
  INVX1 INVX1_670 ( .A(alu__abc_41682_n88), .Y(alu__abc_41682_n90) );
  INVX1 INVX1_671 ( .A(alu__abc_41682_n87), .Y(alu__abc_41682_n94) );
  INVX1 INVX1_672 ( .A(alu_oprb_7_), .Y(alu__abc_41682_n96) );
  INVX1 INVX1_673 ( .A(alu_opra_7_), .Y(alu__abc_41682_n97) );
  INVX1 INVX1_674 ( .A(alu__abc_41682_n101), .Y(alu__abc_41682_n102) );
  INVX1 INVX1_675 ( .A(alu_sel_0_), .Y(alu__abc_41682_n104) );
  INVX1 INVX1_676 ( .A(alu__abc_41682_n105), .Y(alu__abc_41682_n106) );
  INVX1 INVX1_677 ( .A(alu__abc_41682_n99), .Y(alu__abc_41682_n108) );
  INVX1 INVX1_678 ( .A(alu__abc_41682_n109), .Y(alu__abc_41682_n110) );
  INVX1 INVX1_679 ( .A(alu__abc_41682_n84), .Y(alu__abc_41682_n114) );
  INVX1 INVX1_68 ( .A(_abc_42016_n654), .Y(_abc_42016_n655_1) );
  INVX1 INVX1_680 ( .A(alu_opra_5_), .Y(alu__abc_41682_n115) );
  INVX1 INVX1_681 ( .A(alu__abc_41682_n116), .Y(alu__abc_41682_n117) );
  INVX1 INVX1_682 ( .A(alu_opra_4_), .Y(alu__abc_41682_n118) );
  INVX1 INVX1_683 ( .A(alu__abc_41682_n59), .Y(alu__abc_41682_n120) );
  INVX1 INVX1_684 ( .A(alu_opra_2_), .Y(alu__abc_41682_n121) );
  INVX1 INVX1_685 ( .A(alu_opra_1_), .Y(alu__abc_41682_n123) );
  INVX1 INVX1_686 ( .A(alu_oprb_0_), .Y(alu__abc_41682_n125) );
  INVX1 INVX1_687 ( .A(alu__abc_41682_n119), .Y(alu__abc_41682_n134) );
  INVX1 INVX1_688 ( .A(alu__abc_41682_n62), .Y(alu__abc_41682_n135) );
  INVX1 INVX1_689 ( .A(alu__abc_41682_n122), .Y(alu__abc_41682_n136) );
  INVX1 INVX1_69 ( .A(_abc_42016_n656), .Y(_abc_42016_n657) );
  INVX1 INVX1_690 ( .A(alu_opra_0_), .Y(alu__abc_41682_n139) );
  INVX1 INVX1_691 ( .A(alu__abc_41682_n132), .Y(alu__abc_41682_n147) );
  INVX1 INVX1_692 ( .A(alu_sel_1_), .Y(alu__abc_41682_n149) );
  INVX1 INVX1_693 ( .A(alu_sel_2_), .Y(alu__abc_41682_n153) );
  INVX1 INVX1_694 ( .A(alu__abc_41682_n154), .Y(alu__abc_41682_n155) );
  INVX1 INVX1_695 ( .A(alu__abc_41682_n150), .Y(alu__abc_41682_n158) );
  INVX1 INVX1_696 ( .A(alu__abc_41682_n161), .Y(alu__abc_41682_n162) );
  INVX1 INVX1_697 ( .A(alu__abc_41682_n52), .Y(alu__abc_41682_n169_1) );
  INVX1 INVX1_698 ( .A(alu__abc_41682_n173), .Y(alu__abc_41682_n174) );
  INVX1 INVX1_699 ( .A(alu__abc_41682_n181), .Y(alu__abc_41682_n182) );
  INVX1 INVX1_7 ( .A(_abc_42016_n510), .Y(_abc_42016_n511) );
  INVX1 INVX1_70 ( .A(_abc_42016_n659_1), .Y(_abc_42016_n660) );
  INVX1 INVX1_700 ( .A(alu__abc_41682_n193), .Y(alu__abc_41682_n194) );
  INVX1 INVX1_701 ( .A(alu__abc_41682_n196), .Y(alu_sout) );
  INVX1 INVX1_702 ( .A(alu__abc_41682_n107), .Y(alu__abc_41682_n198) );
  INVX1 INVX1_703 ( .A(alu__abc_41682_n163), .Y(alu__abc_41682_n202) );
  INVX1 INVX1_704 ( .A(alu__abc_41682_n224), .Y(alu__abc_41682_n226) );
  INVX1 INVX1_705 ( .A(alu__abc_41682_n40), .Y(alu__abc_41682_n232) );
  INVX1 INVX1_706 ( .A(alu__abc_41682_n179), .Y(alu__abc_41682_n240) );
  INVX1 INVX1_707 ( .A(alu__abc_41682_n80), .Y(alu__abc_41682_n247) );
  INVX1 INVX1_708 ( .A(alu__abc_41682_n259_1), .Y(alu__abc_41682_n260) );
  INVX1 INVX1_709 ( .A(alu__abc_41682_n159), .Y(alu__abc_41682_n265) );
  INVX1 INVX1_71 ( .A(_abc_42016_n663), .Y(_abc_42016_n664_1) );
  INVX1 INVX1_710 ( .A(alu__abc_41682_n288), .Y(alu__abc_41682_n289) );
  INVX1 INVX1_711 ( .A(alu__abc_41682_n291), .Y(alu__abc_41682_n292) );
  INVX1 INVX1_712 ( .A(alu__abc_41682_n246), .Y(alu__abc_41682_n320) );
  INVX1 INVX1_713 ( .A(alu__abc_41682_n225), .Y(alu__abc_41682_n329) );
  INVX1 INVX1_714 ( .A(alu__abc_41682_n133), .Y(alu__abc_41682_n362) );
  INVX1 INVX1_72 ( .A(_abc_42016_n666), .Y(_abc_42016_n667) );
  INVX1 INVX1_73 ( .A(_abc_42016_n668), .Y(_abc_42016_n669) );
  INVX1 INVX1_74 ( .A(_abc_42016_n670), .Y(_abc_42016_n671_1) );
  INVX1 INVX1_75 ( .A(opcode_7_), .Y(_abc_42016_n672_1) );
  INVX1 INVX1_76 ( .A(_abc_42016_n673), .Y(_abc_42016_n674) );
  INVX1 INVX1_77 ( .A(_abc_42016_n675), .Y(_abc_42016_n676) );
  INVX1 INVX1_78 ( .A(_abc_42016_n677), .Y(_abc_42016_n678) );
  INVX1 INVX1_79 ( .A(_abc_42016_n679), .Y(_abc_42016_n680) );
  INVX1 INVX1_8 ( .A(_abc_42016_n512), .Y(_abc_42016_n513) );
  INVX1 INVX1_80 ( .A(_abc_42016_n573), .Y(_abc_42016_n682) );
  INVX1 INVX1_81 ( .A(popdes_0_), .Y(_abc_42016_n686) );
  INVX1 INVX1_82 ( .A(_abc_42016_n688), .Y(_abc_42016_n689) );
  INVX1 INVX1_83 ( .A(_abc_42016_n691), .Y(_abc_42016_n692) );
  INVX1 INVX1_84 ( .A(regfil_5__0_), .Y(_abc_42016_n695) );
  INVX1 INVX1_85 ( .A(_abc_42016_n696), .Y(_abc_42016_n697) );
  INVX1 INVX1_86 ( .A(_abc_42016_n694), .Y(_abc_42016_n701) );
  INVX1 INVX1_87 ( .A(regfil_3__1_), .Y(_abc_42016_n703) );
  INVX1 INVX1_88 ( .A(regfil_5__1_), .Y(_abc_42016_n709) );
  INVX1 INVX1_89 ( .A(regfil_0__1_), .Y(_abc_42016_n712) );
  INVX1 INVX1_9 ( .A(state_4_), .Y(_abc_42016_n514) );
  INVX1 INVX1_90 ( .A(_abc_42016_n715), .Y(_abc_42016_n716) );
  INVX1 INVX1_91 ( .A(rdatahold_1_), .Y(_abc_42016_n719) );
  INVX1 INVX1_92 ( .A(_abc_42016_n588_1), .Y(_abc_42016_n720) );
  INVX1 INVX1_93 ( .A(regfil_4__1_), .Y(_abc_42016_n722) );
  INVX1 INVX1_94 ( .A(regfil_6__1_), .Y(_abc_42016_n723) );
  INVX1 INVX1_95 ( .A(_abc_42016_n630), .Y(_abc_42016_n727) );
  INVX1 INVX1_96 ( .A(regfil_2__1_), .Y(_abc_42016_n728) );
  INVX1 INVX1_97 ( .A(_abc_42016_n738), .Y(_abc_42016_n739) );
  INVX1 INVX1_98 ( .A(regfil_0__2_), .Y(_abc_42016_n743) );
  INVX1 INVX1_99 ( .A(_abc_42016_n746), .Y(_abc_42016_n747) );
  MUX2X1 MUX2X1_1 ( .A(_abc_42016_n739), .B(regfil_5__1_), .S(_abc_42016_n989), .Y(_abc_42016_n1092) );
  MUX2X1 MUX2X1_10 ( .A(_abc_42016_n530), .B(_abc_42016_n2246), .S(_abc_42016_n2230), .Y(opcode_5__FF_INPUT) );
  MUX2X1 MUX2X1_11 ( .A(_abc_42016_n540), .B(_abc_42016_n2248), .S(_abc_42016_n2230), .Y(opcode_6__FF_INPUT) );
  MUX2X1 MUX2X1_12 ( .A(_abc_42016_n891), .B(_abc_42016_n2246), .S(_abc_42016_n2462), .Y(rdatahold_5__FF_INPUT) );
  MUX2X1 MUX2X1_13 ( .A(_abc_42016_n757), .B(_abc_42016_n3078_1), .S(_abc_42016_n2279), .Y(_abc_42016_n3087) );
  MUX2X1 MUX2X1_14 ( .A(_abc_42016_n3314), .B(_abc_42016_n3291), .S(_abc_42016_n3072), .Y(waddrhold_11__FF_INPUT) );
  MUX2X1 MUX2X1_15 ( .A(_abc_42016_n1488), .B(_abc_42016_n4395), .S(_abc_42016_n4394), .Y(_abc_42016_n4396) );
  MUX2X1 MUX2X1_16 ( .A(alu__abc_41682_n311), .B(alu__abc_41682_n139), .S(alu__abc_41682_n339), .Y(alu_res_0_) );
  MUX2X1 MUX2X1_17 ( .A(alu__abc_41682_n303), .B(alu__abc_41682_n123), .S(alu__abc_41682_n339), .Y(alu_res_1_) );
  MUX2X1 MUX2X1_18 ( .A(alu__abc_41682_n321), .B(alu__abc_41682_n115), .S(alu__abc_41682_n339), .Y(alu_res_5_) );
  MUX2X1 MUX2X1_2 ( .A(_abc_42016_n858), .B(regfil_5__4_), .S(_abc_42016_n989), .Y(_abc_42016_n1221_1) );
  MUX2X1 MUX2X1_3 ( .A(_abc_42016_n909), .B(regfil_5__5_), .S(_abc_42016_n989), .Y(_abc_42016_n1257) );
  MUX2X1 MUX2X1_4 ( .A(_abc_42016_n1586_1), .B(pc_15_), .S(pc_0_), .Y(_abc_42016_n1587) );
  MUX2X1 MUX2X1_5 ( .A(_abc_42016_n1626), .B(_abc_42016_n1643), .S(_abc_42016_n720), .Y(_abc_36783_n3554) );
  MUX2X1 MUX2X1_6 ( .A(_abc_42016_n739), .B(regfil_2__1_), .S(_abc_42016_n1767_1), .Y(_abc_42016_n1771) );
  MUX2X1 MUX2X1_7 ( .A(_abc_42016_n819), .B(regfil_2__3_), .S(_abc_42016_n1767_1), .Y(_abc_42016_n1777) );
  MUX2X1 MUX2X1_8 ( .A(_abc_42016_n1456), .B(_abc_42016_n1949), .S(_abc_42016_n566), .Y(_abc_42016_n1950_1) );
  MUX2X1 MUX2X1_9 ( .A(_abc_42016_n2076), .B(_abc_42016_n2064), .S(_abc_42016_n2065), .Y(auxcar_FF_INPUT) );
  NAND2X1 NAND2X1_1 ( .A(_abc_42016_n605_1), .B(_abc_42016_n561), .Y(_abc_42016_n606) );
  NAND2X1 NAND2X1_10 ( .A(_abc_42016_n657), .B(_abc_42016_n658), .Y(_abc_42016_n659_1) );
  NAND2X1 NAND2X1_100 ( .A(regfil_5__6_), .B(_abc_42016_n1006), .Y(_abc_42016_n1320) );
  NAND2X1 NAND2X1_101 ( .A(_abc_42016_n1326), .B(_abc_42016_n1329_1), .Y(_abc_42016_n1330) );
  NAND2X1 NAND2X1_102 ( .A(pc_5_), .B(_abc_42016_n1361), .Y(_abc_42016_n1362) );
  NAND2X1 NAND2X1_103 ( .A(pc_7_), .B(_abc_42016_n1363), .Y(_abc_42016_n1366) );
  NAND2X1 NAND2X1_104 ( .A(_abc_42016_n1365), .B(_abc_42016_n1368), .Y(_abc_42016_n1369) );
  NAND2X1 NAND2X1_105 ( .A(opcode_3_), .B(_abc_42016_n1373), .Y(_abc_42016_n1374) );
  NAND2X1 NAND2X1_106 ( .A(opcode_2_), .B(_abc_42016_n564), .Y(_abc_42016_n1380) );
  NAND2X1 NAND2X1_107 ( .A(pc_3_), .B(_abc_42016_n1384), .Y(_abc_42016_n1385) );
  NAND2X1 NAND2X1_108 ( .A(pc_5_), .B(_abc_42016_n1386_1), .Y(_abc_42016_n1387) );
  NAND2X1 NAND2X1_109 ( .A(pc_7_), .B(_abc_42016_n1388), .Y(_abc_42016_n1389) );
  NAND2X1 NAND2X1_11 ( .A(_abc_42016_n687), .B(_abc_42016_n582_1), .Y(_abc_42016_n688) );
  NAND2X1 NAND2X1_110 ( .A(pc_9_), .B(_abc_42016_n1391), .Y(_abc_42016_n1424) );
  NAND2X1 NAND2X1_111 ( .A(_abc_42016_n1399), .B(_abc_42016_n1429), .Y(_abc_42016_n1430) );
  NAND2X1 NAND2X1_112 ( .A(pc_9_), .B(_abc_42016_n1367), .Y(_abc_42016_n1435) );
  NAND2X1 NAND2X1_113 ( .A(_abc_42016_n1434), .B(_abc_42016_n1435), .Y(_abc_42016_n1436) );
  NAND2X1 NAND2X1_114 ( .A(opcode_4_), .B(_abc_42016_n753), .Y(_abc_42016_n1455) );
  NAND2X1 NAND2X1_115 ( .A(opcode_3_), .B(_abc_42016_n564), .Y(_abc_42016_n1461) );
  NAND2X1 NAND2X1_116 ( .A(pc_11_), .B(_abc_42016_n1466), .Y(_abc_42016_n1480) );
  NAND2X1 NAND2X1_117 ( .A(pc_11_), .B(_abc_42016_n1483), .Y(_abc_42016_n1484) );
  NAND2X1 NAND2X1_118 ( .A(_abc_42016_n1482), .B(_abc_42016_n1484), .Y(_abc_42016_n1485) );
  NAND2X1 NAND2X1_119 ( .A(_abc_42016_n1399), .B(_abc_42016_n1490), .Y(_abc_42016_n1491) );
  NAND2X1 NAND2X1_12 ( .A(regfil_0__1_), .B(_abc_42016_n619), .Y(_abc_42016_n717) );
  NAND2X1 NAND2X1_120 ( .A(pc_11_), .B(_abc_42016_n1505), .Y(_abc_42016_n1506) );
  NAND2X1 NAND2X1_121 ( .A(opcode_4_), .B(_abc_42016_n847), .Y(_abc_42016_n1514) );
  NAND2X1 NAND2X1_122 ( .A(pc_13_), .B(_abc_42016_n1510), .Y(_abc_42016_n1532) );
  NAND2X1 NAND2X1_123 ( .A(opcode_4_), .B(_abc_42016_n895), .Y(_abc_42016_n1534) );
  NAND2X1 NAND2X1_124 ( .A(pc_13_), .B(_abc_42016_n1543), .Y(_abc_42016_n1544) );
  NAND2X1 NAND2X1_125 ( .A(_abc_42016_n1542), .B(_abc_42016_n1544), .Y(_abc_42016_n1545) );
  NAND2X1 NAND2X1_126 ( .A(pc_14_), .B(_abc_42016_n1560), .Y(_abc_42016_n1561) );
  NAND2X1 NAND2X1_127 ( .A(pc_13_), .B(_abc_42016_n1565), .Y(_abc_42016_n1566) );
  NAND2X1 NAND2X1_128 ( .A(opcode_4_), .B(_abc_42016_n919), .Y(_abc_42016_n1572) );
  NAND2X1 NAND2X1_129 ( .A(opcode_4_), .B(regfil_2__7_), .Y(_abc_42016_n1592_1) );
  NAND2X1 NAND2X1_13 ( .A(alu_res_1_), .B(_abc_42016_n552), .Y(_abc_42016_n733) );
  NAND2X1 NAND2X1_130 ( .A(_abc_42016_n530), .B(_abc_42016_n1593), .Y(_abc_42016_n1594_1) );
  NAND2X1 NAND2X1_131 ( .A(_abc_42016_n554), .B(_abc_42016_n1603_1), .Y(_abc_42016_n1604_1) );
  NAND2X1 NAND2X1_132 ( .A(_abc_42016_n1606_1), .B(_abc_42016_n769), .Y(_abc_42016_n1611) );
  NAND2X1 NAND2X1_133 ( .A(_abc_42016_n1606_1), .B(_abc_42016_n858), .Y(_abc_42016_n1615) );
  NAND2X1 NAND2X1_134 ( .A(_abc_42016_n1606_1), .B(_abc_42016_n909), .Y(_abc_42016_n1617) );
  NAND2X1 NAND2X1_135 ( .A(_abc_42016_n1606_1), .B(_abc_42016_n934), .Y(_abc_42016_n1619) );
  NAND2X1 NAND2X1_136 ( .A(regfil_2__0_), .B(_abc_42016_n980), .Y(_abc_42016_n1627) );
  NAND2X1 NAND2X1_137 ( .A(regfil_4__0_), .B(_abc_42016_n696), .Y(_abc_42016_n1635) );
  NAND2X1 NAND2X1_138 ( .A(_abc_42016_n728), .B(_abc_42016_n1633), .Y(_abc_42016_n1651) );
  NAND2X1 NAND2X1_139 ( .A(regfil_4__1_), .B(_abc_42016_n696), .Y(_abc_42016_n1654) );
  NAND2X1 NAND2X1_14 ( .A(regfil_0__1_), .B(_abc_42016_n654), .Y(_abc_42016_n744) );
  NAND2X1 NAND2X1_140 ( .A(_abc_42016_n1623), .B(_abc_42016_n769), .Y(_abc_42016_n1663) );
  NAND2X1 NAND2X1_141 ( .A(_abc_42016_n720), .B(_abc_42016_n1664_1), .Y(_abc_42016_n1665) );
  NAND2X1 NAND2X1_142 ( .A(regfil_2__2_), .B(_abc_42016_n1647_1), .Y(_abc_42016_n1666) );
  NAND2X1 NAND2X1_143 ( .A(_abc_42016_n1680), .B(_abc_42016_n613), .Y(_abc_42016_n1681_1) );
  NAND2X1 NAND2X1_144 ( .A(_abc_42016_n643_1), .B(_abc_42016_n647), .Y(_abc_42016_n1688) );
  NAND2X1 NAND2X1_145 ( .A(regfil_1__3_), .B(_abc_42016_n613), .Y(_abc_42016_n1691) );
  NAND2X1 NAND2X1_146 ( .A(_abc_42016_n1693), .B(_abc_42016_n1689_1), .Y(_abc_42016_n1694) );
  NAND2X1 NAND2X1_147 ( .A(_abc_42016_n796), .B(_abc_42016_n1672), .Y(_abc_42016_n1700) );
  NAND2X1 NAND2X1_148 ( .A(_abc_42016_n1623), .B(_abc_42016_n858), .Y(_abc_42016_n1706_1) );
  NAND2X1 NAND2X1_149 ( .A(_abc_42016_n720), .B(_abc_42016_n1707), .Y(_abc_42016_n1708) );
  NAND2X1 NAND2X1_15 ( .A(_abc_42016_n743), .B(_abc_42016_n715), .Y(_abc_42016_n748) );
  NAND2X1 NAND2X1_150 ( .A(_abc_42016_n1721_1), .B(_abc_42016_n615), .Y(_abc_42016_n1722_1) );
  NAND2X1 NAND2X1_151 ( .A(_abc_42016_n895), .B(_abc_42016_n1715), .Y(_abc_42016_n1733) );
  NAND2X1 NAND2X1_152 ( .A(regfil_2__4_), .B(_abc_42016_n1711), .Y(_abc_42016_n1736) );
  NAND2X1 NAND2X1_153 ( .A(regfil_2__6_), .B(_abc_42016_n1737), .Y(_abc_42016_n1805) );
  NAND2X1 NAND2X1_154 ( .A(_abc_42016_n1815), .B(_abc_42016_n769), .Y(_abc_42016_n1820_1) );
  NAND2X1 NAND2X1_155 ( .A(_abc_42016_n1815), .B(_abc_42016_n909), .Y(_abc_42016_n1827) );
  NAND2X1 NAND2X1_156 ( .A(_abc_42016_n1815), .B(_abc_42016_n934), .Y(_abc_42016_n1830) );
  NAND2X1 NAND2X1_157 ( .A(alu_sel_0_), .B(_abc_42016_n1839), .Y(_abc_42016_n1840) );
  NAND2X1 NAND2X1_158 ( .A(_abc_42016_n1856_1), .B(_abc_42016_n1838_1), .Y(_abc_42016_n1857) );
  NAND2X1 NAND2X1_159 ( .A(alu_sel_2_), .B(_abc_42016_n1857), .Y(_abc_42016_n1858) );
  NAND2X1 NAND2X1_16 ( .A(_abc_42016_n749), .B(_abc_42016_n748), .Y(_abc_42016_n750) );
  NAND2X1 NAND2X1_160 ( .A(_abc_42016_n1851), .B(_abc_42016_n637), .Y(_abc_42016_n1864) );
  NAND2X1 NAND2X1_161 ( .A(opcode_4_), .B(_abc_42016_n634), .Y(_abc_42016_n1903_1) );
  NAND2X1 NAND2X1_162 ( .A(opcode_3_), .B(_abc_42016_n1904), .Y(_abc_42016_n1905_1) );
  NAND2X1 NAND2X1_163 ( .A(regfil_6__0_), .B(_abc_42016_n532_1), .Y(_abc_42016_n1913) );
  NAND2X1 NAND2X1_164 ( .A(_abc_42016_n557), .B(_abc_42016_n1921), .Y(_abc_42016_n1922_1) );
  NAND2X1 NAND2X1_165 ( .A(alu_opra_0_), .B(_abc_42016_n1928), .Y(_abc_42016_n1929) );
  NAND2X1 NAND2X1_166 ( .A(rdatahold_0_), .B(_abc_42016_n1930), .Y(_abc_42016_n1931) );
  NAND2X1 NAND2X1_167 ( .A(regfil_1__2_), .B(_abc_42016_n531), .Y(_abc_42016_n1949) );
  NAND2X1 NAND2X1_168 ( .A(_abc_42016_n557), .B(_abc_42016_n1956), .Y(_abc_42016_n1957_1) );
  NAND2X1 NAND2X1_169 ( .A(alu_opra_2_), .B(_abc_42016_n1928), .Y(_abc_42016_n1958) );
  NAND2X1 NAND2X1_17 ( .A(_abc_42016_n536), .B(_abc_42016_n754), .Y(_abc_42016_n755) );
  NAND2X1 NAND2X1_170 ( .A(rdatahold_2_), .B(_abc_42016_n1930), .Y(_abc_42016_n1959) );
  NAND2X1 NAND2X1_171 ( .A(_abc_42016_n2014), .B(_abc_42016_n2018), .Y(_abc_42016_n2019) );
  NAND2X1 NAND2X1_172 ( .A(_abc_42016_n510), .B(_abc_42016_n1871), .Y(_abc_42016_n2024) );
  NAND2X1 NAND2X1_173 ( .A(alu_res_7_), .B(_abc_42016_n2059), .Y(_abc_42016_n2060) );
  NAND2X1 NAND2X1_174 ( .A(regfil_7__5_), .B(_abc_42016_n2067), .Y(_abc_42016_n2068) );
  NAND2X1 NAND2X1_175 ( .A(regfil_4__6_), .B(sp_14_), .Y(_abc_42016_n2104) );
  NAND2X1 NAND2X1_176 ( .A(_abc_42016_n1554), .B(_abc_42016_n2103), .Y(_abc_42016_n2105) );
  NAND2X1 NAND2X1_177 ( .A(regfil_4__4_), .B(sp_12_), .Y(_abc_42016_n2112) );
  NAND2X1 NAND2X1_178 ( .A(_abc_42016_n842), .B(_abc_42016_n2113), .Y(_abc_42016_n2114) );
  NAND2X1 NAND2X1_179 ( .A(regfil_4__2_), .B(sp_10_), .Y(_abc_42016_n2121) );
  NAND2X1 NAND2X1_18 ( .A(_abc_42016_n761), .B(_abc_42016_n624), .Y(_abc_42016_n762) );
  NAND2X1 NAND2X1_180 ( .A(_abc_42016_n1446), .B(_abc_42016_n2122), .Y(_abc_42016_n2123_1) );
  NAND2X1 NAND2X1_181 ( .A(regfil_4__0_), .B(sp_8_), .Y(_abc_42016_n2130) );
  NAND2X1 NAND2X1_182 ( .A(_abc_42016_n629), .B(_abc_42016_n2131_1), .Y(_abc_42016_n2132_1) );
  NAND2X1 NAND2X1_183 ( .A(regfil_5__6_), .B(sp_6_), .Y(_abc_42016_n2134) );
  NAND2X1 NAND2X1_184 ( .A(regfil_2__6_), .B(regfil_4__6_), .Y(_abc_42016_n2148) );
  NAND2X1 NAND2X1_185 ( .A(_abc_42016_n895), .B(_abc_42016_n1527), .Y(_abc_42016_n2150) );
  NAND2X1 NAND2X1_186 ( .A(regfil_2__4_), .B(regfil_4__4_), .Y(_abc_42016_n2153) );
  NAND2X1 NAND2X1_187 ( .A(regfil_2__2_), .B(regfil_4__2_), .Y(_abc_42016_n2159) );
  NAND2X1 NAND2X1_188 ( .A(_abc_42016_n753), .B(_abc_42016_n1446), .Y(_abc_42016_n2160) );
  NAND2X1 NAND2X1_189 ( .A(_abc_42016_n728), .B(_abc_42016_n722), .Y(_abc_42016_n2162) );
  NAND2X1 NAND2X1_19 ( .A(_abc_42016_n763_1), .B(_abc_42016_n762), .Y(_abc_42016_n764) );
  NAND2X1 NAND2X1_190 ( .A(regfil_2__0_), .B(regfil_4__0_), .Y(_abc_42016_n2165) );
  NAND2X1 NAND2X1_191 ( .A(_abc_42016_n2148), .B(_abc_42016_n2176), .Y(_abc_42016_n2177) );
  NAND2X1 NAND2X1_192 ( .A(regfil_0__6_), .B(regfil_4__6_), .Y(_abc_42016_n2180) );
  NAND2X1 NAND2X1_193 ( .A(_abc_42016_n913), .B(_abc_42016_n1554), .Y(_abc_42016_n2181) );
  NAND2X1 NAND2X1_194 ( .A(_abc_42016_n893), .B(_abc_42016_n1527), .Y(_abc_42016_n2183) );
  NAND2X1 NAND2X1_195 ( .A(regfil_0__4_), .B(regfil_4__4_), .Y(_abc_42016_n2186) );
  NAND2X1 NAND2X1_196 ( .A(_abc_42016_n812), .B(_abc_42016_n800), .Y(_abc_42016_n2188) );
  NAND2X1 NAND2X1_197 ( .A(regfil_0__2_), .B(regfil_4__2_), .Y(_abc_42016_n2191) );
  NAND2X1 NAND2X1_198 ( .A(_abc_42016_n743), .B(_abc_42016_n1446), .Y(_abc_42016_n2192) );
  NAND2X1 NAND2X1_199 ( .A(_abc_42016_n712), .B(_abc_42016_n722), .Y(_abc_42016_n2194) );
  NAND2X1 NAND2X1_2 ( .A(_abc_42016_n611), .B(_abc_42016_n612), .Y(_abc_42016_n613) );
  NAND2X1 NAND2X1_20 ( .A(_abc_42016_n683), .B(_abc_42016_n658), .Y(_abc_42016_n772) );
  NAND2X1 NAND2X1_200 ( .A(regfil_0__0_), .B(regfil_4__0_), .Y(_abc_42016_n2197) );
  NAND2X1 NAND2X1_201 ( .A(_abc_42016_n608), .B(_abc_42016_n629), .Y(_abc_42016_n2199) );
  NAND2X1 NAND2X1_202 ( .A(alu_cout), .B(_abc_42016_n2034), .Y(_abc_42016_n2219) );
  NAND2X1 NAND2X1_203 ( .A(_abc_42016_n510), .B(_abc_42016_n2227), .Y(_abc_42016_n2228) );
  NAND2X1 NAND2X1_204 ( .A(_abc_42016_n2226), .B(_abc_42016_n2229), .Y(_abc_42016_n2230) );
  NAND2X1 NAND2X1_205 ( .A(_abc_42016_n2030), .B(_abc_42016_n2260), .Y(_abc_42016_n2261) );
  NAND2X1 NAND2X1_206 ( .A(_abc_42016_n2030), .B(_abc_42016_n2266), .Y(_abc_42016_n2267) );
  NAND2X1 NAND2X1_207 ( .A(_abc_42016_n2265), .B(_abc_42016_n2274), .Y(_abc_42016_n2275) );
  NAND2X1 NAND2X1_208 ( .A(_abc_42016_n529), .B(_abc_42016_n2277), .Y(_abc_42016_n2278) );
  NAND2X1 NAND2X1_209 ( .A(_abc_42016_n2279), .B(_abc_42016_n2297_1), .Y(_abc_42016_n2298) );
  NAND2X1 NAND2X1_21 ( .A(regfil_3__2_), .B(_abc_42016_n704), .Y(_abc_42016_n775) );
  NAND2X1 NAND2X1_210 ( .A(_abc_42016_n673), .B(_abc_42016_n2330), .Y(_abc_42016_n2331) );
  NAND2X1 NAND2X1_211 ( .A(_abc_42016_n2305), .B(_abc_42016_n2331), .Y(_abc_42016_n2332) );
  NAND2X1 NAND2X1_212 ( .A(_abc_42016_n2370), .B(_abc_42016_n1835), .Y(_abc_42016_n2371) );
  NAND2X1 NAND2X1_213 ( .A(statesel_2_), .B(_abc_42016_n2387), .Y(_abc_42016_n2388) );
  NAND2X1 NAND2X1_214 ( .A(_abc_42016_n2386), .B(_abc_42016_n2388), .Y(_abc_42016_n2389) );
  NAND2X1 NAND2X1_215 ( .A(_abc_42016_n2397), .B(_abc_42016_n2282), .Y(_abc_42016_n2398_1) );
  NAND2X1 NAND2X1_216 ( .A(_abc_42016_n2322), .B(_abc_42016_n2318), .Y(_abc_42016_n2418) );
  NAND2X1 NAND2X1_217 ( .A(_abc_42016_n2430), .B(_abc_42016_n2428), .Y(_abc_42016_n2431) );
  NAND2X1 NAND2X1_218 ( .A(_abc_42016_n2347_1), .B(_abc_42016_n677), .Y(_abc_42016_n2457) );
  NAND2X1 NAND2X1_219 ( .A(_abc_42016_n2226), .B(_abc_42016_n2334), .Y(_abc_42016_n2462) );
  NAND2X1 NAND2X1_22 ( .A(_abc_42016_n774), .B(_abc_42016_n775), .Y(_abc_42016_n776) );
  NAND2X1 NAND2X1_220 ( .A(_abc_42016_n1015), .B(_abc_42016_n1013), .Y(_abc_42016_n2497) );
  NAND2X1 NAND2X1_221 ( .A(opcode_4_), .B(regfil_3__1_), .Y(_abc_42016_n2527) );
  NAND2X1 NAND2X1_222 ( .A(_abc_42016_n540), .B(_abc_42016_n1346), .Y(_abc_42016_n2542) );
  NAND2X1 NAND2X1_223 ( .A(wdatahold_1_), .B(_abc_42016_n2499), .Y(_abc_42016_n2553) );
  NAND2X1 NAND2X1_224 ( .A(pc_0_), .B(_abc_42016_n1384), .Y(_abc_42016_n2559) );
  NAND2X1 NAND2X1_225 ( .A(regfil_5__2_), .B(_abc_42016_n668), .Y(_abc_42016_n2566) );
  NAND2X1 NAND2X1_226 ( .A(_abc_42016_n2576), .B(_abc_42016_n2512), .Y(_abc_42016_n2577) );
  NAND2X1 NAND2X1_227 ( .A(_abc_42016_n1357), .B(_abc_42016_n2559), .Y(_abc_42016_n2591) );
  NAND2X1 NAND2X1_228 ( .A(opcode_4_), .B(_abc_42016_n795), .Y(_abc_42016_n2596) );
  NAND2X1 NAND2X1_229 ( .A(_abc_42016_n2598), .B(_abc_42016_n1401), .Y(_abc_42016_n2599) );
  NAND2X1 NAND2X1_23 ( .A(_abc_42016_n681), .B(_abc_42016_n561), .Y(_abc_42016_n778_1) );
  NAND2X1 NAND2X1_230 ( .A(wdatahold_3_), .B(_abc_42016_n2582), .Y(_abc_42016_n2604) );
  NAND2X1 NAND2X1_231 ( .A(_abc_42016_n2299), .B(_abc_42016_n805), .Y(_abc_42016_n2605) );
  NAND2X1 NAND2X1_232 ( .A(opcode_4_), .B(_abc_42016_n861), .Y(_abc_42016_n2621) );
  NAND2X1 NAND2X1_233 ( .A(pc_4_), .B(_abc_42016_n1404), .Y(_abc_42016_n2627) );
  NAND2X1 NAND2X1_234 ( .A(_abc_42016_n1245), .B(_abc_42016_n573), .Y(_abc_42016_n2628) );
  NAND2X1 NAND2X1_235 ( .A(_abc_42016_n2634), .B(_abc_42016_n2633), .Y(_abc_42016_n2635) );
  NAND2X1 NAND2X1_236 ( .A(wdatahold_4_), .B(_abc_42016_n2582), .Y(_abc_42016_n2638) );
  NAND2X1 NAND2X1_237 ( .A(opcode_4_), .B(regfil_3__5_), .Y(_abc_42016_n2654) );
  NAND2X1 NAND2X1_238 ( .A(_abc_42016_n2655), .B(_abc_42016_n1401), .Y(_abc_42016_n2656) );
  NAND2X1 NAND2X1_239 ( .A(_abc_42016_n2666), .B(_abc_42016_n2662), .Y(_abc_42016_n2667) );
  NAND2X1 NAND2X1_24 ( .A(_abc_42016_n798), .B(_abc_42016_n804), .Y(_abc_42016_n805) );
  NAND2X1 NAND2X1_240 ( .A(regfil_5__6_), .B(_abc_42016_n668), .Y(_abc_42016_n2680) );
  NAND2X1 NAND2X1_241 ( .A(_abc_42016_n927), .B(_abc_42016_n2299), .Y(_abc_42016_n2691) );
  NAND2X1 NAND2X1_242 ( .A(wdatahold_7_), .B(_abc_42016_n2702), .Y(_abc_42016_n2703) );
  NAND2X1 NAND2X1_243 ( .A(wdatahold2_7_), .B(_abc_42016_n2519), .Y(_abc_42016_n2705) );
  NAND2X1 NAND2X1_244 ( .A(opcode_4_), .B(_abc_42016_n974), .Y(_abc_42016_n2717) );
  NAND2X1 NAND2X1_245 ( .A(_abc_42016_n2500), .B(_abc_42016_n2728), .Y(_abc_42016_n2729) );
  NAND2X1 NAND2X1_246 ( .A(_abc_42016_n2703), .B(_abc_42016_n2729), .Y(wdatahold_7__FF_INPUT) );
  NAND2X1 NAND2X1_247 ( .A(_abc_42016_n529), .B(_abc_42016_n2734), .Y(_abc_42016_n2735) );
  NAND2X1 NAND2X1_248 ( .A(_abc_42016_n2742), .B(_abc_42016_n2315), .Y(_abc_42016_n2743) );
  NAND2X1 NAND2X1_249 ( .A(_abc_42016_n2502), .B(_abc_42016_n2281), .Y(_abc_42016_n2751) );
  NAND2X1 NAND2X1_25 ( .A(_abc_42016_n808), .B(_abc_42016_n720), .Y(_abc_42016_n809) );
  NAND2X1 NAND2X1_250 ( .A(_abc_42016_n1344), .B(_abc_42016_n2357), .Y(_abc_42016_n2754) );
  NAND2X1 NAND2X1_251 ( .A(_abc_42016_n2736), .B(_abc_42016_n2762), .Y(_abc_42016_n2763) );
  NAND2X1 NAND2X1_252 ( .A(_abc_42016_n547), .B(_abc_42016_n2773), .Y(_abc_42016_n2774) );
  NAND2X1 NAND2X1_253 ( .A(_abc_42016_n2781), .B(_abc_42016_n2782), .Y(_abc_42016_n2783) );
  NAND2X1 NAND2X1_254 ( .A(raddrhold_2_), .B(_abc_42016_n2777), .Y(_abc_42016_n2787) );
  NAND2X1 NAND2X1_255 ( .A(_abc_42016_n2564), .B(_abc_42016_n2309), .Y(_abc_42016_n2795) );
  NAND2X1 NAND2X1_256 ( .A(_abc_42016_n2799), .B(_abc_42016_n2797), .Y(_abc_42016_n2800) );
  NAND2X1 NAND2X1_257 ( .A(raddrhold_4_), .B(_abc_42016_n2804), .Y(_abc_42016_n2828) );
  NAND2X1 NAND2X1_258 ( .A(_abc_42016_n2655), .B(_abc_42016_n2309), .Y(_abc_42016_n2842) );
  NAND2X1 NAND2X1_259 ( .A(_abc_42016_n2844), .B(_abc_42016_n2840), .Y(_abc_42016_n2845) );
  NAND2X1 NAND2X1_26 ( .A(regfil_0__3_), .B(_abc_42016_n814), .Y(_abc_42016_n815) );
  NAND2X1 NAND2X1_260 ( .A(raddrhold_6_), .B(_abc_42016_n2847), .Y(_abc_42016_n2880) );
  NAND2X1 NAND2X1_261 ( .A(_abc_42016_n629), .B(_abc_42016_n2279), .Y(_abc_42016_n2893) );
  NAND2X1 NAND2X1_262 ( .A(_abc_42016_n2910), .B(_abc_42016_n2906), .Y(_abc_42016_n2911) );
  NAND2X1 NAND2X1_263 ( .A(raddrhold_9_), .B(_abc_42016_n2888), .Y(_abc_42016_n2912) );
  NAND2X1 NAND2X1_264 ( .A(raddrhold_9_), .B(_abc_42016_n2917), .Y(_abc_42016_n2918) );
  NAND2X1 NAND2X1_265 ( .A(raddrhold_11_), .B(_abc_42016_n2917), .Y(_abc_42016_n2940) );
  NAND2X1 NAND2X1_266 ( .A(_abc_42016_n2940), .B(_abc_42016_n2954), .Y(raddrhold_11__FF_INPUT) );
  NAND2X1 NAND2X1_267 ( .A(_abc_42016_n842), .B(_abc_42016_n2279), .Y(_abc_42016_n2957) );
  NAND2X1 NAND2X1_268 ( .A(raddrhold_12_), .B(_abc_42016_n2951), .Y(_abc_42016_n2983) );
  NAND2X1 NAND2X1_269 ( .A(raddrhold_15_), .B(_abc_42016_n2732), .Y(_abc_42016_n3023) );
  NAND2X1 NAND2X1_27 ( .A(_abc_42016_n795), .B(_abc_42016_n775), .Y(_abc_42016_n823) );
  NAND2X1 NAND2X1_270 ( .A(_abc_42016_n2261), .B(_abc_42016_n3029), .Y(_abc_42016_n3030) );
  NAND2X1 NAND2X1_271 ( .A(_abc_42016_n529), .B(_abc_42016_n3030), .Y(_abc_42016_n3031) );
  NAND2X1 NAND2X1_272 ( .A(_abc_42016_n3053), .B(_abc_42016_n3055), .Y(_abc_42016_n3056) );
  NAND2X1 NAND2X1_273 ( .A(_abc_42016_n2528), .B(_abc_42016_n3033), .Y(_abc_42016_n3062) );
  NAND2X1 NAND2X1_274 ( .A(waddrhold_2_), .B(_abc_42016_n3073), .Y(_abc_42016_n3082) );
  NAND2X1 NAND2X1_275 ( .A(_abc_42016_n1841), .B(_abc_42016_n3087), .Y(_abc_42016_n3088) );
  NAND2X1 NAND2X1_276 ( .A(_abc_42016_n1346), .B(_abc_42016_n2565), .Y(_abc_42016_n3089) );
  NAND2X1 NAND2X1_277 ( .A(waddrhold_2_), .B(_abc_42016_n3090), .Y(_abc_42016_n3091) );
  NAND2X1 NAND2X1_278 ( .A(_abc_42016_n3122), .B(_abc_42016_n3121), .Y(_abc_42016_n3123) );
  NAND2X1 NAND2X1_279 ( .A(_abc_42016_n1210), .B(_abc_42016_n3120), .Y(_abc_42016_n3131) );
  NAND2X1 NAND2X1_28 ( .A(_abc_42016_n795), .B(_abc_42016_n783), .Y(_abc_42016_n828) );
  NAND2X1 NAND2X1_280 ( .A(_abc_42016_n3132), .B(_abc_42016_n3131), .Y(_abc_42016_n3133) );
  NAND2X1 NAND2X1_281 ( .A(_abc_42016_n843), .B(_abc_42016_n2279), .Y(_abc_42016_n3138) );
  NAND2X1 NAND2X1_282 ( .A(_abc_42016_n559), .B(_abc_42016_n3156), .Y(_abc_42016_n3157) );
  NAND2X1 NAND2X1_283 ( .A(waddrhold_6_), .B(_abc_42016_n3170_1), .Y(_abc_42016_n3194) );
  NAND2X1 NAND2X1_284 ( .A(_abc_42016_n2131_1), .B(_abc_42016_n3202), .Y(_abc_42016_n3224) );
  NAND2X1 NAND2X1_285 ( .A(_abc_42016_n3241), .B(_abc_42016_n3072), .Y(_abc_42016_n3242) );
  NAND2X1 NAND2X1_286 ( .A(_abc_42016_n1841), .B(_abc_42016_n3252), .Y(_abc_42016_n3253) );
  NAND2X1 NAND2X1_287 ( .A(waddrhold_9_), .B(_abc_42016_n3238), .Y(_abc_42016_n3264) );
  NAND2X1 NAND2X1_288 ( .A(_abc_42016_n2122), .B(_abc_42016_n3248), .Y(_abc_42016_n3269) );
  NAND2X1 NAND2X1_289 ( .A(_abc_42016_n3291), .B(_abc_42016_n1851), .Y(_abc_42016_n3292) );
  NAND2X1 NAND2X1_29 ( .A(_abc_42016_n827), .B(_abc_42016_n828), .Y(_abc_42016_n829) );
  NAND2X1 NAND2X1_290 ( .A(_abc_42016_n3294), .B(_abc_42016_n3296_1), .Y(_abc_42016_n3297) );
  NAND2X1 NAND2X1_291 ( .A(_abc_42016_n559), .B(_abc_42016_n3303), .Y(_abc_42016_n3304) );
  NAND2X1 NAND2X1_292 ( .A(_abc_42016_n3305), .B(_abc_42016_n3304), .Y(_abc_42016_n3306) );
  NAND2X1 NAND2X1_293 ( .A(waddrhold_11_), .B(_abc_42016_n3285), .Y(_abc_42016_n3309) );
  NAND2X1 NAND2X1_294 ( .A(_abc_42016_n2113), .B(_abc_42016_n3295_1), .Y(_abc_42016_n3319_1) );
  NAND2X1 NAND2X1_295 ( .A(_abc_42016_n673), .B(_abc_42016_n3323), .Y(_abc_42016_n3324) );
  NAND2X1 NAND2X1_296 ( .A(_abc_42016_n1516), .B(_abc_42016_n1346), .Y(_abc_42016_n3325) );
  NAND2X1 NAND2X1_297 ( .A(_abc_42016_n3338), .B(_abc_42016_n3340), .Y(_abc_42016_n3341) );
  NAND2X1 NAND2X1_298 ( .A(_abc_42016_n3364), .B(_abc_42016_n3363), .Y(_abc_42016_n3365) );
  NAND2X1 NAND2X1_299 ( .A(waddrhold_13_), .B(_abc_42016_n3354), .Y(_abc_42016_n3380) );
  NAND2X1 NAND2X1_3 ( .A(_abc_42016_n610), .B(_abc_42016_n614), .Y(_abc_42016_n615) );
  NAND2X1 NAND2X1_30 ( .A(_abc_42016_n834), .B(_abc_42016_n789), .Y(_abc_42016_n838) );
  NAND2X1 NAND2X1_300 ( .A(_abc_42016_n3056), .B(_abc_42016_n3389), .Y(_abc_42016_n3390) );
  NAND2X1 NAND2X1_301 ( .A(_abc_42016_n1801_1), .B(_abc_42016_n2279), .Y(_abc_42016_n3395) );
  NAND2X1 NAND2X1_302 ( .A(_abc_42016_n3393), .B(_abc_42016_n3398_1), .Y(_abc_42016_n3399) );
  NAND2X1 NAND2X1_303 ( .A(_abc_42016_n510), .B(_abc_42016_n3457), .Y(_abc_42016_n3458) );
  NAND2X1 NAND2X1_304 ( .A(_abc_42016_n547), .B(_abc_42016_n3463), .Y(_abc_42016_n3464) );
  NAND2X1 NAND2X1_305 ( .A(_abc_42016_n1868), .B(_abc_42016_n2227), .Y(_abc_42016_n3503) );
  NAND2X1 NAND2X1_306 ( .A(sp_3_), .B(_abc_42016_n3098), .Y(_abc_42016_n3509) );
  NAND2X1 NAND2X1_307 ( .A(_abc_42016_n3548), .B(_abc_42016_n3540), .Y(_abc_42016_n3549) );
  NAND2X1 NAND2X1_308 ( .A(_abc_42016_n3550), .B(_abc_42016_n3501), .Y(_abc_42016_n3551) );
  NAND2X1 NAND2X1_309 ( .A(_abc_42016_n3557), .B(_abc_42016_n3556), .Y(_abc_42016_n3558) );
  NAND2X1 NAND2X1_31 ( .A(_abc_42016_n839), .B(_abc_42016_n838), .Y(_abc_42016_n840) );
  NAND2X1 NAND2X1_310 ( .A(_abc_42016_n3542), .B(_abc_42016_n2255), .Y(_abc_42016_n3562) );
  NAND2X1 NAND2X1_311 ( .A(sp_6_), .B(_abc_42016_n3555), .Y(_abc_42016_n3583) );
  NAND2X1 NAND2X1_312 ( .A(_abc_42016_n3582), .B(_abc_42016_n3583), .Y(_abc_42016_n3584) );
  NAND2X1 NAND2X1_313 ( .A(_abc_42016_n3177), .B(_abc_42016_n3542), .Y(_abc_42016_n3589) );
  NAND2X1 NAND2X1_314 ( .A(_abc_42016_n3588), .B(_abc_42016_n3598), .Y(_abc_42016_n3599) );
  NAND2X1 NAND2X1_315 ( .A(_abc_42016_n673), .B(_abc_42016_n3621), .Y(_abc_42016_n3622) );
  NAND2X1 NAND2X1_316 ( .A(sp_8_), .B(_abc_42016_n3606_1), .Y(_abc_42016_n3629) );
  NAND2X1 NAND2X1_317 ( .A(sp_7_), .B(_abc_42016_n3594), .Y(_abc_42016_n3633) );
  NAND2X1 NAND2X1_318 ( .A(_abc_42016_n3639), .B(_abc_42016_n3629), .Y(_abc_42016_n3640) );
  NAND2X1 NAND2X1_319 ( .A(sp_10_), .B(_abc_42016_n3652), .Y(_abc_42016_n3672) );
  NAND2X1 NAND2X1_32 ( .A(_abc_42016_n850), .B(_abc_42016_n624), .Y(_abc_42016_n851_1) );
  NAND2X1 NAND2X1_320 ( .A(_abc_42016_n3670_1), .B(_abc_42016_n3676), .Y(_abc_42016_n3677) );
  NAND2X1 NAND2X1_321 ( .A(_abc_42016_n3501), .B(_abc_42016_n3683), .Y(_abc_42016_n3684) );
  NAND2X1 NAND2X1_322 ( .A(_abc_42016_n2122), .B(_abc_42016_n3572), .Y(_abc_42016_n3685) );
  NAND2X1 NAND2X1_323 ( .A(sp_12_), .B(_abc_42016_n3702), .Y(_abc_42016_n3718) );
  NAND2X1 NAND2X1_324 ( .A(_abc_42016_n3474), .B(_abc_42016_n3718), .Y(_abc_42016_n3719) );
  NAND2X1 NAND2X1_325 ( .A(_abc_42016_n3724), .B(_abc_42016_n3726), .Y(_abc_42016_n3727) );
  NAND2X1 NAND2X1_326 ( .A(sp_13_), .B(_abc_42016_n3738), .Y(_abc_42016_n3739) );
  NAND2X1 NAND2X1_327 ( .A(_abc_42016_n3748), .B(_abc_42016_n3749), .Y(_abc_42016_n3750) );
  NAND2X1 NAND2X1_328 ( .A(_abc_42016_n3502), .B(_abc_42016_n3747), .Y(_abc_42016_n3753) );
  NAND2X1 NAND2X1_329 ( .A(_abc_42016_n3501), .B(_abc_42016_n3755_1), .Y(_abc_42016_n3756) );
  NAND2X1 NAND2X1_33 ( .A(_abc_42016_n852), .B(_abc_42016_n851_1), .Y(_abc_42016_n853) );
  NAND2X1 NAND2X1_330 ( .A(sp_14_), .B(_abc_42016_n3746), .Y(_abc_42016_n3762) );
  NAND2X1 NAND2X1_331 ( .A(_abc_42016_n3768), .B(_abc_42016_n3762), .Y(_abc_42016_n3769) );
  NAND2X1 NAND2X1_332 ( .A(_abc_42016_n3785), .B(_abc_42016_n3782), .Y(_abc_42016_n3786) );
  NAND2X1 NAND2X1_333 ( .A(_abc_42016_n3527), .B(_abc_42016_n3389), .Y(_abc_42016_n3794) );
  NAND2X1 NAND2X1_334 ( .A(_abc_42016_n3795), .B(_abc_42016_n3794), .Y(_abc_42016_n3796) );
  NAND2X1 NAND2X1_335 ( .A(_abc_42016_n997), .B(_abc_42016_n3804), .Y(_abc_42016_n3805) );
  NAND2X1 NAND2X1_336 ( .A(_abc_42016_n629), .B(_abc_42016_n1335_1), .Y(_abc_42016_n3806) );
  NAND2X1 NAND2X1_337 ( .A(regfil_4__0_), .B(_abc_42016_n1337_1), .Y(_abc_42016_n3810) );
  NAND2X1 NAND2X1_338 ( .A(_abc_42016_n2136_1), .B(_abc_42016_n3815), .Y(_abc_42016_n3816) );
  NAND2X1 NAND2X1_339 ( .A(_abc_42016_n2203), .B(_abc_42016_n3820), .Y(_abc_42016_n3821) );
  NAND2X1 NAND2X1_34 ( .A(regfil_3__4_), .B(_abc_42016_n824), .Y(_abc_42016_n863) );
  NAND2X1 NAND2X1_340 ( .A(_abc_42016_n2194), .B(_abc_42016_n2196), .Y(_abc_42016_n3847) );
  NAND2X1 NAND2X1_341 ( .A(_abc_42016_n2162), .B(_abc_42016_n2164), .Y(_abc_42016_n3850) );
  NAND2X1 NAND2X1_342 ( .A(_abc_42016_n1446), .B(_abc_42016_n3856), .Y(_abc_42016_n3867) );
  NAND2X1 NAND2X1_343 ( .A(regfil_4__2_), .B(_abc_42016_n3838), .Y(_abc_42016_n3872) );
  NAND2X1 NAND2X1_344 ( .A(_abc_42016_n3871), .B(_abc_42016_n3872), .Y(_abc_42016_n3873) );
  NAND2X1 NAND2X1_345 ( .A(_abc_42016_n3881), .B(_abc_42016_n3882), .Y(_abc_42016_n3883) );
  NAND2X1 NAND2X1_346 ( .A(_abc_42016_n673), .B(_abc_42016_n557), .Y(_abc_42016_n3890) );
  NAND2X1 NAND2X1_347 ( .A(_abc_42016_n2188), .B(_abc_42016_n2190), .Y(_abc_42016_n3903) );
  NAND2X1 NAND2X1_348 ( .A(regfil_4__2_), .B(_abc_42016_n1047_1), .Y(_abc_42016_n3906) );
  NAND2X1 NAND2X1_349 ( .A(_abc_42016_n842), .B(_abc_42016_n3898), .Y(_abc_42016_n3947) );
  NAND2X1 NAND2X1_35 ( .A(regfil_5__4_), .B(_abc_42016_n696), .Y(_abc_42016_n868) );
  NAND2X1 NAND2X1_350 ( .A(_abc_42016_n3800), .B(_abc_42016_n909), .Y(_abc_42016_n3955) );
  NAND2X1 NAND2X1_351 ( .A(_abc_42016_n2150), .B(_abc_42016_n2152), .Y(_abc_42016_n3962) );
  NAND2X1 NAND2X1_352 ( .A(_abc_42016_n1031_1), .B(_abc_42016_n3963), .Y(_abc_42016_n3964) );
  NAND2X1 NAND2X1_353 ( .A(_abc_42016_n2183), .B(_abc_42016_n2185), .Y(_abc_42016_n3966) );
  NAND2X1 NAND2X1_354 ( .A(regfil_4__4_), .B(_abc_42016_n1047_1), .Y(_abc_42016_n3969) );
  NAND2X1 NAND2X1_355 ( .A(regfil_4__5_), .B(_abc_42016_n3933), .Y(_abc_42016_n3976) );
  NAND2X1 NAND2X1_356 ( .A(rdatahold_6_), .B(_abc_42016_n1019), .Y(_abc_42016_n3987) );
  NAND2X1 NAND2X1_357 ( .A(_abc_42016_n3990), .B(_abc_42016_n3991), .Y(_abc_42016_n3992) );
  NAND2X1 NAND2X1_358 ( .A(_abc_42016_n1031_1), .B(_abc_42016_n2176), .Y(_abc_42016_n3999) );
  NAND2X1 NAND2X1_359 ( .A(_abc_42016_n4016), .B(_abc_42016_n2210), .Y(_abc_42016_n4019) );
  NAND2X1 NAND2X1_36 ( .A(_abc_42016_n874), .B(_abc_42016_n866), .Y(_abc_42016_n877) );
  NAND2X1 NAND2X1_360 ( .A(_abc_42016_n4021), .B(_abc_42016_n2177), .Y(_abc_42016_n4022) );
  NAND2X1 NAND2X1_361 ( .A(_abc_42016_n561), .B(_abc_42016_n4026), .Y(_abc_42016_n4027) );
  NAND2X1 NAND2X1_362 ( .A(_abc_42016_n4029), .B(_abc_42016_n2143_1), .Y(_abc_42016_n4032) );
  NAND2X1 NAND2X1_363 ( .A(_abc_42016_n4031), .B(_abc_42016_n4032), .Y(_abc_42016_n4033) );
  NAND2X1 NAND2X1_364 ( .A(regfil_4__7_), .B(_abc_42016_n4000), .Y(_abc_42016_n4034) );
  NAND2X1 NAND2X1_365 ( .A(_abc_42016_n1554), .B(_abc_42016_n3958), .Y(_abc_42016_n4039) );
  NAND2X1 NAND2X1_366 ( .A(_abc_42016_n4053), .B(_abc_42016_n4054), .Y(_abc_42016_n4055) );
  NAND2X1 NAND2X1_367 ( .A(_abc_42016_n4070), .B(_abc_42016_n4062), .Y(_abc_42016_n4071) );
  NAND2X1 NAND2X1_368 ( .A(_abc_42016_n4012), .B(_abc_42016_n4073), .Y(_abc_36783_n4538) );
  NAND2X1 NAND2X1_369 ( .A(_abc_42016_n2286), .B(_abc_42016_n2284), .Y(_abc_42016_n4075) );
  NAND2X1 NAND2X1_37 ( .A(regfil_0__5_), .B(_abc_42016_n883), .Y(_abc_42016_n885) );
  NAND2X1 NAND2X1_370 ( .A(_abc_42016_n4103), .B(_abc_42016_n4112), .Y(_abc_42016_n4113) );
  NAND2X1 NAND2X1_371 ( .A(_abc_42016_n2526), .B(_abc_42016_n4113), .Y(_abc_42016_n4124) );
  NAND2X1 NAND2X1_372 ( .A(_abc_42016_n4142), .B(_abc_42016_n1841), .Y(_abc_42016_n4143) );
  NAND2X1 NAND2X1_373 ( .A(_abc_42016_n4160), .B(_abc_42016_n1385), .Y(_abc_42016_n4161) );
  NAND2X1 NAND2X1_374 ( .A(_abc_42016_n1841), .B(_abc_42016_n4173), .Y(_abc_42016_n4174) );
  NAND2X1 NAND2X1_375 ( .A(_abc_42016_n4186), .B(_abc_42016_n1387), .Y(_abc_42016_n4187) );
  NAND2X1 NAND2X1_376 ( .A(_abc_42016_n1841), .B(_abc_42016_n4200), .Y(_abc_42016_n4201) );
  NAND2X1 NAND2X1_377 ( .A(_abc_42016_n547), .B(_abc_42016_n4219), .Y(_abc_42016_n4220) );
  NAND2X1 NAND2X1_378 ( .A(_abc_42016_n4224), .B(_abc_42016_n1392), .Y(_abc_42016_n4225) );
  NAND2X1 NAND2X1_379 ( .A(_abc_42016_n4237), .B(_abc_42016_n1424), .Y(_abc_42016_n4238) );
  NAND2X1 NAND2X1_38 ( .A(_abc_42016_n660), .B(_abc_42016_n885), .Y(_abc_42016_n886) );
  NAND2X1 NAND2X1_380 ( .A(_abc_42016_n4262), .B(_abc_42016_n1480), .Y(_abc_42016_n4263) );
  NAND2X1 NAND2X1_381 ( .A(_abc_42016_n4275), .B(_abc_42016_n1511), .Y(_abc_42016_n4276) );
  NAND2X1 NAND2X1_382 ( .A(_abc_42016_n4287), .B(_abc_42016_n1532), .Y(_abc_42016_n4288) );
  NAND2X1 NAND2X1_383 ( .A(_abc_42016_n4293), .B(_abc_42016_n4294), .Y(_abc_42016_n4295) );
  NAND2X1 NAND2X1_384 ( .A(_abc_42016_n1558), .B(_abc_42016_n4299), .Y(_abc_42016_n4300) );
  NAND2X1 NAND2X1_385 ( .A(_abc_42016_n547), .B(_abc_42016_n4210), .Y(_abc_42016_n4310) );
  NAND2X1 NAND2X1_386 ( .A(ei), .B(intr), .Y(_abc_42016_n4323) );
  NAND2X1 NAND2X1_387 ( .A(_abc_42016_n517), .B(_abc_42016_n2078), .Y(_abc_42016_n4330) );
  NAND2X1 NAND2X1_388 ( .A(_abc_42016_n517), .B(_abc_42016_n1017), .Y(_abc_42016_n4332) );
  NAND2X1 NAND2X1_389 ( .A(_abc_42016_n2030), .B(_abc_42016_n3457), .Y(_abc_42016_n4333) );
  NAND2X1 NAND2X1_39 ( .A(_abc_42016_n889_1), .B(_abc_42016_n888), .Y(_abc_42016_n890) );
  NAND2X1 NAND2X1_390 ( .A(_auto_iopadmap_cc_313_execute_46280), .B(_abc_42016_n529), .Y(_abc_42016_n4335) );
  NAND2X1 NAND2X1_391 ( .A(_abc_42016_n517), .B(_abc_42016_n1872), .Y(_abc_42016_n4337) );
  NAND2X1 NAND2X1_392 ( .A(opcode_4_), .B(_abc_42016_n4050), .Y(_abc_42016_n4345) );
  NAND2X1 NAND2X1_393 ( .A(_abc_42016_n559), .B(_abc_42016_n1911), .Y(_abc_42016_n4346) );
  NAND2X1 NAND2X1_394 ( .A(alu_res_1_), .B(_abc_42016_n4057), .Y(_abc_42016_n4359) );
  NAND2X1 NAND2X1_395 ( .A(alu_res_2_), .B(_abc_42016_n4057), .Y(_abc_42016_n4374) );
  NAND2X1 NAND2X1_396 ( .A(alu_res_3_), .B(_abc_42016_n4057), .Y(_abc_42016_n4389) );
  NAND2X1 NAND2X1_397 ( .A(_abc_42016_n1454), .B(_abc_42016_n1427), .Y(_abc_42016_n4393) );
  NAND2X1 NAND2X1_398 ( .A(_abc_42016_n2066), .B(_abc_42016_n4350), .Y(_abc_42016_n4405) );
  NAND2X1 NAND2X1_399 ( .A(rdatahold_6_), .B(_abc_42016_n4382), .Y(_abc_42016_n4431_1) );
  NAND2X1 NAND2X1_4 ( .A(_abc_42016_n609), .B(_abc_42016_n616), .Y(_abc_42016_n617) );
  NAND2X1 NAND2X1_40 ( .A(alu_res_5_), .B(_abc_42016_n552), .Y(_abc_42016_n904) );
  NAND2X1 NAND2X1_400 ( .A(_abc_42016_n960), .B(_abc_42016_n4052), .Y(_abc_42016_n4441) );
  NAND2X1 NAND2X1_401 ( .A(_abc_42016_n531), .B(_abc_42016_n628), .Y(_abc_42016_n4449) );
  NAND2X1 NAND2X1_402 ( .A(_abc_42016_n512), .B(_abc_42016_n2260), .Y(_abc_42016_n4458) );
  NAND2X1 NAND2X1_403 ( .A(_abc_42016_n4551), .B(_abc_42016_n4550), .Y(_abc_42016_n4552) );
  NAND2X1 NAND2X1_404 ( .A(_abc_42016_n4578), .B(_abc_42016_n4550), .Y(_abc_42016_n4593) );
  NAND2X1 NAND2X1_405 ( .A(_abc_42016_n4323), .B(_abc_42016_n512), .Y(_abc_42016_n4604) );
  NAND2X1 NAND2X1_406 ( .A(_abc_42016_n4549), .B(_abc_42016_n4553), .Y(_abc_42016_n4611) );
  NAND2X1 NAND2X1_407 ( .A(_abc_42016_n4580), .B(_abc_42016_n4551), .Y(_abc_42016_n4614) );
  NAND2X1 NAND2X1_408 ( .A(_abc_42016_n4615_1), .B(_abc_42016_n4550), .Y(_abc_42016_n4616) );
  NAND2X1 NAND2X1_409 ( .A(_abc_42016_n4626), .B(_abc_42016_n4559), .Y(_abc_42016_n4627) );
  NAND2X1 NAND2X1_41 ( .A(_abc_42016_n913), .B(_abc_42016_n887), .Y(_abc_42016_n914) );
  NAND2X1 NAND2X1_410 ( .A(opcode_3_), .B(_abc_42016_n4640), .Y(_abc_42016_n4641) );
  NAND2X1 NAND2X1_411 ( .A(opcode_5_), .B(_abc_42016_n2056), .Y(_abc_42016_n4643) );
  NAND2X1 NAND2X1_412 ( .A(_abc_42016_n4648), .B(_abc_42016_n4652), .Y(_abc_42016_n4653) );
  NAND2X1 NAND2X1_413 ( .A(_abc_42016_n2369), .B(_abc_42016_n2364), .Y(_abc_42016_n4657_1) );
  NAND2X1 NAND2X1_414 ( .A(_abc_42016_n2450_1), .B(_abc_42016_n4661_1), .Y(_abc_42016_n4662) );
  NAND2X1 NAND2X1_415 ( .A(_abc_42016_n2369), .B(_abc_42016_n4664), .Y(_abc_42016_n4665) );
  NAND2X1 NAND2X1_416 ( .A(_abc_42016_n4677), .B(_abc_42016_n4559), .Y(_abc_42016_n4687) );
  NAND2X1 NAND2X1_417 ( .A(_abc_42016_n4689_1), .B(_abc_42016_n4687), .Y(_abc_42016_n4690) );
  NAND2X1 NAND2X1_418 ( .A(_abc_42016_n4709), .B(_abc_42016_n4684_1), .Y(_abc_42016_n4710) );
  NAND2X1 NAND2X1_419 ( .A(_abc_42016_n4570_1), .B(_abc_42016_n4594), .Y(_abc_42016_n4712) );
  NAND2X1 NAND2X1_42 ( .A(_abc_42016_n915), .B(_abc_42016_n914), .Y(_abc_42016_n916) );
  NAND2X1 NAND2X1_420 ( .A(_abc_42016_n4625), .B(_abc_42016_n4715), .Y(_abc_42016_n4716) );
  NAND2X1 NAND2X1_421 ( .A(_abc_42016_n4722), .B(_abc_42016_n4572), .Y(_abc_42016_n4723_1) );
  NAND2X1 NAND2X1_422 ( .A(_abc_42016_n4584), .B(_abc_42016_n4550), .Y(_abc_42016_n4726) );
  NAND2X1 NAND2X1_423 ( .A(alu_oprb_1_), .B(alu_opra_1_), .Y(alu__abc_41682_n42) );
  NAND2X1 NAND2X1_424 ( .A(alu_oprb_0_), .B(alu_opra_0_), .Y(alu__abc_41682_n43) );
  NAND2X1 NAND2X1_425 ( .A(alu_oprb_3_), .B(alu__abc_41682_n48), .Y(alu__abc_41682_n49) );
  NAND2X1 NAND2X1_426 ( .A(alu_opra_3_), .B(alu__abc_41682_n50_1), .Y(alu__abc_41682_n51) );
  NAND2X1 NAND2X1_427 ( .A(alu__abc_41682_n49), .B(alu__abc_41682_n51), .Y(alu__abc_41682_n52) );
  NAND2X1 NAND2X1_428 ( .A(alu_oprb_2_), .B(alu_opra_2_), .Y(alu__abc_41682_n53) );
  NAND2X1 NAND2X1_429 ( .A(alu_oprb_4_), .B(alu_opra_4_), .Y(alu__abc_41682_n60) );
  NAND2X1 NAND2X1_43 ( .A(alu_res_6_), .B(_abc_42016_n552), .Y(_abc_42016_n917) );
  NAND2X1 NAND2X1_430 ( .A(alu__abc_41682_n44), .B(alu__abc_41682_n41), .Y(alu__abc_41682_n65) );
  NAND2X1 NAND2X1_431 ( .A(alu_oprb_3_), .B(alu_opra_3_), .Y(alu__abc_41682_n66) );
  NAND2X1 NAND2X1_432 ( .A(alu_oprb_5_), .B(alu_opra_5_), .Y(alu__abc_41682_n75) );
  NAND2X1 NAND2X1_433 ( .A(alu__abc_41682_n75), .B(alu__abc_41682_n74), .Y(alu__abc_41682_n76) );
  NAND2X1 NAND2X1_434 ( .A(alu__abc_41682_n60), .B(alu__abc_41682_n68), .Y(alu__abc_41682_n78) );
  NAND2X1 NAND2X1_435 ( .A(alu__abc_41682_n77), .B(alu__abc_41682_n78), .Y(alu__abc_41682_n79) );
  NAND2X1 NAND2X1_436 ( .A(alu__abc_41682_n89), .B(alu__abc_41682_n91), .Y(alu__abc_41682_n92) );
  NAND2X1 NAND2X1_437 ( .A(alu_oprb_0_), .B(alu__abc_41682_n139), .Y(alu__abc_41682_n163) );
  NAND2X1 NAND2X1_438 ( .A(alu__abc_41682_n148), .B(alu__abc_41682_n133), .Y(alu__abc_41682_n177) );
  NAND2X1 NAND2X1_439 ( .A(alu__abc_41682_n149), .B(alu__abc_41682_n178), .Y(alu__abc_41682_n179) );
  NAND2X1 NAND2X1_44 ( .A(_abc_42016_n536), .B(_abc_42016_n920), .Y(_abc_42016_n921) );
  NAND2X1 NAND2X1_440 ( .A(alu_sel_1_), .B(alu__abc_41682_n180), .Y(alu__abc_41682_n181) );
  NAND2X1 NAND2X1_441 ( .A(alu__abc_41682_n156), .B(alu__abc_41682_n130), .Y(alu__abc_41682_n188) );
  NAND2X1 NAND2X1_442 ( .A(alu__abc_41682_n153), .B(alu__abc_41682_n184), .Y(alu__abc_41682_n193) );
  NAND2X1 NAND2X1_443 ( .A(alu__abc_41682_n195), .B(alu__abc_41682_n192), .Y(alu__abc_41682_n196) );
  NAND2X1 NAND2X1_444 ( .A(alu__abc_41682_n202), .B(alu__abc_41682_n36), .Y(alu__abc_41682_n203) );
  NAND2X1 NAND2X1_445 ( .A(alu__abc_41682_n150), .B(alu__abc_41682_n210), .Y(alu__abc_41682_n211) );
  NAND2X1 NAND2X1_446 ( .A(alu__abc_41682_n146), .B(alu__abc_41682_n151), .Y(alu__abc_41682_n214) );
  NAND2X1 NAND2X1_447 ( .A(alu__abc_41682_n144), .B(alu__abc_41682_n160), .Y(alu__abc_41682_n215) );
  NAND2X1 NAND2X1_448 ( .A(alu_sel_2_), .B(alu__abc_41682_n184), .Y(alu__abc_41682_n218) );
  NAND2X1 NAND2X1_449 ( .A(alu__abc_41682_n226), .B(alu__abc_41682_n196), .Y(alu__abc_41682_n227) );
  NAND2X1 NAND2X1_45 ( .A(_abc_42016_n917), .B(_abc_42016_n928), .Y(_abc_42016_n929) );
  NAND2X1 NAND2X1_450 ( .A(alu__abc_41682_n68), .B(alu__abc_41682_n228), .Y(alu__abc_41682_n229) );
  NAND2X1 NAND2X1_451 ( .A(alu__abc_41682_n52), .B(alu__abc_41682_n55), .Y(alu__abc_41682_n236) );
  NAND2X1 NAND2X1_452 ( .A(alu__abc_41682_n180), .B(alu__abc_41682_n263), .Y(alu__abc_41682_n264) );
  NAND2X1 NAND2X1_453 ( .A(alu__abc_41682_n65), .B(alu__abc_41682_n233), .Y(alu__abc_41682_n273_1) );
  NAND2X1 NAND2X1_454 ( .A(alu__abc_41682_n278), .B(alu__abc_41682_n281), .Y(alu__abc_41682_n282) );
  NAND2X1 NAND2X1_455 ( .A(alu__abc_41682_n206), .B(alu__abc_41682_n284), .Y(alu__abc_41682_n285) );
  NAND2X1 NAND2X1_456 ( .A(alu__abc_41682_n276), .B(alu__abc_41682_n286_1), .Y(alu__abc_41682_n287) );
  NAND2X1 NAND2X1_457 ( .A(alu__abc_41682_n36), .B(alu__abc_41682_n240), .Y(alu__abc_41682_n296) );
  NAND2X1 NAND2X1_458 ( .A(alu_cin), .B(alu__abc_41682_n39), .Y(alu__abc_41682_n299) );
  NAND2X1 NAND2X1_459 ( .A(alu__abc_41682_n184), .B(alu__abc_41682_n37), .Y(alu__abc_41682_n304) );
  NAND2X1 NAND2X1_46 ( .A(_abc_42016_n930), .B(_abc_42016_n933), .Y(_abc_42016_n934) );
  NAND2X1 NAND2X1_460 ( .A(alu__abc_41682_n317), .B(alu__abc_41682_n313), .Y(alu__abc_41682_n318) );
  NAND2X1 NAND2X1_461 ( .A(alu__abc_41682_n248), .B(alu__abc_41682_n257), .Y(alu__abc_41682_n321) );
  NAND2X1 NAND2X1_462 ( .A(alu__abc_41682_n320), .B(alu__abc_41682_n321), .Y(alu__abc_41682_n322) );
  NAND2X1 NAND2X1_463 ( .A(alu__abc_41682_n323), .B(alu__abc_41682_n324), .Y(alu__abc_41682_n325) );
  NAND2X1 NAND2X1_464 ( .A(alu__abc_41682_n326), .B(alu__abc_41682_n319), .Y(alu__abc_41682_n327) );
  NAND2X1 NAND2X1_465 ( .A(alu__abc_41682_n332), .B(alu__abc_41682_n331), .Y(alu__abc_41682_n333) );
  NAND2X1 NAND2X1_466 ( .A(alu__abc_41682_n328), .B(alu__abc_41682_n334), .Y(alu_parity) );
  NAND2X1 NAND2X1_467 ( .A(alu_sel_1_), .B(alu__abc_41682_n178), .Y(alu__abc_41682_n339) );
  NAND2X1 NAND2X1_468 ( .A(alu__abc_41682_n339), .B(alu__abc_41682_n287), .Y(alu__abc_41682_n342) );
  NAND2X1 NAND2X1_469 ( .A(alu__abc_41682_n339), .B(alu__abc_41682_n246), .Y(alu__abc_41682_n346) );
  NAND2X1 NAND2X1_47 ( .A(regfil_3__6_), .B(_abc_42016_n937), .Y(_abc_42016_n938) );
  NAND2X1 NAND2X1_470 ( .A(alu__abc_41682_n339), .B(alu__abc_41682_n224), .Y(alu__abc_41682_n349) );
  NAND2X1 NAND2X1_471 ( .A(alu__abc_41682_n339), .B(alu_sout), .Y(alu__abc_41682_n351) );
  NAND2X1 NAND2X1_472 ( .A(alu__abc_41682_n150), .B(alu__abc_41682_n209), .Y(alu__abc_41682_n355) );
  NAND2X1 NAND2X1_48 ( .A(_abc_42016_n940), .B(_abc_42016_n938), .Y(_abc_42016_n941_1) );
  NAND2X1 NAND2X1_49 ( .A(regfil_0__7_), .B(_abc_42016_n952), .Y(_abc_42016_n953) );
  NAND2X1 NAND2X1_5 ( .A(_abc_42016_n608), .B(_abc_42016_n618), .Y(_abc_42016_n619) );
  NAND2X1 NAND2X1_50 ( .A(_abc_42016_n536), .B(_abc_42016_n965), .Y(_abc_42016_n966) );
  NAND2X1 NAND2X1_51 ( .A(_abc_42016_n974), .B(_abc_42016_n943), .Y(_abc_42016_n976) );
  NAND2X1 NAND2X1_52 ( .A(regfil_5__7_), .B(_abc_42016_n696), .Y(_abc_42016_n983) );
  NAND2X1 NAND2X1_53 ( .A(_abc_42016_n1007), .B(_abc_42016_n1002), .Y(_abc_42016_n1008) );
  NAND2X1 NAND2X1_54 ( .A(_abc_42016_n997), .B(_abc_42016_n1009), .Y(_abc_42016_n1010) );
  NAND2X1 NAND2X1_55 ( .A(_abc_42016_n543), .B(_abc_42016_n1013), .Y(_abc_42016_n1014) );
  NAND2X1 NAND2X1_56 ( .A(_abc_42016_n512), .B(_abc_42016_n1017), .Y(_abc_42016_n1018) );
  NAND2X1 NAND2X1_57 ( .A(regfil_5__0_), .B(sp_0_), .Y(_abc_42016_n1024) );
  NAND2X1 NAND2X1_58 ( .A(regfil_1__0_), .B(regfil_5__0_), .Y(_abc_42016_n1028) );
  NAND2X1 NAND2X1_59 ( .A(_abc_42016_n1000), .B(_abc_42016_n561), .Y(_abc_42016_n1030) );
  NAND2X1 NAND2X1_6 ( .A(alu_res_0_), .B(_abc_42016_n552), .Y(_abc_42016_n638) );
  NAND2X1 NAND2X1_60 ( .A(_abc_42016_n634), .B(_abc_42016_n695), .Y(_abc_42016_n1032) );
  NAND2X1 NAND2X1_61 ( .A(regfil_3__0_), .B(regfil_5__0_), .Y(_abc_42016_n1033) );
  NAND2X1 NAND2X1_62 ( .A(_abc_42016_n1042), .B(_abc_42016_n1039), .Y(_abc_42016_n1043) );
  NAND2X1 NAND2X1_63 ( .A(regfil_5__1_), .B(sp_1_), .Y(_abc_42016_n1069) );
  NAND2X1 NAND2X1_64 ( .A(_abc_42016_n1088), .B(_abc_42016_n1059), .Y(_abc_42016_n1089) );
  NAND2X1 NAND2X1_65 ( .A(regfil_3__1_), .B(regfil_5__1_), .Y(_abc_42016_n1099) );
  NAND2X1 NAND2X1_66 ( .A(regfil_1__1_), .B(regfil_5__1_), .Y(_abc_42016_n1106_1) );
  NAND2X1 NAND2X1_67 ( .A(_abc_42016_n1107_1), .B(_abc_42016_n1108), .Y(_abc_42016_n1109) );
  NAND2X1 NAND2X1_68 ( .A(_abc_42016_n1114_1), .B(_abc_42016_n1115), .Y(_abc_42016_n1117) );
  NAND2X1 NAND2X1_69 ( .A(_abc_42016_n1117), .B(_abc_42016_n1116), .Y(_abc_42016_n1118) );
  NAND2X1 NAND2X1_7 ( .A(regfil_1__2_), .B(_abc_42016_n646), .Y(_abc_42016_n647) );
  NAND2X1 NAND2X1_70 ( .A(regfil_5__2_), .B(_abc_42016_n1063), .Y(_abc_42016_n1120) );
  NAND2X1 NAND2X1_71 ( .A(_abc_42016_n1121_1), .B(_abc_42016_n1120), .Y(_abc_42016_n1122) );
  NAND2X1 NAND2X1_72 ( .A(_abc_42016_n757), .B(_abc_42016_n1062), .Y(_abc_42016_n1126) );
  NAND2X1 NAND2X1_73 ( .A(_abc_42016_n1139), .B(_abc_42016_n1120), .Y(_abc_42016_n1141) );
  NAND2X1 NAND2X1_74 ( .A(regfil_3__3_), .B(regfil_5__3_), .Y(_abc_42016_n1143) );
  NAND2X1 NAND2X1_75 ( .A(_abc_42016_n795), .B(_abc_42016_n1139), .Y(_abc_42016_n1144) );
  NAND2X1 NAND2X1_76 ( .A(_abc_42016_n643_1), .B(_abc_42016_n1139), .Y(_abc_42016_n1153) );
  NAND2X1 NAND2X1_77 ( .A(regfil_1__3_), .B(regfil_5__3_), .Y(_abc_42016_n1154) );
  NAND2X1 NAND2X1_78 ( .A(_abc_42016_n1154), .B(_abc_42016_n1153), .Y(_abc_42016_n1155) );
  NAND2X1 NAND2X1_79 ( .A(regfil_5__3_), .B(sp_3_), .Y(_abc_42016_n1163) );
  NAND2X1 NAND2X1_8 ( .A(regfil_1__6_), .B(_abc_42016_n650), .Y(_abc_42016_n651_1) );
  NAND2X1 NAND2X1_80 ( .A(_abc_42016_n1163), .B(_abc_42016_n1162), .Y(_abc_42016_n1166) );
  NAND2X1 NAND2X1_81 ( .A(_abc_42016_n1179), .B(_abc_42016_n993), .Y(_abc_42016_n1180) );
  NAND2X1 NAND2X1_82 ( .A(_abc_42016_n843), .B(_abc_42016_n1183), .Y(_abc_42016_n1184) );
  NAND2X1 NAND2X1_83 ( .A(_abc_42016_n1182), .B(_abc_42016_n1184), .Y(_abc_42016_n1185) );
  NAND2X1 NAND2X1_84 ( .A(_abc_42016_n1189), .B(_abc_42016_n1188), .Y(_abc_42016_n1190) );
  NAND2X1 NAND2X1_85 ( .A(_abc_42016_n610), .B(_abc_42016_n843), .Y(_abc_42016_n1192) );
  NAND2X1 NAND2X1_86 ( .A(regfil_1__4_), .B(regfil_5__4_), .Y(_abc_42016_n1193) );
  NAND2X1 NAND2X1_87 ( .A(regfil_1__2_), .B(regfil_5__2_), .Y(_abc_42016_n1195) );
  NAND2X1 NAND2X1_88 ( .A(_abc_42016_n1198), .B(_abc_42016_n1199_1), .Y(_abc_42016_n1200) );
  NAND2X1 NAND2X1_89 ( .A(_abc_42016_n1203), .B(_abc_42016_n1202), .Y(_abc_42016_n1204) );
  NAND2X1 NAND2X1_9 ( .A(_abc_42016_n570), .B(_abc_42016_n573), .Y(_abc_42016_n656) );
  NAND2X1 NAND2X1_90 ( .A(regfil_5__2_), .B(sp_2_), .Y(_abc_42016_n1213) );
  NAND2X1 NAND2X1_91 ( .A(_abc_42016_n1232), .B(_abc_42016_n1234), .Y(_abc_42016_n1235) );
  NAND2X1 NAND2X1_92 ( .A(regfil_3__4_), .B(regfil_5__4_), .Y(_abc_42016_n1241) );
  NAND2X1 NAND2X1_93 ( .A(_abc_42016_n1245), .B(_abc_42016_n998), .Y(_abc_42016_n1246) );
  NAND2X1 NAND2X1_94 ( .A(_abc_42016_n1008), .B(_abc_42016_n1286), .Y(_abc_42016_n1287) );
  NAND2X1 NAND2X1_95 ( .A(regfil_5__6_), .B(_abc_42016_n1226), .Y(_abc_42016_n1290) );
  NAND2X1 NAND2X1_96 ( .A(_abc_42016_n1290), .B(_abc_42016_n1138), .Y(_abc_42016_n1291) );
  NAND2X1 NAND2X1_97 ( .A(_abc_42016_n923), .B(_abc_42016_n1251), .Y(_abc_42016_n1295) );
  NAND2X1 NAND2X1_98 ( .A(regfil_1__6_), .B(regfil_5__6_), .Y(_abc_42016_n1305) );
  NAND2X1 NAND2X1_99 ( .A(regfil_3__6_), .B(regfil_5__6_), .Y(_abc_42016_n1313) );
  NAND3X1 NAND3X1_1 ( .A(_abc_42016_n652), .B(_abc_42016_n660), .C(_abc_42016_n655_1), .Y(_abc_42016_n661_1) );
  NAND3X1 NAND3X1_10 ( .A(_abc_42016_n1032), .B(_abc_42016_n1033), .C(_abc_42016_n1031_1), .Y(_abc_42016_n1034) );
  NAND3X1 NAND3X1_100 ( .A(_abc_42016_n3502), .B(_abc_42016_n3694), .C(_abc_42016_n3695), .Y(_abc_42016_n3708) );
  NAND3X1 NAND3X1_101 ( .A(_abc_42016_n2256), .B(_abc_42016_n3737), .C(_abc_42016_n3739), .Y(_abc_42016_n3740) );
  NAND3X1 NAND3X1_102 ( .A(_abc_42016_n559), .B(_abc_42016_n3740), .C(_abc_42016_n3743), .Y(_abc_42016_n3744) );
  NAND3X1 NAND3X1_103 ( .A(_abc_42016_n3750), .B(_abc_42016_n3751), .C(_abc_42016_n3744), .Y(_abc_42016_n3752) );
  NAND3X1 NAND3X1_104 ( .A(_abc_42016_n3753), .B(_abc_42016_n3754), .C(_abc_42016_n3752), .Y(_abc_42016_n3755_1) );
  NAND3X1 NAND3X1_105 ( .A(_abc_42016_n559), .B(_abc_42016_n3760), .C(_abc_42016_n3766), .Y(_abc_42016_n3767) );
  NAND3X1 NAND3X1_106 ( .A(_abc_42016_n3772), .B(_abc_42016_n3773), .C(_abc_42016_n3767), .Y(_abc_42016_n3774) );
  NAND3X1 NAND3X1_107 ( .A(_abc_42016_n2129), .B(_abc_42016_n2126), .C(_abc_42016_n3842), .Y(_abc_42016_n3843) );
  NAND3X1 NAND3X1_108 ( .A(_abc_42016_n1023), .B(_abc_42016_n3844), .C(_abc_42016_n3843), .Y(_abc_42016_n3845) );
  NAND3X1 NAND3X1_109 ( .A(_abc_42016_n2156), .B(_abc_42016_n2158), .C(_abc_42016_n3910), .Y(_abc_42016_n3911) );
  NAND3X1 NAND3X1_11 ( .A(_abc_42016_n1045), .B(_abc_42016_n1040), .C(_abc_42016_n1049), .Y(_abc_42016_n1050) );
  NAND3X1 NAND3X1_110 ( .A(_abc_42016_n1031_1), .B(_abc_42016_n3911), .C(_abc_42016_n3913), .Y(_abc_42016_n3914) );
  NAND3X1 NAND3X1_111 ( .A(_abc_42016_n3905), .B(_abc_42016_n3906), .C(_abc_42016_n3919), .Y(_abc_42016_n3920) );
  NAND3X1 NAND3X1_112 ( .A(_abc_42016_n3941), .B(_abc_42016_n3938), .C(_abc_42016_n3944), .Y(_abc_42016_n3945) );
  NAND3X1 NAND3X1_113 ( .A(_abc_42016_n3969), .B(_abc_42016_n3968), .C(_abc_42016_n3964), .Y(_abc_42016_n3970) );
  NAND3X1 NAND3X1_114 ( .A(_abc_42016_n1036), .B(_abc_42016_n2209), .C(_abc_42016_n3992), .Y(_abc_42016_n3993) );
  NAND3X1 NAND3X1_115 ( .A(_abc_42016_n3986), .B(_abc_42016_n3987), .C(_abc_42016_n4009), .Y(_abc_36783_n4537) );
  NAND3X1 NAND3X1_116 ( .A(_abc_42016_n2180), .B(_abc_42016_n4017), .C(_abc_42016_n2209), .Y(_abc_42016_n4018) );
  NAND3X1 NAND3X1_117 ( .A(_abc_42016_n1036), .B(_abc_42016_n4018), .C(_abc_42016_n4019), .Y(_abc_42016_n4020) );
  NAND3X1 NAND3X1_118 ( .A(_abc_42016_n2148), .B(_abc_42016_n4023), .C(_abc_42016_n2176), .Y(_abc_42016_n4024) );
  NAND3X1 NAND3X1_119 ( .A(_abc_42016_n1031_1), .B(_abc_42016_n4024), .C(_abc_42016_n4022), .Y(_abc_42016_n4025) );
  NAND3X1 NAND3X1_12 ( .A(_abc_42016_n1109), .B(_abc_42016_n1110_1), .C(_abc_42016_n1001_1), .Y(_abc_42016_n1111_1) );
  NAND3X1 NAND3X1_120 ( .A(_abc_42016_n4020), .B(_abc_42016_n4027), .C(_abc_42016_n4025), .Y(_abc_42016_n4028) );
  NAND3X1 NAND3X1_121 ( .A(_abc_42016_n2104), .B(_abc_42016_n4030), .C(_abc_42016_n2142), .Y(_abc_42016_n4031) );
  NAND3X1 NAND3X1_122 ( .A(_abc_42016_n4051), .B(_abc_42016_n4060), .C(_abc_42016_n4058), .Y(_abc_42016_n4061) );
  NAND3X1 NAND3X1_123 ( .A(_abc_42016_n2256), .B(_abc_42016_n4083), .C(_abc_42016_n4084), .Y(_abc_42016_n4085) );
  NAND3X1 NAND3X1_124 ( .A(_abc_42016_n1046), .B(_abc_42016_n1380), .C(_abc_42016_n4091), .Y(_abc_42016_n4092_1) );
  NAND3X1 NAND3X1_125 ( .A(_abc_42016_n574), .B(_abc_42016_n2322), .C(_abc_42016_n2256), .Y(_abc_42016_n4102) );
  NAND3X1 NAND3X1_126 ( .A(_abc_42016_n671_1), .B(_abc_42016_n1061), .C(_abc_42016_n1035), .Y(_abc_42016_n4104) );
  NAND3X1 NAND3X1_127 ( .A(_abc_42016_n4078), .B(_abc_42016_n4109), .C(_abc_42016_n4107), .Y(_abc_42016_n4110) );
  NAND3X1 NAND3X1_128 ( .A(_abc_42016_n4147), .B(_abc_42016_n4148), .C(_abc_42016_n4149), .Y(_abc_42016_n4150_1) );
  NAND3X1 NAND3X1_129 ( .A(_abc_42016_n531), .B(_abc_42016_n561), .C(_abc_42016_n2095), .Y(_abc_42016_n4352) );
  NAND3X1 NAND3X1_13 ( .A(_abc_42016_n561), .B(_abc_42016_n1010), .C(_abc_42016_n1128), .Y(_abc_42016_n1129) );
  NAND3X1 NAND3X1_130 ( .A(_abc_42016_n4356), .B(_abc_42016_n4357), .C(_abc_42016_n4342), .Y(_abc_36783_n4579) );
  NAND3X1 NAND3X1_131 ( .A(_abc_42016_n4376), .B(_abc_42016_n4385), .C(_abc_42016_n4373), .Y(_abc_36783_n4581) );
  NAND3X1 NAND3X1_132 ( .A(_abc_42016_n4391), .B(_abc_42016_n4400), .C(_abc_42016_n4388), .Y(_abc_36783_n4582) );
  NAND3X1 NAND3X1_133 ( .A(_abc_42016_n4433), .B(_abc_42016_n4437), .C(_abc_42016_n4430), .Y(_abc_42016_n4438) );
  NAND3X1 NAND3X1_134 ( .A(_abc_42016_n2218), .B(_abc_42016_n4441), .C(_abc_42016_n4056), .Y(_abc_42016_n4442) );
  NAND3X1 NAND3X1_135 ( .A(_abc_42016_n1860), .B(_abc_42016_n679), .C(_abc_42016_n4063), .Y(_abc_42016_n4447_1) );
  NAND3X1 NAND3X1_136 ( .A(_abc_42016_n4600_1), .B(_abc_42016_n4608), .C(_abc_42016_n4576), .Y(_abc_42016_n4609) );
  NAND3X1 NAND3X1_137 ( .A(_abc_42016_n2363), .B(_abc_42016_n2408_1), .C(_abc_42016_n2450_1), .Y(_abc_42016_n4613) );
  NAND3X1 NAND3X1_138 ( .A(_abc_42016_n4618), .B(_abc_42016_n4619), .C(_abc_42016_n4616), .Y(_abc_42016_n4620) );
  NAND3X1 NAND3X1_139 ( .A(_abc_42016_n2230), .B(_abc_42016_n4628), .C(_abc_42016_n4627), .Y(_abc_42016_n4629) );
  NAND3X1 NAND3X1_14 ( .A(_abc_42016_n1140), .B(_abc_42016_n1141), .C(_abc_42016_n1138), .Y(_abc_42016_n1142) );
  NAND3X1 NAND3X1_140 ( .A(_abc_42016_n4103), .B(_abc_42016_n4105), .C(_abc_42016_n4634), .Y(_abc_42016_n4635) );
  NAND3X1 NAND3X1_141 ( .A(_abc_42016_n4622), .B(_abc_42016_n4625), .C(_abc_42016_n4637), .Y(_abc_42016_n4638) );
  NAND3X1 NAND3X1_142 ( .A(_abc_42016_n1061), .B(_abc_42016_n1374), .C(_abc_42016_n4650_1), .Y(_abc_42016_n4651) );
  NAND3X1 NAND3X1_143 ( .A(_abc_42016_n2259), .B(_abc_42016_n4578), .C(_abc_42016_n4655), .Y(_abc_42016_n4663) );
  NAND3X1 NAND3X1_144 ( .A(_abc_42016_n4659), .B(_abc_42016_n4662), .C(_abc_42016_n4666_1), .Y(_abc_42016_n4667) );
  NAND3X1 NAND3X1_145 ( .A(_abc_42016_n4654_1), .B(_abc_42016_n4670_1), .C(_abc_42016_n4668_1), .Y(_abc_42016_n4671) );
  NAND3X1 NAND3X1_146 ( .A(_abc_42016_n4557), .B(_abc_42016_n4569), .C(_abc_42016_n4679), .Y(_abc_42016_n4680_1) );
  NAND3X1 NAND3X1_147 ( .A(_abc_42016_n4678_1), .B(_abc_42016_n4680_1), .C(_abc_42016_n4676_1), .Y(_abc_42016_n4681) );
  NAND3X1 NAND3X1_148 ( .A(_abc_42016_n2408_1), .B(_abc_42016_n4664), .C(_abc_42016_n4550), .Y(_abc_42016_n4685) );
  NAND3X1 NAND3X1_149 ( .A(_abc_42016_n4686), .B(_abc_42016_n4693), .C(_abc_42016_n4674_1), .Y(_abc_42016_n4694) );
  NAND3X1 NAND3X1_15 ( .A(_abc_42016_n1142), .B(_abc_42016_n1168), .C(_abc_42016_n1158), .Y(_abc_42016_n1169) );
  NAND3X1 NAND3X1_150 ( .A(_abc_42016_n4576), .B(_abc_42016_n4693), .C(_abc_42016_n4699), .Y(_abc_36783_n4645) );
  NAND3X1 NAND3X1_151 ( .A(_abc_42016_n4689_1), .B(_abc_42016_n4703), .C(_abc_42016_n4687), .Y(_abc_42016_n4704) );
  NAND3X1 NAND3X1_152 ( .A(_abc_42016_n4592), .B(_abc_42016_n4705_1), .C(_abc_42016_n4706), .Y(_abc_36783_n4646) );
  NAND3X1 NAND3X1_153 ( .A(_abc_42016_n4711_1), .B(_abc_42016_n4714), .C(_abc_42016_n4717_1), .Y(_abc_36783_n4647) );
  NAND3X1 NAND3X1_154 ( .A(_abc_42016_n3418), .B(_abc_42016_n4628), .C(_abc_42016_n4618), .Y(_abc_42016_n4719_1) );
  NAND3X1 NAND3X1_155 ( .A(_abc_42016_n4726), .B(_abc_42016_n4685), .C(_abc_42016_n4715), .Y(_abc_42016_n4727) );
  NAND3X1 NAND3X1_156 ( .A(_abc_42016_n4672_1), .B(_abc_42016_n4725_1), .C(_abc_42016_n4728), .Y(_abc_36783_n4648) );
  NAND3X1 NAND3X1_157 ( .A(_abc_42016_n4611), .B(_abc_42016_n4730), .C(_abc_42016_n4733), .Y(_abc_36783_n4649) );
  NAND3X1 NAND3X1_158 ( .A(alu_cin), .B(alu__abc_41682_n36), .C(alu__abc_41682_n39), .Y(alu__abc_41682_n40) );
  NAND3X1 NAND3X1_159 ( .A(alu__abc_41682_n53), .B(alu__abc_41682_n66), .C(alu__abc_41682_n65), .Y(alu__abc_41682_n67) );
  NAND3X1 NAND3X1_16 ( .A(_abc_42016_n1195), .B(_abc_42016_n1154), .C(_abc_42016_n1109), .Y(_abc_42016_n1196_1) );
  NAND3X1 NAND3X1_160 ( .A(alu__abc_41682_n62), .B(alu__abc_41682_n64), .C(alu__abc_41682_n67), .Y(alu__abc_41682_n68) );
  NAND3X1 NAND3X1_161 ( .A(alu__abc_41682_n60), .B(alu__abc_41682_n76), .C(alu__abc_41682_n68), .Y(alu__abc_41682_n80) );
  NAND3X1 NAND3X1_162 ( .A(alu__abc_41682_n79), .B(alu__abc_41682_n80), .C(alu__abc_41682_n72), .Y(alu__abc_41682_n81) );
  NAND3X1 NAND3X1_163 ( .A(alu__abc_41682_n75), .B(alu__abc_41682_n90), .C(alu__abc_41682_n79), .Y(alu__abc_41682_n91) );
  NAND3X1 NAND3X1_164 ( .A(alu__abc_41682_n94), .B(alu__abc_41682_n99), .C(alu__abc_41682_n89), .Y(alu__abc_41682_n101) );
  NAND3X1 NAND3X1_165 ( .A(alu__abc_41682_n94), .B(alu__abc_41682_n108), .C(alu__abc_41682_n89), .Y(alu__abc_41682_n109) );
  NAND3X1 NAND3X1_166 ( .A(alu__abc_41682_n107), .B(alu__abc_41682_n112), .C(alu__abc_41682_n103), .Y(alu__abc_41682_n113) );
  NAND3X1 NAND3X1_167 ( .A(alu__abc_41682_n136), .B(alu__abc_41682_n51), .C(alu__abc_41682_n142), .Y(alu__abc_41682_n143) );
  NAND3X1 NAND3X1_168 ( .A(alu__abc_41682_n49), .B(alu__abc_41682_n135), .C(alu__abc_41682_n143), .Y(alu__abc_41682_n144) );
  NAND3X1 NAND3X1_169 ( .A(alu__abc_41682_n99), .B(alu__abc_41682_n147), .C(alu__abc_41682_n146), .Y(alu__abc_41682_n148) );
  NAND3X1 NAND3X1_17 ( .A(_abc_42016_n1153), .B(_abc_42016_n1194), .C(_abc_42016_n1196_1), .Y(_abc_42016_n1197_1) );
  NAND3X1 NAND3X1_170 ( .A(alu__abc_41682_n88), .B(alu__abc_41682_n117), .C(alu__abc_41682_n130), .Y(alu__abc_41682_n151) );
  NAND3X1 NAND3X1_171 ( .A(alu__abc_41682_n150), .B(alu__abc_41682_n146), .C(alu__abc_41682_n151), .Y(alu__abc_41682_n152) );
  NAND3X1 NAND3X1_172 ( .A(alu__abc_41682_n77), .B(alu__abc_41682_n134), .C(alu__abc_41682_n144), .Y(alu__abc_41682_n156) );
  NAND3X1 NAND3X1_173 ( .A(alu__abc_41682_n155), .B(alu__abc_41682_n156), .C(alu__abc_41682_n130), .Y(alu__abc_41682_n157) );
  NAND3X1 NAND3X1_174 ( .A(alu__abc_41682_n51), .B(alu__abc_41682_n62), .C(alu__abc_41682_n128), .Y(alu__abc_41682_n160) );
  NAND3X1 NAND3X1_175 ( .A(alu__abc_41682_n124_1), .B(alu__abc_41682_n41), .C(alu__abc_41682_n126), .Y(alu__abc_41682_n166) );
  NAND3X1 NAND3X1_176 ( .A(alu__abc_41682_n136), .B(alu__abc_41682_n169_1), .C(alu__abc_41682_n142), .Y(alu__abc_41682_n170) );
  NAND3X1 NAND3X1_177 ( .A(alu__abc_41682_n168), .B(alu__abc_41682_n170), .C(alu__abc_41682_n167), .Y(alu__abc_41682_n171) );
  NAND3X1 NAND3X1_178 ( .A(alu__abc_41682_n157), .B(alu__abc_41682_n174), .C(alu__abc_41682_n152), .Y(alu__abc_41682_n175) );
  NAND3X1 NAND3X1_179 ( .A(alu__abc_41682_n133), .B(alu__abc_41682_n148), .C(alu__abc_41682_n175), .Y(alu__abc_41682_n176) );
  NAND3X1 NAND3X1_18 ( .A(_abc_42016_n1197_1), .B(_abc_42016_n1200), .C(_abc_42016_n1036), .Y(_abc_42016_n1201) );
  NAND3X1 NAND3X1_180 ( .A(alu__abc_41682_n150), .B(alu__abc_41682_n172), .C(alu__abc_41682_n188), .Y(alu__abc_41682_n189) );
  NAND3X1 NAND3X1_181 ( .A(alu__abc_41682_n176), .B(alu__abc_41682_n191), .C(alu__abc_41682_n113), .Y(alu__abc_41682_n192) );
  NAND3X1 NAND3X1_182 ( .A(alu__abc_41682_n136), .B(alu__abc_41682_n52), .C(alu__abc_41682_n142), .Y(alu__abc_41682_n207) );
  NAND3X1 NAND3X1_183 ( .A(alu__abc_41682_n159), .B(alu__abc_41682_n211), .C(alu__abc_41682_n157), .Y(alu__abc_41682_n212) );
  NAND3X1 NAND3X1_184 ( .A(alu__abc_41682_n146), .B(alu__abc_41682_n151), .C(alu__abc_41682_n212), .Y(alu__abc_41682_n213) );
  NAND3X1 NAND3X1_185 ( .A(alu__abc_41682_n150), .B(alu__abc_41682_n209), .C(alu__abc_41682_n215), .Y(alu__abc_41682_n216) );
  NAND3X1 NAND3X1_186 ( .A(alu__abc_41682_n195), .B(alu__abc_41682_n224), .C(alu__abc_41682_n192), .Y(alu__abc_41682_n225) );
  NAND3X1 NAND3X1_187 ( .A(alu__abc_41682_n65), .B(alu__abc_41682_n233), .C(alu__abc_41682_n232), .Y(alu__abc_41682_n234) );
  NAND3X1 NAND3X1_188 ( .A(alu__abc_41682_n68), .B(alu__abc_41682_n228), .C(alu__abc_41682_n237), .Y(alu__abc_41682_n238) );
  NAND3X1 NAND3X1_189 ( .A(alu__abc_41682_n107), .B(alu__abc_41682_n249), .C(alu__abc_41682_n81), .Y(alu__abc_41682_n250) );
  NAND3X1 NAND3X1_19 ( .A(_abc_42016_n1204), .B(_abc_42016_n1205), .C(_abc_42016_n1031_1), .Y(_abc_42016_n1206) );
  NAND3X1 NAND3X1_190 ( .A(alu__abc_41682_n130), .B(alu__abc_41682_n156), .C(alu__abc_41682_n173), .Y(alu__abc_41682_n251) );
  NAND3X1 NAND3X1_191 ( .A(alu__abc_41682_n250), .B(alu__abc_41682_n251), .C(alu__abc_41682_n256), .Y(alu__abc_41682_n257) );
  NAND3X1 NAND3X1_192 ( .A(alu__abc_41682_n248), .B(alu__abc_41682_n246), .C(alu__abc_41682_n257), .Y(alu__abc_41682_n259_1) );
  NAND3X1 NAND3X1_193 ( .A(alu__abc_41682_n47), .B(alu__abc_41682_n107), .C(alu__abc_41682_n261), .Y(alu__abc_41682_n262) );
  NAND3X1 NAND3X1_194 ( .A(alu__abc_41682_n262), .B(alu__abc_41682_n264), .C(alu__abc_41682_n267), .Y(alu__abc_41682_n268_1) );
  NAND3X1 NAND3X1_195 ( .A(alu__abc_41682_n294), .B(alu__abc_41682_n298), .C(alu__abc_41682_n301), .Y(alu__abc_41682_n302) );
  NAND3X1 NAND3X1_196 ( .A(alu__abc_41682_n105), .B(alu__abc_41682_n307), .C(alu__abc_41682_n299), .Y(alu__abc_41682_n308) );
  NAND3X1 NAND3X1_197 ( .A(alu__abc_41682_n276), .B(alu__abc_41682_n286_1), .C(alu__abc_41682_n314_1), .Y(alu__abc_41682_n315) );
  NAND3X1 NAND3X1_198 ( .A(alu__abc_41682_n288), .B(alu__abc_41682_n316), .C(alu__abc_41682_n315), .Y(alu__abc_41682_n317) );
  NAND3X1 NAND3X1_199 ( .A(alu__abc_41682_n288), .B(alu__abc_41682_n312), .C(alu__abc_41682_n315), .Y(alu__abc_41682_n323) );
  NAND3X1 NAND3X1_2 ( .A(_abc_42016_n660), .B(_abc_42016_n813), .C(_abc_42016_n815), .Y(_abc_42016_n816) );
  NAND3X1 NAND3X1_20 ( .A(_abc_42016_n1201), .B(_abc_42016_n1206), .C(_abc_42016_n1207), .Y(_abc_42016_n1208) );
  NAND3X1 NAND3X1_200 ( .A(alu__abc_41682_n259_1), .B(alu__abc_41682_n322), .C(alu__abc_41682_n325), .Y(alu__abc_41682_n326) );
  NAND3X1 NAND3X1_201 ( .A(alu__abc_41682_n225), .B(alu__abc_41682_n227), .C(alu__abc_41682_n327), .Y(alu__abc_41682_n328) );
  NAND3X1 NAND3X1_202 ( .A(alu__abc_41682_n259_1), .B(alu__abc_41682_n322), .C(alu__abc_41682_n318), .Y(alu__abc_41682_n332) );
  NAND3X1 NAND3X1_203 ( .A(alu__abc_41682_n303), .B(alu__abc_41682_n311), .C(alu__abc_41682_n290), .Y(alu__abc_41682_n336) );
  NAND3X1 NAND3X1_204 ( .A(alu__abc_41682_n360), .B(alu__abc_41682_n365), .C(alu__abc_41682_n364), .Y(alu_cout) );
  NAND3X1 NAND3X1_21 ( .A(_abc_42016_n1213), .B(_abc_42016_n1163), .C(_abc_42016_n1117), .Y(_abc_42016_n1214) );
  NAND3X1 NAND3X1_22 ( .A(_abc_42016_n1162), .B(_abc_42016_n1212), .C(_abc_42016_n1214), .Y(_abc_42016_n1230) );
  NAND3X1 NAND3X1_23 ( .A(_abc_42016_n1229), .B(_abc_42016_n1231), .C(_abc_42016_n1230), .Y(_abc_42016_n1232) );
  NAND3X1 NAND3X1_24 ( .A(_abc_42016_n1193), .B(_abc_42016_n1236), .C(_abc_42016_n1197_1), .Y(_abc_42016_n1239) );
  NAND3X1 NAND3X1_25 ( .A(_abc_42016_n1238), .B(_abc_42016_n1239), .C(_abc_42016_n1036), .Y(_abc_42016_n1240) );
  NAND3X1 NAND3X1_26 ( .A(_abc_42016_n1036), .B(_abc_42016_n1266), .C(_abc_42016_n1268), .Y(_abc_42016_n1269) );
  NAND3X1 NAND3X1_27 ( .A(_abc_42016_n1305), .B(_abc_42016_n1308), .C(_abc_42016_n1266), .Y(_abc_42016_n1310) );
  NAND3X1 NAND3X1_28 ( .A(_abc_42016_n1336), .B(_abc_42016_n1340), .C(_abc_42016_n1059), .Y(_abc_42016_n1341_1) );
  NAND3X1 NAND3X1_29 ( .A(pc_8_), .B(pc_9_), .C(pc_10_), .Y(_abc_42016_n1451) );
  NAND3X1 NAND3X1_3 ( .A(_abc_42016_n823), .B(_abc_42016_n825), .C(_abc_42016_n822), .Y(_abc_42016_n826_1) );
  NAND3X1 NAND3X1_30 ( .A(_abc_42016_n1634), .B(_abc_42016_n1635), .C(_abc_42016_n1630_1), .Y(_abc_42016_n1636) );
  NAND3X1 NAND3X1_31 ( .A(_abc_42016_n1653), .B(_abc_42016_n1654), .C(_abc_42016_n1649_1), .Y(_abc_42016_n1655) );
  NAND3X1 NAND3X1_32 ( .A(_abc_42016_n1670), .B(_abc_42016_n1673_1), .C(_abc_42016_n1669), .Y(_abc_42016_n1674_1) );
  NAND3X1 NAND3X1_33 ( .A(_abc_42016_n647), .B(_abc_42016_n1677), .C(_abc_42016_n660), .Y(_abc_42016_n1678) );
  NAND3X1 NAND3X1_34 ( .A(_abc_42016_n1679), .B(_abc_42016_n1682_1), .C(_abc_42016_n1678), .Y(_abc_42016_n1683) );
  NAND3X1 NAND3X1_35 ( .A(_abc_42016_n648_1), .B(_abc_42016_n1688), .C(_abc_42016_n660), .Y(_abc_42016_n1689_1) );
  NAND3X1 NAND3X1_36 ( .A(_abc_42016_n1717), .B(_abc_42016_n1713_1), .C(_abc_42016_n1716), .Y(_abc_42016_n1718) );
  NAND3X1 NAND3X1_37 ( .A(_abc_42016_n1720), .B(_abc_42016_n1723), .C(_abc_42016_n1719), .Y(_abc_42016_n1724) );
  NAND3X1 NAND3X1_38 ( .A(_abc_42016_n688), .B(_abc_42016_n1740), .C(_abc_42016_n1735), .Y(_abc_42016_n1741) );
  NAND3X1 NAND3X1_39 ( .A(_abc_42016_n1743), .B(_abc_42016_n1745), .C(_abc_42016_n1742), .Y(_abc_42016_n1746) );
  NAND3X1 NAND3X1_4 ( .A(_abc_42016_n831), .B(_abc_42016_n832), .C(_abc_42016_n821), .Y(_abc_36783_n3370) );
  NAND3X1 NAND3X1_40 ( .A(_abc_42016_n919), .B(_abc_42016_n779), .C(_abc_42016_n1734), .Y(_abc_42016_n1789) );
  NAND3X1 NAND3X1_41 ( .A(regfil_2__6_), .B(_abc_42016_n779), .C(_abc_42016_n1733), .Y(_abc_42016_n1790) );
  NAND3X1 NAND3X1_42 ( .A(_abc_42016_n1790), .B(_abc_42016_n1791), .C(_abc_42016_n1789), .Y(_abc_42016_n1792) );
  NAND3X1 NAND3X1_43 ( .A(_abc_42016_n1922_1), .B(_abc_42016_n1931), .C(_abc_42016_n1929), .Y(aluopra_0__FF_INPUT) );
  NAND3X1 NAND3X1_44 ( .A(_abc_42016_n1957_1), .B(_abc_42016_n1959), .C(_abc_42016_n1958), .Y(aluopra_2__FF_INPUT) );
  NAND3X1 NAND3X1_45 ( .A(_abc_42016_n559), .B(_abc_42016_n668), .C(_abc_42016_n1463), .Y(_abc_42016_n2070) );
  NAND3X1 NAND3X1_46 ( .A(_abc_42016_n548), .B(_abc_42016_n2040), .C(_abc_42016_n2035), .Y(_abc_42016_n2081) );
  NAND3X1 NAND3X1_47 ( .A(_abc_42016_n1916), .B(_abc_42016_n2089), .C(_abc_42016_n1508), .Y(_abc_42016_n2090) );
  NAND3X1 NAND3X1_48 ( .A(_abc_42016_n2134), .B(_abc_42016_n1329_1), .C(_abc_42016_n1284), .Y(_abc_42016_n2135_1) );
  NAND3X1 NAND3X1_49 ( .A(_abc_42016_n1326), .B(_abc_42016_n2133), .C(_abc_42016_n2135_1), .Y(_abc_42016_n2136_1) );
  NAND3X1 NAND3X1_5 ( .A(_abc_42016_n862), .B(_abc_42016_n863), .C(_abc_42016_n822), .Y(_abc_42016_n864) );
  NAND3X1 NAND3X1_50 ( .A(_abc_42016_n2129), .B(_abc_42016_n2130), .C(_abc_42016_n2136_1), .Y(_abc_42016_n2137) );
  NAND3X1 NAND3X1_51 ( .A(_abc_42016_n2124_1), .B(_abc_42016_n2126), .C(_abc_42016_n2137), .Y(_abc_42016_n2138) );
  NAND3X1 NAND3X1_52 ( .A(_abc_42016_n2120_1), .B(_abc_42016_n2121), .C(_abc_42016_n2138), .Y(_abc_42016_n2139_1) );
  NAND3X1 NAND3X1_53 ( .A(_abc_42016_n2115_1), .B(_abc_42016_n2117), .C(_abc_42016_n2139_1), .Y(_abc_42016_n2140_1) );
  NAND3X1 NAND3X1_54 ( .A(_abc_42016_n2111), .B(_abc_42016_n2112), .C(_abc_42016_n2140_1), .Y(_abc_42016_n2141) );
  NAND3X1 NAND3X1_55 ( .A(_abc_42016_n2106), .B(_abc_42016_n2108), .C(_abc_42016_n2141), .Y(_abc_42016_n2142) );
  NAND3X1 NAND3X1_56 ( .A(_abc_42016_n1313), .B(_abc_42016_n2168), .C(_abc_42016_n1314), .Y(_abc_42016_n2169) );
  NAND3X1 NAND3X1_57 ( .A(_abc_42016_n2166), .B(_abc_42016_n2167), .C(_abc_42016_n2169), .Y(_abc_42016_n2170) );
  NAND3X1 NAND3X1_58 ( .A(_abc_42016_n2164), .B(_abc_42016_n2165), .C(_abc_42016_n2170), .Y(_abc_42016_n2171) );
  NAND3X1 NAND3X1_59 ( .A(_abc_42016_n2161), .B(_abc_42016_n2162), .C(_abc_42016_n2171), .Y(_abc_42016_n2172_1) );
  NAND3X1 NAND3X1_6 ( .A(_abc_42016_n867_1), .B(_abc_42016_n864), .C(_abc_42016_n868), .Y(_abc_42016_n869) );
  NAND3X1 NAND3X1_60 ( .A(_abc_42016_n2158), .B(_abc_42016_n2159), .C(_abc_42016_n2172_1), .Y(_abc_42016_n2173) );
  NAND3X1 NAND3X1_61 ( .A(_abc_42016_n2154), .B(_abc_42016_n2156), .C(_abc_42016_n2173), .Y(_abc_42016_n2174) );
  NAND3X1 NAND3X1_62 ( .A(_abc_42016_n2152), .B(_abc_42016_n2153), .C(_abc_42016_n2174), .Y(_abc_42016_n2175) );
  NAND3X1 NAND3X1_63 ( .A(_abc_42016_n2149), .B(_abc_42016_n2150), .C(_abc_42016_n2175), .Y(_abc_42016_n2176) );
  NAND3X1 NAND3X1_64 ( .A(_abc_42016_n1305), .B(_abc_42016_n2201), .C(_abc_42016_n1266), .Y(_abc_42016_n2202) );
  NAND3X1 NAND3X1_65 ( .A(_abc_42016_n2198), .B(_abc_42016_n2200), .C(_abc_42016_n2202), .Y(_abc_42016_n2203) );
  NAND3X1 NAND3X1_66 ( .A(_abc_42016_n2196), .B(_abc_42016_n2197), .C(_abc_42016_n2203), .Y(_abc_42016_n2204) );
  NAND3X1 NAND3X1_67 ( .A(_abc_42016_n2193), .B(_abc_42016_n2194), .C(_abc_42016_n2204), .Y(_abc_42016_n2205) );
  NAND3X1 NAND3X1_68 ( .A(_abc_42016_n2190), .B(_abc_42016_n2191), .C(_abc_42016_n2205), .Y(_abc_42016_n2206) );
  NAND3X1 NAND3X1_69 ( .A(_abc_42016_n2187), .B(_abc_42016_n2188), .C(_abc_42016_n2206), .Y(_abc_42016_n2207) );
  NAND3X1 NAND3X1_7 ( .A(_abc_42016_n660), .B(_abc_42016_n955), .C(_abc_42016_n953), .Y(_abc_42016_n956) );
  NAND3X1 NAND3X1_70 ( .A(_abc_42016_n2185), .B(_abc_42016_n2186), .C(_abc_42016_n2207), .Y(_abc_42016_n2208) );
  NAND3X1 NAND3X1_71 ( .A(_abc_42016_n2182), .B(_abc_42016_n2183), .C(_abc_42016_n2208), .Y(_abc_42016_n2209) );
  NAND3X1 NAND3X1_72 ( .A(_abc_42016_n529), .B(eienb), .C(_abc_42016_n2024), .Y(_abc_42016_n2257) );
  NAND3X1 NAND3X1_73 ( .A(_abc_42016_n2284), .B(_abc_42016_n2313), .C(_abc_42016_n2312), .Y(_abc_42016_n2314) );
  NAND3X1 NAND3X1_74 ( .A(_abc_42016_n2350), .B(_abc_42016_n2360), .C(_abc_42016_n2354), .Y(_abc_42016_n2361) );
  NAND3X1 NAND3X1_75 ( .A(_abc_42016_n2538), .B(_abc_42016_n2546), .C(_abc_42016_n2541), .Y(_abc_42016_n2547_1) );
  NAND3X1 NAND3X1_76 ( .A(_abc_42016_n2605), .B(_abc_42016_n2608_1), .C(_abc_42016_n2604), .Y(_abc_42016_n2609_1) );
  NAND3X1 NAND3X1_77 ( .A(_abc_42016_n2626), .B(_abc_42016_n2628), .C(_abc_42016_n2627), .Y(_abc_42016_n2629) );
  NAND3X1 NAND3X1_78 ( .A(_abc_42016_n2637), .B(_abc_42016_n2642), .C(_abc_42016_n2638), .Y(_abc_42016_n2643) );
  NAND3X1 NAND3X1_79 ( .A(_abc_42016_n2691), .B(_abc_42016_n2693), .C(_abc_42016_n2690), .Y(_abc_42016_n2694) );
  NAND3X1 NAND3X1_8 ( .A(_abc_42016_n957_1), .B(_abc_42016_n969), .C(_abc_42016_n956), .Y(_abc_42016_n970) );
  NAND3X1 NAND3X1_80 ( .A(_abc_42016_n2272), .B(_abc_42016_n548), .C(_abc_42016_n2733), .Y(_abc_42016_n2734) );
  NAND3X1 NAND3X1_81 ( .A(_abc_42016_n1879_1), .B(_abc_42016_n2958), .C(_abc_42016_n2957), .Y(_abc_42016_n2959) );
  NAND3X1 NAND3X1_82 ( .A(_abc_42016_n3009), .B(_abc_42016_n2732), .C(_abc_42016_n3003), .Y(_abc_42016_n3010) );
  NAND3X1 NAND3X1_83 ( .A(_abc_42016_n3021), .B(_abc_42016_n3020), .C(_abc_42016_n3017), .Y(_abc_42016_n3022) );
  NAND3X1 NAND3X1_84 ( .A(sp_0_), .B(_abc_42016_n673), .C(_abc_42016_n1411), .Y(_abc_42016_n3038) );
  NAND3X1 NAND3X1_85 ( .A(_abc_42016_n3037), .B(_abc_42016_n3041), .C(_abc_42016_n3038), .Y(_abc_42016_n3042) );
  NAND3X1 NAND3X1_86 ( .A(_abc_42016_n3088), .B(_abc_42016_n3089), .C(_abc_42016_n3091), .Y(_abc_42016_n3092) );
  NAND3X1 NAND3X1_87 ( .A(_abc_42016_n1863), .B(_abc_42016_n3212), .C(_abc_42016_n3211), .Y(_abc_42016_n3213) );
  NAND3X1 NAND3X1_88 ( .A(_abc_42016_n1863), .B(_abc_42016_n3234), .C(_abc_42016_n3233), .Y(_abc_42016_n3235) );
  NAND3X1 NAND3X1_89 ( .A(_abc_42016_n1863), .B(_abc_42016_n3280), .C(_abc_42016_n3279), .Y(_abc_42016_n3281) );
  NAND3X1 NAND3X1_9 ( .A(_abc_42016_n978), .B(_abc_42016_n983), .C(_abc_42016_n982), .Y(_abc_42016_n984) );
  NAND3X1 NAND3X1_90 ( .A(_abc_42016_n1863), .B(_abc_42016_n3330), .C(_abc_42016_n3324), .Y(_abc_42016_n3331) );
  NAND3X1 NAND3X1_91 ( .A(_abc_42016_n529), .B(rdatahold2_0_), .C(_abc_42016_n3459), .Y(_abc_42016_n3465) );
  NAND3X1 NAND3X1_92 ( .A(_abc_42016_n3465), .B(_abc_42016_n3467), .C(_abc_42016_n3464), .Y(sp_0__FF_INPUT) );
  NAND3X1 NAND3X1_93 ( .A(_abc_42016_n3473), .B(_abc_42016_n3481), .C(_abc_42016_n3480), .Y(_abc_42016_n3482_1) );
  NAND3X1 NAND3X1_94 ( .A(_abc_42016_n3518_1), .B(_abc_42016_n3520), .C(_abc_42016_n3474), .Y(_abc_42016_n3521) );
  NAND3X1 NAND3X1_95 ( .A(sp_4_), .B(_abc_42016_n3519), .C(_abc_42016_n2255), .Y(_abc_42016_n3545) );
  NAND3X1 NAND3X1_96 ( .A(_abc_42016_n3561), .B(_abc_42016_n3573), .C(_abc_42016_n3570), .Y(_abc_42016_n3574) );
  NAND3X1 NAND3X1_97 ( .A(_abc_42016_n3685), .B(_abc_42016_n3677), .C(_abc_42016_n3684), .Y(_abc_42016_n3686) );
  NAND3X1 NAND3X1_98 ( .A(sp_11_), .B(sp_10_), .C(sp_9_), .Y(_abc_42016_n3692) );
  NAND3X1 NAND3X1_99 ( .A(_abc_42016_n2347_1), .B(_abc_42016_n3694), .C(_abc_42016_n3695), .Y(_abc_42016_n3696) );
  NOR2X1 NOR2X1_1 ( .A(state_3_), .B(_abc_42016_n501), .Y(_abc_42016_n502) );
  NOR2X1 NOR2X1_10 ( .A(_abc_42016_n520), .B(_abc_42016_n523_1), .Y(_abc_42016_n524_1) );
  NOR2X1 NOR2X1_100 ( .A(_abc_42016_n664_1), .B(_abc_42016_n990), .Y(_abc_42016_n991) );
  NOR2X1 NOR2X1_101 ( .A(_abc_42016_n992), .B(_abc_42016_n585), .Y(_abc_42016_n993) );
  NOR2X1 NOR2X1_102 ( .A(_abc_42016_n669), .B(_abc_42016_n682), .Y(_abc_42016_n996) );
  NOR2X1 NOR2X1_103 ( .A(_abc_42016_n568), .B(_abc_42016_n626), .Y(_abc_42016_n998) );
  NOR2X1 NOR2X1_104 ( .A(_abc_42016_n680), .B(_abc_42016_n999), .Y(_abc_42016_n1000) );
  NOR2X1 NOR2X1_105 ( .A(_abc_42016_n604_1), .B(_abc_42016_n999), .Y(_abc_42016_n1001_1) );
  NOR2X1 NOR2X1_106 ( .A(_abc_42016_n531), .B(_abc_42016_n530), .Y(_abc_42016_n1003) );
  NOR2X1 NOR2X1_107 ( .A(_abc_42016_n1004), .B(_abc_42016_n999), .Y(_abc_42016_n1005) );
  NOR2X1 NOR2X1_108 ( .A(_abc_42016_n669), .B(_abc_42016_n999), .Y(_abc_42016_n1006) );
  NOR2X1 NOR2X1_109 ( .A(_abc_42016_n1010), .B(_abc_42016_n995), .Y(_abc_42016_n1011) );
  NOR2X1 NOR2X1_11 ( .A(_abc_42016_n518_1), .B(_abc_42016_n525), .Y(_abc_42016_n526_1) );
  NOR2X1 NOR2X1_110 ( .A(_abc_42016_n511), .B(_abc_42016_n523_1), .Y(_abc_42016_n1013) );
  NOR2X1 NOR2X1_111 ( .A(state_0_), .B(_abc_42016_n504), .Y(_abc_42016_n1015) );
  NOR2X1 NOR2X1_112 ( .A(_abc_42016_n576_1), .B(_abc_42016_n1016), .Y(_abc_42016_n1017) );
  NOR2X1 NOR2X1_113 ( .A(_abc_42016_n1019), .B(_abc_42016_n1012), .Y(_abc_42016_n1020) );
  NOR2X1 NOR2X1_114 ( .A(_abc_42016_n1022), .B(_abc_42016_n562), .Y(_abc_42016_n1023) );
  NOR2X1 NOR2X1_115 ( .A(regfil_5__0_), .B(sp_0_), .Y(_abc_42016_n1026) );
  NOR2X1 NOR2X1_116 ( .A(_abc_42016_n1035), .B(_abc_42016_n562), .Y(_abc_42016_n1036) );
  NOR2X1 NOR2X1_117 ( .A(_abc_42016_n1046), .B(_abc_42016_n562), .Y(_abc_42016_n1047_1) );
  NOR2X1 NOR2X1_118 ( .A(_abc_42016_n995), .B(_abc_42016_n1050), .Y(_abc_42016_n1051) );
  NOR2X1 NOR2X1_119 ( .A(_abc_42016_n695), .B(_abc_42016_n1046), .Y(_abc_42016_n1060) );
  NOR2X1 NOR2X1_12 ( .A(opcode_3_), .B(_abc_42016_n531), .Y(_abc_42016_n532_1) );
  NOR2X1 NOR2X1_120 ( .A(regfil_5__0_), .B(regfil_5__1_), .Y(_abc_42016_n1062) );
  NOR2X1 NOR2X1_121 ( .A(_abc_42016_n695), .B(_abc_42016_n709), .Y(_abc_42016_n1063) );
  NOR2X1 NOR2X1_122 ( .A(_abc_42016_n1062), .B(_abc_42016_n1063), .Y(_abc_42016_n1064) );
  NOR2X1 NOR2X1_123 ( .A(_abc_42016_n1060), .B(_abc_42016_n1066), .Y(_abc_42016_n1067) );
  NOR2X1 NOR2X1_124 ( .A(regfil_5__1_), .B(sp_1_), .Y(_abc_42016_n1068) );
  NOR2X1 NOR2X1_125 ( .A(_abc_42016_n1068), .B(_abc_42016_n1070_1), .Y(_abc_42016_n1072) );
  NOR2X1 NOR2X1_126 ( .A(regfil_1__1_), .B(regfil_5__1_), .Y(_abc_42016_n1074) );
  NOR2X1 NOR2X1_127 ( .A(_abc_42016_n645), .B(_abc_42016_n709), .Y(_abc_42016_n1075) );
  NOR2X1 NOR2X1_128 ( .A(_abc_42016_n1074), .B(_abc_42016_n1075), .Y(_abc_42016_n1076) );
  NOR2X1 NOR2X1_129 ( .A(_abc_42016_n703), .B(_abc_42016_n709), .Y(_abc_42016_n1079) );
  NOR2X1 NOR2X1_13 ( .A(opcode_0_), .B(_abc_42016_n537_1), .Y(_abc_42016_n538_1) );
  NOR2X1 NOR2X1_130 ( .A(regfil_3__1_), .B(regfil_5__1_), .Y(_abc_42016_n1080) );
  NOR2X1 NOR2X1_131 ( .A(_abc_42016_n1080), .B(_abc_42016_n1079), .Y(_abc_42016_n1081) );
  NOR2X1 NOR2X1_132 ( .A(reset), .B(_abc_42016_n1014), .Y(_abc_42016_n1096) );
  NOR2X1 NOR2X1_133 ( .A(_abc_42016_n1096), .B(_abc_42016_n993), .Y(_abc_42016_n1097) );
  NOR2X1 NOR2X1_134 ( .A(_abc_42016_n773), .B(_abc_42016_n757), .Y(_abc_42016_n1101_1) );
  NOR2X1 NOR2X1_135 ( .A(regfil_3__2_), .B(regfil_5__2_), .Y(_abc_42016_n1102) );
  NOR2X1 NOR2X1_136 ( .A(_abc_42016_n1102), .B(_abc_42016_n1101_1), .Y(_abc_42016_n1103_1) );
  NOR2X1 NOR2X1_137 ( .A(_abc_42016_n671_1), .B(_abc_42016_n562), .Y(_abc_42016_n1125) );
  NOR2X1 NOR2X1_138 ( .A(_abc_42016_n1061), .B(_abc_42016_n562), .Y(_abc_42016_n1138) );
  NOR2X1 NOR2X1_139 ( .A(regfil_5__3_), .B(sp_3_), .Y(_abc_42016_n1161) );
  NOR2X1 NOR2X1_14 ( .A(opcode_7_), .B(_abc_42016_n540), .Y(_abc_42016_n541) );
  NOR2X1 NOR2X1_140 ( .A(regfil_5__3_), .B(_abc_42016_n1126), .Y(_abc_42016_n1183) );
  NOR2X1 NOR2X1_141 ( .A(_abc_42016_n1185), .B(_abc_42016_n1170), .Y(_abc_42016_n1186) );
  NOR2X1 NOR2X1_142 ( .A(regfil_5__4_), .B(sp_4_), .Y(_abc_42016_n1209) );
  NOR2X1 NOR2X1_143 ( .A(_abc_42016_n843), .B(_abc_42016_n1210), .Y(_abc_42016_n1211) );
  NOR2X1 NOR2X1_144 ( .A(_abc_42016_n1209), .B(_abc_42016_n1211), .Y(_abc_42016_n1212) );
  NOR2X1 NOR2X1_145 ( .A(_abc_42016_n874), .B(_abc_42016_n697), .Y(_abc_42016_n1223) );
  NOR2X1 NOR2X1_146 ( .A(_abc_42016_n872), .B(_abc_42016_n1188), .Y(_abc_42016_n1226) );
  NOR2X1 NOR2X1_147 ( .A(_abc_42016_n843), .B(_abc_42016_n669), .Y(_abc_42016_n1245) );
  NOR2X1 NOR2X1_148 ( .A(regfil_5__5_), .B(_abc_42016_n1184), .Y(_abc_42016_n1251) );
  NOR2X1 NOR2X1_149 ( .A(_abc_42016_n642), .B(_abc_42016_n872), .Y(_abc_42016_n1264) );
  NOR2X1 NOR2X1_15 ( .A(state_1_), .B(state_0_), .Y(_abc_42016_n543) );
  NOR2X1 NOR2X1_150 ( .A(_abc_42016_n874), .B(_abc_42016_n872), .Y(_abc_42016_n1270) );
  NOR2X1 NOR2X1_151 ( .A(_abc_42016_n872), .B(_abc_42016_n1046), .Y(_abc_42016_n1276) );
  NOR2X1 NOR2X1_152 ( .A(_abc_42016_n1281), .B(_abc_42016_n1280), .Y(_abc_42016_n1282) );
  NOR2X1 NOR2X1_153 ( .A(_abc_42016_n872), .B(_abc_42016_n1279), .Y(_abc_42016_n1283) );
  NOR2X1 NOR2X1_154 ( .A(regfil_5__6_), .B(_abc_42016_n1226), .Y(_abc_42016_n1289) );
  NOR2X1 NOR2X1_155 ( .A(_abc_42016_n1296_1), .B(_abc_42016_n1170), .Y(_abc_42016_n1297_1) );
  NOR2X1 NOR2X1_156 ( .A(regfil_1__7_), .B(regfil_5__7_), .Y(_abc_42016_n1306) );
  NOR2X1 NOR2X1_157 ( .A(_abc_42016_n641), .B(_abc_42016_n959), .Y(_abc_42016_n1307) );
  NOR2X1 NOR2X1_158 ( .A(_abc_42016_n1306), .B(_abc_42016_n1307), .Y(_abc_42016_n1308) );
  NOR2X1 NOR2X1_159 ( .A(_abc_42016_n974), .B(_abc_42016_n959), .Y(_abc_42016_n1316) );
  NOR2X1 NOR2X1_16 ( .A(_abc_42016_n544_1), .B(_abc_42016_n503), .Y(_abc_42016_n545_1) );
  NOR2X1 NOR2X1_160 ( .A(regfil_3__7_), .B(regfil_5__7_), .Y(_abc_42016_n1317) );
  NOR2X1 NOR2X1_161 ( .A(_abc_42016_n1317), .B(_abc_42016_n1316), .Y(_abc_42016_n1318) );
  NOR2X1 NOR2X1_162 ( .A(regfil_5__7_), .B(sp_7_), .Y(_abc_42016_n1325) );
  NOR2X1 NOR2X1_163 ( .A(_abc_42016_n959), .B(_abc_42016_n1327_1), .Y(_abc_42016_n1328) );
  NOR2X1 NOR2X1_164 ( .A(_abc_42016_n959), .B(_abc_42016_n1296_1), .Y(_abc_42016_n1334) );
  NOR2X1 NOR2X1_165 ( .A(regfil_5__7_), .B(_abc_42016_n1295), .Y(_abc_42016_n1335_1) );
  NOR2X1 NOR2X1_166 ( .A(_abc_42016_n959), .B(_abc_42016_n1290), .Y(_abc_42016_n1337_1) );
  NOR2X1 NOR2X1_167 ( .A(_abc_42016_n559), .B(_abc_42016_n673), .Y(_abc_42016_n1344) );
  NOR2X1 NOR2X1_168 ( .A(_abc_42016_n1344), .B(_abc_42016_n558), .Y(_abc_42016_n1345) );
  NOR2X1 NOR2X1_169 ( .A(_abc_42016_n572), .B(_abc_42016_n539), .Y(_abc_42016_n1346) );
  NOR2X1 NOR2X1_17 ( .A(_abc_42016_n511), .B(_abc_42016_n546), .Y(_abc_42016_n547) );
  NOR2X1 NOR2X1_170 ( .A(_abc_42016_n669), .B(_abc_42016_n1347), .Y(_abc_42016_n1348) );
  NOR2X1 NOR2X1_171 ( .A(_abc_42016_n1350), .B(_abc_42016_n562), .Y(_abc_42016_n1351) );
  NOR2X1 NOR2X1_172 ( .A(_abc_42016_n1357), .B(_abc_42016_n1358), .Y(_abc_42016_n1359) );
  NOR2X1 NOR2X1_173 ( .A(_abc_42016_n1356), .B(_abc_42016_n1360), .Y(_abc_42016_n1361) );
  NOR2X1 NOR2X1_174 ( .A(_abc_42016_n1355), .B(_abc_42016_n1362), .Y(_abc_42016_n1363) );
  NOR2X1 NOR2X1_175 ( .A(_abc_42016_n1353), .B(_abc_42016_n1366), .Y(_abc_42016_n1367) );
  NOR2X1 NOR2X1_176 ( .A(_abc_42016_n536), .B(_abc_42016_n626), .Y(_abc_42016_n1371) );
  NOR2X1 NOR2X1_177 ( .A(_abc_42016_n604_1), .B(_abc_42016_n1372), .Y(_abc_42016_n1373) );
  NOR2X1 NOR2X1_178 ( .A(_abc_42016_n536), .B(_abc_42016_n727), .Y(_abc_42016_n1376) );
  NOR2X1 NOR2X1_179 ( .A(_abc_42016_n1382), .B(_abc_42016_n1383), .Y(_abc_42016_n1384) );
  NOR2X1 NOR2X1_18 ( .A(_abc_42016_n542), .B(_abc_42016_n548), .Y(_abc_42016_n549) );
  NOR2X1 NOR2X1_180 ( .A(_abc_42016_n1356), .B(_abc_42016_n1385), .Y(_abc_42016_n1386_1) );
  NOR2X1 NOR2X1_181 ( .A(_abc_42016_n1355), .B(_abc_42016_n1387), .Y(_abc_42016_n1388) );
  NOR2X1 NOR2X1_182 ( .A(_abc_42016_n1353), .B(_abc_42016_n1389), .Y(_abc_42016_n1391) );
  NOR2X1 NOR2X1_183 ( .A(opcode_4_), .B(_abc_42016_n608), .Y(_abc_42016_n1394) );
  NOR2X1 NOR2X1_184 ( .A(opcode_3_), .B(_abc_42016_n536), .Y(_abc_42016_n1397) );
  NOR2X1 NOR2X1_185 ( .A(_abc_42016_n1398), .B(_abc_42016_n626), .Y(_abc_42016_n1399) );
  NOR2X1 NOR2X1_186 ( .A(opcode_5_), .B(_abc_42016_n1400), .Y(_abc_42016_n1401) );
  NOR2X1 NOR2X1_187 ( .A(_abc_42016_n1004), .B(_abc_42016_n1400), .Y(_abc_42016_n1402) );
  NOR2X1 NOR2X1_188 ( .A(_abc_42016_n1375), .B(_abc_42016_n1374), .Y(_abc_42016_n1404) );
  NOR2X1 NOR2X1_189 ( .A(_abc_42016_n1409), .B(_abc_42016_n1377), .Y(_abc_42016_n1410_1) );
  NOR2X1 NOR2X1_19 ( .A(_abc_42016_n513), .B(_abc_42016_n509), .Y(_abc_42016_n552) );
  NOR2X1 NOR2X1_190 ( .A(_abc_42016_n1406), .B(_abc_42016_n1413), .Y(_abc_42016_n1414) );
  NOR2X1 NOR2X1_191 ( .A(_abc_42016_n1410_1), .B(_abc_42016_n1459), .Y(_abc_42016_n1460) );
  NOR2X1 NOR2X1_192 ( .A(_abc_42016_n536), .B(_abc_42016_n1461), .Y(_abc_42016_n1462) );
  NOR2X1 NOR2X1_193 ( .A(_abc_42016_n1398), .B(_abc_42016_n565), .Y(_abc_42016_n1463) );
  NOR2X1 NOR2X1_194 ( .A(_abc_42016_n1449), .B(_abc_42016_n1424), .Y(_abc_42016_n1466) );
  NOR2X1 NOR2X1_195 ( .A(_abc_42016_n1451), .B(_abc_42016_n1366), .Y(_abc_42016_n1483) );
  NOR2X1 NOR2X1_196 ( .A(_abc_42016_n1492), .B(_abc_42016_n1410_1), .Y(_abc_42016_n1493) );
  NOR2X1 NOR2X1_197 ( .A(_abc_42016_n1449), .B(_abc_42016_n1435), .Y(_abc_42016_n1505) );
  NOR2X1 NOR2X1_198 ( .A(_abc_42016_n1503), .B(_abc_42016_n1480), .Y(_abc_42016_n1510) );
  NOR2X1 NOR2X1_199 ( .A(opcode_5_), .B(_abc_42016_n1515), .Y(_abc_42016_n1516) );
  NOR2X1 NOR2X1_2 ( .A(_abc_42016_n504), .B(_abc_42016_n505), .Y(_abc_42016_n506) );
  NOR2X1 NOR2X1_20 ( .A(_abc_42016_n554), .B(_abc_42016_n550), .Y(_abc_42016_n555) );
  NOR2X1 NOR2X1_200 ( .A(opcode_5_), .B(_abc_42016_n1535), .Y(_abc_42016_n1536) );
  NOR2X1 NOR2X1_201 ( .A(_abc_42016_n1503), .B(_abc_42016_n1484), .Y(_abc_42016_n1543) );
  NOR2X1 NOR2X1_202 ( .A(_abc_42016_n1381), .B(_abc_42016_n1532), .Y(_abc_42016_n1560) );
  NOR2X1 NOR2X1_203 ( .A(_abc_42016_n1559), .B(_abc_42016_n1562), .Y(_abc_42016_n1563) );
  NOR2X1 NOR2X1_204 ( .A(_abc_42016_n1503), .B(_abc_42016_n1506), .Y(_abc_42016_n1565) );
  NOR2X1 NOR2X1_205 ( .A(_abc_42016_n1557), .B(_abc_42016_n1566), .Y(_abc_42016_n1570) );
  NOR2X1 NOR2X1_206 ( .A(opcode_5_), .B(_abc_42016_n1573), .Y(_abc_42016_n1574) );
  NOR2X1 NOR2X1_207 ( .A(_abc_42016_n1557), .B(_abc_42016_n1532), .Y(_abc_42016_n1585) );
  NOR2X1 NOR2X1_208 ( .A(_abc_42016_n1410_1), .B(_abc_42016_n1597), .Y(_abc_42016_n1598) );
  NOR2X1 NOR2X1_209 ( .A(_abc_42016_n556), .B(_abc_42016_n1605_1), .Y(_abc_42016_n1623) );
  NOR2X1 NOR2X1_21 ( .A(_abc_42016_n513), .B(_abc_42016_n546), .Y(_abc_42016_n557) );
  NOR2X1 NOR2X1_210 ( .A(_abc_42016_n1628), .B(_abc_42016_n772), .Y(_abc_42016_n1629_1) );
  NOR2X1 NOR2X1_211 ( .A(_abc_42016_n1631), .B(_abc_42016_n977), .Y(_abc_42016_n1632) );
  NOR2X1 NOR2X1_212 ( .A(regfil_2__0_), .B(_abc_42016_n976), .Y(_abc_42016_n1633) );
  NOR2X1 NOR2X1_213 ( .A(_abc_42016_n1044), .B(_abc_42016_n587), .Y(_abc_42016_n1637) );
  NOR2X1 NOR2X1_214 ( .A(_abc_42016_n513), .B(_abc_42016_n667), .Y(_abc_42016_n1639_1) );
  NOR2X1 NOR2X1_215 ( .A(_abc_42016_n728), .B(_abc_42016_n1627), .Y(_abc_42016_n1647_1) );
  NOR2X1 NOR2X1_216 ( .A(_abc_42016_n1647_1), .B(_abc_42016_n772), .Y(_abc_42016_n1648) );
  NOR2X1 NOR2X1_217 ( .A(_abc_42016_n728), .B(_abc_42016_n1633), .Y(_abc_42016_n1650) );
  NOR2X1 NOR2X1_218 ( .A(_abc_42016_n612), .B(_abc_42016_n646), .Y(_abc_42016_n1656) );
  NOR2X1 NOR2X1_219 ( .A(_abc_42016_n772), .B(_abc_42016_n1667), .Y(_abc_42016_n1668) );
  NOR2X1 NOR2X1_22 ( .A(opcode_7_), .B(opcode_6_), .Y(_abc_42016_n559) );
  NOR2X1 NOR2X1_220 ( .A(_abc_42016_n753), .B(_abc_42016_n1652_1), .Y(_abc_42016_n1671) );
  NOR2X1 NOR2X1_221 ( .A(regfil_2__2_), .B(_abc_42016_n1651), .Y(_abc_42016_n1672) );
  NOR2X1 NOR2X1_222 ( .A(regfil_2__3_), .B(_abc_42016_n1667), .Y(_abc_42016_n1697_1) );
  NOR2X1 NOR2X1_223 ( .A(_abc_42016_n796), .B(_abc_42016_n1666), .Y(_abc_42016_n1711) );
  NOR2X1 NOR2X1_224 ( .A(regfil_2__4_), .B(_abc_42016_n1700), .Y(_abc_42016_n1715) );
  NOR2X1 NOR2X1_225 ( .A(_abc_42016_n895), .B(_abc_42016_n1715), .Y(_abc_42016_n1732_1) );
  NOR2X1 NOR2X1_226 ( .A(_abc_42016_n895), .B(_abc_42016_n1736), .Y(_abc_42016_n1737) );
  NOR2X1 NOR2X1_227 ( .A(regfil_1__6_), .B(_abc_42016_n1623), .Y(_abc_42016_n1749_1) );
  NOR2X1 NOR2X1_228 ( .A(_abc_42016_n609), .B(_abc_42016_n616), .Y(_abc_42016_n1752) );
  NOR2X1 NOR2X1_229 ( .A(_abc_42016_n641), .B(_abc_42016_n1751), .Y(_abc_42016_n1760) );
  NOR2X1 NOR2X1_23 ( .A(_abc_42016_n560), .B(_abc_42016_n558), .Y(_abc_42016_n561) );
  NOR2X1 NOR2X1_230 ( .A(_abc_42016_n1762), .B(_abc_42016_n1759), .Y(_abc_42016_n1763) );
  NOR2X1 NOR2X1_231 ( .A(regfil_1__7_), .B(_abc_42016_n1623), .Y(_abc_42016_n1764) );
  NOR2X1 NOR2X1_232 ( .A(_abc_42016_n1604_1), .B(_abc_42016_n599), .Y(_abc_42016_n1767_1) );
  NOR2X1 NOR2X1_233 ( .A(_abc_42016_n684), .B(_abc_42016_n1807), .Y(_abc_42016_n1808) );
  NOR2X1 NOR2X1_234 ( .A(_abc_42016_n596), .B(_abc_42016_n593), .Y(_abc_42016_n1813) );
  NOR2X1 NOR2X1_235 ( .A(_abc_42016_n1604_1), .B(_abc_42016_n1814), .Y(_abc_42016_n1815) );
  NOR2X1 NOR2X1_236 ( .A(regfil_6__0_), .B(_abc_42016_n1815), .Y(_abc_42016_n1816) );
  NOR2X1 NOR2X1_237 ( .A(regfil_6__4_), .B(_abc_42016_n1815), .Y(_abc_42016_n1824) );
  NOR2X1 NOR2X1_238 ( .A(_abc_42016_n539), .B(_abc_42016_n1398), .Y(_abc_42016_n1835) );
  NOR2X1 NOR2X1_239 ( .A(_abc_42016_n536), .B(_abc_42016_n539), .Y(_abc_42016_n1841) );
  NOR2X1 NOR2X1_24 ( .A(_abc_42016_n563), .B(_abc_42016_n537_1), .Y(_abc_42016_n564) );
  NOR2X1 NOR2X1_240 ( .A(_abc_42016_n1842), .B(_abc_42016_n558), .Y(_abc_42016_n1843) );
  NOR2X1 NOR2X1_241 ( .A(opcode_4_), .B(_abc_42016_n1848), .Y(_abc_42016_n1849) );
  NOR2X1 NOR2X1_242 ( .A(opcode_6_), .B(_abc_42016_n672_1), .Y(_abc_42016_n1851) );
  NOR2X1 NOR2X1_243 ( .A(state_4_), .B(_abc_42016_n1867), .Y(_abc_42016_n1868) );
  NOR2X1 NOR2X1_244 ( .A(state_2_), .B(state_3_), .Y(_abc_42016_n1869) );
  NOR2X1 NOR2X1_245 ( .A(_abc_42016_n1870), .B(_abc_42016_n520), .Y(_abc_42016_n1871) );
  NOR2X1 NOR2X1_246 ( .A(_abc_42016_n503), .B(_abc_42016_n1016), .Y(_abc_42016_n1872) );
  NOR2X1 NOR2X1_247 ( .A(reset), .B(_abc_42016_n1873_1), .Y(_abc_42016_n1874_1) );
  NOR2X1 NOR2X1_248 ( .A(_abc_42016_n557), .B(_abc_42016_n1874_1), .Y(_abc_42016_n1875_1) );
  NOR2X1 NOR2X1_249 ( .A(_abc_42016_n1863), .B(_abc_42016_n558), .Y(_abc_42016_n1882) );
  NOR2X1 NOR2X1_25 ( .A(opcode_2_), .B(_abc_42016_n566), .Y(_abc_42016_n567) );
  NOR2X1 NOR2X1_250 ( .A(opcode_4_), .B(opcode_3_), .Y(_abc_42016_n1911) );
  NOR2X1 NOR2X1_251 ( .A(opcode_4_), .B(_abc_42016_n566), .Y(_abc_42016_n1915) );
  NOR2X1 NOR2X1_252 ( .A(_abc_42016_n531), .B(_abc_42016_n566), .Y(_abc_42016_n1917) );
  NOR2X1 NOR2X1_253 ( .A(_abc_42016_n1923), .B(_abc_42016_n581_1), .Y(_abc_42016_n1924) );
  NOR2X1 NOR2X1_254 ( .A(_abc_42016_n1950_1), .B(_abc_42016_n1948), .Y(_abc_42016_n1951) );
  NOR2X1 NOR2X1_255 ( .A(_abc_42016_n2012), .B(_abc_42016_n2011), .Y(_abc_42016_n2013) );
  NOR2X1 NOR2X1_256 ( .A(_abc_42016_n2025), .B(_abc_42016_n2027), .Y(intcyc_FF_INPUT) );
  NOR2X1 NOR2X1_257 ( .A(state_5_), .B(_abc_42016_n514), .Y(_abc_42016_n2030) );
  NOR2X1 NOR2X1_258 ( .A(_abc_42016_n2031), .B(_abc_42016_n581_1), .Y(_abc_42016_n2032) );
  NOR2X1 NOR2X1_259 ( .A(_abc_42016_n511), .B(_abc_42016_n2033), .Y(_abc_42016_n2034) );
  NOR2X1 NOR2X1_26 ( .A(_abc_42016_n568), .B(_abc_42016_n565), .Y(_abc_42016_n569) );
  NOR2X1 NOR2X1_260 ( .A(_abc_42016_n686), .B(_abc_42016_n992), .Y(_abc_42016_n2041) );
  NOR2X1 NOR2X1_261 ( .A(_abc_42016_n2042), .B(_abc_42016_n2040), .Y(_abc_42016_n2043) );
  NOR2X1 NOR2X1_262 ( .A(_abc_42016_n1130), .B(_abc_42016_n2044), .Y(_abc_42016_n2045) );
  NOR2X1 NOR2X1_263 ( .A(_abc_42016_n2041), .B(_abc_42016_n2040), .Y(_abc_42016_n2047) );
  NOR2X1 NOR2X1_264 ( .A(_abc_42016_n2047), .B(_abc_42016_n2037), .Y(_abc_42016_n2048) );
  NOR2X1 NOR2X1_265 ( .A(_abc_42016_n1302), .B(_abc_42016_n2044), .Y(_abc_42016_n2057) );
  NOR2X1 NOR2X1_266 ( .A(state_4_), .B(_abc_42016_n509), .Y(_abc_42016_n2059) );
  NOR2X1 NOR2X1_267 ( .A(_abc_42016_n1974), .B(_abc_42016_n2066), .Y(_abc_42016_n2067) );
  NOR2X1 NOR2X1_268 ( .A(_abc_42016_n924), .B(_abc_42016_n2068), .Y(_abc_42016_n2069) );
  NOR2X1 NOR2X1_269 ( .A(_abc_42016_n1870), .B(_abc_42016_n1016), .Y(_abc_42016_n2078) );
  NOR2X1 NOR2X1_27 ( .A(opcode_4_), .B(opcode_5_), .Y(_abc_42016_n570) );
  NOR2X1 NOR2X1_270 ( .A(_abc_42016_n1923), .B(_abc_42016_n2079), .Y(_abc_42016_n2080) );
  NOR2X1 NOR2X1_271 ( .A(regfil_4__7_), .B(sp_15_), .Y(_abc_42016_n2083) );
  NOR2X1 NOR2X1_272 ( .A(opcode_5_), .B(_abc_42016_n2085), .Y(_abc_42016_n2086) );
  NOR2X1 NOR2X1_273 ( .A(_abc_42016_n668), .B(_abc_42016_n679), .Y(_abc_42016_n2089) );
  NOR2X1 NOR2X1_274 ( .A(opcode_5_), .B(_abc_42016_n2084), .Y(_abc_42016_n2093) );
  NOR2X1 NOR2X1_275 ( .A(_abc_42016_n960), .B(_abc_42016_n2094), .Y(_abc_42016_n2095) );
  NOR2X1 NOR2X1_276 ( .A(_abc_42016_n2095), .B(_abc_42016_n2097), .Y(_abc_42016_n2098) );
  NOR2X1 NOR2X1_277 ( .A(_abc_42016_n2092), .B(_abc_42016_n2099), .Y(_abc_42016_n2100) );
  NOR2X1 NOR2X1_278 ( .A(_abc_42016_n1801_1), .B(_abc_42016_n2101), .Y(_abc_42016_n2102_1) );
  NOR2X1 NOR2X1_279 ( .A(regfil_4__5_), .B(sp_13_), .Y(_abc_42016_n2107) );
  NOR2X1 NOR2X1_28 ( .A(opcode_3_), .B(opcode_2_), .Y(_abc_42016_n571) );
  NOR2X1 NOR2X1_280 ( .A(_abc_42016_n1527), .B(_abc_42016_n2109_1), .Y(_abc_42016_n2110_1) );
  NOR2X1 NOR2X1_281 ( .A(regfil_4__3_), .B(sp_11_), .Y(_abc_42016_n2116_1) );
  NOR2X1 NOR2X1_282 ( .A(_abc_42016_n800), .B(_abc_42016_n2118), .Y(_abc_42016_n2119_1) );
  NOR2X1 NOR2X1_283 ( .A(regfil_4__1_), .B(sp_9_), .Y(_abc_42016_n2125) );
  NOR2X1 NOR2X1_284 ( .A(_abc_42016_n722), .B(_abc_42016_n2127_1), .Y(_abc_42016_n2128_1) );
  NOR2X1 NOR2X1_285 ( .A(regfil_2__7_), .B(regfil_4__7_), .Y(_abc_42016_n2146) );
  NOR2X1 NOR2X1_286 ( .A(_abc_42016_n964), .B(_abc_42016_n1801_1), .Y(_abc_42016_n2147) );
  NOR2X1 NOR2X1_287 ( .A(_abc_42016_n895), .B(_abc_42016_n1527), .Y(_abc_42016_n2151_1) );
  NOR2X1 NOR2X1_288 ( .A(regfil_2__3_), .B(regfil_4__3_), .Y(_abc_42016_n2155) );
  NOR2X1 NOR2X1_289 ( .A(_abc_42016_n796), .B(_abc_42016_n800), .Y(_abc_42016_n2157) );
  NOR2X1 NOR2X1_29 ( .A(_abc_42016_n572), .B(_abc_42016_n565), .Y(_abc_42016_n573) );
  NOR2X1 NOR2X1_290 ( .A(_abc_42016_n728), .B(_abc_42016_n722), .Y(_abc_42016_n2163) );
  NOR2X1 NOR2X1_291 ( .A(_abc_42016_n954), .B(_abc_42016_n1801_1), .Y(_abc_42016_n2179) );
  NOR2X1 NOR2X1_292 ( .A(_abc_42016_n893), .B(_abc_42016_n1527), .Y(_abc_42016_n2184) );
  NOR2X1 NOR2X1_293 ( .A(_abc_42016_n812), .B(_abc_42016_n800), .Y(_abc_42016_n2189) );
  NOR2X1 NOR2X1_294 ( .A(_abc_42016_n712), .B(_abc_42016_n722), .Y(_abc_42016_n2195) );
  NOR2X1 NOR2X1_295 ( .A(regfil_0__7_), .B(regfil_4__7_), .Y(_abc_42016_n2211) );
  NOR2X1 NOR2X1_296 ( .A(_abc_42016_n2211), .B(_abc_42016_n1035), .Y(_abc_42016_n2212) );
  NOR2X1 NOR2X1_297 ( .A(_abc_42016_n2082), .B(_abc_42016_n2222), .Y(_abc_42016_n2223) );
  NOR2X1 NOR2X1_298 ( .A(reset), .B(waitr), .Y(_abc_42016_n2226) );
  NOR2X1 NOR2X1_299 ( .A(_abc_42016_n1870), .B(_abc_42016_n507), .Y(_abc_42016_n2227) );
  NOR2X1 NOR2X1_3 ( .A(_abc_42016_n503), .B(_abc_42016_n507), .Y(_abc_42016_n508) );
  NOR2X1 NOR2X1_30 ( .A(state_2_), .B(_abc_42016_n521), .Y(_abc_42016_n575) );
  NOR2X1 NOR2X1_300 ( .A(opcode_2_), .B(_abc_42016_n1004), .Y(_abc_42016_n2253) );
  NOR2X1 NOR2X1_301 ( .A(_abc_42016_n565), .B(_abc_42016_n2254), .Y(_abc_42016_n2255) );
  NOR2X1 NOR2X1_302 ( .A(_abc_42016_n507), .B(_abc_42016_n523_1), .Y(_abc_42016_n2260) );
  NOR2X1 NOR2X1_303 ( .A(_abc_42016_n2264), .B(_abc_42016_n2262), .Y(_abc_42016_n2265) );
  NOR2X1 NOR2X1_304 ( .A(_abc_42016_n1016), .B(_abc_42016_n523_1), .Y(_abc_42016_n2266) );
  NOR2X1 NOR2X1_305 ( .A(_abc_42016_n544_1), .B(_abc_42016_n1870), .Y(_abc_42016_n2269) );
  NOR2X1 NOR2X1_306 ( .A(_abc_42016_n1923), .B(_abc_42016_n2270_1), .Y(_abc_42016_n2271_1) );
  NOR2X1 NOR2X1_307 ( .A(_abc_42016_n2268), .B(_abc_42016_n2273), .Y(_abc_42016_n2274) );
  NOR2X1 NOR2X1_308 ( .A(_abc_42016_n530), .B(_abc_42016_n533), .Y(_abc_42016_n2279) );
  NOR2X1 NOR2X1_309 ( .A(_abc_42016_n539), .B(_abc_42016_n568), .Y(_abc_42016_n2281) );
  NOR2X1 NOR2X1_31 ( .A(_abc_42016_n544_1), .B(_abc_42016_n576_1), .Y(_abc_42016_n577) );
  NOR2X1 NOR2X1_310 ( .A(_abc_42016_n2287), .B(_abc_42016_n2285), .Y(_abc_42016_n2288) );
  NOR2X1 NOR2X1_311 ( .A(_abc_42016_n2306), .B(_abc_42016_n2307), .Y(_abc_42016_n2308) );
  NOR2X1 NOR2X1_312 ( .A(opcode_5_), .B(_abc_42016_n2291), .Y(_abc_42016_n2309) );
  NOR2X1 NOR2X1_313 ( .A(opcode_2_), .B(_abc_42016_n727), .Y(_abc_42016_n2317) );
  NOR2X1 NOR2X1_314 ( .A(_abc_42016_n2317), .B(_abc_42016_n1001_1), .Y(_abc_42016_n2318) );
  NOR2X1 NOR2X1_315 ( .A(_abc_42016_n2319), .B(_abc_42016_n2316), .Y(_abc_42016_n2320) );
  NOR2X1 NOR2X1_316 ( .A(_abc_42016_n2306), .B(_abc_42016_n2323_1), .Y(_abc_42016_n2324_1) );
  NOR2X1 NOR2X1_317 ( .A(_abc_42016_n1377), .B(_abc_42016_n2325), .Y(_abc_42016_n2326) );
  NOR2X1 NOR2X1_318 ( .A(_abc_42016_n2327), .B(_abc_42016_n2321), .Y(_abc_42016_n2328) );
  NOR2X1 NOR2X1_319 ( .A(_abc_42016_n2031), .B(_abc_42016_n546), .Y(_abc_42016_n2334) );
  NOR2X1 NOR2X1_32 ( .A(_abc_42016_n513), .B(_abc_42016_n578), .Y(_abc_42016_n579) );
  NOR2X1 NOR2X1_320 ( .A(_abc_42016_n2338), .B(_abc_42016_n2335), .Y(_abc_42016_n2339) );
  NOR2X1 NOR2X1_321 ( .A(_abc_42016_n572), .B(_abc_42016_n626), .Y(_abc_42016_n2347_1) );
  NOR2X1 NOR2X1_322 ( .A(statesel_0_), .B(_abc_42016_n2344), .Y(_abc_42016_n2363) );
  NOR2X1 NOR2X1_323 ( .A(statesel_1_), .B(_abc_42016_n2259), .Y(_abc_42016_n2364) );
  NOR2X1 NOR2X1_324 ( .A(_abc_42016_n2278), .B(_abc_42016_n2366), .Y(_abc_42016_n2367) );
  NOR2X1 NOR2X1_325 ( .A(_abc_42016_n2355), .B(_abc_42016_n1004), .Y(_abc_42016_n2370) );
  NOR2X1 NOR2X1_326 ( .A(_abc_42016_n2325), .B(_abc_42016_n2316), .Y(_abc_42016_n2383) );
  NOR2X1 NOR2X1_327 ( .A(_abc_42016_n2259), .B(_abc_42016_n2344), .Y(_abc_42016_n2387) );
  NOR2X1 NOR2X1_328 ( .A(_abc_42016_n1863), .B(_abc_42016_n1848), .Y(_abc_42016_n2403) );
  NOR2X1 NOR2X1_329 ( .A(statesel_3_), .B(_abc_42016_n2369), .Y(_abc_42016_n2408_1) );
  NOR2X1 NOR2X1_33 ( .A(_abc_42016_n503), .B(_abc_42016_n520), .Y(_abc_42016_n580) );
  NOR2X1 NOR2X1_330 ( .A(_abc_42016_n2409), .B(_abc_42016_n2407), .Y(_abc_42016_n2410) );
  NOR2X1 NOR2X1_331 ( .A(_abc_42016_n1377), .B(_abc_42016_n2418), .Y(_abc_42016_n2419) );
  NOR2X1 NOR2X1_332 ( .A(_abc_42016_n2369), .B(_abc_42016_n2394_1), .Y(_abc_42016_n2436) );
  NOR2X1 NOR2X1_333 ( .A(_abc_42016_n2407), .B(_abc_42016_n2437), .Y(_abc_42016_n2438_1) );
  NOR2X1 NOR2X1_334 ( .A(statesel_4_), .B(_abc_42016_n2438_1), .Y(_abc_42016_n2439) );
  NOR2X1 NOR2X1_335 ( .A(_abc_42016_n2417_1), .B(_abc_42016_n2440), .Y(_abc_42016_n2441_1) );
  NOR2X1 NOR2X1_336 ( .A(_abc_42016_n2439), .B(_abc_42016_n2441_1), .Y(_abc_42016_n2442) );
  NOR2X1 NOR2X1_337 ( .A(statesel_5_), .B(_abc_42016_n2417_1), .Y(_abc_42016_n2450_1) );
  NOR2X1 NOR2X1_338 ( .A(_abc_42016_n2451), .B(_abc_42016_n2440), .Y(_abc_42016_n2452) );
  NOR2X1 NOR2X1_339 ( .A(_abc_42016_n1508), .B(_abc_42016_n1438), .Y(_abc_42016_n2501) );
  NOR2X1 NOR2X1_34 ( .A(_abc_42016_n518_1), .B(_abc_42016_n581_1), .Y(_abc_42016_n582_1) );
  NOR2X1 NOR2X1_340 ( .A(opcode_5_), .B(_abc_42016_n1904), .Y(_abc_42016_n2502) );
  NOR2X1 NOR2X1_341 ( .A(_abc_42016_n2496), .B(_abc_42016_n1411), .Y(_abc_42016_n2507) );
  NOR2X1 NOR2X1_342 ( .A(_abc_42016_n560), .B(_abc_42016_n1347), .Y(_abc_42016_n2512) );
  NOR2X1 NOR2X1_343 ( .A(_abc_42016_n1923), .B(_abc_42016_n509), .Y(_abc_42016_n2518_1) );
  NOR2X1 NOR2X1_344 ( .A(pc_1_), .B(pc_0_), .Y(_abc_42016_n2524) );
  NOR2X1 NOR2X1_345 ( .A(_abc_42016_n1383), .B(_abc_42016_n1381), .Y(_abc_42016_n2525) );
  NOR2X1 NOR2X1_346 ( .A(_abc_42016_n2524), .B(_abc_42016_n2525), .Y(_abc_42016_n2526) );
  NOR2X1 NOR2X1_347 ( .A(regfil_5__1_), .B(_abc_42016_n669), .Y(_abc_42016_n2529) );
  NOR2X1 NOR2X1_348 ( .A(_abc_42016_n2529), .B(_abc_42016_n1400), .Y(_abc_42016_n2530) );
  NOR2X1 NOR2X1_349 ( .A(_abc_42016_n2526), .B(_abc_42016_n1378), .Y(_abc_42016_n2535) );
  NOR2X1 NOR2X1_35 ( .A(popdes_0_), .B(_abc_42016_n583), .Y(_abc_42016_n584_1) );
  NOR2X1 NOR2X1_350 ( .A(_abc_42016_n674), .B(_abc_42016_n1411), .Y(_abc_42016_n2539) );
  NOR2X1 NOR2X1_351 ( .A(pc_2_), .B(pc_1_), .Y(_abc_42016_n2572) );
  NOR2X1 NOR2X1_352 ( .A(pc_3_), .B(_abc_42016_n2571), .Y(_abc_42016_n2588) );
  NOR2X1 NOR2X1_353 ( .A(_abc_42016_n1359), .B(_abc_42016_n2588), .Y(_abc_42016_n2589) );
  NOR2X1 NOR2X1_354 ( .A(_abc_42016_n1139), .B(_abc_42016_n669), .Y(_abc_42016_n2593) );
  NOR2X1 NOR2X1_355 ( .A(_abc_42016_n2595), .B(_abc_42016_n2600), .Y(_abc_42016_n2601) );
  NOR2X1 NOR2X1_356 ( .A(_abc_42016_n2499), .B(_abc_42016_n2616), .Y(_abc_42016_n2617) );
  NOR2X1 NOR2X1_357 ( .A(opcode_5_), .B(_abc_42016_n2622), .Y(_abc_42016_n2623) );
  NOR2X1 NOR2X1_358 ( .A(_abc_42016_n2536), .B(_abc_42016_n2660), .Y(_abc_42016_n2661) );
  NOR2X1 NOR2X1_359 ( .A(_abc_42016_n2499), .B(_abc_42016_n2671), .Y(_abc_42016_n2672_1) );
  NOR2X1 NOR2X1_36 ( .A(popdes_1_), .B(_abc_42016_n585), .Y(_abc_42016_n586) );
  NOR2X1 NOR2X1_360 ( .A(_abc_42016_n1380), .B(_abc_42016_n2676), .Y(_abc_42016_n2677) );
  NOR2X1 NOR2X1_361 ( .A(_abc_42016_n2031), .B(_abc_42016_n2079), .Y(_abc_42016_n2732) );
  NOR2X1 NOR2X1_362 ( .A(_abc_42016_n1879_1), .B(_abc_42016_n2426_1), .Y(_abc_42016_n2737) );
  NOR2X1 NOR2X1_363 ( .A(_abc_42016_n2347_1), .B(_abc_42016_n2319), .Y(_abc_42016_n2739) );
  NOR2X1 NOR2X1_364 ( .A(_abc_42016_n2323_1), .B(_abc_42016_n2741), .Y(_abc_42016_n2742) );
  NOR2X1 NOR2X1_365 ( .A(_abc_42016_n2740), .B(_abc_42016_n2743), .Y(_abc_42016_n2744) );
  NOR2X1 NOR2X1_366 ( .A(_abc_42016_n2280), .B(_abc_42016_n2748_1), .Y(_abc_42016_n2750) );
  NOR2X1 NOR2X1_367 ( .A(_abc_42016_n2731), .B(_abc_42016_n2765), .Y(_abc_42016_n2777) );
  NOR2X1 NOR2X1_368 ( .A(_abc_42016_n2731), .B(_abc_42016_n2733), .Y(_abc_42016_n2779) );
  NOR2X1 NOR2X1_369 ( .A(_abc_42016_n2765), .B(_abc_42016_n2733), .Y(_abc_42016_n2780) );
  NOR2X1 NOR2X1_37 ( .A(_abc_42016_n579), .B(_abc_42016_n586), .Y(_abc_42016_n587) );
  NOR2X1 NOR2X1_370 ( .A(_abc_42016_n2562), .B(_abc_42016_n2425), .Y(_abc_42016_n2794) );
  NOR2X1 NOR2X1_371 ( .A(_abc_42016_n2803), .B(_abc_42016_n2787), .Y(_abc_42016_n2804) );
  NOR2X1 NOR2X1_372 ( .A(_abc_42016_n2804), .B(_abc_42016_n2733), .Y(_abc_42016_n2805) );
  NOR2X1 NOR2X1_373 ( .A(_abc_42016_n2735), .B(_abc_42016_n2807), .Y(_abc_42016_n2808) );
  NOR2X1 NOR2X1_374 ( .A(regfil_5__3_), .B(_abc_42016_n2280), .Y(_abc_42016_n2810_1) );
  NOR2X1 NOR2X1_375 ( .A(_abc_42016_n2622), .B(_abc_42016_n2310), .Y(_abc_42016_n2823) );
  NOR2X1 NOR2X1_376 ( .A(regfil_5__5_), .B(_abc_42016_n2280), .Y(_abc_42016_n2838) );
  NOR2X1 NOR2X1_377 ( .A(_abc_42016_n1909_1), .B(_abc_42016_n2838), .Y(_abc_42016_n2839) );
  NOR2X1 NOR2X1_378 ( .A(_abc_42016_n2836), .B(_abc_42016_n2828), .Y(_abc_42016_n2847) );
  NOR2X1 NOR2X1_379 ( .A(_abc_42016_n2852), .B(_abc_42016_n2747_1), .Y(_abc_42016_n2853) );
  NOR2X1 NOR2X1_38 ( .A(_abc_42016_n591), .B(_abc_42016_n588_1), .Y(_abc_42016_n592_1) );
  NOR2X1 NOR2X1_380 ( .A(_abc_42016_n2678), .B(_abc_42016_n2291), .Y(_abc_42016_n2854) );
  NOR2X1 NOR2X1_381 ( .A(regfil_5__6_), .B(_abc_42016_n2280), .Y(_abc_42016_n2855_1) );
  NOR2X1 NOR2X1_382 ( .A(_abc_42016_n1837_1), .B(_abc_42016_n2855_1), .Y(_abc_42016_n2856_1) );
  NOR2X1 NOR2X1_383 ( .A(_abc_42016_n2869), .B(_abc_42016_n2880), .Y(_abc_42016_n2881) );
  NOR2X1 NOR2X1_384 ( .A(_abc_42016_n2887), .B(_abc_42016_n2882), .Y(_abc_42016_n2888) );
  NOR2X1 NOR2X1_385 ( .A(_abc_42016_n2887), .B(_abc_42016_n2747_1), .Y(_abc_42016_n2892) );
  NOR2X1 NOR2X1_386 ( .A(_abc_42016_n1428), .B(_abc_42016_n2291), .Y(_abc_42016_n2902) );
  NOR2X1 NOR2X1_387 ( .A(regfil_4__1_), .B(_abc_42016_n2280), .Y(_abc_42016_n2903) );
  NOR2X1 NOR2X1_388 ( .A(regfil_4__2_), .B(_abc_42016_n2280), .Y(_abc_42016_n2922) );
  NOR2X1 NOR2X1_389 ( .A(_abc_42016_n2924_1), .B(_abc_42016_n2737), .Y(_abc_42016_n2925_1) );
  NOR2X1 NOR2X1_39 ( .A(_abc_42016_n596), .B(_abc_42016_n588_1), .Y(_abc_42016_n597_1) );
  NOR2X1 NOR2X1_390 ( .A(_abc_42016_n1446), .B(_abc_42016_n2754), .Y(_abc_42016_n2930) );
  NOR2X1 NOR2X1_391 ( .A(_abc_42016_n2920), .B(_abc_42016_n2912), .Y(_abc_42016_n2934) );
  NOR2X1 NOR2X1_392 ( .A(_abc_42016_n2425), .B(_abc_42016_n1481), .Y(_abc_42016_n2941) );
  NOR2X1 NOR2X1_393 ( .A(regfil_4__3_), .B(_abc_42016_n2280), .Y(_abc_42016_n2943) );
  NOR2X1 NOR2X1_394 ( .A(_abc_42016_n2942), .B(_abc_42016_n2935), .Y(_abc_42016_n2951) );
  NOR2X1 NOR2X1_395 ( .A(_abc_42016_n2427), .B(_abc_42016_n2961), .Y(_abc_42016_n2962) );
  NOR2X1 NOR2X1_396 ( .A(_abc_42016_n2969_1), .B(_abc_42016_n2968), .Y(_abc_42016_n2970_1) );
  NOR2X1 NOR2X1_397 ( .A(_abc_42016_n2972), .B(_abc_42016_n2983), .Y(_abc_42016_n2984) );
  NOR2X1 NOR2X1_398 ( .A(_abc_42016_n1554), .B(_abc_42016_n2754), .Y(_abc_42016_n2991_1) );
  NOR2X1 NOR2X1_399 ( .A(_abc_42016_n2995), .B(_abc_42016_n2737), .Y(_abc_42016_n2996) );
  NOR2X1 NOR2X1_4 ( .A(state_5_), .B(state_4_), .Y(_abc_42016_n510) );
  NOR2X1 NOR2X1_40 ( .A(_abc_42016_n597_1), .B(_abc_42016_n593), .Y(_abc_42016_n598_1) );
  NOR2X1 NOR2X1_400 ( .A(_abc_42016_n2990_1), .B(_abc_42016_n2985), .Y(_abc_42016_n3003) );
  NOR2X1 NOR2X1_401 ( .A(_abc_42016_n2101), .B(_abc_42016_n2739), .Y(_abc_42016_n3018) );
  NOR2X1 NOR2X1_402 ( .A(_abc_42016_n2759), .B(_abc_42016_n1587), .Y(_abc_42016_n3019) );
  NOR2X1 NOR2X1_403 ( .A(_abc_42016_n2518_1), .B(_abc_42016_n2498), .Y(_abc_42016_n3029) );
  NOR2X1 NOR2X1_404 ( .A(opcode_5_), .B(_abc_42016_n1347), .Y(_abc_42016_n3033) );
  NOR2X1 NOR2X1_405 ( .A(_abc_42016_n1904), .B(_abc_42016_n3034), .Y(_abc_42016_n3035_1) );
  NOR2X1 NOR2X1_406 ( .A(_abc_42016_n695), .B(_abc_42016_n2280), .Y(_abc_42016_n3039) );
  NOR2X1 NOR2X1_407 ( .A(_abc_42016_n3047), .B(_abc_42016_n3031), .Y(_abc_42016_n3048) );
  NOR2X1 NOR2X1_408 ( .A(_abc_42016_n3054), .B(_abc_42016_n1402), .Y(_abc_42016_n3055) );
  NOR2X1 NOR2X1_409 ( .A(_abc_42016_n1851), .B(_abc_42016_n3065), .Y(_abc_42016_n3066) );
  NOR2X1 NOR2X1_41 ( .A(_abc_42016_n556), .B(_abc_42016_n599), .Y(_abc_42016_n600) );
  NOR2X1 NOR2X1_410 ( .A(_abc_42016_n3028), .B(_abc_42016_n3050), .Y(_abc_42016_n3073) );
  NOR2X1 NOR2X1_411 ( .A(_abc_42016_n3071), .B(_abc_42016_n3075), .Y(_abc_42016_n3076) );
  NOR2X1 NOR2X1_412 ( .A(_abc_42016_n1841), .B(_abc_42016_n3087), .Y(_abc_42016_n3093) );
  NOR2X1 NOR2X1_413 ( .A(sp_1_), .B(sp_2_), .Y(_abc_42016_n3097) );
  NOR2X1 NOR2X1_414 ( .A(_abc_42016_n2775), .B(_abc_42016_n1159), .Y(_abc_42016_n3098) );
  NOR2X1 NOR2X1_415 ( .A(_abc_42016_n3097), .B(_abc_42016_n3098), .Y(_abc_42016_n3099) );
  NOR2X1 NOR2X1_416 ( .A(_abc_42016_n3105_1), .B(_abc_42016_n3082), .Y(_abc_42016_n3107) );
  NOR2X1 NOR2X1_417 ( .A(_abc_42016_n3105_1), .B(_abc_42016_n2293), .Y(_abc_42016_n3111) );
  NOR2X1 NOR2X1_418 ( .A(_abc_42016_n1851), .B(_abc_42016_n3117), .Y(_abc_42016_n3118) );
  NOR2X1 NOR2X1_419 ( .A(sp_3_), .B(_abc_42016_n3119), .Y(_abc_42016_n3120) );
  NOR2X1 NOR2X1_42 ( .A(_abc_42016_n604_1), .B(_abc_42016_n603), .Y(_abc_42016_n605_1) );
  NOR2X1 NOR2X1_420 ( .A(_abc_42016_n3128), .B(_abc_42016_n1411), .Y(_abc_42016_n3129) );
  NOR2X1 NOR2X1_421 ( .A(waddrhold_4_), .B(_abc_42016_n2279), .Y(_abc_42016_n3137) );
  NOR2X1 NOR2X1_422 ( .A(_abc_42016_n3128), .B(_abc_42016_n3146), .Y(_abc_42016_n3147_1) );
  NOR2X1 NOR2X1_423 ( .A(_abc_42016_n1841), .B(_abc_42016_n3154), .Y(_abc_42016_n3158) );
  NOR2X1 NOR2X1_424 ( .A(_abc_42016_n1851), .B(_abc_42016_n3160), .Y(_abc_42016_n3161) );
  NOR2X1 NOR2X1_425 ( .A(sp_5_), .B(_abc_42016_n3131), .Y(_abc_42016_n3163) );
  NOR2X1 NOR2X1_426 ( .A(_abc_42016_n3162), .B(_abc_42016_n3163), .Y(_abc_42016_n3164) );
  NOR2X1 NOR2X1_427 ( .A(_abc_42016_n3164), .B(_abc_42016_n3130), .Y(_abc_42016_n3165) );
  NOR2X1 NOR2X1_428 ( .A(_abc_42016_n1279), .B(_abc_42016_n1061), .Y(_abc_42016_n3166) );
  NOR2X1 NOR2X1_429 ( .A(_abc_42016_n3175), .B(_abc_42016_n1411), .Y(_abc_42016_n3176) );
  NOR2X1 NOR2X1_43 ( .A(regfil_1__0_), .B(regfil_1__1_), .Y(_abc_42016_n612) );
  NOR2X1 NOR2X1_430 ( .A(sp_5_), .B(sp_6_), .Y(_abc_42016_n3177) );
  NOR2X1 NOR2X1_431 ( .A(_abc_42016_n3178), .B(_abc_42016_n3131), .Y(_abc_42016_n3179) );
  NOR2X1 NOR2X1_432 ( .A(waddrhold_6_), .B(_abc_42016_n2279), .Y(_abc_42016_n3185) );
  NOR2X1 NOR2X1_433 ( .A(_abc_42016_n1848), .B(_abc_42016_n2855_1), .Y(_abc_42016_n3186) );
  NOR2X1 NOR2X1_434 ( .A(sp_7_), .B(_abc_42016_n3180), .Y(_abc_42016_n3202) );
  NOR2X1 NOR2X1_435 ( .A(_abc_42016_n1327_1), .B(_abc_42016_n3179), .Y(_abc_42016_n3203) );
  NOR2X1 NOR2X1_436 ( .A(_abc_42016_n2718), .B(_abc_42016_n3034), .Y(_abc_42016_n3207) );
  NOR2X1 NOR2X1_437 ( .A(_abc_42016_n3201), .B(_abc_42016_n3194), .Y(_abc_42016_n3216) );
  NOR2X1 NOR2X1_438 ( .A(_abc_42016_n2131_1), .B(_abc_42016_n3202), .Y(_abc_42016_n3226) );
  NOR2X1 NOR2X1_439 ( .A(_abc_42016_n1395), .B(_abc_42016_n3034), .Y(_abc_42016_n3230) );
  NOR2X1 NOR2X1_44 ( .A(regfil_1__3_), .B(_abc_42016_n613), .Y(_abc_42016_n614) );
  NOR2X1 NOR2X1_440 ( .A(_abc_42016_n3223), .B(_abc_42016_n3217_1), .Y(_abc_42016_n3238) );
  NOR2X1 NOR2X1_441 ( .A(_abc_42016_n2127_1), .B(_abc_42016_n3225), .Y(_abc_42016_n3247) );
  NOR2X1 NOR2X1_442 ( .A(sp_9_), .B(_abc_42016_n3224), .Y(_abc_42016_n3248) );
  NOR2X1 NOR2X1_443 ( .A(_abc_42016_n3248), .B(_abc_42016_n3247), .Y(_abc_42016_n3249) );
  NOR2X1 NOR2X1_444 ( .A(_abc_42016_n1428), .B(_abc_42016_n1347), .Y(_abc_42016_n3255) );
  NOR2X1 NOR2X1_445 ( .A(_abc_42016_n1456), .B(_abc_42016_n3034), .Y(_abc_42016_n3275) );
  NOR2X1 NOR2X1_446 ( .A(_abc_42016_n1848), .B(_abc_42016_n2922), .Y(_abc_42016_n3276) );
  NOR2X1 NOR2X1_447 ( .A(_abc_42016_n3268), .B(_abc_42016_n3264), .Y(_abc_42016_n3285) );
  NOR2X1 NOR2X1_448 ( .A(_abc_42016_n2497), .B(_abc_42016_n3285), .Y(_abc_42016_n3286) );
  NOR2X1 NOR2X1_449 ( .A(sp_11_), .B(_abc_42016_n3269), .Y(_abc_42016_n3295_1) );
  NOR2X1 NOR2X1_45 ( .A(regfil_1__5_), .B(_abc_42016_n615), .Y(_abc_42016_n616) );
  NOR2X1 NOR2X1_450 ( .A(waddrhold_12_), .B(_abc_42016_n2279), .Y(_abc_42016_n3326) );
  NOR2X1 NOR2X1_451 ( .A(sp_13_), .B(_abc_42016_n3319_1), .Y(_abc_42016_n3339) );
  NOR2X1 NOR2X1_452 ( .A(_abc_42016_n3316), .B(_abc_42016_n3309), .Y(_abc_42016_n3354) );
  NOR2X1 NOR2X1_453 ( .A(_abc_42016_n3358), .B(_abc_42016_n3356), .Y(_abc_42016_n3359) );
  NOR2X1 NOR2X1_454 ( .A(sp_14_), .B(_abc_42016_n3340), .Y(_abc_42016_n3362) );
  NOR2X1 NOR2X1_455 ( .A(_abc_42016_n3371), .B(_abc_42016_n3373), .Y(_abc_42016_n3374) );
  NOR2X1 NOR2X1_456 ( .A(_abc_42016_n3361), .B(_abc_42016_n3380), .Y(_abc_42016_n3381) );
  NOR2X1 NOR2X1_457 ( .A(waddrhold_15_), .B(_abc_42016_n2279), .Y(_abc_42016_n3394) );
  NOR2X1 NOR2X1_458 ( .A(reset), .B(_abc_42016_n2497), .Y(_abc_42016_n3407) );
  NOR2X1 NOR2X1_459 ( .A(_abc_42016_n518_1), .B(_abc_42016_n667), .Y(_abc_42016_n3409) );
  NOR2X1 NOR2X1_46 ( .A(regfil_1__7_), .B(_abc_42016_n617), .Y(_abc_42016_n618) );
  NOR2X1 NOR2X1_460 ( .A(_abc_42016_n2031), .B(_abc_42016_n667), .Y(_abc_42016_n3410) );
  NOR2X1 NOR2X1_461 ( .A(opcode_7_), .B(_abc_42016_n558), .Y(_abc_42016_n3429) );
  NOR2X1 NOR2X1_462 ( .A(_abc_42016_n1849), .B(_abc_42016_n3442), .Y(_abc_42016_n3443) );
  NOR2X1 NOR2X1_463 ( .A(_abc_42016_n674), .B(_abc_42016_n1022), .Y(_abc_42016_n3452) );
  NOR2X1 NOR2X1_464 ( .A(_abc_42016_n560), .B(_abc_42016_n3453), .Y(_abc_42016_n3455) );
  NOR2X1 NOR2X1_465 ( .A(_abc_42016_n576_1), .B(_abc_42016_n507), .Y(_abc_42016_n3457) );
  NOR2X1 NOR2X1_466 ( .A(_abc_42016_n2306), .B(_abc_42016_n1005), .Y(_abc_42016_n3469) );
  NOR2X1 NOR2X1_467 ( .A(_abc_42016_n1004), .B(_abc_42016_n682), .Y(_abc_42016_n3474) );
  NOR2X1 NOR2X1_468 ( .A(_abc_42016_n3483), .B(_abc_42016_n3462), .Y(_abc_42016_n3484) );
  NOR2X1 NOR2X1_469 ( .A(_abc_42016_n1923), .B(_abc_42016_n546), .Y(_abc_42016_n3502) );
  NOR2X1 NOR2X1_47 ( .A(_abc_42016_n608), .B(_abc_42016_n618), .Y(_abc_42016_n621) );
  NOR2X1 NOR2X1_470 ( .A(sp_0_), .B(_abc_42016_n3121), .Y(_abc_42016_n3514) );
  NOR2X1 NOR2X1_471 ( .A(_abc_42016_n2758), .B(_abc_42016_n3509), .Y(_abc_42016_n3519) );
  NOR2X1 NOR2X1_472 ( .A(_abc_42016_n3462), .B(_abc_42016_n3529), .Y(_abc_42016_n3530) );
  NOR2X1 NOR2X1_473 ( .A(_abc_42016_n1210), .B(_abc_42016_n3509), .Y(_abc_42016_n3533) );
  NOR2X1 NOR2X1_474 ( .A(_abc_42016_n1210), .B(_abc_42016_n3514), .Y(_abc_42016_n3541) );
  NOR2X1 NOR2X1_475 ( .A(sp_0_), .B(_abc_42016_n3131), .Y(_abc_42016_n3542) );
  NOR2X1 NOR2X1_476 ( .A(_abc_42016_n1279), .B(_abc_42016_n3534), .Y(_abc_42016_n3555) );
  NOR2X1 NOR2X1_477 ( .A(_abc_42016_n3554), .B(_abc_42016_n3559), .Y(_abc_42016_n3560) );
  NOR2X1 NOR2X1_478 ( .A(_abc_42016_n566), .B(_abc_42016_n3562), .Y(_abc_42016_n3566) );
  NOR2X1 NOR2X1_479 ( .A(_abc_42016_n3576), .B(_abc_42016_n3578), .Y(_abc_42016_n3579) );
  NOR2X1 NOR2X1_48 ( .A(opcode_1_), .B(_abc_42016_n563), .Y(_abc_42016_n625) );
  NOR2X1 NOR2X1_480 ( .A(_abc_42016_n2758), .B(_abc_42016_n3583), .Y(_abc_42016_n3594) );
  NOR2X1 NOR2X1_481 ( .A(_abc_42016_n3475), .B(_abc_42016_n3594), .Y(_abc_42016_n3595) );
  NOR2X1 NOR2X1_482 ( .A(_abc_42016_n3575), .B(_abc_42016_n3584), .Y(_abc_42016_n3600) );
  NOR2X1 NOR2X1_483 ( .A(_abc_42016_n3600), .B(_abc_42016_n3602), .Y(_abc_42016_n3603) );
  NOR2X1 NOR2X1_484 ( .A(_abc_42016_n3203), .B(_abc_42016_n3202), .Y(_abc_42016_n3605) );
  NOR2X1 NOR2X1_485 ( .A(_abc_42016_n1327_1), .B(_abc_42016_n3583), .Y(_abc_42016_n3606_1) );
  NOR2X1 NOR2X1_486 ( .A(_abc_42016_n1327_1), .B(_abc_42016_n3590), .Y(_abc_42016_n3613) );
  NOR2X1 NOR2X1_487 ( .A(sp_7_), .B(_abc_42016_n3589), .Y(_abc_42016_n3614) );
  NOR2X1 NOR2X1_488 ( .A(sp_0_), .B(_abc_42016_n3224), .Y(_abc_42016_n3627) );
  NOR2X1 NOR2X1_489 ( .A(_abc_42016_n3475), .B(_abc_42016_n3630), .Y(_abc_42016_n3631) );
  NOR2X1 NOR2X1_49 ( .A(opcode_0_), .B(opcode_1_), .Y(_abc_42016_n630) );
  NOR2X1 NOR2X1_490 ( .A(sp_0_), .B(_abc_42016_n3293), .Y(_abc_42016_n3649) );
  NOR2X1 NOR2X1_491 ( .A(_abc_42016_n2127_1), .B(_abc_42016_n3627), .Y(_abc_42016_n3650) );
  NOR2X1 NOR2X1_492 ( .A(_abc_42016_n2127_1), .B(_abc_42016_n3629), .Y(_abc_42016_n3652) );
  NOR2X1 NOR2X1_493 ( .A(_abc_42016_n2376), .B(_abc_42016_n3659), .Y(_abc_42016_n3660) );
  NOR2X1 NOR2X1_494 ( .A(sp_0_), .B(_abc_42016_n3269), .Y(_abc_42016_n3671) );
  NOR2X1 NOR2X1_495 ( .A(_abc_42016_n3692), .B(_abc_42016_n3629), .Y(_abc_42016_n3693) );
  NOR2X1 NOR2X1_496 ( .A(_abc_42016_n2118), .B(_abc_42016_n3671), .Y(_abc_42016_n3698) );
  NOR2X1 NOR2X1_497 ( .A(sp_0_), .B(_abc_42016_n3296_1), .Y(_abc_42016_n3699) );
  NOR2X1 NOR2X1_498 ( .A(_abc_42016_n2758), .B(_abc_42016_n3694), .Y(_abc_42016_n3702) );
  NOR2X1 NOR2X1_499 ( .A(sp_0_), .B(_abc_42016_n3319_1), .Y(_abc_42016_n3713_1) );
  NOR2X1 NOR2X1_5 ( .A(reset), .B(_abc_42016_n511), .Y(_abc_42016_n512) );
  NOR2X1 NOR2X1_50 ( .A(_abc_42016_n644), .B(_abc_42016_n645), .Y(_abc_42016_n646) );
  NOR2X1 NOR2X1_500 ( .A(sp_12_), .B(_abc_42016_n3702), .Y(_abc_42016_n3717) );
  NOR2X1 NOR2X1_501 ( .A(_abc_42016_n3717), .B(_abc_42016_n3719), .Y(_abc_42016_n3720) );
  NOR2X1 NOR2X1_502 ( .A(_abc_42016_n1408), .B(_abc_42016_n3321), .Y(_abc_42016_n3723) );
  NOR2X1 NOR2X1_503 ( .A(_abc_42016_n2113), .B(_abc_42016_n3694), .Y(_abc_42016_n3725) );
  NOR2X1 NOR2X1_504 ( .A(_abc_42016_n3453), .B(_abc_42016_n3718), .Y(_abc_42016_n3738) );
  NOR2X1 NOR2X1_505 ( .A(sp_0_), .B(_abc_42016_n3340), .Y(_abc_42016_n3741) );
  NOR2X1 NOR2X1_506 ( .A(_abc_42016_n2109_1), .B(_abc_42016_n3713_1), .Y(_abc_42016_n3742) );
  NOR2X1 NOR2X1_507 ( .A(sp_13_), .B(_abc_42016_n3725), .Y(_abc_42016_n3745) );
  NOR2X1 NOR2X1_508 ( .A(_abc_42016_n2109_1), .B(_abc_42016_n3726), .Y(_abc_42016_n3746) );
  NOR2X1 NOR2X1_509 ( .A(_abc_42016_n3745), .B(_abc_42016_n3746), .Y(_abc_42016_n3747) );
  NOR2X1 NOR2X1_51 ( .A(_abc_42016_n642), .B(_abc_42016_n649_1), .Y(_abc_42016_n650) );
  NOR2X1 NOR2X1_510 ( .A(sp_0_), .B(_abc_42016_n3363), .Y(_abc_42016_n3758) );
  NOR2X1 NOR2X1_511 ( .A(_abc_42016_n2103), .B(_abc_42016_n3741), .Y(_abc_42016_n3759) );
  NOR2X1 NOR2X1_512 ( .A(_abc_42016_n2758), .B(_abc_42016_n3762), .Y(_abc_42016_n3763) );
  NOR2X1 NOR2X1_513 ( .A(_abc_42016_n3475), .B(_abc_42016_n3763), .Y(_abc_42016_n3764) );
  NOR2X1 NOR2X1_514 ( .A(_abc_42016_n2103), .B(_abc_42016_n2255), .Y(_abc_42016_n3765) );
  NOR2X1 NOR2X1_515 ( .A(_abc_42016_n3775_1), .B(_abc_42016_n3776), .Y(_abc_42016_n3777) );
  NOR2X1 NOR2X1_516 ( .A(_abc_42016_n2101), .B(_abc_42016_n3758), .Y(_abc_42016_n3781) );
  NOR2X1 NOR2X1_517 ( .A(_abc_42016_n2101), .B(_abc_42016_n3763), .Y(_abc_42016_n3784) );
  NOR2X1 NOR2X1_518 ( .A(_abc_42016_n1604_1), .B(_abc_42016_n988), .Y(_abc_42016_n3800) );
  NOR2X1 NOR2X1_519 ( .A(_abc_42016_n1047_1), .B(_abc_42016_n3803), .Y(_abc_42016_n3804) );
  NOR2X1 NOR2X1_52 ( .A(_abc_42016_n608), .B(_abc_42016_n653), .Y(_abc_42016_n654) );
  NOR2X1 NOR2X1_520 ( .A(_abc_42016_n722), .B(_abc_42016_n3810), .Y(_abc_42016_n3838) );
  NOR2X1 NOR2X1_521 ( .A(regfil_4__1_), .B(_abc_42016_n3806), .Y(_abc_42016_n3856) );
  NOR2X1 NOR2X1_522 ( .A(_abc_42016_n3836), .B(_abc_42016_n3859_1), .Y(_abc_42016_n3860) );
  NOR2X1 NOR2X1_523 ( .A(rdatahold_2_), .B(_abc_42016_n994), .Y(_abc_42016_n3866) );
  NOR2X1 NOR2X1_524 ( .A(_abc_42016_n3879), .B(_abc_42016_n3878), .Y(_abc_42016_n3880) );
  NOR2X1 NOR2X1_525 ( .A(_abc_42016_n1125), .B(_abc_42016_n3888), .Y(_abc_42016_n3889) );
  NOR2X1 NOR2X1_526 ( .A(_abc_42016_n671_1), .B(_abc_42016_n3890), .Y(_abc_42016_n3891) );
  NOR2X1 NOR2X1_527 ( .A(regfil_4__3_), .B(_abc_42016_n3800), .Y(_abc_42016_n3896) );
  NOR2X1 NOR2X1_528 ( .A(regfil_4__3_), .B(_abc_42016_n3867), .Y(_abc_42016_n3898) );
  NOR2X1 NOR2X1_529 ( .A(_abc_42016_n1170), .B(_abc_42016_n3898), .Y(_abc_42016_n3899) );
  NOR2X1 NOR2X1_53 ( .A(_abc_42016_n569), .B(_abc_42016_n562), .Y(_abc_42016_n658) );
  NOR2X1 NOR2X1_530 ( .A(_abc_42016_n800), .B(_abc_42016_n3872), .Y(_abc_42016_n3907) );
  NOR2X1 NOR2X1_531 ( .A(_abc_42016_n2116_1), .B(_abc_42016_n2119_1), .Y(_abc_42016_n3916) );
  NOR2X1 NOR2X1_532 ( .A(rdatahold_4_), .B(_abc_42016_n994), .Y(_abc_42016_n3928) );
  NOR2X1 NOR2X1_533 ( .A(_abc_42016_n800), .B(_abc_42016_n1046), .Y(_abc_42016_n3935_1) );
  NOR2X1 NOR2X1_534 ( .A(_abc_42016_n1170), .B(_abc_42016_n3948), .Y(_abc_42016_n3949) );
  NOR2X1 NOR2X1_535 ( .A(regfil_4__5_), .B(_abc_42016_n3947), .Y(_abc_42016_n3958) );
  NOR2X1 NOR2X1_536 ( .A(_abc_42016_n2107), .B(_abc_42016_n2110_1), .Y(_abc_42016_n3972) );
  NOR2X1 NOR2X1_537 ( .A(regfil_4__5_), .B(_abc_42016_n3933), .Y(_abc_42016_n3977) );
  NOR2X1 NOR2X1_538 ( .A(_abc_42016_n1187), .B(_abc_42016_n3977), .Y(_abc_42016_n3978) );
  NOR2X1 NOR2X1_539 ( .A(_abc_42016_n3995), .B(_abc_42016_n3994), .Y(_abc_42016_n3996) );
  NOR2X1 NOR2X1_54 ( .A(_abc_42016_n623), .B(_abc_42016_n662), .Y(_abc_42016_n663) );
  NOR2X1 NOR2X1_540 ( .A(_abc_42016_n2149), .B(_abc_42016_n3997), .Y(_abc_42016_n3998) );
  NOR2X1 NOR2X1_541 ( .A(_abc_42016_n1554), .B(_abc_42016_n3976), .Y(_abc_42016_n4000) );
  NOR2X1 NOR2X1_542 ( .A(_abc_42016_n2211), .B(_abc_42016_n2179), .Y(_abc_42016_n4016) );
  NOR2X1 NOR2X1_543 ( .A(_abc_42016_n2146), .B(_abc_42016_n2147), .Y(_abc_42016_n4021) );
  NOR2X1 NOR2X1_544 ( .A(_abc_42016_n1554), .B(_abc_42016_n1046), .Y(_abc_42016_n4026) );
  NOR2X1 NOR2X1_545 ( .A(_abc_42016_n2083), .B(_abc_42016_n2102_1), .Y(_abc_42016_n4029) );
  NOR2X1 NOR2X1_546 ( .A(regfil_4__7_), .B(_abc_42016_n4000), .Y(_abc_42016_n4035) );
  NOR2X1 NOR2X1_547 ( .A(_abc_42016_n1187), .B(_abc_42016_n4035), .Y(_abc_42016_n4036) );
  NOR2X1 NOR2X1_548 ( .A(_abc_42016_n2031), .B(_abc_42016_n578), .Y(_abc_42016_n4045) );
  NOR2X1 NOR2X1_549 ( .A(_abc_42016_n2231), .B(_abc_42016_n4046), .Y(_abc_42016_n4047) );
  NOR2X1 NOR2X1_55 ( .A(_abc_42016_n664_1), .B(_abc_42016_n601), .Y(_abc_42016_n665_1) );
  NOR2X1 NOR2X1_550 ( .A(_abc_42016_n2094), .B(_abc_42016_n562), .Y(_abc_42016_n4050) );
  NOR2X1 NOR2X1_551 ( .A(regfil_7__5_), .B(regfil_7__6_), .Y(_abc_42016_n4052) );
  NOR2X1 NOR2X1_552 ( .A(reset), .B(_abc_42016_n2217), .Y(_abc_42016_n4054) );
  NOR2X1 NOR2X1_553 ( .A(_abc_42016_n513), .B(_abc_42016_n2033), .Y(_abc_42016_n4057) );
  NOR2X1 NOR2X1_554 ( .A(_abc_42016_n4057), .B(_abc_42016_n4056), .Y(_abc_42016_n4058) );
  NOR2X1 NOR2X1_555 ( .A(_abc_42016_n2087), .B(_abc_42016_n562), .Y(_abc_42016_n4059) );
  NOR2X1 NOR2X1_556 ( .A(_abc_42016_n4049), .B(_abc_42016_n4061), .Y(_abc_42016_n4062) );
  NOR2X1 NOR2X1_557 ( .A(_abc_42016_n2085), .B(_abc_42016_n562), .Y(_abc_42016_n4063) );
  NOR2X1 NOR2X1_558 ( .A(_abc_42016_n669), .B(_abc_42016_n4064), .Y(_abc_42016_n4065) );
  NOR2X1 NOR2X1_559 ( .A(_abc_42016_n2070), .B(_abc_42016_n558), .Y(_abc_42016_n4067) );
  NOR2X1 NOR2X1_56 ( .A(_abc_42016_n520), .B(_abc_42016_n576_1), .Y(_abc_42016_n666) );
  NOR2X1 NOR2X1_560 ( .A(_abc_42016_n4069), .B(_abc_42016_n4065), .Y(_abc_42016_n4070) );
  NOR2X1 NOR2X1_561 ( .A(_abc_42016_n1376), .B(_abc_42016_n4075), .Y(_abc_42016_n4076) );
  NOR2X1 NOR2X1_562 ( .A(_abc_42016_n2317), .B(_abc_42016_n2347_1), .Y(_abc_42016_n4080) );
  NOR2X1 NOR2X1_563 ( .A(_abc_42016_n1000), .B(_abc_42016_n996), .Y(_abc_42016_n4084) );
  NOR2X1 NOR2X1_564 ( .A(_abc_42016_n4082), .B(_abc_42016_n4085), .Y(_abc_42016_n4086) );
  NOR2X1 NOR2X1_565 ( .A(_abc_42016_n4077), .B(_abc_42016_n4087), .Y(_abc_42016_n4088) );
  NOR2X1 NOR2X1_566 ( .A(_abc_42016_n4092_1), .B(_abc_42016_n4090), .Y(_abc_42016_n4093) );
  NOR2X1 NOR2X1_567 ( .A(pc_0_), .B(_abc_42016_n3497_1), .Y(_abc_42016_n4097) );
  NOR2X1 NOR2X1_568 ( .A(_abc_42016_n4101), .B(_abc_42016_n4102), .Y(_abc_42016_n4103) );
  NOR2X1 NOR2X1_569 ( .A(_abc_42016_n2088), .B(_abc_42016_n4104), .Y(_abc_42016_n4105) );
  NOR2X1 NOR2X1_57 ( .A(opcode_4_), .B(_abc_42016_n530), .Y(_abc_42016_n668) );
  NOR2X1 NOR2X1_570 ( .A(_abc_42016_n1376), .B(_abc_42016_n1373), .Y(_abc_42016_n4107) );
  NOR2X1 NOR2X1_571 ( .A(_abc_42016_n566), .B(_abc_42016_n626), .Y(_abc_42016_n4108) );
  NOR2X1 NOR2X1_572 ( .A(_abc_42016_n4106), .B(_abc_42016_n4110), .Y(_abc_42016_n4111) );
  NOR2X1 NOR2X1_573 ( .A(_abc_42016_n2285), .B(_abc_42016_n4113), .Y(_abc_42016_n4114) );
  NOR2X1 NOR2X1_574 ( .A(_abc_42016_n547), .B(_abc_42016_n4119), .Y(_abc_42016_n4120) );
  NOR2X1 NOR2X1_575 ( .A(_abc_42016_n2572), .B(_abc_42016_n1384), .Y(_abc_42016_n4142) );
  NOR2X1 NOR2X1_576 ( .A(_abc_42016_n2592), .B(_abc_42016_n4158), .Y(_abc_42016_n4159) );
  NOR2X1 NOR2X1_577 ( .A(_abc_42016_n4161), .B(_abc_42016_n4091), .Y(_abc_42016_n4163) );
  NOR2X1 NOR2X1_578 ( .A(_abc_42016_n4164), .B(_abc_42016_n4163), .Y(_abc_42016_n4165) );
  NOR2X1 NOR2X1_579 ( .A(_abc_42016_n2632), .B(_abc_42016_n4158), .Y(_abc_42016_n4172) );
  NOR2X1 NOR2X1_58 ( .A(_abc_42016_n669), .B(_abc_42016_n603), .Y(_abc_42016_n670) );
  NOR2X1 NOR2X1_580 ( .A(_abc_42016_n2653), .B(_abc_42016_n4158), .Y(_abc_42016_n4184) );
  NOR2X1 NOR2X1_581 ( .A(_abc_42016_n4187), .B(_abc_42016_n4091), .Y(_abc_42016_n4189) );
  NOR2X1 NOR2X1_582 ( .A(_abc_42016_n4190), .B(_abc_42016_n4189), .Y(_abc_42016_n4191) );
  NOR2X1 NOR2X1_583 ( .A(_abc_42016_n2676), .B(_abc_42016_n4158), .Y(_abc_42016_n4198) );
  NOR2X1 NOR2X1_584 ( .A(_abc_42016_n1353), .B(_abc_42016_n4130), .Y(_abc_42016_n4223) );
  NOR2X1 NOR2X1_585 ( .A(_abc_42016_n4227), .B(_abc_42016_n4226), .Y(_abc_42016_n4228) );
  NOR2X1 NOR2X1_586 ( .A(_abc_42016_n4239), .B(_abc_42016_n4236), .Y(_abc_42016_n4240) );
  NOR2X1 NOR2X1_587 ( .A(_abc_42016_n4131), .B(_abc_42016_n4240), .Y(_abc_42016_n4241) );
  NOR2X1 NOR2X1_588 ( .A(pc_10_), .B(_abc_42016_n1464), .Y(_abc_42016_n4250) );
  NOR2X1 NOR2X1_589 ( .A(_abc_42016_n1466), .B(_abc_42016_n4250), .Y(_abc_42016_n4251) );
  NOR2X1 NOR2X1_59 ( .A(_abc_42016_n672_1), .B(_abc_42016_n540), .Y(_abc_42016_n673) );
  NOR2X1 NOR2X1_590 ( .A(_abc_42016_n4131), .B(_abc_42016_n4267), .Y(_abc_42016_n4268) );
  NOR2X1 NOR2X1_591 ( .A(_abc_42016_n1527), .B(_abc_42016_n1046), .Y(_abc_42016_n4291) );
  NOR2X1 NOR2X1_592 ( .A(_abc_42016_n1848), .B(_abc_42016_n4300), .Y(_abc_42016_n4306) );
  NOR2X1 NOR2X1_593 ( .A(_abc_42016_n4323), .B(_abc_42016_n2024), .Y(_abc_42016_n4324) );
  NOR2X1 NOR2X1_594 ( .A(reset), .B(_abc_42016_n2338), .Y(_abc_42016_n4325) );
  NOR2X1 NOR2X1_595 ( .A(waitr), .B(_abc_42016_n4333), .Y(_abc_42016_n4334) );
  NOR2X1 NOR2X1_596 ( .A(_abc_42016_n556), .B(_abc_42016_n1814), .Y(_abc_42016_n4340) );
  NOR2X1 NOR2X1_597 ( .A(_abc_42016_n4346), .B(_abc_42016_n4098), .Y(_abc_42016_n4347) );
  NOR2X1 NOR2X1_598 ( .A(regfil_7__0_), .B(_abc_42016_n4350), .Y(_abc_42016_n4351) );
  NOR2X1 NOR2X1_599 ( .A(_abc_42016_n2042), .B(_abc_42016_n583), .Y(_abc_42016_n4362) );
  NOR2X1 NOR2X1_6 ( .A(reset), .B(state_5_), .Y(_abc_42016_n515) );
  NOR2X1 NOR2X1_60 ( .A(_abc_42016_n674), .B(_abc_42016_n548), .Y(_abc_42016_n675) );
  NOR2X1 NOR2X1_600 ( .A(_abc_42016_n4367), .B(_abc_42016_n739), .Y(_abc_42016_n4368) );
  NOR2X1 NOR2X1_601 ( .A(opcode_5_), .B(_abc_42016_n4064), .Y(_abc_42016_n4381) );
  NOR2X1 NOR2X1_602 ( .A(reset), .B(_abc_42016_n2044), .Y(_abc_42016_n4382) );
  NOR2X1 NOR2X1_603 ( .A(_abc_42016_n4393), .B(_abc_42016_n4068), .Y(_abc_42016_n4394) );
  NOR2X1 NOR2X1_604 ( .A(_abc_42016_n4397), .B(_abc_42016_n4396), .Y(_abc_42016_n4398) );
  NOR2X1 NOR2X1_605 ( .A(regfil_7__4_), .B(_abc_42016_n4340), .Y(_abc_42016_n4402) );
  NOR2X1 NOR2X1_606 ( .A(_abc_42016_n4411), .B(_abc_42016_n4409), .Y(_abc_42016_n4412) );
  NOR2X1 NOR2X1_607 ( .A(_abc_42016_n4421), .B(_abc_42016_n4419), .Y(_abc_42016_n4422) );
  NOR2X1 NOR2X1_608 ( .A(_abc_42016_n4367), .B(_abc_42016_n909), .Y(_abc_42016_n4423) );
  NOR2X1 NOR2X1_609 ( .A(regfil_7__6_), .B(_abc_42016_n4340), .Y(_abc_42016_n4426) );
  NOR2X1 NOR2X1_61 ( .A(reset), .B(_abc_42016_n676), .Y(_abc_42016_n677) );
  NOR2X1 NOR2X1_610 ( .A(_abc_42016_n898), .B(_abc_42016_n924), .Y(_abc_42016_n4434) );
  NOR2X1 NOR2X1_611 ( .A(_abc_42016_n4452), .B(_abc_42016_n4070), .Y(_abc_42016_n4453) );
  NOR2X1 NOR2X1_612 ( .A(_abc_42016_n2031), .B(_abc_42016_n2270_1), .Y(_abc_42016_n4459) );
  NOR2X1 NOR2X1_613 ( .A(_auto_iopadmap_cc_313_execute_46278), .B(_abc_42016_n2025), .Y(_abc_42016_n4463_1) );
  NOR2X1 NOR2X1_614 ( .A(_abc_42016_n3028), .B(_abc_42016_n2497), .Y(_abc_42016_n4473) );
  NOR2X1 NOR2X1_615 ( .A(_abc_42016_n3223), .B(_abc_42016_n2497), .Y(_abc_42016_n4515) );
  NOR2X1 NOR2X1_616 ( .A(_auto_iopadmap_cc_313_execute_46257_9_), .B(_abc_42016_n4471), .Y(_abc_42016_n4521) );
  NOR2X1 NOR2X1_617 ( .A(_auto_iopadmap_cc_313_execute_46257_10_), .B(_abc_42016_n4471), .Y(_abc_42016_n4525) );
  NOR2X1 NOR2X1_618 ( .A(_auto_iopadmap_cc_313_execute_46257_11_), .B(_abc_42016_n4471), .Y(_abc_42016_n4529) );
  NOR2X1 NOR2X1_619 ( .A(_auto_iopadmap_cc_313_execute_46257_12_), .B(_abc_42016_n4471), .Y(_abc_42016_n4533) );
  NOR2X1 NOR2X1_62 ( .A(opcode_5_), .B(_abc_42016_n531), .Y(_abc_42016_n679) );
  NOR2X1 NOR2X1_620 ( .A(_abc_42016_n1530), .B(_abc_42016_n2024), .Y(_abc_42016_n4536) );
  NOR2X1 NOR2X1_621 ( .A(_auto_iopadmap_cc_313_execute_46257_14_), .B(_abc_42016_n4471), .Y(_abc_42016_n4542) );
  NOR2X1 NOR2X1_622 ( .A(_auto_iopadmap_cc_313_execute_46257_15_), .B(_abc_42016_n4471), .Y(_abc_42016_n4546) );
  NOR2X1 NOR2X1_623 ( .A(_abc_42016_n4548), .B(_abc_42016_n2437), .Y(_abc_42016_n4549) );
  NOR2X1 NOR2X1_624 ( .A(statesel_4_), .B(_abc_42016_n2446), .Y(_abc_42016_n4551) );
  NOR2X1 NOR2X1_625 ( .A(_abc_42016_n2417_1), .B(_abc_42016_n2446), .Y(_abc_42016_n4557) );
  NOR2X1 NOR2X1_626 ( .A(_abc_42016_n4558), .B(_abc_42016_n4556), .Y(_abc_42016_n4559) );
  NOR2X1 NOR2X1_627 ( .A(_abc_42016_n1909_1), .B(_abc_42016_n548), .Y(_abc_42016_n4561) );
  NOR2X1 NOR2X1_628 ( .A(statesel_2_), .B(statesel_3_), .Y(_abc_42016_n4565) );
  NOR2X1 NOR2X1_629 ( .A(_abc_42016_n4566), .B(_abc_42016_n4564), .Y(_abc_42016_n4567) );
  NOR2X1 NOR2X1_63 ( .A(_abc_42016_n680), .B(_abc_42016_n603), .Y(_abc_42016_n681) );
  NOR2X1 NOR2X1_630 ( .A(statesel_2_), .B(_abc_42016_n2394_1), .Y(_abc_42016_n4568) );
  NOR2X1 NOR2X1_631 ( .A(_abc_42016_n4569), .B(_abc_42016_n2407), .Y(_abc_42016_n4570_1) );
  NOR2X1 NOR2X1_632 ( .A(_abc_42016_n2451), .B(_abc_42016_n4556), .Y(_abc_42016_n4571) );
  NOR2X1 NOR2X1_633 ( .A(_abc_42016_n4573), .B(_abc_42016_n4563), .Y(_abc_42016_n4574) );
  NOR2X1 NOR2X1_634 ( .A(_abc_42016_n4554_1), .B(_abc_42016_n4575), .Y(_abc_42016_n4576) );
  NOR2X1 NOR2X1_635 ( .A(statesel_4_), .B(statesel_5_), .Y(_abc_42016_n4578) );
  NOR2X1 NOR2X1_636 ( .A(statesel_0_), .B(statesel_1_), .Y(_abc_42016_n4580) );
  NOR2X1 NOR2X1_637 ( .A(_abc_42016_n4581), .B(_abc_42016_n4569), .Y(_abc_42016_n4582) );
  NOR2X1 NOR2X1_638 ( .A(_abc_42016_n4581), .B(_abc_42016_n2437), .Y(_abc_42016_n4587) );
  NOR2X1 NOR2X1_639 ( .A(_abc_42016_n4583), .B(_abc_42016_n4552), .Y(_abc_42016_n4589) );
  NOR2X1 NOR2X1_64 ( .A(_abc_42016_n680), .B(_abc_42016_n682), .Y(_abc_42016_n683) );
  NOR2X1 NOR2X1_640 ( .A(_abc_42016_n4591), .B(_abc_42016_n4586), .Y(_abc_42016_n4592) );
  NOR2X1 NOR2X1_641 ( .A(_abc_42016_n4566), .B(_abc_42016_n2407), .Y(_abc_42016_n4595) );
  NOR2X1 NOR2X1_642 ( .A(_abc_42016_n4548), .B(_abc_42016_n2409), .Y(_abc_42016_n4601) );
  NOR2X1 NOR2X1_643 ( .A(_abc_42016_n4602), .B(_abc_42016_n4560), .Y(_abc_42016_n4603) );
  NOR2X1 NOR2X1_644 ( .A(_abc_42016_n4607), .B(_abc_42016_n4603), .Y(_abc_42016_n4608) );
  NOR2X1 NOR2X1_645 ( .A(_abc_42016_n4588), .B(_abc_42016_n4593), .Y(_abc_42016_n4612) );
  NOR2X1 NOR2X1_646 ( .A(_abc_42016_n4620), .B(_abc_42016_n4612), .Y(_abc_42016_n4621) );
  NOR2X1 NOR2X1_647 ( .A(_abc_42016_n4548), .B(_abc_42016_n4569), .Y(_abc_42016_n4626) );
  NOR2X1 NOR2X1_648 ( .A(_abc_42016_n4596), .B(_abc_42016_n4552), .Y(_abc_42016_n4630) );
  NOR2X1 NOR2X1_649 ( .A(_abc_42016_n4632_1), .B(_abc_42016_n562), .Y(_abc_42016_n4633) );
  NOR2X1 NOR2X1_65 ( .A(popdes_1_), .B(_abc_42016_n686), .Y(_abc_42016_n687) );
  NOR2X1 NOR2X1_650 ( .A(_abc_42016_n4636), .B(_abc_42016_n4629), .Y(_abc_42016_n4637) );
  NOR2X1 NOR2X1_651 ( .A(_abc_42016_n2347_1), .B(_abc_42016_n1001_1), .Y(_abc_42016_n4650_1) );
  NOR2X1 NOR2X1_652 ( .A(_abc_42016_n4649), .B(_abc_42016_n4651), .Y(_abc_42016_n4652) );
  NOR2X1 NOR2X1_653 ( .A(_abc_42016_n4565), .B(_abc_42016_n2436), .Y(_abc_42016_n4655) );
  NOR2X1 NOR2X1_654 ( .A(_abc_42016_n4564), .B(_abc_42016_n4655), .Y(_abc_42016_n4656) );
  NOR2X1 NOR2X1_655 ( .A(_abc_42016_n4581), .B(_abc_42016_n4558), .Y(_abc_42016_n4664) );
  NOR2X1 NOR2X1_656 ( .A(reset), .B(_abc_42016_n2280), .Y(_abc_42016_n4669) );
  NOR2X1 NOR2X1_657 ( .A(_abc_42016_n2344), .B(_abc_42016_n4569), .Y(_abc_42016_n4677) );
  NOR2X1 NOR2X1_658 ( .A(reset), .B(_abc_42016_n1923), .Y(_abc_42016_n4688_1) );
  NOR2X1 NOR2X1_659 ( .A(_abc_42016_n4692), .B(_abc_42016_n4690), .Y(_abc_42016_n4693) );
  NOR2X1 NOR2X1_66 ( .A(_abc_42016_n689), .B(_abc_42016_n685), .Y(_abc_42016_n690) );
  NOR2X1 NOR2X1_660 ( .A(_abc_42016_n4696), .B(_abc_42016_n4697), .Y(_abc_42016_n4698_1) );
  NOR2X1 NOR2X1_661 ( .A(_abc_42016_n2231), .B(_abc_42016_n4333), .Y(_abc_42016_n4702) );
  NOR2X1 NOR2X1_662 ( .A(_abc_42016_n4702), .B(_abc_42016_n4605), .Y(_abc_42016_n4703) );
  NOR2X1 NOR2X1_663 ( .A(_abc_42016_n4704), .B(_abc_42016_n4701), .Y(_abc_42016_n4705_1) );
  NOR2X1 NOR2X1_664 ( .A(_abc_42016_n4696), .B(_abc_42016_n4575), .Y(_abc_42016_n4706) );
  NOR2X1 NOR2X1_665 ( .A(_abc_42016_n4702), .B(_abc_42016_n4554_1), .Y(_abc_42016_n4709) );
  NOR2X1 NOR2X1_666 ( .A(_abc_42016_n4710), .B(_abc_42016_n4708), .Y(_abc_42016_n4711_1) );
  NOR2X1 NOR2X1_667 ( .A(_abc_42016_n4713_1), .B(_abc_42016_n4573), .Y(_abc_42016_n4714) );
  NOR2X1 NOR2X1_668 ( .A(_abc_42016_n4612), .B(_abc_42016_n4603), .Y(_abc_42016_n4715) );
  NOR2X1 NOR2X1_669 ( .A(_abc_42016_n4586), .B(_abc_42016_n4716), .Y(_abc_42016_n4717_1) );
  NOR2X1 NOR2X1_67 ( .A(_abc_42016_n671_1), .B(_abc_42016_n678), .Y(_abc_42016_n696) );
  NOR2X1 NOR2X1_670 ( .A(_abc_42016_n4719_1), .B(_abc_42016_n4721), .Y(_abc_42016_n4722) );
  NOR2X1 NOR2X1_671 ( .A(_abc_42016_n4724), .B(_abc_42016_n4723_1), .Y(_abc_42016_n4725_1) );
  NOR2X1 NOR2X1_672 ( .A(_abc_42016_n4589), .B(_abc_42016_n4727), .Y(_abc_42016_n4728) );
  NOR2X1 NOR2X1_673 ( .A(alu_oprb_1_), .B(alu_opra_1_), .Y(alu__abc_41682_n34) );
  NOR2X1 NOR2X1_674 ( .A(alu__abc_41682_n34), .B(alu__abc_41682_n35), .Y(alu__abc_41682_n36) );
  NOR2X1 NOR2X1_675 ( .A(alu_oprb_0_), .B(alu_opra_0_), .Y(alu__abc_41682_n38) );
  NOR2X1 NOR2X1_676 ( .A(alu__abc_41682_n38), .B(alu__abc_41682_n37), .Y(alu__abc_41682_n39) );
  NOR2X1 NOR2X1_677 ( .A(alu__abc_41682_n44), .B(alu__abc_41682_n41), .Y(alu__abc_41682_n46_1) );
  NOR2X1 NOR2X1_678 ( .A(alu__abc_41682_n52), .B(alu__abc_41682_n55), .Y(alu__abc_41682_n56) );
  NOR2X1 NOR2X1_679 ( .A(alu_oprb_4_), .B(alu_opra_4_), .Y(alu__abc_41682_n59) );
  NOR2X1 NOR2X1_68 ( .A(regfil_3__0_), .B(regfil_3__1_), .Y(_abc_42016_n702_1) );
  NOR2X1 NOR2X1_680 ( .A(alu__abc_41682_n59), .B(alu__abc_41682_n61), .Y(alu__abc_41682_n62) );
  NOR2X1 NOR2X1_681 ( .A(alu_oprb_3_), .B(alu_opra_3_), .Y(alu__abc_41682_n63) );
  NOR2X1 NOR2X1_682 ( .A(alu__abc_41682_n62), .B(alu__abc_41682_n70), .Y(alu__abc_41682_n71) );
  NOR2X1 NOR2X1_683 ( .A(alu_oprb_5_), .B(alu_opra_5_), .Y(alu__abc_41682_n73) );
  NOR2X1 NOR2X1_684 ( .A(alu_oprb_6_), .B(alu_opra_6_), .Y(alu__abc_41682_n84) );
  NOR2X1 NOR2X1_685 ( .A(alu__abc_41682_n85), .B(alu__abc_41682_n86), .Y(alu__abc_41682_n87) );
  NOR2X1 NOR2X1_686 ( .A(alu__abc_41682_n84), .B(alu__abc_41682_n87), .Y(alu__abc_41682_n88) );
  NOR2X1 NOR2X1_687 ( .A(alu__abc_41682_n81), .B(alu__abc_41682_n92), .Y(alu__abc_41682_n93) );
  NOR2X1 NOR2X1_688 ( .A(alu_oprb_7_), .B(alu_opra_7_), .Y(alu__abc_41682_n95) );
  NOR2X1 NOR2X1_689 ( .A(alu__abc_41682_n96), .B(alu__abc_41682_n97), .Y(alu__abc_41682_n98) );
  NOR2X1 NOR2X1_69 ( .A(_abc_42016_n634), .B(_abc_42016_n703), .Y(_abc_42016_n704) );
  NOR2X1 NOR2X1_690 ( .A(alu__abc_41682_n95), .B(alu__abc_41682_n98), .Y(alu__abc_41682_n99) );
  NOR2X1 NOR2X1_691 ( .A(alu_sel_2_), .B(alu__abc_41682_n104), .Y(alu__abc_41682_n105) );
  NOR2X1 NOR2X1_692 ( .A(alu_sel_1_), .B(alu__abc_41682_n106), .Y(alu__abc_41682_n107) );
  NOR2X1 NOR2X1_693 ( .A(alu_oprb_5_), .B(alu__abc_41682_n115), .Y(alu__abc_41682_n116) );
  NOR2X1 NOR2X1_694 ( .A(alu_oprb_4_), .B(alu__abc_41682_n118), .Y(alu__abc_41682_n119) );
  NOR2X1 NOR2X1_695 ( .A(alu_oprb_2_), .B(alu__abc_41682_n121), .Y(alu__abc_41682_n122) );
  NOR2X1 NOR2X1_696 ( .A(alu_oprb_6_), .B(alu__abc_41682_n86), .Y(alu__abc_41682_n132) );
  NOR2X1 NOR2X1_697 ( .A(alu_oprb_1_), .B(alu__abc_41682_n123), .Y(alu__abc_41682_n138) );
  NOR2X1 NOR2X1_698 ( .A(alu__abc_41682_n149), .B(alu__abc_41682_n106), .Y(alu__abc_41682_n150) );
  NOR2X1 NOR2X1_699 ( .A(alu__abc_41682_n104), .B(alu__abc_41682_n153), .Y(alu__abc_41682_n178) );
  NOR2X1 NOR2X1_7 ( .A(_abc_42016_n514), .B(_abc_42016_n516), .Y(_abc_42016_n517) );
  NOR2X1 NOR2X1_70 ( .A(_abc_42016_n702_1), .B(_abc_42016_n704), .Y(_abc_42016_n706) );
  NOR2X1 NOR2X1_700 ( .A(alu_sel_0_), .B(alu__abc_41682_n153), .Y(alu__abc_41682_n180) );
  NOR2X1 NOR2X1_701 ( .A(alu_sel_1_), .B(alu_sel_0_), .Y(alu__abc_41682_n184) );
  NOR2X1 NOR2X1_702 ( .A(alu__abc_41682_n194), .B(alu__abc_41682_n219), .Y(alu__abc_41682_n220) );
  NOR2X1 NOR2X1_703 ( .A(alu__abc_41682_n209), .B(alu__abc_41682_n215), .Y(alu__abc_41682_n230) );
  NOR2X1 NOR2X1_704 ( .A(alu__abc_41682_n255), .B(alu__abc_41682_n217), .Y(alu__abc_41682_n256) );
  NOR2X1 NOR2X1_705 ( .A(alu__abc_41682_n56), .B(alu__abc_41682_n57), .Y(alu__abc_41682_n261) );
  NOR2X1 NOR2X1_706 ( .A(alu__abc_41682_n193), .B(alu__abc_41682_n273_1), .Y(alu__abc_41682_n274) );
  NOR2X1 NOR2X1_707 ( .A(alu__abc_41682_n198), .B(alu__abc_41682_n47), .Y(alu__abc_41682_n275_1) );
  NOR2X1 NOR2X1_708 ( .A(alu__abc_41682_n127), .B(alu__abc_41682_n205), .Y(alu__abc_41682_n279_1) );
  NOR2X1 NOR2X1_709 ( .A(alu__abc_41682_n53), .B(alu__abc_41682_n218), .Y(alu__abc_41682_n280_1) );
  NOR2X1 NOR2X1_71 ( .A(regfil_0__1_), .B(_abc_42016_n619), .Y(_abc_42016_n715) );
  NOR2X1 NOR2X1_710 ( .A(alu__abc_41682_n141), .B(alu__abc_41682_n164), .Y(alu__abc_41682_n283) );
  NOR2X1 NOR2X1_711 ( .A(alu__abc_41682_n295), .B(alu__abc_41682_n297), .Y(alu__abc_41682_n298) );
  NOR2X1 NOR2X1_712 ( .A(alu__abc_41682_n268_1), .B(alu__abc_41682_n271_1), .Y(alu__abc_41682_n314_1) );
  NOR2X1 NOR2X1_713 ( .A(alu__abc_41682_n336), .B(alu__abc_41682_n322), .Y(alu__abc_41682_n337) );
  NOR2X1 NOR2X1_72 ( .A(_abc_42016_n714), .B(_abc_42016_n737), .Y(_abc_42016_n738) );
  NOR2X1 NOR2X1_73 ( .A(_abc_42016_n601), .B(_abc_42016_n739), .Y(_abc_42016_n740) );
  NOR2X1 NOR2X1_74 ( .A(_abc_42016_n601), .B(_abc_42016_n769), .Y(_abc_42016_n770) );
  NOR2X1 NOR2X1_75 ( .A(_abc_42016_n776), .B(_abc_42016_n772), .Y(_abc_42016_n777) );
  NOR2X1 NOR2X1_76 ( .A(regfil_3__2_), .B(_abc_42016_n782), .Y(_abc_42016_n783) );
  NOR2X1 NOR2X1_77 ( .A(regfil_0__3_), .B(_abc_42016_n748), .Y(_abc_42016_n789) );
  NOR2X1 NOR2X1_78 ( .A(_abc_42016_n743), .B(_abc_42016_n744), .Y(_abc_42016_n814) );
  NOR2X1 NOR2X1_79 ( .A(_abc_42016_n810_1), .B(_abc_42016_n817), .Y(_abc_42016_n818) );
  NOR2X1 NOR2X1_8 ( .A(state_1_), .B(_abc_42016_n505), .Y(_abc_42016_n519) );
  NOR2X1 NOR2X1_80 ( .A(_abc_42016_n795), .B(_abc_42016_n775), .Y(_abc_42016_n824) );
  NOR2X1 NOR2X1_81 ( .A(_abc_42016_n601), .B(_abc_42016_n858), .Y(_abc_42016_n859) );
  NOR2X1 NOR2X1_82 ( .A(regfil_3__4_), .B(_abc_42016_n828), .Y(_abc_42016_n866) );
  NOR2X1 NOR2X1_83 ( .A(_abc_42016_n872), .B(_abc_42016_n697), .Y(_abc_42016_n873) );
  NOR2X1 NOR2X1_84 ( .A(_abc_42016_n874), .B(_abc_42016_n866), .Y(_abc_42016_n876) );
  NOR2X1 NOR2X1_85 ( .A(_abc_42016_n834), .B(_abc_42016_n815), .Y(_abc_42016_n883) );
  NOR2X1 NOR2X1_86 ( .A(regfil_0__5_), .B(_abc_42016_n883), .Y(_abc_42016_n884) );
  NOR2X1 NOR2X1_87 ( .A(regfil_0__5_), .B(_abc_42016_n838), .Y(_abc_42016_n887) );
  NOR2X1 NOR2X1_88 ( .A(regfil_6__5_), .B(_abc_42016_n539), .Y(_abc_42016_n892) );
  NOR2X1 NOR2X1_89 ( .A(_abc_42016_n601), .B(_abc_42016_n909), .Y(_abc_42016_n910_1) );
  NOR2X1 NOR2X1_9 ( .A(_abc_42016_n501), .B(_abc_42016_n521), .Y(_abc_42016_n522) );
  NOR2X1 NOR2X1_90 ( .A(_abc_42016_n601), .B(_abc_42016_n934), .Y(_abc_42016_n935) );
  NOR2X1 NOR2X1_91 ( .A(_abc_42016_n874), .B(_abc_42016_n863), .Y(_abc_42016_n937) );
  NOR2X1 NOR2X1_92 ( .A(_abc_42016_n939), .B(_abc_42016_n878), .Y(_abc_42016_n942) );
  NOR2X1 NOR2X1_93 ( .A(regfil_3__6_), .B(_abc_42016_n877), .Y(_abc_42016_n943) );
  NOR2X1 NOR2X1_94 ( .A(_abc_42016_n913), .B(_abc_42016_n885), .Y(_abc_42016_n952) );
  NOR2X1 NOR2X1_95 ( .A(_abc_42016_n601), .B(_abc_42016_n971), .Y(_abc_42016_n972) );
  NOR2X1 NOR2X1_96 ( .A(_abc_42016_n974), .B(_abc_42016_n943), .Y(_abc_42016_n975) );
  NOR2X1 NOR2X1_97 ( .A(_abc_42016_n974), .B(_abc_42016_n938), .Y(_abc_42016_n980) );
  NOR2X1 NOR2X1_98 ( .A(_abc_42016_n980), .B(_abc_42016_n772), .Y(_abc_42016_n981) );
  NOR2X1 NOR2X1_99 ( .A(_abc_42016_n556), .B(_abc_42016_n988), .Y(_abc_42016_n989) );
  NOR3X1 NOR3X1_1 ( .A(alu__abc_41682_n40), .B(alu__abc_41682_n46_1), .C(alu__abc_41682_n45_1), .Y(alu__abc_41682_n47) );
  NOR3X1 NOR3X1_2 ( .A(alu__abc_41682_n71), .B(alu__abc_41682_n69), .C(alu__abc_41682_n58), .Y(alu__abc_41682_n72) );
  NOR3X1 NOR3X1_3 ( .A(alu__abc_41682_n34), .B(alu__abc_41682_n35), .C(alu__abc_41682_n163), .Y(alu__abc_41682_n164) );
  NOR3X1 NOR3X1_4 ( .A(alu__abc_41682_n138), .B(alu__abc_41682_n137), .C(alu__abc_41682_n141), .Y(alu__abc_41682_n205) );
  NOR3X1 NOR3X1_5 ( .A(alu__abc_41682_n271_1), .B(alu__abc_41682_n268_1), .C(alu__abc_41682_n287), .Y(alu__abc_41682_n290) );
  OAI21X1 OAI21X1_1 ( .A(_abc_42016_n509), .B(_abc_42016_n513), .C(_abc_42016_n527), .Y(_abc_42016_n528_1) );
  OAI21X1 OAI21X1_10 ( .A(_abc_42016_n552), .B(_abc_42016_n526_1), .C(_abc_42016_n594_1), .Y(_abc_42016_n595) );
  OAI21X1 OAI21X1_100 ( .A(_abc_42016_n973), .B(_abc_42016_n972), .C(_abc_42016_n985), .Y(_abc_36783_n3382) );
  OAI21X1 OAI21X1_1000 ( .A(_abc_42016_n3807), .B(_abc_42016_n3808), .C(_abc_42016_n3805), .Y(_abc_42016_n3809) );
  OAI21X1 OAI21X1_1001 ( .A(_abc_42016_n959), .B(_abc_42016_n1290), .C(_abc_42016_n629), .Y(_abc_42016_n3811) );
  OAI21X1 OAI21X1_1002 ( .A(_abc_42016_n1325), .B(_abc_42016_n3814), .C(_abc_42016_n3813), .Y(_abc_42016_n3815) );
  OAI21X1 OAI21X1_1003 ( .A(_abc_42016_n1306), .B(_abc_42016_n3819), .C(_abc_42016_n3818), .Y(_abc_42016_n3820) );
  OAI21X1 OAI21X1_1004 ( .A(_abc_42016_n1317), .B(_abc_42016_n1315), .C(_abc_42016_n2168), .Y(_abc_42016_n3822) );
  OAI21X1 OAI21X1_1005 ( .A(_abc_42016_n2167), .B(_abc_42016_n3822), .C(_abc_42016_n1031_1), .Y(_abc_42016_n3823) );
  OAI21X1 OAI21X1_1006 ( .A(_abc_42016_n1045), .B(_abc_42016_n3816), .C(_abc_42016_n3825), .Y(_abc_42016_n3826) );
  OAI21X1 OAI21X1_1007 ( .A(_abc_42016_n3802), .B(_abc_42016_n3828), .C(_abc_42016_n3829), .Y(_abc_42016_n3830) );
  OAI21X1 OAI21X1_1008 ( .A(_abc_42016_n714), .B(_abc_42016_n737), .C(_abc_42016_n3800), .Y(_abc_42016_n3833) );
  OAI21X1 OAI21X1_1009 ( .A(_abc_42016_n728), .B(_abc_42016_n697), .C(_abc_42016_n994), .Y(_abc_42016_n3836) );
  OAI21X1 OAI21X1_101 ( .A(_abc_42016_n671_1), .B(_abc_42016_n678), .C(_abc_42016_n994), .Y(_abc_42016_n995) );
  OAI21X1 OAI21X1_1010 ( .A(_abc_42016_n3837), .B(_abc_42016_n3838), .C(_abc_42016_n1170), .Y(_abc_42016_n3839_1) );
  OAI21X1 OAI21X1_1011 ( .A(_abc_42016_n1125), .B(_abc_42016_n1138), .C(_abc_42016_n3839_1), .Y(_abc_42016_n3840) );
  OAI21X1 OAI21X1_1012 ( .A(_abc_42016_n629), .B(_abc_42016_n2131_1), .C(_abc_42016_n2136_1), .Y(_abc_42016_n3841) );
  OAI21X1 OAI21X1_1013 ( .A(_abc_42016_n2128_1), .B(_abc_42016_n2125), .C(_abc_42016_n3841), .Y(_abc_42016_n3844) );
  OAI21X1 OAI21X1_1014 ( .A(_abc_42016_n608), .B(_abc_42016_n629), .C(_abc_42016_n2203), .Y(_abc_42016_n3846) );
  OAI21X1 OAI21X1_1015 ( .A(_abc_42016_n3849), .B(_abc_42016_n3850), .C(_abc_42016_n3851), .Y(_abc_42016_n3852) );
  OAI21X1 OAI21X1_1016 ( .A(_abc_42016_n1151), .B(_abc_42016_n3848), .C(_abc_42016_n3852), .Y(_abc_42016_n3853) );
  OAI21X1 OAI21X1_1017 ( .A(_abc_42016_n629), .B(_abc_42016_n1048), .C(_abc_42016_n1045), .Y(_abc_42016_n3854) );
  OAI21X1 OAI21X1_1018 ( .A(_abc_42016_n3854), .B(_abc_42016_n3853), .C(_abc_42016_n3845), .Y(_abc_42016_n3855) );
  OAI21X1 OAI21X1_1019 ( .A(_abc_42016_n722), .B(_abc_42016_n3807), .C(_abc_42016_n1125), .Y(_abc_42016_n3857) );
  OAI21X1 OAI21X1_102 ( .A(_abc_42016_n670), .B(_abc_42016_n996), .C(_abc_42016_n561), .Y(_abc_42016_n997) );
  OAI21X1 OAI21X1_1020 ( .A(_abc_42016_n3856), .B(_abc_42016_n3857), .C(_abc_42016_n3805), .Y(_abc_42016_n3858) );
  OAI21X1 OAI21X1_1021 ( .A(_abc_42016_n719), .B(_abc_42016_n1056), .C(_abc_42016_n3860), .Y(_abc_42016_n3861) );
  OAI21X1 OAI21X1_1022 ( .A(rdatahold_1_), .B(_abc_42016_n1097), .C(_abc_42016_n3861), .Y(_abc_42016_n3862) );
  OAI21X1 OAI21X1_1023 ( .A(_abc_42016_n769), .B(_abc_42016_n3834), .C(_abc_42016_n3864), .Y(_abc_42016_n3865) );
  OAI21X1 OAI21X1_1024 ( .A(_abc_42016_n1446), .B(_abc_42016_n3856), .C(_abc_42016_n1125), .Y(_abc_42016_n3869) );
  OAI21X1 OAI21X1_1025 ( .A(_abc_42016_n3869), .B(_abc_42016_n3868), .C(_abc_42016_n3805), .Y(_abc_42016_n3870) );
  OAI21X1 OAI21X1_1026 ( .A(_abc_42016_n722), .B(_abc_42016_n3810), .C(_abc_42016_n1446), .Y(_abc_42016_n3871) );
  OAI21X1 OAI21X1_1027 ( .A(_abc_42016_n2125), .B(_abc_42016_n3875), .C(_abc_42016_n3874), .Y(_abc_42016_n3876) );
  OAI21X1 OAI21X1_1028 ( .A(regfil_2__1_), .B(regfil_4__1_), .C(_abc_42016_n2171), .Y(_abc_42016_n3882) );
  OAI21X1 OAI21X1_1029 ( .A(_abc_42016_n722), .B(_abc_42016_n1048), .C(_abc_42016_n3885), .Y(_abc_42016_n3886) );
  OAI21X1 OAI21X1_103 ( .A(_abc_42016_n1000), .B(_abc_42016_n1001_1), .C(_abc_42016_n561), .Y(_abc_42016_n1002) );
  OAI21X1 OAI21X1_1030 ( .A(_abc_42016_n1187), .B(_abc_42016_n3873), .C(_abc_42016_n3887), .Y(_abc_42016_n3888) );
  OAI21X1 OAI21X1_1031 ( .A(_abc_42016_n3870), .B(_abc_42016_n3889), .C(_abc_42016_n3892), .Y(_abc_42016_n3893) );
  OAI21X1 OAI21X1_1032 ( .A(_abc_42016_n3866), .B(_abc_42016_n3894), .C(_abc_42016_n3865), .Y(_abc_36783_n4533) );
  OAI21X1 OAI21X1_1033 ( .A(_abc_42016_n3834), .B(_abc_42016_n819), .C(_abc_42016_n1020), .Y(_abc_42016_n3897) );
  OAI21X1 OAI21X1_1034 ( .A(_abc_42016_n800), .B(_abc_42016_n3868), .C(_abc_42016_n3899), .Y(_abc_42016_n3900) );
  OAI21X1 OAI21X1_1035 ( .A(_abc_42016_n743), .B(_abc_42016_n1446), .C(_abc_42016_n2205), .Y(_abc_42016_n3901) );
  OAI21X1 OAI21X1_1036 ( .A(_abc_42016_n3902), .B(_abc_42016_n3903), .C(_abc_42016_n3904), .Y(_abc_42016_n3905) );
  OAI21X1 OAI21X1_1037 ( .A(_abc_42016_n3908), .B(_abc_42016_n3907), .C(_abc_42016_n1170), .Y(_abc_42016_n3909) );
  OAI21X1 OAI21X1_1038 ( .A(_abc_42016_n753), .B(_abc_42016_n1446), .C(_abc_42016_n2172_1), .Y(_abc_42016_n3910) );
  OAI21X1 OAI21X1_1039 ( .A(_abc_42016_n2155), .B(_abc_42016_n2157), .C(_abc_42016_n3912), .Y(_abc_42016_n3913) );
  OAI21X1 OAI21X1_104 ( .A(_abc_42016_n1005), .B(_abc_42016_n1006), .C(_abc_42016_n561), .Y(_abc_42016_n1007) );
  OAI21X1 OAI21X1_1040 ( .A(_abc_42016_n1446), .B(_abc_42016_n2122), .C(_abc_42016_n2138), .Y(_abc_42016_n3915) );
  OAI21X1 OAI21X1_1041 ( .A(_abc_42016_n1045), .B(_abc_42016_n3917), .C(_abc_42016_n3914), .Y(_abc_42016_n3918) );
  OAI21X1 OAI21X1_1042 ( .A(_abc_42016_n796), .B(_abc_42016_n697), .C(_abc_42016_n994), .Y(_abc_42016_n3921) );
  OAI21X1 OAI21X1_1043 ( .A(_abc_42016_n811), .B(_abc_42016_n1056), .C(_abc_42016_n3922), .Y(_abc_42016_n3923) );
  OAI21X1 OAI21X1_1044 ( .A(rdatahold_3_), .B(_abc_42016_n994), .C(_abc_42016_n3923), .Y(_abc_42016_n3924) );
  OAI21X1 OAI21X1_1045 ( .A(_abc_42016_n3896), .B(_abc_42016_n3897), .C(_abc_42016_n3924), .Y(_abc_36783_n4534) );
  OAI21X1 OAI21X1_1046 ( .A(_abc_42016_n3834), .B(_abc_42016_n858), .C(_abc_42016_n3926), .Y(_abc_42016_n3927) );
  OAI21X1 OAI21X1_1047 ( .A(_abc_42016_n2116_1), .B(_abc_42016_n3930), .C(_abc_42016_n3929), .Y(_abc_42016_n3931) );
  OAI21X1 OAI21X1_1048 ( .A(regfil_4__4_), .B(_abc_42016_n3907), .C(_abc_42016_n1138), .Y(_abc_42016_n3934) );
  OAI21X1 OAI21X1_1049 ( .A(_abc_42016_n670), .B(_abc_42016_n3935_1), .C(_abc_42016_n561), .Y(_abc_42016_n3936) );
  OAI21X1 OAI21X1_105 ( .A(reset), .B(_abc_42016_n1014), .C(_abc_42016_n1018), .Y(_abc_42016_n1019) );
  OAI21X1 OAI21X1_1050 ( .A(_abc_42016_n3933), .B(_abc_42016_n3934), .C(_abc_42016_n3936), .Y(_abc_42016_n3937) );
  OAI21X1 OAI21X1_1051 ( .A(_abc_42016_n2187), .B(_abc_42016_n3939), .C(_abc_42016_n3940), .Y(_abc_42016_n3941) );
  OAI21X1 OAI21X1_1052 ( .A(_abc_42016_n2154), .B(_abc_42016_n3942), .C(_abc_42016_n3943), .Y(_abc_42016_n3944) );
  OAI21X1 OAI21X1_1053 ( .A(regfil_4__3_), .B(_abc_42016_n3867), .C(regfil_4__4_), .Y(_abc_42016_n3946) );
  OAI21X1 OAI21X1_1054 ( .A(_abc_42016_n847), .B(_abc_42016_n697), .C(_abc_42016_n3951), .Y(_abc_42016_n3952) );
  OAI21X1 OAI21X1_1055 ( .A(_abc_42016_n3928), .B(_abc_42016_n3953), .C(_abc_42016_n3927), .Y(_abc_36783_n4535) );
  OAI21X1 OAI21X1_1056 ( .A(_abc_42016_n895), .B(_abc_42016_n697), .C(_abc_42016_n994), .Y(_abc_42016_n3957) );
  OAI21X1 OAI21X1_1057 ( .A(_abc_42016_n1527), .B(_abc_42016_n3948), .C(_abc_42016_n1125), .Y(_abc_42016_n3959) );
  OAI21X1 OAI21X1_1058 ( .A(_abc_42016_n3958), .B(_abc_42016_n3959), .C(_abc_42016_n3805), .Y(_abc_42016_n3960) );
  OAI21X1 OAI21X1_1059 ( .A(_abc_42016_n847), .B(_abc_42016_n842), .C(_abc_42016_n2174), .Y(_abc_42016_n3961) );
  OAI21X1 OAI21X1_106 ( .A(regfil_5__0_), .B(_abc_42016_n989), .C(_abc_42016_n1020), .Y(_abc_42016_n1021) );
  OAI21X1 OAI21X1_1060 ( .A(_abc_42016_n3965), .B(_abc_42016_n3966), .C(_abc_42016_n3967), .Y(_abc_42016_n3968) );
  OAI21X1 OAI21X1_1061 ( .A(_abc_42016_n842), .B(_abc_42016_n2113), .C(_abc_42016_n2140_1), .Y(_abc_42016_n3971) );
  OAI21X1 OAI21X1_1062 ( .A(_abc_42016_n1023), .B(_abc_42016_n3970), .C(_abc_42016_n3974), .Y(_abc_42016_n3975) );
  OAI21X1 OAI21X1_1063 ( .A(_abc_42016_n3957), .B(_abc_42016_n3980), .C(_abc_42016_n3981), .Y(_abc_42016_n3982) );
  OAI21X1 OAI21X1_1064 ( .A(_abc_42016_n3834), .B(_abc_42016_n934), .C(_abc_42016_n3985), .Y(_abc_42016_n3986) );
  OAI21X1 OAI21X1_1065 ( .A(regfil_4__5_), .B(_abc_42016_n3947), .C(regfil_4__6_), .Y(_abc_42016_n3988) );
  OAI21X1 OAI21X1_1066 ( .A(regfil_0__5_), .B(regfil_4__5_), .C(_abc_42016_n2208), .Y(_abc_42016_n3991) );
  OAI21X1 OAI21X1_1067 ( .A(_abc_42016_n4001), .B(_abc_42016_n4000), .C(_abc_42016_n1170), .Y(_abc_42016_n4002) );
  OAI21X1 OAI21X1_1068 ( .A(_abc_42016_n3999), .B(_abc_42016_n3998), .C(_abc_42016_n4003), .Y(_abc_42016_n4004) );
  OAI21X1 OAI21X1_1069 ( .A(_abc_42016_n919), .B(_abc_42016_n697), .C(_abc_42016_n994), .Y(_abc_42016_n4007) );
  OAI21X1 OAI21X1_107 ( .A(_abc_42016_n1025), .B(_abc_42016_n1026), .C(_abc_42016_n1023), .Y(_abc_42016_n1027) );
  OAI21X1 OAI21X1_1070 ( .A(_abc_42016_n4007), .B(_abc_42016_n4006), .C(_abc_42016_n4008), .Y(_abc_42016_n4009) );
  OAI21X1 OAI21X1_1071 ( .A(_abc_42016_n3834), .B(_abc_42016_n971), .C(_abc_42016_n4011), .Y(_abc_42016_n4012) );
  OAI21X1 OAI21X1_1072 ( .A(_abc_42016_n2478), .B(_abc_42016_n1018), .C(_abc_42016_n4013), .Y(_abc_42016_n4014) );
  OAI21X1 OAI21X1_1073 ( .A(regfil_2__7_), .B(_abc_42016_n993), .C(_abc_42016_n995), .Y(_abc_42016_n4015) );
  OAI21X1 OAI21X1_1074 ( .A(_abc_42016_n1045), .B(_abc_42016_n4033), .C(_abc_42016_n4037), .Y(_abc_42016_n4038) );
  OAI21X1 OAI21X1_1075 ( .A(regfil_4__7_), .B(_abc_42016_n4039), .C(_abc_42016_n4040), .Y(_abc_42016_n4041_1) );
  OAI21X1 OAI21X1_1076 ( .A(_abc_42016_n4038), .B(_abc_42016_n4028), .C(_abc_42016_n4042), .Y(_abc_42016_n4043) );
  OAI21X1 OAI21X1_1077 ( .A(_abc_42016_n583), .B(_abc_42016_n2042), .C(_abc_42016_n4048), .Y(_abc_42016_n4049) );
  OAI21X1 OAI21X1_1078 ( .A(_abc_42016_n960), .B(_abc_42016_n4052), .C(_abc_42016_n1860), .Y(_abc_42016_n4053) );
  OAI21X1 OAI21X1_1079 ( .A(auxcar), .B(_abc_42016_n4066), .C(_abc_42016_n4067), .Y(_abc_42016_n4068) );
  OAI21X1 OAI21X1_108 ( .A(regfil_1__0_), .B(regfil_5__0_), .C(_abc_42016_n1036), .Y(_abc_42016_n1037) );
  OAI21X1 OAI21X1_1080 ( .A(_abc_42016_n4014), .B(_abc_42016_n4044), .C(_abc_42016_n4072), .Y(_abc_42016_n4073) );
  OAI21X1 OAI21X1_1081 ( .A(_abc_42016_n573), .B(_abc_42016_n998), .C(_abc_42016_n1003), .Y(_abc_42016_n4078) );
  OAI21X1 OAI21X1_1082 ( .A(_abc_42016_n604_1), .B(_abc_42016_n1400), .C(_abc_42016_n4080), .Y(_abc_42016_n4081) );
  OAI21X1 OAI21X1_1083 ( .A(_abc_42016_n536), .B(_abc_42016_n539), .C(_abc_42016_n2322), .Y(_abc_42016_n4089) );
  OAI21X1 OAI21X1_1084 ( .A(_abc_42016_n4089), .B(_abc_42016_n4093), .C(pc_0_), .Y(_abc_42016_n4094) );
  OAI21X1 OAI21X1_1085 ( .A(pc_0_), .B(_abc_42016_n4088), .C(_abc_42016_n4094), .Y(_abc_42016_n4095) );
  OAI21X1 OAI21X1_1086 ( .A(_abc_42016_n1060), .B(_abc_42016_n4095), .C(_abc_42016_n675), .Y(_abc_42016_n4096) );
  OAI21X1 OAI21X1_1087 ( .A(_abc_42016_n1463), .B(_abc_42016_n1462), .C(opcode_5_), .Y(_abc_42016_n4098) );
  OAI21X1 OAI21X1_1088 ( .A(_abc_42016_n1935), .B(_abc_42016_n3052), .C(_abc_42016_n2317), .Y(_abc_42016_n4099) );
  OAI21X1 OAI21X1_1089 ( .A(_abc_42016_n4098), .B(_abc_42016_n2089), .C(_abc_42016_n4100), .Y(_abc_42016_n4101) );
  OAI21X1 OAI21X1_109 ( .A(_abc_42016_n1029), .B(_abc_42016_n1037), .C(_abc_42016_n1034), .Y(_abc_42016_n1038) );
  OAI21X1 OAI21X1_1090 ( .A(_abc_42016_n1400), .B(_abc_42016_n2089), .C(_abc_42016_n2286), .Y(_abc_42016_n4106) );
  OAI21X1 OAI21X1_1091 ( .A(_abc_42016_n536), .B(_abc_42016_n539), .C(pc_0_), .Y(_abc_42016_n4115) );
  OAI21X1 OAI21X1_1092 ( .A(_abc_42016_n4115), .B(_abc_42016_n4114), .C(_abc_42016_n559), .Y(_abc_42016_n4116) );
  OAI21X1 OAI21X1_1093 ( .A(_abc_42016_n4097), .B(_abc_42016_n4117), .C(_abc_42016_n547), .Y(_abc_42016_n4118) );
  OAI21X1 OAI21X1_1094 ( .A(_abc_42016_n511), .B(_abc_42016_n525), .C(_abc_42016_n3460), .Y(_abc_42016_n4119) );
  OAI21X1 OAI21X1_1095 ( .A(_abc_42016_n536), .B(_abc_42016_n539), .C(_abc_42016_n4114), .Y(_abc_42016_n4128) );
  OAI21X1 OAI21X1_1096 ( .A(_abc_42016_n4092_1), .B(_abc_42016_n4090), .C(_abc_42016_n673), .Y(_abc_42016_n4131) );
  OAI21X1 OAI21X1_1097 ( .A(_abc_42016_n2526), .B(_abc_42016_n4076), .C(_abc_42016_n4134), .Y(_abc_42016_n4135) );
  OAI21X1 OAI21X1_1098 ( .A(_abc_42016_n1383), .B(_abc_42016_n4130), .C(_abc_42016_n4136), .Y(_abc_42016_n4137) );
  OAI21X1 OAI21X1_1099 ( .A(_abc_42016_n4126), .B(_abc_42016_n4137), .C(_abc_42016_n547), .Y(_abc_42016_n4138) );
  OAI21X1 OAI21X1_11 ( .A(opcode_5_), .B(_abc_42016_n528_1), .C(_abc_42016_n595), .Y(_abc_42016_n596) );
  OAI21X1 OAI21X1_110 ( .A(_abc_42016_n1023), .B(_abc_42016_n1038), .C(_abc_42016_n1027), .Y(_abc_42016_n1039) );
  OAI21X1 OAI21X1_1100 ( .A(_abc_42016_n2347_1), .B(_abc_42016_n2283), .C(_abc_42016_n2573), .Y(_abc_42016_n4141) );
  OAI21X1 OAI21X1_1101 ( .A(_abc_42016_n560), .B(_abc_42016_n4145), .C(_abc_42016_n3497_1), .Y(_abc_42016_n4146) );
  OAI21X1 OAI21X1_1102 ( .A(_abc_42016_n1376), .B(_abc_42016_n4075), .C(_abc_42016_n2573), .Y(_abc_42016_n4147) );
  OAI21X1 OAI21X1_1103 ( .A(_abc_42016_n1841), .B(_abc_42016_n2323_1), .C(_abc_42016_n4142), .Y(_abc_42016_n4148) );
  OAI21X1 OAI21X1_1104 ( .A(_abc_42016_n1382), .B(_abc_42016_n4130), .C(_abc_42016_n4151), .Y(_abc_42016_n4152) );
  OAI21X1 OAI21X1_1105 ( .A(_abc_42016_n4144), .B(_abc_42016_n4152), .C(_abc_42016_n547), .Y(_abc_42016_n4153) );
  OAI21X1 OAI21X1_1106 ( .A(_abc_42016_n4086), .B(_abc_42016_n4131), .C(_abc_42016_n4156), .Y(_abc_42016_n4157) );
  OAI21X1 OAI21X1_1107 ( .A(_abc_42016_n1382), .B(_abc_42016_n1383), .C(_abc_42016_n1357), .Y(_abc_42016_n4160) );
  OAI21X1 OAI21X1_1108 ( .A(_abc_42016_n2606), .B(_abc_42016_n999), .C(_abc_42016_n2085), .Y(_abc_42016_n4164) );
  OAI21X1 OAI21X1_1109 ( .A(_abc_42016_n2590), .B(_abc_42016_n4076), .C(_abc_42016_n4165), .Y(_abc_42016_n4166) );
  OAI21X1 OAI21X1_111 ( .A(_abc_42016_n670), .B(_abc_42016_n996), .C(_abc_42016_n561), .Y(_abc_42016_n1040) );
  OAI21X1 OAI21X1_1110 ( .A(_abc_42016_n1357), .B(_abc_42016_n4130), .C(_abc_42016_n4167), .Y(_abc_42016_n4168) );
  OAI21X1 OAI21X1_1111 ( .A(_abc_42016_n4168), .B(_abc_42016_n4159), .C(_abc_42016_n547), .Y(_abc_42016_n4169) );
  OAI21X1 OAI21X1_1112 ( .A(_abc_42016_n2635), .B(_abc_42016_n2423_1), .C(_abc_42016_n4174), .Y(_abc_42016_n4175) );
  OAI21X1 OAI21X1_1113 ( .A(_abc_42016_n531), .B(_abc_42016_n1380), .C(_abc_42016_n1246), .Y(_abc_42016_n4176) );
  OAI21X1 OAI21X1_1114 ( .A(_abc_42016_n2635), .B(_abc_42016_n4076), .C(_abc_42016_n4177), .Y(_abc_42016_n4178) );
  OAI21X1 OAI21X1_1115 ( .A(_abc_42016_n1356), .B(_abc_42016_n4130), .C(_abc_42016_n4179), .Y(_abc_42016_n4180) );
  OAI21X1 OAI21X1_1116 ( .A(_abc_42016_n4180), .B(_abc_42016_n4172), .C(_abc_42016_n547), .Y(_abc_42016_n4181) );
  OAI21X1 OAI21X1_1117 ( .A(_abc_42016_n1356), .B(_abc_42016_n1385), .C(_abc_42016_n2649), .Y(_abc_42016_n4186) );
  OAI21X1 OAI21X1_1118 ( .A(_abc_42016_n872), .B(_abc_42016_n1046), .C(_abc_42016_n4098), .Y(_abc_42016_n4190) );
  OAI21X1 OAI21X1_1119 ( .A(_abc_42016_n4185), .B(_abc_42016_n4076), .C(_abc_42016_n4191), .Y(_abc_42016_n4192) );
  OAI21X1 OAI21X1_112 ( .A(regfil_5__0_), .B(_abc_42016_n1040), .C(_abc_42016_n994), .Y(_abc_42016_n1041) );
  OAI21X1 OAI21X1_1120 ( .A(_abc_42016_n2649), .B(_abc_42016_n4130), .C(_abc_42016_n4193), .Y(_abc_42016_n4194) );
  OAI21X1 OAI21X1_1121 ( .A(_abc_42016_n4194), .B(_abc_42016_n4184), .C(_abc_42016_n547), .Y(_abc_42016_n4195) );
  OAI21X1 OAI21X1_1122 ( .A(_abc_42016_n2649), .B(_abc_42016_n2630), .C(_abc_42016_n1355), .Y(_abc_42016_n4199) );
  OAI21X1 OAI21X1_1123 ( .A(_abc_42016_n2423_1), .B(_abc_42016_n2688), .C(_abc_42016_n4201), .Y(_abc_42016_n4202) );
  OAI21X1 OAI21X1_1124 ( .A(_abc_42016_n4076), .B(_abc_42016_n2688), .C(_abc_42016_n4203), .Y(_abc_42016_n4204_1) );
  OAI21X1 OAI21X1_1125 ( .A(_abc_42016_n1355), .B(_abc_42016_n4130), .C(_abc_42016_n4205), .Y(_abc_42016_n4206) );
  OAI21X1 OAI21X1_1126 ( .A(_abc_42016_n4206), .B(_abc_42016_n4198), .C(_abc_42016_n547), .Y(_abc_42016_n4207) );
  OAI21X1 OAI21X1_1127 ( .A(_abc_42016_n1355), .B(_abc_42016_n1387), .C(_abc_42016_n1354), .Y(_abc_42016_n4211) );
  OAI21X1 OAI21X1_1128 ( .A(_abc_42016_n1841), .B(_abc_42016_n2323_1), .C(_abc_42016_n4212), .Y(_abc_42016_n4214) );
  OAI21X1 OAI21X1_1129 ( .A(_abc_42016_n959), .B(_abc_42016_n1046), .C(_abc_42016_n4214), .Y(_abc_42016_n4215) );
  OAI21X1 OAI21X1_113 ( .A(_abc_42016_n1021), .B(_abc_42016_n991), .C(_abc_42016_n1053), .Y(_abc_36783_n3435) );
  OAI21X1 OAI21X1_1130 ( .A(_abc_42016_n2716), .B(_abc_42016_n4158), .C(_abc_42016_n4218), .Y(_abc_42016_n4219) );
  OAI21X1 OAI21X1_1131 ( .A(_abc_42016_n1354), .B(_abc_42016_n2674), .C(_abc_42016_n1353), .Y(_abc_42016_n4224) );
  OAI21X1 OAI21X1_1132 ( .A(_abc_42016_n4131), .B(_abc_42016_n4228), .C(_abc_42016_n4231), .Y(_abc_42016_n4232) );
  OAI21X1 OAI21X1_1133 ( .A(_abc_42016_n4232), .B(_abc_42016_n4223), .C(_abc_42016_n547), .Y(_abc_42016_n4233) );
  OAI21X1 OAI21X1_1134 ( .A(_abc_42016_n1353), .B(_abc_42016_n1389), .C(_abc_42016_n1422), .Y(_abc_42016_n4237) );
  OAI21X1 OAI21X1_1135 ( .A(_abc_42016_n1422), .B(_abc_42016_n4130), .C(_abc_42016_n4244), .Y(_abc_42016_n4245) );
  OAI21X1 OAI21X1_1136 ( .A(_abc_42016_n4241), .B(_abc_42016_n4245), .C(_abc_42016_n547), .Y(_abc_42016_n4246) );
  OAI21X1 OAI21X1_1137 ( .A(_abc_42016_n560), .B(_abc_42016_n4255), .C(_abc_42016_n4256), .Y(_abc_42016_n4257) );
  OAI21X1 OAI21X1_1138 ( .A(_abc_42016_n4254), .B(_abc_42016_n4257), .C(_abc_42016_n547), .Y(_abc_42016_n4258) );
  OAI21X1 OAI21X1_1139 ( .A(_abc_42016_n1449), .B(_abc_42016_n1424), .C(_abc_42016_n1477), .Y(_abc_42016_n4262) );
  OAI21X1 OAI21X1_114 ( .A(_abc_42016_n992), .B(_abc_42016_n585), .C(_abc_42016_n1056), .Y(_abc_42016_n1057) );
  OAI21X1 OAI21X1_1140 ( .A(_abc_42016_n1485), .B(_abc_42016_n4076), .C(_abc_42016_n4265), .Y(_abc_42016_n4266_1) );
  OAI21X1 OAI21X1_1141 ( .A(_abc_42016_n1481), .B(_abc_42016_n4156), .C(_abc_42016_n4270), .Y(_abc_42016_n4271) );
  OAI21X1 OAI21X1_1142 ( .A(_abc_42016_n4268), .B(_abc_42016_n4271), .C(_abc_42016_n547), .Y(_abc_42016_n4272) );
  OAI21X1 OAI21X1_1143 ( .A(_abc_42016_n1477), .B(_abc_42016_n1478), .C(_abc_42016_n1503), .Y(_abc_42016_n4275) );
  OAI21X1 OAI21X1_1144 ( .A(_abc_42016_n842), .B(_abc_42016_n1046), .C(_abc_42016_n4278), .Y(_abc_42016_n4279) );
  OAI21X1 OAI21X1_1145 ( .A(_abc_42016_n1503), .B(_abc_42016_n4130), .C(_abc_42016_n4282), .Y(_abc_42016_n4283) );
  OAI21X1 OAI21X1_1146 ( .A(_abc_42016_n4283), .B(_abc_42016_n4280), .C(_abc_42016_n547), .Y(_abc_42016_n4284) );
  OAI21X1 OAI21X1_1147 ( .A(_abc_42016_n1503), .B(_abc_42016_n1480), .C(_abc_42016_n1530), .Y(_abc_42016_n4287) );
  OAI21X1 OAI21X1_1148 ( .A(_abc_42016_n4291), .B(_abc_42016_n4292), .C(_abc_42016_n4132), .Y(_abc_42016_n4293) );
  OAI21X1 OAI21X1_1149 ( .A(_abc_42016_n4290), .B(_abc_42016_n4295), .C(_abc_42016_n547), .Y(_abc_42016_n4296) );
  OAI21X1 OAI21X1_115 ( .A(_abc_42016_n1010), .B(_abc_42016_n696), .C(_abc_42016_n994), .Y(_abc_42016_n1058) );
  OAI21X1 OAI21X1_1150 ( .A(_abc_42016_n4091), .B(_abc_42016_n4300), .C(_abc_42016_n4302), .Y(_abc_42016_n4303) );
  OAI21X1 OAI21X1_1151 ( .A(_abc_42016_n2424), .B(_abc_42016_n4113), .C(_abc_42016_n559), .Y(_abc_42016_n4305) );
  OAI21X1 OAI21X1_1152 ( .A(_abc_42016_n4304), .B(_abc_42016_n4308), .C(_abc_42016_n547), .Y(_abc_42016_n4309) );
  OAI21X1 OAI21X1_1153 ( .A(_abc_42016_n547), .B(_abc_42016_n4119), .C(_abc_42016_n4310), .Y(_abc_42016_n4311) );
  OAI21X1 OAI21X1_1154 ( .A(_abc_42016_n1376), .B(_abc_42016_n4075), .C(_abc_42016_n1589), .Y(_abc_42016_n4314) );
  OAI21X1 OAI21X1_1155 ( .A(_abc_42016_n4305), .B(_abc_42016_n4317), .C(_abc_42016_n4318), .Y(_abc_42016_n4319) );
  OAI21X1 OAI21X1_1156 ( .A(_abc_42016_n4316), .B(_abc_42016_n4319), .C(_abc_42016_n547), .Y(_abc_42016_n4320_1) );
  OAI21X1 OAI21X1_1157 ( .A(_abc_42016_n2031), .B(_abc_42016_n546), .C(_abc_42016_n2228), .Y(_abc_42016_n4327) );
  OAI21X1 OAI21X1_1158 ( .A(reset), .B(_abc_42016_n4327), .C(_abc_42016_n4326), .Y(_abc_42016_n4328) );
  OAI21X1 OAI21X1_1159 ( .A(_auto_iopadmap_cc_313_execute_46274), .B(_abc_42016_n4324), .C(_abc_42016_n4328), .Y(_abc_42016_n4329) );
  OAI21X1 OAI21X1_116 ( .A(_abc_42016_n1065), .B(_abc_42016_n1061), .C(_abc_42016_n671_1), .Y(_abc_42016_n1066) );
  OAI21X1 OAI21X1_1160 ( .A(_abc_42016_n1375), .B(_abc_42016_n4330), .C(_abc_42016_n4329), .Y(inta_FF_INPUT) );
  OAI21X1 OAI21X1_1161 ( .A(_abc_42016_n4335), .B(_abc_42016_n4334), .C(_abc_42016_n4332), .Y(writeio_FF_INPUT) );
  OAI21X1 OAI21X1_1162 ( .A(waitr), .B(_abc_42016_n4046), .C(_auto_iopadmap_cc_313_execute_46276), .Y(_abc_42016_n4338) );
  OAI21X1 OAI21X1_1163 ( .A(reset), .B(_abc_42016_n4338), .C(_abc_42016_n4337), .Y(readio_FF_INPUT) );
  OAI21X1 OAI21X1_1164 ( .A(regfil_7__0_), .B(_abc_42016_n4340), .C(_abc_42016_n4341), .Y(_abc_42016_n4342) );
  OAI21X1 OAI21X1_1165 ( .A(rdatahold_0_), .B(_abc_42016_n4047), .C(_abc_42016_n4049), .Y(_abc_42016_n4343) );
  OAI21X1 OAI21X1_1166 ( .A(_abc_42016_n1427), .B(_abc_42016_n4060), .C(_abc_42016_n4343), .Y(_abc_42016_n4344) );
  OAI21X1 OAI21X1_1167 ( .A(auxcar), .B(_abc_42016_n4066), .C(_abc_42016_n4348), .Y(_abc_42016_n4349) );
  OAI21X1 OAI21X1_1168 ( .A(_abc_42016_n628), .B(_abc_42016_n4349), .C(_abc_42016_n4352), .Y(_abc_42016_n4353) );
  OAI21X1 OAI21X1_1169 ( .A(_abc_42016_n1860), .B(_abc_42016_n4345), .C(_abc_42016_n4354), .Y(_abc_42016_n4355) );
  OAI21X1 OAI21X1_117 ( .A(_abc_42016_n1068), .B(_abc_42016_n1070_1), .C(_abc_42016_n1024), .Y(_abc_42016_n1071) );
  OAI21X1 OAI21X1_1170 ( .A(_abc_42016_n2234), .B(_abc_42016_n4048), .C(_abc_42016_n4359), .Y(_abc_42016_n4360) );
  OAI21X1 OAI21X1_1171 ( .A(regfil_7__1_), .B(_abc_42016_n4070), .C(_abc_42016_n4363), .Y(_abc_42016_n4364) );
  OAI21X1 OAI21X1_1172 ( .A(regfil_7__1_), .B(_abc_42016_n4340), .C(_abc_42016_n4369), .Y(_abc_42016_n4370) );
  OAI21X1 OAI21X1_1173 ( .A(_abc_42016_n4370), .B(_abc_42016_n4368), .C(_abc_42016_n4366), .Y(_abc_36783_n4580) );
  OAI21X1 OAI21X1_1174 ( .A(regfil_7__2_), .B(_abc_42016_n4340), .C(_abc_42016_n4372), .Y(_abc_42016_n4373) );
  OAI21X1 OAI21X1_1175 ( .A(_abc_42016_n2237), .B(_abc_42016_n4048), .C(_abc_42016_n4374), .Y(_abc_42016_n4375) );
  OAI21X1 OAI21X1_1176 ( .A(_abc_42016_n1454), .B(_abc_42016_n4349), .C(_abc_42016_n4051), .Y(_abc_42016_n4377) );
  OAI21X1 OAI21X1_1177 ( .A(_abc_42016_n669), .B(_abc_42016_n4064), .C(_abc_42016_n4349), .Y(_abc_42016_n4378) );
  OAI21X1 OAI21X1_1178 ( .A(_abc_42016_n1427), .B(_abc_42016_n4349), .C(_abc_42016_n1454), .Y(_abc_42016_n4380) );
  OAI21X1 OAI21X1_1179 ( .A(_abc_42016_n4380), .B(_abc_42016_n4379), .C(_abc_42016_n4383), .Y(_abc_42016_n4384) );
  OAI21X1 OAI21X1_118 ( .A(_abc_42016_n1078), .B(_abc_42016_n1081), .C(_abc_42016_n1083), .Y(_abc_42016_n1084) );
  OAI21X1 OAI21X1_1180 ( .A(regfil_7__3_), .B(_abc_42016_n4340), .C(_abc_42016_n4387), .Y(_abc_42016_n4388) );
  OAI21X1 OAI21X1_1181 ( .A(_abc_42016_n2240), .B(_abc_42016_n4048), .C(_abc_42016_n4389), .Y(_abc_42016_n4390) );
  OAI21X1 OAI21X1_1182 ( .A(_abc_42016_n4069), .B(_abc_42016_n4065), .C(_abc_42016_n1488), .Y(_abc_42016_n4395) );
  OAI21X1 OAI21X1_1183 ( .A(_abc_42016_n811), .B(_abc_42016_n4392), .C(_abc_42016_n4398), .Y(_abc_42016_n4399) );
  OAI21X1 OAI21X1_1184 ( .A(_abc_42016_n4367), .B(_abc_42016_n858), .C(_abc_42016_n4369), .Y(_abc_42016_n4403_1) );
  OAI21X1 OAI21X1_1185 ( .A(_abc_42016_n4066), .B(_abc_42016_n4068), .C(_abc_42016_n1974), .Y(_abc_42016_n4404) );
  OAI21X1 OAI21X1_1186 ( .A(_abc_42016_n1974), .B(_abc_42016_n4405), .C(_abc_42016_n4406), .Y(_abc_42016_n4407) );
  OAI21X1 OAI21X1_1187 ( .A(_abc_42016_n4379), .B(_abc_42016_n4404), .C(_abc_42016_n4408), .Y(_abc_42016_n4409) );
  OAI21X1 OAI21X1_1188 ( .A(_abc_42016_n1974), .B(_abc_42016_n4055), .C(_abc_42016_n4410), .Y(_abc_42016_n4411) );
  OAI21X1 OAI21X1_1189 ( .A(_abc_42016_n4402), .B(_abc_42016_n4403_1), .C(_abc_42016_n4412), .Y(_abc_36783_n4583) );
  OAI21X1 OAI21X1_119 ( .A(_abc_42016_n1035), .B(_abc_42016_n1077), .C(_abc_42016_n1084), .Y(_abc_42016_n1085) );
  OAI21X1 OAI21X1_1190 ( .A(_abc_42016_n2067), .B(_abc_42016_n4068), .C(_abc_42016_n898), .Y(_abc_42016_n4414) );
  OAI21X1 OAI21X1_1191 ( .A(_abc_42016_n1974), .B(_abc_42016_n2066), .C(_abc_42016_n4350), .Y(_abc_42016_n4415) );
  OAI21X1 OAI21X1_1192 ( .A(_abc_42016_n898), .B(_abc_42016_n4415), .C(_abc_42016_n4416_1), .Y(_abc_42016_n4417) );
  OAI21X1 OAI21X1_1193 ( .A(_abc_42016_n4379), .B(_abc_42016_n4414), .C(_abc_42016_n4418), .Y(_abc_42016_n4419) );
  OAI21X1 OAI21X1_1194 ( .A(regfil_7__5_), .B(_abc_42016_n4055), .C(_abc_42016_n4420), .Y(_abc_42016_n4421) );
  OAI21X1 OAI21X1_1195 ( .A(regfil_7__5_), .B(_abc_42016_n4340), .C(_abc_42016_n4369), .Y(_abc_42016_n4424) );
  OAI21X1 OAI21X1_1196 ( .A(_abc_42016_n4424), .B(_abc_42016_n4423), .C(_abc_42016_n4422), .Y(_abc_36783_n4584) );
  OAI21X1 OAI21X1_1197 ( .A(_abc_42016_n4367), .B(_abc_42016_n934), .C(_abc_42016_n4369), .Y(_abc_42016_n4427) );
  OAI21X1 OAI21X1_1198 ( .A(regfil_7__5_), .B(_abc_42016_n4349), .C(_abc_42016_n4415), .Y(_abc_42016_n4428) );
  OAI21X1 OAI21X1_1199 ( .A(_abc_42016_n924), .B(_abc_42016_n4428), .C(_abc_42016_n4429), .Y(_abc_42016_n4430) );
  OAI21X1 OAI21X1_12 ( .A(_abc_42016_n621), .B(_abc_42016_n620), .C(_abc_42016_n607), .Y(_abc_42016_n622) );
  OAI21X1 OAI21X1_120 ( .A(_abc_42016_n671_1), .B(_abc_42016_n1065), .C(_abc_42016_n561), .Y(_abc_42016_n1087) );
  OAI21X1 OAI21X1_1200 ( .A(_abc_42016_n898), .B(_abc_42016_n4051), .C(_abc_42016_n4431_1), .Y(_abc_42016_n4432) );
  OAI21X1 OAI21X1_1201 ( .A(_abc_42016_n4434), .B(_abc_42016_n4052), .C(_abc_42016_n4056), .Y(_abc_42016_n4435) );
  OAI21X1 OAI21X1_1202 ( .A(_abc_42016_n4426), .B(_abc_42016_n4427), .C(_abc_42016_n4439), .Y(_abc_36783_n4585) );
  OAI21X1 OAI21X1_1203 ( .A(_abc_42016_n2478), .B(_abc_42016_n4392), .C(_abc_42016_n4442), .Y(_abc_42016_n4443) );
  OAI21X1 OAI21X1_1204 ( .A(_abc_42016_n924), .B(_abc_42016_n2068), .C(_abc_42016_n4069), .Y(_abc_42016_n4448) );
  OAI21X1 OAI21X1_1205 ( .A(_abc_42016_n960), .B(_abc_42016_n4448), .C(_abc_42016_n4450), .Y(_abc_42016_n4451) );
  OAI21X1 OAI21X1_1206 ( .A(_abc_42016_n2069), .B(_abc_42016_n4068), .C(_abc_42016_n960), .Y(_abc_42016_n4452) );
  OAI21X1 OAI21X1_1207 ( .A(_abc_42016_n4451), .B(_abc_42016_n4453), .C(_abc_42016_n4447_1), .Y(_abc_42016_n4454) );
  OAI21X1 OAI21X1_1208 ( .A(_abc_42016_n556), .B(_abc_42016_n1814), .C(_abc_42016_n960), .Y(_abc_42016_n4455) );
  OAI21X1 OAI21X1_1209 ( .A(_abc_42016_n4367), .B(_abc_42016_n971), .C(_abc_42016_n4455), .Y(_abc_42016_n4456) );
  OAI21X1 OAI21X1_121 ( .A(_abc_42016_n703), .B(_abc_42016_n697), .C(_abc_42016_n1089), .Y(_abc_42016_n1090) );
  OAI21X1 OAI21X1_1210 ( .A(waitr), .B(_abc_42016_n4460), .C(_auto_iopadmap_cc_313_execute_46282), .Y(_abc_42016_n4461) );
  OAI21X1 OAI21X1_1211 ( .A(reset), .B(_abc_42016_n4461), .C(_abc_42016_n4458), .Y(writemem_FF_INPUT) );
  OAI21X1 OAI21X1_1212 ( .A(intcyc), .B(_abc_42016_n2733), .C(_abc_42016_n4463_1), .Y(_abc_42016_n4464) );
  OAI21X1 OAI21X1_1213 ( .A(_abc_42016_n2031), .B(_abc_42016_n2079), .C(_abc_42016_n2024), .Y(_abc_42016_n4467) );
  OAI21X1 OAI21X1_1214 ( .A(_abc_42016_n2031), .B(_abc_42016_n2033), .C(_abc_42016_n4468), .Y(_abc_42016_n4469) );
  OAI21X1 OAI21X1_1215 ( .A(_abc_42016_n4467), .B(_abc_42016_n4469), .C(_abc_42016_n529), .Y(_abc_42016_n4470) );
  OAI21X1 OAI21X1_1216 ( .A(reset), .B(_abc_42016_n2497), .C(_abc_42016_n4470), .Y(_abc_42016_n4471) );
  OAI21X1 OAI21X1_1217 ( .A(_abc_42016_n602), .B(_abc_42016_n4472), .C(_abc_42016_n4474), .Y(_abc_42016_n4475) );
  OAI21X1 OAI21X1_1218 ( .A(_abc_42016_n2779), .B(_abc_42016_n4475), .C(_abc_42016_n4471), .Y(_abc_42016_n4476) );
  OAI21X1 OAI21X1_1219 ( .A(_abc_42016_n4466), .B(_abc_42016_n4471), .C(_abc_42016_n4476), .Y(addr_0__FF_INPUT) );
  OAI21X1 OAI21X1_122 ( .A(_abc_42016_n1055), .B(_abc_42016_n1092), .C(_abc_42016_n1091), .Y(_abc_36783_n3438) );
  OAI21X1 OAI21X1_1220 ( .A(_abc_42016_n1383), .B(_abc_42016_n2024), .C(_abc_42016_n4479_1), .Y(_abc_42016_n4480) );
  OAI21X1 OAI21X1_1221 ( .A(_abc_42016_n4480), .B(_abc_42016_n4481), .C(_abc_42016_n4471), .Y(_abc_42016_n4482) );
  OAI21X1 OAI21X1_1222 ( .A(_abc_42016_n4478), .B(_abc_42016_n4471), .C(_abc_42016_n4482), .Y(addr_1__FF_INPUT) );
  OAI21X1 OAI21X1_1223 ( .A(_abc_42016_n4485), .B(_abc_42016_n4486), .C(_abc_42016_n4471), .Y(_abc_42016_n4487) );
  OAI21X1 OAI21X1_1224 ( .A(_abc_42016_n4484), .B(_abc_42016_n4471), .C(_abc_42016_n4487), .Y(addr_2__FF_INPUT) );
  OAI21X1 OAI21X1_1225 ( .A(_abc_42016_n4490), .B(_abc_42016_n4491), .C(_abc_42016_n4471), .Y(_abc_42016_n4492) );
  OAI21X1 OAI21X1_1226 ( .A(_abc_42016_n4489), .B(_abc_42016_n4471), .C(_abc_42016_n4492), .Y(addr_3__FF_INPUT) );
  OAI21X1 OAI21X1_1227 ( .A(_abc_42016_n4495), .B(_abc_42016_n4496), .C(_abc_42016_n4471), .Y(_abc_42016_n4497) );
  OAI21X1 OAI21X1_1228 ( .A(_abc_42016_n4494_1), .B(_abc_42016_n4471), .C(_abc_42016_n4497), .Y(addr_4__FF_INPUT) );
  OAI21X1 OAI21X1_1229 ( .A(_abc_42016_n4500), .B(_abc_42016_n4501), .C(_abc_42016_n4471), .Y(_abc_42016_n4502) );
  OAI21X1 OAI21X1_123 ( .A(_abc_42016_n556), .B(_abc_42016_n988), .C(regfil_5__2_), .Y(_abc_42016_n1094) );
  OAI21X1 OAI21X1_1230 ( .A(_abc_42016_n4499), .B(_abc_42016_n4471), .C(_abc_42016_n4502), .Y(addr_5__FF_INPUT) );
  OAI21X1 OAI21X1_1231 ( .A(_abc_42016_n4505), .B(_abc_42016_n4506), .C(_abc_42016_n4471), .Y(_abc_42016_n4507) );
  OAI21X1 OAI21X1_1232 ( .A(_abc_42016_n4504), .B(_abc_42016_n4471), .C(_abc_42016_n4507), .Y(addr_6__FF_INPUT) );
  OAI21X1 OAI21X1_1233 ( .A(_abc_42016_n4510), .B(_abc_42016_n4511), .C(_abc_42016_n4471), .Y(_abc_42016_n4512) );
  OAI21X1 OAI21X1_1234 ( .A(_abc_42016_n4509_1), .B(_abc_42016_n4471), .C(_abc_42016_n4512), .Y(addr_7__FF_INPUT) );
  OAI21X1 OAI21X1_1235 ( .A(_abc_42016_n4515), .B(_abc_42016_n4516), .C(_abc_42016_n4471), .Y(_abc_42016_n4517) );
  OAI21X1 OAI21X1_1236 ( .A(_abc_42016_n4514), .B(_abc_42016_n4471), .C(_abc_42016_n4517), .Y(addr_8__FF_INPUT) );
  OAI21X1 OAI21X1_1237 ( .A(_abc_42016_n4536), .B(_abc_42016_n4537), .C(_abc_42016_n4471), .Y(_abc_42016_n4538) );
  OAI21X1 OAI21X1_1238 ( .A(_abc_42016_n4535), .B(_abc_42016_n4471), .C(_abc_42016_n4538), .Y(addr_13__FF_INPUT) );
  OAI21X1 OAI21X1_1239 ( .A(_abc_42016_n3388), .B(_abc_42016_n2497), .C(_abc_42016_n3023), .Y(_abc_42016_n4544) );
  OAI21X1 OAI21X1_124 ( .A(_abc_42016_n709), .B(_abc_42016_n1046), .C(_abc_42016_n1022), .Y(_abc_42016_n1098) );
  OAI21X1 OAI21X1_1240 ( .A(reset), .B(_abc_42016_n2276), .C(_abc_42016_n2462), .Y(_abc_42016_n4550) );
  OAI21X1 OAI21X1_1241 ( .A(_abc_42016_n4326), .B(_abc_42016_n4333), .C(_abc_42016_n4332), .Y(_abc_42016_n4554_1) );
  OAI21X1 OAI21X1_1242 ( .A(_abc_42016_n4555), .B(_abc_42016_n4560), .C(_abc_42016_n4562), .Y(_abc_42016_n4563) );
  OAI21X1 OAI21X1_1243 ( .A(_abc_42016_n4567), .B(_abc_42016_n4570_1), .C(_abc_42016_n4571), .Y(_abc_42016_n4572) );
  OAI21X1 OAI21X1_1244 ( .A(reset), .B(_abc_42016_n2497), .C(_abc_42016_n4572), .Y(_abc_42016_n4573) );
  OAI21X1 OAI21X1_1245 ( .A(_abc_42016_n4567), .B(_abc_42016_n2438_1), .C(_abc_42016_n4578), .Y(_abc_42016_n4579) );
  OAI21X1 OAI21X1_1246 ( .A(_abc_42016_n2451), .B(_abc_42016_n4583), .C(_abc_42016_n4579), .Y(_abc_42016_n4584) );
  OAI21X1 OAI21X1_1247 ( .A(_abc_42016_n4577), .B(_abc_42016_n4560), .C(_abc_42016_n4585_1), .Y(_abc_42016_n4586) );
  OAI21X1 OAI21X1_1248 ( .A(_abc_42016_n4588), .B(_abc_42016_n4560), .C(_abc_42016_n4590), .Y(_abc_42016_n4591) );
  OAI21X1 OAI21X1_1249 ( .A(_abc_42016_n4596), .B(_abc_42016_n4560), .C(_abc_42016_n4597), .Y(_abc_42016_n4598) );
  OAI21X1 OAI21X1_125 ( .A(_abc_42016_n1033), .B(_abc_42016_n1080), .C(_abc_42016_n1099), .Y(_abc_42016_n1100) );
  OAI21X1 OAI21X1_1250 ( .A(_abc_42016_n4577), .B(_abc_42016_n4593), .C(_abc_42016_n4606), .Y(_abc_42016_n4607) );
  OAI21X1 OAI21X1_1251 ( .A(_abc_42016_n4566), .B(_abc_42016_n4614), .C(_abc_42016_n4613), .Y(_abc_42016_n4615_1) );
  OAI21X1 OAI21X1_1252 ( .A(_abc_42016_n4326), .B(_abc_42016_n4460), .C(_abc_42016_n4458), .Y(_abc_42016_n4617) );
  OAI21X1 OAI21X1_1253 ( .A(_abc_42016_n2026), .B(_abc_42016_n4334), .C(_abc_42016_n529), .Y(_abc_42016_n4619) );
  OAI21X1 OAI21X1_1254 ( .A(_abc_42016_n4602), .B(_abc_42016_n4593), .C(_abc_42016_n4623), .Y(_abc_42016_n4624) );
  OAI21X1 OAI21X1_1255 ( .A(_abc_42016_n999), .B(_abc_42016_n2089), .C(_abc_42016_n3034), .Y(_abc_42016_n4632_1) );
  OAI21X1 OAI21X1_1256 ( .A(_abc_42016_n2738), .B(_abc_42016_n4635), .C(_abc_42016_n4631_1), .Y(_abc_42016_n4636) );
  OAI21X1 OAI21X1_1257 ( .A(opcode_5_), .B(carry), .C(_abc_42016_n4643), .Y(_abc_42016_n4644) );
  OAI21X1 OAI21X1_1258 ( .A(opcode_5_), .B(_abc_42016_n4639), .C(_abc_42016_n4646_1), .Y(_abc_42016_n4647) );
  OAI21X1 OAI21X1_1259 ( .A(_abc_42016_n630), .B(_abc_42016_n4075), .C(_abc_42016_n4647), .Y(_abc_42016_n4648) );
  OAI21X1 OAI21X1_126 ( .A(_abc_42016_n1100), .B(_abc_42016_n1103_1), .C(_abc_42016_n1000), .Y(_abc_42016_n1105) );
  OAI21X1 OAI21X1_1260 ( .A(_abc_42016_n604_1), .B(_abc_42016_n682), .C(_abc_42016_n4091), .Y(_abc_42016_n4649) );
  OAI21X1 OAI21X1_1261 ( .A(_abc_42016_n2309), .B(_abc_42016_n2424), .C(_abc_42016_n561), .Y(_abc_42016_n4654_1) );
  OAI21X1 OAI21X1_1262 ( .A(_abc_42016_n2409), .B(_abc_42016_n2407), .C(_abc_42016_n4657_1), .Y(_abc_42016_n4658) );
  OAI21X1 OAI21X1_1263 ( .A(_abc_42016_n4658), .B(_abc_42016_n4656), .C(_abc_42016_n4551), .Y(_abc_42016_n4659) );
  OAI21X1 OAI21X1_1264 ( .A(_abc_42016_n4548), .B(_abc_42016_n4566), .C(_abc_42016_n4660), .Y(_abc_42016_n4661_1) );
  OAI21X1 OAI21X1_1265 ( .A(_abc_42016_n2452), .B(_abc_42016_n4667), .C(_abc_42016_n4550), .Y(_abc_42016_n4668_1) );
  OAI21X1 OAI21X1_1266 ( .A(_abc_42016_n558), .B(_abc_42016_n2070), .C(_abc_42016_n4672_1), .Y(_abc_42016_n4673) );
  OAI21X1 OAI21X1_1267 ( .A(statesel_1_), .B(_abc_42016_n2437), .C(_abc_42016_n4596), .Y(_abc_42016_n4675) );
  OAI21X1 OAI21X1_1268 ( .A(_abc_42016_n4677), .B(_abc_42016_n4601), .C(_abc_42016_n4551), .Y(_abc_42016_n4678_1) );
  OAI21X1 OAI21X1_1269 ( .A(statesel_0_), .B(_abc_42016_n2344), .C(_abc_42016_n4657_1), .Y(_abc_42016_n4679) );
  OAI21X1 OAI21X1_127 ( .A(_abc_42016_n1028), .B(_abc_42016_n1074), .C(_abc_42016_n1106_1), .Y(_abc_42016_n1107_1) );
  OAI21X1 OAI21X1_1270 ( .A(_abc_42016_n1408), .B(_abc_42016_n678), .C(_abc_42016_n4682), .Y(_abc_42016_n4683) );
  OAI21X1 OAI21X1_1271 ( .A(_abc_42016_n4691), .B(_abc_42016_n4556), .C(_abc_42016_n3418), .Y(_abc_42016_n4692) );
  OAI21X1 OAI21X1_1272 ( .A(_abc_42016_n4638), .B(_abc_42016_n4694), .C(_abc_42016_n4610), .Y(_abc_36783_n4644) );
  OAI21X1 OAI21X1_1273 ( .A(_abc_42016_n4588), .B(_abc_42016_n4593), .C(_abc_42016_n4686), .Y(_abc_42016_n4696) );
  OAI21X1 OAI21X1_1274 ( .A(reset), .B(_abc_42016_n2024), .C(_abc_42016_n4599), .Y(_abc_42016_n4697) );
  OAI21X1 OAI21X1_1275 ( .A(_abc_42016_n4577), .B(_abc_42016_n4593), .C(_abc_42016_n4712), .Y(_abc_42016_n4713_1) );
  OAI21X1 OAI21X1_1276 ( .A(_abc_42016_n2231), .B(_abc_42016_n4460), .C(_abc_42016_n4720), .Y(_abc_42016_n4721) );
  OAI21X1 OAI21X1_1277 ( .A(reset), .B(_abc_42016_n2733), .C(_abc_42016_n4709), .Y(_abc_42016_n4724) );
  OAI21X1 OAI21X1_1278 ( .A(_abc_42016_n4564), .B(_abc_42016_n4569), .C(_abc_42016_n4731_1), .Y(_abc_42016_n4732) );
  OAI21X1 OAI21X1_1279 ( .A(_abc_42016_n4626), .B(_abc_42016_n4732), .C(_abc_42016_n4559), .Y(_abc_42016_n4733) );
  OAI21X1 OAI21X1_128 ( .A(_abc_42016_n1104_1), .B(_abc_42016_n1105), .C(_abc_42016_n1111_1), .Y(_abc_42016_n1112) );
  OAI21X1 OAI21X1_1280 ( .A(_abc_42016_n3475), .B(_abc_42016_n676), .C(ei), .Y(_abc_42016_n4735_1) );
  OAI21X1 OAI21X1_1281 ( .A(intr), .B(_abc_42016_n4736), .C(_abc_42016_n4737_1), .Y(_abc_42016_n4738) );
  OAI21X1 OAI21X1_1282 ( .A(_abc_42016_n2026), .B(_abc_42016_n4735_1), .C(_abc_42016_n4739), .Y(ei_FF_INPUT) );
  OAI21X1 OAI21X1_1283 ( .A(alu__abc_41682_n43), .B(alu__abc_41682_n34), .C(alu__abc_41682_n42), .Y(alu__abc_41682_n44) );
  OAI21X1 OAI21X1_1284 ( .A(alu__abc_41682_n56), .B(alu__abc_41682_n57), .C(alu__abc_41682_n47), .Y(alu__abc_41682_n58) );
  OAI21X1 OAI21X1_1285 ( .A(alu__abc_41682_n63), .B(alu__abc_41682_n55), .C(alu__abc_41682_n66), .Y(alu__abc_41682_n70) );
  OAI21X1 OAI21X1_1286 ( .A(alu__abc_41682_n82), .B(alu__abc_41682_n83), .C(alu__abc_41682_n88), .Y(alu__abc_41682_n89) );
  OAI21X1 OAI21X1_1287 ( .A(alu__abc_41682_n100), .B(alu__abc_41682_n102), .C(alu__abc_41682_n93), .Y(alu__abc_41682_n103) );
  OAI21X1 OAI21X1_1288 ( .A(alu__abc_41682_n122), .B(alu__abc_41682_n127), .C(alu__abc_41682_n49), .Y(alu__abc_41682_n128) );
  OAI21X1 OAI21X1_1289 ( .A(alu__abc_41682_n119), .B(alu__abc_41682_n129), .C(alu__abc_41682_n76), .Y(alu__abc_41682_n130) );
  OAI21X1 OAI21X1_129 ( .A(_abc_42016_n1024), .B(_abc_42016_n1068), .C(_abc_42016_n1069), .Y(_abc_42016_n1114_1) );
  OAI21X1 OAI21X1_1290 ( .A(alu__abc_41682_n132), .B(alu__abc_41682_n131), .C(alu__abc_41682_n108), .Y(alu__abc_41682_n133) );
  OAI21X1 OAI21X1_1291 ( .A(alu__abc_41682_n138), .B(alu__abc_41682_n141), .C(alu__abc_41682_n137), .Y(alu__abc_41682_n142) );
  OAI21X1 OAI21X1_1292 ( .A(alu__abc_41682_n116), .B(alu__abc_41682_n145), .C(alu__abc_41682_n90), .Y(alu__abc_41682_n146) );
  OAI21X1 OAI21X1_1293 ( .A(alu_sel_0_), .B(alu__abc_41682_n153), .C(alu_sel_1_), .Y(alu__abc_41682_n154) );
  OAI21X1 OAI21X1_1294 ( .A(alu__abc_41682_n104), .B(alu_sel_2_), .C(alu__abc_41682_n155), .Y(alu__abc_41682_n159) );
  OAI21X1 OAI21X1_1295 ( .A(alu__abc_41682_n38), .B(alu__abc_41682_n37), .C(alu_cin), .Y(alu__abc_41682_n161) );
  OAI21X1 OAI21X1_1296 ( .A(alu__abc_41682_n141), .B(alu__abc_41682_n164), .C(alu__abc_41682_n162), .Y(alu__abc_41682_n165) );
  OAI21X1 OAI21X1_1297 ( .A(alu__abc_41682_n122), .B(alu__abc_41682_n127), .C(alu__abc_41682_n52), .Y(alu__abc_41682_n168) );
  OAI21X1 OAI21X1_1298 ( .A(alu__abc_41682_n158), .B(alu__abc_41682_n172), .C(alu__abc_41682_n159), .Y(alu__abc_41682_n173) );
  OAI21X1 OAI21X1_1299 ( .A(alu_oprb_7_), .B(alu_opra_7_), .C(alu__abc_41682_n182), .Y(alu__abc_41682_n183) );
  OAI21X1 OAI21X1_13 ( .A(_abc_42016_n602), .B(_abc_42016_n587), .C(_abc_42016_n622), .Y(_abc_42016_n623) );
  OAI21X1 OAI21X1_130 ( .A(_abc_42016_n695), .B(_abc_42016_n709), .C(_abc_42016_n757), .Y(_abc_42016_n1121_1) );
  OAI21X1 OAI21X1_1300 ( .A(alu__abc_41682_n153), .B(alu__abc_41682_n98), .C(alu__abc_41682_n184), .Y(alu__abc_41682_n185) );
  OAI21X1 OAI21X1_1301 ( .A(alu__abc_41682_n108), .B(alu__abc_41682_n179), .C(alu__abc_41682_n186), .Y(alu__abc_41682_n187) );
  OAI21X1 OAI21X1_1302 ( .A(alu__abc_41682_n111), .B(alu__abc_41682_n110), .C(alu__abc_41682_n194), .Y(alu__abc_41682_n195) );
  OAI21X1 OAI21X1_1303 ( .A(alu__abc_41682_n81), .B(alu__abc_41682_n92), .C(alu__abc_41682_n199), .Y(alu__abc_41682_n200) );
  OAI21X1 OAI21X1_1304 ( .A(alu__abc_41682_n127), .B(alu__abc_41682_n205), .C(alu__abc_41682_n204), .Y(alu__abc_41682_n206) );
  OAI21X1 OAI21X1_1305 ( .A(alu__abc_41682_n122), .B(alu__abc_41682_n127), .C(alu__abc_41682_n169_1), .Y(alu__abc_41682_n208) );
  OAI21X1 OAI21X1_1306 ( .A(alu__abc_41682_n129), .B(alu__abc_41682_n201), .C(alu__abc_41682_n209), .Y(alu__abc_41682_n210) );
  OAI21X1 OAI21X1_1307 ( .A(alu__abc_41682_n84), .B(alu__abc_41682_n181), .C(alu__abc_41682_n220), .Y(alu__abc_41682_n221) );
  OAI21X1 OAI21X1_1308 ( .A(alu__abc_41682_n172), .B(alu__abc_41682_n230), .C(alu__abc_41682_n150), .Y(alu__abc_41682_n231) );
  OAI21X1 OAI21X1_1309 ( .A(alu__abc_41682_n54), .B(alu__abc_41682_n45_1), .C(alu__abc_41682_n169_1), .Y(alu__abc_41682_n235) );
  OAI21X1 OAI21X1_131 ( .A(_abc_42016_n1122), .B(_abc_42016_n1061), .C(_abc_42016_n671_1), .Y(_abc_42016_n1123) );
  OAI21X1 OAI21X1_1310 ( .A(alu__abc_41682_n153), .B(alu__abc_41682_n61), .C(alu__abc_41682_n184), .Y(alu__abc_41682_n241) );
  OAI21X1 OAI21X1_1311 ( .A(alu__abc_41682_n59), .B(alu__abc_41682_n181), .C(alu__abc_41682_n241), .Y(alu__abc_41682_n242) );
  OAI21X1 OAI21X1_1312 ( .A(alu__abc_41682_n159), .B(alu__abc_41682_n215), .C(alu__abc_41682_n243), .Y(alu__abc_41682_n244) );
  OAI21X1 OAI21X1_1313 ( .A(alu__abc_41682_n83), .B(alu__abc_41682_n247), .C(alu__abc_41682_n194), .Y(alu__abc_41682_n248) );
  OAI21X1 OAI21X1_1314 ( .A(alu__abc_41682_n83), .B(alu__abc_41682_n247), .C(alu__abc_41682_n238), .Y(alu__abc_41682_n249) );
  OAI21X1 OAI21X1_1315 ( .A(alu_oprb_5_), .B(alu_opra_5_), .C(alu__abc_41682_n182), .Y(alu__abc_41682_n252) );
  OAI21X1 OAI21X1_1316 ( .A(alu__abc_41682_n153), .B(alu__abc_41682_n82), .C(alu__abc_41682_n184), .Y(alu__abc_41682_n253) );
  OAI21X1 OAI21X1_1317 ( .A(alu__abc_41682_n76), .B(alu__abc_41682_n179), .C(alu__abc_41682_n254), .Y(alu__abc_41682_n255) );
  OAI21X1 OAI21X1_1318 ( .A(alu__abc_41682_n149), .B(alu__abc_41682_n63), .C(alu__abc_41682_n66), .Y(alu__abc_41682_n263) );
  OAI21X1 OAI21X1_1319 ( .A(alu__abc_41682_n265), .B(alu__abc_41682_n206), .C(alu__abc_41682_n266_1), .Y(alu__abc_41682_n267) );
  OAI21X1 OAI21X1_132 ( .A(_abc_42016_n757), .B(_abc_42016_n1062), .C(_abc_42016_n1127), .Y(_abc_42016_n1128) );
  OAI21X1 OAI21X1_1320 ( .A(alu__abc_41682_n261), .B(alu__abc_41682_n269), .C(alu__abc_41682_n270_1), .Y(alu__abc_41682_n271_1) );
  OAI21X1 OAI21X1_1321 ( .A(alu__abc_41682_n46_1), .B(alu__abc_41682_n45_1), .C(alu__abc_41682_n40), .Y(alu__abc_41682_n272) );
  OAI21X1 OAI21X1_1322 ( .A(alu__abc_41682_n274), .B(alu__abc_41682_n275_1), .C(alu__abc_41682_n272), .Y(alu__abc_41682_n276) );
  OAI21X1 OAI21X1_1323 ( .A(alu__abc_41682_n54), .B(alu__abc_41682_n179), .C(alu__abc_41682_n181), .Y(alu__abc_41682_n277_1) );
  OAI21X1 OAI21X1_1324 ( .A(alu_oprb_2_), .B(alu_opra_2_), .C(alu__abc_41682_n277_1), .Y(alu__abc_41682_n278) );
  OAI21X1 OAI21X1_1325 ( .A(alu__abc_41682_n161), .B(alu__abc_41682_n283), .C(alu__abc_41682_n279_1), .Y(alu__abc_41682_n284) );
  OAI21X1 OAI21X1_1326 ( .A(alu__abc_41682_n271_1), .B(alu__abc_41682_n268_1), .C(alu__abc_41682_n287), .Y(alu__abc_41682_n288) );
  OAI21X1 OAI21X1_1327 ( .A(alu__abc_41682_n204), .B(alu__abc_41682_n293), .C(alu__abc_41682_n150), .Y(alu__abc_41682_n294) );
  OAI21X1 OAI21X1_1328 ( .A(alu__abc_41682_n34), .B(alu__abc_41682_n181), .C(alu__abc_41682_n193), .Y(alu__abc_41682_n295) );
  OAI21X1 OAI21X1_1329 ( .A(alu__abc_41682_n42), .B(alu__abc_41682_n218), .C(alu__abc_41682_n296), .Y(alu__abc_41682_n297) );
  OAI21X1 OAI21X1_133 ( .A(_abc_42016_n1130), .B(_abc_42016_n1056), .C(_abc_42016_n994), .Y(_abc_42016_n1131) );
  OAI21X1 OAI21X1_1330 ( .A(alu__abc_41682_n193), .B(alu__abc_41682_n292), .C(alu__abc_41682_n302), .Y(alu__abc_41682_n303) );
  OAI21X1 OAI21X1_1331 ( .A(alu__abc_41682_n38), .B(alu__abc_41682_n181), .C(alu__abc_41682_n304), .Y(alu__abc_41682_n305) );
  OAI21X1 OAI21X1_1332 ( .A(alu_sel_1_), .B(alu_sel_0_), .C(alu_cin), .Y(alu__abc_41682_n306) );
  OAI21X1 OAI21X1_1333 ( .A(alu__abc_41682_n38), .B(alu__abc_41682_n37), .C(alu__abc_41682_n306), .Y(alu__abc_41682_n307) );
  OAI21X1 OAI21X1_1334 ( .A(alu__abc_41682_n104), .B(alu_sel_2_), .C(alu__abc_41682_n39), .Y(alu__abc_41682_n309) );
  OAI21X1 OAI21X1_1335 ( .A(alu__abc_41682_n180), .B(alu__abc_41682_n309), .C(alu__abc_41682_n308), .Y(alu__abc_41682_n310) );
  OAI21X1 OAI21X1_1336 ( .A(alu__abc_41682_n290), .B(alu__abc_41682_n289), .C(alu__abc_41682_n312), .Y(alu__abc_41682_n313) );
  OAI21X1 OAI21X1_1337 ( .A(alu__abc_41682_n258), .B(alu__abc_41682_n260), .C(alu__abc_41682_n318), .Y(alu__abc_41682_n319) );
  OAI21X1 OAI21X1_1338 ( .A(alu__abc_41682_n290), .B(alu__abc_41682_n289), .C(alu__abc_41682_n316), .Y(alu__abc_41682_n324) );
  OAI21X1 OAI21X1_1339 ( .A(alu__abc_41682_n258), .B(alu__abc_41682_n260), .C(alu__abc_41682_n325), .Y(alu__abc_41682_n331) );
  OAI21X1 OAI21X1_134 ( .A(_abc_42016_n1124), .B(_abc_42016_n1129), .C(_abc_42016_n1132), .Y(_abc_42016_n1133) );
  OAI21X1 OAI21X1_1340 ( .A(alu__abc_41682_n330), .B(alu__abc_41682_n329), .C(alu__abc_41682_n333), .Y(alu__abc_41682_n334) );
  OAI21X1 OAI21X1_1341 ( .A(alu__abc_41682_n121), .B(alu__abc_41682_n339), .C(alu__abc_41682_n342), .Y(alu_res_2_) );
  OAI21X1 OAI21X1_1342 ( .A(alu__abc_41682_n268_1), .B(alu__abc_41682_n271_1), .C(alu__abc_41682_n339), .Y(alu__abc_41682_n344) );
  OAI21X1 OAI21X1_1343 ( .A(alu__abc_41682_n48), .B(alu__abc_41682_n339), .C(alu__abc_41682_n344), .Y(alu_res_3_) );
  OAI21X1 OAI21X1_1344 ( .A(alu__abc_41682_n118), .B(alu__abc_41682_n339), .C(alu__abc_41682_n346), .Y(alu_res_4_) );
  OAI21X1 OAI21X1_1345 ( .A(alu__abc_41682_n86), .B(alu__abc_41682_n339), .C(alu__abc_41682_n349), .Y(alu_res_6_) );
  OAI21X1 OAI21X1_1346 ( .A(alu__abc_41682_n97), .B(alu__abc_41682_n339), .C(alu__abc_41682_n351), .Y(alu_res_7_) );
  OAI21X1 OAI21X1_1347 ( .A(alu_oprb_3_), .B(alu_opra_3_), .C(alu__abc_41682_n67), .Y(alu__abc_41682_n353) );
  OAI21X1 OAI21X1_1348 ( .A(alu_oprb_3_), .B(alu__abc_41682_n48), .C(alu__abc_41682_n128), .Y(alu__abc_41682_n354) );
  OAI21X1 OAI21X1_1349 ( .A(alu__abc_41682_n354), .B(alu__abc_41682_n154), .C(alu__abc_41682_n355), .Y(alu__abc_41682_n356) );
  OAI21X1 OAI21X1_135 ( .A(rdatahold2_2_), .B(_abc_42016_n1097), .C(_abc_42016_n1133), .Y(_abc_42016_n1134) );
  OAI21X1 OAI21X1_1350 ( .A(alu__abc_41682_n353), .B(alu__abc_41682_n269), .C(alu__abc_41682_n357), .Y(alu_auxcar) );
  OAI21X1 OAI21X1_1351 ( .A(alu__abc_41682_n363), .B(alu__abc_41682_n361), .C(alu__abc_41682_n155), .Y(alu__abc_41682_n364) );
  OAI21X1 OAI21X1_136 ( .A(_abc_42016_n556), .B(_abc_42016_n988), .C(regfil_5__3_), .Y(_abc_42016_n1136) );
  OAI21X1 OAI21X1_137 ( .A(_abc_42016_n1101_1), .B(_abc_42016_n1104_1), .C(_abc_42016_n1145), .Y(_abc_42016_n1146_1) );
  OAI21X1 OAI21X1_138 ( .A(_abc_42016_n611), .B(_abc_42016_n757), .C(_abc_42016_n1109), .Y(_abc_42016_n1152) );
  OAI21X1 OAI21X1_139 ( .A(_abc_42016_n757), .B(_abc_42016_n1159), .C(_abc_42016_n1117), .Y(_abc_42016_n1160) );
  OAI21X1 OAI21X1_14 ( .A(regfil_5__0_), .B(_abc_42016_n626), .C(opcode_2_), .Y(_abc_42016_n627) );
  OAI21X1 OAI21X1_140 ( .A(_abc_42016_n1165), .B(_abc_42016_n1166), .C(_abc_42016_n1023), .Y(_abc_42016_n1167) );
  OAI21X1 OAI21X1_141 ( .A(_abc_42016_n1170), .B(_abc_42016_n1172_1), .C(_abc_42016_n1171_1), .Y(_abc_42016_n1173) );
  OAI21X1 OAI21X1_142 ( .A(_abc_42016_n1173), .B(_abc_42016_n1169), .C(_abc_42016_n1175), .Y(_abc_42016_n1176) );
  OAI21X1 OAI21X1_143 ( .A(regfil_3__4_), .B(_abc_42016_n993), .C(_abc_42016_n995), .Y(_abc_42016_n1181) );
  OAI21X1 OAI21X1_144 ( .A(regfil_5__3_), .B(_abc_42016_n1126), .C(regfil_5__4_), .Y(_abc_42016_n1182) );
  OAI21X1 OAI21X1_145 ( .A(_abc_42016_n1139), .B(_abc_42016_n1120), .C(_abc_42016_n843), .Y(_abc_42016_n1189) );
  OAI21X1 OAI21X1_146 ( .A(_abc_42016_n1190), .B(_abc_42016_n1187), .C(_abc_42016_n1170), .Y(_abc_42016_n1191) );
  OAI21X1 OAI21X1_147 ( .A(regfil_1__3_), .B(regfil_5__3_), .C(_abc_42016_n1196_1), .Y(_abc_42016_n1199_1) );
  OAI21X1 OAI21X1_148 ( .A(_abc_42016_n1149_1), .B(_abc_42016_n1148), .C(_abc_42016_n1143), .Y(_abc_42016_n1202) );
  OAI21X1 OAI21X1_149 ( .A(regfil_5__3_), .B(sp_3_), .C(_abc_42016_n1214), .Y(_abc_42016_n1215) );
  OAI21X1 OAI21X1_15 ( .A(regfil_6__0_), .B(_abc_42016_n539), .C(_abc_42016_n631), .Y(_abc_42016_n632) );
  OAI21X1 OAI21X1_150 ( .A(_abc_42016_n1186), .B(_abc_42016_n1218), .C(_abc_42016_n1181), .Y(_abc_42016_n1219) );
  OAI21X1 OAI21X1_151 ( .A(_abc_42016_n1055), .B(_abc_42016_n1221_1), .C(_abc_42016_n1220), .Y(_abc_36783_n3447) );
  OAI21X1 OAI21X1_152 ( .A(rdatahold2_5_), .B(_abc_42016_n993), .C(_abc_42016_n1057), .Y(_abc_42016_n1224_1) );
  OAI21X1 OAI21X1_153 ( .A(_abc_42016_n1226), .B(_abc_42016_n1227), .C(_abc_42016_n1170), .Y(_abc_42016_n1228) );
  OAI21X1 OAI21X1_154 ( .A(_abc_42016_n562), .B(_abc_42016_n1246), .C(_abc_42016_n1045), .Y(_abc_42016_n1247_1) );
  OAI21X1 OAI21X1_155 ( .A(_abc_42016_n872), .B(_abc_42016_n1252), .C(_abc_42016_n1125), .Y(_abc_42016_n1253) );
  OAI21X1 OAI21X1_156 ( .A(_abc_42016_n1251), .B(_abc_42016_n1253), .C(_abc_42016_n1050), .Y(_abc_42016_n1254) );
  OAI21X1 OAI21X1_157 ( .A(_abc_42016_n1254), .B(_abc_42016_n1250_1), .C(_abc_42016_n1224_1), .Y(_abc_42016_n1255) );
  OAI21X1 OAI21X1_158 ( .A(_abc_42016_n1055), .B(_abc_42016_n1257), .C(_abc_42016_n1256), .Y(_abc_36783_n3450) );
  OAI21X1 OAI21X1_159 ( .A(_abc_42016_n923), .B(_abc_42016_n989), .C(_abc_42016_n1020), .Y(_abc_42016_n1260) );
  OAI21X1 OAI21X1_16 ( .A(regfil_1__0_), .B(_abc_42016_n626), .C(_abc_42016_n536), .Y(_abc_42016_n633) );
  OAI21X1 OAI21X1_160 ( .A(_abc_42016_n1019), .B(_abc_42016_n993), .C(_abc_42016_n1261), .Y(_abc_42016_n1262) );
  OAI21X1 OAI21X1_161 ( .A(_abc_42016_n1260), .B(_abc_42016_n1259), .C(_abc_42016_n1262), .Y(_abc_42016_n1263) );
  OAI21X1 OAI21X1_162 ( .A(_abc_42016_n1264), .B(_abc_42016_n1237), .C(_abc_42016_n1265), .Y(_abc_42016_n1266) );
  OAI21X1 OAI21X1_163 ( .A(_abc_42016_n642), .B(_abc_42016_n872), .C(_abc_42016_n1238), .Y(_abc_42016_n1267) );
  OAI21X1 OAI21X1_164 ( .A(_abc_42016_n1272_1), .B(_abc_42016_n1273), .C(_abc_42016_n1274_1), .Y(_abc_42016_n1275) );
  OAI21X1 OAI21X1_165 ( .A(_abc_42016_n1005), .B(_abc_42016_n1276), .C(_abc_42016_n561), .Y(_abc_42016_n1277) );
  OAI21X1 OAI21X1_166 ( .A(_abc_42016_n872), .B(_abc_42016_n1279), .C(_abc_42016_n1234), .Y(_abc_42016_n1280) );
  OAI21X1 OAI21X1_167 ( .A(_abc_42016_n1283), .B(_abc_42016_n1233), .C(_abc_42016_n1281), .Y(_abc_42016_n1284) );
  OAI21X1 OAI21X1_168 ( .A(_abc_42016_n1285), .B(_abc_42016_n1282), .C(_abc_42016_n1023), .Y(_abc_42016_n1286) );
  OAI21X1 OAI21X1_169 ( .A(_abc_42016_n1289), .B(_abc_42016_n1291), .C(_abc_42016_n1170), .Y(_abc_42016_n1292) );
  OAI21X1 OAI21X1_17 ( .A(regfil_2__0_), .B(_abc_42016_n539), .C(_abc_42016_n635), .Y(_abc_42016_n636) );
  OAI21X1 OAI21X1_170 ( .A(regfil_5__5_), .B(_abc_42016_n1184), .C(regfil_5__6_), .Y(_abc_42016_n1294) );
  OAI21X1 OAI21X1_171 ( .A(_abc_42016_n1292), .B(_abc_42016_n1288), .C(_abc_42016_n1298), .Y(_abc_42016_n1299_1) );
  OAI21X1 OAI21X1_172 ( .A(_abc_42016_n959), .B(_abc_42016_n989), .C(_abc_42016_n1011), .Y(_abc_42016_n1304) );
  OAI21X1 OAI21X1_173 ( .A(_abc_42016_n1309), .B(_abc_42016_n1311), .C(_abc_42016_n1036), .Y(_abc_42016_n1312) );
  OAI21X1 OAI21X1_174 ( .A(_abc_42016_n1270), .B(_abc_42016_n1271_1), .C(_abc_42016_n1273), .Y(_abc_42016_n1314) );
  OAI21X1 OAI21X1_175 ( .A(_abc_42016_n562), .B(_abc_42016_n1320), .C(_abc_42016_n1045), .Y(_abc_42016_n1321_1) );
  OAI21X1 OAI21X1_176 ( .A(_abc_42016_n923), .B(_abc_42016_n1323), .C(_abc_42016_n1284), .Y(_abc_42016_n1324) );
  OAI21X1 OAI21X1_177 ( .A(_abc_42016_n1335_1), .B(_abc_42016_n1334), .C(_abc_42016_n1125), .Y(_abc_42016_n1336) );
  OAI21X1 OAI21X1_178 ( .A(_abc_42016_n1348), .B(_abc_42016_n562), .C(_abc_42016_n1345), .Y(_abc_42016_n1349) );
  OAI21X1 OAI21X1_179 ( .A(pc_1_), .B(pc_0_), .C(pc_2_), .Y(_abc_42016_n1358) );
  OAI21X1 OAI21X1_18 ( .A(_abc_42016_n602), .B(_abc_42016_n527), .C(_abc_42016_n638), .Y(_abc_42016_n639) );
  OAI21X1 OAI21X1_180 ( .A(_abc_42016_n1354), .B(_abc_42016_n1364), .C(_abc_42016_n1353), .Y(_abc_42016_n1365) );
  OAI21X1 OAI21X1_181 ( .A(_abc_42016_n536), .B(_abc_42016_n727), .C(_abc_42016_n1374), .Y(_abc_42016_n1377) );
  OAI21X1 OAI21X1_182 ( .A(_abc_42016_n1375), .B(_abc_42016_n1376), .C(_abc_42016_n1377), .Y(_abc_42016_n1378) );
  OAI21X1 OAI21X1_183 ( .A(_abc_42016_n1353), .B(_abc_42016_n1374), .C(_abc_42016_n1378), .Y(_abc_42016_n1379) );
  OAI21X1 OAI21X1_184 ( .A(_abc_42016_n1381), .B(_abc_42016_n1389), .C(_abc_42016_n1353), .Y(_abc_42016_n1390) );
  OAI21X1 OAI21X1_185 ( .A(_abc_42016_n1381), .B(_abc_42016_n1392), .C(_abc_42016_n1390), .Y(_abc_42016_n1393) );
  OAI21X1 OAI21X1_186 ( .A(_abc_42016_n1353), .B(_abc_42016_n1405), .C(_abc_42016_n1403), .Y(_abc_42016_n1406) );
  OAI21X1 OAI21X1_187 ( .A(_abc_42016_n1398), .B(_abc_42016_n626), .C(_abc_42016_n1380), .Y(_abc_42016_n1407) );
  OAI21X1 OAI21X1_188 ( .A(_abc_42016_n669), .B(_abc_42016_n682), .C(_abc_42016_n1408), .Y(_abc_42016_n1409) );
  OAI21X1 OAI21X1_189 ( .A(_abc_42016_n573), .B(_abc_42016_n1399), .C(_abc_42016_n668), .Y(_abc_42016_n1412) );
  OAI21X1 OAI21X1_19 ( .A(_abc_42016_n641), .B(_abc_42016_n651_1), .C(_abc_42016_n608), .Y(_abc_42016_n652) );
  OAI21X1 OAI21X1_190 ( .A(_abc_42016_n629), .B(_abc_42016_n1412), .C(_abc_42016_n1411), .Y(_abc_42016_n1413) );
  OAI21X1 OAI21X1_191 ( .A(_abc_42016_n1380), .B(_abc_42016_n1393), .C(_abc_42016_n1414), .Y(_abc_42016_n1415) );
  OAI21X1 OAI21X1_192 ( .A(wdatahold2_0_), .B(_abc_42016_n1411), .C(_abc_42016_n677), .Y(_abc_42016_n1417) );
  OAI21X1 OAI21X1_193 ( .A(_abc_42016_n1417), .B(_abc_42016_n1416), .C(_abc_42016_n1352), .Y(wdatahold2_0__FF_INPUT) );
  OAI21X1 OAI21X1_194 ( .A(_abc_42016_n669), .B(_abc_42016_n1347), .C(wdatahold2_1_), .Y(_abc_42016_n1420) );
  OAI21X1 OAI21X1_195 ( .A(_abc_42016_n722), .B(_abc_42016_n1350), .C(_abc_42016_n1420), .Y(_abc_42016_n1421) );
  OAI21X1 OAI21X1_196 ( .A(_abc_42016_n1381), .B(_abc_42016_n1392), .C(_abc_42016_n1422), .Y(_abc_42016_n1423) );
  OAI21X1 OAI21X1_197 ( .A(_abc_42016_n1381), .B(_abc_42016_n1424), .C(_abc_42016_n1423), .Y(_abc_42016_n1425) );
  OAI21X1 OAI21X1_198 ( .A(_abc_42016_n1427), .B(_abc_42016_n1004), .C(_abc_42016_n1428), .Y(_abc_42016_n1429) );
  OAI21X1 OAI21X1_199 ( .A(_abc_42016_n1422), .B(_abc_42016_n1405), .C(_abc_42016_n1430), .Y(_abc_42016_n1431) );
  OAI21X1 OAI21X1_2 ( .A(_abc_42016_n530), .B(_abc_42016_n533), .C(_abc_42016_n529), .Y(_abc_42016_n534_1) );
  OAI21X1 OAI21X1_20 ( .A(_abc_42016_n588_1), .B(_abc_42016_n640), .C(_abc_42016_n661_1), .Y(_abc_42016_n662) );
  OAI21X1 OAI21X1_200 ( .A(_abc_42016_n1380), .B(_abc_42016_n1425), .C(_abc_42016_n1432), .Y(_abc_42016_n1433) );
  OAI21X1 OAI21X1_201 ( .A(_abc_42016_n1353), .B(_abc_42016_n1366), .C(_abc_42016_n1422), .Y(_abc_42016_n1434) );
  OAI21X1 OAI21X1_202 ( .A(_abc_42016_n1436), .B(_abc_42016_n1439_1), .C(_abc_42016_n1411), .Y(_abc_42016_n1440) );
  OAI21X1 OAI21X1_203 ( .A(_abc_42016_n669), .B(_abc_42016_n1347), .C(wdatahold2_2_), .Y(_abc_42016_n1447) );
  OAI21X1 OAI21X1_204 ( .A(_abc_42016_n1446), .B(_abc_42016_n1350), .C(_abc_42016_n1447), .Y(_abc_42016_n1448) );
  OAI21X1 OAI21X1_205 ( .A(_abc_42016_n1422), .B(_abc_42016_n1368), .C(_abc_42016_n1449), .Y(_abc_42016_n1450) );
  OAI21X1 OAI21X1_206 ( .A(_abc_42016_n1366), .B(_abc_42016_n1451), .C(_abc_42016_n1450), .Y(_abc_42016_n1452) );
  OAI21X1 OAI21X1_207 ( .A(opcode_4_), .B(regfil_0__2_), .C(_abc_42016_n1455), .Y(_abc_42016_n1456) );
  OAI21X1 OAI21X1_208 ( .A(_abc_42016_n1449), .B(_abc_42016_n1405), .C(_abc_42016_n1458), .Y(_abc_42016_n1459) );
  OAI21X1 OAI21X1_209 ( .A(_abc_42016_n1462), .B(_abc_42016_n1463), .C(_abc_42016_n1467), .Y(_abc_42016_n1468) );
  OAI21X1 OAI21X1_21 ( .A(_abc_42016_n681), .B(_abc_42016_n683), .C(_abc_42016_n561), .Y(_abc_42016_n684) );
  OAI21X1 OAI21X1_210 ( .A(_abc_42016_n1452), .B(_abc_42016_n1453), .C(_abc_42016_n1469), .Y(_abc_42016_n1470) );
  OAI21X1 OAI21X1_211 ( .A(_abc_42016_n669), .B(_abc_42016_n1347), .C(wdatahold2_3_), .Y(_abc_42016_n1475) );
  OAI21X1 OAI21X1_212 ( .A(_abc_42016_n800), .B(_abc_42016_n1350), .C(_abc_42016_n1475), .Y(_abc_42016_n1476) );
  OAI21X1 OAI21X1_213 ( .A(_abc_42016_n1381), .B(_abc_42016_n1478), .C(_abc_42016_n1477), .Y(_abc_42016_n1479) );
  OAI21X1 OAI21X1_214 ( .A(_abc_42016_n1381), .B(_abc_42016_n1480), .C(_abc_42016_n1479), .Y(_abc_42016_n1481) );
  OAI21X1 OAI21X1_215 ( .A(_abc_42016_n1451), .B(_abc_42016_n1366), .C(_abc_42016_n1477), .Y(_abc_42016_n1482) );
  OAI21X1 OAI21X1_216 ( .A(_abc_42016_n1374), .B(_abc_42016_n1483), .C(_abc_42016_n1378), .Y(_abc_42016_n1487) );
  OAI21X1 OAI21X1_217 ( .A(_abc_42016_n1488), .B(_abc_42016_n1004), .C(_abc_42016_n1489), .Y(_abc_42016_n1490) );
  OAI21X1 OAI21X1_218 ( .A(_abc_42016_n800), .B(_abc_42016_n1412), .C(_abc_42016_n1491), .Y(_abc_42016_n1492) );
  OAI21X1 OAI21X1_219 ( .A(_abc_42016_n1477), .B(_abc_42016_n1405), .C(_abc_42016_n1493), .Y(_abc_42016_n1494) );
  OAI21X1 OAI21X1_22 ( .A(_abc_42016_n671_1), .B(_abc_42016_n678), .C(_abc_42016_n684), .Y(_abc_42016_n685) );
  OAI21X1 OAI21X1_220 ( .A(_abc_42016_n1380), .B(_abc_42016_n1481), .C(_abc_42016_n1495), .Y(_abc_42016_n1496_1) );
  OAI21X1 OAI21X1_221 ( .A(_abc_42016_n669), .B(_abc_42016_n1347), .C(wdatahold2_4_), .Y(_abc_42016_n1501) );
  OAI21X1 OAI21X1_222 ( .A(_abc_42016_n842), .B(_abc_42016_n1350), .C(_abc_42016_n1501), .Y(_abc_42016_n1502) );
  OAI21X1 OAI21X1_223 ( .A(_abc_42016_n1381), .B(_abc_42016_n1480), .C(_abc_42016_n1503), .Y(_abc_42016_n1509) );
  OAI21X1 OAI21X1_224 ( .A(_abc_42016_n1381), .B(_abc_42016_n1511), .C(_abc_42016_n1509), .Y(_abc_42016_n1512) );
  OAI21X1 OAI21X1_225 ( .A(opcode_4_), .B(regfil_0__4_), .C(_abc_42016_n1514), .Y(_abc_42016_n1515) );
  OAI21X1 OAI21X1_226 ( .A(_abc_42016_n1503), .B(_abc_42016_n1405), .C(_abc_42016_n1517), .Y(_abc_42016_n1518) );
  OAI21X1 OAI21X1_227 ( .A(_abc_42016_n842), .B(_abc_42016_n1412), .C(_abc_42016_n1411), .Y(_abc_42016_n1519) );
  OAI21X1 OAI21X1_228 ( .A(_abc_42016_n1504), .B(_abc_42016_n1507), .C(_abc_42016_n1521), .Y(_abc_42016_n1522_1) );
  OAI21X1 OAI21X1_229 ( .A(_abc_42016_n669), .B(_abc_42016_n1347), .C(wdatahold2_5_), .Y(_abc_42016_n1528) );
  OAI21X1 OAI21X1_23 ( .A(_abc_42016_n513), .B(_abc_42016_n667), .C(_abc_42016_n690), .Y(_abc_42016_n691) );
  OAI21X1 OAI21X1_230 ( .A(_abc_42016_n1527), .B(_abc_42016_n1350), .C(_abc_42016_n1528), .Y(_abc_42016_n1529) );
  OAI21X1 OAI21X1_231 ( .A(_abc_42016_n1381), .B(_abc_42016_n1511), .C(_abc_42016_n1530), .Y(_abc_42016_n1531) );
  OAI21X1 OAI21X1_232 ( .A(_abc_42016_n1381), .B(_abc_42016_n1532), .C(_abc_42016_n1531), .Y(_abc_42016_n1533) );
  OAI21X1 OAI21X1_233 ( .A(opcode_4_), .B(regfil_0__5_), .C(_abc_42016_n1534), .Y(_abc_42016_n1535) );
  OAI21X1 OAI21X1_234 ( .A(_abc_42016_n898), .B(_abc_42016_n1004), .C(_abc_42016_n1537), .Y(_abc_42016_n1538) );
  OAI21X1 OAI21X1_235 ( .A(_abc_42016_n1530), .B(_abc_42016_n1405), .C(_abc_42016_n1539), .Y(_abc_42016_n1540) );
  OAI21X1 OAI21X1_236 ( .A(_abc_42016_n1503), .B(_abc_42016_n1484), .C(_abc_42016_n1530), .Y(_abc_42016_n1542) );
  OAI21X1 OAI21X1_237 ( .A(_abc_42016_n1530), .B(_abc_42016_n1374), .C(_abc_42016_n1378), .Y(_abc_42016_n1547) );
  OAI21X1 OAI21X1_238 ( .A(_abc_42016_n1380), .B(_abc_42016_n1533), .C(_abc_42016_n1548), .Y(_abc_42016_n1549) );
  OAI21X1 OAI21X1_239 ( .A(_abc_42016_n669), .B(_abc_42016_n1347), .C(wdatahold2_6_), .Y(_abc_42016_n1555) );
  OAI21X1 OAI21X1_24 ( .A(regfil_3__0_), .B(_abc_42016_n600), .C(_abc_42016_n692), .Y(_abc_42016_n693) );
  OAI21X1 OAI21X1_240 ( .A(_abc_42016_n1554), .B(_abc_42016_n1350), .C(_abc_42016_n1555), .Y(_abc_42016_n1556) );
  OAI21X1 OAI21X1_241 ( .A(_abc_42016_n1530), .B(_abc_42016_n1511), .C(_abc_42016_n1557), .Y(_abc_42016_n1558) );
  OAI21X1 OAI21X1_242 ( .A(pc_0_), .B(pc_14_), .C(_abc_42016_n1558), .Y(_abc_42016_n1559) );
  OAI21X1 OAI21X1_243 ( .A(pc_14_), .B(_abc_42016_n1567), .C(_abc_42016_n1438), .Y(_abc_42016_n1568) );
  OAI21X1 OAI21X1_244 ( .A(_abc_42016_n1557), .B(_abc_42016_n1374), .C(_abc_42016_n1568), .Y(_abc_42016_n1569) );
  OAI21X1 OAI21X1_245 ( .A(_abc_42016_n1375), .B(_abc_42016_n1374), .C(_abc_42016_n1570), .Y(_abc_42016_n1571) );
  OAI21X1 OAI21X1_246 ( .A(opcode_4_), .B(regfil_0__6_), .C(_abc_42016_n1572), .Y(_abc_42016_n1573) );
  OAI21X1 OAI21X1_247 ( .A(_abc_42016_n1400), .B(_abc_42016_n1575), .C(_abc_42016_n1576), .Y(_abc_42016_n1577) );
  OAI21X1 OAI21X1_248 ( .A(_abc_42016_n1380), .B(_abc_42016_n1564), .C(_abc_42016_n1578_1), .Y(_abc_42016_n1579) );
  OAI21X1 OAI21X1_249 ( .A(opcode_4_), .B(_abc_42016_n954), .C(_abc_42016_n1592_1), .Y(_abc_42016_n1593) );
  OAI21X1 OAI21X1_25 ( .A(_abc_42016_n513), .B(_abc_42016_n667), .C(_abc_42016_n688), .Y(_abc_42016_n694) );
  OAI21X1 OAI21X1_250 ( .A(_abc_42016_n960), .B(_abc_42016_n1004), .C(_abc_42016_n1594_1), .Y(_abc_42016_n1595) );
  OAI21X1 OAI21X1_251 ( .A(_abc_42016_n1584_1), .B(_abc_42016_n1405), .C(_abc_42016_n1596_1), .Y(_abc_42016_n1597) );
  OAI21X1 OAI21X1_252 ( .A(_abc_42016_n1591), .B(_abc_42016_n1590_1), .C(_abc_42016_n1598), .Y(_abc_42016_n1599_1) );
  OAI21X1 OAI21X1_253 ( .A(wdatahold2_7_), .B(_abc_42016_n1411), .C(_abc_42016_n677), .Y(_abc_42016_n1601_1) );
  OAI21X1 OAI21X1_254 ( .A(_abc_42016_n1601_1), .B(_abc_42016_n1600_1), .C(_abc_42016_n1583), .Y(wdatahold2_7__FF_INPUT) );
  OAI21X1 OAI21X1_255 ( .A(_abc_42016_n588_1), .B(_abc_42016_n596), .C(_abc_42016_n593), .Y(_abc_42016_n1605_1) );
  OAI21X1 OAI21X1_256 ( .A(_abc_42016_n623), .B(_abc_42016_n662), .C(_abc_42016_n1606_1), .Y(_abc_42016_n1607_1) );
  OAI21X1 OAI21X1_257 ( .A(_abc_42016_n608), .B(_abc_42016_n1606_1), .C(_abc_42016_n1607_1), .Y(_abc_36783_n3520) );
  OAI21X1 OAI21X1_258 ( .A(_abc_42016_n714), .B(_abc_42016_n737), .C(_abc_42016_n1606_1), .Y(_abc_42016_n1609) );
  OAI21X1 OAI21X1_259 ( .A(_abc_42016_n712), .B(_abc_42016_n1606_1), .C(_abc_42016_n1609), .Y(_abc_36783_n3523) );
  OAI21X1 OAI21X1_26 ( .A(_abc_42016_n693), .B(_abc_42016_n665_1), .C(_abc_42016_n699), .Y(_abc_36783_n3361) );
  OAI21X1 OAI21X1_260 ( .A(_abc_42016_n743), .B(_abc_42016_n1606_1), .C(_abc_42016_n1611), .Y(_abc_36783_n3526) );
  OAI21X1 OAI21X1_261 ( .A(_abc_42016_n810_1), .B(_abc_42016_n817), .C(_abc_42016_n1606_1), .Y(_abc_42016_n1613) );
  OAI21X1 OAI21X1_262 ( .A(_abc_42016_n812), .B(_abc_42016_n1606_1), .C(_abc_42016_n1613), .Y(_abc_36783_n3529) );
  OAI21X1 OAI21X1_263 ( .A(_abc_42016_n834), .B(_abc_42016_n1606_1), .C(_abc_42016_n1615), .Y(_abc_36783_n3532) );
  OAI21X1 OAI21X1_264 ( .A(_abc_42016_n893), .B(_abc_42016_n1606_1), .C(_abc_42016_n1617), .Y(_abc_36783_n3535) );
  OAI21X1 OAI21X1_265 ( .A(_abc_42016_n913), .B(_abc_42016_n1606_1), .C(_abc_42016_n1619), .Y(_abc_36783_n3538) );
  OAI21X1 OAI21X1_266 ( .A(_abc_42016_n951), .B(_abc_42016_n970), .C(_abc_42016_n1606_1), .Y(_abc_42016_n1621) );
  OAI21X1 OAI21X1_267 ( .A(_abc_42016_n954), .B(_abc_42016_n1606_1), .C(_abc_42016_n1621), .Y(_abc_36783_n3541) );
  OAI21X1 OAI21X1_268 ( .A(_abc_42016_n556), .B(_abc_42016_n1605_1), .C(_abc_42016_n644), .Y(_abc_42016_n1625) );
  OAI21X1 OAI21X1_269 ( .A(_abc_42016_n664_1), .B(_abc_42016_n1624), .C(_abc_42016_n1625), .Y(_abc_42016_n1626) );
  OAI21X1 OAI21X1_27 ( .A(_abc_42016_n702_1), .B(_abc_42016_n704), .C(_abc_42016_n681), .Y(_abc_42016_n705) );
  OAI21X1 OAI21X1_270 ( .A(regfil_2__0_), .B(_abc_42016_n980), .C(_abc_42016_n1629_1), .Y(_abc_42016_n1630_1) );
  OAI21X1 OAI21X1_271 ( .A(_abc_42016_n1633), .B(_abc_42016_n1632), .C(_abc_42016_n779), .Y(_abc_42016_n1634) );
  OAI21X1 OAI21X1_272 ( .A(_abc_42016_n605_1), .B(_abc_42016_n657), .C(_abc_42016_n561), .Y(_abc_42016_n1638_1) );
  OAI21X1 OAI21X1_273 ( .A(_abc_42016_n1639_1), .B(_abc_42016_n689), .C(rdatahold_0_), .Y(_abc_42016_n1640) );
  OAI21X1 OAI21X1_274 ( .A(regfil_1__0_), .B(_abc_42016_n1638_1), .C(_abc_42016_n1640), .Y(_abc_42016_n1641) );
  OAI21X1 OAI21X1_275 ( .A(_abc_42016_n556), .B(_abc_42016_n1605_1), .C(_abc_42016_n645), .Y(_abc_42016_n1645) );
  OAI21X1 OAI21X1_276 ( .A(_abc_42016_n1624), .B(_abc_42016_n739), .C(_abc_42016_n1645), .Y(_abc_42016_n1646) );
  OAI21X1 OAI21X1_277 ( .A(regfil_2__1_), .B(_abc_42016_n1628), .C(_abc_42016_n1648), .Y(_abc_42016_n1649_1) );
  OAI21X1 OAI21X1_278 ( .A(_abc_42016_n1650), .B(_abc_42016_n1652_1), .C(_abc_42016_n779), .Y(_abc_42016_n1653) );
  OAI21X1 OAI21X1_279 ( .A(_abc_42016_n659_1), .B(_abc_42016_n1657), .C(_abc_42016_n1659), .Y(_abc_42016_n1660) );
  OAI21X1 OAI21X1_28 ( .A(_abc_42016_n680), .B(_abc_42016_n603), .C(_abc_42016_n706), .Y(_abc_42016_n707_1) );
  OAI21X1 OAI21X1_280 ( .A(_abc_42016_n1655), .B(_abc_42016_n1660), .C(_abc_42016_n588_1), .Y(_abc_42016_n1661) );
  OAI21X1 OAI21X1_281 ( .A(_abc_42016_n588_1), .B(_abc_42016_n1646), .C(_abc_42016_n1661), .Y(_abc_36783_n3557) );
  OAI21X1 OAI21X1_282 ( .A(_abc_42016_n611), .B(_abc_42016_n1623), .C(_abc_42016_n1663), .Y(_abc_42016_n1664_1) );
  OAI21X1 OAI21X1_283 ( .A(regfil_2__2_), .B(_abc_42016_n1647_1), .C(_abc_42016_n1668), .Y(_abc_42016_n1669) );
  OAI21X1 OAI21X1_284 ( .A(_abc_42016_n1672), .B(_abc_42016_n1671), .C(_abc_42016_n779), .Y(_abc_42016_n1673_1) );
  OAI21X1 OAI21X1_285 ( .A(_abc_42016_n644), .B(_abc_42016_n645), .C(_abc_42016_n611), .Y(_abc_42016_n1677) );
  OAI21X1 OAI21X1_286 ( .A(_abc_42016_n579), .B(_abc_42016_n586), .C(rdatahold2_2_), .Y(_abc_42016_n1679) );
  OAI21X1 OAI21X1_287 ( .A(regfil_1__0_), .B(regfil_1__1_), .C(regfil_1__2_), .Y(_abc_42016_n1680) );
  OAI21X1 OAI21X1_288 ( .A(_abc_42016_n720), .B(_abc_42016_n1684), .C(_abc_42016_n1665), .Y(_abc_36783_n3560) );
  OAI21X1 OAI21X1_289 ( .A(_abc_42016_n556), .B(_abc_42016_n1605_1), .C(_abc_42016_n643_1), .Y(_abc_42016_n1686) );
  OAI21X1 OAI21X1_29 ( .A(_abc_42016_n709), .B(_abc_42016_n697), .C(_abc_42016_n701), .Y(_abc_42016_n710) );
  OAI21X1 OAI21X1_290 ( .A(_abc_42016_n1624), .B(_abc_42016_n819), .C(_abc_42016_n1686), .Y(_abc_42016_n1687) );
  OAI21X1 OAI21X1_291 ( .A(_abc_42016_n796), .B(_abc_42016_n1666), .C(_abc_42016_n822), .Y(_abc_42016_n1698_1) );
  OAI21X1 OAI21X1_292 ( .A(regfil_2__2_), .B(_abc_42016_n1651), .C(regfil_2__3_), .Y(_abc_42016_n1699) );
  OAI21X1 OAI21X1_293 ( .A(_abc_42016_n1697_1), .B(_abc_42016_n1698_1), .C(_abc_42016_n1702), .Y(_abc_42016_n1703) );
  OAI21X1 OAI21X1_294 ( .A(_abc_42016_n1696), .B(_abc_42016_n1703), .C(_abc_42016_n588_1), .Y(_abc_42016_n1704) );
  OAI21X1 OAI21X1_295 ( .A(_abc_42016_n588_1), .B(_abc_42016_n1687), .C(_abc_42016_n1704), .Y(_abc_36783_n3563) );
  OAI21X1 OAI21X1_296 ( .A(_abc_42016_n610), .B(_abc_42016_n1623), .C(_abc_42016_n1706_1), .Y(_abc_42016_n1707) );
  OAI21X1 OAI21X1_297 ( .A(_abc_42016_n643_1), .B(_abc_42016_n647), .C(_abc_42016_n610), .Y(_abc_42016_n1709) );
  OAI21X1 OAI21X1_298 ( .A(regfil_2__4_), .B(_abc_42016_n1711), .C(_abc_42016_n1712), .Y(_abc_42016_n1713_1) );
  OAI21X1 OAI21X1_299 ( .A(_abc_42016_n1714_1), .B(_abc_42016_n1715), .C(_abc_42016_n779), .Y(_abc_42016_n1716) );
  OAI21X1 OAI21X1_3 ( .A(_abc_42016_n536), .B(_abc_42016_n539), .C(_abc_42016_n541), .Y(_abc_42016_n542) );
  OAI21X1 OAI21X1_30 ( .A(_abc_42016_n712), .B(_abc_42016_n655_1), .C(_abc_42016_n660), .Y(_abc_42016_n713) );
  OAI21X1 OAI21X1_300 ( .A(rdatahold_4_), .B(_abc_42016_n688), .C(_abc_42016_n1718), .Y(_abc_42016_n1719) );
  OAI21X1 OAI21X1_301 ( .A(_abc_42016_n579), .B(_abc_42016_n586), .C(rdatahold2_4_), .Y(_abc_42016_n1720) );
  OAI21X1 OAI21X1_302 ( .A(regfil_1__3_), .B(_abc_42016_n613), .C(regfil_1__4_), .Y(_abc_42016_n1721_1) );
  OAI21X1 OAI21X1_303 ( .A(_abc_42016_n720), .B(_abc_42016_n1725), .C(_abc_42016_n1708), .Y(_abc_36783_n3566) );
  OAI21X1 OAI21X1_304 ( .A(_abc_42016_n1624), .B(_abc_42016_n909), .C(_abc_42016_n1727), .Y(_abc_42016_n1728) );
  OAI21X1 OAI21X1_305 ( .A(_abc_42016_n610), .B(_abc_42016_n648_1), .C(_abc_42016_n642), .Y(_abc_42016_n1730) );
  OAI21X1 OAI21X1_306 ( .A(_abc_42016_n1732_1), .B(_abc_42016_n1734), .C(_abc_42016_n779), .Y(_abc_42016_n1735) );
  OAI21X1 OAI21X1_307 ( .A(rdatahold_5_), .B(_abc_42016_n688), .C(_abc_42016_n1741), .Y(_abc_42016_n1742) );
  OAI21X1 OAI21X1_308 ( .A(_abc_42016_n579), .B(_abc_42016_n586), .C(rdatahold2_5_), .Y(_abc_42016_n1743) );
  OAI21X1 OAI21X1_309 ( .A(_abc_42016_n720), .B(_abc_42016_n1747), .C(_abc_42016_n1728), .Y(_abc_36783_n3569) );
  OAI21X1 OAI21X1_31 ( .A(regfil_7__1_), .B(_abc_42016_n565), .C(opcode_2_), .Y(_abc_42016_n721) );
  OAI21X1 OAI21X1_310 ( .A(_abc_42016_n1624), .B(_abc_42016_n934), .C(_abc_42016_n720), .Y(_abc_42016_n1750_1) );
  OAI21X1 OAI21X1_311 ( .A(_abc_42016_n1752), .B(_abc_42016_n1751), .C(_abc_42016_n607), .Y(_abc_42016_n1753) );
  OAI21X1 OAI21X1_312 ( .A(_abc_42016_n1261), .B(_abc_42016_n587), .C(_abc_42016_n1753), .Y(_abc_42016_n1754) );
  OAI21X1 OAI21X1_313 ( .A(_abc_42016_n1749_1), .B(_abc_42016_n1750_1), .C(_abc_42016_n1756), .Y(_abc_36783_n3572) );
  OAI21X1 OAI21X1_314 ( .A(_abc_42016_n641), .B(_abc_42016_n651_1), .C(_abc_42016_n660), .Y(_abc_42016_n1758) );
  OAI21X1 OAI21X1_315 ( .A(_abc_42016_n618), .B(_abc_42016_n1760), .C(_abc_42016_n607), .Y(_abc_42016_n1761) );
  OAI21X1 OAI21X1_316 ( .A(_abc_42016_n1302), .B(_abc_42016_n587), .C(_abc_42016_n1761), .Y(_abc_42016_n1762) );
  OAI21X1 OAI21X1_317 ( .A(_abc_42016_n1624), .B(_abc_42016_n971), .C(_abc_42016_n720), .Y(_abc_42016_n1765) );
  OAI21X1 OAI21X1_318 ( .A(_abc_42016_n1764), .B(_abc_42016_n1765), .C(_abc_42016_n1763), .Y(_abc_36783_n3575) );
  OAI21X1 OAI21X1_319 ( .A(_abc_42016_n1631), .B(_abc_42016_n1767_1), .C(_abc_42016_n692), .Y(_abc_42016_n1768) );
  OAI21X1 OAI21X1_32 ( .A(regfil_5__1_), .B(_abc_42016_n626), .C(_abc_42016_n724), .Y(_abc_42016_n725) );
  OAI21X1 OAI21X1_320 ( .A(_abc_42016_n1655), .B(_abc_42016_n1660), .C(_abc_42016_n691), .Y(_abc_42016_n1772) );
  OAI21X1 OAI21X1_321 ( .A(_abc_42016_n691), .B(_abc_42016_n1771), .C(_abc_42016_n1772), .Y(_abc_36783_n3640) );
  OAI21X1 OAI21X1_322 ( .A(_abc_42016_n753), .B(_abc_42016_n1767_1), .C(_abc_42016_n692), .Y(_abc_42016_n1774) );
  OAI21X1 OAI21X1_323 ( .A(_abc_42016_n1696), .B(_abc_42016_n1703), .C(_abc_42016_n691), .Y(_abc_42016_n1778) );
  OAI21X1 OAI21X1_324 ( .A(_abc_42016_n691), .B(_abc_42016_n1777), .C(_abc_42016_n1778), .Y(_abc_36783_n3644) );
  OAI21X1 OAI21X1_325 ( .A(_abc_42016_n847), .B(_abc_42016_n1767_1), .C(_abc_42016_n692), .Y(_abc_42016_n1780) );
  OAI21X1 OAI21X1_326 ( .A(_abc_42016_n1783_1), .B(_abc_42016_n909), .C(_abc_42016_n1784_1), .Y(_abc_42016_n1785) );
  OAI21X1 OAI21X1_327 ( .A(_abc_42016_n692), .B(_abc_42016_n1747), .C(_abc_42016_n1785), .Y(_abc_36783_n3648) );
  OAI21X1 OAI21X1_328 ( .A(_abc_42016_n919), .B(_abc_42016_n1738), .C(_abc_42016_n822), .Y(_abc_42016_n1787) );
  OAI21X1 OAI21X1_329 ( .A(_abc_42016_n1792), .B(_abc_42016_n1788), .C(_abc_42016_n1794), .Y(_abc_42016_n1795) );
  OAI21X1 OAI21X1_33 ( .A(regfil_3__1_), .B(_abc_42016_n565), .C(_abc_42016_n536), .Y(_abc_42016_n726) );
  OAI21X1 OAI21X1_330 ( .A(_abc_42016_n1604_1), .B(_abc_42016_n599), .C(_abc_42016_n919), .Y(_abc_42016_n1797) );
  OAI21X1 OAI21X1_331 ( .A(_abc_42016_n1783_1), .B(_abc_42016_n934), .C(_abc_42016_n1797), .Y(_abc_42016_n1798) );
  OAI21X1 OAI21X1_332 ( .A(_abc_42016_n1801_1), .B(_abc_42016_n697), .C(_abc_42016_n688), .Y(_abc_42016_n1802_1) );
  OAI21X1 OAI21X1_333 ( .A(regfil_2__6_), .B(_abc_42016_n1733), .C(_abc_42016_n779), .Y(_abc_42016_n1803) );
  OAI21X1 OAI21X1_334 ( .A(_abc_42016_n772), .B(_abc_42016_n1805), .C(_abc_42016_n1789), .Y(_abc_42016_n1806) );
  OAI21X1 OAI21X1_335 ( .A(_abc_42016_n1604_1), .B(_abc_42016_n599), .C(_abc_42016_n964), .Y(_abc_42016_n1810) );
  OAI21X1 OAI21X1_336 ( .A(_abc_42016_n1783_1), .B(_abc_42016_n971), .C(_abc_42016_n1810), .Y(_abc_42016_n1811) );
  OAI21X1 OAI21X1_337 ( .A(_abc_42016_n714), .B(_abc_42016_n737), .C(_abc_42016_n1815), .Y(_abc_42016_n1818) );
  OAI21X1 OAI21X1_338 ( .A(_abc_42016_n723), .B(_abc_42016_n1815), .C(_abc_42016_n1818), .Y(_abc_36783_n3732) );
  OAI21X1 OAI21X1_339 ( .A(_abc_42016_n758), .B(_abc_42016_n1815), .C(_abc_42016_n1820_1), .Y(_abc_36783_n3733) );
  OAI21X1 OAI21X1_34 ( .A(regfil_0__1_), .B(_abc_42016_n727), .C(_abc_42016_n729), .Y(_abc_42016_n730) );
  OAI21X1 OAI21X1_340 ( .A(_abc_42016_n810_1), .B(_abc_42016_n817), .C(_abc_42016_n1815), .Y(_abc_42016_n1822) );
  OAI21X1 OAI21X1_341 ( .A(_abc_42016_n799), .B(_abc_42016_n1815), .C(_abc_42016_n1822), .Y(_abc_36783_n3734) );
  OAI21X1 OAI21X1_342 ( .A(_abc_42016_n1826), .B(_abc_42016_n1815), .C(_abc_42016_n1827), .Y(_abc_36783_n3736) );
  OAI21X1 OAI21X1_343 ( .A(_abc_42016_n1829), .B(_abc_42016_n1815), .C(_abc_42016_n1830), .Y(_abc_36783_n3737) );
  OAI21X1 OAI21X1_344 ( .A(_abc_42016_n951), .B(_abc_42016_n970), .C(_abc_42016_n1815), .Y(_abc_42016_n1833) );
  OAI21X1 OAI21X1_345 ( .A(_abc_42016_n1832), .B(_abc_42016_n1815), .C(_abc_42016_n1833), .Y(_abc_36783_n3738) );
  OAI21X1 OAI21X1_346 ( .A(opcode_7_), .B(_abc_42016_n540), .C(_abc_42016_n557), .Y(_abc_42016_n1836) );
  OAI21X1 OAI21X1_347 ( .A(_abc_42016_n630), .B(_abc_42016_n625), .C(opcode_2_), .Y(_abc_42016_n1837_1) );
  OAI21X1 OAI21X1_348 ( .A(_abc_42016_n1835), .B(_abc_42016_n674), .C(_abc_42016_n1838_1), .Y(_abc_42016_n1839) );
  OAI21X1 OAI21X1_349 ( .A(_abc_42016_n540), .B(_abc_42016_n1841), .C(opcode_7_), .Y(_abc_42016_n1842) );
  OAI21X1 OAI21X1_35 ( .A(_abc_42016_n719), .B(_abc_42016_n527), .C(_abc_42016_n733), .Y(_abc_42016_n734) );
  OAI21X1 OAI21X1_350 ( .A(_abc_42016_n566), .B(_abc_42016_n1844), .C(_abc_42016_n1840), .Y(alusel_0__FF_INPUT) );
  OAI21X1 OAI21X1_351 ( .A(_abc_42016_n1846), .B(_abc_42016_n1376), .C(_abc_42016_n1372), .Y(_abc_42016_n1847) );
  OAI21X1 OAI21X1_352 ( .A(alu_sel_1_), .B(_abc_42016_n1841), .C(_abc_42016_n673), .Y(_abc_42016_n1850) );
  OAI21X1 OAI21X1_353 ( .A(_abc_42016_n1849), .B(_abc_42016_n1850), .C(_abc_42016_n1852), .Y(_abc_42016_n1853) );
  OAI21X1 OAI21X1_354 ( .A(opcode_5_), .B(_abc_42016_n1848), .C(_abc_42016_n673), .Y(_abc_42016_n1856_1) );
  OAI21X1 OAI21X1_355 ( .A(_abc_42016_n530), .B(_abc_42016_n1844), .C(_abc_42016_n1858), .Y(alusel_2__FF_INPUT) );
  OAI21X1 OAI21X1_356 ( .A(_abc_42016_n1842), .B(_abc_42016_n558), .C(alu_cin), .Y(_abc_42016_n1861) );
  OAI21X1 OAI21X1_357 ( .A(_abc_42016_n1860), .B(_abc_42016_n1844), .C(_abc_42016_n1861), .Y(alucin_FF_INPUT) );
  OAI21X1 OAI21X1_358 ( .A(_abc_42016_n560), .B(_abc_42016_n1837_1), .C(_abc_42016_n1864), .Y(_abc_42016_n1865) );
  OAI21X1 OAI21X1_359 ( .A(_abc_42016_n1871), .B(_abc_42016_n1872), .C(_abc_42016_n1868), .Y(_abc_42016_n1873_1) );
  OAI21X1 OAI21X1_36 ( .A(_abc_42016_n732), .B(_abc_42016_n734), .C(_abc_42016_n720), .Y(_abc_42016_n735) );
  OAI21X1 OAI21X1_360 ( .A(_abc_42016_n558), .B(_abc_42016_n1866), .C(_abc_42016_n1876), .Y(aluoprb_0__FF_INPUT) );
  OAI21X1 OAI21X1_361 ( .A(opcode_7_), .B(_abc_42016_n1879_1), .C(_abc_42016_n540), .Y(_abc_42016_n1880) );
  OAI21X1 OAI21X1_362 ( .A(_abc_42016_n1878), .B(_abc_42016_n1881), .C(_abc_42016_n1883), .Y(aluoprb_1__FF_INPUT) );
  OAI21X1 OAI21X1_363 ( .A(_abc_42016_n1885), .B(_abc_42016_n1881), .C(_abc_42016_n1886_1), .Y(aluoprb_2__FF_INPUT) );
  OAI21X1 OAI21X1_364 ( .A(_abc_42016_n1888_1), .B(_abc_42016_n1881), .C(_abc_42016_n1889), .Y(aluoprb_3__FF_INPUT) );
  OAI21X1 OAI21X1_365 ( .A(_abc_42016_n1891), .B(_abc_42016_n1881), .C(_abc_42016_n1892), .Y(aluoprb_4__FF_INPUT) );
  OAI21X1 OAI21X1_366 ( .A(_abc_42016_n1894_1), .B(_abc_42016_n1881), .C(_abc_42016_n1895), .Y(aluoprb_5__FF_INPUT) );
  OAI21X1 OAI21X1_367 ( .A(_abc_42016_n1897), .B(_abc_42016_n1881), .C(_abc_42016_n1898), .Y(aluoprb_6__FF_INPUT) );
  OAI21X1 OAI21X1_368 ( .A(_abc_42016_n558), .B(_abc_42016_n1900), .C(_abc_42016_n1901_1), .Y(aluoprb_7__FF_INPUT) );
  OAI21X1 OAI21X1_369 ( .A(opcode_4_), .B(regfil_1__0_), .C(_abc_42016_n1903_1), .Y(_abc_42016_n1904) );
  OAI21X1 OAI21X1_37 ( .A(_abc_42016_n719), .B(_abc_42016_n587), .C(_abc_42016_n735), .Y(_abc_42016_n736) );
  OAI21X1 OAI21X1_370 ( .A(opcode_4_), .B(_abc_42016_n608), .C(_abc_42016_n566), .Y(_abc_42016_n1906) );
  OAI21X1 OAI21X1_371 ( .A(_abc_42016_n1631), .B(_abc_42016_n533), .C(_abc_42016_n530), .Y(_abc_42016_n1907) );
  OAI21X1 OAI21X1_372 ( .A(_abc_42016_n1376), .B(_abc_42016_n1371), .C(_abc_42016_n559), .Y(_abc_42016_n1909_1) );
  OAI21X1 OAI21X1_373 ( .A(_abc_42016_n629), .B(_abc_42016_n1912), .C(_abc_42016_n1913), .Y(_abc_42016_n1914) );
  OAI21X1 OAI21X1_374 ( .A(_abc_42016_n695), .B(_abc_42016_n1916), .C(_abc_42016_n1918), .Y(_abc_42016_n1919) );
  OAI21X1 OAI21X1_375 ( .A(_abc_42016_n1914), .B(_abc_42016_n1919), .C(_abc_42016_n1910), .Y(_abc_42016_n1920) );
  OAI21X1 OAI21X1_376 ( .A(_abc_42016_n547), .B(_abc_42016_n1924), .C(_abc_42016_n529), .Y(_abc_42016_n1925) );
  OAI21X1 OAI21X1_377 ( .A(opcode_6_), .B(_abc_42016_n1837_1), .C(_abc_42016_n1842), .Y(_abc_42016_n1927) );
  OAI21X1 OAI21X1_378 ( .A(_abc_42016_n558), .B(_abc_42016_n1927), .C(_abc_42016_n1926_1), .Y(_abc_42016_n1928) );
  OAI21X1 OAI21X1_379 ( .A(_abc_42016_n709), .B(_abc_42016_n1916), .C(opcode_5_), .Y(_abc_42016_n1934) );
  OAI21X1 OAI21X1_38 ( .A(regfil_3__1_), .B(_abc_42016_n600), .C(_abc_42016_n692), .Y(_abc_42016_n741) );
  OAI21X1 OAI21X1_380 ( .A(_abc_42016_n1427), .B(_abc_42016_n1935), .C(_abc_42016_n1936), .Y(_abc_42016_n1937) );
  OAI21X1 OAI21X1_381 ( .A(_abc_42016_n712), .B(_abc_42016_n1912), .C(_abc_42016_n530), .Y(_abc_42016_n1938) );
  OAI21X1 OAI21X1_382 ( .A(_abc_42016_n703), .B(_abc_42016_n1935), .C(_abc_42016_n1939), .Y(_abc_42016_n1940) );
  OAI21X1 OAI21X1_383 ( .A(_abc_42016_n1938), .B(_abc_42016_n1940), .C(_abc_42016_n1910), .Y(_abc_42016_n1941) );
  OAI21X1 OAI21X1_384 ( .A(_abc_42016_n1934), .B(_abc_42016_n1937), .C(_abc_42016_n1942), .Y(_abc_42016_n1943) );
  OAI21X1 OAI21X1_385 ( .A(_abc_42016_n1427), .B(_abc_42016_n1842), .C(_abc_42016_n1943), .Y(_abc_42016_n1944) );
  OAI21X1 OAI21X1_386 ( .A(_abc_42016_n558), .B(_abc_42016_n1945), .C(_abc_42016_n1946), .Y(aluopra_1__FF_INPUT) );
  OAI21X1 OAI21X1_387 ( .A(_abc_42016_n773), .B(_abc_42016_n1935), .C(_abc_42016_n530), .Y(_abc_42016_n1948) );
  OAI21X1 OAI21X1_388 ( .A(_abc_42016_n757), .B(_abc_42016_n1916), .C(opcode_5_), .Y(_abc_42016_n1952_1) );
  OAI21X1 OAI21X1_389 ( .A(_abc_42016_n758), .B(_abc_42016_n533), .C(_abc_42016_n1953), .Y(_abc_42016_n1954) );
  OAI21X1 OAI21X1_39 ( .A(_abc_42016_n741), .B(_abc_42016_n740), .C(_abc_42016_n711), .Y(_abc_36783_n3364) );
  OAI21X1 OAI21X1_390 ( .A(_abc_42016_n1952_1), .B(_abc_42016_n1954), .C(_abc_42016_n1910), .Y(_abc_42016_n1955_1) );
  OAI21X1 OAI21X1_391 ( .A(_abc_42016_n799), .B(_abc_42016_n533), .C(opcode_5_), .Y(_abc_42016_n1961_1) );
  OAI21X1 OAI21X1_392 ( .A(_abc_42016_n1488), .B(_abc_42016_n1935), .C(_abc_42016_n1962), .Y(_abc_42016_n1963_1) );
  OAI21X1 OAI21X1_393 ( .A(_abc_42016_n812), .B(_abc_42016_n1912), .C(_abc_42016_n530), .Y(_abc_42016_n1964) );
  OAI21X1 OAI21X1_394 ( .A(_abc_42016_n795), .B(_abc_42016_n1935), .C(_abc_42016_n1965), .Y(_abc_42016_n1966_1) );
  OAI21X1 OAI21X1_395 ( .A(_abc_42016_n1964), .B(_abc_42016_n1966_1), .C(_abc_42016_n1910), .Y(_abc_42016_n1967) );
  OAI21X1 OAI21X1_396 ( .A(_abc_42016_n1961_1), .B(_abc_42016_n1963_1), .C(_abc_42016_n1968_1), .Y(_abc_42016_n1969) );
  OAI21X1 OAI21X1_397 ( .A(_abc_42016_n1488), .B(_abc_42016_n1842), .C(_abc_42016_n1969), .Y(_abc_42016_n1970) );
  OAI21X1 OAI21X1_398 ( .A(_abc_42016_n558), .B(_abc_42016_n1971), .C(_abc_42016_n1972), .Y(aluopra_3__FF_INPUT) );
  OAI21X1 OAI21X1_399 ( .A(_abc_42016_n1974), .B(_abc_42016_n1935), .C(opcode_5_), .Y(_abc_42016_n1975) );
  OAI21X1 OAI21X1_4 ( .A(_abc_42016_n552), .B(_abc_42016_n526_1), .C(_abc_42016_n551), .Y(_abc_42016_n553) );
  OAI21X1 OAI21X1_40 ( .A(_abc_42016_n743), .B(_abc_42016_n744), .C(_abc_42016_n660), .Y(_abc_42016_n745) );
  OAI21X1 OAI21X1_400 ( .A(_abc_42016_n842), .B(_abc_42016_n1912), .C(_abc_42016_n1976), .Y(_abc_42016_n1977) );
  OAI21X1 OAI21X1_401 ( .A(_abc_42016_n861), .B(_abc_42016_n1935), .C(_abc_42016_n530), .Y(_abc_42016_n1978) );
  OAI21X1 OAI21X1_402 ( .A(opcode_3_), .B(_abc_42016_n1515), .C(_abc_42016_n1979), .Y(_abc_42016_n1980) );
  OAI21X1 OAI21X1_403 ( .A(_abc_42016_n1975), .B(_abc_42016_n1977), .C(_abc_42016_n1981), .Y(_abc_42016_n1982) );
  OAI21X1 OAI21X1_404 ( .A(_abc_42016_n1974), .B(_abc_42016_n1842), .C(_abc_42016_n1982), .Y(_abc_42016_n1983) );
  OAI21X1 OAI21X1_405 ( .A(_abc_42016_n558), .B(_abc_42016_n1984), .C(_abc_42016_n1985), .Y(aluopra_4__FF_INPUT) );
  OAI21X1 OAI21X1_406 ( .A(_abc_42016_n895), .B(_abc_42016_n533), .C(_abc_42016_n530), .Y(_abc_42016_n1987) );
  OAI21X1 OAI21X1_407 ( .A(_abc_42016_n874), .B(_abc_42016_n1935), .C(_abc_42016_n1988), .Y(_abc_42016_n1989) );
  OAI21X1 OAI21X1_408 ( .A(_abc_42016_n898), .B(_abc_42016_n1935), .C(_abc_42016_n1990), .Y(_abc_42016_n1991) );
  OAI21X1 OAI21X1_409 ( .A(_abc_42016_n872), .B(_abc_42016_n1916), .C(_abc_42016_n1992), .Y(_abc_42016_n1993) );
  OAI21X1 OAI21X1_41 ( .A(regfil_0__1_), .B(_abc_42016_n619), .C(regfil_0__2_), .Y(_abc_42016_n749) );
  OAI21X1 OAI21X1_410 ( .A(_abc_42016_n1987), .B(_abc_42016_n1989), .C(_abc_42016_n1994), .Y(_abc_42016_n1995) );
  OAI21X1 OAI21X1_411 ( .A(_abc_42016_n898), .B(_abc_42016_n1842), .C(_abc_42016_n1995), .Y(_abc_42016_n1996) );
  OAI21X1 OAI21X1_412 ( .A(_abc_42016_n558), .B(_abc_42016_n1997), .C(_abc_42016_n1998), .Y(aluopra_5__FF_INPUT) );
  OAI21X1 OAI21X1_413 ( .A(opcode_3_), .B(_abc_42016_n1573), .C(_abc_42016_n2000), .Y(_abc_42016_n2001) );
  OAI21X1 OAI21X1_414 ( .A(_abc_42016_n1829), .B(_abc_42016_n533), .C(opcode_5_), .Y(_abc_42016_n2003) );
  OAI21X1 OAI21X1_415 ( .A(_abc_42016_n1554), .B(_abc_42016_n1912), .C(_abc_42016_n2004), .Y(_abc_42016_n2005) );
  OAI21X1 OAI21X1_416 ( .A(_abc_42016_n2003), .B(_abc_42016_n2005), .C(_abc_42016_n1910), .Y(_abc_42016_n2006) );
  OAI21X1 OAI21X1_417 ( .A(_abc_42016_n558), .B(_abc_42016_n2008), .C(_abc_42016_n2009), .Y(aluopra_6__FF_INPUT) );
  OAI21X1 OAI21X1_418 ( .A(_abc_42016_n960), .B(_abc_42016_n1935), .C(opcode_5_), .Y(_abc_42016_n2011) );
  OAI21X1 OAI21X1_419 ( .A(_abc_42016_n959), .B(_abc_42016_n1916), .C(_abc_42016_n2013), .Y(_abc_42016_n2014) );
  OAI21X1 OAI21X1_42 ( .A(regfil_4__2_), .B(_abc_42016_n727), .C(opcode_2_), .Y(_abc_42016_n756) );
  OAI21X1 OAI21X1_420 ( .A(_abc_42016_n974), .B(_abc_42016_n1935), .C(_abc_42016_n530), .Y(_abc_42016_n2016) );
  OAI21X1 OAI21X1_421 ( .A(_abc_42016_n960), .B(_abc_42016_n1842), .C(_abc_42016_n2019), .Y(_abc_42016_n2020) );
  OAI21X1 OAI21X1_422 ( .A(_abc_42016_n558), .B(_abc_42016_n2021), .C(_abc_42016_n2022), .Y(aluopra_7__FF_INPUT) );
  OAI21X1 OAI21X1_423 ( .A(intcyc), .B(_abc_42016_n2026), .C(_abc_42016_n529), .Y(_abc_42016_n2027) );
  OAI21X1 OAI21X1_424 ( .A(state_4_), .B(_abc_42016_n509), .C(_abc_42016_n2035), .Y(_abc_42016_n2036) );
  OAI21X1 OAI21X1_425 ( .A(_abc_42016_n2032), .B(_abc_42016_n2036), .C(_abc_42016_n529), .Y(_abc_42016_n2037) );
  OAI21X1 OAI21X1_426 ( .A(_abc_42016_n2039), .B(_abc_42016_n2045), .C(_abc_42016_n2038), .Y(_abc_42016_n2046) );
  OAI21X1 OAI21X1_427 ( .A(_abc_42016_n2029), .B(_abc_42016_n2048), .C(_abc_42016_n2046), .Y(parity_FF_INPUT) );
  OAI21X1 OAI21X1_428 ( .A(_abc_42016_n686), .B(_abc_42016_n992), .C(zero), .Y(_abc_42016_n2052) );
  OAI21X1 OAI21X1_429 ( .A(_abc_42016_n1261), .B(_abc_42016_n2042), .C(_abc_42016_n2052), .Y(_abc_42016_n2053) );
  OAI21X1 OAI21X1_43 ( .A(regfil_7__2_), .B(_abc_42016_n565), .C(_abc_42016_n759), .Y(_abc_42016_n760) );
  OAI21X1 OAI21X1_430 ( .A(_abc_42016_n2050), .B(_abc_42016_n2038), .C(_abc_42016_n2054), .Y(zero_FF_INPUT) );
  OAI21X1 OAI21X1_431 ( .A(_abc_42016_n2058), .B(_abc_42016_n2035), .C(_abc_42016_n2060), .Y(_abc_42016_n2061) );
  OAI21X1 OAI21X1_432 ( .A(_abc_42016_n2061), .B(_abc_42016_n2057), .C(_abc_42016_n2038), .Y(_abc_42016_n2062) );
  OAI21X1 OAI21X1_433 ( .A(_abc_42016_n2056), .B(_abc_42016_n2048), .C(_abc_42016_n2062), .Y(sign_FF_INPUT) );
  OAI21X1 OAI21X1_434 ( .A(reset), .B(_abc_42016_n548), .C(_abc_42016_n2037), .Y(_abc_42016_n2065) );
  OAI21X1 OAI21X1_435 ( .A(regfil_7__2_), .B(regfil_7__1_), .C(regfil_7__3_), .Y(_abc_42016_n2066) );
  OAI21X1 OAI21X1_436 ( .A(auxcar), .B(_abc_42016_n2072), .C(_abc_42016_n547), .Y(_abc_42016_n2073) );
  OAI21X1 OAI21X1_437 ( .A(_abc_42016_n2071), .B(_abc_42016_n2073), .C(_abc_42016_n2074), .Y(_abc_42016_n2075) );
  OAI21X1 OAI21X1_438 ( .A(_abc_42016_n2080), .B(_abc_42016_n2081), .C(_abc_42016_n529), .Y(_abc_42016_n2082) );
  OAI21X1 OAI21X1_439 ( .A(_abc_42016_n680), .B(_abc_42016_n2084), .C(_abc_42016_n2087), .Y(_abc_42016_n2088) );
  OAI21X1 OAI21X1_44 ( .A(regfil_3__2_), .B(_abc_42016_n600), .C(_abc_42016_n692), .Y(_abc_42016_n771) );
  OAI21X1 OAI21X1_440 ( .A(_abc_42016_n568), .B(_abc_42016_n626), .C(_abc_42016_n2090), .Y(_abc_42016_n2091) );
  OAI21X1 OAI21X1_441 ( .A(_abc_42016_n2091), .B(_abc_42016_n2088), .C(_abc_42016_n559), .Y(_abc_42016_n2092) );
  OAI21X1 OAI21X1_442 ( .A(_abc_42016_n566), .B(_abc_42016_n1860), .C(_abc_42016_n1003), .Y(_abc_42016_n2096) );
  OAI21X1 OAI21X1_443 ( .A(_abc_42016_n628), .B(_abc_42016_n2087), .C(_abc_42016_n2098), .Y(_abc_42016_n2099) );
  OAI21X1 OAI21X1_444 ( .A(_abc_42016_n1554), .B(_abc_42016_n2103), .C(_abc_42016_n2142), .Y(_abc_42016_n2143_1) );
  OAI21X1 OAI21X1_445 ( .A(_abc_42016_n2102_1), .B(_abc_42016_n2143_1), .C(_abc_42016_n1005), .Y(_abc_42016_n2144_1) );
  OAI21X1 OAI21X1_446 ( .A(_abc_42016_n2083), .B(_abc_42016_n2144_1), .C(_abc_42016_n2100), .Y(_abc_42016_n2145) );
  OAI21X1 OAI21X1_447 ( .A(_abc_42016_n2147), .B(_abc_42016_n2177), .C(_abc_42016_n1000), .Y(_abc_42016_n2178) );
  OAI21X1 OAI21X1_448 ( .A(_abc_42016_n913), .B(_abc_42016_n1554), .C(_abc_42016_n2209), .Y(_abc_42016_n2210) );
  OAI21X1 OAI21X1_449 ( .A(_abc_42016_n2179), .B(_abc_42016_n2210), .C(_abc_42016_n2212), .Y(_abc_42016_n2213) );
  OAI21X1 OAI21X1_45 ( .A(_abc_42016_n634), .B(_abc_42016_n703), .C(_abc_42016_n773), .Y(_abc_42016_n774) );
  OAI21X1 OAI21X1_450 ( .A(_abc_42016_n2146), .B(_abc_42016_n2178), .C(_abc_42016_n2213), .Y(_abc_42016_n2214) );
  OAI21X1 OAI21X1_451 ( .A(_abc_42016_n2145), .B(_abc_42016_n2214), .C(_abc_42016_n2215), .Y(_abc_42016_n2216) );
  OAI21X1 OAI21X1_452 ( .A(regfil_7__5_), .B(regfil_7__6_), .C(regfil_7__7_), .Y(_abc_42016_n2218) );
  OAI21X1 OAI21X1_453 ( .A(_abc_42016_n2218), .B(_abc_42016_n2217), .C(_abc_42016_n2219), .Y(_abc_42016_n2220) );
  OAI21X1 OAI21X1_454 ( .A(_abc_42016_n1044), .B(_abc_42016_n2044), .C(_abc_42016_n2221), .Y(_abc_42016_n2222) );
  OAI21X1 OAI21X1_455 ( .A(_abc_42016_n2231), .B(_abc_42016_n2228), .C(opcode_0_), .Y(_abc_42016_n2232) );
  OAI21X1 OAI21X1_456 ( .A(_abc_42016_n2225), .B(_abc_42016_n2230), .C(_abc_42016_n2232), .Y(opcode_0__FF_INPUT) );
  OAI21X1 OAI21X1_457 ( .A(_abc_42016_n2231), .B(_abc_42016_n2228), .C(opcode_1_), .Y(_abc_42016_n2235) );
  OAI21X1 OAI21X1_458 ( .A(_abc_42016_n2234), .B(_abc_42016_n2230), .C(_abc_42016_n2235), .Y(opcode_1__FF_INPUT) );
  OAI21X1 OAI21X1_459 ( .A(_abc_42016_n2231), .B(_abc_42016_n2228), .C(opcode_2_), .Y(_abc_42016_n2238) );
  OAI21X1 OAI21X1_46 ( .A(regfil_3__0_), .B(regfil_3__1_), .C(regfil_3__2_), .Y(_abc_42016_n780) );
  OAI21X1 OAI21X1_460 ( .A(_abc_42016_n2237), .B(_abc_42016_n2230), .C(_abc_42016_n2238), .Y(opcode_2__FF_INPUT) );
  OAI21X1 OAI21X1_461 ( .A(_abc_42016_n2231), .B(_abc_42016_n2228), .C(opcode_3_), .Y(_abc_42016_n2241) );
  OAI21X1 OAI21X1_462 ( .A(_abc_42016_n2240), .B(_abc_42016_n2230), .C(_abc_42016_n2241), .Y(opcode_3__FF_INPUT) );
  OAI21X1 OAI21X1_463 ( .A(_abc_42016_n2231), .B(_abc_42016_n2228), .C(opcode_4_), .Y(_abc_42016_n2244) );
  OAI21X1 OAI21X1_464 ( .A(_abc_42016_n2243), .B(_abc_42016_n2230), .C(_abc_42016_n2244), .Y(opcode_4__FF_INPUT) );
  OAI21X1 OAI21X1_465 ( .A(_abc_42016_n2231), .B(_abc_42016_n2228), .C(opcode_7_), .Y(_abc_42016_n2251) );
  OAI21X1 OAI21X1_466 ( .A(_abc_42016_n2250), .B(_abc_42016_n2230), .C(_abc_42016_n2251), .Y(opcode_7__FF_INPUT) );
  OAI21X1 OAI21X1_467 ( .A(_abc_42016_n1004), .B(_abc_42016_n682), .C(_abc_42016_n2255), .Y(_abc_42016_n2256) );
  OAI21X1 OAI21X1_468 ( .A(_abc_42016_n2256), .B(_abc_42016_n678), .C(_abc_42016_n2257), .Y(eienb_FF_INPUT) );
  OAI21X1 OAI21X1_469 ( .A(_abc_42016_n1923), .B(_abc_42016_n2033), .C(_abc_42016_n2261), .Y(_abc_42016_n2262) );
  OAI21X1 OAI21X1_47 ( .A(_abc_42016_n781), .B(_abc_42016_n783), .C(_abc_42016_n779), .Y(_abc_42016_n784) );
  OAI21X1 OAI21X1_470 ( .A(_abc_42016_n1869), .B(_abc_42016_n522), .C(_abc_42016_n519), .Y(_abc_42016_n2263) );
  OAI21X1 OAI21X1_471 ( .A(_abc_42016_n2031), .B(_abc_42016_n2263), .C(_abc_42016_n1014), .Y(_abc_42016_n2264) );
  OAI21X1 OAI21X1_472 ( .A(_abc_42016_n1923), .B(_abc_42016_n509), .C(_abc_42016_n2267), .Y(_abc_42016_n2268) );
  OAI21X1 OAI21X1_473 ( .A(_abc_42016_n581_1), .B(_abc_42016_n1923), .C(_abc_42016_n2272), .Y(_abc_42016_n2273) );
  OAI21X1 OAI21X1_474 ( .A(state_5_), .B(_abc_42016_n546), .C(_abc_42016_n2276), .Y(_abc_42016_n2277) );
  OAI21X1 OAI21X1_475 ( .A(_abc_42016_n1346), .B(_abc_42016_n2281), .C(_abc_42016_n668), .Y(_abc_42016_n2282) );
  OAI21X1 OAI21X1_476 ( .A(_abc_42016_n539), .B(_abc_42016_n2254), .C(_abc_42016_n2282), .Y(_abc_42016_n2283) );
  OAI21X1 OAI21X1_477 ( .A(_abc_42016_n572), .B(_abc_42016_n626), .C(_abc_42016_n2284), .Y(_abc_42016_n2285) );
  OAI21X1 OAI21X1_478 ( .A(_abc_42016_n1346), .B(_abc_42016_n2281), .C(_abc_42016_n530), .Y(_abc_42016_n2286) );
  OAI21X1 OAI21X1_479 ( .A(_abc_42016_n536), .B(_abc_42016_n564), .C(_abc_42016_n2286), .Y(_abc_42016_n2287) );
  OAI21X1 OAI21X1_48 ( .A(_abc_42016_n757), .B(_abc_42016_n697), .C(_abc_42016_n785), .Y(_abc_42016_n786) );
  OAI21X1 OAI21X1_480 ( .A(_abc_42016_n2287), .B(_abc_42016_n2285), .C(_abc_42016_n1837_1), .Y(_abc_42016_n2289) );
  OAI21X1 OAI21X1_481 ( .A(_abc_42016_n2280), .B(_abc_42016_n2288), .C(_abc_42016_n2289), .Y(_abc_42016_n2290) );
  OAI21X1 OAI21X1_482 ( .A(opcode_5_), .B(_abc_42016_n1347), .C(_abc_42016_n1848), .Y(_abc_42016_n2293) );
  OAI21X1 OAI21X1_483 ( .A(_abc_42016_n2259), .B(_abc_42016_n2290), .C(_abc_42016_n2294), .Y(_abc_42016_n2295) );
  OAI21X1 OAI21X1_484 ( .A(opcode_3_), .B(_abc_42016_n1004), .C(_abc_42016_n1841), .Y(_abc_42016_n2300) );
  OAI21X1 OAI21X1_485 ( .A(_abc_42016_n536), .B(_abc_42016_n539), .C(_abc_42016_n1851), .Y(_abc_42016_n2301) );
  OAI21X1 OAI21X1_486 ( .A(_abc_42016_n541), .B(_abc_42016_n2302), .C(_abc_42016_n2300), .Y(_abc_42016_n2303) );
  OAI21X1 OAI21X1_487 ( .A(statesel_0_), .B(_abc_42016_n2299), .C(_abc_42016_n2304), .Y(_abc_42016_n2305) );
  OAI21X1 OAI21X1_488 ( .A(_abc_42016_n572), .B(_abc_42016_n626), .C(_abc_42016_n1408), .Y(_abc_42016_n2306) );
  OAI21X1 OAI21X1_489 ( .A(_abc_42016_n2089), .B(_abc_42016_n682), .C(_abc_42016_n1848), .Y(_abc_42016_n2307) );
  OAI21X1 OAI21X1_49 ( .A(_abc_42016_n771), .B(_abc_42016_n770), .C(_abc_42016_n787), .Y(_abc_36783_n3367) );
  OAI21X1 OAI21X1_490 ( .A(_abc_42016_n680), .B(_abc_42016_n1347), .C(_abc_42016_n2310), .Y(_abc_42016_n2311) );
  OAI21X1 OAI21X1_491 ( .A(_abc_42016_n1346), .B(_abc_42016_n573), .C(_abc_42016_n570), .Y(_abc_42016_n2313) );
  OAI21X1 OAI21X1_492 ( .A(_abc_42016_n536), .B(_abc_42016_n539), .C(_abc_42016_n2315), .Y(_abc_42016_n2316) );
  OAI21X1 OAI21X1_493 ( .A(_abc_42016_n682), .B(_abc_42016_n669), .C(_abc_42016_n2318), .Y(_abc_42016_n2319) );
  OAI21X1 OAI21X1_494 ( .A(_abc_42016_n569), .B(_abc_42016_n573), .C(_abc_42016_n679), .Y(_abc_42016_n2322) );
  OAI21X1 OAI21X1_495 ( .A(_abc_42016_n2259), .B(_abc_42016_n2329), .C(_abc_42016_n2308), .Y(_abc_42016_n2330) );
  OAI21X1 OAI21X1_496 ( .A(_abc_42016_n2296_1), .B(_abc_42016_n2332), .C(_abc_42016_n547), .Y(_abc_42016_n2333) );
  OAI21X1 OAI21X1_497 ( .A(waitr), .B(_abc_42016_n2335), .C(_abc_42016_n2276), .Y(_abc_42016_n2336) );
  OAI21X1 OAI21X1_498 ( .A(_abc_42016_n2259), .B(_abc_42016_n2340), .C(_abc_42016_n2337), .Y(_abc_42016_n2341) );
  OAI21X1 OAI21X1_499 ( .A(_abc_42016_n2279), .B(_abc_42016_n1848), .C(_abc_42016_n2282), .Y(_abc_42016_n2346) );
  OAI21X1 OAI21X1_5 ( .A(opcode_3_), .B(_abc_42016_n528_1), .C(_abc_42016_n553), .Y(_abc_42016_n554) );
  OAI21X1 OAI21X1_50 ( .A(regfil_0__2_), .B(_abc_42016_n716), .C(regfil_0__3_), .Y(_abc_42016_n791_1) );
  OAI21X1 OAI21X1_500 ( .A(_abc_42016_n2344), .B(_abc_42016_n2290), .C(_abc_42016_n2348_1), .Y(_abc_42016_n2349) );
  OAI21X1 OAI21X1_501 ( .A(_abc_42016_n2346), .B(_abc_42016_n2349), .C(_abc_42016_n559), .Y(_abc_42016_n2350) );
  OAI21X1 OAI21X1_502 ( .A(_abc_42016_n2327), .B(_abc_42016_n2321), .C(_abc_42016_n2315), .Y(_abc_42016_n2351) );
  OAI21X1 OAI21X1_503 ( .A(_abc_42016_n2327), .B(_abc_42016_n2321), .C(_abc_42016_n673), .Y(_abc_42016_n2352) );
  OAI21X1 OAI21X1_504 ( .A(_abc_42016_n2344), .B(_abc_42016_n674), .C(_abc_42016_n2352), .Y(_abc_42016_n2353) );
  OAI21X1 OAI21X1_505 ( .A(_abc_42016_n2347_1), .B(_abc_42016_n2351), .C(_abc_42016_n2353), .Y(_abc_42016_n2354) );
  OAI21X1 OAI21X1_506 ( .A(_abc_42016_n1004), .B(_abc_42016_n2355), .C(_abc_42016_n1841), .Y(_abc_42016_n2356) );
  OAI21X1 OAI21X1_507 ( .A(_abc_42016_n566), .B(_abc_42016_n1848), .C(_abc_42016_n2356), .Y(_abc_42016_n2357) );
  OAI21X1 OAI21X1_508 ( .A(_abc_42016_n1841), .B(_abc_42016_n2280), .C(_abc_42016_n541), .Y(_abc_42016_n2358) );
  OAI21X1 OAI21X1_509 ( .A(statesel_1_), .B(_abc_42016_n2357), .C(_abc_42016_n2359), .Y(_abc_42016_n2360) );
  OAI21X1 OAI21X1_51 ( .A(_abc_42016_n794), .B(_abc_42016_n797), .C(_abc_42016_n536), .Y(_abc_42016_n798) );
  OAI21X1 OAI21X1_510 ( .A(_abc_42016_n2345), .B(_abc_42016_n2361), .C(_abc_42016_n547), .Y(_abc_42016_n2362) );
  OAI21X1 OAI21X1_511 ( .A(_abc_42016_n2363), .B(_abc_42016_n2364), .C(_abc_42016_n2336), .Y(_abc_42016_n2365) );
  OAI21X1 OAI21X1_512 ( .A(_abc_42016_n2344), .B(_abc_42016_n2340), .C(_abc_42016_n2365), .Y(_abc_42016_n2366) );
  OAI21X1 OAI21X1_513 ( .A(_abc_42016_n2279), .B(_abc_42016_n542), .C(_abc_42016_n2371), .Y(_abc_42016_n2372_1) );
  OAI21X1 OAI21X1_514 ( .A(statesel_2_), .B(_abc_42016_n2279), .C(_abc_42016_n2289), .Y(_abc_42016_n2375) );
  OAI21X1 OAI21X1_515 ( .A(opcode_5_), .B(_abc_42016_n2376), .C(_abc_42016_n2377), .Y(_abc_42016_n2378) );
  OAI21X1 OAI21X1_516 ( .A(_abc_42016_n2374), .B(_abc_42016_n2380), .C(_abc_42016_n2381), .Y(_abc_42016_n2382) );
  OAI21X1 OAI21X1_517 ( .A(_abc_42016_n2369), .B(_abc_42016_n2329), .C(_abc_42016_n2383), .Y(_abc_42016_n2384) );
  OAI21X1 OAI21X1_518 ( .A(_abc_42016_n2259), .B(_abc_42016_n2344), .C(_abc_42016_n2369), .Y(_abc_42016_n2386) );
  OAI21X1 OAI21X1_519 ( .A(_abc_42016_n2385), .B(_abc_42016_n2389), .C(_abc_42016_n2390), .Y(_abc_42016_n2391) );
  OAI21X1 OAI21X1_52 ( .A(regfil_7__3_), .B(_abc_42016_n565), .C(_abc_42016_n801), .Y(_abc_42016_n802) );
  OAI21X1 OAI21X1_520 ( .A(_abc_42016_n2398_1), .B(_abc_42016_n2396), .C(_abc_42016_n559), .Y(_abc_42016_n2399) );
  OAI21X1 OAI21X1_521 ( .A(_abc_42016_n672_1), .B(opcode_6_), .C(_abc_42016_n2373_1), .Y(_abc_42016_n2402_1) );
  OAI21X1 OAI21X1_522 ( .A(statesel_3_), .B(_abc_42016_n2403), .C(_abc_42016_n2402_1), .Y(_abc_42016_n2404) );
  OAI21X1 OAI21X1_523 ( .A(_abc_42016_n674), .B(_abc_42016_n2401), .C(_abc_42016_n2404), .Y(_abc_42016_n2405_1) );
  OAI21X1 OAI21X1_524 ( .A(_abc_42016_n2400), .B(_abc_42016_n2405_1), .C(_abc_42016_n547), .Y(_abc_42016_n2406) );
  OAI21X1 OAI21X1_525 ( .A(_abc_42016_n2031), .B(_abc_42016_n546), .C(_abc_42016_n2276), .Y(_abc_42016_n2411_1) );
  OAI21X1 OAI21X1_526 ( .A(_abc_42016_n2388), .B(_abc_42016_n2339), .C(statesel_3_), .Y(_abc_42016_n2413) );
  OAI21X1 OAI21X1_527 ( .A(_abc_42016_n2412), .B(_abc_42016_n2413), .C(_abc_42016_n2337), .Y(_abc_42016_n2414_1) );
  OAI21X1 OAI21X1_528 ( .A(statesel_4_), .B(_abc_42016_n2329), .C(_abc_42016_n673), .Y(_abc_42016_n2420_1) );
  OAI21X1 OAI21X1_529 ( .A(_abc_42016_n536), .B(_abc_42016_n539), .C(_abc_42016_n2423_1), .Y(_abc_42016_n2424) );
  OAI21X1 OAI21X1_53 ( .A(regfil_5__3_), .B(_abc_42016_n626), .C(_abc_42016_n803), .Y(_abc_42016_n804) );
  OAI21X1 OAI21X1_530 ( .A(opcode_5_), .B(_abc_42016_n2291), .C(_abc_42016_n2425), .Y(_abc_42016_n2426_1) );
  OAI21X1 OAI21X1_531 ( .A(_abc_42016_n1879_1), .B(_abc_42016_n2426_1), .C(_abc_42016_n559), .Y(_abc_42016_n2427) );
  OAI21X1 OAI21X1_532 ( .A(_abc_42016_n1376), .B(_abc_42016_n1371), .C(_abc_42016_n2279), .Y(_abc_42016_n2429_1) );
  OAI21X1 OAI21X1_533 ( .A(_abc_42016_n2417_1), .B(_abc_42016_n2422), .C(_abc_42016_n2433), .Y(_abc_42016_n2434) );
  OAI21X1 OAI21X1_534 ( .A(_abc_42016_n2434), .B(_abc_42016_n2421), .C(_abc_42016_n547), .Y(_abc_42016_n2435_1) );
  OAI21X1 OAI21X1_535 ( .A(_abc_42016_n2417_1), .B(_abc_42016_n2340), .C(_abc_42016_n2337), .Y(_abc_42016_n2443) );
  OAI21X1 OAI21X1_536 ( .A(_abc_42016_n1848), .B(_abc_42016_n1863), .C(_abc_42016_n2352), .Y(_abc_42016_n2448) );
  OAI21X1 OAI21X1_537 ( .A(_abc_42016_n2448), .B(_abc_42016_n2447_1), .C(_abc_42016_n547), .Y(_abc_42016_n2449) );
  OAI21X1 OAI21X1_538 ( .A(_abc_42016_n2376), .B(_abc_42016_n678), .C(popdes_0_), .Y(_abc_42016_n2458) );
  OAI21X1 OAI21X1_539 ( .A(_abc_42016_n531), .B(_abc_42016_n2457), .C(_abc_42016_n2458), .Y(popdes_0__FF_INPUT) );
  OAI21X1 OAI21X1_54 ( .A(_abc_42016_n528_1), .B(_abc_42016_n806), .C(_abc_42016_n807), .Y(_abc_42016_n808) );
  OAI21X1 OAI21X1_540 ( .A(_abc_42016_n2376), .B(_abc_42016_n678), .C(popdes_1_), .Y(_abc_42016_n2460) );
  OAI21X1 OAI21X1_541 ( .A(_abc_42016_n530), .B(_abc_42016_n2457), .C(_abc_42016_n2460), .Y(popdes_1__FF_INPUT) );
  OAI21X1 OAI21X1_542 ( .A(_abc_42016_n2231), .B(_abc_42016_n2335), .C(rdatahold2_0_), .Y(_abc_42016_n2463) );
  OAI21X1 OAI21X1_543 ( .A(_abc_42016_n602), .B(_abc_42016_n2462), .C(_abc_42016_n2463), .Y(rdatahold2_0__FF_INPUT) );
  OAI21X1 OAI21X1_544 ( .A(_abc_42016_n2231), .B(_abc_42016_n2335), .C(rdatahold2_1_), .Y(_abc_42016_n2465) );
  OAI21X1 OAI21X1_545 ( .A(_abc_42016_n719), .B(_abc_42016_n2462), .C(_abc_42016_n2465), .Y(rdatahold2_1__FF_INPUT) );
  OAI21X1 OAI21X1_546 ( .A(_abc_42016_n2231), .B(_abc_42016_n2335), .C(rdatahold2_2_), .Y(_abc_42016_n2467) );
  OAI21X1 OAI21X1_547 ( .A(_abc_42016_n1675), .B(_abc_42016_n2462), .C(_abc_42016_n2467), .Y(rdatahold2_2__FF_INPUT) );
  OAI21X1 OAI21X1_548 ( .A(_abc_42016_n2231), .B(_abc_42016_n2335), .C(rdatahold2_3_), .Y(_abc_42016_n2469) );
  OAI21X1 OAI21X1_549 ( .A(_abc_42016_n811), .B(_abc_42016_n2462), .C(_abc_42016_n2469), .Y(rdatahold2_3__FF_INPUT) );
  OAI21X1 OAI21X1_55 ( .A(_abc_42016_n606), .B(_abc_42016_n792), .C(_abc_42016_n809), .Y(_abc_42016_n810_1) );
  OAI21X1 OAI21X1_550 ( .A(_abc_42016_n2231), .B(_abc_42016_n2335), .C(rdatahold2_4_), .Y(_abc_42016_n2472) );
  OAI21X1 OAI21X1_551 ( .A(_abc_42016_n2471), .B(_abc_42016_n2462), .C(_abc_42016_n2472), .Y(rdatahold2_4__FF_INPUT) );
  OAI21X1 OAI21X1_552 ( .A(_abc_42016_n2231), .B(_abc_42016_n2335), .C(rdatahold2_5_), .Y(_abc_42016_n2474) );
  OAI21X1 OAI21X1_553 ( .A(_abc_42016_n891), .B(_abc_42016_n2462), .C(_abc_42016_n2474), .Y(rdatahold2_5__FF_INPUT) );
  OAI21X1 OAI21X1_554 ( .A(_abc_42016_n2231), .B(_abc_42016_n2335), .C(rdatahold2_6_), .Y(_abc_42016_n2476) );
  OAI21X1 OAI21X1_555 ( .A(_abc_42016_n1793), .B(_abc_42016_n2462), .C(_abc_42016_n2476), .Y(rdatahold2_6__FF_INPUT) );
  OAI21X1 OAI21X1_556 ( .A(_abc_42016_n2231), .B(_abc_42016_n2335), .C(rdatahold2_7_), .Y(_abc_42016_n2479) );
  OAI21X1 OAI21X1_557 ( .A(_abc_42016_n2478), .B(_abc_42016_n2462), .C(_abc_42016_n2479), .Y(rdatahold2_7__FF_INPUT) );
  OAI21X1 OAI21X1_558 ( .A(_abc_42016_n2231), .B(_abc_42016_n2335), .C(rdatahold_0_), .Y(_abc_42016_n2481) );
  OAI21X1 OAI21X1_559 ( .A(_abc_42016_n2225), .B(_abc_42016_n2462), .C(_abc_42016_n2481), .Y(rdatahold_0__FF_INPUT) );
  OAI21X1 OAI21X1_56 ( .A(_abc_42016_n743), .B(_abc_42016_n744), .C(_abc_42016_n812), .Y(_abc_42016_n813) );
  OAI21X1 OAI21X1_560 ( .A(_abc_42016_n2231), .B(_abc_42016_n2335), .C(rdatahold_1_), .Y(_abc_42016_n2483) );
  OAI21X1 OAI21X1_561 ( .A(_abc_42016_n2234), .B(_abc_42016_n2462), .C(_abc_42016_n2483), .Y(rdatahold_1__FF_INPUT) );
  OAI21X1 OAI21X1_562 ( .A(_abc_42016_n2231), .B(_abc_42016_n2335), .C(rdatahold_2_), .Y(_abc_42016_n2485) );
  OAI21X1 OAI21X1_563 ( .A(_abc_42016_n2237), .B(_abc_42016_n2462), .C(_abc_42016_n2485), .Y(rdatahold_2__FF_INPUT) );
  OAI21X1 OAI21X1_564 ( .A(_abc_42016_n2231), .B(_abc_42016_n2335), .C(rdatahold_3_), .Y(_abc_42016_n2487_1) );
  OAI21X1 OAI21X1_565 ( .A(_abc_42016_n2240), .B(_abc_42016_n2462), .C(_abc_42016_n2487_1), .Y(rdatahold_3__FF_INPUT) );
  OAI21X1 OAI21X1_566 ( .A(_abc_42016_n2231), .B(_abc_42016_n2335), .C(rdatahold_4_), .Y(_abc_42016_n2489) );
  OAI21X1 OAI21X1_567 ( .A(_abc_42016_n2243), .B(_abc_42016_n2462), .C(_abc_42016_n2489), .Y(rdatahold_4__FF_INPUT) );
  OAI21X1 OAI21X1_568 ( .A(_abc_42016_n2231), .B(_abc_42016_n2335), .C(rdatahold_6_), .Y(_abc_42016_n2492) );
  OAI21X1 OAI21X1_569 ( .A(_abc_42016_n2248), .B(_abc_42016_n2462), .C(_abc_42016_n2492), .Y(rdatahold_6__FF_INPUT) );
  OAI21X1 OAI21X1_57 ( .A(_abc_42016_n811), .B(_abc_42016_n587), .C(_abc_42016_n816), .Y(_abc_42016_n817) );
  OAI21X1 OAI21X1_570 ( .A(_abc_42016_n2231), .B(_abc_42016_n2335), .C(rdatahold_7_), .Y(_abc_42016_n2494) );
  OAI21X1 OAI21X1_571 ( .A(_abc_42016_n2250), .B(_abc_42016_n2462), .C(_abc_42016_n2494), .Y(rdatahold_7__FF_INPUT) );
  OAI21X1 OAI21X1_572 ( .A(_abc_42016_n511), .B(_abc_42016_n546), .C(_abc_42016_n2497), .Y(_abc_42016_n2498) );
  OAI21X1 OAI21X1_573 ( .A(_abc_42016_n2498), .B(_abc_42016_n2268), .C(_abc_42016_n529), .Y(_abc_42016_n2499) );
  OAI21X1 OAI21X1_574 ( .A(pc_0_), .B(_abc_42016_n2501), .C(_abc_42016_n2505), .Y(_abc_42016_n2506) );
  OAI21X1 OAI21X1_575 ( .A(_abc_42016_n2507), .B(_abc_42016_n2506), .C(_abc_42016_n673), .Y(_abc_42016_n2508) );
  OAI21X1 OAI21X1_576 ( .A(opcode_4_), .B(_abc_42016_n530), .C(regfil_7__0_), .Y(_abc_42016_n2510) );
  OAI21X1 OAI21X1_577 ( .A(_abc_42016_n695), .B(_abc_42016_n669), .C(_abc_42016_n2510), .Y(_abc_42016_n2511) );
  OAI21X1 OAI21X1_578 ( .A(_abc_42016_n2496), .B(_abc_42016_n2509), .C(_abc_42016_n2513), .Y(_abc_42016_n2514) );
  OAI21X1 OAI21X1_579 ( .A(wdatahold_0_), .B(_abc_42016_n1863), .C(_abc_42016_n547), .Y(_abc_42016_n2516) );
  OAI21X1 OAI21X1_58 ( .A(_abc_42016_n601), .B(_abc_42016_n819), .C(_abc_42016_n820), .Y(_abc_42016_n821) );
  OAI21X1 OAI21X1_580 ( .A(_abc_42016_n602), .B(_abc_42016_n2267), .C(_abc_42016_n2520), .Y(_abc_42016_n2521) );
  OAI21X1 OAI21X1_581 ( .A(_abc_42016_n2521), .B(_abc_42016_n2517_1), .C(_abc_42016_n2500), .Y(_abc_42016_n2522) );
  OAI21X1 OAI21X1_582 ( .A(_abc_42016_n2496), .B(_abc_42016_n2500), .C(_abc_42016_n2522), .Y(wdatahold_0__FF_INPUT) );
  OAI21X1 OAI21X1_583 ( .A(opcode_4_), .B(_abc_42016_n645), .C(_abc_42016_n2527), .Y(_abc_42016_n2528) );
  OAI21X1 OAI21X1_584 ( .A(opcode_5_), .B(_abc_42016_n2528), .C(_abc_42016_n2530), .Y(_abc_42016_n2531) );
  OAI21X1 OAI21X1_585 ( .A(_abc_42016_n709), .B(_abc_42016_n1061), .C(_abc_42016_n2531), .Y(_abc_42016_n2532) );
  OAI21X1 OAI21X1_586 ( .A(_abc_42016_n1383), .B(_abc_42016_n1405), .C(_abc_42016_n2533), .Y(_abc_42016_n2534) );
  OAI21X1 OAI21X1_587 ( .A(_abc_42016_n1409), .B(_abc_42016_n1377), .C(_abc_42016_n673), .Y(_abc_42016_n2536) );
  OAI21X1 OAI21X1_588 ( .A(_abc_42016_n2535), .B(_abc_42016_n2534), .C(_abc_42016_n2537), .Y(_abc_42016_n2538) );
  OAI21X1 OAI21X1_589 ( .A(opcode_6_), .B(_abc_42016_n1346), .C(_abc_42016_n2358), .Y(_abc_42016_n2540) );
  OAI21X1 OAI21X1_59 ( .A(regfil_3__2_), .B(_abc_42016_n782), .C(regfil_3__3_), .Y(_abc_42016_n827) );
  OAI21X1 OAI21X1_590 ( .A(_abc_42016_n2540), .B(_abc_42016_n2539), .C(wdatahold_1_), .Y(_abc_42016_n2541) );
  OAI21X1 OAI21X1_591 ( .A(regfil_7__1_), .B(_abc_42016_n668), .C(_abc_42016_n2543), .Y(_abc_42016_n2544) );
  OAI21X1 OAI21X1_592 ( .A(_abc_42016_n2542), .B(_abc_42016_n2544), .C(_abc_42016_n1863), .Y(_abc_42016_n2545) );
  OAI21X1 OAI21X1_593 ( .A(_abc_42016_n719), .B(_abc_42016_n2267), .C(_abc_42016_n2550), .Y(_abc_42016_n2551) );
  OAI21X1 OAI21X1_594 ( .A(_abc_42016_n2499), .B(_abc_42016_n2552), .C(_abc_42016_n2553), .Y(wdatahold_1__FF_INPUT) );
  OAI21X1 OAI21X1_595 ( .A(_abc_42016_n1675), .B(_abc_42016_n2267), .C(_abc_42016_n2556), .Y(_abc_42016_n2557) );
  OAI21X1 OAI21X1_596 ( .A(wdatahold_2_), .B(_abc_42016_n1863), .C(_abc_42016_n547), .Y(_abc_42016_n2558) );
  OAI21X1 OAI21X1_597 ( .A(_abc_42016_n1383), .B(_abc_42016_n1381), .C(_abc_42016_n1382), .Y(_abc_42016_n2560) );
  OAI21X1 OAI21X1_598 ( .A(_abc_42016_n531), .B(_abc_42016_n773), .C(_abc_42016_n1949), .Y(_abc_42016_n2564) );
  OAI21X1 OAI21X1_599 ( .A(_abc_42016_n2029), .B(_abc_42016_n1004), .C(_abc_42016_n2566), .Y(_abc_42016_n2567) );
  OAI21X1 OAI21X1_6 ( .A(_abc_42016_n569), .B(_abc_42016_n573), .C(_abc_42016_n570), .Y(_abc_42016_n574) );
  OAI21X1 OAI21X1_60 ( .A(rdatahold2_3_), .B(_abc_42016_n685), .C(_abc_42016_n694), .Y(_abc_42016_n832) );
  OAI21X1 OAI21X1_600 ( .A(_abc_42016_n2565), .B(_abc_42016_n2567), .C(_abc_42016_n1399), .Y(_abc_42016_n2568) );
  OAI21X1 OAI21X1_601 ( .A(_abc_42016_n1382), .B(_abc_42016_n1405), .C(_abc_42016_n2568), .Y(_abc_42016_n2569) );
  OAI21X1 OAI21X1_602 ( .A(_abc_42016_n2574), .B(_abc_42016_n2570), .C(_abc_42016_n2537), .Y(_abc_42016_n2575) );
  OAI21X1 OAI21X1_603 ( .A(_abc_42016_n1454), .B(_abc_42016_n668), .C(_abc_42016_n2566), .Y(_abc_42016_n2576) );
  OAI21X1 OAI21X1_604 ( .A(_abc_42016_n672_1), .B(opcode_6_), .C(_abc_42016_n2577), .Y(_abc_42016_n2578_1) );
  OAI21X1 OAI21X1_605 ( .A(_abc_42016_n2557), .B(_abc_42016_n2580), .C(_abc_42016_n2500), .Y(_abc_42016_n2581) );
  OAI21X1 OAI21X1_606 ( .A(_abc_42016_n674), .B(_abc_42016_n1411), .C(_abc_42016_n2509), .Y(_abc_42016_n2582) );
  OAI21X1 OAI21X1_607 ( .A(_abc_42016_n2555), .B(_abc_42016_n2585), .C(_abc_42016_n2581), .Y(wdatahold_2__FF_INPUT) );
  OAI21X1 OAI21X1_608 ( .A(_abc_42016_n1381), .B(_abc_42016_n1385), .C(_abc_42016_n2591), .Y(_abc_42016_n2592) );
  OAI21X1 OAI21X1_609 ( .A(_abc_42016_n573), .B(_abc_42016_n1399), .C(_abc_42016_n2593), .Y(_abc_42016_n2594) );
  OAI21X1 OAI21X1_61 ( .A(_abc_42016_n834), .B(_abc_42016_n815), .C(_abc_42016_n660), .Y(_abc_42016_n835) );
  OAI21X1 OAI21X1_610 ( .A(_abc_42016_n1380), .B(_abc_42016_n2592), .C(_abc_42016_n2594), .Y(_abc_42016_n2595) );
  OAI21X1 OAI21X1_611 ( .A(opcode_4_), .B(regfil_1__3_), .C(_abc_42016_n2596), .Y(_abc_42016_n2597) );
  OAI21X1 OAI21X1_612 ( .A(_abc_42016_n1357), .B(_abc_42016_n1405), .C(_abc_42016_n2599), .Y(_abc_42016_n2600) );
  OAI21X1 OAI21X1_613 ( .A(_abc_42016_n1378), .B(_abc_42016_n2590), .C(_abc_42016_n2601), .Y(_abc_42016_n2602) );
  OAI21X1 OAI21X1_614 ( .A(_abc_42016_n1488), .B(_abc_42016_n668), .C(_abc_42016_n2606), .Y(_abc_42016_n2607) );
  OAI21X1 OAI21X1_615 ( .A(_abc_42016_n2609_1), .B(_abc_42016_n2603), .C(_abc_42016_n2610), .Y(_abc_42016_n2611) );
  OAI21X1 OAI21X1_616 ( .A(_abc_42016_n2612), .B(_abc_42016_n2613), .C(_abc_42016_n2615), .Y(_abc_42016_n2616) );
  OAI21X1 OAI21X1_617 ( .A(opcode_4_), .B(regfil_1__4_), .C(_abc_42016_n2621), .Y(_abc_42016_n2622) );
  OAI21X1 OAI21X1_618 ( .A(_abc_42016_n2064), .B(_abc_42016_n1004), .C(_abc_42016_n2624), .Y(_abc_42016_n2625) );
  OAI21X1 OAI21X1_619 ( .A(_abc_42016_n2623), .B(_abc_42016_n2625), .C(_abc_42016_n1399), .Y(_abc_42016_n2626) );
  OAI21X1 OAI21X1_62 ( .A(regfil_0__3_), .B(_abc_42016_n748), .C(regfil_0__4_), .Y(_abc_42016_n839) );
  OAI21X1 OAI21X1_620 ( .A(_abc_42016_n1381), .B(_abc_42016_n1385), .C(_abc_42016_n1356), .Y(_abc_42016_n2631) );
  OAI21X1 OAI21X1_621 ( .A(_abc_42016_n1381), .B(_abc_42016_n2630), .C(_abc_42016_n2631), .Y(_abc_42016_n2632) );
  OAI21X1 OAI21X1_622 ( .A(_abc_42016_n1357), .B(_abc_42016_n1358), .C(_abc_42016_n1356), .Y(_abc_42016_n2634) );
  OAI21X1 OAI21X1_623 ( .A(_abc_42016_n2629), .B(_abc_42016_n2636), .C(_abc_42016_n2537), .Y(_abc_42016_n2637) );
  OAI21X1 OAI21X1_624 ( .A(_abc_42016_n2640_1), .B(_abc_42016_n2639_1), .C(_abc_42016_n1863), .Y(_abc_42016_n2641) );
  OAI21X1 OAI21X1_625 ( .A(_abc_42016_n2471), .B(_abc_42016_n2267), .C(_abc_42016_n2500), .Y(_abc_42016_n2645) );
  OAI21X1 OAI21X1_626 ( .A(_abc_42016_n1356), .B(_abc_42016_n1360), .C(_abc_42016_n2649), .Y(_abc_42016_n2650) );
  OAI21X1 OAI21X1_627 ( .A(_abc_42016_n1381), .B(_abc_42016_n2630), .C(_abc_42016_n2649), .Y(_abc_42016_n2652) );
  OAI21X1 OAI21X1_628 ( .A(_abc_42016_n1381), .B(_abc_42016_n1387), .C(_abc_42016_n2652), .Y(_abc_42016_n2653) );
  OAI21X1 OAI21X1_629 ( .A(opcode_4_), .B(_abc_42016_n642), .C(_abc_42016_n2654), .Y(_abc_42016_n2655) );
  OAI21X1 OAI21X1_63 ( .A(regfil_7__4_), .B(_abc_42016_n565), .C(opcode_2_), .Y(_abc_42016_n841) );
  OAI21X1 OAI21X1_630 ( .A(_abc_42016_n2649), .B(_abc_42016_n1405), .C(_abc_42016_n2656), .Y(_abc_42016_n2657) );
  OAI21X1 OAI21X1_631 ( .A(_abc_42016_n1380), .B(_abc_42016_n2653), .C(_abc_42016_n2658), .Y(_abc_42016_n2659) );
  OAI21X1 OAI21X1_632 ( .A(_abc_42016_n2540), .B(_abc_42016_n2539), .C(wdatahold_5_), .Y(_abc_42016_n2662) );
  OAI21X1 OAI21X1_633 ( .A(opcode_4_), .B(_abc_42016_n530), .C(_abc_42016_n898), .Y(_abc_42016_n2663) );
  OAI21X1 OAI21X1_634 ( .A(regfil_5__5_), .B(_abc_42016_n669), .C(_abc_42016_n2663), .Y(_abc_42016_n2664) );
  OAI21X1 OAI21X1_635 ( .A(_abc_42016_n2664), .B(_abc_42016_n2542), .C(_abc_42016_n1863), .Y(_abc_42016_n2665) );
  OAI21X1 OAI21X1_636 ( .A(_abc_42016_n2667), .B(_abc_42016_n2661), .C(_abc_42016_n2668), .Y(_abc_42016_n2669) );
  OAI21X1 OAI21X1_637 ( .A(_abc_42016_n1526), .B(_abc_42016_n2497), .C(_abc_42016_n2670), .Y(_abc_42016_n2671) );
  OAI21X1 OAI21X1_638 ( .A(_abc_42016_n1381), .B(_abc_42016_n1387), .C(_abc_42016_n1355), .Y(_abc_42016_n2675) );
  OAI21X1 OAI21X1_639 ( .A(_abc_42016_n1381), .B(_abc_42016_n2674), .C(_abc_42016_n2675), .Y(_abc_42016_n2676) );
  OAI21X1 OAI21X1_64 ( .A(regfil_6__4_), .B(_abc_42016_n539), .C(_abc_42016_n844), .Y(_abc_42016_n845) );
  OAI21X1 OAI21X1_640 ( .A(_abc_42016_n2050), .B(_abc_42016_n1004), .C(_abc_42016_n2680), .Y(_abc_42016_n2681) );
  OAI21X1 OAI21X1_641 ( .A(_abc_42016_n1355), .B(_abc_42016_n1405), .C(_abc_42016_n2683), .Y(_abc_42016_n2684) );
  OAI21X1 OAI21X1_642 ( .A(_abc_42016_n2649), .B(_abc_42016_n2633), .C(_abc_42016_n1355), .Y(_abc_42016_n2686) );
  OAI21X1 OAI21X1_643 ( .A(_abc_42016_n1378), .B(_abc_42016_n2688), .C(_abc_42016_n2685), .Y(_abc_42016_n2689) );
  OAI21X1 OAI21X1_644 ( .A(_abc_42016_n2677), .B(_abc_42016_n2689), .C(_abc_42016_n2537), .Y(_abc_42016_n2690) );
  OAI21X1 OAI21X1_645 ( .A(_abc_42016_n924), .B(_abc_42016_n668), .C(_abc_42016_n2680), .Y(_abc_42016_n2692) );
  OAI21X1 OAI21X1_646 ( .A(_abc_42016_n2695), .B(_abc_42016_n2613), .C(_abc_42016_n2696), .Y(_abc_42016_n2697) );
  OAI21X1 OAI21X1_647 ( .A(waddrhold_5_), .B(_abc_42016_n1863), .C(_abc_42016_n547), .Y(_abc_42016_n2701) );
  OAI21X1 OAI21X1_648 ( .A(_abc_42016_n2701), .B(_abc_42016_n2700), .C(_abc_42016_n2500), .Y(_abc_42016_n2702) );
  OAI21X1 OAI21X1_649 ( .A(wdatahold_7_), .B(_abc_42016_n1863), .C(_abc_42016_n547), .Y(_abc_42016_n2704) );
  OAI21X1 OAI21X1_65 ( .A(regfil_3__4_), .B(_abc_42016_n565), .C(_abc_42016_n536), .Y(_abc_42016_n846) );
  OAI21X1 OAI21X1_650 ( .A(_abc_42016_n2478), .B(_abc_42016_n2267), .C(_abc_42016_n2705), .Y(_abc_42016_n2706_1) );
  OAI21X1 OAI21X1_651 ( .A(opcode_4_), .B(_abc_42016_n530), .C(regfil_7__7_), .Y(_abc_42016_n2710) );
  OAI21X1 OAI21X1_652 ( .A(_abc_42016_n959), .B(_abc_42016_n669), .C(_abc_42016_n2710), .Y(_abc_42016_n2711_1) );
  OAI21X1 OAI21X1_653 ( .A(_abc_42016_n2709), .B(_abc_42016_n2509), .C(_abc_42016_n2712), .Y(_abc_42016_n2713) );
  OAI21X1 OAI21X1_654 ( .A(_abc_42016_n1381), .B(_abc_42016_n2674), .C(_abc_42016_n1354), .Y(_abc_42016_n2715) );
  OAI21X1 OAI21X1_655 ( .A(_abc_42016_n1381), .B(_abc_42016_n1389), .C(_abc_42016_n2715), .Y(_abc_42016_n2716) );
  OAI21X1 OAI21X1_656 ( .A(opcode_4_), .B(regfil_1__7_), .C(_abc_42016_n2717), .Y(_abc_42016_n2718) );
  OAI21X1 OAI21X1_657 ( .A(opcode_5_), .B(_abc_42016_n2718), .C(_abc_42016_n2719), .Y(_abc_42016_n2720) );
  OAI21X1 OAI21X1_658 ( .A(_abc_42016_n1354), .B(_abc_42016_n1405), .C(_abc_42016_n2721), .Y(_abc_42016_n2722) );
  OAI21X1 OAI21X1_659 ( .A(_abc_42016_n1355), .B(_abc_42016_n1362), .C(_abc_42016_n1354), .Y(_abc_42016_n2723) );
  OAI21X1 OAI21X1_66 ( .A(regfil_1__4_), .B(_abc_42016_n626), .C(_abc_42016_n848), .Y(_abc_42016_n849) );
  OAI21X1 OAI21X1_660 ( .A(_abc_42016_n1380), .B(_abc_42016_n2716), .C(_abc_42016_n2725), .Y(_abc_42016_n2726) );
  OAI21X1 OAI21X1_661 ( .A(_abc_42016_n2704), .B(_abc_42016_n2727), .C(_abc_42016_n2707), .Y(_abc_42016_n2728) );
  OAI21X1 OAI21X1_662 ( .A(opcode_0_), .B(_abc_42016_n536), .C(_abc_42016_n1374), .Y(_abc_42016_n2741) );
  OAI21X1 OAI21X1_663 ( .A(_abc_42016_n560), .B(_abc_42016_n2738), .C(_abc_42016_n2745), .Y(_abc_42016_n2746) );
  OAI21X1 OAI21X1_664 ( .A(regfil_5__0_), .B(_abc_42016_n2280), .C(_abc_42016_n1879_1), .Y(_abc_42016_n2748_1) );
  OAI21X1 OAI21X1_665 ( .A(_abc_42016_n560), .B(_abc_42016_n2748_1), .C(_abc_42016_n2747_1), .Y(_abc_42016_n2749) );
  OAI21X1 OAI21X1_666 ( .A(pc_0_), .B(_abc_42016_n2425), .C(_abc_42016_n2751), .Y(_abc_42016_n2752) );
  OAI21X1 OAI21X1_667 ( .A(_abc_42016_n2750), .B(_abc_42016_n2752), .C(_abc_42016_n2428), .Y(_abc_42016_n2753) );
  OAI21X1 OAI21X1_668 ( .A(_abc_42016_n695), .B(_abc_42016_n2754), .C(_abc_42016_n2753), .Y(_abc_42016_n2755) );
  OAI21X1 OAI21X1_669 ( .A(_abc_42016_n548), .B(_abc_42016_n2756), .C(_abc_42016_n2761), .Y(_abc_42016_n2762) );
  OAI21X1 OAI21X1_67 ( .A(regfil_3__4_), .B(_abc_42016_n600), .C(_abc_42016_n692), .Y(_abc_42016_n860) );
  OAI21X1 OAI21X1_670 ( .A(_abc_42016_n2731), .B(_abc_42016_n2736), .C(_abc_42016_n2763), .Y(raddrhold_0__FF_INPUT) );
  OAI21X1 OAI21X1_671 ( .A(regfil_5__1_), .B(_abc_42016_n2280), .C(_abc_42016_n1910), .Y(_abc_42016_n2766) );
  OAI21X1 OAI21X1_672 ( .A(_abc_42016_n2769), .B(_abc_42016_n2425), .C(_abc_42016_n2770), .Y(_abc_42016_n2771) );
  OAI21X1 OAI21X1_673 ( .A(_abc_42016_n2765), .B(_abc_42016_n2767_1), .C(_abc_42016_n2772), .Y(_abc_42016_n2773) );
  OAI21X1 OAI21X1_674 ( .A(_abc_42016_n2779), .B(_abc_42016_n2780), .C(_abc_42016_n2778), .Y(_abc_42016_n2781) );
  OAI21X1 OAI21X1_675 ( .A(raddrhold_2_), .B(_abc_42016_n2777), .C(_abc_42016_n2732), .Y(_abc_42016_n2789_1) );
  OAI21X1 OAI21X1_676 ( .A(_abc_42016_n2788_1), .B(_abc_42016_n2789_1), .C(_abc_42016_n2736), .Y(_abc_42016_n2790) );
  OAI21X1 OAI21X1_677 ( .A(regfil_5__2_), .B(_abc_42016_n2280), .C(_abc_42016_n1910), .Y(_abc_42016_n2792) );
  OAI21X1 OAI21X1_678 ( .A(_abc_42016_n757), .B(_abc_42016_n2429_1), .C(_abc_42016_n2795), .Y(_abc_42016_n2796) );
  OAI21X1 OAI21X1_679 ( .A(_abc_42016_n2794), .B(_abc_42016_n2796), .C(_abc_42016_n2428), .Y(_abc_42016_n2797) );
  OAI21X1 OAI21X1_68 ( .A(_abc_42016_n795), .B(_abc_42016_n775), .C(_abc_42016_n861), .Y(_abc_42016_n862) );
  OAI21X1 OAI21X1_680 ( .A(_abc_42016_n2800), .B(_abc_42016_n2793), .C(_abc_42016_n547), .Y(_abc_42016_n2801) );
  OAI21X1 OAI21X1_681 ( .A(raddrhold_3_), .B(_abc_42016_n2788_1), .C(_abc_42016_n2805), .Y(_abc_42016_n2806) );
  OAI21X1 OAI21X1_682 ( .A(_abc_42016_n1174_1), .B(_abc_42016_n2272), .C(_abc_42016_n2806), .Y(_abc_42016_n2807) );
  OAI21X1 OAI21X1_683 ( .A(_abc_42016_n2803), .B(_abc_42016_n2812), .C(_abc_42016_n2816), .Y(_abc_42016_n2817) );
  OAI21X1 OAI21X1_684 ( .A(_abc_42016_n2809), .B(_abc_42016_n2817), .C(_abc_42016_n547), .Y(_abc_42016_n2818) );
  OAI21X1 OAI21X1_685 ( .A(regfil_5__4_), .B(_abc_42016_n2280), .C(_abc_42016_n1910), .Y(_abc_42016_n2821) );
  OAI21X1 OAI21X1_686 ( .A(_abc_42016_n2823), .B(_abc_42016_n2824), .C(_abc_42016_n2428), .Y(_abc_42016_n2825) );
  OAI21X1 OAI21X1_687 ( .A(_abc_42016_n843), .B(_abc_42016_n2754), .C(_abc_42016_n2825), .Y(_abc_42016_n2826) );
  OAI21X1 OAI21X1_688 ( .A(_abc_42016_n2826), .B(_abc_42016_n2822), .C(_abc_42016_n547), .Y(_abc_42016_n2827) );
  OAI21X1 OAI21X1_689 ( .A(raddrhold_4_), .B(_abc_42016_n2804), .C(_abc_42016_n2732), .Y(_abc_42016_n2830) );
  OAI21X1 OAI21X1_69 ( .A(_abc_42016_n865), .B(_abc_42016_n866), .C(_abc_42016_n779), .Y(_abc_42016_n867_1) );
  OAI21X1 OAI21X1_690 ( .A(_abc_42016_n2839), .B(_abc_42016_n2746), .C(raddrhold_5_), .Y(_abc_42016_n2840) );
  OAI21X1 OAI21X1_691 ( .A(_abc_42016_n2653), .B(_abc_42016_n2425), .C(_abc_42016_n2842), .Y(_abc_42016_n2843) );
  OAI21X1 OAI21X1_692 ( .A(_abc_42016_n2837), .B(_abc_42016_n2845), .C(_abc_42016_n547), .Y(_abc_42016_n2846) );
  OAI21X1 OAI21X1_693 ( .A(raddrhold_5_), .B(_abc_42016_n2829), .C(_abc_42016_n2732), .Y(_abc_42016_n2848) );
  OAI21X1 OAI21X1_694 ( .A(_abc_42016_n2847), .B(_abc_42016_n2848), .C(_abc_42016_n2736), .Y(_abc_42016_n2849) );
  OAI21X1 OAI21X1_695 ( .A(raddrhold_6_), .B(_abc_42016_n2279), .C(_abc_42016_n2856_1), .Y(_abc_42016_n2857) );
  OAI21X1 OAI21X1_696 ( .A(_abc_42016_n2676), .B(_abc_42016_n2425), .C(_abc_42016_n2857), .Y(_abc_42016_n2858) );
  OAI21X1 OAI21X1_697 ( .A(_abc_42016_n2854), .B(_abc_42016_n2858), .C(_abc_42016_n2428), .Y(_abc_42016_n2859) );
  OAI21X1 OAI21X1_698 ( .A(_abc_42016_n923), .B(_abc_42016_n2754), .C(_abc_42016_n2859), .Y(_abc_42016_n2860) );
  OAI21X1 OAI21X1_699 ( .A(_abc_42016_n2860), .B(_abc_42016_n2853), .C(_abc_42016_n547), .Y(_abc_42016_n2861) );
  OAI21X1 OAI21X1_7 ( .A(_abc_42016_n562), .B(_abc_42016_n574), .C(_abc_42016_n587), .Y(_abc_42016_n588_1) );
  OAI21X1 OAI21X1_70 ( .A(_abc_42016_n860), .B(_abc_42016_n859), .C(_abc_42016_n870), .Y(_abc_36783_n3373) );
  OAI21X1 OAI21X1_700 ( .A(raddrhold_6_), .B(_abc_42016_n2847), .C(_abc_42016_n2862), .Y(_abc_42016_n2863) );
  OAI21X1 OAI21X1_701 ( .A(_abc_42016_n1261), .B(_abc_42016_n2272), .C(_abc_42016_n2863), .Y(_abc_42016_n2864) );
  OAI21X1 OAI21X1_702 ( .A(_abc_42016_n2870), .B(_abc_42016_n2737), .C(raddrhold_7_), .Y(_abc_42016_n2871) );
  OAI21X1 OAI21X1_703 ( .A(_abc_42016_n2869), .B(_abc_42016_n2745), .C(_abc_42016_n2877), .Y(_abc_42016_n2878_1) );
  OAI21X1 OAI21X1_704 ( .A(_abc_42016_n2875), .B(_abc_42016_n2878_1), .C(_abc_42016_n547), .Y(_abc_42016_n2879_1) );
  OAI21X1 OAI21X1_705 ( .A(_abc_42016_n1302), .B(_abc_42016_n2272), .C(_abc_42016_n2736), .Y(_abc_42016_n2884) );
  OAI21X1 OAI21X1_706 ( .A(raddrhold_8_), .B(_abc_42016_n2881), .C(_abc_42016_n2732), .Y(_abc_42016_n2889) );
  OAI21X1 OAI21X1_707 ( .A(_abc_42016_n2889), .B(_abc_42016_n2888), .C(_abc_42016_n2736), .Y(_abc_42016_n2890) );
  OAI21X1 OAI21X1_708 ( .A(_abc_42016_n1393), .B(_abc_42016_n2425), .C(_abc_42016_n2895), .Y(_abc_42016_n2896) );
  OAI21X1 OAI21X1_709 ( .A(_abc_42016_n629), .B(_abc_42016_n2754), .C(_abc_42016_n2898), .Y(_abc_42016_n2899) );
  OAI21X1 OAI21X1_71 ( .A(_abc_42016_n876), .B(_abc_42016_n878), .C(_abc_42016_n779), .Y(_abc_42016_n879) );
  OAI21X1 OAI21X1_710 ( .A(_abc_42016_n2899), .B(_abc_42016_n2892), .C(_abc_42016_n547), .Y(_abc_42016_n2900_1) );
  OAI21X1 OAI21X1_711 ( .A(raddrhold_9_), .B(_abc_42016_n2279), .C(_abc_42016_n1879_1), .Y(_abc_42016_n2904) );
  OAI21X1 OAI21X1_712 ( .A(_abc_42016_n2902), .B(_abc_42016_n2905), .C(_abc_42016_n2428), .Y(_abc_42016_n2906) );
  OAI21X1 OAI21X1_713 ( .A(_abc_42016_n2740), .B(_abc_42016_n2743), .C(_abc_42016_n673), .Y(_abc_42016_n2908) );
  OAI21X1 OAI21X1_714 ( .A(raddrhold_9_), .B(_abc_42016_n2888), .C(_abc_42016_n2732), .Y(_abc_42016_n2914) );
  OAI21X1 OAI21X1_715 ( .A(_abc_42016_n548), .B(_abc_42016_n2747_1), .C(_abc_42016_n2736), .Y(_abc_42016_n2917) );
  OAI21X1 OAI21X1_716 ( .A(_abc_42016_n2735), .B(_abc_42016_n2916), .C(_abc_42016_n2918), .Y(raddrhold_9__FF_INPUT) );
  OAI21X1 OAI21X1_717 ( .A(_abc_42016_n1841), .B(_abc_42016_n2285), .C(_abc_42016_n1467), .Y(_abc_42016_n2921) );
  OAI21X1 OAI21X1_718 ( .A(raddrhold_10_), .B(_abc_42016_n2279), .C(_abc_42016_n1879_1), .Y(_abc_42016_n2923) );
  OAI21X1 OAI21X1_719 ( .A(raddrhold_10_), .B(_abc_42016_n2738), .C(_abc_42016_n559), .Y(_abc_42016_n2926) );
  OAI21X1 OAI21X1_72 ( .A(_abc_42016_n772), .B(_abc_42016_n875), .C(_abc_42016_n880), .Y(_abc_42016_n881) );
  OAI21X1 OAI21X1_720 ( .A(_abc_42016_n2908), .B(_abc_42016_n2928), .C(_abc_42016_n2931), .Y(_abc_42016_n2932) );
  OAI21X1 OAI21X1_721 ( .A(_abc_42016_n2927), .B(_abc_42016_n2932), .C(_abc_42016_n547), .Y(_abc_42016_n2933) );
  OAI21X1 OAI21X1_722 ( .A(_abc_42016_n1675), .B(_abc_42016_n2272), .C(_abc_42016_n2736), .Y(_abc_42016_n2937) );
  OAI21X1 OAI21X1_723 ( .A(_abc_42016_n1371), .B(_abc_42016_n1376), .C(_abc_42016_n2944), .Y(_abc_42016_n2945) );
  OAI21X1 OAI21X1_724 ( .A(_abc_42016_n1489), .B(_abc_42016_n2291), .C(_abc_42016_n2945), .Y(_abc_42016_n2946_1) );
  OAI21X1 OAI21X1_725 ( .A(_abc_42016_n2946_1), .B(_abc_42016_n2941), .C(_abc_42016_n2428), .Y(_abc_42016_n2947_1) );
  OAI21X1 OAI21X1_726 ( .A(raddrhold_11_), .B(_abc_42016_n2934), .C(_abc_42016_n2732), .Y(_abc_42016_n2952) );
  OAI21X1 OAI21X1_727 ( .A(_abc_42016_n2953), .B(_abc_42016_n2950), .C(_abc_42016_n2736), .Y(_abc_42016_n2954) );
  OAI21X1 OAI21X1_728 ( .A(_abc_42016_n530), .B(_abc_42016_n533), .C(_abc_42016_n2956), .Y(_abc_42016_n2958) );
  OAI21X1 OAI21X1_729 ( .A(_abc_42016_n1515), .B(_abc_42016_n2310), .C(_abc_42016_n2959), .Y(_abc_42016_n2960) );
  OAI21X1 OAI21X1_73 ( .A(regfil_0__4_), .B(_abc_42016_n790), .C(regfil_0__5_), .Y(_abc_42016_n889_1) );
  OAI21X1 OAI21X1_730 ( .A(_abc_42016_n2908), .B(_abc_42016_n2963), .C(_abc_42016_n2964), .Y(_abc_42016_n2965) );
  OAI21X1 OAI21X1_731 ( .A(_abc_42016_n2962), .B(_abc_42016_n2965), .C(_abc_42016_n547), .Y(_abc_42016_n2966) );
  OAI21X1 OAI21X1_732 ( .A(raddrhold_12_), .B(_abc_42016_n2951), .C(_abc_42016_n2732), .Y(_abc_42016_n2967) );
  OAI21X1 OAI21X1_733 ( .A(_abc_42016_n2471), .B(_abc_42016_n2272), .C(_abc_42016_n2736), .Y(_abc_42016_n2969_1) );
  OAI21X1 OAI21X1_734 ( .A(raddrhold_13_), .B(_abc_42016_n2279), .C(_abc_42016_n1879_1), .Y(_abc_42016_n2974) );
  OAI21X1 OAI21X1_735 ( .A(_abc_42016_n1535), .B(_abc_42016_n2310), .C(_abc_42016_n2976), .Y(_abc_42016_n2977) );
  OAI21X1 OAI21X1_736 ( .A(_abc_42016_n2908), .B(_abc_42016_n2979), .C(_abc_42016_n2980), .Y(_abc_42016_n2981) );
  OAI21X1 OAI21X1_737 ( .A(_abc_42016_n2981), .B(_abc_42016_n2978), .C(_abc_42016_n547), .Y(_abc_42016_n2982) );
  OAI21X1 OAI21X1_738 ( .A(_abc_42016_n891), .B(_abc_42016_n2272), .C(_abc_42016_n2736), .Y(_abc_42016_n2987) );
  OAI21X1 OAI21X1_739 ( .A(raddrhold_14_), .B(_abc_42016_n2279), .C(_abc_42016_n2993), .Y(_abc_42016_n2994) );
  OAI21X1 OAI21X1_74 ( .A(_abc_42016_n894), .B(_abc_42016_n896), .C(_abc_42016_n536), .Y(_abc_42016_n897) );
  OAI21X1 OAI21X1_740 ( .A(_abc_42016_n1573), .B(_abc_42016_n2310), .C(_abc_42016_n2994), .Y(_abc_42016_n2995) );
  OAI21X1 OAI21X1_741 ( .A(_abc_42016_n2425), .B(_abc_42016_n1564), .C(_abc_42016_n2996), .Y(_abc_42016_n2997) );
  OAI21X1 OAI21X1_742 ( .A(raddrhold_14_), .B(_abc_42016_n2738), .C(_abc_42016_n559), .Y(_abc_42016_n2998) );
  OAI21X1 OAI21X1_743 ( .A(_abc_42016_n2908), .B(_abc_42016_n2992), .C(_abc_42016_n3000), .Y(_abc_42016_n3001) );
  OAI21X1 OAI21X1_744 ( .A(_abc_42016_n2991_1), .B(_abc_42016_n3001), .C(_abc_42016_n547), .Y(_abc_42016_n3002) );
  OAI21X1 OAI21X1_745 ( .A(_abc_42016_n1793), .B(_abc_42016_n2272), .C(_abc_42016_n2736), .Y(_abc_42016_n3006) );
  OAI21X1 OAI21X1_746 ( .A(raddrhold_15_), .B(_abc_42016_n2279), .C(_abc_42016_n1879_1), .Y(_abc_42016_n3011) );
  OAI21X1 OAI21X1_747 ( .A(_abc_42016_n2425), .B(_abc_42016_n1587), .C(_abc_42016_n3013), .Y(_abc_42016_n3014_1) );
  OAI21X1 OAI21X1_748 ( .A(raddrhold_15_), .B(_abc_42016_n2738), .C(_abc_42016_n559), .Y(_abc_42016_n3015_1) );
  OAI21X1 OAI21X1_749 ( .A(_abc_42016_n3012), .B(_abc_42016_n3014_1), .C(_abc_42016_n3016), .Y(_abc_42016_n3017) );
  OAI21X1 OAI21X1_75 ( .A(regfil_4__5_), .B(_abc_42016_n727), .C(opcode_2_), .Y(_abc_42016_n899) );
  OAI21X1 OAI21X1_750 ( .A(_abc_42016_n3018), .B(_abc_42016_n3019), .C(_abc_42016_n2909), .Y(_abc_42016_n3020) );
  OAI21X1 OAI21X1_751 ( .A(_abc_42016_n3023), .B(_abc_42016_n3003), .C(_abc_42016_n3024), .Y(_abc_42016_n3025) );
  OAI21X1 OAI21X1_752 ( .A(_abc_42016_n3036_1), .B(_abc_42016_n3035_1), .C(_abc_42016_n559), .Y(_abc_42016_n3037) );
  OAI21X1 OAI21X1_753 ( .A(_abc_42016_n560), .B(_abc_42016_n1848), .C(_abc_42016_n542), .Y(_abc_42016_n3040) );
  OAI21X1 OAI21X1_754 ( .A(_abc_42016_n3042), .B(_abc_42016_n3032), .C(_abc_42016_n3043), .Y(_abc_42016_n3044) );
  OAI21X1 OAI21X1_755 ( .A(_abc_42016_n695), .B(_abc_42016_n2613), .C(_abc_42016_n3046), .Y(_abc_42016_n3047) );
  OAI21X1 OAI21X1_756 ( .A(_abc_42016_n669), .B(_abc_42016_n682), .C(sp_1_), .Y(_abc_42016_n3051) );
  OAI21X1 OAI21X1_757 ( .A(_abc_42016_n536), .B(_abc_42016_n727), .C(_abc_42016_n1380), .Y(_abc_42016_n3054) );
  OAI21X1 OAI21X1_758 ( .A(sp_1_), .B(_abc_42016_n3056), .C(_abc_42016_n3051), .Y(_abc_42016_n3057_1) );
  OAI21X1 OAI21X1_759 ( .A(_abc_42016_n3050), .B(_abc_42016_n1411), .C(_abc_42016_n3057_1), .Y(_abc_42016_n3058_1) );
  OAI21X1 OAI21X1_76 ( .A(regfil_5__5_), .B(_abc_42016_n626), .C(_abc_42016_n900), .Y(_abc_42016_n901) );
  OAI21X1 OAI21X1_760 ( .A(regfil_5__1_), .B(_abc_42016_n2280), .C(_abc_42016_n1841), .Y(_abc_42016_n3060) );
  OAI21X1 OAI21X1_761 ( .A(_abc_42016_n3050), .B(_abc_42016_n2293), .C(_abc_42016_n3062), .Y(_abc_42016_n3063) );
  OAI21X1 OAI21X1_762 ( .A(_abc_42016_n3061), .B(_abc_42016_n3063), .C(_abc_42016_n559), .Y(_abc_42016_n3064) );
  OAI21X1 OAI21X1_763 ( .A(_abc_42016_n709), .B(_abc_42016_n2298), .C(_abc_42016_n3064), .Y(_abc_42016_n3065) );
  OAI21X1 OAI21X1_764 ( .A(_abc_42016_n3050), .B(_abc_42016_n2358), .C(_abc_42016_n3066), .Y(_abc_42016_n3067) );
  OAI21X1 OAI21X1_765 ( .A(_abc_42016_n3067), .B(_abc_42016_n3059), .C(_abc_42016_n3068), .Y(_abc_42016_n3069) );
  OAI21X1 OAI21X1_766 ( .A(waddrhold_0_), .B(waddrhold_1_), .C(_abc_42016_n2519), .Y(_abc_42016_n3074) );
  OAI21X1 OAI21X1_767 ( .A(_abc_42016_n3073), .B(_abc_42016_n3074), .C(_abc_42016_n3072), .Y(_abc_42016_n3075) );
  OAI21X1 OAI21X1_768 ( .A(_abc_42016_n2701), .B(_abc_42016_n2700), .C(_abc_42016_n3072), .Y(_abc_42016_n3079) );
  OAI21X1 OAI21X1_769 ( .A(waddrhold_2_), .B(_abc_42016_n3073), .C(_abc_42016_n2519), .Y(_abc_42016_n3084) );
  OAI21X1 OAI21X1_77 ( .A(_abc_42016_n892), .B(_abc_42016_n901), .C(_abc_42016_n897), .Y(_abc_42016_n902) );
  OAI21X1 OAI21X1_770 ( .A(_abc_42016_n3083), .B(_abc_42016_n3084), .C(_abc_42016_n3085), .Y(_abc_42016_n3086) );
  OAI21X1 OAI21X1_771 ( .A(waddrhold_2_), .B(_abc_42016_n1848), .C(_abc_42016_n541), .Y(_abc_42016_n3094) );
  OAI21X1 OAI21X1_772 ( .A(_abc_42016_n3094), .B(_abc_42016_n3093), .C(_abc_42016_n1863), .Y(_abc_42016_n3095) );
  OAI21X1 OAI21X1_773 ( .A(_abc_42016_n674), .B(_abc_42016_n3101), .C(_abc_42016_n3096), .Y(_abc_42016_n3102) );
  OAI21X1 OAI21X1_774 ( .A(waddrhold_3_), .B(_abc_42016_n3083), .C(_abc_42016_n2519), .Y(_abc_42016_n3108) );
  OAI21X1 OAI21X1_775 ( .A(_abc_42016_n3107), .B(_abc_42016_n3108), .C(_abc_42016_n3109), .Y(_abc_42016_n3110) );
  OAI21X1 OAI21X1_776 ( .A(waddrhold_3_), .B(_abc_42016_n2279), .C(_abc_42016_n2811_1), .Y(_abc_42016_n3112) );
  OAI21X1 OAI21X1_777 ( .A(_abc_42016_n3111), .B(_abc_42016_n3113), .C(_abc_42016_n559), .Y(_abc_42016_n3114) );
  OAI21X1 OAI21X1_778 ( .A(waddrhold_3_), .B(_abc_42016_n1848), .C(_abc_42016_n541), .Y(_abc_42016_n3116) );
  OAI21X1 OAI21X1_779 ( .A(_abc_42016_n3115), .B(_abc_42016_n3116), .C(_abc_42016_n3114), .Y(_abc_42016_n3117) );
  OAI21X1 OAI21X1_78 ( .A(_abc_42016_n891), .B(_abc_42016_n527), .C(_abc_42016_n904), .Y(_abc_42016_n905) );
  OAI21X1 OAI21X1_780 ( .A(sp_1_), .B(sp_2_), .C(sp_3_), .Y(_abc_42016_n3122) );
  OAI21X1 OAI21X1_781 ( .A(_abc_42016_n674), .B(_abc_42016_n3124), .C(_abc_42016_n3118), .Y(_abc_42016_n3125_1) );
  OAI21X1 OAI21X1_782 ( .A(sp_3_), .B(_abc_42016_n3119), .C(sp_4_), .Y(_abc_42016_n3132) );
  OAI21X1 OAI21X1_783 ( .A(_abc_42016_n3135), .B(_abc_42016_n3129), .C(_abc_42016_n673), .Y(_abc_42016_n3136) );
  OAI21X1 OAI21X1_784 ( .A(_abc_42016_n843), .B(_abc_42016_n2298), .C(_abc_42016_n3141), .Y(_abc_42016_n3142) );
  OAI21X1 OAI21X1_785 ( .A(waddrhold_4_), .B(_abc_42016_n1863), .C(_abc_42016_n547), .Y(_abc_42016_n3144) );
  OAI21X1 OAI21X1_786 ( .A(waddrhold_4_), .B(_abc_42016_n3107), .C(_abc_42016_n2519), .Y(_abc_42016_n3148_1) );
  OAI21X1 OAI21X1_787 ( .A(_abc_42016_n3147_1), .B(_abc_42016_n3148_1), .C(_abc_42016_n3149), .Y(_abc_42016_n3150) );
  OAI21X1 OAI21X1_788 ( .A(_abc_42016_n3150), .B(_abc_42016_n3145), .C(_abc_42016_n3072), .Y(_abc_42016_n3151) );
  OAI21X1 OAI21X1_789 ( .A(_abc_42016_n3128), .B(_abc_42016_n3072), .C(_abc_42016_n3151), .Y(waddrhold_4__FF_INPUT) );
  OAI21X1 OAI21X1_79 ( .A(_abc_42016_n903), .B(_abc_42016_n905), .C(_abc_42016_n720), .Y(_abc_42016_n906) );
  OAI21X1 OAI21X1_790 ( .A(_abc_42016_n3153), .B(_abc_42016_n2293), .C(_abc_42016_n3155), .Y(_abc_42016_n3156) );
  OAI21X1 OAI21X1_791 ( .A(waddrhold_5_), .B(_abc_42016_n1848), .C(_abc_42016_n541), .Y(_abc_42016_n3159) );
  OAI21X1 OAI21X1_792 ( .A(_abc_42016_n3158), .B(_abc_42016_n3159), .C(_abc_42016_n3157), .Y(_abc_42016_n3160) );
  OAI21X1 OAI21X1_793 ( .A(_abc_42016_n3166), .B(_abc_42016_n3165), .C(_abc_42016_n673), .Y(_abc_42016_n3167) );
  OAI21X1 OAI21X1_794 ( .A(waddrhold_5_), .B(_abc_42016_n3147_1), .C(_abc_42016_n2519), .Y(_abc_42016_n3171) );
  OAI21X1 OAI21X1_795 ( .A(_abc_42016_n3170_1), .B(_abc_42016_n3171), .C(_abc_42016_n3169_1), .Y(_abc_42016_n3172) );
  OAI21X1 OAI21X1_796 ( .A(_abc_42016_n3172), .B(_abc_42016_n3168), .C(_abc_42016_n3072), .Y(_abc_42016_n3173) );
  OAI21X1 OAI21X1_797 ( .A(_abc_42016_n3153), .B(_abc_42016_n3080_1), .C(_abc_42016_n3173), .Y(waddrhold_5__FF_INPUT) );
  OAI21X1 OAI21X1_798 ( .A(sp_5_), .B(_abc_42016_n3131), .C(sp_6_), .Y(_abc_42016_n3181) );
  OAI21X1 OAI21X1_799 ( .A(_abc_42016_n3183), .B(_abc_42016_n3176), .C(_abc_42016_n673), .Y(_abc_42016_n3184) );
  OAI21X1 OAI21X1_8 ( .A(_abc_42016_n552), .B(_abc_42016_n526_1), .C(_abc_42016_n589), .Y(_abc_42016_n590) );
  OAI21X1 OAI21X1_80 ( .A(_abc_42016_n891), .B(_abc_42016_n587), .C(_abc_42016_n906), .Y(_abc_42016_n907) );
  OAI21X1 OAI21X1_800 ( .A(_abc_42016_n923), .B(_abc_42016_n2298), .C(_abc_42016_n3189), .Y(_abc_42016_n3190) );
  OAI21X1 OAI21X1_801 ( .A(waddrhold_6_), .B(_abc_42016_n1863), .C(_abc_42016_n547), .Y(_abc_42016_n3192) );
  OAI21X1 OAI21X1_802 ( .A(waddrhold_6_), .B(_abc_42016_n3170_1), .C(_abc_42016_n2519), .Y(_abc_42016_n3196_1) );
  OAI21X1 OAI21X1_803 ( .A(_abc_42016_n3196_1), .B(_abc_42016_n3195_1), .C(_abc_42016_n3197), .Y(_abc_42016_n3198) );
  OAI21X1 OAI21X1_804 ( .A(_abc_42016_n3198), .B(_abc_42016_n3193), .C(_abc_42016_n3072), .Y(_abc_42016_n3199) );
  OAI21X1 OAI21X1_805 ( .A(_abc_42016_n3175), .B(_abc_42016_n3072), .C(_abc_42016_n3199), .Y(waddrhold_6__FF_INPUT) );
  OAI21X1 OAI21X1_806 ( .A(_abc_42016_n3202), .B(_abc_42016_n3203), .C(_abc_42016_n3056), .Y(_abc_42016_n3204) );
  OAI21X1 OAI21X1_807 ( .A(waddrhold_7_), .B(_abc_42016_n2279), .C(_abc_42016_n3208), .Y(_abc_42016_n3209) );
  OAI21X1 OAI21X1_808 ( .A(_abc_42016_n3201), .B(_abc_42016_n2293), .C(_abc_42016_n3209), .Y(_abc_42016_n3210) );
  OAI21X1 OAI21X1_809 ( .A(_abc_42016_n3207), .B(_abc_42016_n3210), .C(_abc_42016_n559), .Y(_abc_42016_n3211) );
  OAI21X1 OAI21X1_81 ( .A(_abc_42016_n884), .B(_abc_42016_n886), .C(_abc_42016_n908), .Y(_abc_42016_n909) );
  OAI21X1 OAI21X1_810 ( .A(_abc_42016_n3213), .B(_abc_42016_n3206), .C(_abc_42016_n3214), .Y(_abc_42016_n3215) );
  OAI21X1 OAI21X1_811 ( .A(_abc_42016_n1302), .B(_abc_42016_n2261), .C(_abc_42016_n3219), .Y(_abc_42016_n3220) );
  OAI21X1 OAI21X1_812 ( .A(_abc_42016_n3226), .B(_abc_42016_n3225), .C(_abc_42016_n3056), .Y(_abc_42016_n3227) );
  OAI21X1 OAI21X1_813 ( .A(waddrhold_8_), .B(_abc_42016_n2279), .C(_abc_42016_n2893), .Y(_abc_42016_n3231) );
  OAI21X1 OAI21X1_814 ( .A(_abc_42016_n3232), .B(_abc_42016_n3230), .C(_abc_42016_n559), .Y(_abc_42016_n3233) );
  OAI21X1 OAI21X1_815 ( .A(_abc_42016_n3235), .B(_abc_42016_n3229), .C(_abc_42016_n3236), .Y(_abc_42016_n3237) );
  OAI21X1 OAI21X1_816 ( .A(_abc_42016_n3245_1), .B(_abc_42016_n2293), .C(_abc_42016_n3253), .Y(_abc_42016_n3254) );
  OAI21X1 OAI21X1_817 ( .A(_abc_42016_n3255), .B(_abc_42016_n3254), .C(_abc_42016_n559), .Y(_abc_42016_n3256) );
  OAI21X1 OAI21X1_818 ( .A(_abc_42016_n1841), .B(_abc_42016_n3252), .C(_abc_42016_n3257), .Y(_abc_42016_n3258) );
  OAI21X1 OAI21X1_819 ( .A(_abc_42016_n674), .B(_abc_42016_n3251), .C(_abc_42016_n3259), .Y(_abc_42016_n3260) );
  OAI21X1 OAI21X1_82 ( .A(regfil_3__5_), .B(_abc_42016_n600), .C(_abc_42016_n692), .Y(_abc_42016_n911) );
  OAI21X1 OAI21X1_820 ( .A(_abc_42016_n1851), .B(_abc_42016_n3260), .C(_abc_42016_n3246), .Y(_abc_42016_n3261) );
  OAI21X1 OAI21X1_821 ( .A(_abc_42016_n719), .B(_abc_42016_n2261), .C(_abc_42016_n3262), .Y(_abc_42016_n3263) );
  OAI21X1 OAI21X1_822 ( .A(sp_9_), .B(_abc_42016_n3224), .C(sp_10_), .Y(_abc_42016_n3270) );
  OAI21X1 OAI21X1_823 ( .A(_abc_42016_n3130), .B(_abc_42016_n3271), .C(_abc_42016_n3272), .Y(_abc_42016_n3273) );
  OAI21X1 OAI21X1_824 ( .A(waddrhold_10_), .B(_abc_42016_n2279), .C(_abc_42016_n3276), .Y(_abc_42016_n3277) );
  OAI21X1 OAI21X1_825 ( .A(_abc_42016_n3268), .B(_abc_42016_n2293), .C(_abc_42016_n3277), .Y(_abc_42016_n3278) );
  OAI21X1 OAI21X1_826 ( .A(_abc_42016_n3275), .B(_abc_42016_n3278), .C(_abc_42016_n559), .Y(_abc_42016_n3279) );
  OAI21X1 OAI21X1_827 ( .A(_abc_42016_n3281), .B(_abc_42016_n3274), .C(_abc_42016_n3282), .Y(_abc_42016_n3283) );
  OAI21X1 OAI21X1_828 ( .A(_abc_42016_n3245_1), .B(_abc_42016_n3239), .C(_abc_42016_n3268), .Y(_abc_42016_n3284) );
  OAI21X1 OAI21X1_829 ( .A(_abc_42016_n1675), .B(_abc_42016_n2261), .C(_abc_42016_n3287), .Y(_abc_42016_n3288) );
  OAI21X1 OAI21X1_83 ( .A(_abc_42016_n911), .B(_abc_42016_n910_1), .C(_abc_42016_n882), .Y(_abc_36783_n3376) );
  OAI21X1 OAI21X1_830 ( .A(sp_10_), .B(_abc_42016_n3293), .C(sp_11_), .Y(_abc_42016_n3294) );
  OAI21X1 OAI21X1_831 ( .A(_abc_42016_n3130), .B(_abc_42016_n3298), .C(_abc_42016_n3299), .Y(_abc_42016_n3300) );
  OAI21X1 OAI21X1_832 ( .A(waddrhold_11_), .B(_abc_42016_n2279), .C(_abc_42016_n3301), .Y(_abc_42016_n3302) );
  OAI21X1 OAI21X1_833 ( .A(_abc_42016_n1347), .B(_abc_42016_n1489), .C(_abc_42016_n3302), .Y(_abc_42016_n3303) );
  OAI21X1 OAI21X1_834 ( .A(waddrhold_11_), .B(_abc_42016_n3285), .C(_abc_42016_n2519), .Y(_abc_42016_n3311) );
  OAI21X1 OAI21X1_835 ( .A(_abc_42016_n3311), .B(_abc_42016_n3310), .C(_abc_42016_n3312), .Y(_abc_42016_n3313) );
  OAI21X1 OAI21X1_836 ( .A(_abc_42016_n3316), .B(_abc_42016_n3309), .C(_abc_42016_n3317), .Y(_abc_42016_n3318_1) );
  OAI21X1 OAI21X1_837 ( .A(sp_11_), .B(_abc_42016_n3269), .C(sp_12_), .Y(_abc_42016_n3320) );
  OAI21X1 OAI21X1_838 ( .A(_abc_42016_n3130), .B(_abc_42016_n3321), .C(_abc_42016_n3322), .Y(_abc_42016_n3323) );
  OAI21X1 OAI21X1_839 ( .A(_abc_42016_n3326), .B(_abc_42016_n3327), .C(_abc_42016_n3325), .Y(_abc_42016_n3328) );
  OAI21X1 OAI21X1_84 ( .A(regfil_0__5_), .B(_abc_42016_n838), .C(regfil_0__6_), .Y(_abc_42016_n915) );
  OAI21X1 OAI21X1_840 ( .A(_abc_42016_n842), .B(_abc_42016_n2613), .C(_abc_42016_n3333), .Y(_abc_42016_n3334) );
  OAI21X1 OAI21X1_841 ( .A(sp_12_), .B(_abc_42016_n3296_1), .C(sp_13_), .Y(_abc_42016_n3338) );
  OAI21X1 OAI21X1_842 ( .A(_abc_42016_n3337), .B(_abc_42016_n1411), .C(_abc_42016_n3342), .Y(_abc_42016_n3343) );
  OAI21X1 OAI21X1_843 ( .A(waddrhold_13_), .B(_abc_42016_n2293), .C(_abc_42016_n559), .Y(_abc_42016_n3345_1) );
  OAI21X1 OAI21X1_844 ( .A(regfil_4__5_), .B(_abc_42016_n2280), .C(_abc_42016_n1841), .Y(_abc_42016_n3346_1) );
  OAI21X1 OAI21X1_845 ( .A(_abc_42016_n1527), .B(_abc_42016_n2298), .C(_abc_42016_n1863), .Y(_abc_42016_n3349) );
  OAI21X1 OAI21X1_846 ( .A(_abc_42016_n3345_1), .B(_abc_42016_n3348), .C(_abc_42016_n3350), .Y(_abc_42016_n3351) );
  OAI21X1 OAI21X1_847 ( .A(_abc_42016_n3351), .B(_abc_42016_n3344), .C(_abc_42016_n3352), .Y(_abc_42016_n3353) );
  OAI21X1 OAI21X1_848 ( .A(waddrhold_13_), .B(_abc_42016_n3354), .C(_abc_42016_n2519), .Y(_abc_42016_n3355) );
  OAI21X1 OAI21X1_849 ( .A(_abc_42016_n891), .B(_abc_42016_n2261), .C(_abc_42016_n3357), .Y(_abc_42016_n3358) );
  OAI21X1 OAI21X1_85 ( .A(regfil_6__6_), .B(_abc_42016_n539), .C(opcode_2_), .Y(_abc_42016_n922) );
  OAI21X1 OAI21X1_850 ( .A(sp_13_), .B(_abc_42016_n3319_1), .C(sp_14_), .Y(_abc_42016_n3364) );
  OAI21X1 OAI21X1_851 ( .A(_abc_42016_n3130), .B(_abc_42016_n3366), .C(_abc_42016_n3367), .Y(_abc_42016_n3368_1) );
  OAI21X1 OAI21X1_852 ( .A(waddrhold_14_), .B(_abc_42016_n2293), .C(_abc_42016_n559), .Y(_abc_42016_n3370) );
  OAI21X1 OAI21X1_853 ( .A(regfil_4__6_), .B(_abc_42016_n2280), .C(_abc_42016_n1841), .Y(_abc_42016_n3372) );
  OAI21X1 OAI21X1_854 ( .A(_abc_42016_n1554), .B(_abc_42016_n2298), .C(_abc_42016_n1863), .Y(_abc_42016_n3375) );
  OAI21X1 OAI21X1_855 ( .A(_abc_42016_n3370), .B(_abc_42016_n3374), .C(_abc_42016_n3376), .Y(_abc_42016_n3377) );
  OAI21X1 OAI21X1_856 ( .A(_abc_42016_n3377), .B(_abc_42016_n3369_1), .C(_abc_42016_n3378), .Y(_abc_42016_n3379) );
  OAI21X1 OAI21X1_857 ( .A(_abc_42016_n1793), .B(_abc_42016_n2261), .C(_abc_42016_n3384), .Y(_abc_42016_n3385) );
  OAI21X1 OAI21X1_858 ( .A(opcode_7_), .B(_abc_42016_n3397_1), .C(_abc_42016_n540), .Y(_abc_42016_n3398_1) );
  OAI21X1 OAI21X1_859 ( .A(_abc_42016_n3399), .B(_abc_42016_n3392), .C(_abc_42016_n3400), .Y(_abc_42016_n3401) );
  OAI21X1 OAI21X1_86 ( .A(regfil_4__6_), .B(_abc_42016_n727), .C(_abc_42016_n925), .Y(_abc_42016_n926) );
  OAI21X1 OAI21X1_860 ( .A(_abc_42016_n1801_1), .B(_abc_42016_n2613), .C(_abc_42016_n3402), .Y(_abc_42016_n3403) );
  OAI21X1 OAI21X1_861 ( .A(_abc_42016_n2519), .B(_abc_42016_n3410), .C(_abc_42016_n529), .Y(_abc_42016_n3411) );
  OAI21X1 OAI21X1_862 ( .A(_abc_42016_n2496), .B(_abc_42016_n3408), .C(_abc_42016_n3412), .Y(datao_0__FF_INPUT) );
  OAI21X1 OAI21X1_863 ( .A(_abc_42016_n2548_1), .B(_abc_42016_n3408), .C(_abc_42016_n3414), .Y(datao_1__FF_INPUT) );
  OAI21X1 OAI21X1_864 ( .A(_abc_42016_n2555), .B(_abc_42016_n3408), .C(_abc_42016_n3416), .Y(datao_2__FF_INPUT) );
  OAI21X1 OAI21X1_865 ( .A(_abc_42016_n1488), .B(_abc_42016_n3418), .C(_abc_42016_n3419), .Y(datao_3__FF_INPUT) );
  OAI21X1 OAI21X1_866 ( .A(_abc_42016_n2619), .B(_abc_42016_n3408), .C(_abc_42016_n3421_1), .Y(datao_4__FF_INPUT) );
  OAI21X1 OAI21X1_867 ( .A(_abc_42016_n2648), .B(_abc_42016_n3408), .C(_abc_42016_n3423), .Y(datao_5__FF_INPUT) );
  OAI21X1 OAI21X1_868 ( .A(_abc_42016_n924), .B(_abc_42016_n3418), .C(_abc_42016_n3425), .Y(datao_6__FF_INPUT) );
  OAI21X1 OAI21X1_869 ( .A(_abc_42016_n2709), .B(_abc_42016_n3408), .C(_abc_42016_n3427), .Y(datao_7__FF_INPUT) );
  OAI21X1 OAI21X1_87 ( .A(_abc_42016_n913), .B(_abc_42016_n885), .C(_abc_42016_n660), .Y(_abc_42016_n931) );
  OAI21X1 OAI21X1_870 ( .A(_abc_42016_n563), .B(_abc_42016_n537_1), .C(opcode_2_), .Y(_abc_42016_n3431) );
  OAI21X1 OAI21X1_871 ( .A(_abc_42016_n668), .B(_abc_42016_n2291), .C(_abc_42016_n3431), .Y(_abc_42016_n3432) );
  OAI21X1 OAI21X1_872 ( .A(regd_0_), .B(_abc_42016_n3432), .C(_abc_42016_n3434), .Y(_abc_42016_n3435) );
  OAI21X1 OAI21X1_873 ( .A(_abc_42016_n2370), .B(_abc_42016_n1848), .C(regd_0_), .Y(_abc_42016_n3436) );
  OAI21X1 OAI21X1_874 ( .A(_abc_42016_n566), .B(_abc_42016_n1848), .C(_abc_42016_n3436), .Y(_abc_42016_n3437) );
  OAI21X1 OAI21X1_875 ( .A(_abc_42016_n3437), .B(_abc_42016_n3430), .C(_abc_42016_n562), .Y(_abc_42016_n3438) );
  OAI21X1 OAI21X1_876 ( .A(regd_1_), .B(_abc_42016_n3432), .C(_abc_42016_n559), .Y(_abc_42016_n3440) );
  OAI21X1 OAI21X1_877 ( .A(regd_1_), .B(_abc_42016_n2357), .C(_abc_42016_n541), .Y(_abc_42016_n3442) );
  OAI21X1 OAI21X1_878 ( .A(_abc_42016_n3443), .B(_abc_42016_n3441), .C(_abc_42016_n3429), .Y(_abc_42016_n3444) );
  OAI21X1 OAI21X1_879 ( .A(_abc_42016_n589), .B(_abc_42016_n3429), .C(_abc_42016_n3444), .Y(regd_1__FF_INPUT) );
  OAI21X1 OAI21X1_88 ( .A(regfil_3__6_), .B(_abc_42016_n600), .C(_abc_42016_n692), .Y(_abc_42016_n936) );
  OAI21X1 OAI21X1_880 ( .A(regd_2_), .B(_abc_42016_n3432), .C(_abc_42016_n559), .Y(_abc_42016_n3446) );
  OAI21X1 OAI21X1_881 ( .A(regd_2_), .B(_abc_42016_n2357), .C(_abc_42016_n541), .Y(_abc_42016_n3448_1) );
  OAI21X1 OAI21X1_882 ( .A(_abc_42016_n3449), .B(_abc_42016_n3447_1), .C(_abc_42016_n557), .Y(_abc_42016_n3450) );
  OAI21X1 OAI21X1_883 ( .A(_abc_42016_n594_1), .B(_abc_42016_n3429), .C(_abc_42016_n3450), .Y(regd_2__FF_INPUT) );
  OAI21X1 OAI21X1_884 ( .A(_abc_42016_n560), .B(_abc_42016_n3453), .C(sp_0_), .Y(_abc_42016_n3454) );
  OAI21X1 OAI21X1_885 ( .A(_abc_42016_n545_1), .B(_abc_42016_n2227), .C(_abc_42016_n1868), .Y(_abc_42016_n3460) );
  OAI21X1 OAI21X1_886 ( .A(_abc_42016_n511), .B(_abc_42016_n546), .C(_abc_42016_n3460), .Y(_abc_42016_n3461) );
  OAI21X1 OAI21X1_887 ( .A(_abc_42016_n3459), .B(_abc_42016_n3461), .C(_abc_42016_n529), .Y(_abc_42016_n3462) );
  OAI21X1 OAI21X1_888 ( .A(_abc_42016_n3466), .B(_abc_42016_n3462), .C(sp_0_), .Y(_abc_42016_n3467) );
  OAI21X1 OAI21X1_889 ( .A(_abc_42016_n709), .B(_abc_42016_n1022), .C(_abc_42016_n673), .Y(_abc_42016_n3471) );
  OAI21X1 OAI21X1_89 ( .A(_abc_42016_n874), .B(_abc_42016_n863), .C(_abc_42016_n939), .Y(_abc_42016_n940) );
  OAI21X1 OAI21X1_890 ( .A(_abc_42016_n2775), .B(_abc_42016_n3470_1), .C(_abc_42016_n3472), .Y(_abc_42016_n3473) );
  OAI21X1 OAI21X1_891 ( .A(_abc_42016_n3476_1), .B(_abc_42016_n2256), .C(_abc_42016_n559), .Y(_abc_42016_n3478) );
  OAI21X1 OAI21X1_892 ( .A(_abc_42016_n3475), .B(_abc_42016_n3477), .C(_abc_42016_n3479_1), .Y(_abc_42016_n3480) );
  OAI21X1 OAI21X1_893 ( .A(_abc_42016_n3097), .B(_abc_42016_n3098), .C(_abc_42016_n1407), .Y(_abc_42016_n3486) );
  OAI21X1 OAI21X1_894 ( .A(_abc_42016_n2376), .B(_abc_42016_n3100), .C(_abc_42016_n3486), .Y(_abc_42016_n3487) );
  OAI21X1 OAI21X1_895 ( .A(_abc_42016_n1159), .B(_abc_42016_n3470_1), .C(_abc_42016_n3488_1), .Y(_abc_42016_n3489) );
  OAI21X1 OAI21X1_896 ( .A(sp_0_), .B(sp_1_), .C(sp_2_), .Y(_abc_42016_n3491_1) );
  OAI21X1 OAI21X1_897 ( .A(sp_0_), .B(_abc_42016_n3119), .C(_abc_42016_n3491_1), .Y(_abc_42016_n3492) );
  OAI21X1 OAI21X1_898 ( .A(_abc_42016_n2758), .B(_abc_42016_n2775), .C(_abc_42016_n1159), .Y(_abc_42016_n3494_1) );
  OAI21X1 OAI21X1_899 ( .A(sp_2_), .B(_abc_42016_n3497_1), .C(_abc_42016_n547), .Y(_abc_42016_n3498) );
  OAI21X1 OAI21X1_9 ( .A(opcode_4_), .B(_abc_42016_n528_1), .C(_abc_42016_n590), .Y(_abc_42016_n591) );
  OAI21X1 OAI21X1_90 ( .A(_abc_42016_n772), .B(_abc_42016_n941_1), .C(_abc_42016_n945), .Y(_abc_42016_n946) );
  OAI21X1 OAI21X1_900 ( .A(_abc_42016_n3487), .B(_abc_42016_n3489), .C(_abc_42016_n3499), .Y(_abc_42016_n3500) );
  OAI21X1 OAI21X1_901 ( .A(_abc_42016_n2775), .B(_abc_42016_n1159), .C(_abc_42016_n2813), .Y(_abc_42016_n3508) );
  OAI21X1 OAI21X1_902 ( .A(_abc_42016_n1139), .B(_abc_42016_n1022), .C(_abc_42016_n3511), .Y(_abc_42016_n3512) );
  OAI21X1 OAI21X1_903 ( .A(_abc_42016_n2813), .B(_abc_42016_n3470_1), .C(_abc_42016_n673), .Y(_abc_42016_n3513) );
  OAI21X1 OAI21X1_904 ( .A(_abc_42016_n3514), .B(_abc_42016_n3515), .C(_abc_42016_n3490), .Y(_abc_42016_n3516) );
  OAI21X1 OAI21X1_905 ( .A(_abc_42016_n2758), .B(_abc_42016_n3517), .C(_abc_42016_n2813), .Y(_abc_42016_n3518_1) );
  OAI21X1 OAI21X1_906 ( .A(sp_3_), .B(_abc_42016_n3497_1), .C(_abc_42016_n547), .Y(_abc_42016_n3524) );
  OAI21X1 OAI21X1_907 ( .A(_abc_42016_n3512), .B(_abc_42016_n3513), .C(_abc_42016_n3525), .Y(_abc_42016_n3526_1) );
  OAI21X1 OAI21X1_908 ( .A(_abc_42016_n1174_1), .B(_abc_42016_n3458), .C(_abc_42016_n3528), .Y(_abc_42016_n3529) );
  OAI21X1 OAI21X1_909 ( .A(_abc_42016_n2813), .B(_abc_42016_n3517), .C(_abc_42016_n1210), .Y(_abc_42016_n3532) );
  OAI21X1 OAI21X1_91 ( .A(_abc_42016_n936), .B(_abc_42016_n935), .C(_abc_42016_n947), .Y(_abc_36783_n3379) );
  OAI21X1 OAI21X1_910 ( .A(_abc_42016_n843), .B(_abc_42016_n1022), .C(_abc_42016_n673), .Y(_abc_42016_n3536) );
  OAI21X1 OAI21X1_911 ( .A(_abc_42016_n1408), .B(_abc_42016_n3134), .C(_abc_42016_n3537), .Y(_abc_42016_n3538) );
  OAI21X1 OAI21X1_912 ( .A(sp_4_), .B(_abc_42016_n3497_1), .C(_abc_42016_n3538), .Y(_abc_42016_n3539) );
  OAI21X1 OAI21X1_913 ( .A(_abc_42016_n1210), .B(_abc_42016_n3470_1), .C(_abc_42016_n3539), .Y(_abc_42016_n3540) );
  OAI21X1 OAI21X1_914 ( .A(_abc_42016_n3541), .B(_abc_42016_n3542), .C(_abc_42016_n3490), .Y(_abc_42016_n3543) );
  OAI21X1 OAI21X1_915 ( .A(_abc_42016_n3520), .B(_abc_42016_n3453), .C(_abc_42016_n1210), .Y(_abc_42016_n3544) );
  OAI21X1 OAI21X1_916 ( .A(_abc_42016_n2306), .B(_abc_42016_n1005), .C(_abc_42016_n673), .Y(_abc_42016_n3554) );
  OAI21X1 OAI21X1_917 ( .A(_abc_42016_n1210), .B(_abc_42016_n3509), .C(_abc_42016_n1279), .Y(_abc_42016_n3557) );
  OAI21X1 OAI21X1_918 ( .A(_abc_42016_n872), .B(_abc_42016_n1022), .C(_abc_42016_n3560), .Y(_abc_42016_n3561) );
  OAI21X1 OAI21X1_919 ( .A(_abc_42016_n1004), .B(_abc_42016_n682), .C(_abc_42016_n3562), .Y(_abc_42016_n3563) );
  OAI21X1 OAI21X1_92 ( .A(regfil_0__6_), .B(_abc_42016_n888), .C(regfil_0__7_), .Y(_abc_42016_n949) );
  OAI21X1 OAI21X1_920 ( .A(_abc_42016_n2758), .B(_abc_42016_n3556), .C(_abc_42016_n3474), .Y(_abc_42016_n3565) );
  OAI21X1 OAI21X1_921 ( .A(_abc_42016_n3564), .B(_abc_42016_n3565), .C(_abc_42016_n3567_1), .Y(_abc_42016_n3568) );
  OAI21X1 OAI21X1_922 ( .A(_abc_42016_n1279), .B(_abc_42016_n3563), .C(_abc_42016_n3569), .Y(_abc_42016_n3570) );
  OAI21X1 OAI21X1_923 ( .A(opcode_7_), .B(opcode_6_), .C(_abc_42016_n3554), .Y(_abc_42016_n3571) );
  OAI21X1 OAI21X1_924 ( .A(_abc_42016_n3577), .B(_abc_42016_n3458), .C(_abc_42016_n3501), .Y(_abc_42016_n3578) );
  OAI21X1 OAI21X1_925 ( .A(_abc_42016_n1279), .B(_abc_42016_n3534), .C(_abc_42016_n1323), .Y(_abc_42016_n3582) );
  OAI21X1 OAI21X1_926 ( .A(_abc_42016_n1408), .B(_abc_42016_n3182), .C(opcode_7_), .Y(_abc_42016_n3586_1) );
  OAI21X1 OAI21X1_927 ( .A(_abc_42016_n3586_1), .B(_abc_42016_n3585), .C(_abc_42016_n3497_1), .Y(_abc_42016_n3587) );
  OAI21X1 OAI21X1_928 ( .A(_abc_42016_n1323), .B(_abc_42016_n3581), .C(_abc_42016_n3587), .Y(_abc_42016_n3588) );
  OAI21X1 OAI21X1_929 ( .A(_abc_42016_n2758), .B(_abc_42016_n1323), .C(_abc_42016_n3181), .Y(_abc_42016_n3591) );
  OAI21X1 OAI21X1_93 ( .A(_abc_42016_n913), .B(_abc_42016_n885), .C(_abc_42016_n954), .Y(_abc_42016_n955) );
  OAI21X1 OAI21X1_930 ( .A(_abc_42016_n3590), .B(_abc_42016_n3591), .C(_abc_42016_n3490), .Y(_abc_42016_n3592) );
  OAI21X1 OAI21X1_931 ( .A(_abc_42016_n2758), .B(_abc_42016_n3556), .C(_abc_42016_n1323), .Y(_abc_42016_n3593) );
  OAI21X1 OAI21X1_932 ( .A(_abc_42016_n1323), .B(_abc_42016_n2255), .C(_abc_42016_n559), .Y(_abc_42016_n3596) );
  OAI21X1 OAI21X1_933 ( .A(_abc_42016_n3182), .B(_abc_42016_n3503), .C(_abc_42016_n3601), .Y(_abc_42016_n3602) );
  OAI21X1 OAI21X1_934 ( .A(_abc_42016_n1323), .B(_abc_42016_n3556), .C(_abc_42016_n1327_1), .Y(_abc_42016_n3608) );
  OAI21X1 OAI21X1_935 ( .A(_abc_42016_n3605), .B(_abc_42016_n3503), .C(_abc_42016_n3610), .Y(_abc_42016_n3611) );
  OAI21X1 OAI21X1_936 ( .A(_abc_42016_n3614), .B(_abc_42016_n3613), .C(_abc_42016_n3490), .Y(_abc_42016_n3615) );
  OAI21X1 OAI21X1_937 ( .A(sp_7_), .B(_abc_42016_n3594), .C(_abc_42016_n3616), .Y(_abc_42016_n3617) );
  OAI21X1 OAI21X1_938 ( .A(_abc_42016_n560), .B(_abc_42016_n3453), .C(_abc_42016_n3554), .Y(_abc_42016_n3619) );
  OAI21X1 OAI21X1_939 ( .A(_abc_42016_n1408), .B(_abc_42016_n3605), .C(_abc_42016_n3620), .Y(_abc_42016_n3621) );
  OAI21X1 OAI21X1_94 ( .A(_abc_42016_n526_1), .B(_abc_42016_n751), .C(rdatahold_7_), .Y(_abc_42016_n957_1) );
  OAI21X1 OAI21X1_940 ( .A(_abc_42016_n1327_1), .B(_abc_42016_n3619), .C(_abc_42016_n3622), .Y(_abc_42016_n3623) );
  OAI21X1 OAI21X1_941 ( .A(_abc_42016_n3618), .B(_abc_42016_n3623), .C(_abc_42016_n547), .Y(_abc_42016_n3624) );
  OAI21X1 OAI21X1_942 ( .A(_abc_42016_n3226), .B(_abc_42016_n3225), .C(_abc_42016_n3527), .Y(_abc_42016_n3626) );
  OAI21X1 OAI21X1_943 ( .A(_abc_42016_n3475), .B(_abc_42016_n3633), .C(_abc_42016_n2131_1), .Y(_abc_42016_n3634) );
  OAI21X1 OAI21X1_944 ( .A(_abc_42016_n2256), .B(_abc_42016_n3632), .C(_abc_42016_n3634), .Y(_abc_42016_n3635) );
  OAI21X1 OAI21X1_945 ( .A(_abc_42016_n3635), .B(_abc_42016_n3631), .C(_abc_42016_n3628_1), .Y(_abc_42016_n3636) );
  OAI21X1 OAI21X1_946 ( .A(_abc_42016_n3226), .B(_abc_42016_n3225), .C(_abc_42016_n1407), .Y(_abc_42016_n3637) );
  OAI21X1 OAI21X1_947 ( .A(_abc_42016_n629), .B(_abc_42016_n1022), .C(_abc_42016_n3637), .Y(_abc_42016_n3638) );
  OAI21X1 OAI21X1_948 ( .A(_abc_42016_n1327_1), .B(_abc_42016_n3583), .C(_abc_42016_n2131_1), .Y(_abc_42016_n3639) );
  OAI21X1 OAI21X1_949 ( .A(_abc_42016_n2376), .B(_abc_42016_n3640), .C(_abc_42016_n3581), .Y(_abc_42016_n3641) );
  OAI21X1 OAI21X1_95 ( .A(regfil_4__7_), .B(_abc_42016_n727), .C(opcode_2_), .Y(_abc_42016_n958) );
  OAI21X1 OAI21X1_950 ( .A(_abc_42016_n3575), .B(_abc_42016_n3640), .C(_abc_42016_n3645), .Y(_abc_42016_n3646) );
  OAI21X1 OAI21X1_951 ( .A(_abc_42016_n3650), .B(_abc_42016_n3649), .C(_abc_42016_n3490), .Y(_abc_42016_n3651) );
  OAI21X1 OAI21X1_952 ( .A(_abc_42016_n2758), .B(_abc_42016_n3653), .C(_abc_42016_n3654), .Y(_abc_42016_n3655) );
  OAI21X1 OAI21X1_953 ( .A(_abc_42016_n2131_1), .B(_abc_42016_n3607), .C(_abc_42016_n2127_1), .Y(_abc_42016_n3657) );
  OAI21X1 OAI21X1_954 ( .A(_abc_42016_n3661), .B(_abc_42016_n3660), .C(_abc_42016_n673), .Y(_abc_42016_n3662) );
  OAI21X1 OAI21X1_955 ( .A(_abc_42016_n2127_1), .B(_abc_42016_n3619), .C(_abc_42016_n3662), .Y(_abc_42016_n3663) );
  OAI21X1 OAI21X1_956 ( .A(_abc_42016_n3656), .B(_abc_42016_n3663), .C(_abc_42016_n547), .Y(_abc_42016_n3664) );
  OAI21X1 OAI21X1_957 ( .A(_abc_42016_n3503), .B(_abc_42016_n3249), .C(_abc_42016_n3665), .Y(_abc_42016_n3666) );
  OAI21X1 OAI21X1_958 ( .A(_abc_42016_n566), .B(_abc_42016_n3649), .C(_abc_42016_n3501), .Y(_abc_42016_n3669) );
  OAI21X1 OAI21X1_959 ( .A(_abc_42016_n3453), .B(_abc_42016_n3669), .C(sp_10_), .Y(_abc_42016_n3670_1) );
  OAI21X1 OAI21X1_96 ( .A(regfil_6__7_), .B(_abc_42016_n539), .C(_abc_42016_n961), .Y(_abc_42016_n962) );
  OAI21X1 OAI21X1_960 ( .A(_abc_42016_n2758), .B(_abc_42016_n3672), .C(_abc_42016_n3474), .Y(_abc_42016_n3673) );
  OAI21X1 OAI21X1_961 ( .A(_abc_42016_n3674), .B(_abc_42016_n3673), .C(_abc_42016_n559), .Y(_abc_42016_n3675) );
  OAI21X1 OAI21X1_962 ( .A(_abc_42016_n2127_1), .B(_abc_42016_n3629), .C(_abc_42016_n2122), .Y(_abc_42016_n3678) );
  OAI21X1 OAI21X1_963 ( .A(_abc_42016_n1408), .B(_abc_42016_n3271), .C(_abc_42016_n3681), .Y(_abc_42016_n3682) );
  OAI21X1 OAI21X1_964 ( .A(_abc_42016_n3682), .B(_abc_42016_n3680), .C(_abc_42016_n547), .Y(_abc_42016_n3683) );
  OAI21X1 OAI21X1_965 ( .A(_abc_42016_n2118), .B(_abc_42016_n3470_1), .C(_abc_42016_n3690_1), .Y(_abc_42016_n3691) );
  OAI21X1 OAI21X1_966 ( .A(_abc_42016_n2122), .B(_abc_42016_n3653), .C(_abc_42016_n2118), .Y(_abc_42016_n3695) );
  OAI21X1 OAI21X1_967 ( .A(_abc_42016_n1408), .B(_abc_42016_n3298), .C(_abc_42016_n3696), .Y(_abc_42016_n3697) );
  OAI21X1 OAI21X1_968 ( .A(_abc_42016_n3698), .B(_abc_42016_n3699), .C(_abc_42016_n3490), .Y(_abc_42016_n3700) );
  OAI21X1 OAI21X1_969 ( .A(_abc_42016_n2758), .B(_abc_42016_n3672), .C(_abc_42016_n2118), .Y(_abc_42016_n3701) );
  OAI21X1 OAI21X1_97 ( .A(regfil_3__7_), .B(_abc_42016_n600), .C(_abc_42016_n692), .Y(_abc_42016_n973) );
  OAI21X1 OAI21X1_970 ( .A(sp_11_), .B(_abc_42016_n3497_1), .C(_abc_42016_n547), .Y(_abc_42016_n3705) );
  OAI21X1 OAI21X1_971 ( .A(_abc_42016_n3691), .B(_abc_42016_n3697), .C(_abc_42016_n3706), .Y(_abc_42016_n3707) );
  OAI21X1 OAI21X1_972 ( .A(_abc_42016_n811), .B(_abc_42016_n3458), .C(_abc_42016_n3501), .Y(_abc_42016_n3709) );
  OAI21X1 OAI21X1_973 ( .A(sp_0_), .B(_abc_42016_n3296_1), .C(sp_12_), .Y(_abc_42016_n3715) );
  OAI21X1 OAI21X1_974 ( .A(_abc_42016_n3720), .B(_abc_42016_n3716), .C(_abc_42016_n559), .Y(_abc_42016_n3721) );
  OAI21X1 OAI21X1_975 ( .A(_abc_42016_n3692), .B(_abc_42016_n3629), .C(_abc_42016_n2113), .Y(_abc_42016_n3724) );
  OAI21X1 OAI21X1_976 ( .A(_abc_42016_n3723), .B(_abc_42016_n3728), .C(_abc_42016_n673), .Y(_abc_42016_n3729) );
  OAI21X1 OAI21X1_977 ( .A(_abc_42016_n3575), .B(_abc_42016_n3727), .C(_abc_42016_n3733_1), .Y(_abc_42016_n3734) );
  OAI21X1 OAI21X1_978 ( .A(_abc_42016_n3734), .B(_abc_42016_n3731), .C(_abc_42016_n3501), .Y(_abc_42016_n3735) );
  OAI21X1 OAI21X1_979 ( .A(_abc_42016_n2113), .B(_abc_42016_n3501), .C(_abc_42016_n3735), .Y(sp_12__FF_INPUT) );
  OAI21X1 OAI21X1_98 ( .A(_abc_42016_n977), .B(_abc_42016_n975), .C(_abc_42016_n779), .Y(_abc_42016_n978) );
  OAI21X1 OAI21X1_980 ( .A(_abc_42016_n3453), .B(_abc_42016_n3718), .C(_abc_42016_n2109_1), .Y(_abc_42016_n3737) );
  OAI21X1 OAI21X1_981 ( .A(_abc_42016_n3742), .B(_abc_42016_n3741), .C(_abc_42016_n3490), .Y(_abc_42016_n3743) );
  OAI21X1 OAI21X1_982 ( .A(_abc_42016_n2109_1), .B(_abc_42016_n3501), .C(_abc_42016_n3756), .Y(sp_13__FF_INPUT) );
  OAI21X1 OAI21X1_983 ( .A(_abc_42016_n3759), .B(_abc_42016_n3758), .C(_abc_42016_n3490), .Y(_abc_42016_n3760) );
  OAI21X1 OAI21X1_984 ( .A(_abc_42016_n2109_1), .B(_abc_42016_n3718), .C(_abc_42016_n2103), .Y(_abc_42016_n3761) );
  OAI21X1 OAI21X1_985 ( .A(_abc_42016_n3765), .B(_abc_42016_n3764), .C(_abc_42016_n3761), .Y(_abc_42016_n3766) );
  OAI21X1 OAI21X1_986 ( .A(_abc_42016_n2109_1), .B(_abc_42016_n3726), .C(_abc_42016_n2103), .Y(_abc_42016_n3768) );
  OAI21X1 OAI21X1_987 ( .A(_abc_42016_n1554), .B(_abc_42016_n1022), .C(_abc_42016_n3581), .Y(_abc_42016_n3770) );
  OAI21X1 OAI21X1_988 ( .A(_abc_42016_n2376), .B(_abc_42016_n3769), .C(_abc_42016_n3771), .Y(_abc_42016_n3772) );
  OAI21X1 OAI21X1_989 ( .A(_abc_42016_n1793), .B(_abc_42016_n3458), .C(_abc_42016_n3501), .Y(_abc_42016_n3775_1) );
  OAI21X1 OAI21X1_99 ( .A(regfil_3__7_), .B(_abc_42016_n979_1), .C(_abc_42016_n981), .Y(_abc_42016_n982) );
  OAI21X1 OAI21X1_990 ( .A(_abc_42016_n2101), .B(_abc_42016_n2255), .C(_abc_42016_n559), .Y(_abc_42016_n3779) );
  OAI21X1 OAI21X1_991 ( .A(_abc_42016_n3781), .B(_abc_42016_n3780), .C(_abc_42016_n3490), .Y(_abc_42016_n3782) );
  OAI21X1 OAI21X1_992 ( .A(_abc_42016_n3784), .B(_abc_42016_n3783), .C(_abc_42016_n3474), .Y(_abc_42016_n3785) );
  OAI21X1 OAI21X1_993 ( .A(_abc_42016_n1801_1), .B(_abc_42016_n1022), .C(_abc_42016_n673), .Y(_abc_42016_n3787) );
  OAI21X1 OAI21X1_994 ( .A(sp_15_), .B(_abc_42016_n3497_1), .C(_abc_42016_n547), .Y(_abc_42016_n3791) );
  OAI21X1 OAI21X1_995 ( .A(_abc_42016_n3779), .B(_abc_42016_n3786), .C(_abc_42016_n3792), .Y(_abc_42016_n3793) );
  OAI21X1 OAI21X1_996 ( .A(_abc_42016_n1604_1), .B(_abc_42016_n988), .C(regfil_4__0_), .Y(_abc_42016_n3799) );
  OAI21X1 OAI21X1_997 ( .A(_abc_42016_n1631), .B(_abc_42016_n697), .C(_abc_42016_n994), .Y(_abc_42016_n3802) );
  OAI21X1 OAI21X1_998 ( .A(_abc_42016_n1022), .B(_abc_42016_n562), .C(_abc_42016_n1002), .Y(_abc_42016_n3803) );
  OAI21X1 OAI21X1_999 ( .A(_abc_42016_n629), .B(_abc_42016_n1335_1), .C(_abc_42016_n1125), .Y(_abc_42016_n3808) );
  OAI22X1 OAI22X1_1 ( .A(_abc_42016_n627), .B(_abc_42016_n632), .C(_abc_42016_n633), .D(_abc_42016_n636), .Y(_abc_42016_n637) );
  OAI22X1 OAI22X1_10 ( .A(rdatahold2_5_), .B(_abc_42016_n701), .C(_abc_42016_n881), .D(_abc_42016_n873), .Y(_abc_42016_n882) );
  OAI22X1 OAI22X1_100 ( .A(\data[0] ), .B(_abc_42016_n4048), .C(_abc_42016_n4344), .D(_abc_42016_n4355), .Y(_abc_42016_n4356) );
  OAI22X1 OAI22X1_101 ( .A(_abc_42016_n1454), .B(_abc_42016_n4051), .C(_abc_42016_n1974), .D(_abc_42016_n4060), .Y(_abc_42016_n4397) );
  OAI22X1 OAI22X1_102 ( .A(_abc_42016_n3050), .B(_abc_42016_n2497), .C(_abc_42016_n719), .D(_abc_42016_n4472), .Y(_abc_42016_n4481) );
  OAI22X1 OAI22X1_103 ( .A(_abc_42016_n1382), .B(_abc_42016_n2024), .C(_abc_42016_n2786), .D(_abc_42016_n2733), .Y(_abc_42016_n4485) );
  OAI22X1 OAI22X1_104 ( .A(_abc_42016_n3078_1), .B(_abc_42016_n2497), .C(_abc_42016_n1675), .D(_abc_42016_n4472), .Y(_abc_42016_n4486) );
  OAI22X1 OAI22X1_105 ( .A(_abc_42016_n1357), .B(_abc_42016_n2024), .C(_abc_42016_n2803), .D(_abc_42016_n2733), .Y(_abc_42016_n4490) );
  OAI22X1 OAI22X1_106 ( .A(_abc_42016_n3105_1), .B(_abc_42016_n2497), .C(_abc_42016_n811), .D(_abc_42016_n4472), .Y(_abc_42016_n4491) );
  OAI22X1 OAI22X1_107 ( .A(_abc_42016_n3128), .B(_abc_42016_n2497), .C(_abc_42016_n2820), .D(_abc_42016_n2733), .Y(_abc_42016_n4495) );
  OAI22X1 OAI22X1_108 ( .A(_abc_42016_n1356), .B(_abc_42016_n2024), .C(_abc_42016_n2471), .D(_abc_42016_n4472), .Y(_abc_42016_n4496) );
  OAI22X1 OAI22X1_109 ( .A(_abc_42016_n3153), .B(_abc_42016_n2497), .C(_abc_42016_n2836), .D(_abc_42016_n2733), .Y(_abc_42016_n4500) );
  OAI22X1 OAI22X1_11 ( .A(_abc_42016_n893), .B(_abc_42016_n727), .C(_abc_42016_n642), .D(_abc_42016_n626), .Y(_abc_42016_n894) );
  OAI22X1 OAI22X1_110 ( .A(_abc_42016_n2649), .B(_abc_42016_n2024), .C(_abc_42016_n891), .D(_abc_42016_n4472), .Y(_abc_42016_n4501) );
  OAI22X1 OAI22X1_111 ( .A(_abc_42016_n3175), .B(_abc_42016_n2497), .C(_abc_42016_n2852), .D(_abc_42016_n2733), .Y(_abc_42016_n4505) );
  OAI22X1 OAI22X1_112 ( .A(_abc_42016_n1355), .B(_abc_42016_n2024), .C(_abc_42016_n1793), .D(_abc_42016_n4472), .Y(_abc_42016_n4506) );
  OAI22X1 OAI22X1_113 ( .A(_abc_42016_n3201), .B(_abc_42016_n2497), .C(_abc_42016_n2869), .D(_abc_42016_n2733), .Y(_abc_42016_n4510) );
  OAI22X1 OAI22X1_114 ( .A(_abc_42016_n1354), .B(_abc_42016_n2024), .C(_abc_42016_n2478), .D(_abc_42016_n4472), .Y(_abc_42016_n4511) );
  OAI22X1 OAI22X1_115 ( .A(_abc_42016_n1353), .B(_abc_42016_n2024), .C(_abc_42016_n2887), .D(_abc_42016_n2733), .Y(_abc_42016_n4516) );
  OAI22X1 OAI22X1_116 ( .A(_abc_42016_n1422), .B(_abc_42016_n2024), .C(_abc_42016_n3245_1), .D(_abc_42016_n2497), .Y(_abc_42016_n4519) );
  OAI22X1 OAI22X1_117 ( .A(_abc_42016_n1449), .B(_abc_42016_n2024), .C(_abc_42016_n3268), .D(_abc_42016_n2497), .Y(_abc_42016_n4523) );
  OAI22X1 OAI22X1_118 ( .A(_abc_42016_n1477), .B(_abc_42016_n2024), .C(_abc_42016_n3291), .D(_abc_42016_n2497), .Y(_abc_42016_n4527) );
  OAI22X1 OAI22X1_119 ( .A(_abc_42016_n1503), .B(_abc_42016_n2024), .C(_abc_42016_n3316), .D(_abc_42016_n2497), .Y(_abc_42016_n4531) );
  OAI22X1 OAI22X1_12 ( .A(_abc_42016_n895), .B(_abc_42016_n539), .C(_abc_42016_n874), .D(_abc_42016_n565), .Y(_abc_42016_n896) );
  OAI22X1 OAI22X1_120 ( .A(_abc_42016_n3337), .B(_abc_42016_n2497), .C(_abc_42016_n2972), .D(_abc_42016_n2733), .Y(_abc_42016_n4537) );
  OAI22X1 OAI22X1_121 ( .A(_abc_42016_n1557), .B(_abc_42016_n2024), .C(_abc_42016_n3361), .D(_abc_42016_n2497), .Y(_abc_42016_n4540) );
  OAI22X1 OAI22X1_122 ( .A(_abc_42016_n581_1), .B(_abc_42016_n4604), .C(_abc_42016_n2371), .D(_abc_42016_n558), .Y(_abc_42016_n4605) );
  OAI22X1 OAI22X1_123 ( .A(_abc_42016_n2050), .B(_abc_42016_n604_1), .C(_abc_42016_n2056), .D(_abc_42016_n1004), .Y(_abc_42016_n4640) );
  OAI22X1 OAI22X1_124 ( .A(alu__abc_41682_n81), .B(alu__abc_41682_n92), .C(alu__abc_41682_n111), .D(alu__abc_41682_n110), .Y(alu__abc_41682_n112) );
  OAI22X1 OAI22X1_125 ( .A(alu__abc_41682_n125), .B(alu_opra_0_), .C(alu__abc_41682_n34), .D(alu__abc_41682_n35), .Y(alu__abc_41682_n126) );
  OAI22X1 OAI22X1_126 ( .A(alu__abc_41682_n94), .B(alu__abc_41682_n218), .C(alu__abc_41682_n179), .D(alu__abc_41682_n90), .Y(alu__abc_41682_n219) );
  OAI22X1 OAI22X1_127 ( .A(alu__abc_41682_n107), .B(alu__abc_41682_n194), .C(alu__abc_41682_n98), .D(alu__abc_41682_n359), .Y(alu__abc_41682_n360) );
  OAI22X1 OAI22X1_13 ( .A(regfil_0__6_), .B(_abc_42016_n727), .C(regfil_3__6_), .D(_abc_42016_n565), .Y(_abc_42016_n918) );
  OAI22X1 OAI22X1_14 ( .A(_abc_42016_n918), .B(_abc_42016_n921), .C(_abc_42016_n922), .D(_abc_42016_n926), .Y(_abc_42016_n927) );
  OAI22X1 OAI22X1_15 ( .A(regfil_1__7_), .B(_abc_42016_n626), .C(regfil_3__7_), .D(_abc_42016_n565), .Y(_abc_42016_n963) );
  OAI22X1 OAI22X1_16 ( .A(_abc_42016_n963), .B(_abc_42016_n966), .C(_abc_42016_n958), .D(_abc_42016_n962), .Y(_abc_42016_n967) );
  OAI22X1 OAI22X1_17 ( .A(_abc_42016_n757), .B(_abc_42016_n1048), .C(_abc_42016_n1151), .D(_abc_42016_n1156), .Y(_abc_42016_n1157) );
  OAI22X1 OAI22X1_18 ( .A(rdatahold2_5_), .B(_abc_42016_n1097), .C(_abc_42016_n1223), .D(_abc_42016_n1255), .Y(_abc_42016_n1256) );
  OAI22X1 OAI22X1_19 ( .A(_abc_42016_n1333_1), .B(_abc_42016_n1341_1), .C(_abc_42016_n1304), .D(_abc_42016_n1303), .Y(_abc_42016_n1342) );
  OAI22X1 OAI22X1_2 ( .A(regfil_3__0_), .B(_abc_42016_n684), .C(_abc_42016_n695), .D(_abc_42016_n697), .Y(_abc_42016_n698) );
  OAI22X1 OAI22X1_20 ( .A(_abc_42016_n1419), .B(_abc_42016_n1345), .C(_abc_42016_n558), .D(_abc_42016_n1443), .Y(wdatahold2_1__FF_INPUT) );
  OAI22X1 OAI22X1_21 ( .A(opcode_5_), .B(_abc_42016_n1456), .C(_abc_42016_n1454), .D(_abc_42016_n1004), .Y(_abc_42016_n1457) );
  OAI22X1 OAI22X1_22 ( .A(_abc_42016_n1445), .B(_abc_42016_n1345), .C(_abc_42016_n558), .D(_abc_42016_n1472), .Y(wdatahold2_2__FF_INPUT) );
  OAI22X1 OAI22X1_23 ( .A(_abc_42016_n1474), .B(_abc_42016_n1345), .C(_abc_42016_n558), .D(_abc_42016_n1498), .Y(wdatahold2_3__FF_INPUT) );
  OAI22X1 OAI22X1_24 ( .A(_abc_42016_n1500), .B(_abc_42016_n1345), .C(_abc_42016_n558), .D(_abc_42016_n1524), .Y(wdatahold2_4__FF_INPUT) );
  OAI22X1 OAI22X1_25 ( .A(_abc_42016_n1526), .B(_abc_42016_n1345), .C(_abc_42016_n558), .D(_abc_42016_n1551), .Y(wdatahold2_5__FF_INPUT) );
  OAI22X1 OAI22X1_26 ( .A(_abc_42016_n1553), .B(_abc_42016_n1345), .C(_abc_42016_n558), .D(_abc_42016_n1581), .Y(wdatahold2_6__FF_INPUT) );
  OAI22X1 OAI22X1_27 ( .A(_abc_42016_n719), .B(_abc_42016_n701), .C(_abc_42016_n1656), .D(_abc_42016_n606), .Y(_abc_42016_n1658_1) );
  OAI22X1 OAI22X1_28 ( .A(rdatahold_7_), .B(_abc_42016_n688), .C(_abc_42016_n1802_1), .D(_abc_42016_n1808), .Y(_abc_42016_n1809) );
  OAI22X1 OAI22X1_29 ( .A(_abc_42016_n628), .B(_abc_42016_n1842), .C(_abc_42016_n1908), .D(_abc_42016_n1920), .Y(_abc_42016_n1921) );
  OAI22X1 OAI22X1_3 ( .A(rdatahold2_1_), .B(_abc_42016_n701), .C(_abc_42016_n708), .D(_abc_42016_n710), .Y(_abc_42016_n711) );
  OAI22X1 OAI22X1_30 ( .A(_abc_42016_n1454), .B(_abc_42016_n1842), .C(_abc_42016_n1951), .D(_abc_42016_n1955_1), .Y(_abc_42016_n1956) );
  OAI22X1 OAI22X1_31 ( .A(_abc_42016_n924), .B(_abc_42016_n1842), .C(_abc_42016_n2002), .D(_abc_42016_n2006), .Y(_abc_42016_n2007) );
  OAI22X1 OAI22X1_32 ( .A(_abc_42016_n1801_1), .B(_abc_42016_n1912), .C(_abc_42016_n1832), .D(_abc_42016_n533), .Y(_abc_42016_n2012) );
  OAI22X1 OAI22X1_33 ( .A(_abc_42016_n1380), .B(_abc_42016_n2096), .C(_abc_42016_n1801_1), .D(_abc_42016_n1046), .Y(_abc_42016_n2097) );
  OAI22X1 OAI22X1_34 ( .A(_abc_42016_n539), .B(_abc_42016_n2254), .C(_abc_42016_n669), .D(_abc_42016_n2291), .Y(_abc_42016_n2292) );
  OAI22X1 OAI22X1_35 ( .A(_abc_42016_n1400), .B(_abc_42016_n2503), .C(_abc_42016_n1381), .D(_abc_42016_n1405), .Y(_abc_42016_n2504) );
  OAI22X1 OAI22X1_36 ( .A(_abc_42016_n1380), .B(_abc_42016_n2562), .C(_abc_42016_n757), .D(_abc_42016_n1061), .Y(_abc_42016_n2563) );
  OAI22X1 OAI22X1_37 ( .A(_abc_42016_n1380), .B(_abc_42016_n2632), .C(_abc_42016_n2635), .D(_abc_42016_n1378), .Y(_abc_42016_n2636) );
  OAI22X1 OAI22X1_38 ( .A(_abc_42016_n2583), .B(_abc_42016_n2585), .C(_abc_42016_n2499), .D(_abc_42016_n2698), .Y(wdatahold_6__FF_INPUT) );
  OAI22X1 OAI22X1_39 ( .A(_abc_42016_n1044), .B(_abc_42016_n2272), .C(raddrhold_0_), .D(_abc_42016_n2733), .Y(_abc_42016_n2757) );
  OAI22X1 OAI22X1_4 ( .A(_abc_42016_n721), .B(_abc_42016_n725), .C(_abc_42016_n726), .D(_abc_42016_n730), .Y(_abc_42016_n731) );
  OAI22X1 OAI22X1_40 ( .A(_abc_42016_n2758), .B(_abc_42016_n2739), .C(pc_0_), .D(_abc_42016_n2759), .Y(_abc_42016_n2760) );
  OAI22X1 OAI22X1_41 ( .A(_abc_42016_n2775), .B(_abc_42016_n2739), .C(_abc_42016_n2769), .D(_abc_42016_n2759), .Y(_abc_42016_n2776) );
  OAI22X1 OAI22X1_42 ( .A(_abc_42016_n1159), .B(_abc_42016_n2739), .C(_abc_42016_n2562), .D(_abc_42016_n2759), .Y(_abc_42016_n2798) );
  OAI22X1 OAI22X1_43 ( .A(_abc_42016_n2813), .B(_abc_42016_n2739), .C(_abc_42016_n2592), .D(_abc_42016_n2759), .Y(_abc_42016_n2814) );
  OAI22X1 OAI22X1_44 ( .A(_abc_42016_n2310), .B(_abc_42016_n2597), .C(_abc_42016_n2592), .D(_abc_42016_n2425), .Y(_abc_42016_n2815) );
  OAI22X1 OAI22X1_45 ( .A(_abc_42016_n843), .B(_abc_42016_n2429_1), .C(_abc_42016_n2632), .D(_abc_42016_n2425), .Y(_abc_42016_n2824) );
  OAI22X1 OAI22X1_46 ( .A(_abc_42016_n1179), .B(_abc_42016_n2272), .C(_abc_42016_n2829), .D(_abc_42016_n2830), .Y(_abc_42016_n2831) );
  OAI22X1 OAI22X1_47 ( .A(_abc_42016_n1210), .B(_abc_42016_n2739), .C(_abc_42016_n2632), .D(_abc_42016_n2759), .Y(_abc_42016_n2833_1) );
  OAI22X1 OAI22X1_48 ( .A(_abc_42016_n1279), .B(_abc_42016_n2739), .C(_abc_42016_n2653), .D(_abc_42016_n2759), .Y(_abc_42016_n2841) );
  OAI22X1 OAI22X1_49 ( .A(_abc_42016_n1323), .B(_abc_42016_n2739), .C(_abc_42016_n2676), .D(_abc_42016_n2759), .Y(_abc_42016_n2866) );
  OAI22X1 OAI22X1_5 ( .A(regfil_1__2_), .B(_abc_42016_n626), .C(regfil_3__2_), .D(_abc_42016_n565), .Y(_abc_42016_n752) );
  OAI22X1 OAI22X1_50 ( .A(_abc_42016_n959), .B(_abc_42016_n2429_1), .C(_abc_42016_n2718), .D(_abc_42016_n2310), .Y(_abc_42016_n2873) );
  OAI22X1 OAI22X1_51 ( .A(_abc_42016_n1327_1), .B(_abc_42016_n2739), .C(_abc_42016_n2716), .D(_abc_42016_n2759), .Y(_abc_42016_n2876) );
  OAI22X1 OAI22X1_52 ( .A(_abc_42016_n2131_1), .B(_abc_42016_n2739), .C(_abc_42016_n1393), .D(_abc_42016_n2759), .Y(_abc_42016_n2897) );
  OAI22X1 OAI22X1_53 ( .A(_abc_42016_n2903), .B(_abc_42016_n2904), .C(_abc_42016_n1425), .D(_abc_42016_n2425), .Y(_abc_42016_n2905) );
  OAI22X1 OAI22X1_54 ( .A(_abc_42016_n2127_1), .B(_abc_42016_n2739), .C(_abc_42016_n1425), .D(_abc_42016_n2759), .Y(_abc_42016_n2907) );
  OAI22X1 OAI22X1_55 ( .A(_abc_42016_n719), .B(_abc_42016_n2272), .C(_abc_42016_n2914), .D(_abc_42016_n2913), .Y(_abc_42016_n2915) );
  OAI22X1 OAI22X1_56 ( .A(_abc_42016_n2922), .B(_abc_42016_n2923), .C(_abc_42016_n1456), .D(_abc_42016_n2310), .Y(_abc_42016_n2924_1) );
  OAI22X1 OAI22X1_57 ( .A(_abc_42016_n2118), .B(_abc_42016_n2739), .C(_abc_42016_n2759), .D(_abc_42016_n1481), .Y(_abc_42016_n2948) );
  OAI22X1 OAI22X1_58 ( .A(_abc_42016_n811), .B(_abc_42016_n2272), .C(_abc_42016_n2952), .D(_abc_42016_n2951), .Y(_abc_42016_n2953) );
  OAI22X1 OAI22X1_59 ( .A(_abc_42016_n3070), .B(_abc_42016_n2261), .C(_abc_42016_n709), .D(_abc_42016_n2613), .Y(_abc_42016_n3071) );
  OAI22X1 OAI22X1_6 ( .A(_abc_42016_n752), .B(_abc_42016_n755), .C(_abc_42016_n756), .D(_abc_42016_n760), .Y(_abc_42016_n761) );
  OAI22X1 OAI22X1_60 ( .A(_abc_42016_n3031), .B(_abc_42016_n3103), .C(_abc_42016_n3078_1), .D(_abc_42016_n3080_1), .Y(waddrhold_2__FF_INPUT) );
  OAI22X1 OAI22X1_61 ( .A(_abc_42016_n3034), .B(_abc_42016_n2597), .C(_abc_42016_n1848), .D(_abc_42016_n3112), .Y(_abc_42016_n3113) );
  OAI22X1 OAI22X1_62 ( .A(_abc_42016_n3105_1), .B(_abc_42016_n3080_1), .C(_abc_42016_n3031), .D(_abc_42016_n3126_1), .Y(waddrhold_3__FF_INPUT) );
  OAI22X1 OAI22X1_63 ( .A(_abc_42016_n1210), .B(_abc_42016_n1061), .C(_abc_42016_n3134), .D(_abc_42016_n3130), .Y(_abc_42016_n3135) );
  OAI22X1 OAI22X1_64 ( .A(_abc_42016_n3034), .B(_abc_42016_n2622), .C(_abc_42016_n3137), .D(_abc_42016_n3139), .Y(_abc_42016_n3140) );
  OAI22X1 OAI22X1_65 ( .A(_abc_42016_n1323), .B(_abc_42016_n1061), .C(_abc_42016_n3182), .D(_abc_42016_n3130), .Y(_abc_42016_n3183) );
  OAI22X1 OAI22X1_66 ( .A(_abc_42016_n1347), .B(_abc_42016_n2678), .C(_abc_42016_n3185), .D(_abc_42016_n3187), .Y(_abc_42016_n3188) );
  OAI22X1 OAI22X1_67 ( .A(_abc_42016_n1848), .B(_abc_42016_n3231), .C(_abc_42016_n3223), .D(_abc_42016_n2293), .Y(_abc_42016_n3232) );
  OAI22X1 OAI22X1_68 ( .A(_abc_42016_n2127_1), .B(_abc_42016_n1061), .C(_abc_42016_n3130), .D(_abc_42016_n3249), .Y(_abc_42016_n3250) );
  OAI22X1 OAI22X1_69 ( .A(_abc_42016_n1848), .B(_abc_42016_n2943), .C(_abc_42016_n3291), .D(_abc_42016_n2293), .Y(_abc_42016_n3301) );
  OAI22X1 OAI22X1_7 ( .A(rdatahold2_2_), .B(_abc_42016_n701), .C(_abc_42016_n777), .D(_abc_42016_n786), .Y(_abc_42016_n787) );
  OAI22X1 OAI22X1_70 ( .A(_abc_42016_n842), .B(_abc_42016_n2298), .C(_abc_42016_n3316), .D(_abc_42016_n2358), .Y(_abc_42016_n3329) );
  OAI22X1 OAI22X1_71 ( .A(_abc_42016_n1347), .B(_abc_42016_n1594_1), .C(_abc_42016_n3394), .D(_abc_42016_n3396), .Y(_abc_42016_n3397_1) );
  OAI22X1 OAI22X1_72 ( .A(_abc_42016_n3452), .B(_abc_42016_n3454), .C(_abc_42016_n3462), .D(_abc_42016_n3456), .Y(_abc_42016_n3463) );
  OAI22X1 OAI22X1_73 ( .A(_abc_42016_n3070), .B(_abc_42016_n3458), .C(sp_1_), .D(_abc_42016_n3460), .Y(_abc_42016_n3483) );
  OAI22X1 OAI22X1_74 ( .A(_abc_42016_n1130), .B(_abc_42016_n3458), .C(_abc_42016_n3099), .D(_abc_42016_n3503), .Y(_abc_42016_n3504) );
  OAI22X1 OAI22X1_75 ( .A(_abc_42016_n1408), .B(_abc_42016_n3164), .C(_abc_42016_n2376), .D(_abc_42016_n3558), .Y(_abc_42016_n3559) );
  OAI22X1 OAI22X1_76 ( .A(_abc_42016_n3164), .B(_abc_42016_n3503), .C(_abc_42016_n3575), .D(_abc_42016_n3558), .Y(_abc_42016_n3576) );
  OAI22X1 OAI22X1_77 ( .A(_abc_42016_n923), .B(_abc_42016_n1022), .C(_abc_42016_n2376), .D(_abc_42016_n3584), .Y(_abc_42016_n3585) );
  OAI22X1 OAI22X1_78 ( .A(_abc_42016_n722), .B(_abc_42016_n1022), .C(_abc_42016_n1408), .D(_abc_42016_n3249), .Y(_abc_42016_n3661) );
  OAI22X1 OAI22X1_79 ( .A(_abc_42016_n1675), .B(_abc_42016_n3458), .C(_abc_42016_n3503), .D(_abc_42016_n3271), .Y(_abc_42016_n3687) );
  OAI22X1 OAI22X1_8 ( .A(_abc_42016_n796), .B(_abc_42016_n539), .C(_abc_42016_n795), .D(_abc_42016_n565), .Y(_abc_42016_n797) );
  OAI22X1 OAI22X1_80 ( .A(_abc_42016_n2118), .B(_abc_42016_n2255), .C(_abc_42016_n3475), .D(_abc_42016_n3702), .Y(_abc_42016_n3703) );
  OAI22X1 OAI22X1_81 ( .A(_abc_42016_n842), .B(_abc_42016_n1022), .C(_abc_42016_n2376), .D(_abc_42016_n3727), .Y(_abc_42016_n3728) );
  OAI22X1 OAI22X1_82 ( .A(_abc_42016_n3575), .B(_abc_42016_n3769), .C(_abc_42016_n3503), .D(_abc_42016_n3366), .Y(_abc_42016_n3776) );
  OAI22X1 OAI22X1_83 ( .A(_abc_42016_n1151), .B(_abc_42016_n3821), .C(_abc_42016_n3817_1), .D(_abc_42016_n3823), .Y(_abc_42016_n3824) );
  OAI22X1 OAI22X1_84 ( .A(_abc_42016_n709), .B(_abc_42016_n1046), .C(pc_1_), .D(_abc_42016_n4091), .Y(_abc_42016_n4133) );
  OAI22X1 OAI22X1_85 ( .A(_abc_42016_n1848), .B(_abc_42016_n4161), .C(_abc_42016_n2590), .D(_abc_42016_n2423_1), .Y(_abc_42016_n4162) );
  OAI22X1 OAI22X1_86 ( .A(_abc_42016_n1848), .B(_abc_42016_n4187), .C(_abc_42016_n4185), .D(_abc_42016_n2423_1), .Y(_abc_42016_n4188) );
  OAI22X1 OAI22X1_87 ( .A(_abc_42016_n560), .B(_abc_42016_n4213), .C(_abc_42016_n4216), .D(_abc_42016_n4131), .Y(_abc_42016_n4217) );
  OAI22X1 OAI22X1_88 ( .A(_abc_42016_n4091), .B(_abc_42016_n4225), .C(_abc_42016_n4086), .D(_abc_42016_n1393), .Y(_abc_42016_n4226) );
  OAI22X1 OAI22X1_89 ( .A(_abc_42016_n629), .B(_abc_42016_n1046), .C(_abc_42016_n4076), .D(_abc_42016_n1369), .Y(_abc_42016_n4227) );
  OAI22X1 OAI22X1_9 ( .A(_abc_42016_n841), .B(_abc_42016_n845), .C(_abc_42016_n846), .D(_abc_42016_n849), .Y(_abc_42016_n850) );
  OAI22X1 OAI22X1_90 ( .A(_abc_42016_n1848), .B(_abc_42016_n4225), .C(_abc_42016_n2423_1), .D(_abc_42016_n1369), .Y(_abc_42016_n4230) );
  OAI22X1 OAI22X1_91 ( .A(_abc_42016_n722), .B(_abc_42016_n1046), .C(_abc_42016_n4086), .D(_abc_42016_n1425), .Y(_abc_42016_n4236) );
  OAI22X1 OAI22X1_92 ( .A(_abc_42016_n4091), .B(_abc_42016_n4238), .C(_abc_42016_n4076), .D(_abc_42016_n1436), .Y(_abc_42016_n4239) );
  OAI22X1 OAI22X1_93 ( .A(_abc_42016_n1848), .B(_abc_42016_n4238), .C(_abc_42016_n2423_1), .D(_abc_42016_n1436), .Y(_abc_42016_n4243) );
  OAI22X1 OAI22X1_94 ( .A(_abc_42016_n1485), .B(_abc_42016_n2423_1), .C(_abc_42016_n1848), .D(_abc_42016_n4263), .Y(_abc_42016_n4269) );
  OAI22X1 OAI22X1_95 ( .A(_abc_42016_n1504), .B(_abc_42016_n4076), .C(_abc_42016_n4091), .D(_abc_42016_n4276), .Y(_abc_42016_n4277) );
  OAI22X1 OAI22X1_96 ( .A(_abc_42016_n1504), .B(_abc_42016_n2423_1), .C(_abc_42016_n1848), .D(_abc_42016_n4276), .Y(_abc_42016_n4281) );
  OAI22X1 OAI22X1_97 ( .A(_abc_42016_n1545), .B(_abc_42016_n2423_1), .C(_abc_42016_n1848), .D(_abc_42016_n4288), .Y(_abc_42016_n4289) );
  OAI22X1 OAI22X1_98 ( .A(_abc_42016_n1545), .B(_abc_42016_n4076), .C(_abc_42016_n4091), .D(_abc_42016_n4288), .Y(_abc_42016_n4292) );
  OAI22X1 OAI22X1_99 ( .A(_abc_42016_n1564), .B(_abc_42016_n4158), .C(_abc_42016_n4305), .D(_abc_42016_n4307), .Y(_abc_42016_n4308) );
  OR2X2 OR2X2_1 ( .A(_abc_42016_n647), .B(_abc_42016_n643_1), .Y(_abc_42016_n648_1) );
  OR2X2 OR2X2_10 ( .A(_abc_42016_n1112), .B(_abc_42016_n1098), .Y(_abc_42016_n1113_1) );
  OR2X2 OR2X2_11 ( .A(_abc_42016_n1115), .B(_abc_42016_n1114_1), .Y(_abc_42016_n1116) );
  OR2X2 OR2X2_12 ( .A(_abc_42016_n1120), .B(_abc_42016_n1139), .Y(_abc_42016_n1140) );
  OR2X2 OR2X2_13 ( .A(_abc_42016_n1167), .B(_abc_42016_n1164), .Y(_abc_42016_n1168) );
  OR2X2 OR2X2_14 ( .A(_abc_42016_n1140), .B(_abc_42016_n843), .Y(_abc_42016_n1188) );
  OR2X2 OR2X2_15 ( .A(_abc_42016_n1202), .B(_abc_42016_n1203), .Y(_abc_42016_n1205) );
  OR2X2 OR2X2_16 ( .A(_abc_42016_n1267), .B(_abc_42016_n1265), .Y(_abc_42016_n1268) );
  OR2X2 OR2X2_17 ( .A(_abc_42016_n1271_1), .B(_abc_42016_n1270), .Y(_abc_42016_n1272_1) );
  OR2X2 OR2X2_18 ( .A(_abc_42016_n1324), .B(_abc_42016_n1330), .Y(_abc_42016_n1331_1) );
  OR2X2 OR2X2_19 ( .A(_abc_42016_n1433), .B(_abc_42016_n1440), .Y(_abc_42016_n1441) );
  OR2X2 OR2X2_2 ( .A(_abc_42016_n648_1), .B(_abc_42016_n610), .Y(_abc_42016_n649_1) );
  OR2X2 OR2X2_20 ( .A(_abc_42016_n1519), .B(_abc_42016_n1518), .Y(_abc_42016_n1520) );
  OR2X2 OR2X2_21 ( .A(_abc_42016_n1540), .B(_abc_42016_n1410_1), .Y(_abc_42016_n1541) );
  OR2X2 OR2X2_22 ( .A(_abc_42016_n1637), .B(_abc_42016_n1641), .Y(_abc_42016_n1642) );
  OR2X2 OR2X2_23 ( .A(_abc_42016_n2569), .B(_abc_42016_n2563), .Y(_abc_42016_n2570) );
  OR2X2 OR2X2_24 ( .A(_abc_42016_n2681), .B(_abc_42016_n2679), .Y(_abc_42016_n2682) );
  OR2X2 OR2X2_25 ( .A(_abc_42016_n2713), .B(_abc_42016_n2708), .Y(_abc_42016_n2714) );
  OR2X2 OR2X2_26 ( .A(_abc_42016_n2735), .B(_abc_42016_n2831), .Y(_abc_42016_n2832) );
  OR2X2 OR2X2_27 ( .A(_abc_42016_n2864), .B(_abc_42016_n2735), .Y(_abc_42016_n2865) );
  OR2X2 OR2X2_28 ( .A(_abc_42016_n3629), .B(_abc_42016_n2758), .Y(_abc_42016_n3630) );
  OR2X2 OR2X2_29 ( .A(_abc_42016_n3638), .B(_abc_42016_n3641), .Y(_abc_42016_n3642) );
  OR2X2 OR2X2_3 ( .A(_abc_42016_n651_1), .B(_abc_42016_n641), .Y(_abc_42016_n653) );
  OR2X2 OR2X2_30 ( .A(_abc_42016_n3619), .B(_abc_42016_n2113), .Y(_abc_42016_n3722) );
  OR2X2 OR2X2_31 ( .A(_abc_42016_n4079), .B(_abc_42016_n4081), .Y(_abc_42016_n4082) );
  OR2X2 OR2X2_32 ( .A(_abc_42016_n4692), .B(_abc_42016_n4630), .Y(_abc_42016_n4708) );
  OR2X2 OR2X2_33 ( .A(alu__abc_41682_n123), .B(alu_oprb_1_), .Y(alu__abc_41682_n124_1) );
  OR2X2 OR2X2_34 ( .A(alu_oprb_1_), .B(alu_opra_1_), .Y(alu__abc_41682_n140) );
  OR2X2 OR2X2_35 ( .A(alu__abc_41682_n70), .B(alu__abc_41682_n62), .Y(alu__abc_41682_n228) );
  OR2X2 OR2X2_36 ( .A(alu__abc_41682_n41), .B(alu__abc_41682_n44), .Y(alu__abc_41682_n233) );
  OR2X2 OR2X2_37 ( .A(alu__abc_41682_n103), .B(alu__abc_41682_n198), .Y(alu__abc_41682_n365) );
  OR2X2 OR2X2_4 ( .A(_abc_42016_n736), .B(_abc_42016_n718), .Y(_abc_42016_n737) );
  OR2X2 OR2X2_5 ( .A(_abc_42016_n942), .B(_abc_42016_n943), .Y(_abc_42016_n944) );
  OR2X2 OR2X2_6 ( .A(_abc_42016_n914), .B(regfil_0__7_), .Y(_abc_42016_n950) );
  OR2X2 OR2X2_7 ( .A(_abc_42016_n588_1), .B(_abc_42016_n968), .Y(_abc_42016_n969) );
  OR2X2 OR2X2_8 ( .A(_abc_42016_n970), .B(_abc_42016_n951), .Y(_abc_42016_n971) );
  OR2X2 OR2X2_9 ( .A(_abc_42016_n1108), .B(_abc_42016_n1107_1), .Y(_abc_42016_n1110_1) );
  XNOR2X1 XNOR2X1_1 ( .A(_abc_42016_n863), .B(_abc_42016_n874), .Y(_abc_42016_n875) );
  XNOR2X1 XNOR2X1_10 ( .A(_abc_42016_n1570), .B(_abc_42016_n1584_1), .Y(_abc_42016_n1589) );
  XNOR2X1 XNOR2X1_11 ( .A(_abc_42016_n615), .B(regfil_1__5_), .Y(_abc_42016_n1744) );
  XNOR2X1 XNOR2X1_12 ( .A(_abc_42016_n3362), .B(_abc_42016_n2101), .Y(_abc_42016_n3389) );
  XNOR2X1 XNOR2X1_13 ( .A(_abc_42016_n3381), .B(_abc_42016_n3388), .Y(_abc_42016_n3404) );
  XNOR2X1 XNOR2X1_14 ( .A(_abc_42016_n3762), .B(sp_15_), .Y(_abc_42016_n3789) );
  XNOR2X1 XNOR2X1_15 ( .A(_abc_42016_n3915), .B(_abc_42016_n3916), .Y(_abc_42016_n3917) );
  XNOR2X1 XNOR2X1_16 ( .A(_abc_42016_n3961), .B(_abc_42016_n3962), .Y(_abc_42016_n3963) );
  XNOR2X1 XNOR2X1_17 ( .A(_abc_42016_n3971), .B(_abc_42016_n3972), .Y(_abc_42016_n3973) );
  XNOR2X1 XNOR2X1_18 ( .A(_abc_42016_n1385), .B(pc_4_), .Y(_abc_42016_n4173) );
  XNOR2X1 XNOR2X1_19 ( .A(_abc_42016_n1544), .B(pc_14_), .Y(_abc_42016_n4301) );
  XNOR2X1 XNOR2X1_2 ( .A(_abc_42016_n1076), .B(_abc_42016_n1029), .Y(_abc_42016_n1077) );
  XNOR2X1 XNOR2X1_20 ( .A(opcode_3_), .B(parity), .Y(_abc_42016_n4642) );
  XNOR2X1 XNOR2X1_21 ( .A(alu_oprb_2_), .B(alu_opra_2_), .Y(alu__abc_41682_n137) );
  XNOR2X1 XNOR2X1_22 ( .A(alu__abc_41682_n36), .B(alu__abc_41682_n37), .Y(alu__abc_41682_n291) );
  XNOR2X1 XNOR2X1_23 ( .A(alu__abc_41682_n303), .B(alu__abc_41682_n311), .Y(alu__abc_41682_n316) );
  XNOR2X1 XNOR2X1_3 ( .A(_abc_42016_n1126), .B(_abc_42016_n1139), .Y(_abc_42016_n1172_1) );
  XNOR2X1 XNOR2X1_4 ( .A(regfil_5__5_), .B(sp_5_), .Y(_abc_42016_n1231) );
  XNOR2X1 XNOR2X1_5 ( .A(regfil_1__5_), .B(regfil_5__5_), .Y(_abc_42016_n1236) );
  XNOR2X1 XNOR2X1_6 ( .A(regfil_3__5_), .B(regfil_5__5_), .Y(_abc_42016_n1243) );
  XNOR2X1 XNOR2X1_7 ( .A(_abc_42016_n1315), .B(_abc_42016_n1318), .Y(_abc_42016_n1319) );
  XNOR2X1 XNOR2X1_8 ( .A(_abc_42016_n1484), .B(_abc_42016_n1503), .Y(_abc_42016_n1504) );
  XNOR2X1 XNOR2X1_9 ( .A(_abc_42016_n1585), .B(_abc_42016_n1584_1), .Y(_abc_42016_n1586_1) );
  XOR2X1 XOR2X1_1 ( .A(regfil_1__2_), .B(regfil_5__2_), .Y(_abc_42016_n1108) );
  XOR2X1 XOR2X1_10 ( .A(regfil_2__6_), .B(regfil_4__6_), .Y(_abc_42016_n2149) );
  XOR2X1 XOR2X1_11 ( .A(regfil_2__4_), .B(regfil_4__4_), .Y(_abc_42016_n2154) );
  XOR2X1 XOR2X1_12 ( .A(regfil_2__0_), .B(regfil_4__0_), .Y(_abc_42016_n2167) );
  XOR2X1 XOR2X1_13 ( .A(regfil_0__4_), .B(regfil_4__4_), .Y(_abc_42016_n2187) );
  XOR2X1 XOR2X1_14 ( .A(sp_0_), .B(sp_1_), .Y(_abc_42016_n3476_1) );
  XOR2X1 XOR2X1_15 ( .A(_abc_42016_n3846), .B(_abc_42016_n3847), .Y(_abc_42016_n3848) );
  XOR2X1 XOR2X1_16 ( .A(alu_oprb_2_), .B(alu_opra_2_), .Y(alu__abc_41682_n41) );
  XOR2X1 XOR2X1_17 ( .A(alu__abc_41682_n303), .B(alu__abc_41682_n311), .Y(alu__abc_41682_n312) );
  XOR2X1 XOR2X1_2 ( .A(regfil_5__2_), .B(sp_2_), .Y(_abc_42016_n1115) );
  XOR2X1 XOR2X1_3 ( .A(_abc_42016_n1152), .B(_abc_42016_n1155), .Y(_abc_42016_n1156) );
  XOR2X1 XOR2X1_4 ( .A(regfil_3__4_), .B(regfil_5__4_), .Y(_abc_42016_n1203) );
  XOR2X1 XOR2X1_5 ( .A(_abc_42016_n1215), .B(_abc_42016_n1212), .Y(_abc_42016_n1216) );
  XOR2X1 XOR2X1_6 ( .A(_abc_42016_n1242), .B(_abc_42016_n1243), .Y(_abc_42016_n1244) );
  XOR2X1 XOR2X1_7 ( .A(regfil_1__6_), .B(regfil_5__6_), .Y(_abc_42016_n1265) );
  XOR2X1 XOR2X1_8 ( .A(regfil_3__6_), .B(regfil_5__6_), .Y(_abc_42016_n1273) );
  XOR2X1 XOR2X1_9 ( .A(regfil_5__6_), .B(sp_6_), .Y(_abc_42016_n1281) );
endmodule
